/******** Key Information: *********** 
Key 1:   bin: '1100110000000110011101110000100001000111100011100'    dec: 448656277802780
Key 2:   bin: '1100000010000101001001101001011011011000101001110'    dec: 423356221206862
Key 3:   bin: '1111001101000011111000001111001110110010110011010'    dec: 534945724851610
Key 4:   bin: '0010100101001110100110111100101110110010101101011'    dec: 90835196011883
Key 5:   bin: '0000101011011100100011010010100010000011011011011'    dec: 23884754650843
Key 6:   bin: '0111011011111010111001111001111010100110011111011'    dec: 261639999671547
Key 7:   bin: '1000111101000100000100011111110011000100001110001'    dec: 315045044652145
Key 8:   bin: '0100010010111001100111111000101110000100010000001'    dec: 151128072718465
Key 9:   bin: '1000001000111100110011101110111010111101101101110'    dec: 286395362802542
Key 10:   bin: '0100001100111110100011000001011000100001100011110'    dec: 147871834587934
Key 11:   bin: '1111101000100110111101001110010001110100000100111'    dec: 550090448627751
Key 12:   bin: '0011101010101110111100101010000111100101001101111'    dec: 129046138833519
Key 13:   bin: '0100000110100110110011001110111110001010100010110'    dec: 144369317254422
Key 14:   bin: '0011011001011010011011000101011000001100110001000'    dec: 119523985070472
Key 15:   bin: '1010101001011001111110101111111111110101010100001'    dec: 374606879779489
Key 16:   bin: '1111011010000001010011010101100000110110101100000'    dec: 542070417681760
**************************************/

module cow (keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, clk,rst,
	x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
	x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
	x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45,
	x46, x47, x48, x49, 
	y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24);

input clk, rst, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
	x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
	x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45,
	x46, x47, x48, x49;
input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48;
output y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24;
reg[9:0] counter = 0;
reg y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24;

parameter s1=1, s2=2, s3=3, s4=4, s5=5, s6=6, s7=7, s8=8, s9=9, s10=10,
	s11=11, s12=12, s13=13, s14=14, s15=15, s16=16, s17=17, s18=18, s19=19, s20=20,
	s21=21, s22=22, s23=23, s24=24;
integer pr_state;
integer nx_state;

always @(negedge clk or posedge rst)
begin
	if (rst == 1'b1)
		counter <= 0;
	else
		counter <= (counter >= 319) ? 0 : counter + 1;
end

always@(  negedge clk or posedge rst )
begin
	if (rst == 1'b1)
	 begin
		pr_state = s1;
	end
	else
	begin
		if ( counter <= 19 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b1 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b1 && keyinput5 == 1'b1 && keyinput6 == 1'b0 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b0 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b1 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b0 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b1 && keyinput20 == 1'b0 && keyinput21 == 1'b1 && keyinput22 == 1'b1 && keyinput23 == 1'b1 && keyinput24 == 1'b0 && keyinput25 == 1'b0 && keyinput26 == 1'b0 && keyinput27 == 1'b0 && keyinput28 == 1'b1 && keyinput29 == 1'b0 && keyinput30 == 1'b0 && keyinput31 == 1'b0 && keyinput32 == 1'b0 && keyinput33 == 1'b1 && keyinput34 == 1'b0 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b1 && keyinput39 == 1'b1 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b0 && keyinput43 == 1'b0 && keyinput44 == 1'b1 && keyinput45 == 1'b1 && keyinput46 == 1'b1 && keyinput47 == 1'b0 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s12;
		end
		if ( counter > 19 && counter <= 39 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b1 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b0 && keyinput5 == 1'b0 && keyinput6 == 1'b0 && keyinput7 == 1'b0 && keyinput8 == 1'b1 && keyinput9 == 1'b0 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b1 && keyinput14 == 1'b0 && keyinput15 == 1'b1 && keyinput16 == 1'b0 && keyinput17 == 1'b0 && keyinput18 == 1'b1 && keyinput19 == 1'b0 && keyinput20 == 1'b0 && keyinput21 == 1'b1 && keyinput22 == 1'b1 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b0 && keyinput26 == 1'b0 && keyinput27 == 1'b1 && keyinput28 == 1'b0 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b0 && keyinput32 == 1'b1 && keyinput33 == 1'b1 && keyinput34 == 1'b0 && keyinput35 == 1'b1 && keyinput36 == 1'b1 && keyinput37 == 1'b0 && keyinput38 == 1'b0 && keyinput39 == 1'b0 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b1 && keyinput43 == 1'b0 && keyinput44 == 1'b0 && keyinput45 == 1'b1 && keyinput46 == 1'b1 && keyinput47 == 1'b1 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s4;
		end
		if ( counter > 39 && counter <= 59 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b1 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b0 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b1 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b0 && keyinput14 == 1'b1 && keyinput15 == 1'b1 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b0 && keyinput20 == 1'b0 && keyinput21 == 1'b0 && keyinput22 == 1'b0 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b1 && keyinput27 == 1'b1 && keyinput28 == 1'b0 && keyinput29 == 1'b0 && keyinput30 == 1'b1 && keyinput31 == 1'b1 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b1 && keyinput35 == 1'b1 && keyinput36 == 1'b0 && keyinput37 == 1'b0 && keyinput38 == 1'b1 && keyinput39 == 1'b0 && keyinput40 == 1'b1 && keyinput41 == 1'b1 && keyinput42 == 1'b0 && keyinput43 == 1'b0 && keyinput44 == 1'b1 && keyinput45 == 1'b1 && keyinput46 == 1'b0 && keyinput47 == 1'b1 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s20;
		end
		if ( counter > 59 && counter <= 79 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b0 && keyinput2 == 1'b1 && keyinput3 == 1'b0 && keyinput4 == 1'b1 && keyinput5 == 1'b0 && keyinput6 == 1'b0 && keyinput7 == 1'b1 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b1 && keyinput13 == 1'b1 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b0 && keyinput18 == 1'b0 && keyinput19 == 1'b1 && keyinput20 == 1'b1 && keyinput21 == 1'b0 && keyinput22 == 1'b1 && keyinput23 == 1'b1 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b0 && keyinput27 == 1'b0 && keyinput28 == 1'b1 && keyinput29 == 1'b0 && keyinput30 == 1'b1 && keyinput31 == 1'b1 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b1 && keyinput35 == 1'b1 && keyinput36 == 1'b0 && keyinput37 == 1'b0 && keyinput38 == 1'b1 && keyinput39 == 1'b0 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b1 && keyinput43 == 1'b1 && keyinput44 == 1'b0 && keyinput45 == 1'b1 && keyinput46 == 1'b0 && keyinput47 == 1'b1 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s19;
		end
		if ( counter > 79 && counter <= 99 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b0 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b1 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b1 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b1 && keyinput14 == 1'b0 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b0 && keyinput18 == 1'b0 && keyinput19 == 1'b0 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b0 && keyinput23 == 1'b1 && keyinput24 == 1'b0 && keyinput25 == 1'b0 && keyinput26 == 1'b1 && keyinput27 == 1'b0 && keyinput28 == 1'b1 && keyinput29 == 1'b0 && keyinput30 == 1'b0 && keyinput31 == 1'b0 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b0 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b0 && keyinput38 == 1'b1 && keyinput39 == 1'b1 && keyinput40 == 1'b0 && keyinput41 == 1'b1 && keyinput42 == 1'b1 && keyinput43 == 1'b0 && keyinput44 == 1'b1 && keyinput45 == 1'b1 && keyinput46 == 1'b0 && keyinput47 == 1'b1 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s14;
		end
		if ( counter > 99 && counter <= 119 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b1 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b0 && keyinput5 == 1'b1 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b1 && keyinput9 == 1'b1 && keyinput10 == 1'b1 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b0 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b0 && keyinput20 == 1'b0 && keyinput21 == 1'b1 && keyinput22 == 1'b1 && keyinput23 == 1'b1 && keyinput24 == 1'b1 && keyinput25 == 1'b0 && keyinput26 == 1'b0 && keyinput27 == 1'b1 && keyinput28 == 1'b1 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b0 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b1 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b1 && keyinput39 == 1'b0 && keyinput40 == 1'b0 && keyinput41 == 1'b1 && keyinput42 == 1'b1 && keyinput43 == 1'b1 && keyinput44 == 1'b1 && keyinput45 == 1'b1 && keyinput46 == 1'b0 && keyinput47 == 1'b1 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s1;
		end
		if ( counter > 119 && counter <= 139 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b0 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b1 && keyinput5 == 1'b1 && keyinput6 == 1'b1 && keyinput7 == 1'b1 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b1 && keyinput14 == 1'b0 && keyinput15 == 1'b0 && keyinput16 == 1'b0 && keyinput17 == 1'b0 && keyinput18 == 1'b0 && keyinput19 == 1'b1 && keyinput20 == 1'b0 && keyinput21 == 1'b0 && keyinput22 == 1'b0 && keyinput23 == 1'b1 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b1 && keyinput27 == 1'b1 && keyinput28 == 1'b1 && keyinput29 == 1'b1 && keyinput30 == 1'b0 && keyinput31 == 1'b0 && keyinput32 == 1'b1 && keyinput33 == 1'b1 && keyinput34 == 1'b0 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b0 && keyinput40 == 1'b0 && keyinput41 == 1'b0 && keyinput42 == 1'b1 && keyinput43 == 1'b1 && keyinput44 == 1'b1 && keyinput45 == 1'b0 && keyinput46 == 1'b0 && keyinput47 == 1'b0 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s10;
		end
		if ( counter > 139 && counter <= 159 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b1 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b0 && keyinput5 == 1'b1 && keyinput6 == 1'b0 && keyinput7 == 1'b0 && keyinput8 == 1'b1 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b0 && keyinput14 == 1'b0 && keyinput15 == 1'b1 && keyinput16 == 1'b1 && keyinput17 == 1'b0 && keyinput18 == 1'b0 && keyinput19 == 1'b1 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b1 && keyinput23 == 1'b1 && keyinput24 == 1'b1 && keyinput25 == 1'b0 && keyinput26 == 1'b0 && keyinput27 == 1'b0 && keyinput28 == 1'b1 && keyinput29 == 1'b0 && keyinput30 == 1'b1 && keyinput31 == 1'b1 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b0 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b0 && keyinput40 == 1'b0 && keyinput41 == 1'b1 && keyinput42 == 1'b0 && keyinput43 == 1'b0 && keyinput44 == 1'b0 && keyinput45 == 1'b0 && keyinput46 == 1'b0 && keyinput47 == 1'b0 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s17;
		end
		if ( counter > 159 && counter <= 179 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b0 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b0 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b1 && keyinput14 == 1'b0 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b0 && keyinput19 == 1'b0 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b1 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b1 && keyinput27 == 1'b0 && keyinput28 == 1'b1 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b0 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b1 && keyinput35 == 1'b1 && keyinput36 == 1'b1 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b1 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b1 && keyinput43 == 1'b1 && keyinput44 == 1'b0 && keyinput45 == 1'b1 && keyinput46 == 1'b1 && keyinput47 == 1'b1 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s8;
		end
		if ( counter > 179 && counter <= 199 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b1 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b0 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b1 && keyinput8 == 1'b0 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b1 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b0 && keyinput18 == 1'b0 && keyinput19 == 1'b0 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b0 && keyinput23 == 1'b0 && keyinput24 == 1'b0 && keyinput25 == 1'b0 && keyinput26 == 1'b0 && keyinput27 == 1'b1 && keyinput28 == 1'b0 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b0 && keyinput32 == 1'b0 && keyinput33 == 1'b0 && keyinput34 == 1'b1 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b0 && keyinput38 == 1'b0 && keyinput39 == 1'b1 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b0 && keyinput43 == 1'b0 && keyinput44 == 1'b1 && keyinput45 == 1'b1 && keyinput46 == 1'b1 && keyinput47 == 1'b1 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s16;
		end
		if ( counter > 199 && counter <= 219 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b1 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b1 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b1 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b1 && keyinput20 == 1'b0 && keyinput21 == 1'b1 && keyinput22 == 1'b0 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b1 && keyinput27 == 1'b0 && keyinput28 == 1'b0 && keyinput29 == 1'b1 && keyinput30 == 1'b0 && keyinput31 == 1'b0 && keyinput32 == 1'b0 && keyinput33 == 1'b1 && keyinput34 == 1'b1 && keyinput35 == 1'b1 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b0 && keyinput40 == 1'b0 && keyinput41 == 1'b0 && keyinput42 == 1'b0 && keyinput43 == 1'b1 && keyinput44 == 1'b0 && keyinput45 == 1'b0 && keyinput46 == 1'b1 && keyinput47 == 1'b1 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s22;
		end
		if ( counter > 219 && counter <= 239 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b0 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b1 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b1 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b0 && keyinput12 == 1'b1 && keyinput13 == 1'b1 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b1 && keyinput20 == 1'b0 && keyinput21 == 1'b0 && keyinput22 == 1'b1 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b0 && keyinput26 == 1'b1 && keyinput27 == 1'b0 && keyinput28 == 1'b0 && keyinput29 == 1'b0 && keyinput30 == 1'b0 && keyinput31 == 1'b1 && keyinput32 == 1'b1 && keyinput33 == 1'b1 && keyinput34 == 1'b1 && keyinput35 == 1'b0 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b1 && keyinput40 == 1'b0 && keyinput41 == 1'b0 && keyinput42 == 1'b1 && keyinput43 == 1'b1 && keyinput44 == 1'b0 && keyinput45 == 1'b1 && keyinput46 == 1'b1 && keyinput47 == 1'b1 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s2;
		end
		if ( counter > 239 && counter <= 259 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b1 && keyinput2 == 1'b0 && keyinput3 == 1'b0 && keyinput4 == 1'b0 && keyinput5 == 1'b0 && keyinput6 == 1'b0 && keyinput7 == 1'b1 && keyinput8 == 1'b1 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b1 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b0 && keyinput19 == 1'b0 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b0 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b1 && keyinput27 == 1'b0 && keyinput28 == 1'b1 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b1 && keyinput32 == 1'b1 && keyinput33 == 1'b0 && keyinput34 == 1'b0 && keyinput35 == 1'b0 && keyinput36 == 1'b1 && keyinput37 == 1'b0 && keyinput38 == 1'b1 && keyinput39 == 1'b0 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b0 && keyinput43 == 1'b0 && keyinput44 == 1'b1 && keyinput45 == 1'b0 && keyinput46 == 1'b1 && keyinput47 == 1'b1 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s13;
		end
		if ( counter > 259 && counter <= 279 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b0 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b0 && keyinput5 == 1'b1 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b0 && keyinput14 == 1'b1 && keyinput15 == 1'b0 && keyinput16 == 1'b0 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b0 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b0 && keyinput23 == 1'b0 && keyinput24 == 1'b0 && keyinput25 == 1'b1 && keyinput26 == 1'b0 && keyinput27 == 1'b1 && keyinput28 == 1'b0 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b0 && keyinput32 == 1'b0 && keyinput33 == 1'b0 && keyinput34 == 1'b0 && keyinput35 == 1'b0 && keyinput36 == 1'b1 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b0 && keyinput40 == 1'b1 && keyinput41 == 1'b1 && keyinput42 == 1'b0 && keyinput43 == 1'b0 && keyinput44 == 1'b0 && keyinput45 == 1'b1 && keyinput46 == 1'b0 && keyinput47 == 1'b0 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s15;
		end
		if ( counter > 279 && counter <= 299 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b0 && keyinput2 == 1'b1 && keyinput3 == 1'b0 && keyinput4 == 1'b1 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b1 && keyinput12 == 1'b1 && keyinput13 == 1'b0 && keyinput14 == 1'b0 && keyinput15 == 1'b1 && keyinput16 == 1'b1 && keyinput17 == 1'b1 && keyinput18 == 1'b1 && keyinput19 == 1'b1 && keyinput20 == 1'b1 && keyinput21 == 1'b0 && keyinput22 == 1'b1 && keyinput23 == 1'b0 && keyinput24 == 1'b1 && keyinput25 == 1'b1 && keyinput26 == 1'b1 && keyinput27 == 1'b1 && keyinput28 == 1'b1 && keyinput29 == 1'b1 && keyinput30 == 1'b1 && keyinput31 == 1'b1 && keyinput32 == 1'b1 && keyinput33 == 1'b1 && keyinput34 == 1'b1 && keyinput35 == 1'b1 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b0 && keyinput39 == 1'b1 && keyinput40 == 1'b0 && keyinput41 == 1'b1 && keyinput42 == 1'b0 && keyinput43 == 1'b1 && keyinput44 == 1'b0 && keyinput45 == 1'b0 && keyinput46 == 1'b0 && keyinput47 == 1'b0 && keyinput48 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s9;
		end
		if ( counter > 299 && counter <= 319 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b1 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b0 && keyinput5 == 1'b1 && keyinput6 == 1'b1 && keyinput7 == 1'b0 && keyinput8 == 1'b1 && keyinput9 == 1'b0 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b0 && keyinput14 == 1'b0 && keyinput15 == 1'b1 && keyinput16 == 1'b0 && keyinput17 == 1'b1 && keyinput18 == 1'b0 && keyinput19 == 1'b0 && keyinput20 == 1'b1 && keyinput21 == 1'b1 && keyinput22 == 1'b0 && keyinput23 == 1'b1 && keyinput24 == 1'b0 && keyinput25 == 1'b1 && keyinput26 == 1'b0 && keyinput27 == 1'b1 && keyinput28 == 1'b1 && keyinput29 == 1'b0 && keyinput30 == 1'b0 && keyinput31 == 1'b0 && keyinput32 == 1'b0 && keyinput33 == 1'b0 && keyinput34 == 1'b1 && keyinput35 == 1'b1 && keyinput36 == 1'b0 && keyinput37 == 1'b1 && keyinput38 == 1'b1 && keyinput39 == 1'b0 && keyinput40 == 1'b1 && keyinput41 == 1'b0 && keyinput42 == 1'b1 && keyinput43 == 1'b1 && keyinput44 == 1'b0 && keyinput45 == 1'b0 && keyinput46 == 1'b0 && keyinput47 == 1'b0 && keyinput48 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s3;
		end
	end
end


always@ ( pr_state or x1 or x2 or x3 or x4 or x5 or x6 or x7 or x8 or x9 or x10 or x11 or x12 or x13 or x14 or x15 or 
	x16 or x17 or x18 or x19 or x20 or x21 or x22 or x23 or x24 or x25 or x26 or x27 or x28 or x29 or x30 or 
	x31 or x32 or x33 or x34 or x35 or x36 or x37 or x38 or x39 or x40 or x41 or x42 or x43 or x44 or x45 or 
	x46 or x47 or x48 or x49)
	begin
			y1 = 1'b0;	y2 = 1'b0;	y3 = 1'b0;	y4 = 1'b0;	
			y5 = 1'b0;	y6 = 1'b0;	y7 = 1'b0;	y8 = 1'b0;	
			y9 = 1'b0;	y10 = 1'b0;	y11 = 1'b0;	y12 = 1'b0;	
			y13 = 1'b0;	y14 = 1'b0;	y15 = 1'b0;	y16 = 1'b0;	
			y17 = 1'b0;	y18 = 1'b0;	y19 = 1'b0;	y20 = 1'b0;	
			y21 = 1'b0;	y22 = 1'b0;	y23 = 1'b0;	y24 = 1'b0;	
		case ( pr_state )
				s1 : if( x15 && x10 && x12 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s2;
						end
					else if( x15 && x10 && x12 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( x15 && x10 && x12 && ~x23 && ~x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && x10 && ~x12 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s5;
						end
					else if( x15 && ~x10 && x1 && x22 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s6;
						end
					else if( x15 && ~x10 && x1 && ~x22 && x2 && x3 && x11 )
						nx_state = s1;
					else if( x15 && ~x10 && x1 && ~x22 && x2 && x3 && ~x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x15 && ~x10 && x1 && ~x22 && x2 && ~x3 && x11 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && ~x10 && x1 && ~x22 && x2 && ~x3 && x11 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( x15 && ~x10 && x1 && ~x22 && x2 && ~x3 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( x15 && ~x10 && x1 && ~x22 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && ~x10 && ~x1 && x11 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && ~x10 && ~x1 && x11 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x15 && ~x10 && ~x1 && ~x11 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x10 && x39 && x36 )
						nx_state = s1;
					else if( ~x15 && x10 && x39 && ~x36 && x46 && x48 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && x10 && x39 && ~x36 && x46 && ~x48 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x15 && x10 && x39 && ~x36 && ~x46 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && x10 && ~x39 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x15 && ~x10 && x11 && x34 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x15 && ~x10 && x11 && x34 && ~x8 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && ~x10 && x11 && x34 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x10 && x11 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x15 && ~x10 && x11 && ~x34 && x32 && ~x7 && x43 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && ~x10 && x11 && ~x34 && x32 && ~x7 && x43 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x10 && x11 && ~x34 && x32 && ~x7 && ~x43 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && ~x10 && x11 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x15 && ~x10 && ~x11 && x12 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && ~x10 && ~x11 && x12 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && ~x10 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && ~x10 && ~x11 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x15 && ~x10 && ~x11 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x10 && ~x11 && ~x12 && x13 && x1 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x10 && ~x11 && ~x12 && x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && ~x10 && ~x11 && ~x12 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s1;
				s2 : if( x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s2;
				s3 : if( x15 && x19 && x28 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s16;
						end
					else if( x15 && x19 && x28 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x19 && x28 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( x15 && x19 && ~x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x15 && ~x19 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x15 && x13 && x23 && x48 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && x13 && x23 && ~x48 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x15 && x13 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && ~x13 && x28 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && ~x13 && x28 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x13 && x28 && ~x35 && x21 )
						nx_state = s1;
					else if( ~x15 && ~x13 && x28 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x13 && ~x28 && x6 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x15 && ~x13 && ~x28 && x6 && ~x35 && x21 )
						nx_state = s1;
					else if( ~x15 && ~x13 && ~x28 && x6 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else nx_state = s3;
				s4 : if( x15 && x30 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s18;
						end
					else if( x15 && x30 && x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s14;
						end
					else if( x15 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( x15 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( x15 && x30 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s16;
						end
					else if( x15 && x30 && x16 && ~x6 && ~x8 )
						nx_state = s1;
					else if( x15 && x30 && ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x30 && ~x16 && ~x10 )
						nx_state = s1;
					else if( x15 && ~x30 && x5 && x9 )
						nx_state = s1;
					else if( x15 && ~x30 && x5 && ~x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && ~x30 && ~x5 && x3 && x11 )
						nx_state = s4;
					else if( x15 && ~x30 && ~x5 && x3 && ~x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x15 && ~x30 && ~x5 && ~x3 && x11 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( x15 && ~x30 && ~x5 && ~x3 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && x48 && x24 && x5 && x36 )
						nx_state = s4;
					else if( ~x15 && x48 && x24 && x5 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && x48 && x24 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && x48 && ~x24 && x31 && x29 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && x48 && ~x24 && x31 && ~x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && x48 && ~x24 && ~x31 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && ~x48 && x11 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x15 && ~x48 && x11 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x48 && x11 && ~x35 && x21 )
						nx_state = s1;
					else if( ~x15 && ~x48 && x11 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x48 && ~x11 && x45 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x15 && ~x48 && ~x11 && x45 && ~x35 && x21 )
						nx_state = s1;
					else if( ~x15 && ~x48 && ~x11 && x45 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x48 && ~x11 && ~x45 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x15 && ~x48 && ~x11 && ~x45 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && ~x48 && ~x11 && ~x45 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else nx_state = s4;
				s5 : if( x15 && x12 && x27 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( x15 && x12 && x27 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && x12 && x27 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x12 && ~x27 && x1 && x29 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x15 && x12 && ~x27 && x1 && ~x29 )
						nx_state = s5;
					else if( x15 && x12 && ~x27 && ~x1 )
						nx_state = s5;
					else if( x15 && ~x12 && x29 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s14;
						end
					else if( x15 && ~x12 && ~x29 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x15 && x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x15 && ~x17 && x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x15 && ~x17 && ~x41 )
						nx_state = s5;
					else nx_state = s5;
				s6 : if( x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else nx_state = s6;
				s7 : if( x15 && x14 && x8 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x14 && x8 && ~x10 )
						nx_state = s1;
					else if( x15 && x14 && ~x8 && x30 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x15 && x14 && ~x8 && x30 && ~x1 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( x15 && x14 && ~x8 && x30 && ~x1 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( x15 && x14 && ~x8 && ~x30 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && ~x14 && x3 && x32 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( x15 && ~x14 && x3 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && ~x14 && ~x3 )
						nx_state = s7;
					else if( ~x15 && x16 && x43 && x27 && x29 && x40 )
						begin
							y13 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x15 && x16 && x43 && x27 && x29 && ~x40 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x16 && x43 && x27 && ~x29 && x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x16 && x43 && x27 && ~x29 && ~x33 && x41 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x15 && x16 && x43 && x27 && ~x29 && ~x33 && ~x41 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x16 && x43 && ~x27 )
						nx_state = s7;
					else if( ~x15 && x16 && ~x43 )
						nx_state = s1;
					else if( ~x15 && ~x16 && x37 && x42 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && ~x16 && x37 && x42 && ~x1 )
						nx_state = s7;
					else if( ~x15 && ~x16 && x37 && ~x42 )
						nx_state = s1;
					else if( ~x15 && ~x16 && ~x37 && x25 )
						nx_state = s1;
					else if( ~x15 && ~x16 && ~x37 && ~x25 && x4 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x15 && ~x16 && ~x37 && ~x25 && x4 && ~x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && ~x16 && ~x37 && ~x25 && ~x4 )
						nx_state = s7;
					else nx_state = s7;
				s8 : if( x15 && x24 && x26 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( x15 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s24;
						end
					else if( x15 && x24 && ~x26 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( x15 && ~x24 && x28 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s5;
						end
					else if( x15 && ~x24 && ~x28 )
						nx_state = s1;
					else if( ~x15 && x31 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x15 && x31 && x19 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x15 && x31 && ~x19 )
						nx_state = s8;
					else if( ~x15 && ~x31 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else nx_state = s8;
				s9 : if( x15 && x19 && x13 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && x19 && ~x13 && x32 && x18 && x12 )
						nx_state = s9;
					else if( x15 && x19 && ~x13 && x32 && x18 && ~x12 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( x15 && x19 && ~x13 && x32 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x15 && x19 && ~x13 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && ~x19 )
						nx_state = s1;
					else if( ~x15 && x17 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x15 && x17 && x19 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x15 && x17 && ~x19 )
						nx_state = s9;
					else if( ~x15 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && ~x17 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && ~x17 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else nx_state = s9;
				s10 : if( x15 && x11 && x25 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( x15 && x11 && x25 && ~x3 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && x11 && x25 && ~x3 && ~x5 )
						nx_state = s10;
					else if( x15 && x11 && ~x25 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( x15 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && x44 && x47 )
						nx_state = s10;
					else if( ~x15 && x44 && ~x47 && x40 && x48 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && x44 && ~x47 && x40 && ~x48 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x44 && ~x47 && ~x40 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x44 && ~x47 && ~x40 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && ~x44 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else nx_state = s10;
				s11 : if( x15 && x7 && x35 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s16;
						end
					else if( x15 && x7 && x35 && ~x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x7 && ~x35 && x1 )
						nx_state = s11;
					else if( x15 && x7 && ~x35 && ~x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( x15 && ~x7 )
						nx_state = s11;
					else if( ~x15 && x3 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x15 && ~x3 && x2 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x15 && ~x3 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && ~x3 && ~x2 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else nx_state = s11;
				s12 : if( x15 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x15 && ~x5 && x34 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( x15 && ~x5 && ~x34 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x15 && x35 )
						nx_state = s1;
					else if( ~x15 && ~x35 && x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x15 && ~x35 && ~x13 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s14;
						end
					else nx_state = s12;
				s13 : if( x15 && x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( x15 && ~x10 && x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s11;
						end
					else if( x15 && ~x10 && ~x25 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x15 && x8 && x44 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x15 && x8 && ~x44 && x37 )
						nx_state = s1;
					else if( ~x15 && x8 && ~x44 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x15 && ~x8 && x48 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x15 && ~x8 && ~x48 && x37 )
						nx_state = s1;
					else if( ~x15 && ~x8 && ~x48 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else nx_state = s13;
				s14 : if( x15 && x2 && x8 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s16;
						end
					else if( x15 && x2 && x8 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x2 && x8 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( x15 && x2 && ~x8 && x32 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x15 && x2 && ~x8 && x32 && ~x1 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( x15 && x2 && ~x8 && x32 && ~x1 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s22;
						end
					else if( x15 && x2 && ~x8 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else if( x15 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x15 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && x37 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && ~x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else nx_state = s14;
				s15 : if( x15 && x16 && x19 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( x15 && x16 && x19 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && x16 && x19 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x16 && ~x19 && x1 && x26 && x30 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x15 && x16 && ~x19 && x1 && x26 && ~x30 )
						nx_state = s15;
					else if( x15 && x16 && ~x19 && x1 && ~x26 && x3 )
						nx_state = s15;
					else if( x15 && x16 && ~x19 && x1 && ~x26 && ~x3 && x30 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x15 && x16 && ~x19 && x1 && ~x26 && ~x3 && ~x30 )
						nx_state = s15;
					else if( x15 && x16 && ~x19 && ~x1 )
						nx_state = s15;
					else if( x15 && ~x16 )
						nx_state = s1;
					else if( ~x15 && x28 && x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x15 && x28 && ~x41 )
						nx_state = s15;
					else if( ~x15 && ~x28 && x27 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x15 && ~x28 && x27 && ~x8 && x37 )
						nx_state = s1;
					else if( ~x15 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x15 && ~x28 && ~x27 && x49 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && ~x28 && ~x27 && ~x49 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else nx_state = s15;
				s16 : if( x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s9;
						end
					else nx_state = s16;
				s17 : if( x15 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s23;
						end
					else if( x15 && ~x9 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && ~x9 && ~x3 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x15 && x29 && x49 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x15 && x29 && ~x49 )
						nx_state = s17;
					else if( ~x15 && ~x29 && x21 )
						nx_state = s1;
					else if( ~x15 && ~x29 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s7;
						end
					else nx_state = s17;
				s18 : if( x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s18;
						end
					else if( x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s14;
						end
					else if( x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else if( x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s16;
						end
					else if( x16 && ~x6 && ~x8 )
						nx_state = s1;
					else if( ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x16 && ~x10 )
						nx_state = s1;
					else nx_state = s18;
				s19 : if( x15 && x22 && x2 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( x15 && x22 && x2 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && x22 && x2 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( x15 && x22 && ~x2 )
						nx_state = s1;
					else if( x15 && ~x22 && x31 )
						nx_state = s1;
					else if( x15 && ~x22 && ~x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x15 && x46 && x3 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x15 && x46 && x3 && ~x23 )
						nx_state = s19;
					else if( ~x15 && x46 && ~x3 )
						nx_state = s1;
					else if( ~x15 && ~x46 && x2 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x15 && ~x46 && x2 && ~x23 )
						nx_state = s19;
					else if( ~x15 && ~x46 && ~x2 )
						nx_state = s1;
					else nx_state = s19;
				s20 : if( x9 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x9 && x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x9 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else nx_state = s20;
				s21 : if( 1'b1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s21;
				s22 : if( x15 && x25 && x22 )
						nx_state = s1;
					else if( x15 && x25 && ~x22 && x6 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( x15 && x25 && ~x22 && x6 && ~x8 )
						nx_state = s1;
					else if( x15 && x25 && ~x22 && ~x6 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( x15 && ~x25 && x29 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s6;
						end
					else if( x15 && ~x25 && ~x29 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x15 && x38 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x15 && ~x38 && x49 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x15 && ~x38 && ~x49 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s15;
						end
					else nx_state = s22;
				s23 : if( x15 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s19;
						end
					else if( x15 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s4;
						end
					else if( x15 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x15 && x49 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x15 && ~x49 )
						nx_state = s23;
					else nx_state = s23;
				s24 : if( x16 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s18;
						end
					else if( x16 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s5;
						end
					else nx_state = s24;

			default : nx_state = 0;
		endcase
	end
endmodule
