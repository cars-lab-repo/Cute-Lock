/******** Key Information: *********** 
Key 1:   bin: '11010000010001'    dec: 13329
Key 2:   bin: '01111011111011'    dec: 7931
Key 3:   bin: '01111100011100'    dec: 7964
Key 4:   bin: '00110101001101'    dec: 3405
**************************************/

module v1120 (keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, clk,rst,
	x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, 
	y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29);

input clk, rst, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14;
input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13;
output y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29;
reg[6:0] counter = 0;
reg y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29;

parameter s1=1, s2=2, s3=3, s4=4, s5=5, s6=6, s7=7, s8=8, s9=9, s10=10,
	s11=11, s12=12, s13=13, s14=14, s15=15, s16=16, s17=17, s18=18;
integer pr_state;
integer nx_state;

always @(negedge clk or posedge rst)
begin
	if (rst == 1'b1)
		counter <= 0;
	else
		counter <= (counter >= 35) ? 0 : counter + 1;
end

always@(  negedge clk or posedge rst )
begin
	if (rst == 1'b1)
	 begin
		pr_state = s1;
	end
	else
	begin
		if ( counter <= 8 ) begin 
			if ( keyinput0 == 1'b1 && keyinput1 == 1'b1 && keyinput2 == 1'b0 && keyinput3 == 1'b1 && keyinput4 == 1'b0 && keyinput5 == 1'b0 && keyinput6 == 1'b0 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b0 && keyinput11 == 1'b0 && keyinput12 == 1'b0 && keyinput13 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s15;
		end
		if ( counter > 8 && counter <= 17 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b1 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b1 && keyinput5 == 1'b0 && keyinput6 == 1'b1 && keyinput7 == 1'b1 && keyinput8 == 1'b1 && keyinput9 == 1'b1 && keyinput10 == 1'b1 && keyinput11 == 1'b0 && keyinput12 == 1'b1 && keyinput13 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s16;
		end
		if ( counter > 17 && counter <= 26 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b1 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b1 && keyinput5 == 1'b1 && keyinput6 == 1'b0 && keyinput7 == 1'b0 && keyinput8 == 1'b0 && keyinput9 == 1'b1 && keyinput10 == 1'b1 && keyinput11 == 1'b1 && keyinput12 == 1'b0 && keyinput13 == 1'b0 )
				pr_state = nx_state;
			else
				pr_state = s18;
		end
		if ( counter > 26 && counter <= 35 ) begin 
			if ( keyinput0 == 1'b0 && keyinput1 == 1'b0 && keyinput2 == 1'b1 && keyinput3 == 1'b1 && keyinput4 == 1'b0 && keyinput5 == 1'b1 && keyinput6 == 1'b0 && keyinput7 == 1'b1 && keyinput8 == 1'b0 && keyinput9 == 1'b0 && keyinput10 == 1'b1 && keyinput11 == 1'b1 && keyinput12 == 1'b0 && keyinput13 == 1'b1 )
				pr_state = nx_state;
			else
				pr_state = s14;
		end
	end
end


always@ ( pr_state or x1 or x2 or x3 or x4 or x5 or x6 or x7 or x8 or x9 or x10 or x11 or x12 or x13 or x14)
	begin
			y1 = 1'b0;	y2 = 1'b0;	y3 = 1'b0;	y4 = 1'b0;	
			y5 = 1'b0;	y6 = 1'b0;	y7 = 1'b0;	y8 = 1'b0;	
			y9 = 1'b0;	y10 = 1'b0;	y11 = 1'b0;	y12 = 1'b0;	
			y13 = 1'b0;	y14 = 1'b0;	y15 = 1'b0;	y16 = 1'b0;	
			y17 = 1'b0;	y18 = 1'b0;	y19 = 1'b0;	y20 = 1'b0;	
			y21 = 1'b0;	y22 = 1'b0;	y23 = 1'b0;	y24 = 1'b0;	
			y25 = 1'b0;	y26 = 1'b0;	y27 = 1'b0;	y28 = 1'b0;	
			y29 = 1'b0;	
		case ( pr_state )
				s1 : if( x10 && x12 && x11 && x13 && x1 && x3 && x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s2;
						end
					else if( x10 && x12 && x11 && x13 && x1 && x3 && ~x6 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x12 && x11 && x13 && x1 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x12 && x11 && x13 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( x10 && x12 && x11 && ~x13 && x5 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s4;
						end
					else if( x10 && x12 && x11 && ~x13 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x12 && ~x11 && x8 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( x10 && x12 && ~x11 && ~x8 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && x12 && ~x11 && ~x8 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && x13 && x11 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x1 && x5 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x1 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( x10 && ~x12 && ~x13 && x11 && x14 && x7 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( x10 && ~x12 && ~x13 && x11 && x14 && ~x7 && x1 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x12 && ~x13 && x11 && x14 && ~x7 && x1 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && ~x13 && x11 && x14 && ~x7 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( x10 && ~x12 && ~x13 && x11 && ~x14 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x10 && ~x12 && ~x13 && ~x11 && x1 && x14 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x12 && ~x13 && ~x11 && x1 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && ~x13 && ~x11 && x1 && ~x14 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && ~x12 && ~x13 && ~x11 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x10 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s1;
				s2 : if( x13 && x10 && x11 && x12 && x4 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( x13 && x10 && x11 && x12 && ~x4 )
						nx_state = s2;
					else if( x13 && x10 && x11 && ~x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && x10 && x11 && ~x12 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x13 && x10 && x11 && ~x12 && ~x3 && ~x2 )
						nx_state = s2;
					else if( x13 && x10 && ~x11 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && x10 && ~x11 && x12 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x13 && x10 && ~x11 && x12 && ~x3 && ~x2 )
						nx_state = s2;
					else if( x13 && x10 && ~x11 && ~x12 && x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && x10 && ~x11 && ~x12 && x14 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x13 && x10 && ~x11 && ~x12 && x14 && ~x3 && ~x2 )
						nx_state = s2;
					else if( x13 && x10 && ~x11 && ~x12 && ~x14 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x13 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && ~x10 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x13 && ~x10 && ~x3 && ~x2 )
						nx_state = s2;
					else if( ~x13 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x13 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x13 && ~x3 && ~x2 )
						nx_state = s2;
					else nx_state = s2;
				s3 : if( x10 && x12 && x11 && x3 && x4 && x13 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x10 && x12 && x11 && x3 && x4 && ~x13 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s13;
						end
					else if( x10 && x12 && x11 && x3 && ~x4 )
						nx_state = s3;
					else if( x10 && x12 && x11 && ~x3 && x4 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && x12 && x11 && ~x3 && ~x4 )
						nx_state = s3;
					else if( x10 && x12 && ~x11 && x4 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && x12 && ~x11 && ~x4 )
						nx_state = s3;
					else if( x10 && ~x12 && x13 && x11 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s2;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x3 && x4 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x3 && ~x4 )
						nx_state = s3;
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x3 && x4 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x3 && ~x4 )
						nx_state = s3;
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 )
						nx_state = s1;
					else if( x10 && ~x12 && ~x13 && x14 && x4 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && ~x12 && ~x13 && x14 && ~x4 )
						nx_state = s3;
					else if( x10 && ~x12 && ~x13 && ~x14 )
						nx_state = s1;
					else if( ~x10 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s2;
						end
					else nx_state = s3;
				s4 : if( x11 && x12 && x2 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( x11 && x12 && ~x2 )
						nx_state = s4;
					else if( x11 && ~x12 && x3 )
						nx_state = s1;
					else if( x11 && ~x12 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x11 && x3 )
						nx_state = s1;
					else if( ~x11 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else nx_state = s4;
				s5 : if( x12 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && x11 && x13 && x7 )
						nx_state = s1;
					else if( ~x12 && x11 && x13 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && ~x11 && x14 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && ~x11 && ~x14 && x7 )
						nx_state = s1;
					else if( ~x12 && ~x11 && ~x14 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else nx_state = s5;
				s6 : if( x12 && x11 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x12 && x11 && ~x3 && x2 )
						nx_state = s1;
					else if( x12 && x11 && ~x3 && ~x2 )
						nx_state = s6;
					else if( x12 && ~x11 && x10 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( x12 && ~x11 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x12 && ~x11 && ~x10 && ~x3 && x2 )
						nx_state = s1;
					else if( x12 && ~x11 && ~x10 && ~x3 && ~x2 )
						nx_state = s6;
					else if( ~x12 && x13 && x11 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && x13 && x11 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && x13 && x11 && ~x3 && ~x2 )
						nx_state = s6;
					else if( ~x12 && x13 && ~x11 && x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && x13 && ~x11 && x14 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && x13 && ~x11 && x14 && ~x3 && ~x2 )
						nx_state = s6;
					else if( ~x12 && x13 && ~x11 && ~x14 && x10 && x5 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && x10 && ~x5 && x1 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && x10 && ~x5 && ~x1 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && ~x10 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && x13 && ~x11 && ~x14 && ~x10 && ~x3 && ~x2 )
						nx_state = s6;
					else if( ~x12 && ~x13 && x14 && x10 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && ~x13 && x14 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && ~x13 && x14 && ~x10 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && ~x13 && x14 && ~x10 && ~x3 && ~x2 )
						nx_state = s6;
					else if( ~x12 && ~x13 && ~x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && ~x13 && ~x14 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && ~x13 && ~x14 && ~x3 && ~x2 )
						nx_state = s6;
					else nx_state = s6;
				s7 : if( x12 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x12 && x10 && x13 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && x2 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && x2 && ~x6 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && ~x2 )
						nx_state = s7;
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x12 && x10 && ~x13 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x12 && ~x10 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else nx_state = s7;
				s8 : if( x10 && x12 )
						nx_state = s1;
					else if( x10 && ~x12 && x13 && x11 && x2 && x4 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( x10 && ~x12 && x13 && x11 && x2 && ~x4 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x10 && ~x12 && x13 && x11 && ~x2 )
						nx_state = s8;
					else if( x10 && ~x12 && x13 && ~x11 && x14 )
						nx_state = s1;
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && x1 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s2;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && ~x1 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x10 && ~x12 && ~x13 && x14 )
						nx_state = s1;
					else if( x10 && ~x12 && ~x13 && ~x14 && x2 && x4 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( x10 && ~x12 && ~x13 && ~x14 && x2 && ~x4 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( x10 && ~x12 && ~x13 && ~x14 && ~x2 )
						nx_state = s8;
					else if( ~x10 && x2 && x4 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x10 && x2 && ~x4 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x10 && ~x2 )
						nx_state = s8;
					else nx_state = s8;
				s9 : if( x10 && x12 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x10 && ~x12 && x13 && x11 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x2 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x2 && ~x6 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x2 )
						nx_state = s9;
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x10 && ~x12 && ~x13 && x11 && x14 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( x10 && ~x12 && ~x13 && x11 && ~x14 && x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s11;
						end
					else if( x10 && ~x12 && ~x13 && x11 && ~x14 && ~x1 && x2 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && ~x12 && ~x13 && x11 && ~x14 && ~x1 && ~x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( x10 && ~x12 && ~x13 && ~x11 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x10 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s9;
				s10 : if( x10 && x12 && x11 && x13 && x3 && x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s2;
						end
					else if( x10 && x12 && x11 && x13 && x3 && ~x6 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x12 && x11 && x13 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x12 && x11 && ~x13 && x5 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s4;
						end
					else if( x10 && x12 && x11 && ~x13 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x12 && ~x11 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && x12 && ~x11 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && x13 && x11 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x5 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && x8 && x1 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && x8 && ~x1 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && ~x8 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x12 && ~x13 && x14 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x12 && ~x13 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x12 && ~x13 && ~x14 && x1 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s4;
						end
					else if( x10 && ~x12 && ~x13 && ~x14 && ~x1 && x3 )
						nx_state = s1;
					else if( x10 && ~x12 && ~x13 && ~x14 && ~x1 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x10 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s10;
				s11 : if( x12 && x11 && x10 && x13 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( x12 && x11 && x10 && x13 && ~x2 )
						nx_state = s11;
					else if( x12 && x11 && x10 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( x12 && x11 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( x12 && ~x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x14 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x14 && ~x11 && x10 && x13 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x14 && ~x11 && x10 && x13 && ~x2 )
						nx_state = s11;
					else if( ~x12 && x14 && ~x11 && x10 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x14 && ~x11 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && ~x14 && x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && ~x14 && ~x13 && x10 && x2 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && ~x14 && ~x13 && x10 && ~x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && ~x14 && ~x13 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s11;
				s12 : if( x13 && x10 && x11 && x12 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( x13 && x10 && x11 && ~x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && x10 && x11 && ~x12 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x13 && x10 && x11 && ~x12 && ~x3 && ~x6 )
						nx_state = s12;
					else if( x13 && x10 && ~x11 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && x10 && ~x11 && x12 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x13 && x10 && ~x11 && x12 && ~x3 && ~x6 )
						nx_state = s12;
					else if( x13 && x10 && ~x11 && ~x12 && x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && x10 && ~x11 && ~x12 && x14 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x13 && x10 && ~x11 && ~x12 && x14 && ~x3 && ~x6 )
						nx_state = s12;
					else if( x13 && x10 && ~x11 && ~x12 && ~x14 && x1 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( x13 && x10 && ~x11 && ~x12 && ~x14 && ~x1 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x13 && ~x10 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x13 && ~x10 && ~x3 && ~x6 )
						nx_state = s12;
					else if( ~x13 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x13 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x13 && ~x3 && ~x6 )
						nx_state = s12;
					else nx_state = s12;
				s13 : if( x2 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x2 )
						nx_state = s13;
					else nx_state = s13;
				s14 : if( x12 && x11 && x10 && x13 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && x11 && x10 && x13 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && x11 && x10 && x13 && ~x8 && ~x1 )
						nx_state = s14;
					else if( x12 && x11 && x10 && ~x13 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( x12 && x11 && ~x10 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && x11 && ~x10 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && x11 && ~x10 && ~x8 && ~x1 )
						nx_state = s14;
					else if( x12 && ~x11 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && ~x11 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && ~x11 && ~x8 && ~x1 )
						nx_state = s14;
					else if( ~x12 && x11 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x11 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x11 && ~x8 && ~x1 )
						nx_state = s14;
					else if( ~x12 && ~x11 && x14 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x11 && x14 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x11 && x14 && ~x8 && ~x1 )
						nx_state = s14;
					else if( ~x12 && ~x11 && ~x14 && x13 && x10 && x9 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && x10 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x12 && ~x11 && ~x14 && x13 && x10 && ~x9 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && ~x10 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && ~x10 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && ~x10 && ~x8 && ~x1 )
						nx_state = s14;
					else if( ~x12 && ~x11 && ~x14 && ~x13 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x11 && ~x14 && ~x13 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x11 && ~x14 && ~x13 && ~x8 && ~x1 )
						nx_state = s14;
					else nx_state = s14;
				s15 : if( x11 && x12 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( x11 && x12 && ~x4 )
						nx_state = s15;
					else if( x11 && ~x12 && x13 )
						nx_state = s1;
					else if( x11 && ~x12 && ~x13 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( x11 && ~x12 && ~x13 && ~x4 )
						nx_state = s15;
					else if( ~x11 && x14 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x11 && x14 && ~x4 )
						nx_state = s15;
					else if( ~x11 && ~x14 && x12 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x11 && ~x14 && x12 && ~x4 )
						nx_state = s15;
					else if( ~x11 && ~x14 && ~x12 && x13 )
						nx_state = s1;
					else if( ~x11 && ~x14 && ~x12 && ~x13 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x11 && ~x14 && ~x12 && ~x13 && ~x4 )
						nx_state = s15;
					else nx_state = s15;
				s16 : if( x10 && x13 && x11 && x12 && x3 && x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s2;
						end
					else if( x10 && x13 && x11 && x12 && x3 && ~x6 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x13 && x11 && x12 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x13 && x11 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x10 && x13 && ~x11 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && x13 && ~x11 && x12 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( x10 && x13 && ~x11 && x12 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( x10 && x13 && ~x11 && x12 && ~x3 && ~x1 && ~x7 )
						nx_state = s16;
					else if( x10 && x13 && ~x11 && ~x12 && x14 && x5 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s7;
						end
					else if( x10 && x13 && ~x11 && ~x12 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && x13 && ~x11 && ~x12 && ~x14 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x13 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x10 && ~x13 && x12 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( x10 && ~x13 && x12 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( x10 && ~x13 && x12 && ~x3 && ~x1 && ~x7 )
						nx_state = s16;
					else if( x10 && ~x13 && ~x12 && x14 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s6;
						end
					else if( x10 && ~x13 && ~x12 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( x10 && ~x13 && ~x12 && ~x14 && x1 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s4;
						end
					else if( x10 && ~x13 && ~x12 && ~x14 && ~x1 && x3 )
						nx_state = s1;
					else if( x10 && ~x13 && ~x12 && ~x14 && ~x1 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x10 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x10 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x10 && ~x3 && ~x1 && ~x7 )
						nx_state = s16;
					else nx_state = s16;
				s17 : if( x12 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( x12 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( x12 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( x12 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( x12 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s17;
					else if( ~x12 && x10 && x13 && x11 && x4 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x10 && x13 && x11 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s17;
					else if( ~x12 && x10 && ~x13 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x10 && ~x13 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && x10 && ~x13 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x12 && x10 && ~x13 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x10 && ~x13 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s17;
					else if( ~x12 && ~x10 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && ~x10 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x12 && ~x10 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x12 && ~x10 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && ~x10 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s17;
					else nx_state = s17;
				s18 : if( x12 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x12 && x10 && x13 && x11 && x5 && x6 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x12 && x10 && x13 && x11 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( ~x12 && x10 && x13 && x11 && x5 && ~x6 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x12 && x10 && x13 && x11 && ~x5 && x4 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x12 && x10 && x13 && x11 && ~x5 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && x4 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && ~x4 )
						nx_state = s18;
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x12 && x10 && ~x13 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x12 && ~x10 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s3;
						end
					else nx_state = s18;

			default : nx_state = 0;
		endcase
	end
endmodule
