// Benchmark "./test_runs/structural2_16keys_5bits--s-120240927_165426/ITC99/b20_encrypted" written by ABC on Fri Sep 27 18:24:09 2024

module b20_encrypted  ( clock, 
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, keyinput0, keyinput1, keyinput2,
    keyinput3, keyinput4,
    ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123  );
  input  clock;
  input  SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_,
    SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_,
    SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_,
    SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, keyinput0, keyinput1,
    keyinput2, keyinput3, keyinput4;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123;
  reg P1_IR_REG_0_, P1_IR_REG_1_, P1_IR_REG_2_, P1_IR_REG_3_, P1_IR_REG_4_,
    P1_IR_REG_5_, P1_IR_REG_6_, P1_IR_REG_7_, P1_IR_REG_8_, P1_IR_REG_9_,
    P1_IR_REG_10_, P1_IR_REG_11_, P1_IR_REG_12_, P1_IR_REG_13_,
    P1_IR_REG_14_, P1_IR_REG_15_, P1_IR_REG_16_, P1_IR_REG_17_,
    P1_IR_REG_18_, P1_IR_REG_19_, P1_IR_REG_20_, P1_IR_REG_21_,
    P1_IR_REG_22_, P1_IR_REG_23_, P1_IR_REG_24_, P1_IR_REG_25_,
    P1_IR_REG_26_, P1_IR_REG_27_, P1_IR_REG_28_, P1_IR_REG_29_,
    P1_IR_REG_30_, P1_IR_REG_31_, P1_D_REG_0_, P1_D_REG_1_, P1_D_REG_2_,
    P1_D_REG_3_, P1_D_REG_4_, P1_D_REG_5_, P1_D_REG_6_, P1_D_REG_7_,
    P1_D_REG_8_, P1_D_REG_9_, P1_D_REG_10_, P1_D_REG_11_, P1_D_REG_12_,
    P1_D_REG_13_, P1_D_REG_14_, P1_D_REG_15_, P1_D_REG_16_, P1_D_REG_17_,
    P1_D_REG_18_, P1_D_REG_19_, P1_D_REG_20_, P1_D_REG_21_, P1_D_REG_22_,
    P1_D_REG_23_, P1_D_REG_24_, P1_D_REG_25_, P1_D_REG_26_, P1_D_REG_27_,
    P1_D_REG_28_, P1_D_REG_29_, P1_D_REG_30_, P1_D_REG_31_, P1_REG0_REG_0_,
    P1_REG0_REG_1_, P1_REG0_REG_2_, P1_REG0_REG_3_, P1_REG0_REG_4_,
    P1_REG0_REG_5_, P1_REG0_REG_6_, P1_REG0_REG_7_, P1_REG0_REG_8_,
    P1_REG0_REG_9_, P1_REG0_REG_10_, P1_REG0_REG_11_, P1_REG0_REG_12_,
    P1_REG0_REG_13_, P1_REG0_REG_14_, P1_REG0_REG_15_, P1_REG0_REG_16_,
    P1_REG0_REG_17_, P1_REG0_REG_18_, P1_REG0_REG_19_, P1_REG0_REG_20_,
    P1_REG0_REG_21_, P1_REG0_REG_22_, P1_REG0_REG_23_, P1_REG0_REG_24_,
    P1_REG0_REG_25_, P1_REG0_REG_26_, P1_REG0_REG_27_, P1_REG0_REG_28_,
    P1_REG0_REG_29_, P1_REG0_REG_30_, P1_REG0_REG_31_, P1_REG1_REG_0_,
    P1_REG1_REG_1_, P1_REG1_REG_2_, P1_REG1_REG_3_, P1_REG1_REG_4_,
    P1_REG1_REG_5_, P1_REG1_REG_6_, P1_REG1_REG_7_, P1_REG1_REG_8_,
    P1_REG1_REG_9_, P1_REG1_REG_10_, P1_REG1_REG_11_, P1_REG1_REG_12_,
    P1_REG1_REG_13_, P1_REG1_REG_14_, P1_REG1_REG_15_, P1_REG1_REG_16_,
    P1_REG1_REG_17_, P1_REG1_REG_18_, P1_REG1_REG_19_, P1_REG1_REG_20_,
    P1_REG1_REG_21_, P1_REG1_REG_22_, P1_REG1_REG_23_, P1_REG1_REG_24_,
    P1_REG1_REG_25_, P1_REG1_REG_26_, P1_REG1_REG_27_, P1_REG1_REG_28_,
    P1_REG1_REG_29_, P1_REG1_REG_30_, P1_REG1_REG_31_, P1_REG2_REG_0_,
    P1_REG2_REG_1_, P1_REG2_REG_2_, P1_REG2_REG_3_, P1_REG2_REG_4_,
    P1_REG2_REG_5_, P1_REG2_REG_6_, P1_REG2_REG_7_, P1_REG2_REG_8_,
    P1_REG2_REG_9_, P1_REG2_REG_10_, P1_REG2_REG_11_, P1_REG2_REG_12_,
    P1_REG2_REG_13_, P1_REG2_REG_14_, P1_REG2_REG_15_, P1_REG2_REG_16_,
    P1_REG2_REG_17_, P1_REG2_REG_18_, P1_REG2_REG_19_, P1_REG2_REG_20_,
    P1_REG2_REG_21_, P1_REG2_REG_22_, P1_REG2_REG_23_, P1_REG2_REG_24_,
    P1_REG2_REG_25_, P1_REG2_REG_26_, P1_REG2_REG_27_, P1_REG2_REG_28_,
    P1_REG2_REG_29_, P1_REG2_REG_30_, P1_REG2_REG_31_, P1_ADDR_REG_19_,
    P1_ADDR_REG_18_, P1_ADDR_REG_17_, P1_ADDR_REG_16_, P1_ADDR_REG_15_,
    P1_ADDR_REG_14_, P1_ADDR_REG_13_, P1_ADDR_REG_12_, P1_ADDR_REG_11_,
    P1_ADDR_REG_10_, P1_ADDR_REG_9_, P1_ADDR_REG_8_, P1_ADDR_REG_7_,
    P1_ADDR_REG_6_, P1_ADDR_REG_5_, P1_ADDR_REG_4_, P1_ADDR_REG_3_,
    P1_ADDR_REG_2_, P1_ADDR_REG_1_, P1_ADDR_REG_0_, P1_DATAO_REG_0_,
    P1_DATAO_REG_1_, P1_DATAO_REG_2_, P1_DATAO_REG_3_, P1_DATAO_REG_4_,
    P1_DATAO_REG_5_, P1_DATAO_REG_6_, P1_DATAO_REG_7_, P1_DATAO_REG_8_,
    P1_DATAO_REG_9_, P1_DATAO_REG_10_, P1_DATAO_REG_11_, P1_DATAO_REG_12_,
    P1_DATAO_REG_13_, P1_DATAO_REG_14_, P1_DATAO_REG_15_, P1_DATAO_REG_16_,
    P1_DATAO_REG_17_, P1_DATAO_REG_18_, P1_DATAO_REG_19_, P1_DATAO_REG_20_,
    P1_DATAO_REG_21_, P1_DATAO_REG_22_, P1_DATAO_REG_23_, P1_DATAO_REG_24_,
    P1_DATAO_REG_25_, P1_DATAO_REG_26_, P1_DATAO_REG_27_, P1_DATAO_REG_28_,
    P1_DATAO_REG_29_, P1_DATAO_REG_30_, P1_DATAO_REG_31_, P1_B_REG,
    P1_REG3_REG_15_, P1_REG3_REG_26_, P1_REG3_REG_6_, P1_REG3_REG_18_,
    P1_REG3_REG_2_, P1_REG3_REG_11_, P1_REG3_REG_22_, P1_REG3_REG_13_,
    P1_REG3_REG_20_, P1_REG3_REG_0_, P1_REG3_REG_9_, P1_REG3_REG_4_,
    P1_REG3_REG_24_, P1_REG3_REG_17_, P1_REG3_REG_5_, P1_REG3_REG_16_,
    P1_REG3_REG_25_, P1_REG3_REG_12_, P1_REG3_REG_21_, P1_REG3_REG_1_,
    P1_REG3_REG_8_, P1_REG3_REG_28_, P1_REG3_REG_19_, P1_REG3_REG_3_,
    P1_REG3_REG_10_, P1_REG3_REG_23_, P1_REG3_REG_14_, P1_REG3_REG_27_,
    P1_REG3_REG_7_, P1_STATE_REG, P1_RD_REG, P1_WR_REG, P2_IR_REG_0_,
    P2_IR_REG_1_, P2_IR_REG_2_, P2_IR_REG_3_, P2_IR_REG_4_, P2_IR_REG_5_,
    P2_IR_REG_6_, P2_IR_REG_7_, P2_IR_REG_8_, P2_IR_REG_9_, P2_IR_REG_10_,
    P2_IR_REG_11_, P2_IR_REG_12_, P2_IR_REG_13_, P2_IR_REG_14_,
    P2_IR_REG_15_, P2_IR_REG_16_, P2_IR_REG_17_, P2_IR_REG_18_,
    P2_IR_REG_19_, P2_IR_REG_20_, P2_IR_REG_21_, P2_IR_REG_22_,
    P2_IR_REG_23_, P2_IR_REG_24_, P2_IR_REG_25_, P2_IR_REG_26_,
    P2_IR_REG_27_, P2_IR_REG_28_, P2_IR_REG_29_, P2_IR_REG_30_,
    P2_IR_REG_31_, P2_D_REG_0_, P2_D_REG_1_, P2_D_REG_2_, P2_D_REG_3_,
    P2_D_REG_4_, P2_D_REG_5_, P2_D_REG_6_, P2_D_REG_7_, P2_D_REG_8_,
    P2_D_REG_9_, P2_D_REG_10_, P2_D_REG_11_, P2_D_REG_12_, P2_D_REG_13_,
    P2_D_REG_14_, P2_D_REG_15_, P2_D_REG_16_, P2_D_REG_17_, P2_D_REG_18_,
    P2_D_REG_19_, P2_D_REG_20_, P2_D_REG_21_, P2_D_REG_22_, P2_D_REG_23_,
    P2_D_REG_24_, P2_D_REG_25_, P2_D_REG_26_, P2_D_REG_27_, P2_D_REG_28_,
    P2_D_REG_29_, P2_D_REG_30_, P2_D_REG_31_, P2_REG0_REG_0_,
    P2_REG0_REG_1_, P2_REG0_REG_2_, P2_REG0_REG_3_, P2_REG0_REG_4_,
    P2_REG0_REG_5_, P2_REG0_REG_6_, P2_REG0_REG_7_, P2_REG0_REG_8_,
    P2_REG0_REG_9_, P2_REG0_REG_10_, P2_REG0_REG_11_, P2_REG0_REG_12_,
    P2_REG0_REG_13_, P2_REG0_REG_14_, P2_REG0_REG_15_, P2_REG0_REG_16_,
    P2_REG0_REG_17_, P2_REG0_REG_18_, P2_REG0_REG_19_, P2_REG0_REG_20_,
    P2_REG0_REG_21_, P2_REG0_REG_22_, P2_REG0_REG_23_, P2_REG0_REG_24_,
    P2_REG0_REG_25_, P2_REG0_REG_26_, P2_REG0_REG_27_, P2_REG0_REG_28_,
    P2_REG0_REG_29_, P2_REG0_REG_30_, P2_REG0_REG_31_, P2_REG1_REG_0_,
    P2_REG1_REG_1_, P2_REG1_REG_2_, P2_REG1_REG_3_, P2_REG1_REG_4_,
    P2_REG1_REG_5_, P2_REG1_REG_6_, P2_REG1_REG_7_, P2_REG1_REG_8_,
    P2_REG1_REG_9_, P2_REG1_REG_10_, P2_REG1_REG_11_, P2_REG1_REG_12_,
    P2_REG1_REG_13_, P2_REG1_REG_14_, P2_REG1_REG_15_, P2_REG1_REG_16_,
    P2_REG1_REG_17_, P2_REG1_REG_18_, P2_REG1_REG_19_, P2_REG1_REG_20_,
    P2_REG1_REG_21_, P2_REG1_REG_22_, P2_REG1_REG_23_, P2_REG1_REG_24_,
    P2_REG1_REG_25_, P2_REG1_REG_26_, P2_REG1_REG_27_, P2_REG1_REG_28_,
    P2_REG1_REG_29_, P2_REG1_REG_30_, P2_REG1_REG_31_, P2_REG2_REG_0_,
    P2_REG2_REG_1_, P2_REG2_REG_2_, P2_REG2_REG_3_, P2_REG2_REG_4_,
    P2_REG2_REG_5_, P2_REG2_REG_6_, P2_REG2_REG_7_, P2_REG2_REG_8_,
    P2_REG2_REG_9_, P2_REG2_REG_10_, P2_REG2_REG_11_, P2_REG2_REG_12_,
    P2_REG2_REG_13_, P2_REG2_REG_14_, P2_REG2_REG_15_, P2_REG2_REG_16_,
    P2_REG2_REG_17_, P2_REG2_REG_18_, P2_REG2_REG_19_, P2_REG2_REG_20_,
    P2_REG2_REG_21_, P2_REG2_REG_22_, P2_REG2_REG_23_, P2_REG2_REG_24_,
    P2_REG2_REG_25_, P2_REG2_REG_26_, P2_REG2_REG_27_, P2_REG2_REG_28_,
    P2_REG2_REG_29_, P2_REG2_REG_30_, P2_REG2_REG_31_, P2_ADDR_REG_19_,
    P2_ADDR_REG_18_, P2_ADDR_REG_17_, P2_ADDR_REG_16_, P2_ADDR_REG_15_,
    P2_ADDR_REG_14_, P2_ADDR_REG_13_, P2_ADDR_REG_12_, P2_ADDR_REG_11_,
    P2_ADDR_REG_10_, P2_ADDR_REG_9_, P2_ADDR_REG_8_, P2_ADDR_REG_7_,
    P2_ADDR_REG_6_, P2_ADDR_REG_5_, P2_ADDR_REG_4_, P2_ADDR_REG_3_,
    P2_ADDR_REG_2_, P2_ADDR_REG_1_, P2_ADDR_REG_0_, P2_DATAO_REG_0_,
    P2_DATAO_REG_1_, P2_DATAO_REG_2_, P2_DATAO_REG_3_, P2_DATAO_REG_4_,
    P2_DATAO_REG_5_, P2_DATAO_REG_6_, P2_DATAO_REG_7_, P2_DATAO_REG_8_,
    P2_DATAO_REG_9_, P2_DATAO_REG_10_, P2_DATAO_REG_11_, P2_DATAO_REG_12_,
    P2_DATAO_REG_13_, P2_DATAO_REG_14_, P2_DATAO_REG_15_, P2_DATAO_REG_16_,
    P2_DATAO_REG_17_, P2_DATAO_REG_18_, P2_DATAO_REG_19_, P2_DATAO_REG_20_,
    P2_DATAO_REG_21_, P2_DATAO_REG_22_, P2_DATAO_REG_23_, P2_DATAO_REG_24_,
    P2_DATAO_REG_25_, P2_DATAO_REG_26_, P2_DATAO_REG_27_, P2_DATAO_REG_28_,
    P2_DATAO_REG_29_, P2_DATAO_REG_30_, P2_DATAO_REG_31_, P2_B_REG,
    P2_REG3_REG_15_, P2_REG3_REG_26_, P2_REG3_REG_6_, P2_REG3_REG_18_,
    P2_REG3_REG_2_, P2_REG3_REG_11_, P2_REG3_REG_22_, P2_REG3_REG_13_,
    P2_REG3_REG_20_, P2_REG3_REG_0_, P2_REG3_REG_9_, P2_REG3_REG_4_,
    P2_REG3_REG_24_, P2_REG3_REG_17_, P2_REG3_REG_5_, P2_REG3_REG_16_,
    P2_REG3_REG_25_, P2_REG3_REG_12_, P2_REG3_REG_21_, P2_REG3_REG_1_,
    P2_REG3_REG_8_, P2_REG3_REG_28_, P2_REG3_REG_19_, P2_REG3_REG_3_,
    P2_REG3_REG_10_, P2_REG3_REG_23_, P2_REG3_REG_14_, P2_REG3_REG_27_,
    P2_REG3_REG_7_, P2_STATE_REG, P2_RD_REG, P2_WR_REG, Q_0, Q_1, Q_2, Q_3;
  wire new_P2_R1161_U504, new_P2_R1161_U503, new_P2_R1161_U502, new_U25,
    new_U26, new_U27, new_U28, new_U29, new_U30, new_U31, new_U32, new_U33,
    new_U34, new_U35, new_U36, new_U37, new_U38, new_U39, new_U40, new_U41,
    new_U42, new_U43, new_U44, new_U45, new_U46, new_U47, new_U48, new_U49,
    new_U50, new_U51, new_U52, new_U53, new_U54, new_U55, new_U56, new_U57,
    new_U58, new_U59, new_U60, new_U61, new_U62, new_U63, new_U64, new_U65,
    new_U66, new_U67, new_U68, new_U69, new_U70, new_U71, new_U72, new_U73,
    new_U74, new_U75, new_U76, new_U77, new_U78, new_U79, new_U80, new_U81,
    new_U82, new_U83, new_U84, new_U85, new_U86, new_U87, new_U88, new_U89,
    new_U90, new_U91, new_U92, new_U93, new_U94, new_U95, new_U96, new_U97,
    new_U98, new_U99, new_U100, new_U101, new_U102, new_U103, new_U104,
    new_U105, new_U106, new_U107, new_U108, new_U109, new_U110, new_U111,
    new_U112, new_U113, new_U114, new_U115, new_U116, new_U117, new_U118,
    new_U119, new_U120, new_U121, new_U122, new_U124, new_U125, new_U127,
    new_U128, new_U129, new_U130, new_U131, new_U132, new_U133, new_U134,
    new_U135, new_U136, new_U137, new_U138, new_U139, new_U140, new_U141,
    new_U142, new_U143, new_U144, new_U145, new_U146, new_U147, new_U148,
    new_U149, new_U150, new_U151, new_U152, new_U153, new_U154, new_U155,
    new_U156, new_U157, new_U158, new_U159, new_U160, new_U161, new_U162,
    new_U163, new_U164, new_U165, new_U166, new_U167, new_U168, new_U169,
    new_U170, new_U171, new_U172, new_U173, new_U174, new_U175, new_U176,
    new_U177, new_U178, new_U179, new_U180, new_U181, new_U182, new_U183,
    new_U184, new_U185, new_U186, new_U187, new_U188, new_U189, new_U190,
    new_U191, new_U192, new_U193, new_U194, new_U195, new_U196, new_U197,
    new_U198, new_U199, new_U200, new_U201, new_U202, new_U203, new_U204,
    new_U205, new_U206, new_U207, new_U208, new_U209, new_U210, new_U211,
    new_U212, new_U213, new_U214, new_U215, new_U216, new_U217, new_U218,
    new_U219, new_U220, new_U221, new_U222, new_U223, new_U224, new_U225,
    new_U226, new_U227, new_U228, new_U229, new_U230, new_U231, new_U232,
    new_U233, new_U234, new_U235, new_U236, new_U237, new_U238, new_U239,
    new_U240, new_U241, new_U242, new_U243, new_U244, new_U245, new_U246,
    new_U247, new_U248, new_U249, new_U250, new_U251, new_U252, new_U253,
    new_U254, new_U255, new_U256, new_U257, new_U258, new_U259, new_U260,
    new_U261, new_U262, new_U263, new_U264, new_U265, new_U266, new_U267,
    new_U268, new_U269, new_U270, new_U271, new_U272, new_U273, new_U274,
    new_U275, new_U276, new_U277, new_U278, new_U279, new_U280, new_U281,
    new_U282, new_U283, new_U284, new_U285, new_U286, new_U287, new_U288,
    new_U289, new_U290, new_U291, new_U292, new_U293, new_U294, new_U295,
    new_U296, new_U297, new_U298, new_U299, new_U300, new_U301, new_U302,
    new_U303, new_U304, new_U305, new_U306, new_U307, new_U308, new_U309,
    new_U310, new_U311, new_U312, new_U313, new_U314, new_U315, new_U316,
    new_U317, new_U318, new_U319, new_U320, new_U321, new_U322, new_U323,
    new_U324, new_U325, new_U326, new_P2_R1161_U501, new_P2_R1161_U500,
    new_P2_R1161_U499, new_P2_R1161_U498, new_P2_R1161_U497,
    new_P2_R1161_U496, new_P2_R1161_U495, new_P2_R1161_U494,
    new_P2_R1161_U493, new_P2_R1161_U492, new_P2_R1161_U491,
    new_P2_R1161_U490, new_P1_U3014, new_P1_U3015, new_P1_U3016,
    new_P1_U3017, new_P1_U3018, new_P1_U3019, new_P1_U3020, new_P1_U3021,
    new_P1_U3022, new_P1_U3023, new_P1_U3024, new_P1_U3025, new_P1_U3026,
    new_P1_U3027, new_P1_U3028, new_P1_U3029, new_P1_U3030, new_P1_U3031,
    new_P1_U3032, new_P1_U3033, new_P1_U3034, new_P1_U3035, new_P1_U3036,
    new_P1_U3037, new_P1_U3038, new_P1_U3039, new_P1_U3040, new_P1_U3041,
    new_P1_U3042, new_P1_U3043, new_P1_U3044, new_P1_U3045, new_P1_U3046,
    new_P1_U3047, new_P1_U3048, new_P1_U3049, new_P1_U3050, new_P1_U3051,
    new_P1_U3052, new_P1_U3053, new_P1_U3054, new_P1_U3055, new_P1_U3056,
    new_P1_U3057, new_P1_U3058, new_P1_U3059, new_P1_U3060, new_P1_U3061,
    new_P1_U3062, new_P1_U3063, new_P1_U3064, new_P1_U3065, new_P1_U3066,
    new_P1_U3067, new_P1_U3068, new_P1_U3069, new_P1_U3070, new_P1_U3071,
    new_P1_U3072, new_P1_U3073, new_P1_U3074, new_P1_U3075, new_P1_U3076,
    new_P1_U3077, new_P1_U3078, new_P1_U3079, new_P1_U3080, new_P1_U3081,
    new_P1_U3082, new_P1_U3083, new_P1_U3084, new_P1_U3087, new_P1_U3088,
    new_P1_U3089, new_P1_U3090, new_P1_U3091, new_P1_U3092, new_P1_U3093,
    new_P1_U3094, new_P1_U3095, new_P1_U3096, new_P1_U3097, new_P1_U3098,
    new_P1_U3099, new_P1_U3100, new_P1_U3101, new_P1_U3102, new_P1_U3103,
    new_P1_U3104, new_P1_U3105, new_P1_U3106, new_P1_U3107, new_P1_U3108,
    new_P1_U3109, new_P1_U3110, new_P1_U3111, new_P1_U3112, new_P1_U3113,
    new_P1_U3114, new_P1_U3115, new_P1_U3116, new_P1_U3117, new_P1_U3118,
    new_P1_U3119, new_P1_U3120, new_P1_U3121, new_P1_U3122, new_P1_U3123,
    new_P1_U3124, new_P1_U3125, new_P1_U3126, new_P1_U3127, new_P1_U3128,
    new_P1_U3129, new_P1_U3130, new_P1_U3131, new_P1_U3132, new_P1_U3133,
    new_P1_U3134, new_P1_U3135, new_P1_U3136, new_P1_U3137, new_P1_U3138,
    new_P1_U3139, new_P1_U3140, new_P1_U3141, new_P1_U3142, new_P1_U3143,
    new_P1_U3144, new_P1_U3145, new_P1_U3146, new_P1_U3147, new_P1_U3148,
    new_P1_U3149, new_P1_U3150, new_P1_U3151, new_P1_U3152, new_P1_U3153,
    new_P1_U3154, new_P1_U3155, new_P1_U3156, new_P1_U3157, new_P1_U3158,
    new_P1_U3159, new_P1_U3160, new_P1_U3161, new_P1_U3162, new_P1_U3163,
    new_P1_U3164, new_P1_U3165, new_P1_U3166, new_P1_U3167, new_P1_U3168,
    new_P1_U3169, new_P1_U3170, new_P1_U3171, new_P1_U3172, new_P1_U3173,
    new_P1_U3174, new_P1_U3175, new_P1_U3176, new_P1_U3177, new_P1_U3178,
    new_P1_U3179, new_P1_U3180, new_P1_U3181, new_P1_U3182, new_P1_U3183,
    new_P1_U3184, new_P1_U3185, new_P1_U3186, new_P1_U3187, new_P1_U3188,
    new_P1_U3189, new_P1_U3190, new_P1_U3191, new_P1_U3192, new_P1_U3193,
    new_P1_U3194, new_P1_U3195, new_P1_U3196, new_P1_U3197, new_P1_U3198,
    new_P1_U3199, new_P1_U3200, new_P1_U3201, new_P1_U3202, new_P1_U3203,
    new_P1_U3204, new_P1_U3205, new_P1_U3206, new_P1_U3207, new_P1_U3208,
    new_P1_U3209, new_P1_U3210, new_P1_U3211, new_P1_U3212, new_P1_U3355,
    new_P1_U3357, new_P1_U3358, new_P1_U3359, new_P1_U3360, new_P1_U3361,
    new_P1_U3362, new_P1_U3363, new_P1_U3364, new_P1_U3365, new_P1_U3366,
    new_P1_U3367, new_P1_U3368, new_P1_U3369, new_P1_U3370, new_P1_U3371,
    new_P1_U3372, new_P1_U3373, new_P1_U3374, new_P1_U3375, new_P1_U3376,
    new_P1_U3377, new_P1_U3378, new_P1_U3379, new_P1_U3380, new_P1_U3381,
    new_P1_U3382, new_P1_U3383, new_P1_U3384, new_P1_U3385, new_P1_U3386,
    new_P1_U3387, new_P1_U3388, new_P1_U3389, new_P1_U3390, new_P1_U3391,
    new_P1_U3392, new_P1_U3393, new_P1_U3394, new_P1_U3395, new_P1_U3396,
    new_P1_U3397, new_P1_U3398, new_P1_U3399, new_P1_U3400, new_P1_U3401,
    new_P1_U3402, new_P1_U3403, new_P1_U3404, new_P1_U3405, new_P1_U3406,
    new_P1_U3407, new_P1_U3408, new_P1_U3409, new_P1_U3410, new_P1_U3411,
    new_P1_U3412, new_P1_U3413, new_P1_U3414, new_P1_U3415, new_P1_U3416,
    new_P1_U3417, new_P1_U3418, new_P1_U3419, new_P1_U3420, new_P1_U3421,
    new_P1_U3422, new_P1_U3423, new_P1_U3424, new_P1_U3425, new_P1_U3426,
    new_P1_U3427, new_P1_U3428, new_P1_U3429, new_P1_U3430, new_P1_U3431,
    new_P1_U3432, new_P1_U3433, new_P1_U3434, new_P1_U3435, new_P1_U3436,
    new_P1_U3437, new_P1_U3438, new_P1_U3441, new_P1_U3442, new_P1_U3443,
    new_P1_U3444, new_P1_U3445, new_P1_U3446, new_P1_U3447, new_P1_U3448,
    new_P1_U3449, new_P1_U3450, new_P1_U3451, new_P1_U3452, new_P1_U3454,
    new_P1_U3455, new_P1_U3457, new_P1_U3458, new_P1_U3460, new_P1_U3461,
    new_P1_U3463, new_P1_U3464, new_P1_U3466, new_P1_U3467, new_P1_U3469,
    new_P1_U3470, new_P1_U3472, new_P1_U3473, new_P1_U3475, new_P1_U3476,
    new_P1_U3478, new_P1_U3479, new_P1_U3481, new_P1_U3482, new_P1_U3484,
    new_P1_U3485, new_P1_U3487, new_P1_U3488, new_P1_U3490, new_P1_U3491,
    new_P1_U3493, new_P1_U3494, new_P1_U3496, new_P1_U3497, new_P1_U3499,
    new_P1_U3500, new_P1_U3502, new_P1_U3503, new_P1_U3505, new_P1_U3506,
    new_P1_U3508, new_P1_U3586, new_P1_U3587, new_P1_U3588, new_P1_U3589,
    new_P1_U3590, new_P1_U3591, new_P1_U3592, new_P1_U3593, new_P1_U3594,
    new_P1_U3595, new_P1_U3596, new_P1_U3597, new_P1_U3598, new_P1_U3599,
    new_P1_U3600, new_P1_U3601, new_P1_U3602, new_P1_U3603, new_P1_U3604,
    new_P1_U3605, new_P1_U3606, new_P1_U3607, new_P1_U3608, new_P1_U3609,
    new_P1_U3610, new_P1_U3611, new_P1_U3612, new_P1_U3613, new_P1_U3614,
    new_P1_U3615, new_P1_U3616, new_P1_U3617, new_P1_U3618, new_P1_U3619,
    new_P1_U3620, new_P1_U3621, new_P1_U3622, new_P1_U3623, new_P1_U3624,
    new_P1_U3625, new_P1_U3626, new_P1_U3627, new_P1_U3628, new_P1_U3629,
    new_P1_U3630, new_P1_U3631, new_P1_U3632, new_P1_U3633, new_P1_U3634,
    new_P1_U3635, new_P1_U3636, new_P1_U3637, new_P1_U3638, new_P1_U3639,
    new_P1_U3640, new_P1_U3641, new_P1_U3642, new_P1_U3643, new_P1_U3644,
    new_P1_U3645, new_P1_U3646, new_P1_U3647, new_P1_U3648, new_P1_U3649,
    new_P1_U3650, new_P1_U3651, new_P1_U3652, new_P1_U3653, new_P1_U3654,
    new_P1_U3655, new_P1_U3656, new_P1_U3657, new_P1_U3658, new_P1_U3659,
    new_P1_U3660, new_P1_U3661, new_P1_U3662, new_P1_U3663, new_P1_U3664,
    new_P1_U3665, new_P1_U3666, new_P1_U3667, new_P1_U3668, new_P1_U3669,
    new_P1_U3670, new_P1_U3671, new_P1_U3672, new_P1_U3673, new_P1_U3674,
    new_P1_U3675, new_P1_U3676, new_P1_U3677, new_P1_U3678, new_P1_U3679,
    new_P1_U3680, new_P1_U3681, new_P1_U3682, new_P1_U3683, new_P1_U3684,
    new_P1_U3685, new_P1_U3686, new_P1_U3687, new_P1_U3688, new_P1_U3689,
    new_P1_U3690, new_P1_U3691, new_P1_U3692, new_P1_U3693, new_P1_U3694,
    new_P1_U3695, new_P1_U3696, new_P1_U3697, new_P1_U3698, new_P1_U3699,
    new_P1_U3700, new_P1_U3701, new_P1_U3702, new_P1_U3703, new_P1_U3704,
    new_P1_U3705, new_P1_U3706, new_P1_U3707, new_P1_U3708, new_P1_U3709,
    new_P1_U3710, new_P1_U3711, new_P1_U3712, new_P1_U3713, new_P1_U3714,
    new_P1_U3715, new_P1_U3716, new_P1_U3717, new_P1_U3718, new_P1_U3719,
    new_P1_U3720, new_P1_U3721, new_P1_U3722, new_P1_U3723, new_P1_U3724,
    new_P1_U3725, new_P1_U3726, new_P1_U3727, new_P1_U3728, new_P1_U3729,
    new_P1_U3730, new_P1_U3731, new_P1_U3732, new_P1_U3733, new_P1_U3734,
    new_P1_U3735, new_P1_U3736, new_P1_U3737, new_P1_U3738, new_P1_U3739,
    new_P1_U3740, new_P1_U3741, new_P1_U3742, new_P1_U3743, new_P1_U3744,
    new_P1_U3745, new_P1_U3746, new_P1_U3747, new_P1_U3748, new_P1_U3749,
    new_P1_U3750, new_P1_U3751, new_P1_U3752, new_P1_U3753, new_P1_U3754,
    new_P1_U3755, new_P1_U3756, new_P1_U3757, new_P1_U3758, new_P1_U3759,
    new_P1_U3760, new_P1_U3761, new_P1_U3762, new_P1_U3763, new_P1_U3764,
    new_P1_U3765, new_P1_U3766, new_P1_U3767, new_P1_U3768, new_P1_U3769,
    new_P1_U3770, new_P1_U3771, new_P1_U3772, new_P1_U3773, new_P1_U3774,
    new_P1_U3775, new_P1_U3776, new_P1_U3777, new_P1_U3778, new_P1_U3779,
    new_P1_U3780, new_P1_U3781, new_P1_U3782, new_P1_U3783, new_P1_U3784,
    new_P1_U3785, new_P1_U3786, new_P1_U3787, new_P1_U3788, new_P1_U3789,
    new_P1_U3790, new_P1_U3791, new_P1_U3792, new_P1_U3793, new_P1_U3794,
    new_P1_U3795, new_P1_U3796, new_P1_U3797, new_P1_U3798, new_P1_U3799,
    new_P1_U3800, new_P1_U3801, new_P1_U3802, new_P1_U3803, new_P1_U3804,
    new_P1_U3805, new_P1_U3806, new_P1_U3807, new_P1_U3808, new_P1_U3809,
    new_P1_U3810, new_P1_U3811, new_P1_U3812, new_P1_U3813, new_P1_U3814,
    new_P1_U3815, new_P1_U3816, new_P1_U3817, new_P1_U3818, new_P1_U3819,
    new_P1_U3820, new_P1_U3821, new_P1_U3822, new_P1_U3823, new_P1_U3824,
    new_P1_U3825, new_P1_U3826, new_P1_U3827, new_P1_U3828, new_P1_U3829,
    new_P1_U3830, new_P1_U3831, new_P1_U3832, new_P1_U3833, new_P1_U3834,
    new_P1_U3835, new_P1_U3836, new_P1_U3837, new_P1_U3838, new_P1_U3839,
    new_P1_U3840, new_P1_U3841, new_P1_U3842, new_P1_U3843, new_P1_U3844,
    new_P1_U3845, new_P1_U3846, new_P1_U3847, new_P1_U3848, new_P1_U3849,
    new_P1_U3850, new_P1_U3851, new_P1_U3852, new_P1_U3853, new_P1_U3854,
    new_P1_U3855, new_P1_U3856, new_P1_U3857, new_P1_U3858, new_P1_U3859,
    new_P1_U3860, new_P1_U3861, new_P1_U3862, new_P1_U3863, new_P1_U3864,
    new_P1_U3865, new_P1_U3866, new_P1_U3867, new_P1_U3868, new_P1_U3869,
    new_P1_U3870, new_P1_U3871, new_P1_U3872, new_P1_U3873, new_P1_U3874,
    new_P1_U3875, new_P1_U3876, new_P1_U3877, new_P1_U3878, new_P1_U3879,
    new_P1_U3880, new_P1_U3881, new_P1_U3882, new_P1_U3883, new_P1_U3884,
    new_P1_U3885, new_P1_U3886, new_P1_U3887, new_P1_U3888, new_P1_U3889,
    new_P1_U3890, new_P1_U3891, new_P1_U3892, new_P1_U3893, new_P1_U3894,
    new_P1_U3895, new_P1_U3896, new_P1_U3897, new_P1_U3898, new_P1_U3899,
    new_P1_U3900, new_P1_U3901, new_P1_U3902, new_P1_U3903, new_P1_U3904,
    new_P1_U3905, new_P1_U3906, new_P1_U3907, new_P1_U3908, new_P1_U3909,
    new_P1_U3910, new_P1_U3911, new_P1_U3912, new_P1_U3913, new_P1_U3914,
    new_P1_U3915, new_P1_U3916, new_P1_U3917, new_P1_U3918, new_P1_U3919,
    new_P1_U3920, new_P1_U3921, new_P1_U3922, new_P1_U3923, new_P1_U3924,
    new_P1_U3925, new_P1_U3926, new_P1_U3927, new_P1_U3928, new_P1_U3929,
    new_P1_U3930, new_P1_U3931, new_P1_U3932, new_P1_U3933, new_P1_U3934,
    new_P1_U3935, new_P1_U3936, new_P1_U3937, new_P1_U3938, new_P1_U3939,
    new_P1_U3940, new_P1_U3941, new_P1_U3942, new_P1_U3943, new_P1_U3944,
    new_P1_U3945, new_P1_U3946, new_P1_U3947, new_P1_U3948, new_P1_U3949,
    new_P1_U3950, new_P1_U3951, new_P1_U3952, new_P1_U3953, new_P1_U3954,
    new_P1_U3955, new_P1_U3956, new_P1_U3957, new_P1_U3958, new_P1_U3959,
    new_P1_U3960, new_P1_U3961, new_P1_U3962, new_P1_U3963, new_P1_U3964,
    new_P1_U3965, new_P1_U3966, new_P1_U3967, new_P1_U3968, new_P1_U3969,
    new_P1_U3970, new_P1_U3971, new_P1_U3972, new_P1_U3974, new_P1_U3975,
    new_P1_U3976, new_P1_U3977, new_P1_U3978, new_P1_U3979, new_P1_U3980,
    new_P1_U3981, new_P1_U3982, new_P1_U3983, new_P1_U3984, new_P1_U3985,
    new_P1_U3986, new_P1_U3987, new_P1_U3988, new_P1_U3989, new_P1_U3990,
    new_P1_U3991, new_P1_U3992, new_P1_U3993, new_P1_U3994, new_P1_U3995,
    new_P1_U3996, new_P1_U3997, new_P1_U3998, new_P1_U3999, new_P1_U4000,
    new_P1_U4001, new_P1_U4002, new_P1_U4003, new_P1_U4004, new_P1_U4005,
    new_P1_U4006, new_P1_U4007, new_P1_U4008, new_P1_U4009, new_P1_U4010,
    new_P1_U4011, new_P1_U4012, new_P1_U4013, new_P1_U4014, new_P1_U4015,
    new_P1_U4016, new_P1_U4017, new_P1_U4018, new_P1_U4019, new_P1_U4020,
    new_P1_U4021, new_P1_U4022, new_P1_U4023, new_P1_U4024, new_P1_U4025,
    new_P1_U4026, new_P1_U4027, new_P1_U4028, new_P1_U4029, new_P1_U4030,
    new_P1_U4031, new_P1_U4032, new_P1_U4033, new_P1_U4034, new_P1_U4035,
    new_P1_U4036, new_P1_U4037, new_P1_U4038, new_P1_U4039, new_P1_U4040,
    new_P1_U4041, new_P1_U4042, new_P1_U4043, new_P1_U4044, new_P1_U4045,
    new_P1_U4046, new_P1_U4047, new_P1_U4048, new_P1_U4049, new_P1_U4050,
    new_P1_U4051, new_P1_U4052, new_P1_U4053, new_P1_U4054, new_P1_U4055,
    new_P1_U4056, new_P1_U4057, new_P1_U4058, new_P1_U4059, new_P1_U4060,
    new_P1_U4061, new_P1_U4062, new_P1_U4063, new_P1_U4064, new_P1_U4065,
    new_P1_U4066, new_P1_U4067, new_P1_U4068, new_P1_U4069, new_P1_U4070,
    new_P1_U4071, new_P1_U4072, new_P1_U4073, new_P1_U4074, new_P1_U4075,
    new_P1_U4076, new_P1_U4077, new_P1_U4078, new_P1_U4079, new_P1_U4080,
    new_P1_U4081, new_P1_U4082, new_P1_U4083, new_P1_U4084, new_P1_U4085,
    new_P1_U4086, new_P1_U4087, new_P1_U4088, new_P1_U4089, new_P1_U4090,
    new_P1_U4091, new_P1_U4092, new_P1_U4093, new_P1_U4094, new_P1_U4095,
    new_P1_U4096, new_P1_U4097, new_P1_U4098, new_P1_U4099, new_P1_U4100,
    new_P1_U4101, new_P1_U4102, new_P1_U4103, new_P1_U4104, new_P1_U4105,
    new_P1_U4106, new_P1_U4107, new_P1_U4108, new_P1_U4109, new_P1_U4110,
    new_P1_U4111, new_P1_U4112, new_P1_U4113, new_P1_U4114, new_P1_U4115,
    new_P1_U4116, new_P1_U4117, new_P1_U4118, new_P1_U4119, new_P1_U4120,
    new_P1_U4121, new_P1_U4122, new_P1_U4123, new_P1_U4124, new_P1_U4125,
    new_P1_U4126, new_P1_U4127, new_P1_U4128, new_P1_U4129, new_P1_U4130,
    new_P1_U4131, new_P1_U4132, new_P1_U4133, new_P1_U4134, new_P1_U4135,
    new_P1_U4136, new_P1_U4137, new_P1_U4138, new_P1_U4139, new_P1_U4140,
    new_P1_U4141, new_P1_U4142, new_P1_U4143, new_P1_U4144, new_P1_U4145,
    new_P1_U4146, new_P1_U4147, new_P1_U4148, new_P1_U4149, new_P1_U4150,
    new_P1_U4151, new_P1_U4152, new_P1_U4153, new_P1_U4154, new_P1_U4155,
    new_P1_U4156, new_P1_U4157, new_P1_U4158, new_P1_U4159, new_P1_U4160,
    new_P1_U4161, new_P1_U4162, new_P1_U4163, new_P1_U4164, new_P1_U4165,
    new_P1_U4166, new_P1_U4167, new_P1_U4168, new_P1_U4169, new_P1_U4170,
    new_P1_U4171, new_P1_U4172, new_P1_U4173, new_P1_U4174, new_P1_U4175,
    new_P1_U4176, new_P1_U4177, new_P1_U4178, new_P1_U4179, new_P1_U4180,
    new_P1_U4181, new_P1_U4182, new_P1_U4183, new_P1_U4184, new_P1_U4185,
    new_P1_U4186, new_P1_U4187, new_P1_U4188, new_P1_U4189, new_P1_U4190,
    new_P1_U4191, new_P1_U4192, new_P1_U4193, new_P1_U4194, new_P1_U4195,
    new_P1_U4196, new_P1_U4197, new_P1_U4198, new_P1_U4199, new_P1_U4200,
    new_P1_U4201, new_P1_U4202, new_P1_U4203, new_P1_U4204, new_P1_U4205,
    new_P1_U4206, new_P1_U4207, new_P1_U4208, new_P1_U4209, new_P1_U4210,
    new_P1_U4211, new_P1_U4212, new_P1_U4213, new_P1_U4214, new_P1_U4215,
    new_P1_U4216, new_P1_U4217, new_P1_U4218, new_P1_U4219, new_P1_U4220,
    new_P1_U4221, new_P1_U4222, new_P1_U4223, new_P1_U4224, new_P1_U4225,
    new_P1_U4226, new_P1_U4227, new_P1_U4228, new_P1_U4229, new_P1_U4230,
    new_P1_U4231, new_P1_U4232, new_P1_U4233, new_P1_U4234, new_P1_U4235,
    new_P1_U4236, new_P1_U4237, new_P1_U4238, new_P1_U4239, new_P1_U4240,
    new_P1_U4241, new_P1_U4242, new_P1_U4243, new_P1_U4244, new_P1_U4245,
    new_P1_U4246, new_P1_U4247, new_P1_U4248, new_P1_U4249, new_P1_U4250,
    new_P1_U4251, new_P1_U4252, new_P1_U4253, new_P1_U4254, new_P1_U4255,
    new_P1_U4256, new_P1_U4257, new_P1_U4258, new_P1_U4259, new_P1_U4260,
    new_P1_U4261, new_P1_U4262, new_P1_U4263, new_P1_U4264, new_P1_U4265,
    new_P1_U4266, new_P1_U4267, new_P1_U4268, new_P1_U4269, new_P1_U4270,
    new_P1_U4271, new_P1_U4272, new_P1_U4273, new_P1_U4274, new_P1_U4275,
    new_P1_U4276, new_P1_U4277, new_P1_U4278, new_P1_U4279, new_P1_U4280,
    new_P1_U4281, new_P1_U4282, new_P1_U4283, new_P1_U4284, new_P1_U4285,
    new_P1_U4286, new_P1_U4287, new_P1_U4288, new_P1_U4289, new_P1_U4290,
    new_P1_U4291, new_P1_U4292, new_P1_U4293, new_P1_U4294, new_P1_U4295,
    new_P1_U4296, new_P1_U4297, new_P1_U4298, new_P1_U4299, new_P1_U4300,
    new_P1_U4301, new_P1_U4302, new_P1_U4303, new_P1_U4304, new_P1_U4305,
    new_P1_U4306, new_P1_U4307, new_P1_U4308, new_P1_U4309, new_P1_U4310,
    new_P1_U4311, new_P1_U4312, new_P1_U4313, new_P1_U4314, new_P1_U4315,
    new_P1_U4316, new_P1_U4317, new_P1_U4318, new_P1_U4319, new_P1_U4320,
    new_P1_U4321, new_P1_U4322, new_P1_U4323, new_P1_U4324, new_P1_U4325,
    new_P1_U4326, new_P1_U4327, new_P1_U4328, new_P1_U4329, new_P1_U4330,
    new_P1_U4331, new_P1_U4332, new_P1_U4333, new_P1_U4334, new_P1_U4335,
    new_P1_U4336, new_P1_U4337, new_P1_U4338, new_P1_U4339, new_P1_U4340,
    new_P1_U4341, new_P1_U4342, new_P1_U4343, new_P1_U4344, new_P1_U4345,
    new_P1_U4346, new_P1_U4347, new_P1_U4348, new_P1_U4349, new_P1_U4350,
    new_P1_U4351, new_P1_U4352, new_P1_U4353, new_P1_U4354, new_P1_U4355,
    new_P1_U4356, new_P1_U4357, new_P1_U4358, new_P1_U4359, new_P1_U4360,
    new_P1_U4361, new_P1_U4362, new_P1_U4363, new_P1_U4364, new_P1_U4365,
    new_P1_U4366, new_P1_U4367, new_P1_U4368, new_P1_U4369, new_P1_U4370,
    new_P1_U4371, new_P1_U4372, new_P1_U4373, new_P1_U4374, new_P1_U4375,
    new_P1_U4376, new_P1_U4377, new_P1_U4378, new_P1_U4379, new_P1_U4380,
    new_P1_U4381, new_P1_U4382, new_P1_U4383, new_P1_U4384, new_P1_U4385,
    new_P1_U4386, new_P1_U4387, new_P1_U4388, new_P1_U4389, new_P1_U4390,
    new_P1_U4391, new_P1_U4392, new_P1_U4393, new_P1_U4394, new_P1_U4395,
    new_P1_U4396, new_P1_U4397, new_P1_U4398, new_P1_U4399, new_P1_U4400,
    new_P1_U4401, new_P1_U4402, new_P1_U4403, new_P1_U4404, new_P1_U4405,
    new_P1_U4406, new_P1_U4407, new_P1_U4408, new_P1_U4409, new_P1_U4410,
    new_P1_U4411, new_P1_U4412, new_P1_U4413, new_P1_U4414, new_P1_U4415,
    new_P1_U4416, new_P1_U4417, new_P1_U4418, new_P1_U4419, new_P1_U4420,
    new_P1_U4421, new_P1_U4422, new_P1_U4423, new_P1_U4424, new_P1_U4425,
    new_P1_U4426, new_P1_U4427, new_P1_U4428, new_P1_U4429, new_P1_U4430,
    new_P1_U4431, new_P1_U4432, new_P1_U4433, new_P1_U4434, new_P1_U4435,
    new_P1_U4436, new_P1_U4437, new_P1_U4438, new_P1_U4439, new_P1_U4440,
    new_P1_U4441, new_P1_U4442, new_P1_U4443, new_P1_U4444, new_P1_U4445,
    new_P1_U4446, new_P1_U4447, new_P1_U4448, new_P1_U4449, new_P1_U4450,
    new_P1_U4451, new_P1_U4452, new_P1_U4453, new_P1_U4454, new_P1_U4455,
    new_P1_U4456, new_P1_U4457, new_P1_U4458, new_P1_U4459, new_P1_U4460,
    new_P1_U4461, new_P1_U4462, new_P1_U4463, new_P1_U4464, new_P1_U4465,
    new_P1_U4466, new_P1_U4467, new_P1_U4468, new_P1_U4469, new_P1_U4470,
    new_P1_U4471, new_P1_U4472, new_P1_U4473, new_P1_U4474, new_P1_U4475,
    new_P1_U4476, new_P1_U4477, new_P1_U4478, new_P1_U4479, new_P1_U4480,
    new_P1_U4481, new_P1_U4482, new_P1_U4483, new_P1_U4484, new_P1_U4485,
    new_P1_U4486, new_P1_U4487, new_P1_U4488, new_P1_U4489, new_P1_U4490,
    new_P1_U4491, new_P1_U4492, new_P1_U4493, new_P1_U4494, new_P1_U4495,
    new_P1_U4496, new_P1_U4497, new_P1_U4498, new_P1_U4499, new_P1_U4500,
    new_P1_U4501, new_P1_U4502, new_P1_U4503, new_P1_U4504, new_P1_U4505,
    new_P1_U4506, new_P1_U4507, new_P1_U4508, new_P1_U4509, new_P1_U4510,
    new_P1_U4511, new_P1_U4512, new_P1_U4513, new_P1_U4514, new_P1_U4515,
    new_P1_U4516, new_P1_U4517, new_P1_U4518, new_P1_U4519, new_P1_U4520,
    new_P1_U4521, new_P1_U4522, new_P1_U4523, new_P1_U4524, new_P1_U4525,
    new_P1_U4526, new_P1_U4527, new_P1_U4528, new_P1_U4529, new_P1_U4530,
    new_P1_U4531, new_P1_U4532, new_P1_U4533, new_P1_U4534, new_P1_U4535,
    new_P1_U4536, new_P1_U4537, new_P1_U4538, new_P1_U4539, new_P1_U4540,
    new_P1_U4541, new_P1_U4542, new_P1_U4543, new_P1_U4544, new_P1_U4545,
    new_P1_U4546, new_P1_U4547, new_P1_U4548, new_P1_U4549, new_P1_U4550,
    new_P1_U4551, new_P1_U4552, new_P1_U4553, new_P1_U4554, new_P1_U4555,
    new_P1_U4556, new_P1_U4557, new_P1_U4558, new_P1_U4559, new_P1_U4560,
    new_P1_U4561, new_P1_U4562, new_P1_U4563, new_P1_U4564, new_P1_U4565,
    new_P1_U4566, new_P1_U4567, new_P1_U4568, new_P1_U4569, new_P1_U4570,
    new_P1_U4571, new_P1_U4572, new_P1_U4573, new_P1_U4574, new_P1_U4575,
    new_P1_U4576, new_P1_U4577, new_P1_U4578, new_P1_U4579, new_P1_U4580,
    new_P1_U4581, new_P1_U4582, new_P1_U4583, new_P1_U4584, new_P1_U4585,
    new_P1_U4586, new_P1_U4587, new_P1_U4588, new_P1_U4589, new_P1_U4590,
    new_P1_U4591, new_P1_U4592, new_P1_U4593, new_P1_U4594, new_P1_U4595,
    new_P1_U4596, new_P1_U4597, new_P1_U4598, new_P1_U4599, new_P1_U4600,
    new_P1_U4601, new_P1_U4602, new_P1_U4603, new_P1_U4604, new_P1_U4605,
    new_P1_U4606, new_P1_U4607, new_P1_U4608, new_P1_U4609, new_P1_U4610,
    new_P1_U4611, new_P1_U4612, new_P1_U4613, new_P1_U4614, new_P1_U4615,
    new_P1_U4616, new_P1_U4617, new_P1_U4618, new_P1_U4619, new_P1_U4620,
    new_P1_U4621, new_P1_U4622, new_P1_U4623, new_P1_U4624, new_P1_U4625,
    new_P1_U4626, new_P1_U4627, new_P1_U4628, new_P1_U4629, new_P1_U4630,
    new_P1_U4631, new_P1_U4632, new_P1_U4633, new_P1_U4634, new_P1_U4635,
    new_P1_U4636, new_P1_U4637, new_P1_U4638, new_P1_U4639, new_P1_U4640,
    new_P1_U4641, new_P1_U4642, new_P1_U4643, new_P1_U4644, new_P1_U4645,
    new_P1_U4646, new_P1_U4647, new_P1_U4648, new_P1_U4649, new_P1_U4650,
    new_P1_U4651, new_P1_U4652, new_P1_U4653, new_P1_U4654, new_P1_U4655,
    new_P1_U4656, new_P1_U4657, new_P1_U4658, new_P1_U4659, new_P1_U4660,
    new_P1_U4661, new_P1_U4662, new_P1_U4663, new_P1_U4664, new_P1_U4665,
    new_P1_U4666, new_P1_U4667, new_P1_U4668, new_P1_U4669, new_P1_U4670,
    new_P1_U4671, new_P1_U4672, new_P1_U4673, new_P1_U4674, new_P1_U4675,
    new_P1_U4676, new_P1_U4677, new_P1_U4678, new_P1_U4679, new_P1_U4680,
    new_P1_U4681, new_P1_U4682, new_P1_U4683, new_P1_U4684, new_P1_U4685,
    new_P1_U4686, new_P1_U4687, new_P1_U4688, new_P1_U4689, new_P1_U4690,
    new_P1_U4691, new_P1_U4692, new_P1_U4693, new_P1_U4694, new_P1_U4695,
    new_P1_U4696, new_P1_U4697, new_P1_U4698, new_P1_U4699, new_P1_U4700,
    new_P1_U4701, new_P1_U4702, new_P1_U4703, new_P1_U4704, new_P1_U4705,
    new_P1_U4706, new_P1_U4707, new_P1_U4708, new_P1_U4709, new_P1_U4710,
    new_P1_U4711, new_P1_U4712, new_P1_U4713, new_P1_U4714, new_P1_U4715,
    new_P1_U4716, new_P1_U4717, new_P1_U4718, new_P1_U4719, new_P1_U4720,
    new_P1_U4721, new_P1_U4722, new_P1_U4723, new_P1_U4724, new_P1_U4725,
    new_P1_U4726, new_P1_U4727, new_P1_U4728, new_P1_U4729, new_P1_U4730,
    new_P1_U4731, new_P1_U4732, new_P1_U4733, new_P1_U4734, new_P1_U4735,
    new_P1_U4736, new_P1_U4737, new_P1_U4738, new_P1_U4739, new_P1_U4740,
    new_P1_U4741, new_P1_U4742, new_P1_U4743, new_P1_U4744, new_P1_U4745,
    new_P1_U4746, new_P1_U4747, new_P1_U4748, new_P1_U4749, new_P1_U4750,
    new_P1_U4751, new_P1_U4752, new_P1_U4753, new_P1_U4754, new_P1_U4755,
    new_P1_U4756, new_P1_U4757, new_P1_U4758, new_P1_U4759, new_P1_U4760,
    new_P1_U4761, new_P1_U4762, new_P1_U4763, new_P1_U4764, new_P1_U4765,
    new_P1_U4766, new_P1_U4767, new_P1_U4768, new_P1_U4769, new_P1_U4770,
    new_P1_U4771, new_P1_U4772, new_P1_U4773, new_P1_U4774, new_P1_U4775,
    new_P1_U4776, new_P1_U4777, new_P1_U4778, new_P1_U4779, new_P1_U4780,
    new_P1_U4781, new_P1_U4782, new_P1_U4783, new_P1_U4784, new_P1_U4785,
    new_P1_U4786, new_P1_U4787, new_P1_U4788, new_P1_U4789, new_P1_U4790,
    new_P1_U4791, new_P1_U4792, new_P1_U4793, new_P1_U4794, new_P1_U4795,
    new_P1_U4796, new_P1_U4797, new_P1_U4798, new_P1_U4799, new_P1_U4800,
    new_P1_U4801, new_P1_U4802, new_P1_U4803, new_P1_U4804, new_P1_U4805,
    new_P1_U4806, new_P1_U4807, new_P1_U4808, new_P1_U4809, new_P1_U4810,
    new_P1_U4811, new_P1_U4812, new_P1_U4813, new_P1_U4814, new_P1_U4815,
    new_P1_U4816, new_P1_U4817, new_P1_U4818, new_P1_U4819, new_P1_U4820,
    new_P1_U4821, new_P1_U4822, new_P1_U4823, new_P1_U4824, new_P1_U4825,
    new_P1_U4826, new_P1_U4827, new_P1_U4828, new_P1_U4829, new_P1_U4830,
    new_P1_U4831, new_P1_U4832, new_P1_U4833, new_P1_U4834, new_P1_U4835,
    new_P1_U4836, new_P1_U4837, new_P1_U4838, new_P1_U4839, new_P1_U4840,
    new_P1_U4841, new_P1_U4842, new_P1_U4843, new_P1_U4844, new_P1_U4845,
    new_P1_U4846, new_P1_U4847, new_P1_U4848, new_P1_U4849, new_P1_U4850,
    new_P1_U4851, new_P1_U4852, new_P1_U4853, new_P1_U4854, new_P1_U4855,
    new_P1_U4856, new_P1_U4857, new_P1_U4858, new_P1_U4859, new_P1_U4860,
    new_P1_U4861, new_P1_U4862, new_P1_U4863, new_P1_U4864, new_P1_U4865,
    new_P1_U4866, new_P1_U4867, new_P1_U4868, new_P1_U4869, new_P1_U4870,
    new_P1_U4871, new_P1_U4872, new_P1_U4873, new_P1_U4874, new_P1_U4875,
    new_P1_U4876, new_P1_U4877, new_P1_U4878, new_P1_U4879, new_P1_U4880,
    new_P1_U4881, new_P1_U4882, new_P1_U4883, new_P1_U4884, new_P1_U4885,
    new_P1_U4886, new_P1_U4887, new_P1_U4888, new_P1_U4889, new_P1_U4890,
    new_P1_U4891, new_P1_U4892, new_P1_U4893, new_P1_U4894, new_P1_U4895,
    new_P1_U4896, new_P1_U4897, new_P1_U4898, new_P1_U4899, new_P1_U4900,
    new_P1_U4901, new_P1_U4902, new_P1_U4903, new_P1_U4904, new_P1_U4905,
    new_P1_U4906, new_P1_U4907, new_P1_U4908, new_P1_U4909, new_P1_U4910,
    new_P1_U4911, new_P1_U4912, new_P1_U4913, new_P1_U4914, new_P1_U4915,
    new_P1_U4916, new_P1_U4917, new_P1_U4918, new_P1_U4919, new_P1_U4920,
    new_P1_U4921, new_P1_U4922, new_P1_U4923, new_P1_U4924, new_P1_U4925,
    new_P1_U4926, new_P1_U4927, new_P1_U4928, new_P1_U4929, new_P1_U4930,
    new_P1_U4931, new_P1_U4932, new_P1_U4933, new_P1_U4934, new_P1_U4935,
    new_P1_U4936, new_P1_U4937, new_P1_U4938, new_P1_U4939, new_P1_U4940,
    new_P1_U4941, new_P1_U4942, new_P1_U4943, new_P1_U4944, new_P1_U4945,
    new_P1_U4946, new_P1_U4947, new_P1_U4948, new_P1_U4949, new_P1_U4950,
    new_P1_U4951, new_P1_U4952, new_P1_U4953, new_P1_U4954, new_P1_U4955,
    new_P1_U4956, new_P1_U4957, new_P1_U4958, new_P1_U4959, new_P1_U4960,
    new_P1_U4961, new_P1_U4962, new_P1_U4963, new_P1_U4964, new_P1_U4965,
    new_P1_U4966, new_P1_U4967, new_P1_U4968, new_P1_U4969, new_P1_U4970,
    new_P1_U4971, new_P1_U4972, new_P1_U4973, new_P1_U4974, new_P1_U4975,
    new_P1_U4976, new_P1_U4977, new_P1_U4978, new_P1_U4979, new_P1_U4980,
    new_P1_U4981, new_P1_U4982, new_P1_U4983, new_P1_U4984, new_P1_U4985,
    new_P1_U4986, new_P1_U4987, new_P1_U4988, new_P1_U4989, new_P1_U4990,
    new_P1_U4991, new_P1_U4992, new_P1_U4993, new_P1_U4994, new_P1_U4995,
    new_P1_U4996, new_P1_U4997, new_P1_U4998, new_P1_U4999, new_P1_U5000,
    new_P1_U5001, new_P1_U5002, new_P1_U5003, new_P1_U5004, new_P1_U5005,
    new_P1_U5006, new_P1_U5007, new_P1_U5008, new_P1_U5009, new_P1_U5010,
    new_P1_U5011, new_P1_U5012, new_P1_U5013, new_P1_U5014, new_P1_U5015,
    new_P1_U5016, new_P1_U5017, new_P1_U5018, new_P1_U5019, new_P1_U5020,
    new_P1_U5021, new_P1_U5022, new_P1_U5023, new_P1_U5024, new_P1_U5025,
    new_P1_U5026, new_P1_U5027, new_P1_U5028, new_P1_U5029, new_P1_U5030,
    new_P1_U5031, new_P1_U5032, new_P1_U5033, new_P1_U5034, new_P1_U5035,
    new_P1_U5036, new_P1_U5037, new_P1_U5038, new_P1_U5039, new_P1_U5040,
    new_P1_U5041, new_P1_U5042, new_P1_U5043, new_P1_U5044, new_P1_U5045,
    new_P1_U5046, new_P1_U5047, new_P1_U5048, new_P1_U5049, new_P1_U5050,
    new_P1_U5051, new_P1_U5052, new_P1_U5053, new_P1_U5054, new_P1_U5055,
    new_P1_U5056, new_P1_U5057, new_P1_U5058, new_P1_U5059, new_P1_U5060,
    new_P1_U5061, new_P1_U5062, new_P1_U5063, new_P1_U5064, new_P1_U5065,
    new_P1_U5066, new_P1_U5067, new_P1_U5068, new_P1_U5069, new_P1_U5070,
    new_P1_U5071, new_P1_U5072, new_P1_U5073, new_P1_U5074, new_P1_U5075,
    new_P1_U5076, new_P1_U5077, new_P1_U5078, new_P1_U5079, new_P1_U5080,
    new_P1_U5081, new_P1_U5082, new_P1_U5083, new_P1_U5084, new_P1_U5085,
    new_P1_U5086, new_P1_U5087, new_P1_U5088, new_P1_U5089, new_P1_U5090,
    new_P1_U5091, new_P1_U5092, new_P1_U5093, new_P1_U5094, new_P1_U5095,
    new_P1_U5096, new_P1_U5097, new_P1_U5098, new_P1_U5099, new_P1_U5100,
    new_P1_U5101, new_P1_U5102, new_P1_U5103, new_P1_U5104, new_P1_U5105,
    new_P1_U5106, new_P1_U5107, new_P1_U5108, new_P1_U5109, new_P1_U5110,
    new_P1_U5111, new_P1_U5112, new_P1_U5113, new_P1_U5114, new_P1_U5115,
    new_P1_U5116, new_P1_U5117, new_P1_U5118, new_P1_U5119, new_P1_U5120,
    new_P1_U5121, new_P1_U5122, new_P1_U5123, new_P1_U5124, new_P1_U5125,
    new_P1_U5126, new_P1_U5127, new_P1_U5128, new_P1_U5129, new_P1_U5130,
    new_P1_U5131, new_P1_U5132, new_P1_U5133, new_P1_U5134, new_P1_U5135,
    new_P1_U5136, new_P1_U5137, new_P1_U5138, new_P1_U5139, new_P1_U5140,
    new_P1_U5141, new_P1_U5142, new_P1_U5143, new_P1_U5144, new_P1_U5145,
    new_P1_U5146, new_P1_U5147, new_P1_U5148, new_P1_U5149, new_P1_U5150,
    new_P1_U5151, new_P1_U5152, new_P1_U5153, new_P1_U5154, new_P1_U5155,
    new_P1_U5156, new_P1_U5157, new_P1_U5158, new_P1_U5159, new_P1_U5160,
    new_P1_U5161, new_P1_U5162, new_P1_U5163, new_P1_U5164, new_P1_U5165,
    new_P1_U5166, new_P1_U5167, new_P1_U5168, new_P1_U5169, new_P1_U5170,
    new_P1_U5171, new_P1_U5172, new_P1_U5173, new_P1_U5174, new_P1_U5175,
    new_P1_U5176, new_P1_U5177, new_P1_U5178, new_P1_U5179, new_P1_U5180,
    new_P1_U5181, new_P1_U5182, new_P1_U5183, new_P1_U5184, new_P1_U5185,
    new_P1_U5186, new_P1_U5187, new_P1_U5188, new_P1_U5189, new_P1_U5190,
    new_P1_U5191, new_P1_U5192, new_P1_U5193, new_P1_U5194, new_P1_U5195,
    new_P1_U5196, new_P1_U5197, new_P1_U5198, new_P1_U5199, new_P1_U5200,
    new_P1_U5201, new_P1_U5202, new_P1_U5203, new_P1_U5204, new_P1_U5205,
    new_P1_U5206, new_P1_U5207, new_P1_U5208, new_P1_U5209, new_P1_U5210,
    new_P1_U5211, new_P1_U5212, new_P1_U5213, new_P1_U5214, new_P1_U5215,
    new_P1_U5216, new_P1_U5217, new_P1_U5218, new_P1_U5219, new_P1_U5220,
    new_P1_U5221, new_P1_U5222, new_P1_U5223, new_P1_U5224, new_P1_U5225,
    new_P1_U5226, new_P1_U5227, new_P1_U5228, new_P1_U5229, new_P1_U5230,
    new_P1_U5231, new_P1_U5232, new_P1_U5233, new_P1_U5234, new_P1_U5235,
    new_P1_U5236, new_P1_U5237, new_P1_U5238, new_P1_U5239, new_P1_U5240,
    new_P1_U5241, new_P1_U5242, new_P1_U5243, new_P1_U5244, new_P1_U5245,
    new_P1_U5246, new_P1_U5247, new_P1_U5248, new_P1_U5249, new_P1_U5250,
    new_P1_U5251, new_P1_U5252, new_P1_U5253, new_P1_U5254, new_P1_U5255,
    new_P1_U5256, new_P1_U5257, new_P1_U5258, new_P1_U5259, new_P1_U5260,
    new_P1_U5261, new_P1_U5262, new_P1_U5263, new_P1_U5264, new_P1_U5265,
    new_P1_U5266, new_P1_U5267, new_P1_U5268, new_P1_U5269, new_P1_U5270,
    new_P1_U5271, new_P1_U5272, new_P1_U5273, new_P1_U5274, new_P1_U5275,
    new_P1_U5276, new_P1_U5277, new_P1_U5278, new_P1_U5279, new_P1_U5280,
    new_P1_U5281, new_P1_U5282, new_P1_U5283, new_P1_U5284, new_P1_U5285,
    new_P1_U5286, new_P1_U5287, new_P1_U5288, new_P1_U5289, new_P1_U5290,
    new_P1_U5291, new_P1_U5292, new_P1_U5293, new_P1_U5294, new_P1_U5295,
    new_P1_U5296, new_P1_U5297, new_P1_U5298, new_P1_U5299, new_P1_U5300,
    new_P1_U5301, new_P1_U5302, new_P1_U5303, new_P1_U5304, new_P1_U5305,
    new_P1_U5306, new_P1_U5307, new_P1_U5308, new_P1_U5309, new_P1_U5310,
    new_P1_U5311, new_P1_U5312, new_P1_U5313, new_P1_U5314, new_P1_U5315,
    new_P1_U5316, new_P1_U5317, new_P1_U5318, new_P1_U5319, new_P1_U5320,
    new_P1_U5321, new_P1_U5322, new_P1_U5323, new_P1_U5324, new_P1_U5325,
    new_P1_U5326, new_P1_U5327, new_P1_U5328, new_P1_U5329, new_P1_U5330,
    new_P1_U5331, new_P1_U5332, new_P1_U5333, new_P1_U5334, new_P1_U5335,
    new_P1_U5336, new_P1_U5337, new_P1_U5338, new_P1_U5339, new_P1_U5340,
    new_P1_U5341, new_P1_U5342, new_P1_U5343, new_P1_U5344, new_P1_U5345,
    new_P1_U5346, new_P1_U5347, new_P1_U5348, new_P1_U5349, new_P1_U5350,
    new_P1_U5351, new_P1_U5352, new_P1_U5353, new_P1_U5354, new_P1_U5355,
    new_P1_U5356, new_P1_U5357, new_P1_U5358, new_P1_U5359, new_P1_U5360,
    new_P1_U5361, new_P1_U5362, new_P1_U5363, new_P1_U5364, new_P1_U5365,
    new_P1_U5366, new_P1_U5367, new_P1_U5368, new_P1_U5369, new_P1_U5370,
    new_P1_U5371, new_P1_U5372, new_P1_U5373, new_P1_U5374, new_P1_U5375,
    new_P1_U5376, new_P1_U5377, new_P1_U5378, new_P1_U5379, new_P1_U5380,
    new_P1_U5381, new_P1_U5382, new_P1_U5383, new_P1_U5384, new_P1_U5385,
    new_P1_U5386, new_P1_U5387, new_P1_U5388, new_P1_U5389, new_P1_U5390,
    new_P1_U5391, new_P1_U5392, new_P1_U5393, new_P1_U5394, new_P1_U5395,
    new_P1_U5396, new_P1_U5397, new_P1_U5398, new_P1_U5399, new_P1_U5400,
    new_P1_U5401, new_P1_U5402, new_P1_U5403, new_P1_U5404, new_P1_U5405,
    new_P1_U5406, new_P1_U5407, new_P1_U5408, new_P1_U5409, new_P1_U5410,
    new_P1_U5411, new_P1_U5412, new_P1_U5413, new_P1_U5414, new_P1_U5415,
    new_P1_U5416, new_P1_U5417, new_P1_U5418, new_P1_U5419, new_P1_U5420,
    new_P1_U5421, new_P1_U5422, new_P1_U5423, new_P1_U5424, new_P1_U5425,
    new_P1_U5426, new_P1_U5427, new_P1_U5428, new_P1_U5429, new_P1_U5430,
    new_P1_U5431, new_P1_U5432, new_P1_U5433, new_P1_U5434, new_P1_U5435,
    new_P1_U5436, new_P1_U5437, new_P1_U5438, new_P1_U5439, new_P1_U5440,
    new_P1_U5441, new_P1_U5442, new_P1_U5443, new_P1_U5444, new_P1_U5445,
    new_P1_U5446, new_P1_U5447, new_P1_U5448, new_P1_U5449, new_P1_U5450,
    new_P1_U5451, new_P1_U5452, new_P1_U5453, new_P1_U5454, new_P1_U5455,
    new_P1_U5456, new_P1_U5457, new_P1_U5458, new_P1_U5459, new_P1_U5460,
    new_P1_U5461, new_P1_U5462, new_P1_U5463, new_P1_U5464, new_P1_U5465,
    new_P1_U5466, new_P1_U5467, new_P1_U5468, new_P1_U5469, new_P1_U5470,
    new_P1_U5471, new_P1_U5472, new_P1_U5473, new_P1_U5474, new_P1_U5475,
    new_P1_U5476, new_P1_U5477, new_P1_U5478, new_P1_U5479, new_P1_U5480,
    new_P1_U5481, new_P1_U5482, new_P1_U5483, new_P1_U5484, new_P1_U5485,
    new_P1_U5486, new_P1_U5487, new_P1_U5488, new_P1_U5489, new_P1_U5490,
    new_P1_U5491, new_P1_U5492, new_P1_U5493, new_P1_U5494, new_P1_U5495,
    new_P1_U5496, new_P1_U5497, new_P1_U5498, new_P1_U5499, new_P1_U5500,
    new_P1_U5501, new_P1_U5502, new_P1_U5503, new_P1_U5504, new_P1_U5505,
    new_P1_U5506, new_P1_U5507, new_P1_U5508, new_P1_U5509, new_P1_U5510,
    new_P1_U5511, new_P1_U5512, new_P1_U5513, new_P1_U5514, new_P1_U5515,
    new_P1_U5516, new_P1_U5517, new_P1_U5518, new_P1_U5519, new_P1_U5520,
    new_P1_U5521, new_P1_U5522, new_P1_U5523, new_P1_U5524, new_P1_U5525,
    new_P1_U5526, new_P1_U5527, new_P1_U5528, new_P1_U5529, new_P1_U5530,
    new_P1_U5531, new_P1_U5532, new_P1_U5533, new_P1_U5534, new_P1_U5535,
    new_P1_U5536, new_P1_U5537, new_P1_U5538, new_P1_U5539, new_P1_U5540,
    new_P1_U5541, new_P1_U5542, new_P1_U5543, new_P1_U5544, new_P1_U5545,
    new_P1_U5546, new_P1_U5547, new_P1_U5548, new_P1_U5549, new_P1_U5550,
    new_P1_U5551, new_P1_U5552, new_P1_U5553, new_P1_U5554, new_P1_U5555,
    new_P1_U5556, new_P1_U5557, new_P1_U5558, new_P1_U5559, new_P1_U5560,
    new_P1_U5561, new_P1_U5562, new_P1_U5563, new_P1_U5564, new_P1_U5565,
    new_P1_U5566, new_P1_U5567, new_P1_U5568, new_P1_U5569, new_P1_U5570,
    new_P1_U5571, new_P1_U5572, new_P1_U5573, new_P1_U5574, new_P1_U5575,
    new_P1_U5576, new_P1_U5577, new_P1_U5578, new_P1_U5579, new_P1_U5580,
    new_P1_U5581, new_P1_U5582, new_P1_U5583, new_P1_U5584, new_P1_U5585,
    new_P1_U5586, new_P1_U5587, new_P1_U5588, new_P1_U5589, new_P1_U5590,
    new_P1_U5591, new_P1_U5592, new_P1_U5593, new_P1_U5594, new_P1_U5595,
    new_P1_U5596, new_P1_U5597, new_P1_U5598, new_P1_U5599, new_P1_U5600,
    new_P1_U5601, new_P1_U5602, new_P1_U5603, new_P1_U5604, new_P1_U5605,
    new_P1_U5606, new_P1_U5607, new_P1_U5608, new_P1_U5609, new_P1_U5610,
    new_P1_U5611, new_P1_U5612, new_P1_U5613, new_P1_U5614, new_P1_U5615,
    new_P1_U5616, new_P1_U5617, new_P1_U5618, new_P1_U5619, new_P1_U5620,
    new_P1_U5621, new_P1_U5622, new_P1_U5623, new_P1_U5624, new_P1_U5625,
    new_P1_U5626, new_P1_U5627, new_P1_U5628, new_P1_U5629, new_P1_U5630,
    new_P1_U5631, new_P1_U5632, new_P1_U5633, new_P1_U5634, new_P1_U5635,
    new_P1_U5636, new_P1_U5637, new_P1_U5638, new_P1_U5639, new_P1_U5640,
    new_P1_U5641, new_P1_U5642, new_P1_U5643, new_P1_U5644, new_P1_U5645,
    new_P1_U5646, new_P1_U5647, new_P1_U5648, new_P1_U5649, new_P1_U5650,
    new_P1_U5651, new_P1_U5652, new_P1_U5653, new_P1_U5654, new_P1_U5655,
    new_P1_U5656, new_P1_U5657, new_P1_U5658, new_P1_U5659, new_P1_U5660,
    new_P1_U5661, new_P1_U5662, new_P1_U5663, new_P1_U5664, new_P1_U5665,
    new_P1_U5666, new_P1_U5667, new_P1_U5668, new_P1_U5669, new_P1_U5670,
    new_P1_U5671, new_P1_U5672, new_P1_U5673, new_P1_U5674, new_P1_U5675,
    new_P1_U5676, new_P1_U5677, new_P1_U5678, new_P1_U5679, new_P1_U5680,
    new_P1_U5681, new_P1_U5682, new_P1_U5683, new_P1_U5684, new_P1_U5685,
    new_P1_U5686, new_P1_U5687, new_P1_U5688, new_P1_U5689, new_P1_U5690,
    new_P1_U5691, new_P1_U5692, new_P1_U5693, new_P1_U5694, new_P1_U5695,
    new_P1_U5696, new_P1_U5697, new_P1_U5698, new_P1_U5699, new_P1_U5700,
    new_P1_U5701, new_P1_U5702, new_P1_U5703, new_P1_U5704, new_P1_U5705,
    new_P1_U5706, new_P1_U5707, new_P1_U5708, new_P1_U5709, new_P1_U5710,
    new_P1_U5711, new_P1_U5712, new_P1_U5713, new_P1_U5714, new_P1_U5715,
    new_P1_U5716, new_P1_U5717, new_P1_U5718, new_P1_U5719, new_P1_U5720,
    new_P1_U5721, new_P1_U5722, new_P1_U5723, new_P1_U5724, new_P1_U5725,
    new_P1_U5726, new_P1_U5727, new_P1_U5728, new_P1_U5729, new_P1_U5730,
    new_P1_U5731, new_P1_U5732, new_P1_U5733, new_P1_U5734, new_P1_U5735,
    new_P1_U5736, new_P1_U5737, new_P1_U5738, new_P1_U5739, new_P1_U5740,
    new_P1_U5741, new_P1_U5742, new_P1_U5743, new_P1_U5744, new_P1_U5745,
    new_P1_U5746, new_P1_U5747, new_P1_U5748, new_P1_U5749, new_P1_U5750,
    new_P1_U5751, new_P1_U5752, new_P1_U5753, new_P1_U5754, new_P1_U5755,
    new_P1_U5756, new_P1_U5757, new_P1_U5758, new_P1_U5759, new_P1_U5760,
    new_P1_U5761, new_P1_U5762, new_P1_U5763, new_P1_U5764, new_P1_U5765,
    new_P1_U5766, new_P1_U5767, new_P1_U5768, new_P1_U5769, new_P1_U5770,
    new_P1_U5771, new_P1_U5772, new_P1_U5773, new_P1_U5774, new_P1_U5775,
    new_P1_U5776, new_P1_U5777, new_P1_U5778, new_P1_U5779, new_P1_U5780,
    new_P1_U5781, new_P1_U5782, new_P1_U5783, new_P1_U5784, new_P1_U5785,
    new_P1_U5786, new_P1_U5787, new_P1_U5788, new_P1_U5789, new_P1_U5790,
    new_P1_U5791, new_P1_U5792, new_P1_U5793, new_P1_U5794, new_P1_U5795,
    new_P1_U5796, new_P1_U5797, new_P1_U5798, new_P1_U5799, new_P1_U5800,
    new_P1_U5801, new_P1_U5802, new_P1_U5803, new_P1_U5804, new_P1_U5805,
    new_P1_U5806, new_P1_U5807, new_P1_U5808, new_P1_U5809, new_P1_U5810,
    new_P1_U5811, new_P1_U5812, new_P1_U5813, new_P1_U5814, new_P1_U5815,
    new_P1_U5816, new_P1_U5817, new_P1_U5818, new_P1_U5819, new_P1_U5820,
    new_P1_U5821, new_P1_U5822, new_P1_U5823, new_P1_U5824, new_P1_U5825,
    new_P1_U5826, new_P1_U5827, new_P1_U5828, new_P1_U5829, new_P1_U5830,
    new_P1_U5831, new_P1_U5832, new_P1_U5833, new_P1_U5834, new_P1_U5835,
    new_P1_U5836, new_P1_U5837, new_P1_U5838, new_P1_U5839, new_P1_U5840,
    new_P1_U5841, new_P1_U5842, new_P1_U5843, new_P1_U5844, new_P1_U5845,
    new_P1_U5846, new_P1_U5847, new_P1_U5848, new_P1_U5849, new_P1_U5850,
    new_P1_U5851, new_P1_U5852, new_P1_U5853, new_P1_U5854, new_P1_U5855,
    new_P1_U5856, new_P1_U5857, new_P1_U5858, new_P1_U5859, new_P1_U5860,
    new_P1_U5861, new_P1_U5862, new_P1_U5863, new_P1_U5864, new_P1_U5865,
    new_P1_U5866, new_P1_U5867, new_P1_U5868, new_P1_U5869, new_P1_U5870,
    new_P1_U5871, new_P1_U5872, new_P1_U5873, new_P1_U5874, new_P1_U5875,
    new_P1_U5876, new_P1_U5877, new_P1_U5878, new_P1_U5879, new_P1_U5880,
    new_P1_U5881, new_P1_U5882, new_P1_U5883, new_P1_U5884, new_P1_U5885,
    new_P1_U5886, new_P1_U5887, new_P1_U5888, new_P1_U5889, new_P1_U5890,
    new_P1_U5891, new_P1_U5892, new_P1_U5893, new_P1_U5894, new_P1_U5895,
    new_P1_U5896, new_P1_U5897, new_P1_U5898, new_P1_U5899, new_P1_U5900,
    new_P1_U5901, new_P1_U5902, new_P1_U5903, new_P1_U5904, new_P1_U5905,
    new_P1_U5906, new_P1_U5907, new_P1_U5908, new_P1_U5909, new_P1_U5910,
    new_P1_U5911, new_P1_U5912, new_P1_U5913, new_P1_U5914, new_P1_U5915,
    new_P1_U5916, new_P1_U5917, new_P1_U5918, new_P1_U5919, new_P1_U5920,
    new_P1_U5921, new_P1_U5922, new_P1_U5923, new_P1_U5924, new_P1_U5925,
    new_P1_U5926, new_P1_U5927, new_P1_U5928, new_P1_U5929, new_P1_U5930,
    new_P1_U5931, new_P1_U5932, new_P1_U5933, new_P1_U5934, new_P1_U5935,
    new_P1_U5936, new_P1_U5937, new_P1_U5938, new_P1_U5939, new_P1_U5940,
    new_P1_U5941, new_P1_U5942, new_P1_U5943, new_P1_U5944, new_P1_U5945,
    new_P1_U5946, new_P1_U5947, new_P1_U5948, new_P1_U5949, new_P1_U5950,
    new_P1_U5951, new_P1_U5952, new_P1_U5953, new_P1_U5954, new_P1_U5955,
    new_P1_U5956, new_P1_U5957, new_P1_U5958, new_P1_U5959, new_P1_U5960,
    new_P1_U5961, new_P1_U5962, new_P1_U5963, new_P1_U5964, new_P1_U5965,
    new_P1_U5966, new_P1_U5967, new_P1_U5968, new_P1_U5969, new_P1_U5970,
    new_P1_U5971, new_P1_U5972, new_P1_U5973, new_P1_U5974, new_P1_U5975,
    new_P1_U5976, new_P1_U5977, new_P1_U5978, new_P1_U5979, new_P1_U5980,
    new_P1_U5981, new_P1_U5982, new_P1_U5983, new_P1_U5984, new_P1_U5985,
    new_P1_U5986, new_P1_U5987, new_P1_U5988, new_P1_U5989, new_P1_U5990,
    new_P1_U5991, new_P1_U5992, new_P1_U5993, new_P1_U5994, new_P1_U5995,
    new_P1_U5996, new_P1_U5997, new_P1_U5998, new_P1_U5999, new_P1_U6000,
    new_P1_U6001, new_P1_U6002, new_P1_U6003, new_P1_U6004, new_P1_U6005,
    new_P1_U6006, new_P1_U6007, new_P1_U6008, new_P1_U6009, new_P1_U6010,
    new_P1_U6011, new_P1_U6012, new_P1_U6013, new_P1_U6014, new_P1_U6015,
    new_P1_U6016, new_P1_U6017, new_P1_U6018, new_P1_U6019, new_P1_U6020,
    new_P1_U6021, new_P1_U6022, new_P1_U6023, new_P1_U6024, new_P1_U6025,
    new_P1_U6026, new_P1_U6027, new_P1_U6028, new_P1_U6029, new_P1_U6030,
    new_P1_U6031, new_P1_U6032, new_P1_U6033, new_P1_U6034, new_P1_U6035,
    new_P1_U6036, new_P1_U6037, new_P1_U6038, new_P1_U6039, new_P1_U6040,
    new_P1_U6041, new_P1_U6042, new_P1_U6043, new_P1_U6044, new_P1_U6045,
    new_P1_U6046, new_P1_U6047, new_P1_U6048, new_P1_U6049, new_P1_U6050,
    new_P1_U6051, new_P1_U6052, new_P1_U6053, new_P1_U6054, new_P1_U6055,
    new_P1_U6056, new_P1_U6057, new_P1_U6058, new_P1_U6059, new_P1_U6060,
    new_P1_U6061, new_P1_U6062, new_P1_U6063, new_P1_U6064, new_P1_U6065,
    new_P1_U6066, new_P1_U6067, new_P1_U6068, new_P1_U6069, new_P1_U6070,
    new_P1_U6071, new_P1_U6072, new_P1_U6073, new_P1_U6074, new_P1_U6075,
    new_P1_U6076, new_P1_U6077, new_P1_U6078, new_P1_U6079, new_P1_U6080,
    new_P1_U6081, new_P1_U6082, new_P1_U6083, new_P1_U6084, new_P1_U6085,
    new_P1_U6086, new_P1_U6087, new_P1_U6088, new_P1_U6089, new_P1_U6090,
    new_P1_U6091, new_P1_U6092, new_P1_U6093, new_P1_U6094, new_P1_U6095,
    new_P1_U6096, new_P1_U6097, new_P1_U6098, new_P1_U6099, new_P1_U6100,
    new_P1_U6101, new_P1_U6102, new_P1_U6103, new_P1_U6104, new_P1_U6105,
    new_P1_U6106, new_P1_U6107, new_P1_U6108, new_P1_U6109, new_P1_U6110,
    new_P1_U6111, new_P1_U6112, new_P1_U6113, new_P1_U6114, new_P1_U6115,
    new_P1_U6116, new_P1_U6117, new_P1_U6118, new_P1_U6119, new_P1_U6120,
    new_P1_U6121, new_P1_U6122, new_P1_U6123, new_P1_U6124, new_P1_U6125,
    new_P1_U6126, new_P1_U6127, new_P1_U6128, new_P1_U6129, new_P1_U6130,
    new_P1_U6131, new_P1_U6132, new_P1_U6133, new_P1_U6134, new_P1_U6135,
    new_P1_U6136, new_P1_U6137, new_P1_U6138, new_P1_U6139, new_P1_U6140,
    new_P1_U6141, new_P1_U6142, new_P1_U6143, new_P1_U6144, new_P1_U6145,
    new_P1_U6146, new_P1_U6147, new_P1_U6148, new_P1_U6149, new_P1_U6150,
    new_P1_U6151, new_P1_U6152, new_P1_U6153, new_P1_U6154, new_P1_U6155,
    new_P1_U6156, new_P1_U6157, new_P1_U6158, new_P1_U6159, new_P1_U6160,
    new_P1_U6161, new_P1_U6162, new_P1_U6163, new_P1_U6164, new_P1_U6165,
    new_P1_U6166, new_P1_U6167, new_P1_U6168, new_P1_U6169, new_P1_U6170,
    new_P1_U6171, new_P1_U6172, new_P1_U6173, new_P1_U6174, new_P1_U6175,
    new_P1_U6176, new_P1_U6177, new_P1_U6178, new_P1_U6179, new_P1_U6180,
    new_P1_U6181, new_P1_U6182, new_P1_U6183, new_P1_U6184, new_P1_U6185,
    new_P1_U6186, new_P1_U6187, new_P1_U6188, new_P1_U6189, new_P1_U6190,
    new_P1_U6191, new_P1_U6192, new_P1_U6193, new_P1_U6194, new_P1_U6195,
    new_P1_U6196, new_P1_U6197, new_P1_U6198, new_P1_U6199, new_P1_U6200,
    new_P1_U6201, new_P1_U6202, new_P1_U6203, new_P1_U6204, new_P1_U6205,
    new_P1_U6206, new_P1_U6207, new_P1_U6208, new_P1_U6209, new_P1_U6210,
    new_P1_U6211, new_P1_U6212, new_P1_U6213, new_P1_U6214, new_P1_U6215,
    new_P1_U6216, new_P1_U6217, new_P1_U6218, new_P1_U6219, new_P1_U6220,
    new_P1_U6221, new_P1_U6222, new_P1_U6223, new_P1_U6224, new_P1_U6225,
    new_P1_U6226, new_P1_U6227, new_P1_U6228, new_P1_U6229, new_P1_U6230,
    new_P1_U6231, new_P1_U6232, new_P1_U6233, new_P1_U6234, new_P1_U6235,
    new_P1_U6236, new_P2_R1161_U489, new_P2_R1161_U488, new_P2_R1161_U487,
    new_P2_R1161_U486, new_P2_R1161_U485, new_P2_R1161_U484,
    new_P2_R1161_U483, new_P2_R1161_U482, new_P2_R1161_U481,
    new_P2_R1161_U480, new_P2_R1161_U479, new_P2_R1161_U478,
    new_P2_R1161_U477, new_P2_R1161_U476, new_P2_R1161_U475,
    new_P2_R1161_U474, new_P2_R1161_U473, new_P2_R1161_U472,
    new_P2_R1161_U471, new_P2_R1161_U470, new_P2_R1161_U469,
    new_P2_R1161_U468, new_P2_R1161_U467, new_P2_R1161_U466, new_P2_U3013,
    new_P2_U3014, new_P2_U3015, new_P2_U3016, new_P2_U3017, new_P2_U3018,
    new_P2_U3019, new_P2_U3020, new_P2_U3021, new_P2_U3022, new_P2_U3023,
    new_P2_U3024, new_P2_U3025, new_P2_U3026, new_P2_U3027, new_P2_U3028,
    new_P2_U3029, new_P2_U3030, new_P2_U3031, new_P2_U3032, new_P2_U3033,
    new_P2_U3034, new_P2_U3035, new_P2_U3036, new_P2_U3037, new_P2_U3038,
    new_P2_U3039, new_P2_U3040, new_P2_U3041, new_P2_U3042, new_P2_U3043,
    new_P2_U3044, new_P2_U3045, new_P2_U3046, new_P2_U3047, new_P2_U3048,
    new_P2_U3049, new_P2_U3050, new_P2_U3051, new_P2_U3052, new_P2_U3053,
    new_P2_U3054, new_P2_U3055, new_P2_U3056, new_P2_U3057, new_P2_U3058,
    new_P2_U3059, new_P2_U3060, new_P2_U3061, new_P2_U3062, new_P2_U3063,
    new_P2_U3064, new_P2_U3065, new_P2_U3066, new_P2_U3067, new_P2_U3068,
    new_P2_U3069, new_P2_U3070, new_P2_U3071, new_P2_U3072, new_P2_U3073,
    new_P2_U3074, new_P2_U3075, new_P2_U3076, new_P2_U3077, new_P2_U3078,
    new_P2_U3079, new_P2_U3080, new_P2_U3081, new_P2_U3082, new_P2_U3083,
    new_P2_U3084, new_P2_U3085, new_P2_U3086, new_P2_U3087, new_P2_U3088,
    new_P2_U3089, new_P2_U3090, new_P2_U3091, new_P2_U3092, new_P2_U3093,
    new_P2_U3094, new_P2_U3095, new_P2_U3096, new_P2_U3097, new_P2_U3098,
    new_P2_U3099, new_P2_U3100, new_P2_U3101, new_P2_U3102, new_P2_U3103,
    new_P2_U3104, new_P2_U3105, new_P2_U3106, new_P2_U3107, new_P2_U3108,
    new_P2_U3109, new_P2_U3110, new_P2_U3111, new_P2_U3112, new_P2_U3113,
    new_P2_U3114, new_P2_U3115, new_P2_U3116, new_P2_U3117, new_P2_U3118,
    new_P2_U3119, new_P2_U3120, new_P2_U3121, new_P2_U3122, new_P2_U3123,
    new_P2_U3124, new_P2_U3125, new_P2_U3126, new_P2_U3127, new_P2_U3128,
    new_P2_U3129, new_P2_U3130, new_P2_U3131, new_P2_U3132, new_P2_U3133,
    new_P2_U3134, new_P2_U3135, new_P2_U3136, new_P2_U3137, new_P2_U3138,
    new_P2_U3139, new_P2_U3140, new_P2_U3141, new_P2_U3142, new_P2_U3143,
    new_P2_U3144, new_P2_U3145, new_P2_U3146, new_P2_U3147, new_P2_U3148,
    new_P2_U3149, new_P2_U3152, new_P2_U3297, new_P2_U3298, new_P2_U3299,
    new_P2_U3300, new_P2_U3301, new_P2_U3302, new_P2_U3303, new_P2_U3304,
    new_P2_U3305, new_P2_U3306, new_P2_U3307, new_P2_U3308, new_P2_U3309,
    new_P2_U3310, new_P2_U3311, new_P2_U3312, new_P2_U3313, new_P2_U3314,
    new_P2_U3315, new_P2_U3316, new_P2_U3317, new_P2_U3318, new_P2_U3319,
    new_P2_U3320, new_P2_U3321, new_P2_U3322, new_P2_U3323, new_P2_U3324,
    new_P2_U3325, new_P2_U3326, new_P2_U3327, new_P2_U3328, new_P2_U3329,
    new_P2_U3330, new_P2_U3331, new_P2_U3332, new_P2_U3333, new_P2_U3334,
    new_P2_U3335, new_P2_U3336, new_P2_U3337, new_P2_U3338, new_P2_U3339,
    new_P2_U3340, new_P2_U3341, new_P2_U3342, new_P2_U3343, new_P2_U3344,
    new_P2_U3345, new_P2_U3346, new_P2_U3347, new_P2_U3348, new_P2_U3349,
    new_P2_U3350, new_P2_U3351, new_P2_U3352, new_P2_U3353, new_P2_U3354,
    new_P2_U3355, new_P2_U3356, new_P2_U3357, new_P2_U3358, new_P2_U3359,
    new_P2_U3360, new_P2_U3361, new_P2_U3362, new_P2_U3363, new_P2_U3364,
    new_P2_U3365, new_P2_U3366, new_P2_U3367, new_P2_U3368, new_P2_U3369,
    new_P2_U3370, new_P2_U3371, new_P2_U3372, new_P2_U3373, new_P2_U3374,
    new_P2_U3375, new_P2_U3378, new_P2_U3379, new_P2_U3380, new_P2_U3381,
    new_P2_U3382, new_P2_U3383, new_P2_U3384, new_P2_U3385, new_P2_U3386,
    new_P2_U3387, new_P2_U3388, new_P2_U3389, new_P2_U3391, new_P2_U3392,
    new_P2_U3394, new_P2_U3395, new_P2_U3397, new_P2_U3398, new_P2_U3400,
    new_P2_U3401, new_P2_U3403, new_P2_U3404, new_P2_U3406, new_P2_U3407,
    new_P2_U3409, new_P2_U3410, new_P2_U3412, new_P2_U3413, new_P2_U3415,
    new_P2_U3416, new_P2_U3418, new_P2_U3419, new_P2_U3421, new_P2_U3422,
    new_P2_U3424, new_P2_U3425, new_P2_U3427, new_P2_U3428, new_P2_U3430,
    new_P2_U3431, new_P2_U3433, new_P2_U3434, new_P2_U3436, new_P2_U3437,
    new_P2_U3439, new_P2_U3440, new_P2_U3442, new_P2_U3443, new_P2_U3445,
    new_P2_U3523, new_P2_U3524, new_P2_U3525, new_P2_U3526, new_P2_U3527,
    new_P2_U3528, new_P2_U3529, new_P2_U3530, new_P2_U3531, new_P2_U3532,
    new_P2_U3533, new_P2_U3534, new_P2_U3535, new_P2_U3536, new_P2_U3537,
    new_P2_U3538, new_P2_U3539, new_P2_U3540, new_P2_U3541, new_P2_U3542,
    new_P2_U3543, new_P2_U3544, new_P2_U3545, new_P2_U3546, new_P2_U3547,
    new_P2_U3548, new_P2_U3549, new_P2_U3550, new_P2_U3551, new_P2_U3552,
    new_P2_U3553, new_P2_U3554, new_P2_U3555, new_P2_U3556, new_P2_U3557,
    new_P2_U3558, new_P2_U3559, new_P2_U3560, new_P2_U3561, new_P2_U3562,
    new_P2_U3563, new_P2_U3564, new_P2_U3565, new_P2_U3566, new_P2_U3567,
    new_P2_U3568, new_P2_U3569, new_P2_U3570, new_P2_U3571, new_P2_U3572,
    new_P2_U3573, new_P2_U3574, new_P2_U3575, new_P2_U3576, new_P2_U3577,
    new_P2_U3578, new_P2_U3579, new_P2_U3580, new_P2_U3581, new_P2_U3582,
    new_P2_U3583, new_P2_U3584, new_P2_U3585, new_P2_U3586, new_P2_U3587,
    new_P2_U3588, new_P2_U3589, new_P2_U3590, new_P2_U3591, new_P2_U3592,
    new_P2_U3593, new_P2_U3594, new_P2_U3595, new_P2_U3596, new_P2_U3597,
    new_P2_U3598, new_P2_U3599, new_P2_U3600, new_P2_U3601, new_P2_U3602,
    new_P2_U3603, new_P2_U3604, new_P2_U3605, new_P2_U3606, new_P2_U3607,
    new_P2_U3608, new_P2_U3609, new_P2_U3610, new_P2_U3611, new_P2_U3612,
    new_P2_U3613, new_P2_U3614, new_P2_U3615, new_P2_U3616, new_P2_U3617,
    new_P2_U3618, new_P2_U3619, new_P2_U3620, new_P2_U3621, new_P2_U3622,
    new_P2_U3623, new_P2_U3624, new_P2_U3625, new_P2_U3626, new_P2_U3627,
    new_P2_U3628, new_P2_U3629, new_P2_U3630, new_P2_U3631, new_P2_U3632,
    new_P2_U3633, new_P2_U3634, new_P2_U3635, new_P2_U3636, new_P2_U3637,
    new_P2_U3638, new_P2_U3639, new_P2_U3640, new_P2_U3641, new_P2_U3642,
    new_P2_U3643, new_P2_U3644, new_P2_U3645, new_P2_U3646, new_P2_U3647,
    new_P2_U3648, new_P2_U3649, new_P2_U3650, new_P2_U3651, new_P2_U3652,
    new_P2_U3653, new_P2_U3654, new_P2_U3655, new_P2_U3656, new_P2_U3657,
    new_P2_U3658, new_P2_U3659, new_P2_U3660, new_P2_U3661, new_P2_U3662,
    new_P2_U3663, new_P2_U3664, new_P2_U3665, new_P2_U3666, new_P2_U3667,
    new_P2_U3668, new_P2_U3669, new_P2_U3670, new_P2_U3671, new_P2_U3672,
    new_P2_U3673, new_P2_U3674, new_P2_U3675, new_P2_U3676, new_P2_U3677,
    new_P2_U3678, new_P2_U3679, new_P2_U3680, new_P2_U3681, new_P2_U3682,
    new_P2_U3683, new_P2_U3684, new_P2_U3685, new_P2_U3686, new_P2_U3687,
    new_P2_U3688, new_P2_U3689, new_P2_U3690, new_P2_U3691, new_P2_U3692,
    new_P2_U3693, new_P2_U3694, new_P2_U3695, new_P2_U3696, new_P2_U3697,
    new_P2_U3698, new_P2_U3699, new_P2_U3700, new_P2_U3701, new_P2_U3702,
    new_P2_U3703, new_P2_U3704, new_P2_U3705, new_P2_U3706, new_P2_U3707,
    new_P2_U3708, new_P2_U3709, new_P2_U3710, new_P2_U3711, new_P2_U3712,
    new_P2_U3713, new_P2_U3714, new_P2_U3715, new_P2_U3716, new_P2_U3717,
    new_P2_U3718, new_P2_U3719, new_P2_U3720, new_P2_U3721, new_P2_U3722,
    new_P2_U3723, new_P2_U3724, new_P2_U3725, new_P2_U3726, new_P2_U3727,
    new_P2_U3728, new_P2_U3729, new_P2_U3730, new_P2_U3731, new_P2_U3732,
    new_P2_U3733, new_P2_U3734, new_P2_U3735, new_P2_U3736, new_P2_U3737,
    new_P2_U3738, new_P2_U3739, new_P2_U3740, new_P2_U3741, new_P2_U3742,
    new_P2_U3743, new_P2_U3744, new_P2_U3745, new_P2_U3746, new_P2_U3747,
    new_P2_U3748, new_P2_U3749, new_P2_U3750, new_P2_U3751, new_P2_U3752,
    new_P2_U3753, new_P2_U3754, new_P2_U3755, new_P2_U3756, new_P2_U3757,
    new_P2_U3758, new_P2_U3759, new_P2_U3760, new_P2_U3761, new_P2_U3762,
    new_P2_U3763, new_P2_U3764, new_P2_U3765, new_P2_U3766, new_P2_U3767,
    new_P2_U3768, new_P2_U3769, new_P2_U3770, new_P2_U3771, new_P2_U3772,
    new_P2_U3773, new_P2_U3774, new_P2_U3775, new_P2_U3776, new_P2_U3777,
    new_P2_U3778, new_P2_U3779, new_P2_U3780, new_P2_U3781, new_P2_U3782,
    new_P2_U3783, new_P2_U3784, new_P2_U3785, new_P2_U3786, new_P2_U3787,
    new_P2_U3788, new_P2_U3789, new_P2_U3790, new_P2_U3791, new_P2_U3792,
    new_P2_U3793, new_P2_U3794, new_P2_U3795, new_P2_U3796, new_P2_U3797,
    new_P2_U3798, new_P2_U3799, new_P2_U3800, new_P2_U3801, new_P2_U3802,
    new_P2_U3803, new_P2_U3804, new_P2_U3805, new_P2_U3806, new_P2_U3807,
    new_P2_U3808, new_P2_U3809, new_P2_U3810, new_P2_U3811, new_P2_U3812,
    new_P2_U3813, new_P2_U3814, new_P2_U3815, new_P2_U3816, new_P2_U3817,
    new_P2_U3818, new_P2_U3819, new_P2_U3820, new_P2_U3821, new_P2_U3822,
    new_P2_U3823, new_P2_U3824, new_P2_U3825, new_P2_U3826, new_P2_U3827,
    new_P2_U3828, new_P2_U3829, new_P2_U3830, new_P2_U3831, new_P2_U3832,
    new_P2_U3833, new_P2_U3834, new_P2_U3835, new_P2_U3836, new_P2_U3837,
    new_P2_U3838, new_P2_U3839, new_P2_U3840, new_P2_U3841, new_P2_U3842,
    new_P2_U3843, new_P2_U3844, new_P2_U3845, new_P2_U3846, new_P2_U3847,
    new_P2_U3848, new_P2_U3849, new_P2_U3850, new_P2_U3851, new_P2_U3852,
    new_P2_U3853, new_P2_U3854, new_P2_U3855, new_P2_U3856, new_P2_U3857,
    new_P2_U3858, new_P2_U3859, new_P2_U3860, new_P2_U3861, new_P2_U3862,
    new_P2_U3863, new_P2_U3864, new_P2_U3865, new_P2_U3866, new_P2_U3867,
    new_P2_U3868, new_P2_U3869, new_P2_U3870, new_P2_U3871, new_P2_U3872,
    new_P2_U3873, new_P2_U3874, new_P2_U3875, new_P2_U3876, new_P2_U3877,
    new_P2_U3878, new_P2_U3879, new_P2_U3880, new_P2_U3881, new_P2_U3882,
    new_P2_U3883, new_P2_U3884, new_P2_U3885, new_P2_U3886, new_P2_U3887,
    new_P2_U3888, new_P2_U3889, new_P2_U3890, new_P2_U3891, new_P2_U3892,
    new_P2_U3894, new_P2_U3895, new_P2_U3896, new_P2_U3897, new_P2_U3898,
    new_P2_U3899, new_P2_U3900, new_P2_U3901, new_P2_U3902, new_P2_U3903,
    new_P2_U3904, new_P2_U3905, new_P2_U3906, new_P2_U3907, new_P2_U3908,
    new_P2_U3909, new_P2_U3910, new_P2_U3911, new_P2_U3912, new_P2_U3913,
    new_P2_U3914, new_P2_U3915, new_P2_U3916, new_P2_U3917, new_P2_U3918,
    new_P2_U3919, new_P2_U3920, new_P2_U3921, new_P2_U3922, new_P2_U3923,
    new_P2_U3924, new_P2_U3925, new_P2_U3926, new_P2_U3927, new_P2_U3928,
    new_P2_U3929, new_P2_U3930, new_P2_U3931, new_P2_U3932, new_P2_U3933,
    new_P2_U3934, new_P2_U3935, new_P2_U3936, new_P2_U3937, new_P2_U3938,
    new_P2_U3939, new_P2_U3940, new_P2_U3941, new_P2_U3942, new_P2_U3943,
    new_P2_U3944, new_P2_U3945, new_P2_U3946, new_P2_U3947, new_P2_U3948,
    new_P2_U3949, new_P2_U3950, new_P2_U3951, new_P2_U3952, new_P2_U3953,
    new_P2_U3954, new_P2_U3955, new_P2_U3956, new_P2_U3957, new_P2_U3958,
    new_P2_U3959, new_P2_U3960, new_P2_U3961, new_P2_U3962, new_P2_U3963,
    new_P2_U3964, new_P2_U3965, new_P2_U3966, new_P2_U3967, new_P2_U3968,
    new_P2_U3969, new_P2_U3970, new_P2_U3971, new_P2_U3972, new_P2_U3973,
    new_P2_U3974, new_P2_U3975, new_P2_U3976, new_P2_U3977, new_P2_U3978,
    new_P2_U3979, new_P2_U3980, new_P2_U3981, new_P2_U3982, new_P2_U3983,
    new_P2_U3984, new_P2_U3985, new_P2_U3986, new_P2_U3987, new_P2_U3988,
    new_P2_U3989, new_P2_U3990, new_P2_U3991, new_P2_U3992, new_P2_U3993,
    new_P2_U3994, new_P2_U3995, new_P2_U3996, new_P2_U3997, new_P2_U3998,
    new_P2_U3999, new_P2_U4000, new_P2_U4001, new_P2_U4002, new_P2_U4003,
    new_P2_U4004, new_P2_U4005, new_P2_U4006, new_P2_U4007, new_P2_U4008,
    new_P2_U4009, new_P2_U4010, new_P2_U4011, new_P2_U4012, new_P2_U4013,
    new_P2_U4014, new_P2_U4015, new_P2_U4016, new_P2_U4017, new_P2_U4018,
    new_P2_U4019, new_P2_U4020, new_P2_U4021, new_P2_U4022, new_P2_U4023,
    new_P2_U4024, new_P2_U4025, new_P2_U4026, new_P2_U4027, new_P2_U4028,
    new_P2_U4029, new_P2_U4030, new_P2_U4031, new_P2_U4032, new_P2_U4033,
    new_P2_U4034, new_P2_U4035, new_P2_U4036, new_P2_U4037, new_P2_U4038,
    new_P2_U4039, new_P2_U4040, new_P2_U4041, new_P2_U4042, new_P2_U4043,
    new_P2_U4044, new_P2_U4045, new_P2_U4046, new_P2_U4047, new_P2_U4048,
    new_P2_U4049, new_P2_U4050, new_P2_U4051, new_P2_U4052, new_P2_U4053,
    new_P2_U4054, new_P2_U4055, new_P2_U4056, new_P2_U4057, new_P2_U4058,
    new_P2_U4059, new_P2_U4060, new_P2_U4061, new_P2_U4062, new_P2_U4063,
    new_P2_U4064, new_P2_U4065, new_P2_U4066, new_P2_U4067, new_P2_U4068,
    new_P2_U4069, new_P2_U4070, new_P2_U4071, new_P2_U4072, new_P2_U4073,
    new_P2_U4074, new_P2_U4075, new_P2_U4076, new_P2_U4077, new_P2_U4078,
    new_P2_U4079, new_P2_U4080, new_P2_U4081, new_P2_U4082, new_P2_U4083,
    new_P2_U4084, new_P2_U4085, new_P2_U4086, new_P2_U4087, new_P2_U4088,
    new_P2_U4089, new_P2_U4090, new_P2_U4091, new_P2_U4092, new_P2_U4093,
    new_P2_U4094, new_P2_U4095, new_P2_U4096, new_P2_U4097, new_P2_U4098,
    new_P2_U4099, new_P2_U4100, new_P2_U4101, new_P2_U4102, new_P2_U4103,
    new_P2_U4104, new_P2_U4105, new_P2_U4106, new_P2_U4107, new_P2_U4108,
    new_P2_U4109, new_P2_U4110, new_P2_U4111, new_P2_U4112, new_P2_U4113,
    new_P2_U4114, new_P2_U4115, new_P2_U4116, new_P2_U4117, new_P2_U4118,
    new_P2_U4119, new_P2_U4120, new_P2_U4121, new_P2_U4122, new_P2_U4123,
    new_P2_U4124, new_P2_U4125, new_P2_U4126, new_P2_U4127, new_P2_U4128,
    new_P2_U4129, new_P2_U4130, new_P2_U4131, new_P2_U4132, new_P2_U4133,
    new_P2_U4134, new_P2_U4135, new_P2_U4136, new_P2_U4137, new_P2_U4138,
    new_P2_U4139, new_P2_U4140, new_P2_U4141, new_P2_U4142, new_P2_U4143,
    new_P2_U4144, new_P2_U4145, new_P2_U4146, new_P2_U4147, new_P2_U4148,
    new_P2_U4149, new_P2_U4150, new_P2_U4151, new_P2_U4152, new_P2_U4153,
    new_P2_U4154, new_P2_U4155, new_P2_U4156, new_P2_U4157, new_P2_U4158,
    new_P2_U4159, new_P2_U4160, new_P2_U4161, new_P2_U4162, new_P2_U4163,
    new_P2_U4164, new_P2_U4165, new_P2_U4166, new_P2_U4167, new_P2_U4168,
    new_P2_U4169, new_P2_U4170, new_P2_U4171, new_P2_U4172, new_P2_U4173,
    new_P2_U4174, new_P2_U4175, new_P2_U4176, new_P2_U4177, new_P2_U4178,
    new_P2_U4179, new_P2_U4180, new_P2_U4181, new_P2_U4182, new_P2_U4183,
    new_P2_U4184, new_P2_U4185, new_P2_U4186, new_P2_U4187, new_P2_U4188,
    new_P2_U4189, new_P2_U4190, new_P2_U4191, new_P2_U4192, new_P2_U4193,
    new_P2_U4194, new_P2_U4195, new_P2_U4196, new_P2_U4197, new_P2_U4198,
    new_P2_U4199, new_P2_U4200, new_P2_U4201, new_P2_U4202, new_P2_U4203,
    new_P2_U4204, new_P2_U4205, new_P2_U4206, new_P2_U4207, new_P2_U4208,
    new_P2_U4209, new_P2_U4210, new_P2_U4211, new_P2_U4212, new_P2_U4213,
    new_P2_U4214, new_P2_U4215, new_P2_U4216, new_P2_U4217, new_P2_U4218,
    new_P2_U4219, new_P2_U4220, new_P2_U4221, new_P2_U4222, new_P2_U4223,
    new_P2_U4224, new_P2_U4225, new_P2_U4226, new_P2_U4227, new_P2_U4228,
    new_P2_U4229, new_P2_U4230, new_P2_U4231, new_P2_U4232, new_P2_U4233,
    new_P2_U4234, new_P2_U4235, new_P2_U4236, new_P2_U4237, new_P2_U4238,
    new_P2_U4239, new_P2_U4240, new_P2_U4241, new_P2_U4242, new_P2_U4243,
    new_P2_U4244, new_P2_U4245, new_P2_U4246, new_P2_U4247, new_P2_U4248,
    new_P2_U4249, new_P2_U4250, new_P2_U4251, new_P2_U4252, new_P2_U4253,
    new_P2_U4254, new_P2_U4255, new_P2_U4256, new_P2_U4257, new_P2_U4258,
    new_P2_U4259, new_P2_U4260, new_P2_U4261, new_P2_U4262, new_P2_U4263,
    new_P2_U4264, new_P2_U4265, new_P2_U4266, new_P2_U4267, new_P2_U4268,
    new_P2_U4269, new_P2_U4270, new_P2_U4271, new_P2_U4272, new_P2_U4273,
    new_P2_U4274, new_P2_U4275, new_P2_U4276, new_P2_U4277, new_P2_U4278,
    new_P2_U4279, new_P2_U4280, new_P2_U4281, new_P2_U4282, new_P2_U4283,
    new_P2_U4284, new_P2_U4285, new_P2_U4286, new_P2_U4287, new_P2_U4288,
    new_P2_U4289, new_P2_U4290, new_P2_U4291, new_P2_U4292, new_P2_U4293,
    new_P2_U4294, new_P2_U4295, new_P2_U4296, new_P2_U4297, new_P2_U4298,
    new_P2_U4299, new_P2_U4300, new_P2_U4301, new_P2_U4302, new_P2_U4303,
    new_P2_U4304, new_P2_U4305, new_P2_U4306, new_P2_U4307, new_P2_U4308,
    new_P2_U4309, new_P2_U4310, new_P2_U4311, new_P2_U4312, new_P2_U4313,
    new_P2_U4314, new_P2_U4315, new_P2_U4316, new_P2_U4317, new_P2_U4318,
    new_P2_U4319, new_P2_U4320, new_P2_U4321, new_P2_U4322, new_P2_U4323,
    new_P2_U4324, new_P2_U4325, new_P2_U4326, new_P2_U4327, new_P2_U4328,
    new_P2_U4329, new_P2_U4330, new_P2_U4331, new_P2_U4332, new_P2_U4333,
    new_P2_U4334, new_P2_U4335, new_P2_U4336, new_P2_U4337, new_P2_U4338,
    new_P2_U4339, new_P2_U4340, new_P2_U4341, new_P2_U4342, new_P2_U4343,
    new_P2_U4344, new_P2_U4345, new_P2_U4346, new_P2_U4347, new_P2_U4348,
    new_P2_U4349, new_P2_U4350, new_P2_U4351, new_P2_U4352, new_P2_U4353,
    new_P2_U4354, new_P2_U4355, new_P2_U4356, new_P2_U4357, new_P2_U4358,
    new_P2_U4359, new_P2_U4360, new_P2_U4361, new_P2_U4362, new_P2_U4363,
    new_P2_U4364, new_P2_U4365, new_P2_U4366, new_P2_U4367, new_P2_U4368,
    new_P2_U4369, new_P2_U4370, new_P2_U4371, new_P2_U4372, new_P2_U4373,
    new_P2_U4374, new_P2_U4375, new_P2_U4376, new_P2_U4377, new_P2_U4378,
    new_P2_U4379, new_P2_U4380, new_P2_U4381, new_P2_U4382, new_P2_U4383,
    new_P2_U4384, new_P2_U4385, new_P2_U4386, new_P2_U4387, new_P2_U4388,
    new_P2_U4389, new_P2_U4390, new_P2_U4391, new_P2_U4392, new_P2_U4393,
    new_P2_U4394, new_P2_U4395, new_P2_U4396, new_P2_U4397, new_P2_U4398,
    new_P2_U4399, new_P2_U4400, new_P2_U4401, new_P2_U4402, new_P2_U4403,
    new_P2_U4404, new_P2_U4405, new_P2_U4406, new_P2_U4407, new_P2_U4408,
    new_P2_U4409, new_P2_U4410, new_P2_U4411, new_P2_U4412, new_P2_U4413,
    new_P2_U4414, new_P2_U4415, new_P2_U4416, new_P2_U4417, new_P2_U4418,
    new_P2_U4419, new_P2_U4420, new_P2_U4421, new_P2_U4422, new_P2_U4423,
    new_P2_U4424, new_P2_U4425, new_P2_U4426, new_P2_U4427, new_P2_U4428,
    new_P2_U4429, new_P2_U4430, new_P2_U4431, new_P2_U4432, new_P2_U4433,
    new_P2_U4434, new_P2_U4435, new_P2_U4436, new_P2_U4437, new_P2_U4438,
    new_P2_U4439, new_P2_U4440, new_P2_U4441, new_P2_U4442, new_P2_U4443,
    new_P2_U4444, new_P2_U4445, new_P2_U4446, new_P2_U4447, new_P2_U4448,
    new_P2_U4449, new_P2_U4450, new_P2_U4451, new_P2_U4452, new_P2_U4453,
    new_P2_U4454, new_P2_U4455, new_P2_U4456, new_P2_U4457, new_P2_U4458,
    new_P2_U4459, new_P2_U4460, new_P2_U4461, new_P2_U4462, new_P2_U4463,
    new_P2_U4464, new_P2_U4465, new_P2_U4466, new_P2_U4467, new_P2_U4468,
    new_P2_U4469, new_P2_U4470, new_P2_U4471, new_P2_U4472, new_P2_U4473,
    new_P2_U4474, new_P2_U4475, new_P2_U4476, new_P2_U4477, new_P2_U4478,
    new_P2_U4479, new_P2_U4480, new_P2_U4481, new_P2_U4482, new_P2_U4483,
    new_P2_U4484, new_P2_U4485, new_P2_U4486, new_P2_U4487, new_P2_U4488,
    new_P2_U4489, new_P2_U4490, new_P2_U4491, new_P2_U4492, new_P2_U4493,
    new_P2_U4494, new_P2_U4495, new_P2_U4496, new_P2_U4497, new_P2_U4498,
    new_P2_U4499, new_P2_U4500, new_P2_U4501, new_P2_U4502, new_P2_U4503,
    new_P2_U4504, new_P2_U4505, new_P2_U4506, new_P2_U4507, new_P2_U4508,
    new_P2_U4509, new_P2_U4510, new_P2_U4511, new_P2_U4512, new_P2_U4513,
    new_P2_U4514, new_P2_U4515, new_P2_U4516, new_P2_U4517, new_P2_U4518,
    new_P2_U4519, new_P2_U4520, new_P2_U4521, new_P2_U4522, new_P2_U4523,
    new_P2_U4524, new_P2_U4525, new_P2_U4526, new_P2_U4527, new_P2_U4528,
    new_P2_U4529, new_P2_U4530, new_P2_U4531, new_P2_U4532, new_P2_U4533,
    new_P2_U4534, new_P2_U4535, new_P2_U4536, new_P2_U4537, new_P2_U4538,
    new_P2_U4539, new_P2_U4540, new_P2_U4541, new_P2_U4542, new_P2_U4543,
    new_P2_U4544, new_P2_U4545, new_P2_U4546, new_P2_U4547, new_P2_U4548,
    new_P2_U4549, new_P2_U4550, new_P2_U4551, new_P2_U4552, new_P2_U4553,
    new_P2_U4554, new_P2_U4555, new_P2_U4556, new_P2_U4557, new_P2_U4558,
    new_P2_U4559, new_P2_U4560, new_P2_U4561, new_P2_U4562, new_P2_U4563,
    new_P2_U4564, new_P2_U4565, new_P2_U4566, new_P2_U4567, new_P2_U4568,
    new_P2_U4569, new_P2_U4570, new_P2_U4571, new_P2_U4572, new_P2_U4573,
    new_P2_U4574, new_P2_U4575, new_P2_U4576, new_P2_U4577, new_P2_U4578,
    new_P2_U4579, new_P2_U4580, new_P2_U4581, new_P2_U4582, new_P2_U4583,
    new_P2_U4584, new_P2_U4585, new_P2_U4586, new_P2_U4587, new_P2_U4588,
    new_P2_U4589, new_P2_U4590, new_P2_U4591, new_P2_U4592, new_P2_U4593,
    new_P2_U4594, new_P2_U4595, new_P2_U4596, new_P2_U4597, new_P2_U4598,
    new_P2_U4599, new_P2_U4600, new_P2_U4601, new_P2_U4602, new_P2_U4603,
    new_P2_U4604, new_P2_U4605, new_P2_U4606, new_P2_U4607, new_P2_U4608,
    new_P2_U4609, new_P2_U4610, new_P2_U4611, new_P2_U4612, new_P2_U4613,
    new_P2_U4614, new_P2_U4615, new_P2_U4616, new_P2_U4617, new_P2_U4618,
    new_P2_U4619, new_P2_U4620, new_P2_U4621, new_P2_U4622, new_P2_U4623,
    new_P2_U4624, new_P2_U4625, new_P2_U4626, new_P2_U4627, new_P2_U4628,
    new_P2_U4629, new_P2_U4630, new_P2_U4631, new_P2_U4632, new_P2_U4633,
    new_P2_U4634, new_P2_U4635, new_P2_U4636, new_P2_U4637, new_P2_U4638,
    new_P2_U4639, new_P2_U4640, new_P2_U4641, new_P2_U4642, new_P2_U4643,
    new_P2_U4644, new_P2_U4645, new_P2_U4646, new_P2_U4647, new_P2_U4648,
    new_P2_U4649, new_P2_U4650, new_P2_U4651, new_P2_U4652, new_P2_U4653,
    new_P2_U4654, new_P2_U4655, new_P2_U4656, new_P2_U4657, new_P2_U4658,
    new_P2_U4659, new_P2_U4660, new_P2_U4661, new_P2_U4662, new_P2_U4663,
    new_P2_U4664, new_P2_U4665, new_P2_U4666, new_P2_U4667, new_P2_U4668,
    new_P2_U4669, new_P2_U4670, new_P2_U4671, new_P2_U4672, new_P2_U4673,
    new_P2_U4674, new_P2_U4675, new_P2_U4676, new_P2_U4677, new_P2_U4678,
    new_P2_U4679, new_P2_U4680, new_P2_U4681, new_P2_U4682, new_P2_U4683,
    new_P2_U4684, new_P2_U4685, new_P2_U4686, new_P2_U4687, new_P2_U4688,
    new_P2_U4689, new_P2_U4690, new_P2_U4691, new_P2_U4692, new_P2_U4693,
    new_P2_U4694, new_P2_U4695, new_P2_U4696, new_P2_U4697, new_P2_U4698,
    new_P2_U4699, new_P2_U4700, new_P2_U4701, new_P2_U4702, new_P2_U4703,
    new_P2_U4704, new_P2_U4705, new_P2_U4706, new_P2_U4707, new_P2_U4708,
    new_P2_U4709, new_P2_U4710, new_P2_U4711, new_P2_U4712, new_P2_U4713,
    new_P2_U4714, new_P2_U4715, new_P2_U4716, new_P2_U4717, new_P2_U4718,
    new_P2_U4719, new_P2_U4720, new_P2_U4721, new_P2_U4722, new_P2_U4723,
    new_P2_U4724, new_P2_U4725, new_P2_U4726, new_P2_U4727, new_P2_U4728,
    new_P2_U4729, new_P2_U4730, new_P2_U4731, new_P2_U4732, new_P2_U4733,
    new_P2_U4734, new_P2_U4735, new_P2_U4736, new_P2_U4737, new_P2_U4738,
    new_P2_U4739, new_P2_U4740, new_P2_U4741, new_P2_U4742, new_P2_U4743,
    new_P2_U4744, new_P2_U4745, new_P2_U4746, new_P2_U4747, new_P2_U4748,
    new_P2_U4749, new_P2_U4750, new_P2_U4751, new_P2_U4752, new_P2_U4753,
    new_P2_U4754, new_P2_U4755, new_P2_U4756, new_P2_U4757, new_P2_U4758,
    new_P2_U4759, new_P2_U4760, new_P2_U4761, new_P2_U4762, new_P2_U4763,
    new_P2_U4764, new_P2_U4765, new_P2_U4766, new_P2_U4767, new_P2_U4768,
    new_P2_U4769, new_P2_U4770, new_P2_U4771, new_P2_U4772, new_P2_U4773,
    new_P2_U4774, new_P2_U4775, new_P2_U4776, new_P2_U4777, new_P2_U4778,
    new_P2_U4779, new_P2_U4780, new_P2_U4781, new_P2_U4782, new_P2_U4783,
    new_P2_U4784, new_P2_U4785, new_P2_U4786, new_P2_U4787, new_P2_U4788,
    new_P2_U4789, new_P2_U4790, new_P2_U4791, new_P2_U4792, new_P2_U4793,
    new_P2_U4794, new_P2_U4795, new_P2_U4796, new_P2_U4797, new_P2_U4798,
    new_P2_U4799, new_P2_U4800, new_P2_U4801, new_P2_U4802, new_P2_U4803,
    new_P2_U4804, new_P2_U4805, new_P2_U4806, new_P2_U4807, new_P2_U4808,
    new_P2_U4809, new_P2_U4810, new_P2_U4811, new_P2_U4812, new_P2_U4813,
    new_P2_U4814, new_P2_U4815, new_P2_U4816, new_P2_U4817, new_P2_U4818,
    new_P2_U4819, new_P2_U4820, new_P2_U4821, new_P2_U4822, new_P2_U4823,
    new_P2_U4824, new_P2_U4825, new_P2_U4826, new_P2_U4827, new_P2_U4828,
    new_P2_U4829, new_P2_U4830, new_P2_U4831, new_P2_U4832, new_P2_U4833,
    new_P2_U4834, new_P2_U4835, new_P2_U4836, new_P2_U4837, new_P2_U4838,
    new_P2_U4839, new_P2_U4840, new_P2_U4841, new_P2_U4842, new_P2_U4843,
    new_P2_U4844, new_P2_U4845, new_P2_U4846, new_P2_U4847, new_P2_U4848,
    new_P2_U4849, new_P2_U4850, new_P2_U4851, new_P2_U4852, new_P2_U4853,
    new_P2_U4854, new_P2_U4855, new_P2_U4856, new_P2_U4857, new_P2_U4858,
    new_P2_U4859, new_P2_U4860, new_P2_U4861, new_P2_U4862, new_P2_U4863,
    new_P2_U4864, new_P2_U4865, new_P2_U4866, new_P2_U4867, new_P2_U4868,
    new_P2_U4869, new_P2_U4870, new_P2_U4871, new_P2_U4872, new_P2_U4873,
    new_P2_U4874, new_P2_U4875, new_P2_U4876, new_P2_U4877, new_P2_U4878,
    new_P2_U4879, new_P2_U4880, new_P2_U4881, new_P2_U4882, new_P2_U4883,
    new_P2_U4884, new_P2_U4885, new_P2_U4886, new_P2_U4887, new_P2_U4888,
    new_P2_U4889, new_P2_U4890, new_P2_U4891, new_P2_U4892, new_P2_U4893,
    new_P2_U4894, new_P2_U4895, new_P2_U4896, new_P2_U4897, new_P2_U4898,
    new_P2_U4899, new_P2_U4900, new_P2_U4901, new_P2_U4902, new_P2_U4903,
    new_P2_U4904, new_P2_U4905, new_P2_U4906, new_P2_U4907, new_P2_U4908,
    new_P2_U4909, new_P2_U4910, new_P2_U4911, new_P2_U4912, new_P2_U4913,
    new_P2_U4914, new_P2_U4915, new_P2_U4916, new_P2_U4917, new_P2_U4918,
    new_P2_U4919, new_P2_U4920, new_P2_U4921, new_P2_U4922, new_P2_U4923,
    new_P2_U4924, new_P2_U4925, new_P2_U4926, new_P2_U4927, new_P2_U4928,
    new_P2_U4929, new_P2_U4930, new_P2_U4931, new_P2_U4932, new_P2_U4933,
    new_P2_U4934, new_P2_U4935, new_P2_U4936, new_P2_U4937, new_P2_U4938,
    new_P2_U4939, new_P2_U4940, new_P2_U4941, new_P2_U4942, new_P2_U4943,
    new_P2_U4944, new_P2_U4945, new_P2_U4946, new_P2_U4947, new_P2_U4948,
    new_P2_U4949, new_P2_U4950, new_P2_U4951, new_P2_U4952, new_P2_U4953,
    new_P2_U4954, new_P2_U4955, new_P2_U4956, new_P2_U4957, new_P2_U4958,
    new_P2_U4959, new_P2_U4960, new_P2_U4961, new_P2_U4962, new_P2_U4963,
    new_P2_U4964, new_P2_U4965, new_P2_U4966, new_P2_U4967, new_P2_U4968,
    new_P2_U4969, new_P2_U4970, new_P2_U4971, new_P2_U4972, new_P2_U4973,
    new_P2_U4974, new_P2_U4975, new_P2_U4976, new_P2_U4977, new_P2_U4978,
    new_P2_U4979, new_P2_U4980, new_P2_U4981, new_P2_U4982, new_P2_U4983,
    new_P2_U4984, new_P2_U4985, new_P2_U4986, new_P2_U4987, new_P2_U4988,
    new_P2_U4989, new_P2_U4990, new_P2_U4991, new_P2_U4992, new_P2_U4993,
    new_P2_U4994, new_P2_U4995, new_P2_U4996, new_P2_U4997, new_P2_U4998,
    new_P2_U4999, new_P2_U5000, new_P2_U5001, new_P2_U5002, new_P2_U5003,
    new_P2_U5004, new_P2_U5005, new_P2_U5006, new_P2_U5007, new_P2_U5008,
    new_P2_U5009, new_P2_U5010, new_P2_U5011, new_P2_U5012, new_P2_U5013,
    new_P2_U5014, new_P2_U5015, new_P2_U5016, new_P2_U5017, new_P2_U5018,
    new_P2_U5019, new_P2_U5020, new_P2_U5021, new_P2_U5022, new_P2_U5023,
    new_P2_U5024, new_P2_U5025, new_P2_U5026, new_P2_U5027, new_P2_U5028,
    new_P2_U5029, new_P2_U5030, new_P2_U5031, new_P2_U5032, new_P2_U5033,
    new_P2_U5034, new_P2_U5035, new_P2_U5036, new_P2_U5037, new_P2_U5038,
    new_P2_U5039, new_P2_U5040, new_P2_U5041, new_P2_U5042, new_P2_U5043,
    new_P2_U5044, new_P2_U5045, new_P2_U5046, new_P2_U5047, new_P2_U5048,
    new_P2_U5049, new_P2_U5050, new_P2_U5051, new_P2_U5052, new_P2_U5053,
    new_P2_U5054, new_P2_U5055, new_P2_U5056, new_P2_U5057, new_P2_U5058,
    new_P2_U5059, new_P2_U5060, new_P2_U5061, new_P2_U5062, new_P2_U5063,
    new_P2_U5064, new_P2_U5065, new_P2_U5066, new_P2_U5067, new_P2_U5068,
    new_P2_U5069, new_P2_U5070, new_P2_U5071, new_P2_U5072, new_P2_U5073,
    new_P2_U5074, new_P2_U5075, new_P2_U5076, new_P2_U5077, new_P2_U5078,
    new_P2_U5079, new_P2_U5080, new_P2_U5081, new_P2_U5082, new_P2_U5083,
    new_P2_U5084, new_P2_U5085, new_P2_U5086, new_P2_U5087, new_P2_U5088,
    new_P2_U5089, new_P2_U5090, new_P2_U5091, new_P2_U5092, new_P2_U5093,
    new_P2_U5094, new_P2_U5095, new_P2_U5096, new_P2_U5097, new_P2_U5098,
    new_P2_U5099, new_P2_U5100, new_P2_U5101, new_P2_U5102, new_P2_U5103,
    new_P2_U5104, new_P2_U5105, new_P2_U5106, new_P2_U5107, new_P2_U5108,
    new_P2_U5109, new_P2_U5110, new_P2_U5111, new_P2_U5112, new_P2_U5113,
    new_P2_U5114, new_P2_U5115, new_P2_U5116, new_P2_U5117, new_P2_U5118,
    new_P2_U5119, new_P2_U5120, new_P2_U5121, new_P2_U5122, new_P2_U5123,
    new_P2_U5124, new_P2_U5125, new_P2_U5126, new_P2_U5127, new_P2_U5128,
    new_P2_U5129, new_P2_U5130, new_P2_U5131, new_P2_U5132, new_P2_U5133,
    new_P2_U5134, new_P2_U5135, new_P2_U5136, new_P2_U5137, new_P2_U5138,
    new_P2_U5139, new_P2_U5140, new_P2_U5141, new_P2_U5142, new_P2_U5143,
    new_P2_U5144, new_P2_U5145, new_P2_U5146, new_P2_U5147, new_P2_U5148,
    new_P2_U5149, new_P2_U5150, new_P2_U5151, new_P2_U5152, new_P2_U5153,
    new_P2_U5154, new_P2_U5155, new_P2_U5156, new_P2_U5157, new_P2_U5158,
    new_P2_U5159, new_P2_U5160, new_P2_U5161, new_P2_U5162, new_P2_U5163,
    new_P2_U5164, new_P2_U5165, new_P2_U5166, new_P2_U5167, new_P2_U5168,
    new_P2_U5169, new_P2_U5170, new_P2_U5171, new_P2_U5172, new_P2_U5173,
    new_P2_U5174, new_P2_U5175, new_P2_U5176, new_P2_U5177, new_P2_U5178,
    new_P2_U5179, new_P2_U5180, new_P2_U5181, new_P2_U5182, new_P2_U5183,
    new_P2_U5184, new_P2_U5185, new_P2_U5186, new_P2_U5187, new_P2_U5188,
    new_P2_U5189, new_P2_U5190, new_P2_U5191, new_P2_U5192, new_P2_U5193,
    new_P2_U5194, new_P2_U5195, new_P2_U5196, new_P2_U5197, new_P2_U5198,
    new_P2_U5199, new_P2_U5200, new_P2_U5201, new_P2_U5202, new_P2_U5203,
    new_P2_U5204, new_P2_U5205, new_P2_U5206, new_P2_U5207, new_P2_U5208,
    new_P2_U5209, new_P2_U5210, new_P2_U5211, new_P2_U5212, new_P2_U5213,
    new_P2_U5214, new_P2_U5215, new_P2_U5216, new_P2_U5217, new_P2_U5218,
    new_P2_U5219, new_P2_U5220, new_P2_U5221, new_P2_U5222, new_P2_U5223,
    new_P2_U5224, new_P2_U5225, new_P2_U5226, new_P2_U5227, new_P2_U5228,
    new_P2_U5229, new_P2_U5230, new_P2_U5231, new_P2_U5232, new_P2_U5233,
    new_P2_U5234, new_P2_U5235, new_P2_U5236, new_P2_U5237, new_P2_U5238,
    new_P2_U5239, new_P2_U5240, new_P2_U5241, new_P2_U5242, new_P2_U5243,
    new_P2_U5244, new_P2_U5245, new_P2_U5246, new_P2_U5247, new_P2_U5248,
    new_P2_U5249, new_P2_U5250, new_P2_U5251, new_P2_U5252, new_P2_U5253,
    new_P2_U5254, new_P2_U5255, new_P2_U5256, new_P2_U5257, new_P2_U5258,
    new_P2_U5259, new_P2_U5260, new_P2_U5261, new_P2_U5262, new_P2_U5263,
    new_P2_U5264, new_P2_U5265, new_P2_U5266, new_P2_U5267, new_P2_U5268,
    new_P2_U5269, new_P2_U5270, new_P2_U5271, new_P2_U5272, new_P2_U5273,
    new_P2_U5274, new_P2_U5275, new_P2_U5276, new_P2_U5277, new_P2_U5278,
    new_P2_U5279, new_P2_U5280, new_P2_U5281, new_P2_U5282, new_P2_U5283,
    new_P2_U5284, new_P2_U5285, new_P2_U5286, new_P2_U5287, new_P2_U5288,
    new_P2_U5289, new_P2_U5290, new_P2_U5291, new_P2_U5292, new_P2_U5293,
    new_P2_U5294, new_P2_U5295, new_P2_U5296, new_P2_U5297, new_P2_U5298,
    new_P2_U5299, new_P2_U5300, new_P2_U5301, new_P2_U5302, new_P2_U5303,
    new_P2_U5304, new_P2_U5305, new_P2_U5306, new_P2_U5307, new_P2_U5308,
    new_P2_U5309, new_P2_U5310, new_P2_U5311, new_P2_U5312, new_P2_U5313,
    new_P2_U5314, new_P2_U5315, new_P2_U5316, new_P2_U5317, new_P2_U5318,
    new_P2_U5319, new_P2_U5320, new_P2_U5321, new_P2_U5322, new_P2_U5323,
    new_P2_U5324, new_P2_U5325, new_P2_U5326, new_P2_U5327, new_P2_U5328,
    new_P2_U5329, new_P2_U5330, new_P2_U5331, new_P2_U5332, new_P2_U5333,
    new_P2_U5334, new_P2_U5335, new_P2_U5336, new_P2_U5337, new_P2_U5338,
    new_P2_U5339, new_P2_U5340, new_P2_U5341, new_P2_U5342, new_P2_U5343,
    new_P2_U5344, new_P2_U5345, new_P2_U5346, new_P2_U5347, new_P2_U5348,
    new_P2_U5349, new_P2_U5350, new_P2_U5351, new_P2_U5352, new_P2_U5353,
    new_P2_U5354, new_P2_U5355, new_P2_U5356, new_P2_U5357, new_P2_U5358,
    new_P2_U5359, new_P2_U5360, new_P2_U5361, new_P2_U5362, new_P2_U5363,
    new_P2_U5364, new_P2_U5365, new_P2_U5366, new_P2_U5367, new_P2_U5368,
    new_P2_U5369, new_P2_U5370, new_P2_U5371, new_P2_U5372, new_P2_U5373,
    new_P2_U5374, new_P2_U5375, new_P2_U5376, new_P2_U5377, new_P2_U5378,
    new_P2_U5379, new_P2_U5380, new_P2_U5381, new_P2_U5382, new_P2_U5383,
    new_P2_U5384, new_P2_U5385, new_P2_U5386, new_P2_U5387, new_P2_U5388,
    new_P2_U5389, new_P2_U5390, new_P2_U5391, new_P2_U5392, new_P2_U5393,
    new_P2_U5394, new_P2_U5395, new_P2_U5396, new_P2_U5397, new_P2_U5398,
    new_P2_U5399, new_P2_U5400, new_P2_U5401, new_P2_U5402, new_P2_U5403,
    new_P2_U5404, new_P2_U5405, new_P2_U5406, new_P2_U5407, new_P2_U5408,
    new_P2_U5409, new_P2_U5410, new_P2_U5411, new_P2_U5412, new_P2_U5413,
    new_P2_U5414, new_P2_U5415, new_P2_U5416, new_P2_U5417, new_P2_U5418,
    new_P2_U5419, new_P2_U5420, new_P2_U5421, new_P2_U5422, new_P2_U5423,
    new_P2_U5424, new_P2_U5425, new_P2_U5426, new_P2_U5427, new_P2_U5428,
    new_P2_U5429, new_P2_U5430, new_P2_U5431, new_P2_U5432, new_P2_U5433,
    new_P2_U5434, new_P2_U5435, new_P2_U5436, new_P2_U5437, new_P2_U5438,
    new_P2_U5439, new_P2_U5440, new_P2_U5441, new_P2_U5442, new_P2_U5443,
    new_P2_U5444, new_P2_U5445, new_P2_U5446, new_P2_U5447, new_P2_U5448,
    new_P2_U5449, new_P2_U5450, new_P2_U5451, new_P2_U5452, new_P2_U5453,
    new_P2_U5454, new_P2_U5455, new_P2_U5456, new_P2_U5457, new_P2_U5458,
    new_P2_U5459, new_P2_U5460, new_P2_U5461, new_P2_U5462, new_P2_U5463,
    new_P2_U5464, new_P2_U5465, new_P2_U5466, new_P2_U5467, new_P2_U5468,
    new_P2_U5469, new_P2_U5470, new_P2_U5471, new_P2_U5472, new_P2_U5473,
    new_P2_U5474, new_P2_U5475, new_P2_U5476, new_P2_U5477, new_P2_U5478,
    new_P2_U5479, new_P2_U5480, new_P2_U5481, new_P2_U5482, new_P2_U5483,
    new_P2_U5484, new_P2_U5485, new_P2_U5486, new_P2_U5487, new_P2_U5488,
    new_P2_U5489, new_P2_U5490, new_P2_U5491, new_P2_U5492, new_P2_U5493,
    new_P2_U5494, new_P2_U5495, new_P2_U5496, new_P2_U5497, new_P2_U5498,
    new_P2_U5499, new_P2_U5500, new_P2_U5501, new_P2_U5502, new_P2_U5503,
    new_P2_U5504, new_P2_U5505, new_P2_U5506, new_P2_U5507, new_P2_U5508,
    new_P2_U5509, new_P2_U5510, new_P2_U5511, new_P2_U5512, new_P2_U5513,
    new_P2_U5514, new_P2_U5515, new_P2_U5516, new_P2_U5517, new_P2_U5518,
    new_P2_U5519, new_P2_U5520, new_P2_U5521, new_P2_U5522, new_P2_U5523,
    new_P2_U5524, new_P2_U5525, new_P2_U5526, new_P2_U5527, new_P2_U5528,
    new_P2_U5529, new_P2_U5530, new_P2_U5531, new_P2_U5532, new_P2_U5533,
    new_P2_U5534, new_P2_U5535, new_P2_U5536, new_P2_U5537, new_P2_U5538,
    new_P2_U5539, new_P2_U5540, new_P2_U5541, new_P2_U5542, new_P2_U5543,
    new_P2_U5544, new_P2_U5545, new_P2_U5546, new_P2_U5547, new_P2_U5548,
    new_P2_U5549, new_P2_U5550, new_P2_U5551, new_P2_U5552, new_P2_U5553,
    new_P2_U5554, new_P2_U5555, new_P2_U5556, new_P2_U5557, new_P2_U5558,
    new_P2_U5559, new_P2_U5560, new_P2_U5561, new_P2_U5562, new_P2_U5563,
    new_P2_U5564, new_P2_U5565, new_P2_U5566, new_P2_U5567, new_P2_U5568,
    new_P2_U5569, new_P2_U5570, new_P2_U5571, new_P2_U5572, new_P2_U5573,
    new_P2_U5574, new_P2_U5575, new_P2_U5576, new_P2_U5577, new_P2_U5578,
    new_P2_U5579, new_P2_U5580, new_P2_U5581, new_P2_U5582, new_P2_U5583,
    new_P2_U5584, new_P2_U5585, new_P2_U5586, new_P2_U5587, new_P2_U5588,
    new_P2_U5589, new_P2_U5590, new_P2_U5591, new_P2_U5592, new_P2_U5593,
    new_P2_U5594, new_P2_U5595, new_P2_U5596, new_P2_U5597, new_P2_U5598,
    new_P2_U5599, new_P2_U5600, new_P2_U5601, new_P2_U5602, new_P2_U5603,
    new_P2_U5604, new_P2_U5605, new_P2_U5606, new_P2_U5607, new_P2_U5608,
    new_P2_U5609, new_P2_U5610, new_P2_U5611, new_P2_U5612, new_P2_U5613,
    new_P2_U5614, new_P2_U5615, new_P2_U5616, new_P2_U5617, new_P2_U5618,
    new_P2_U5619, new_P2_U5620, new_P2_U5621, new_P2_U5622, new_P2_U5623,
    new_P2_U5624, new_P2_U5625, new_P2_U5626, new_P2_U5627, new_P2_U5628,
    new_P2_U5629, new_P2_U5630, new_P2_U5631, new_P2_U5632, new_P2_U5633,
    new_P2_U5634, new_P2_U5635, new_P2_U5636, new_P2_U5637, new_P2_U5638,
    new_P2_U5639, new_P2_U5640, new_P2_U5641, new_P2_U5642, new_P2_U5643,
    new_P2_U5644, new_P2_U5645, new_P2_U5646, new_P2_U5647, new_P2_U5648,
    new_P2_U5649, new_P2_U5650, new_P2_U5651, new_P2_U5652, new_P2_U5653,
    new_P2_U5654, new_P2_U5655, new_P2_U5656, new_P2_U5657, new_P2_U5658,
    new_P2_U5659, new_P2_U5660, new_P2_U5661, new_P2_U5662, new_P2_U5663,
    new_P2_U5664, new_P2_U5665, new_P2_U5666, new_P2_U5667, new_P2_U5668,
    new_P2_U5669, new_P2_U5670, new_P2_U5671, new_P2_U5672, new_P2_U5673,
    new_P2_U5674, new_P2_U5675, new_P2_U5676, new_P2_U5677, new_P2_U5678,
    new_P2_U5679, new_P2_U5680, new_P2_U5681, new_P2_U5682, new_P2_U5683,
    new_P2_U5684, new_P2_U5685, new_P2_U5686, new_P2_U5687, new_P2_U5688,
    new_P2_U5689, new_P2_U5690, new_P2_U5691, new_P2_U5692, new_P2_U5693,
    new_P2_U5694, new_P2_U5695, new_P2_U5696, new_P2_U5697, new_P2_U5698,
    new_P2_U5699, new_P2_U5700, new_P2_U5701, new_P2_U5702, new_P2_U5703,
    new_P2_U5704, new_P2_U5705, new_P2_U5706, new_P2_U5707, new_P2_U5708,
    new_P2_U5709, new_P2_U5710, new_P2_U5711, new_P2_U5712, new_P2_U5713,
    new_P2_U5714, new_P2_U5715, new_P2_U5716, new_P2_U5717, new_P2_U5718,
    new_P2_U5719, new_P2_U5720, new_P2_U5721, new_P2_U5722, new_P2_U5723,
    new_P2_U5724, new_P2_U5725, new_P2_U5726, new_P2_U5727, new_P2_U5728,
    new_P2_U5729, new_P2_U5730, new_P2_U5731, new_P2_U5732, new_P2_U5733,
    new_P2_U5734, new_P2_U5735, new_P2_U5736, new_P2_U5737, new_P2_U5738,
    new_P2_U5739, new_P2_U5740, new_P2_U5741, new_P2_U5742, new_P2_U5743,
    new_P2_U5744, new_P2_U5745, new_P2_U5746, new_P2_U5747, new_P2_U5748,
    new_P2_U5749, new_P2_U5750, new_P2_U5751, new_P2_U5752, new_P2_U5753,
    new_P2_U5754, new_P2_U5755, new_P2_U5756, new_P2_U5757, new_P2_U5758,
    new_P2_U5759, new_P2_U5760, new_P2_U5761, new_P2_U5762, new_P2_U5763,
    new_P2_U5764, new_P2_U5765, new_P2_U5766, new_P2_U5767, new_P2_U5768,
    new_P2_U5769, new_P2_U5770, new_P2_U5771, new_P2_U5772, new_P2_U5773,
    new_P2_U5774, new_P2_U5775, new_P2_U5776, new_P2_U5777, new_P2_U5778,
    new_P2_U5779, new_P2_U5780, new_P2_U5781, new_P2_U5782, new_P2_U5783,
    new_P2_U5784, new_P2_U5785, new_P2_U5786, new_P2_U5787, new_P2_U5788,
    new_P2_U5789, new_P2_U5790, new_P2_U5791, new_P2_U5792, new_P2_U5793,
    new_P2_U5794, new_P2_U5795, new_P2_U5796, new_P2_U5797, new_P2_U5798,
    new_P2_U5799, new_P2_U5800, new_P2_U5801, new_P2_U5802, new_P2_U5803,
    new_P2_U5804, new_P2_U5805, new_P2_U5806, new_P2_U5807, new_P2_U5808,
    new_P2_U5809, new_P2_U5810, new_P2_U5811, new_P2_U5812, new_P2_U5813,
    new_P2_U5814, new_P2_U5815, new_P2_U5816, new_P2_U5817, new_P2_U5818,
    new_P2_U5819, new_P2_U5820, new_P2_U5821, new_P2_U5822, new_P2_U5823,
    new_P2_U5824, new_P2_U5825, new_P2_U5826, new_P2_U5827, new_P2_U5828,
    new_P2_U5829, new_P2_U5830, new_P2_U5831, new_P2_U5832, new_P2_U5833,
    new_P2_U5834, new_P2_U5835, new_P2_U5836, new_P2_U5837, new_P2_U5838,
    new_P2_U5839, new_P2_U5840, new_P2_U5841, new_P2_U5842, new_P2_U5843,
    new_P2_U5844, new_P2_U5845, new_P2_U5846, new_P2_U5847, new_P2_U5848,
    new_P2_U5849, new_P2_U5850, new_P2_U5851, new_P2_U5852, new_P2_U5853,
    new_P2_U5854, new_P2_U5855, new_P2_U5856, new_P2_U5857, new_P2_U5858,
    new_P2_U5859, new_P2_U5860, new_P2_U5861, new_P2_U5862, new_P2_U5863,
    new_P2_U5864, new_P2_U5865, new_P2_U5866, new_P2_U5867, new_P2_U5868,
    new_P2_U5869, new_P2_U5870, new_P2_U5871, new_P2_U5872, new_P2_U5873,
    new_P2_U5874, new_P2_U5875, new_P2_U5876, new_P2_U5877, new_P2_U5878,
    new_P2_U5879, new_P2_U5880, new_P2_U5881, new_P2_U5882, new_P2_U5883,
    new_P2_U5884, new_P2_U5885, new_P2_U5886, new_P2_U5887, new_P2_U5888,
    new_P2_U5889, new_P2_U5890, new_P2_U5891, new_P2_U5892, new_P2_U5893,
    new_P2_U5894, new_P2_U5895, new_P2_U5896, new_P2_U5897, new_P2_U5898,
    new_P2_U5899, new_P2_U5900, new_P2_U5901, new_P2_U5902, new_P2_U5903,
    new_P2_U5904, new_P2_U5905, new_P2_U5906, new_P2_U5907, new_P2_U5908,
    new_P2_U5909, new_P2_U5910, new_P2_U5911, new_P2_U5912, new_P2_U5913,
    new_P2_U5914, new_P2_U5915, new_P2_U5916, new_P2_U5917, new_P2_U5918,
    new_P2_U5919, new_P2_U5920, new_P2_U5921, new_P2_U5922, new_P2_U5923,
    new_P2_U5924, new_P2_U5925, new_P2_U5926, new_P2_U5927, new_P2_U5928,
    new_P2_U5929, new_P2_U5930, new_P2_U5931, new_P2_U5932, new_P2_U5933,
    new_P2_U5934, new_P2_U5935, new_P2_U5936, new_P2_U5937, new_P2_U5938,
    new_P2_U5939, new_P2_U5940, new_P2_U5941, new_P2_U5942, new_P2_U5943,
    new_P2_U5944, new_P2_U5945, new_P2_U5946, new_P2_U5947, new_P2_U5948,
    new_P2_U5949, new_P2_U5950, new_P2_U5951, new_P2_U5952, new_P2_U5953,
    new_P2_U5954, new_P2_U5955, new_P2_U5956, new_P2_U5957, new_P2_U5958,
    new_P2_U5959, new_P2_U5960, new_P2_U5961, new_P2_U5962, new_P2_U5963,
    new_P2_U5964, new_P2_U5965, new_P2_U5966, new_P2_U5967, new_P2_U5968,
    new_P2_U5969, new_P2_U5970, new_P2_U5971, new_P2_U5972, new_P2_U5973,
    new_P2_U5974, new_P2_U5975, new_P2_U5976, new_P2_U5977, new_P2_U5978,
    new_P2_U5979, new_P2_U5980, new_P2_U5981, new_P2_U5982, new_P2_U5983,
    new_P2_U5984, new_P2_U5985, new_P2_U5986, new_P2_U5987, new_P2_U5988,
    new_P2_U5989, new_P2_U5990, new_P2_U5991, new_P2_U5992, new_P2_U5993,
    new_P2_U5994, new_P2_U5995, new_P2_U5996, new_P2_U5997, new_P2_U5998,
    new_P2_U5999, new_P2_U6000, new_P2_U6001, new_P2_U6002, new_P2_U6003,
    new_P2_U6004, new_P2_U6005, new_P2_U6006, new_P2_U6007, new_P2_U6008,
    new_P2_U6009, new_P2_U6010, new_P2_U6011, new_P2_U6012, new_P2_U6013,
    new_P2_U6014, new_P2_U6015, new_P2_U6016, new_P2_U6017, new_P2_U6018,
    new_P2_U6019, new_P2_U6020, new_P2_U6021, new_P2_U6022, new_P2_U6023,
    new_P2_U6024, new_P2_U6025, new_P2_U6026, new_P2_U6027, new_P2_U6028,
    new_P2_U6029, new_P2_U6030, new_P2_U6031, new_P2_U6032, new_P2_U6033,
    new_P2_U6034, new_P2_U6035, new_P2_U6036, new_P2_U6037, new_P2_U6038,
    new_P2_U6039, new_P2_U6040, new_P2_U6041, new_P2_U6042, new_P2_U6043,
    new_P2_U6044, new_P2_R1161_U465, new_P2_R1161_U464, new_P2_R1161_U463,
    new_P2_R1161_U462, new_P2_R1161_U461, new_P2_R1161_U460,
    new_P2_R1161_U459, new_P2_R1161_U458, new_P2_R1161_U457,
    new_P2_R1161_U456, new_P2_R1161_U455, new_P2_R1161_U454,
    new_P2_R1161_U453, new_P2_R1161_U452, new_P2_R1161_U451,
    new_P2_R1161_U450, new_P2_R1161_U449, new_P2_R1161_U448,
    new_P2_R1161_U447, new_LT_1075_U6, new_ADD_1068_U6, new_ADD_1068_U7,
    new_ADD_1068_U8, new_ADD_1068_U9, new_ADD_1068_U10, new_ADD_1068_U11,
    new_ADD_1068_U12, new_ADD_1068_U13, new_ADD_1068_U14, new_ADD_1068_U15,
    new_ADD_1068_U16, new_ADD_1068_U17, new_ADD_1068_U18, new_ADD_1068_U19,
    new_ADD_1068_U20, new_ADD_1068_U21, new_ADD_1068_U22, new_ADD_1068_U23,
    new_ADD_1068_U24, new_ADD_1068_U25, new_ADD_1068_U26, new_ADD_1068_U27,
    new_ADD_1068_U28, new_ADD_1068_U29, new_ADD_1068_U30, new_ADD_1068_U31,
    new_ADD_1068_U32, new_ADD_1068_U33, new_ADD_1068_U34, new_ADD_1068_U35,
    new_ADD_1068_U36, new_ADD_1068_U37, new_ADD_1068_U38, new_ADD_1068_U39,
    new_ADD_1068_U40, new_ADD_1068_U41, new_ADD_1068_U42, new_ADD_1068_U43,
    new_ADD_1068_U44, new_ADD_1068_U45, new_ADD_1068_U64, new_ADD_1068_U65,
    new_ADD_1068_U66, new_ADD_1068_U67, new_ADD_1068_U68, new_ADD_1068_U69,
    new_ADD_1068_U70, new_ADD_1068_U71, new_ADD_1068_U72, new_ADD_1068_U73,
    new_ADD_1068_U74, new_ADD_1068_U75, new_ADD_1068_U76, new_ADD_1068_U77,
    new_ADD_1068_U78, new_ADD_1068_U79, new_ADD_1068_U80, new_ADD_1068_U81,
    new_ADD_1068_U82, new_ADD_1068_U83, new_ADD_1068_U84, new_ADD_1068_U85,
    new_ADD_1068_U86, new_ADD_1068_U87, new_ADD_1068_U88, new_ADD_1068_U89,
    new_ADD_1068_U90, new_ADD_1068_U91, new_ADD_1068_U92, new_ADD_1068_U93,
    new_ADD_1068_U94, new_ADD_1068_U95, new_ADD_1068_U96, new_ADD_1068_U97,
    new_ADD_1068_U98, new_ADD_1068_U99, new_ADD_1068_U100,
    new_ADD_1068_U101, new_ADD_1068_U102, new_ADD_1068_U103,
    new_ADD_1068_U104, new_ADD_1068_U105, new_ADD_1068_U106,
    new_ADD_1068_U107, new_ADD_1068_U108, new_ADD_1068_U109,
    new_ADD_1068_U110, new_ADD_1068_U111, new_ADD_1068_U112,
    new_ADD_1068_U113, new_ADD_1068_U114, new_ADD_1068_U115,
    new_ADD_1068_U116, new_ADD_1068_U117, new_ADD_1068_U118,
    new_ADD_1068_U119, new_ADD_1068_U120, new_ADD_1068_U121,
    new_ADD_1068_U122, new_ADD_1068_U123, new_ADD_1068_U124,
    new_ADD_1068_U125, new_ADD_1068_U126, new_ADD_1068_U127,
    new_ADD_1068_U128, new_ADD_1068_U129, new_ADD_1068_U130,
    new_ADD_1068_U131, new_ADD_1068_U132, new_ADD_1068_U133,
    new_ADD_1068_U134, new_ADD_1068_U135, new_ADD_1068_U136,
    new_ADD_1068_U137, new_ADD_1068_U138, new_ADD_1068_U139,
    new_ADD_1068_U140, new_ADD_1068_U141, new_ADD_1068_U142,
    new_ADD_1068_U143, new_ADD_1068_U144, new_ADD_1068_U145,
    new_ADD_1068_U146, new_ADD_1068_U147, new_ADD_1068_U148,
    new_ADD_1068_U149, new_ADD_1068_U150, new_ADD_1068_U151,
    new_ADD_1068_U152, new_ADD_1068_U153, new_ADD_1068_U154,
    new_ADD_1068_U155, new_ADD_1068_U156, new_ADD_1068_U157,
    new_ADD_1068_U158, new_ADD_1068_U159, new_ADD_1068_U160,
    new_ADD_1068_U161, new_ADD_1068_U162, new_ADD_1068_U163,
    new_ADD_1068_U164, new_ADD_1068_U165, new_ADD_1068_U166,
    new_ADD_1068_U167, new_ADD_1068_U168, new_ADD_1068_U169,
    new_ADD_1068_U170, new_ADD_1068_U171, new_ADD_1068_U172,
    new_ADD_1068_U173, new_ADD_1068_U174, new_ADD_1068_U175,
    new_ADD_1068_U176, new_ADD_1068_U177, new_ADD_1068_U178,
    new_ADD_1068_U179, new_ADD_1068_U180, new_ADD_1068_U181,
    new_ADD_1068_U182, new_ADD_1068_U183, new_ADD_1068_U184,
    new_ADD_1068_U185, new_ADD_1068_U186, new_ADD_1068_U187,
    new_ADD_1068_U188, new_ADD_1068_U189, new_ADD_1068_U190,
    new_ADD_1068_U191, new_ADD_1068_U192, new_ADD_1068_U193,
    new_ADD_1068_U194, new_ADD_1068_U195, new_ADD_1068_U196,
    new_ADD_1068_U197, new_ADD_1068_U198, new_ADD_1068_U199,
    new_ADD_1068_U200, new_ADD_1068_U201, new_ADD_1068_U202,
    new_ADD_1068_U203, new_ADD_1068_U204, new_ADD_1068_U205,
    new_ADD_1068_U206, new_ADD_1068_U207, new_ADD_1068_U208,
    new_ADD_1068_U209, new_ADD_1068_U210, new_ADD_1068_U211,
    new_ADD_1068_U212, new_ADD_1068_U213, new_ADD_1068_U214,
    new_ADD_1068_U215, new_ADD_1068_U216, new_ADD_1068_U217,
    new_ADD_1068_U218, new_ADD_1068_U219, new_ADD_1068_U220,
    new_ADD_1068_U221, new_ADD_1068_U222, new_ADD_1068_U223,
    new_ADD_1068_U224, new_ADD_1068_U225, new_ADD_1068_U226,
    new_ADD_1068_U227, new_ADD_1068_U228, new_ADD_1068_U229,
    new_ADD_1068_U230, new_ADD_1068_U231, new_ADD_1068_U232,
    new_ADD_1068_U233, new_ADD_1068_U234, new_ADD_1068_U235,
    new_ADD_1068_U236, new_ADD_1068_U237, new_ADD_1068_U238,
    new_ADD_1068_U239, new_ADD_1068_U240, new_ADD_1068_U241,
    new_ADD_1068_U242, new_ADD_1068_U243, new_ADD_1068_U244,
    new_ADD_1068_U245, new_ADD_1068_U246, new_ADD_1068_U247,
    new_ADD_1068_U248, new_ADD_1068_U249, new_ADD_1068_U250,
    new_ADD_1068_U251, new_ADD_1068_U252, new_ADD_1068_U253,
    new_ADD_1068_U254, new_ADD_1068_U255, new_ADD_1068_U256,
    new_ADD_1068_U257, new_ADD_1068_U258, new_ADD_1068_U259,
    new_ADD_1068_U260, new_ADD_1068_U261, new_ADD_1068_U262,
    new_ADD_1068_U263, new_ADD_1068_U264, new_ADD_1068_U265,
    new_ADD_1068_U266, new_ADD_1068_U267, new_ADD_1068_U268,
    new_ADD_1068_U269, new_ADD_1068_U270, new_ADD_1068_U271,
    new_ADD_1068_U272, new_ADD_1068_U273, new_ADD_1068_U274,
    new_ADD_1068_U275, new_ADD_1068_U276, new_ADD_1068_U277,
    new_ADD_1068_U278, new_ADD_1068_U279, new_ADD_1068_U280,
    new_ADD_1068_U281, new_ADD_1068_U282, new_ADD_1068_U283,
    new_ADD_1068_U284, new_ADD_1068_U285, new_ADD_1068_U286,
    new_ADD_1068_U287, new_ADD_1068_U288, new_ADD_1068_U289,
    new_ADD_1068_U290, new_ADD_1068_U291, new_R140_U4, new_R140_U5,
    new_R140_U6, new_R140_U7, new_R140_U8, new_R140_U9, new_R140_U10,
    new_R140_U11, new_R140_U12, new_R140_U13, new_R140_U14, new_R140_U15,
    new_R140_U16, new_R140_U17, new_R140_U18, new_R140_U19, new_R140_U20,
    new_R140_U21, new_R140_U22, new_R140_U23, new_R140_U24, new_R140_U25,
    new_R140_U26, new_R140_U27, new_R140_U28, new_R140_U29, new_R140_U30,
    new_R140_U31, new_R140_U32, new_R140_U33, new_R140_U34, new_R140_U35,
    new_R140_U36, new_R140_U37, new_R140_U38, new_R140_U39, new_R140_U40,
    new_R140_U41, new_R140_U42, new_R140_U43, new_R140_U44, new_R140_U45,
    new_R140_U46, new_R140_U47, new_R140_U48, new_R140_U49, new_R140_U50,
    new_R140_U51, new_R140_U52, new_R140_U53, new_R140_U54, new_R140_U55,
    new_R140_U56, new_R140_U57, new_R140_U58, new_R140_U59, new_R140_U60,
    new_R140_U61, new_R140_U62, new_R140_U63, new_R140_U64, new_R140_U65,
    new_R140_U66, new_R140_U67, new_R140_U68, new_R140_U69, new_R140_U70,
    new_R140_U71, new_R140_U72, new_R140_U73, new_R140_U74, new_R140_U75,
    new_R140_U76, new_R140_U77, new_R140_U78, new_R140_U79, new_R140_U80,
    new_R140_U81, new_R140_U82, new_R140_U83, new_R140_U84, new_R140_U85,
    new_R140_U86, new_R140_U87, new_R140_U88, new_R140_U89, new_R140_U90,
    new_R140_U91, new_R140_U92, new_R140_U93, new_R140_U94, new_R140_U95,
    new_R140_U96, new_R140_U97, new_R140_U98, new_R140_U99, new_R140_U100,
    new_R140_U101, new_R140_U102, new_R140_U103, new_R140_U104,
    new_R140_U105, new_R140_U106, new_R140_U107, new_R140_U108,
    new_R140_U109, new_R140_U110, new_R140_U111, new_R140_U112,
    new_R140_U113, new_R140_U114, new_R140_U115, new_R140_U116,
    new_R140_U117, new_R140_U118, new_R140_U119, new_R140_U120,
    new_R140_U121, new_R140_U122, new_R140_U123, new_R140_U124,
    new_R140_U125, new_R140_U126, new_R140_U127, new_R140_U128,
    new_R140_U129, new_R140_U130, new_R140_U131, new_R140_U132,
    new_R140_U133, new_R140_U134, new_R140_U135, new_R140_U136,
    new_R140_U137, new_R140_U138, new_R140_U139, new_R140_U140,
    new_R140_U141, new_R140_U142, new_R140_U143, new_R140_U144,
    new_R140_U145, new_R140_U146, new_R140_U147, new_R140_U148,
    new_R140_U149, new_R140_U150, new_R140_U151, new_R140_U152,
    new_R140_U153, new_R140_U154, new_R140_U155, new_R140_U156,
    new_R140_U157, new_R140_U158, new_R140_U159, new_R140_U160,
    new_R140_U161, new_R140_U162, new_R140_U163, new_R140_U164,
    new_R140_U165, new_R140_U166, new_R140_U167, new_R140_U168,
    new_R140_U169, new_R140_U170, new_R140_U171, new_R140_U172,
    new_R140_U173, new_R140_U174, new_R140_U175, new_R140_U176,
    new_R140_U177, new_R140_U178, new_R140_U179, new_R140_U180,
    new_R140_U181, new_R140_U182, new_R140_U183, new_R140_U184,
    new_R140_U185, new_R140_U186, new_R140_U187, new_R140_U188,
    new_R140_U189, new_R140_U190, new_R140_U191, new_R140_U192,
    new_R140_U193, new_R140_U194, new_R140_U195, new_R140_U196,
    new_R140_U197, new_R140_U198, new_R140_U199, new_R140_U200,
    new_R140_U201, new_R140_U202, new_R140_U203, new_R140_U204,
    new_R140_U205, new_R140_U206, new_R140_U207, new_R140_U208,
    new_R140_U209, new_R140_U210, new_R140_U211, new_R140_U212,
    new_R140_U213, new_R140_U214, new_R140_U215, new_R140_U216,
    new_R140_U217, new_R140_U218, new_R140_U219, new_R140_U220,
    new_R140_U221, new_R140_U222, new_R140_U223, new_R140_U224,
    new_R140_U225, new_R140_U226, new_R140_U227, new_R140_U228,
    new_R140_U229, new_R140_U230, new_R140_U231, new_R140_U232,
    new_R140_U233, new_R140_U234, new_R140_U235, new_R140_U236,
    new_R140_U237, new_R140_U238, new_R140_U239, new_R140_U240,
    new_R140_U241, new_R140_U242, new_R140_U243, new_R140_U244,
    new_R140_U245, new_R140_U246, new_R140_U247, new_R140_U248,
    new_R140_U249, new_R140_U250, new_R140_U251, new_R140_U252,
    new_R140_U253, new_R140_U254, new_R140_U255, new_R140_U256,
    new_R140_U257, new_R140_U258, new_R140_U259, new_R140_U260,
    new_R140_U261, new_R140_U262, new_R140_U263, new_R140_U264,
    new_R140_U265, new_R140_U266, new_R140_U267, new_R140_U268,
    new_R140_U269, new_R140_U270, new_R140_U271, new_R140_U272,
    new_R140_U273, new_R140_U274, new_R140_U275, new_R140_U276,
    new_R140_U277, new_R140_U278, new_R140_U279, new_R140_U280,
    new_R140_U281, new_R140_U282, new_R140_U283, new_R140_U284,
    new_R140_U285, new_R140_U286, new_R140_U287, new_R140_U288,
    new_R140_U289, new_R140_U290, new_R140_U291, new_R140_U292,
    new_R140_U293, new_R140_U294, new_R140_U295, new_R140_U296,
    new_R140_U297, new_R140_U298, new_R140_U299, new_R140_U300,
    new_R140_U301, new_R140_U302, new_R140_U303, new_R140_U304,
    new_R140_U305, new_R140_U306, new_R140_U307, new_R140_U308,
    new_R140_U309, new_R140_U310, new_R140_U311, new_R140_U312,
    new_R140_U313, new_R140_U314, new_R140_U315, new_R140_U316,
    new_R140_U317, new_R140_U318, new_R140_U319, new_R140_U320,
    new_R140_U321, new_R140_U322, new_R140_U323, new_R140_U324,
    new_R140_U325, new_R140_U326, new_R140_U327, new_R140_U328,
    new_R140_U329, new_R140_U330, new_R140_U331, new_R140_U332,
    new_R140_U333, new_R140_U334, new_R140_U335, new_R140_U336,
    new_R140_U337, new_R140_U338, new_R140_U339, new_R140_U340,
    new_R140_U341, new_R140_U342, new_R140_U343, new_R140_U344,
    new_R140_U345, new_R140_U346, new_R140_U347, new_R140_U348,
    new_R140_U349, new_R140_U350, new_R140_U351, new_R140_U352,
    new_R140_U353, new_R140_U354, new_R140_U355, new_R140_U356,
    new_R140_U357, new_R140_U358, new_R140_U359, new_R140_U360,
    new_R140_U361, new_R140_U362, new_R140_U363, new_R140_U364,
    new_R140_U365, new_R140_U366, new_R140_U367, new_R140_U368,
    new_R140_U369, new_R140_U370, new_R140_U371, new_R140_U372,
    new_R140_U373, new_R140_U374, new_R140_U375, new_R140_U376,
    new_R140_U377, new_R140_U378, new_R140_U379, new_R140_U380,
    new_R140_U381, new_R140_U382, new_R140_U383, new_R140_U384,
    new_R140_U385, new_R140_U386, new_R140_U387, new_R140_U388,
    new_R140_U389, new_R140_U390, new_R140_U391, new_R140_U392,
    new_R140_U393, new_R140_U394, new_R140_U395, new_R140_U396,
    new_R140_U397, new_R140_U398, new_R140_U399, new_R140_U400,
    new_R140_U401, new_R140_U402, new_R140_U403, new_R140_U404,
    new_R140_U405, new_R140_U406, new_R140_U407, new_R140_U408,
    new_R140_U409, new_R140_U410, new_R140_U411, new_R140_U412,
    new_R140_U413, new_R140_U414, new_R140_U415, new_R140_U416,
    new_R140_U417, new_R140_U418, new_R140_U419, new_R140_U420,
    new_R140_U421, new_R140_U422, new_R140_U423, new_R140_U424,
    new_R140_U425, new_R140_U426, new_R140_U427, new_R140_U428,
    new_R140_U429, new_R140_U430, new_R140_U431, new_R140_U432,
    new_R140_U433, new_R140_U434, new_R140_U435, new_R140_U436,
    new_R140_U437, new_R140_U438, new_R140_U439, new_R140_U440,
    new_R140_U441, new_R140_U442, new_R140_U443, new_R140_U444,
    new_R140_U445, new_R140_U446, new_R140_U447, new_R140_U448,
    new_R140_U449, new_R140_U450, new_R140_U451, new_R140_U452,
    new_R140_U453, new_R140_U454, new_R140_U455, new_R140_U456,
    new_R140_U457, new_R140_U458, new_R140_U459, new_R140_U460,
    new_R140_U461, new_R140_U462, new_R140_U463, new_R140_U464,
    new_R140_U465, new_R140_U466, new_R140_U467, new_R140_U468,
    new_R140_U469, new_R140_U470, new_R140_U471, new_R140_U472,
    new_R140_U473, new_R140_U474, new_R140_U475, new_R140_U476,
    new_R140_U477, new_R140_U478, new_R140_U479, new_R140_U480,
    new_R140_U481, new_R140_U482, new_R140_U483, new_R140_U484,
    new_R140_U485, new_R140_U486, new_R140_U487, new_R140_U488,
    new_R140_U489, new_R140_U490, new_R140_U491, new_R140_U492,
    new_R140_U493, new_R140_U494, new_R140_U495, new_R140_U496,
    new_R140_U497, new_R140_U498, new_R140_U499, new_R140_U500,
    new_R140_U501, new_R140_U502, new_R140_U503, new_R140_U504,
    new_R140_U505, new_R140_U506, new_R140_U507, new_R140_U508,
    new_R140_U509, new_R140_U510, new_R140_U511, new_R140_U512,
    new_R140_U513, new_R140_U514, new_R140_U515, new_R140_U516,
    new_R140_U517, new_R140_U518, new_R140_U519, new_R140_U520,
    new_R140_U521, new_R140_U522, new_R140_U523, new_R140_U524,
    new_R140_U525, new_R140_U526, new_R140_U527, new_R140_U528,
    new_R140_U529, new_R140_U530, new_R140_U531, new_R140_U532,
    new_R140_U533, new_R140_U534, new_R140_U535, new_R140_U536,
    new_R140_U537, new_R140_U538, new_R140_U539, new_R140_U540,
    new_R140_U541, new_LT_1075_19_U6, new_P1_ADD_95_U4, new_P1_ADD_95_U5,
    new_P1_ADD_95_U6, new_P1_ADD_95_U7, new_P1_ADD_95_U8, new_P1_ADD_95_U9,
    new_P1_ADD_95_U10, new_P1_ADD_95_U11, new_P1_ADD_95_U12,
    new_P1_ADD_95_U13, new_P1_ADD_95_U14, new_P1_ADD_95_U15,
    new_P1_ADD_95_U16, new_P1_ADD_95_U17, new_P1_ADD_95_U18,
    new_P1_ADD_95_U19, new_P1_ADD_95_U20, new_P1_ADD_95_U21,
    new_P1_ADD_95_U22, new_P1_ADD_95_U23, new_P1_ADD_95_U24,
    new_P1_ADD_95_U25, new_P1_ADD_95_U26, new_P1_ADD_95_U27,
    new_P1_ADD_95_U28, new_P1_ADD_95_U29, new_P1_ADD_95_U30,
    new_P1_ADD_95_U31, new_P1_ADD_95_U32, new_P1_ADD_95_U33,
    new_P1_ADD_95_U34, new_P1_ADD_95_U35, new_P1_ADD_95_U36,
    new_P1_ADD_95_U37, new_P1_ADD_95_U38, new_P1_ADD_95_U39,
    new_P1_ADD_95_U40, new_P1_ADD_95_U41, new_P1_ADD_95_U42,
    new_P1_ADD_95_U43, new_P1_ADD_95_U44, new_P1_ADD_95_U45,
    new_P1_ADD_95_U46, new_P1_ADD_95_U47, new_P1_ADD_95_U48,
    new_P1_ADD_95_U49, new_P1_ADD_95_U50, new_P1_ADD_95_U51,
    new_P1_ADD_95_U52, new_P1_ADD_95_U53, new_P1_ADD_95_U54,
    new_P1_ADD_95_U55, new_P1_ADD_95_U56, new_P1_ADD_95_U57,
    new_P1_ADD_95_U58, new_P1_ADD_95_U59, new_P1_ADD_95_U60,
    new_P1_ADD_95_U61, new_P1_ADD_95_U62, new_P1_ADD_95_U63,
    new_P1_ADD_95_U64, new_P1_ADD_95_U65, new_P1_ADD_95_U66,
    new_P1_ADD_95_U67, new_P1_ADD_95_U68, new_P1_ADD_95_U69,
    new_P1_ADD_95_U70, new_P1_ADD_95_U71, new_P1_ADD_95_U72,
    new_P1_ADD_95_U73, new_P1_ADD_95_U74, new_P1_ADD_95_U75,
    new_P1_ADD_95_U76, new_P1_ADD_95_U77, new_P1_ADD_95_U78,
    new_P1_ADD_95_U79, new_P1_ADD_95_U80, new_P1_ADD_95_U81,
    new_P1_ADD_95_U82, new_P1_ADD_95_U83, new_P1_ADD_95_U84,
    new_P1_ADD_95_U85, new_P1_ADD_95_U86, new_P1_ADD_95_U87,
    new_P1_ADD_95_U88, new_P1_ADD_95_U89, new_P1_ADD_95_U90,
    new_P1_ADD_95_U91, new_P1_ADD_95_U92, new_P1_ADD_95_U93,
    new_P1_ADD_95_U94, new_P1_ADD_95_U95, new_P1_ADD_95_U96,
    new_P1_ADD_95_U97, new_P1_ADD_95_U98, new_P1_ADD_95_U99,
    new_P1_ADD_95_U100, new_P1_ADD_95_U101, new_P1_ADD_95_U102,
    new_P1_ADD_95_U103, new_P1_ADD_95_U104, new_P1_ADD_95_U105,
    new_P1_ADD_95_U106, new_P1_ADD_95_U107, new_P1_ADD_95_U108,
    new_P1_ADD_95_U109, new_P1_ADD_95_U110, new_P1_ADD_95_U111,
    new_P1_ADD_95_U112, new_P1_ADD_95_U113, new_P1_ADD_95_U114,
    new_P1_ADD_95_U115, new_P1_ADD_95_U116, new_P1_ADD_95_U117,
    new_P1_ADD_95_U118, new_P1_ADD_95_U119, new_P1_ADD_95_U120,
    new_P1_ADD_95_U121, new_P1_ADD_95_U122, new_P1_ADD_95_U123,
    new_P1_ADD_95_U124, new_P1_ADD_95_U125, new_P1_ADD_95_U126,
    new_P1_ADD_95_U127, new_P1_ADD_95_U128, new_P1_ADD_95_U129,
    new_P1_ADD_95_U130, new_P1_ADD_95_U131, new_P1_ADD_95_U132,
    new_P1_ADD_95_U133, new_P1_ADD_95_U134, new_P1_ADD_95_U135,
    new_P1_ADD_95_U136, new_P1_ADD_95_U137, new_P1_ADD_95_U138,
    new_P1_ADD_95_U139, new_P1_ADD_95_U140, new_P1_ADD_95_U141,
    new_P1_ADD_95_U142, new_P1_ADD_95_U143, new_P1_ADD_95_U144,
    new_P1_ADD_95_U145, new_P1_ADD_95_U146, new_P1_ADD_95_U147,
    new_P1_ADD_95_U148, new_P1_ADD_95_U149, new_P1_ADD_95_U150,
    new_P1_ADD_95_U151, new_P1_ADD_95_U152, new_P1_ADD_95_U153,
    new_P1_R1105_U4, new_P1_R1105_U5, new_P1_R1105_U6, new_P1_R1105_U7,
    new_P1_R1105_U8, new_P1_R1105_U9, new_P1_R1105_U10, new_P1_R1105_U11,
    new_P1_R1105_U12, new_P1_R1105_U13, new_P1_R1105_U14, new_P1_R1105_U15,
    new_P1_R1105_U16, new_P1_R1105_U17, new_P1_R1105_U18, new_P1_R1105_U19,
    new_P1_R1105_U20, new_P1_R1105_U21, new_P1_R1105_U22, new_P1_R1105_U23,
    new_P1_R1105_U24, new_P1_R1105_U25, new_P1_R1105_U26, new_P1_R1105_U27,
    new_P1_R1105_U28, new_P1_R1105_U29, new_P1_R1105_U30, new_P1_R1105_U31,
    new_P1_R1105_U32, new_P1_R1105_U33, new_P1_R1105_U34, new_P1_R1105_U35,
    new_P1_R1105_U36, new_P1_R1105_U37, new_P1_R1105_U38, new_P1_R1105_U39,
    new_P1_R1105_U40, new_P1_R1105_U41, new_P1_R1105_U42, new_P1_R1105_U43,
    new_P1_R1105_U44, new_P1_R1105_U45, new_P1_R1105_U46, new_P1_R1105_U47,
    new_P1_R1105_U48, new_P1_R1105_U49, new_P1_R1105_U50, new_P1_R1105_U51,
    new_P1_R1105_U52, new_P1_R1105_U53, new_P1_R1105_U54, new_P1_R1105_U55,
    new_P1_R1105_U56, new_P1_R1105_U57, new_P1_R1105_U58, new_P1_R1105_U59,
    new_P1_R1105_U60, new_P1_R1105_U61, new_P1_R1105_U62, new_P1_R1105_U63,
    new_P1_R1105_U64, new_P1_R1105_U65, new_P1_R1105_U66, new_P1_R1105_U67,
    new_P1_R1105_U68, new_P1_R1105_U69, new_P1_R1105_U70, new_P1_R1105_U71,
    new_P1_R1105_U72, new_P1_R1105_U73, new_P1_R1105_U74, new_P1_R1105_U75,
    new_P1_R1105_U76, new_P1_R1105_U77, new_P1_R1105_U78, new_P1_R1105_U79,
    new_P1_R1105_U80, new_P1_R1105_U81, new_P1_R1105_U82, new_P1_R1105_U83,
    new_P1_R1105_U84, new_P1_R1105_U85, new_P1_R1105_U86, new_P1_R1105_U87,
    new_P1_R1105_U88, new_P1_R1105_U89, new_P1_R1105_U90, new_P1_R1105_U91,
    new_P1_R1105_U92, new_P1_R1105_U93, new_P1_R1105_U94, new_P1_R1105_U95,
    new_P1_R1105_U96, new_P1_R1105_U97, new_P1_R1105_U98, new_P1_R1105_U99,
    new_P1_R1105_U100, new_P1_R1105_U101, new_P1_R1105_U102,
    new_P1_R1105_U103, new_P1_R1105_U104, new_P1_R1105_U105,
    new_P1_R1105_U106, new_P1_R1105_U107, new_P1_R1105_U108,
    new_P1_R1105_U109, new_P1_R1105_U110, new_P1_R1105_U111,
    new_P1_R1105_U112, new_P1_R1105_U113, new_P1_R1105_U114,
    new_P1_R1105_U115, new_P1_R1105_U116, new_P1_R1105_U117,
    new_P1_R1105_U118, new_P1_R1105_U119, new_P1_R1105_U120,
    new_P1_R1105_U121, new_P1_R1105_U122, new_P1_R1105_U123,
    new_P1_R1105_U124, new_P1_R1105_U125, new_P1_R1105_U126,
    new_P1_R1105_U127, new_P1_R1105_U128, new_P1_R1105_U129,
    new_P1_R1105_U130, new_P1_R1105_U131, new_P1_R1105_U132,
    new_P1_R1105_U133, new_P1_R1105_U134, new_P1_R1105_U135,
    new_P1_R1105_U136, new_P1_R1105_U137, new_P1_R1105_U138,
    new_P1_R1105_U139, new_P1_R1105_U140, new_P1_R1105_U141,
    new_P1_R1105_U142, new_P1_R1105_U143, new_P1_R1105_U144,
    new_P1_R1105_U145, new_P1_R1105_U146, new_P1_R1105_U147,
    new_P1_R1105_U148, new_P1_R1105_U149, new_P1_R1105_U150,
    new_P1_R1105_U151, new_P1_R1105_U152, new_P1_R1105_U153,
    new_P1_R1105_U154, new_P1_R1105_U155, new_P1_R1105_U156,
    new_P1_R1105_U157, new_P1_R1105_U158, new_P1_R1105_U159,
    new_P1_R1105_U160, new_P1_R1105_U161, new_P1_R1105_U162,
    new_P1_R1105_U163, new_P1_R1105_U164, new_P1_R1105_U165,
    new_P1_R1105_U166, new_P1_R1105_U167, new_P1_R1105_U168,
    new_P1_R1105_U169, new_P1_R1105_U170, new_P1_R1105_U171,
    new_P1_R1105_U172, new_P1_R1105_U173, new_P1_R1105_U174,
    new_P1_R1105_U175, new_P1_R1105_U176, new_P1_R1105_U177,
    new_P1_R1105_U178, new_P1_R1105_U179, new_P1_R1105_U180,
    new_P1_R1105_U181, new_P1_R1105_U182, new_P1_R1105_U183,
    new_P1_R1105_U184, new_P1_R1105_U185, new_P1_R1105_U186,
    new_P1_R1105_U187, new_P1_R1105_U188, new_P1_R1105_U189,
    new_P1_R1105_U190, new_P1_R1105_U191, new_P1_R1105_U192,
    new_P1_R1105_U193, new_P1_R1105_U194, new_P1_R1105_U195,
    new_P1_R1105_U196, new_P1_R1105_U197, new_P1_R1105_U198,
    new_P1_R1105_U199, new_P1_R1105_U200, new_P1_R1105_U201,
    new_P1_R1105_U202, new_P1_R1105_U203, new_P1_R1105_U204,
    new_P1_R1105_U205, new_P1_R1105_U206, new_P1_R1105_U207,
    new_P1_R1105_U208, new_P1_R1105_U209, new_P1_R1105_U210,
    new_P1_R1105_U211, new_P1_R1105_U212, new_P1_R1105_U213,
    new_P1_R1105_U214, new_P1_R1105_U215, new_P1_R1105_U216,
    new_P1_R1105_U217, new_P1_R1105_U218, new_P1_R1105_U219,
    new_P1_R1105_U220, new_P1_R1105_U221, new_P1_R1105_U222,
    new_P1_R1105_U223, new_P1_R1105_U224, new_P1_R1105_U225,
    new_P1_R1105_U226, new_P1_R1105_U227, new_P1_R1105_U228,
    new_P1_R1105_U229, new_P1_R1105_U230, new_P1_R1105_U231,
    new_P1_R1105_U232, new_P1_R1105_U233, new_P1_R1105_U234,
    new_P1_R1105_U235, new_P1_R1105_U236, new_P1_R1105_U237,
    new_P1_R1105_U238, new_P1_R1105_U239, new_P1_R1105_U240,
    new_P1_R1105_U241, new_P1_R1105_U242, new_P1_R1105_U243,
    new_P1_R1105_U244, new_P1_R1105_U245, new_P1_R1105_U246,
    new_P1_R1105_U247, new_P1_R1105_U248, new_P1_R1105_U249,
    new_P1_R1105_U250, new_P1_R1105_U251, new_P1_R1105_U252,
    new_P1_R1105_U253, new_P1_R1105_U254, new_P1_R1105_U255,
    new_P1_R1105_U256, new_P1_R1105_U257, new_P1_R1105_U258,
    new_P1_R1105_U259, new_P1_R1105_U260, new_P1_R1105_U261,
    new_P1_R1105_U262, new_P1_R1105_U263, new_P1_R1105_U264,
    new_P1_R1105_U265, new_P1_R1105_U266, new_P1_R1105_U267,
    new_P1_R1105_U268, new_P1_R1105_U269, new_P1_R1105_U270,
    new_P1_R1105_U271, new_P1_R1105_U272, new_P1_R1105_U273,
    new_P1_R1105_U274, new_P1_R1105_U275, new_P1_R1105_U276,
    new_P1_R1105_U277, new_P1_R1105_U278, new_P1_R1105_U279,
    new_P1_R1105_U280, new_P1_R1105_U281, new_P1_R1105_U282,
    new_P1_R1105_U283, new_P1_R1105_U284, new_P1_R1105_U285,
    new_P1_R1105_U286, new_P1_R1105_U287, new_P1_R1105_U288,
    new_P1_R1105_U289, new_P1_R1105_U290, new_P1_R1105_U291,
    new_P1_R1105_U292, new_P1_R1105_U293, new_P1_R1105_U294,
    new_P1_R1105_U295, new_P1_R1105_U296, new_P1_R1105_U297,
    new_P1_R1105_U298, new_P1_R1105_U299, new_P1_R1105_U300,
    new_P1_R1105_U301, new_P1_R1105_U302, new_P1_R1105_U303,
    new_P1_R1105_U304, new_P1_R1105_U305, new_P1_R1105_U306,
    new_P1_R1105_U307, new_P1_R1105_U308, new_P1_SUB_84_U6,
    new_P1_SUB_84_U7, new_P1_SUB_84_U8, new_P1_SUB_84_U9,
    new_P1_SUB_84_U10, new_P1_SUB_84_U11, new_P1_SUB_84_U12,
    new_P1_SUB_84_U13, new_P1_SUB_84_U14, new_P1_SUB_84_U15,
    new_P1_SUB_84_U16, new_P1_SUB_84_U17, new_P1_SUB_84_U18,
    new_P1_SUB_84_U19, new_P1_SUB_84_U20, new_P1_SUB_84_U21,
    new_P1_SUB_84_U22, new_P1_SUB_84_U23, new_P1_SUB_84_U24,
    new_P1_SUB_84_U25, new_P1_SUB_84_U26, new_P1_SUB_84_U27,
    new_P1_SUB_84_U28, new_P1_SUB_84_U29, new_P1_SUB_84_U30,
    new_P1_SUB_84_U31, new_P1_SUB_84_U32, new_P1_SUB_84_U33,
    new_P1_SUB_84_U34, new_P1_SUB_84_U35, new_P1_SUB_84_U36,
    new_P1_SUB_84_U37, new_P1_SUB_84_U38, new_P1_SUB_84_U39,
    new_P1_SUB_84_U40, new_P1_SUB_84_U41, new_P1_SUB_84_U42,
    new_P1_SUB_84_U43, new_P1_SUB_84_U44, new_P1_SUB_84_U45,
    new_P1_SUB_84_U46, new_P1_SUB_84_U47, new_P1_SUB_84_U48,
    new_P1_SUB_84_U49, new_P1_SUB_84_U50, new_P1_SUB_84_U51,
    new_P1_SUB_84_U52, new_P1_SUB_84_U53, new_P1_SUB_84_U54,
    new_P1_SUB_84_U55, new_P1_SUB_84_U56, new_P1_SUB_84_U57,
    new_P1_SUB_84_U58, new_P1_SUB_84_U59, new_P1_SUB_84_U60,
    new_P1_SUB_84_U61, new_P1_SUB_84_U62, new_P1_SUB_84_U63,
    new_P1_SUB_84_U64, new_P1_SUB_84_U65, new_P1_SUB_84_U66,
    new_P1_SUB_84_U67, new_P1_SUB_84_U68, new_P1_SUB_84_U69,
    new_P1_SUB_84_U70, new_P1_SUB_84_U71, new_P1_SUB_84_U72,
    new_P1_SUB_84_U73, new_P1_SUB_84_U74, new_P1_SUB_84_U75,
    new_P1_SUB_84_U76, new_P1_SUB_84_U77, new_P1_SUB_84_U78,
    new_P1_SUB_84_U79, new_P1_SUB_84_U80, new_P1_SUB_84_U81,
    new_P1_SUB_84_U82, new_P1_SUB_84_U83, new_P1_SUB_84_U84,
    new_P1_SUB_84_U85, new_P1_SUB_84_U86, new_P1_SUB_84_U87,
    new_P1_SUB_84_U88, new_P1_SUB_84_U89, new_P1_SUB_84_U90,
    new_P1_SUB_84_U91, new_P1_SUB_84_U92, new_P1_SUB_84_U93,
    new_P1_SUB_84_U94, new_P1_SUB_84_U95, new_P1_SUB_84_U96,
    new_P1_SUB_84_U97, new_P1_SUB_84_U98, new_P1_SUB_84_U99,
    new_P1_SUB_84_U100, new_P1_SUB_84_U101, new_P1_SUB_84_U102,
    new_P1_SUB_84_U103, new_P1_SUB_84_U104, new_P1_SUB_84_U105,
    new_P1_SUB_84_U106, new_P1_SUB_84_U107, new_P1_SUB_84_U108,
    new_P1_SUB_84_U109, new_P1_SUB_84_U110, new_P1_SUB_84_U111,
    new_P1_SUB_84_U112, new_P1_SUB_84_U113, new_P1_SUB_84_U114,
    new_P1_SUB_84_U115, new_P1_SUB_84_U116, new_P1_SUB_84_U117,
    new_P1_SUB_84_U118, new_P1_SUB_84_U119, new_P1_SUB_84_U120,
    new_P1_SUB_84_U121, new_P1_SUB_84_U122, new_P1_SUB_84_U123,
    new_P1_SUB_84_U124, new_P1_SUB_84_U125, new_P1_SUB_84_U126,
    new_P1_SUB_84_U127, new_P1_SUB_84_U128, new_P1_SUB_84_U129,
    new_P1_SUB_84_U130, new_P1_SUB_84_U131, new_P1_SUB_84_U132,
    new_P1_SUB_84_U133, new_P1_SUB_84_U134, new_P1_SUB_84_U135,
    new_P1_SUB_84_U136, new_P1_SUB_84_U137, new_P1_SUB_84_U138,
    new_P1_SUB_84_U139, new_P1_SUB_84_U140, new_P1_SUB_84_U141,
    new_P1_SUB_84_U142, new_P1_SUB_84_U143, new_P1_SUB_84_U144,
    new_P1_SUB_84_U145, new_P1_SUB_84_U146, new_P1_SUB_84_U147,
    new_P1_SUB_84_U148, new_P1_SUB_84_U149, new_P1_SUB_84_U150,
    new_P1_SUB_84_U151, new_P1_SUB_84_U152, new_P1_SUB_84_U153,
    new_P1_SUB_84_U154, new_P1_SUB_84_U155, new_P1_SUB_84_U156,
    new_P1_SUB_84_U157, new_P1_SUB_84_U158, new_P1_SUB_84_U159,
    new_P1_SUB_84_U160, new_P1_SUB_84_U161, new_P1_SUB_84_U162,
    new_P1_SUB_84_U163, new_P1_SUB_84_U164, new_P1_SUB_84_U165,
    new_P1_SUB_84_U166, new_P1_SUB_84_U167, new_P1_SUB_84_U168,
    new_P1_SUB_84_U169, new_P1_SUB_84_U170, new_P1_SUB_84_U171,
    new_P1_SUB_84_U172, new_P1_SUB_84_U173, new_P1_SUB_84_U174,
    new_P1_SUB_84_U175, new_P1_SUB_84_U176, new_P1_SUB_84_U177,
    new_P1_SUB_84_U178, new_P1_SUB_84_U179, new_P1_SUB_84_U180,
    new_P1_SUB_84_U181, new_P1_SUB_84_U182, new_P1_SUB_84_U183,
    new_P1_SUB_84_U184, new_P1_SUB_84_U185, new_P1_SUB_84_U186,
    new_P1_SUB_84_U187, new_P1_SUB_84_U188, new_P1_SUB_84_U189,
    new_P1_SUB_84_U190, new_P1_SUB_84_U191, new_P1_SUB_84_U192,
    new_P1_SUB_84_U193, new_P1_SUB_84_U194, new_P1_SUB_84_U195,
    new_P1_SUB_84_U196, new_P1_SUB_84_U197, new_P1_SUB_84_U198,
    new_P1_SUB_84_U199, new_P1_SUB_84_U200, new_P1_SUB_84_U201,
    new_P1_SUB_84_U202, new_P1_SUB_84_U203, new_P1_SUB_84_U204,
    new_P1_SUB_84_U205, new_P1_SUB_84_U206, new_P1_SUB_84_U207,
    new_P1_SUB_84_U208, new_P1_SUB_84_U209, new_P1_SUB_84_U210,
    new_P1_SUB_84_U211, new_P1_SUB_84_U212, new_P1_SUB_84_U213,
    new_P1_SUB_84_U214, new_P1_SUB_84_U215, new_P1_SUB_84_U216,
    new_P1_SUB_84_U217, new_P1_SUB_84_U218, new_P1_SUB_84_U219,
    new_P1_SUB_84_U220, new_P1_SUB_84_U221, new_P1_SUB_84_U222,
    new_P1_SUB_84_U223, new_P1_SUB_84_U224, new_P1_SUB_84_U225,
    new_P1_SUB_84_U226, new_P1_SUB_84_U227, new_P1_SUB_84_U228,
    new_P1_SUB_84_U229, new_P1_SUB_84_U230, new_P1_SUB_84_U231,
    new_P1_SUB_84_U232, new_P1_SUB_84_U233, new_P1_SUB_84_U234,
    new_P1_SUB_84_U235, new_P1_SUB_84_U236, new_P1_SUB_84_U237,
    new_P1_SUB_84_U238, new_P1_SUB_84_U239, new_P1_SUB_84_U240,
    new_P1_SUB_84_U241, new_P1_SUB_84_U242, new_P1_SUB_84_U243,
    new_P1_SUB_84_U244, new_P1_SUB_84_U245, new_P1_SUB_84_U246,
    new_P1_SUB_84_U247, new_P1_SUB_84_U248, new_P1_SUB_84_U249,
    new_P1_SUB_84_U250, new_P1_SUB_84_U251, new_P1_R1309_U6,
    new_P1_R1309_U7, new_P1_R1309_U8, new_P1_R1309_U9, new_P1_R1309_U10,
    new_P1_R1282_U6, new_P1_R1282_U7, new_P1_R1282_U8, new_P1_R1282_U9,
    new_P1_R1282_U10, new_P1_R1282_U11, new_P1_R1282_U12, new_P1_R1282_U13,
    new_P1_R1282_U14, new_P1_R1282_U15, new_P1_R1282_U16, new_P1_R1282_U17,
    new_P1_R1282_U18, new_P1_R1282_U19, new_P1_R1282_U20, new_P1_R1282_U21,
    new_P1_R1282_U22, new_P1_R1282_U23, new_P1_R1282_U24, new_P1_R1282_U25,
    new_P1_R1282_U26, new_P1_R1282_U27, new_P1_R1282_U28, new_P1_R1282_U29,
    new_P1_R1282_U30, new_P1_R1282_U31, new_P1_R1282_U32, new_P1_R1282_U33,
    new_P1_R1282_U34, new_P1_R1282_U35, new_P1_R1282_U36, new_P1_R1282_U37,
    new_P1_R1282_U38, new_P1_R1282_U39, new_P1_R1282_U40, new_P1_R1282_U41,
    new_P1_R1282_U42, new_P1_R1282_U43, new_P1_R1282_U44, new_P1_R1282_U45,
    new_P1_R1282_U46, new_P1_R1282_U47, new_P1_R1282_U48, new_P1_R1282_U49,
    new_P1_R1282_U50, new_P1_R1282_U51, new_P1_R1282_U52, new_P1_R1282_U53,
    new_P1_R1282_U54, new_P1_R1282_U55, new_P1_R1282_U56, new_P1_R1282_U57,
    new_P1_R1282_U58, new_P1_R1282_U59, new_P1_R1282_U60, new_P1_R1282_U61,
    new_P1_R1282_U62, new_P1_R1282_U63, new_P1_R1282_U64, new_P1_R1282_U65,
    new_P1_R1282_U66, new_P1_R1282_U67, new_P1_R1282_U68, new_P1_R1282_U69,
    new_P1_R1282_U70, new_P1_R1282_U71, new_P1_R1282_U72, new_P1_R1282_U73,
    new_P1_R1282_U74, new_P1_R1282_U75, new_P1_R1282_U76, new_P1_R1282_U77,
    new_P1_R1282_U78, new_P1_R1282_U79, new_P1_R1282_U80, new_P1_R1282_U81,
    new_P1_R1282_U82, new_P1_R1282_U83, new_P1_R1282_U84, new_P1_R1282_U85,
    new_P1_R1282_U86, new_P1_R1282_U87, new_P1_R1282_U88, new_P1_R1282_U89,
    new_P1_R1282_U90, new_P1_R1282_U91, new_P1_R1282_U92, new_P1_R1282_U93,
    new_P1_R1282_U94, new_P1_R1282_U95, new_P1_R1282_U96, new_P1_R1282_U97,
    new_P1_R1282_U98, new_P1_R1282_U99, new_P1_R1282_U100,
    new_P1_R1282_U101, new_P1_R1282_U102, new_P1_R1282_U103,
    new_P1_R1282_U104, new_P1_R1282_U105, new_P1_R1282_U106,
    new_P1_R1282_U107, new_P1_R1282_U108, new_P1_R1282_U109,
    new_P1_R1282_U110, new_P1_R1282_U111, new_P1_R1282_U112,
    new_P1_R1282_U113, new_P1_R1282_U114, new_P1_R1282_U115,
    new_P1_R1282_U116, new_P1_R1282_U117, new_P1_R1282_U118,
    new_P1_R1282_U119, new_P1_R1282_U120, new_P1_R1282_U121,
    new_P1_R1282_U122, new_P1_R1282_U123, new_P1_R1282_U124,
    new_P1_R1282_U125, new_P1_R1282_U126, new_P1_R1282_U127,
    new_P1_R1282_U128, new_P1_R1282_U129, new_P1_R1282_U130,
    new_P1_R1282_U131, new_P1_R1282_U132, new_P1_R1282_U133,
    new_P1_R1282_U134, new_P1_R1282_U135, new_P1_R1282_U136,
    new_P1_R1282_U137, new_P1_R1282_U138, new_P1_R1282_U139,
    new_P1_R1282_U140, new_P1_R1282_U141, new_P1_R1282_U142,
    new_P1_R1282_U143, new_P1_R1282_U144, new_P1_R1282_U145,
    new_P1_R1282_U146, new_P1_R1282_U147, new_P1_R1282_U148,
    new_P1_R1282_U149, new_P1_R1282_U150, new_P1_R1282_U151,
    new_P1_R1282_U152, new_P1_R1282_U153, new_P1_R1282_U154,
    new_P1_R1282_U155, new_P1_R1282_U156, new_P1_R1282_U157,
    new_P1_R1282_U158, new_P1_R1282_U159, new_P1_R1240_U4, new_P1_R1240_U5,
    new_P1_R1240_U6, new_P1_R1240_U7, new_P1_R1240_U8, new_P1_R1240_U9,
    new_P1_R1240_U10, new_P1_R1240_U11, new_P1_R1240_U12, new_P1_R1240_U13,
    new_P1_R1240_U14, new_P1_R1240_U15, new_P1_R1240_U16, new_P1_R1240_U17,
    new_P1_R1240_U18, new_P1_R1240_U19, new_P1_R1240_U20, new_P1_R1240_U21,
    new_P1_R1240_U22, new_P1_R1240_U23, new_P1_R1240_U24, new_P1_R1240_U25,
    new_P1_R1240_U26, new_P1_R1240_U27, new_P1_R1240_U28, new_P1_R1240_U29,
    new_P1_R1240_U30, new_P1_R1240_U31, new_P1_R1240_U32, new_P1_R1240_U33,
    new_P1_R1240_U34, new_P1_R1240_U35, new_P1_R1240_U36, new_P1_R1240_U37,
    new_P1_R1240_U38, new_P1_R1240_U39, new_P1_R1240_U40, new_P1_R1240_U41,
    new_P1_R1240_U42, new_P1_R1240_U43, new_P1_R1240_U44, new_P1_R1240_U45,
    new_P1_R1240_U46, new_P1_R1240_U47, new_P1_R1240_U48, new_P1_R1240_U49,
    new_P1_R1240_U50, new_P1_R1240_U51, new_P1_R1240_U52, new_P1_R1240_U53,
    new_P1_R1240_U54, new_P1_R1240_U55, new_P1_R1240_U56, new_P1_R1240_U57,
    new_P1_R1240_U58, new_P1_R1240_U59, new_P1_R1240_U60, new_P1_R1240_U61,
    new_P1_R1240_U62, new_P1_R1240_U63, new_P1_R1240_U64, new_P1_R1240_U65,
    new_P1_R1240_U66, new_P1_R1240_U67, new_P1_R1240_U68, new_P1_R1240_U69,
    new_P1_R1240_U70, new_P1_R1240_U71, new_P1_R1240_U72, new_P1_R1240_U73,
    new_P1_R1240_U74, new_P1_R1240_U75, new_P1_R1240_U76, new_P1_R1240_U77,
    new_P1_R1240_U78, new_P1_R1240_U79, new_P1_R1240_U80, new_P1_R1240_U81,
    new_P1_R1240_U82, new_P1_R1240_U83, new_P1_R1240_U84, new_P1_R1240_U85,
    new_P1_R1240_U86, new_P1_R1240_U87, new_P1_R1240_U88, new_P1_R1240_U89,
    new_P1_R1240_U90, new_P1_R1240_U91, new_P1_R1240_U92, new_P1_R1240_U93,
    new_P1_R1240_U94, new_P1_R1240_U95, new_P1_R1240_U96, new_P1_R1240_U97,
    new_P1_R1240_U98, new_P1_R1240_U99, new_P1_R1240_U100,
    new_P1_R1240_U101, new_P1_R1240_U102, new_P1_R1240_U103,
    new_P1_R1240_U104, new_P1_R1240_U105, new_P1_R1240_U106,
    new_P1_R1240_U107, new_P1_R1240_U108, new_P1_R1240_U109,
    new_P1_R1240_U110, new_P1_R1240_U111, new_P1_R1240_U112,
    new_P1_R1240_U113, new_P1_R1240_U114, new_P1_R1240_U115,
    new_P1_R1240_U116, new_P1_R1240_U117, new_P1_R1240_U118,
    new_P1_R1240_U119, new_P1_R1240_U120, new_P1_R1240_U121,
    new_P1_R1240_U122, new_P1_R1240_U123, new_P1_R1240_U124,
    new_P1_R1240_U125, new_P1_R1240_U126, new_P1_R1240_U127,
    new_P1_R1240_U128, new_P1_R1240_U129, new_P1_R1240_U130,
    new_P1_R1240_U131, new_P1_R1240_U132, new_P1_R1240_U133,
    new_P1_R1240_U134, new_P1_R1240_U135, new_P1_R1240_U136,
    new_P1_R1240_U137, new_P1_R1240_U138, new_P1_R1240_U139,
    new_P1_R1240_U140, new_P1_R1240_U141, new_P1_R1240_U142,
    new_P1_R1240_U143, new_P1_R1240_U144, new_P1_R1240_U145,
    new_P1_R1240_U146, new_P1_R1240_U147, new_P1_R1240_U148,
    new_P1_R1240_U149, new_P1_R1240_U150, new_P1_R1240_U151,
    new_P1_R1240_U152, new_P1_R1240_U153, new_P1_R1240_U154,
    new_P1_R1240_U155, new_P1_R1240_U156, new_P1_R1240_U157,
    new_P1_R1240_U158, new_P1_R1240_U159, new_P1_R1240_U160,
    new_P1_R1240_U161, new_P1_R1240_U162, new_P1_R1240_U163,
    new_P1_R1240_U164, new_P1_R1240_U165, new_P1_R1240_U166,
    new_P1_R1240_U167, new_P1_R1240_U168, new_P1_R1240_U169,
    new_P1_R1240_U170, new_P1_R1240_U171, new_P1_R1240_U172,
    new_P1_R1240_U173, new_P1_R1240_U174, new_P1_R1240_U175,
    new_P1_R1240_U176, new_P1_R1240_U177, new_P1_R1240_U178,
    new_P1_R1240_U179, new_P1_R1240_U180, new_P1_R1240_U181,
    new_P1_R1240_U182, new_P1_R1240_U183, new_P1_R1240_U184,
    new_P1_R1240_U185, new_P1_R1240_U186, new_P1_R1240_U187,
    new_P1_R1240_U188, new_P1_R1240_U189, new_P1_R1240_U190,
    new_P1_R1240_U191, new_P1_R1240_U192, new_P1_R1240_U193,
    new_P1_R1240_U194, new_P1_R1240_U195, new_P1_R1240_U196,
    new_P1_R1240_U197, new_P1_R1240_U198, new_P1_R1240_U199,
    new_P1_R1240_U200, new_P1_R1240_U201, new_P1_R1240_U202,
    new_P1_R1240_U203, new_P1_R1240_U204, new_P1_R1240_U205,
    new_P1_R1240_U206, new_P1_R1240_U207, new_P1_R1240_U208,
    new_P1_R1240_U209, new_P1_R1240_U210, new_P1_R1240_U211,
    new_P1_R1240_U212, new_P1_R1240_U213, new_P1_R1240_U214,
    new_P1_R1240_U215, new_P1_R1240_U216, new_P1_R1240_U217,
    new_P1_R1240_U218, new_P1_R1240_U219, new_P1_R1240_U220,
    new_P1_R1240_U221, new_P1_R1240_U222, new_P1_R1240_U223,
    new_P1_R1240_U224, new_P1_R1240_U225, new_P1_R1240_U226,
    new_P1_R1240_U227, new_P1_R1240_U228, new_P1_R1240_U229,
    new_P1_R1240_U230, new_P1_R1240_U231, new_P1_R1240_U232,
    new_P1_R1240_U233, new_P1_R1240_U234, new_P1_R1240_U235,
    new_P1_R1240_U236, new_P1_R1240_U237, new_P1_R1240_U238,
    new_P1_R1240_U239, new_P1_R1240_U240, new_P1_R1240_U241,
    new_P1_R1240_U242, new_P1_R1240_U243, new_P1_R1240_U244,
    new_P1_R1240_U245, new_P1_R1240_U246, new_P1_R1240_U247,
    new_P1_R1240_U248, new_P1_R1240_U249, new_P1_R1240_U250,
    new_P1_R1240_U251, new_P1_R1240_U252, new_P1_R1240_U253,
    new_P1_R1240_U254, new_P1_R1240_U255, new_P1_R1240_U256,
    new_P1_R1240_U257, new_P1_R1240_U258, new_P1_R1240_U259,
    new_P1_R1240_U260, new_P1_R1240_U261, new_P1_R1240_U262,
    new_P1_R1240_U263, new_P1_R1240_U264, new_P1_R1240_U265,
    new_P1_R1240_U266, new_P1_R1240_U267, new_P1_R1240_U268,
    new_P1_R1240_U269, new_P1_R1240_U270, new_P1_R1240_U271,
    new_P1_R1240_U272, new_P1_R1240_U273, new_P1_R1240_U274,
    new_P1_R1240_U275, new_P1_R1240_U276, new_P1_R1240_U277,
    new_P1_R1240_U278, new_P1_R1240_U279, new_P1_R1240_U280,
    new_P1_R1240_U281, new_P1_R1240_U282, new_P1_R1240_U283,
    new_P1_R1240_U284, new_P1_R1240_U285, new_P1_R1240_U286,
    new_P1_R1240_U287, new_P1_R1240_U288, new_P1_R1240_U289,
    new_P1_R1240_U290, new_P1_R1240_U291, new_P1_R1240_U292,
    new_P1_R1240_U293, new_P1_R1240_U294, new_P1_R1240_U295,
    new_P1_R1240_U296, new_P1_R1240_U297, new_P1_R1240_U298,
    new_P1_R1240_U299, new_P1_R1240_U300, new_P1_R1240_U301,
    new_P1_R1240_U302, new_P1_R1240_U303, new_P1_R1240_U304,
    new_P1_R1240_U305, new_P1_R1240_U306, new_P1_R1240_U307,
    new_P1_R1240_U308, new_P1_R1240_U309, new_P1_R1240_U310,
    new_P1_R1240_U311, new_P1_R1240_U312, new_P1_R1240_U313,
    new_P1_R1240_U314, new_P1_R1240_U315, new_P1_R1240_U316,
    new_P1_R1240_U317, new_P1_R1240_U318, new_P1_R1240_U319,
    new_P1_R1240_U320, new_P1_R1240_U321, new_P1_R1240_U322,
    new_P1_R1240_U323, new_P1_R1240_U324, new_P1_R1240_U325,
    new_P1_R1240_U326, new_P1_R1240_U327, new_P1_R1240_U328,
    new_P1_R1240_U329, new_P1_R1240_U330, new_P1_R1240_U331,
    new_P1_R1240_U332, new_P1_R1240_U333, new_P1_R1240_U334,
    new_P1_R1240_U335, new_P1_R1240_U336, new_P1_R1240_U337,
    new_P1_R1240_U338, new_P1_R1240_U339, new_P1_R1240_U340,
    new_P1_R1240_U341, new_P1_R1240_U342, new_P1_R1240_U343,
    new_P1_R1240_U344, new_P1_R1240_U345, new_P1_R1240_U346,
    new_P1_R1240_U347, new_P1_R1240_U348, new_P1_R1240_U349,
    new_P1_R1240_U350, new_P1_R1240_U351, new_P1_R1240_U352,
    new_P1_R1240_U353, new_P1_R1240_U354, new_P1_R1240_U355,
    new_P1_R1240_U356, new_P1_R1240_U357, new_P1_R1240_U358,
    new_P1_R1240_U359, new_P1_R1240_U360, new_P1_R1240_U361,
    new_P1_R1240_U362, new_P1_R1240_U363, new_P1_R1240_U364,
    new_P1_R1240_U365, new_P1_R1240_U366, new_P1_R1240_U367,
    new_P1_R1240_U368, new_P1_R1240_U369, new_P1_R1240_U370,
    new_P1_R1240_U371, new_P1_R1240_U372, new_P1_R1240_U373,
    new_P1_R1240_U374, new_P1_R1240_U375, new_P1_R1240_U376,
    new_P1_R1240_U377, new_P1_R1240_U378, new_P1_R1240_U379,
    new_P1_R1240_U380, new_P1_R1240_U381, new_P1_R1240_U382,
    new_P1_R1240_U383, new_P1_R1240_U384, new_P1_R1240_U385,
    new_P1_R1240_U386, new_P1_R1240_U387, new_P1_R1240_U388,
    new_P1_R1240_U389, new_P1_R1240_U390, new_P1_R1240_U391,
    new_P1_R1240_U392, new_P1_R1240_U393, new_P1_R1240_U394,
    new_P1_R1240_U395, new_P1_R1240_U396, new_P1_R1240_U397,
    new_P1_R1240_U398, new_P1_R1240_U399, new_P1_R1240_U400,
    new_P1_R1240_U401, new_P1_R1240_U402, new_P1_R1240_U403,
    new_P1_R1240_U404, new_P1_R1240_U405, new_P1_R1240_U406,
    new_P1_R1240_U407, new_P1_R1240_U408, new_P1_R1240_U409,
    new_P1_R1240_U410, new_P1_R1240_U411, new_P1_R1240_U412,
    new_P1_R1240_U413, new_P1_R1240_U414, new_P1_R1240_U415,
    new_P1_R1240_U416, new_P1_R1240_U417, new_P1_R1240_U418,
    new_P1_R1240_U419, new_P1_R1240_U420, new_P1_R1240_U421,
    new_P1_R1240_U422, new_P1_R1240_U423, new_P1_R1240_U424,
    new_P1_R1240_U425, new_P1_R1240_U426, new_P1_R1240_U427,
    new_P1_R1240_U428, new_P1_R1240_U429, new_P1_R1240_U430,
    new_P1_R1240_U431, new_P1_R1240_U432, new_P1_R1240_U433,
    new_P1_R1240_U434, new_P1_R1240_U435, new_P1_R1240_U436,
    new_P1_R1240_U437, new_P1_R1240_U438, new_P1_R1240_U439,
    new_P1_R1240_U440, new_P1_R1240_U441, new_P1_R1240_U442,
    new_P1_R1240_U443, new_P1_R1240_U444, new_P1_R1240_U445,
    new_P1_R1240_U446, new_P1_R1240_U447, new_P1_R1240_U448,
    new_P1_R1240_U449, new_P1_R1240_U450, new_P1_R1240_U451,
    new_P1_R1240_U452, new_P1_R1240_U453, new_P1_R1240_U454,
    new_P1_R1240_U455, new_P1_R1240_U456, new_P1_R1240_U457,
    new_P1_R1240_U458, new_P1_R1240_U459, new_P1_R1240_U460,
    new_P1_R1240_U461, new_P1_R1240_U462, new_P1_R1240_U463,
    new_P1_R1240_U464, new_P1_R1240_U465, new_P1_R1240_U466,
    new_P1_R1240_U467, new_P1_R1240_U468, new_P1_R1240_U469,
    new_P1_R1240_U470, new_P1_R1240_U471, new_P1_R1240_U472,
    new_P1_R1240_U473, new_P1_R1240_U474, new_P1_R1240_U475,
    new_P1_R1240_U476, new_P1_R1240_U477, new_P1_R1240_U478,
    new_P1_R1240_U479, new_P1_R1240_U480, new_P1_R1240_U481,
    new_P1_R1240_U482, new_P1_R1240_U483, new_P1_R1240_U484,
    new_P1_R1240_U485, new_P1_R1240_U486, new_P1_R1240_U487,
    new_P1_R1240_U488, new_P1_R1240_U489, new_P1_R1240_U490,
    new_P1_R1240_U491, new_P1_R1240_U492, new_P1_R1240_U493,
    new_P1_R1240_U494, new_P1_R1240_U495, new_P1_R1240_U496,
    new_P1_R1240_U497, new_P1_R1240_U498, new_P1_R1240_U499,
    new_P1_R1240_U500, new_P1_R1240_U501, new_P1_R1240_U502,
    new_P1_R1240_U503, new_P1_R1162_U4, new_P1_R1162_U5, new_P1_R1162_U6,
    new_P1_R1162_U7, new_P1_R1162_U8, new_P1_R1162_U9, new_P1_R1162_U10,
    new_P1_R1162_U11, new_P1_R1162_U12, new_P1_R1162_U13, new_P1_R1162_U14,
    new_P1_R1162_U15, new_P1_R1162_U16, new_P1_R1162_U17, new_P1_R1162_U18,
    new_P1_R1162_U19, new_P1_R1162_U20, new_P1_R1162_U21, new_P1_R1162_U22,
    new_P1_R1162_U23, new_P1_R1162_U24, new_P1_R1162_U25, new_P1_R1162_U26,
    new_P1_R1162_U27, new_P1_R1162_U28, new_P1_R1162_U29, new_P1_R1162_U30,
    new_P1_R1162_U31, new_P1_R1162_U32, new_P1_R1162_U33, new_P1_R1162_U34,
    new_P1_R1162_U35, new_P1_R1162_U36, new_P1_R1162_U37, new_P1_R1162_U38,
    new_P1_R1162_U39, new_P1_R1162_U40, new_P1_R1162_U41, new_P1_R1162_U42,
    new_P1_R1162_U43, new_P1_R1162_U44, new_P1_R1162_U45, new_P1_R1162_U46,
    new_P1_R1162_U47, new_P1_R1162_U48, new_P1_R1162_U49, new_P1_R1162_U50,
    new_P1_R1162_U51, new_P1_R1162_U52, new_P1_R1162_U53, new_P1_R1162_U54,
    new_P1_R1162_U55, new_P1_R1162_U56, new_P1_R1162_U57, new_P1_R1162_U58,
    new_P1_R1162_U59, new_P1_R1162_U60, new_P1_R1162_U61, new_P1_R1162_U62,
    new_P1_R1162_U63, new_P1_R1162_U64, new_P1_R1162_U65, new_P1_R1162_U66,
    new_P1_R1162_U67, new_P1_R1162_U68, new_P1_R1162_U69, new_P1_R1162_U70,
    new_P1_R1162_U71, new_P1_R1162_U72, new_P1_R1162_U73, new_P1_R1162_U74,
    new_P1_R1162_U75, new_P1_R1162_U76, new_P1_R1162_U77, new_P1_R1162_U78,
    new_P1_R1162_U79, new_P1_R1162_U80, new_P1_R1162_U81, new_P1_R1162_U82,
    new_P1_R1162_U83, new_P1_R1162_U84, new_P1_R1162_U85, new_P1_R1162_U86,
    new_P1_R1162_U87, new_P1_R1162_U88, new_P1_R1162_U89, new_P1_R1162_U90,
    new_P1_R1162_U91, new_P1_R1162_U92, new_P1_R1162_U93, new_P1_R1162_U94,
    new_P1_R1162_U95, new_P1_R1162_U96, new_P1_R1162_U97, new_P1_R1162_U98,
    new_P1_R1162_U99, new_P1_R1162_U100, new_P1_R1162_U101,
    new_P1_R1162_U102, new_P1_R1162_U103, new_P1_R1162_U104,
    new_P1_R1162_U105, new_P1_R1162_U106, new_P1_R1162_U107,
    new_P1_R1162_U108, new_P1_R1162_U109, new_P1_R1162_U110,
    new_P1_R1162_U111, new_P1_R1162_U112, new_P1_R1162_U113,
    new_P1_R1162_U114, new_P1_R1162_U115, new_P1_R1162_U116,
    new_P1_R1162_U117, new_P1_R1162_U118, new_P1_R1162_U119,
    new_P1_R1162_U120, new_P1_R1162_U121, new_P1_R1162_U122,
    new_P1_R1162_U123, new_P1_R1162_U124, new_P1_R1162_U125,
    new_P1_R1162_U126, new_P1_R1162_U127, new_P1_R1162_U128,
    new_P1_R1162_U129, new_P1_R1162_U130, new_P1_R1162_U131,
    new_P1_R1162_U132, new_P1_R1162_U133, new_P1_R1162_U134,
    new_P1_R1162_U135, new_P1_R1162_U136, new_P1_R1162_U137,
    new_P1_R1162_U138, new_P1_R1162_U139, new_P1_R1162_U140,
    new_P1_R1162_U141, new_P1_R1162_U142, new_P1_R1162_U143,
    new_P1_R1162_U144, new_P1_R1162_U145, new_P1_R1162_U146,
    new_P1_R1162_U147, new_P1_R1162_U148, new_P1_R1162_U149,
    new_P1_R1162_U150, new_P1_R1162_U151, new_P1_R1162_U152,
    new_P1_R1162_U153, new_P1_R1162_U154, new_P1_R1162_U155,
    new_P1_R1162_U156, new_P1_R1162_U157, new_P1_R1162_U158,
    new_P1_R1162_U159, new_P1_R1162_U160, new_P1_R1162_U161,
    new_P1_R1162_U162, new_P1_R1162_U163, new_P1_R1162_U164,
    new_P1_R1162_U165, new_P1_R1162_U166, new_P1_R1162_U167,
    new_P1_R1162_U168, new_P1_R1162_U169, new_P1_R1162_U170,
    new_P1_R1162_U171, new_P1_R1162_U172, new_P1_R1162_U173,
    new_P1_R1162_U174, new_P1_R1162_U175, new_P1_R1162_U176,
    new_P1_R1162_U177, new_P1_R1162_U178, new_P1_R1162_U179,
    new_P1_R1162_U180, new_P1_R1162_U181, new_P1_R1162_U182,
    new_P1_R1162_U183, new_P1_R1162_U184, new_P1_R1162_U185,
    new_P1_R1162_U186, new_P1_R1162_U187, new_P1_R1162_U188,
    new_P1_R1162_U189, new_P1_R1162_U190, new_P1_R1162_U191,
    new_P1_R1162_U192, new_P1_R1162_U193, new_P1_R1162_U194,
    new_P1_R1162_U195, new_P1_R1162_U196, new_P1_R1162_U197,
    new_P1_R1162_U198, new_P1_R1162_U199, new_P1_R1162_U200,
    new_P1_R1162_U201, new_P1_R1162_U202, new_P1_R1162_U203,
    new_P1_R1162_U204, new_P1_R1162_U205, new_P1_R1162_U206,
    new_P1_R1162_U207, new_P1_R1162_U208, new_P1_R1162_U209,
    new_P1_R1162_U210, new_P1_R1162_U211, new_P1_R1162_U212,
    new_P1_R1162_U213, new_P1_R1162_U214, new_P1_R1162_U215,
    new_P1_R1162_U216, new_P1_R1162_U217, new_P1_R1162_U218,
    new_P1_R1162_U219, new_P1_R1162_U220, new_P1_R1162_U221,
    new_P1_R1162_U222, new_P1_R1162_U223, new_P1_R1162_U224,
    new_P1_R1162_U225, new_P1_R1162_U226, new_P1_R1162_U227,
    new_P1_R1162_U228, new_P1_R1162_U229, new_P1_R1162_U230,
    new_P1_R1162_U231, new_P1_R1162_U232, new_P1_R1162_U233,
    new_P1_R1162_U234, new_P1_R1162_U235, new_P1_R1162_U236,
    new_P1_R1162_U237, new_P1_R1162_U238, new_P1_R1162_U239,
    new_P1_R1162_U240, new_P1_R1162_U241, new_P1_R1162_U242,
    new_P1_R1162_U243, new_P1_R1162_U244, new_P1_R1162_U245,
    new_P1_R1162_U246, new_P1_R1162_U247, new_P1_R1162_U248,
    new_P1_R1162_U249, new_P1_R1162_U250, new_P1_R1162_U251,
    new_P1_R1162_U252, new_P1_R1162_U253, new_P1_R1162_U254,
    new_P1_R1162_U255, new_P1_R1162_U256, new_P1_R1162_U257,
    new_P1_R1162_U258, new_P1_R1162_U259, new_P1_R1162_U260,
    new_P1_R1162_U261, new_P1_R1162_U262, new_P1_R1162_U263,
    new_P1_R1162_U264, new_P1_R1162_U265, new_P1_R1162_U266,
    new_P1_R1162_U267, new_P1_R1162_U268, new_P1_R1162_U269,
    new_P1_R1162_U270, new_P1_R1162_U271, new_P1_R1162_U272,
    new_P1_R1162_U273, new_P1_R1162_U274, new_P1_R1162_U275,
    new_P1_R1162_U276, new_P1_R1162_U277, new_P1_R1162_U278,
    new_P1_R1162_U279, new_P1_R1162_U280, new_P1_R1162_U281,
    new_P1_R1162_U282, new_P1_R1162_U283, new_P1_R1162_U284,
    new_P1_R1162_U285, new_P1_R1162_U286, new_P1_R1162_U287,
    new_P1_R1162_U288, new_P1_R1162_U289, new_P1_R1162_U290,
    new_P1_R1162_U291, new_P1_R1162_U292, new_P1_R1162_U293,
    new_P1_R1162_U294, new_P1_R1162_U295, new_P1_R1162_U296,
    new_P1_R1162_U297, new_P1_R1162_U298, new_P1_R1162_U299,
    new_P1_R1162_U300, new_P1_R1162_U301, new_P1_R1162_U302,
    new_P1_R1162_U303, new_P1_R1162_U304, new_P1_R1162_U305,
    new_P1_R1162_U306, new_P1_R1162_U307, new_P1_R1162_U308,
    new_P1_R1117_U6, new_P1_R1117_U7, new_P1_R1117_U8, new_P1_R1117_U9,
    new_P1_R1117_U10, new_P1_R1117_U11, new_P1_R1117_U12, new_P1_R1117_U13,
    new_P1_R1117_U14, new_P1_R1117_U15, new_P1_R1117_U16, new_P1_R1117_U17,
    new_P1_R1117_U18, new_P1_R1117_U19, new_P1_R1117_U20, new_P1_R1117_U21,
    new_P1_R1117_U22, new_P1_R1117_U23, new_P1_R1117_U24, new_P1_R1117_U25,
    new_P1_R1117_U26, new_P1_R1117_U27, new_P1_R1117_U28, new_P1_R1117_U29,
    new_P1_R1117_U30, new_P1_R1117_U31, new_P1_R1117_U32, new_P1_R1117_U33,
    new_P1_R1117_U34, new_P1_R1117_U35, new_P1_R1117_U36, new_P1_R1117_U37,
    new_P1_R1117_U38, new_P1_R1117_U39, new_P1_R1117_U40, new_P1_R1117_U41,
    new_P1_R1117_U42, new_P1_R1117_U43, new_P1_R1117_U44, new_P1_R1117_U45,
    new_P1_R1117_U46, new_P1_R1117_U47, new_P1_R1117_U48, new_P1_R1117_U49,
    new_P1_R1117_U50, new_P1_R1117_U51, new_P1_R1117_U52, new_P1_R1117_U53,
    new_P1_R1117_U54, new_P1_R1117_U55, new_P1_R1117_U56, new_P1_R1117_U57,
    new_P1_R1117_U58, new_P1_R1117_U59, new_P1_R1117_U60, new_P1_R1117_U61,
    new_P1_R1117_U62, new_P1_R1117_U63, new_P1_R1117_U64, new_P1_R1117_U65,
    new_P1_R1117_U66, new_P1_R1117_U67, new_P1_R1117_U68, new_P1_R1117_U69,
    new_P1_R1117_U70, new_P1_R1117_U71, new_P1_R1117_U72, new_P1_R1117_U73,
    new_P1_R1117_U74, new_P1_R1117_U75, new_P1_R1117_U76, new_P1_R1117_U77,
    new_P1_R1117_U78, new_P1_R1117_U79, new_P1_R1117_U80, new_P1_R1117_U81,
    new_P1_R1117_U82, new_P1_R1117_U83, new_P1_R1117_U84, new_P1_R1117_U85,
    new_P1_R1117_U86, new_P1_R1117_U87, new_P1_R1117_U88, new_P1_R1117_U89,
    new_P1_R1117_U90, new_P1_R1117_U91, new_P1_R1117_U92, new_P1_R1117_U93,
    new_P1_R1117_U94, new_P1_R1117_U95, new_P1_R1117_U96, new_P1_R1117_U97,
    new_P1_R1117_U98, new_P1_R1117_U99, new_P1_R1117_U100,
    new_P1_R1117_U101, new_P1_R1117_U102, new_P1_R1117_U103,
    new_P1_R1117_U104, new_P1_R1117_U105, new_P1_R1117_U106,
    new_P1_R1117_U107, new_P1_R1117_U108, new_P1_R1117_U109,
    new_P1_R1117_U110, new_P1_R1117_U111, new_P1_R1117_U112,
    new_P1_R1117_U113, new_P1_R1117_U114, new_P1_R1117_U115,
    new_P1_R1117_U116, new_P1_R1117_U117, new_P1_R1117_U118,
    new_P1_R1117_U119, new_P1_R1117_U120, new_P1_R1117_U121,
    new_P1_R1117_U122, new_P1_R1117_U123, new_P1_R1117_U124,
    new_P1_R1117_U125, new_P1_R1117_U126, new_P1_R1117_U127,
    new_P1_R1117_U128, new_P1_R1117_U129, new_P1_R1117_U130,
    new_P1_R1117_U131, new_P1_R1117_U132, new_P1_R1117_U133,
    new_P1_R1117_U134, new_P1_R1117_U135, new_P1_R1117_U136,
    new_P1_R1117_U137, new_P1_R1117_U138, new_P1_R1117_U139,
    new_P1_R1117_U140, new_P1_R1117_U141, new_P1_R1117_U142,
    new_P1_R1117_U143, new_P1_R1117_U144, new_P1_R1117_U145,
    new_P1_R1117_U146, new_P1_R1117_U147, new_P1_R1117_U148,
    new_P1_R1117_U149, new_P1_R1117_U150, new_P1_R1117_U151,
    new_P1_R1117_U152, new_P1_R1117_U153, new_P1_R1117_U154,
    new_P1_R1117_U155, new_P1_R1117_U156, new_P1_R1117_U157,
    new_P1_R1117_U158, new_P1_R1117_U159, new_P1_R1117_U160,
    new_P1_R1117_U161, new_P1_R1117_U162, new_P1_R1117_U163,
    new_P1_R1117_U164, new_P1_R1117_U165, new_P1_R1117_U166,
    new_P1_R1117_U167, new_P1_R1117_U168, new_P1_R1117_U169,
    new_P1_R1117_U170, new_P1_R1117_U171, new_P1_R1117_U172,
    new_P1_R1117_U173, new_P1_R1117_U174, new_P1_R1117_U175,
    new_P1_R1117_U176, new_P1_R1117_U177, new_P1_R1117_U178,
    new_P1_R1117_U179, new_P1_R1117_U180, new_P1_R1117_U181,
    new_P1_R1117_U182, new_P1_R1117_U183, new_P1_R1117_U184,
    new_P1_R1117_U185, new_P1_R1117_U186, new_P1_R1117_U187,
    new_P1_R1117_U188, new_P1_R1117_U189, new_P1_R1117_U190,
    new_P1_R1117_U191, new_P1_R1117_U192, new_P1_R1117_U193,
    new_P1_R1117_U194, new_P1_R1117_U195, new_P1_R1117_U196,
    new_P1_R1117_U197, new_P1_R1117_U198, new_P1_R1117_U199,
    new_P1_R1117_U200, new_P1_R1117_U201, new_P1_R1117_U202,
    new_P1_R1117_U203, new_P1_R1117_U204, new_P1_R1117_U205,
    new_P1_R1117_U206, new_P1_R1117_U207, new_P1_R1117_U208,
    new_P1_R1117_U209, new_P1_R1117_U210, new_P1_R1117_U211,
    new_P1_R1117_U212, new_P1_R1117_U213, new_P1_R1117_U214,
    new_P1_R1117_U215, new_P1_R1117_U216, new_P1_R1117_U217,
    new_P1_R1117_U218, new_P1_R1117_U219, new_P1_R1117_U220,
    new_P1_R1117_U221, new_P1_R1117_U222, new_P1_R1117_U223,
    new_P1_R1117_U224, new_P1_R1117_U225, new_P1_R1117_U226,
    new_P1_R1117_U227, new_P1_R1117_U228, new_P1_R1117_U229,
    new_P1_R1117_U230, new_P1_R1117_U231, new_P1_R1117_U232,
    new_P1_R1117_U233, new_P1_R1117_U234, new_P1_R1117_U235,
    new_P1_R1117_U236, new_P1_R1117_U237, new_P1_R1117_U238,
    new_P1_R1117_U239, new_P1_R1117_U240, new_P1_R1117_U241,
    new_P1_R1117_U242, new_P1_R1117_U243, new_P1_R1117_U244,
    new_P1_R1117_U245, new_P1_R1117_U246, new_P1_R1117_U247,
    new_P1_R1117_U248, new_P1_R1117_U249, new_P1_R1117_U250,
    new_P1_R1117_U251, new_P1_R1117_U252, new_P1_R1117_U253,
    new_P1_R1117_U254, new_P1_R1117_U255, new_P1_R1117_U256,
    new_P1_R1117_U257, new_P1_R1117_U258, new_P1_R1117_U259,
    new_P1_R1117_U260, new_P1_R1117_U261, new_P1_R1117_U262,
    new_P1_R1117_U263, new_P1_R1117_U264, new_P1_R1117_U265,
    new_P1_R1117_U266, new_P1_R1117_U267, new_P1_R1117_U268,
    new_P1_R1117_U269, new_P1_R1117_U270, new_P1_R1117_U271,
    new_P1_R1117_U272, new_P1_R1117_U273, new_P1_R1117_U274,
    new_P1_R1117_U275, new_P1_R1117_U276, new_P1_R1117_U277,
    new_P1_R1117_U278, new_P1_R1117_U279, new_P1_R1117_U280,
    new_P1_R1117_U281, new_P1_R1117_U282, new_P1_R1117_U283,
    new_P1_R1117_U284, new_P1_R1117_U285, new_P1_R1117_U286,
    new_P1_R1117_U287, new_P1_R1117_U288, new_P1_R1117_U289,
    new_P1_R1117_U290, new_P1_R1117_U291, new_P1_R1117_U292,
    new_P1_R1117_U293, new_P1_R1117_U294, new_P1_R1117_U295,
    new_P1_R1117_U296, new_P1_R1117_U297, new_P1_R1117_U298,
    new_P1_R1117_U299, new_P1_R1117_U300, new_P1_R1117_U301,
    new_P1_R1117_U302, new_P1_R1117_U303, new_P1_R1117_U304,
    new_P1_R1117_U305, new_P1_R1117_U306, new_P1_R1117_U307,
    new_P1_R1117_U308, new_P1_R1117_U309, new_P1_R1117_U310,
    new_P1_R1117_U311, new_P1_R1117_U312, new_P1_R1117_U313,
    new_P1_R1117_U314, new_P1_R1117_U315, new_P1_R1117_U316,
    new_P1_R1117_U317, new_P1_R1117_U318, new_P1_R1117_U319,
    new_P1_R1117_U320, new_P1_R1117_U321, new_P1_R1117_U322,
    new_P1_R1117_U323, new_P1_R1117_U324, new_P1_R1117_U325,
    new_P1_R1117_U326, new_P1_R1117_U327, new_P1_R1117_U328,
    new_P1_R1117_U329, new_P1_R1117_U330, new_P1_R1117_U331,
    new_P1_R1117_U332, new_P1_R1117_U333, new_P1_R1117_U334,
    new_P1_R1117_U335, new_P1_R1117_U336, new_P1_R1117_U337,
    new_P1_R1117_U338, new_P1_R1117_U339, new_P1_R1117_U340,
    new_P1_R1117_U341, new_P1_R1117_U342, new_P1_R1117_U343,
    new_P1_R1117_U344, new_P1_R1117_U345, new_P1_R1117_U346,
    new_P1_R1117_U347, new_P1_R1117_U348, new_P1_R1117_U349,
    new_P1_R1117_U350, new_P1_R1117_U351, new_P1_R1117_U352,
    new_P1_R1117_U353, new_P1_R1117_U354, new_P1_R1117_U355,
    new_P1_R1117_U356, new_P1_R1117_U357, new_P1_R1117_U358,
    new_P1_R1117_U359, new_P1_R1117_U360, new_P1_R1117_U361,
    new_P1_R1117_U362, new_P1_R1117_U363, new_P1_R1117_U364,
    new_P1_R1117_U365, new_P1_R1117_U366, new_P1_R1117_U367,
    new_P1_R1117_U368, new_P1_R1117_U369, new_P1_R1117_U370,
    new_P1_R1117_U371, new_P1_R1117_U372, new_P1_R1117_U373,
    new_P1_R1117_U374, new_P1_R1117_U375, new_P1_R1117_U376,
    new_P1_R1117_U377, new_P1_R1117_U378, new_P1_R1117_U379,
    new_P1_R1117_U380, new_P1_R1117_U381, new_P1_R1117_U382,
    new_P1_R1117_U383, new_P1_R1117_U384, new_P1_R1117_U385,
    new_P1_R1117_U386, new_P1_R1117_U387, new_P1_R1117_U388,
    new_P1_R1117_U389, new_P1_R1117_U390, new_P1_R1117_U391,
    new_P1_R1117_U392, new_P1_R1117_U393, new_P1_R1117_U394,
    new_P1_R1117_U395, new_P1_R1117_U396, new_P1_R1117_U397,
    new_P1_R1117_U398, new_P1_R1117_U399, new_P1_R1117_U400,
    new_P1_R1117_U401, new_P1_R1117_U402, new_P1_R1117_U403,
    new_P1_R1117_U404, new_P1_R1117_U405, new_P1_R1117_U406,
    new_P1_R1117_U407, new_P1_R1117_U408, new_P1_R1117_U409,
    new_P1_R1117_U410, new_P1_R1117_U411, new_P1_R1117_U412,
    new_P1_R1117_U413, new_P1_R1117_U414, new_P1_R1117_U415,
    new_P1_R1117_U416, new_P1_R1117_U417, new_P1_R1117_U418,
    new_P1_R1117_U419, new_P1_R1117_U420, new_P1_R1117_U421,
    new_P1_R1117_U422, new_P1_R1117_U423, new_P1_R1117_U424,
    new_P1_R1117_U425, new_P1_R1117_U426, new_P1_R1117_U427,
    new_P1_R1117_U428, new_P1_R1117_U429, new_P1_R1117_U430,
    new_P1_R1117_U431, new_P1_R1117_U432, new_P1_R1117_U433,
    new_P1_R1117_U434, new_P1_R1117_U435, new_P1_R1117_U436,
    new_P1_R1117_U437, new_P1_R1117_U438, new_P1_R1117_U439,
    new_P1_R1117_U440, new_P1_R1117_U441, new_P1_R1117_U442,
    new_P1_R1117_U443, new_P1_R1117_U444, new_P1_R1117_U445,
    new_P1_R1117_U446, new_P1_R1117_U447, new_P1_R1117_U448,
    new_P1_R1117_U449, new_P1_R1117_U450, new_P1_R1117_U451,
    new_P1_R1117_U452, new_P1_R1117_U453, new_P1_R1117_U454,
    new_P1_R1117_U455, new_P1_R1117_U456, new_P1_R1117_U457,
    new_P1_R1117_U458, new_P1_R1117_U459, new_P1_R1117_U460,
    new_P1_R1117_U461, new_P1_R1117_U462, new_P1_R1117_U463,
    new_P1_R1117_U464, new_P1_R1117_U465, new_P1_R1117_U466,
    new_P1_R1117_U467, new_P1_R1117_U468, new_P1_R1117_U469,
    new_P1_R1117_U470, new_P1_R1117_U471, new_P1_R1117_U472,
    new_P1_R1117_U473, new_P1_R1375_U6, new_P1_R1375_U7, new_P1_R1375_U8,
    new_P1_R1375_U9, new_P1_R1375_U10, new_P1_R1375_U11, new_P1_R1375_U12,
    new_P1_R1375_U13, new_P1_R1375_U14, new_P1_R1375_U15, new_P1_R1375_U16,
    new_P1_R1375_U17, new_P1_R1375_U18, new_P1_R1375_U19, new_P1_R1375_U20,
    new_P1_R1375_U21, new_P1_R1375_U22, new_P1_R1375_U23, new_P1_R1375_U24,
    new_P1_R1375_U25, new_P1_R1375_U26, new_P1_R1375_U27, new_P1_R1375_U28,
    new_P1_R1375_U29, new_P1_R1375_U30, new_P1_R1375_U31, new_P1_R1375_U32,
    new_P1_R1375_U33, new_P1_R1375_U34, new_P1_R1375_U35, new_P1_R1375_U36,
    new_P1_R1375_U37, new_P1_R1375_U38, new_P1_R1375_U39, new_P1_R1375_U40,
    new_P1_R1375_U41, new_P1_R1375_U42, new_P1_R1375_U43, new_P1_R1375_U44,
    new_P1_R1375_U45, new_P1_R1375_U46, new_P1_R1375_U47, new_P1_R1375_U48,
    new_P1_R1375_U49, new_P1_R1375_U50, new_P1_R1375_U51, new_P1_R1375_U52,
    new_P1_R1375_U53, new_P1_R1375_U54, new_P1_R1375_U55, new_P1_R1375_U56,
    new_P1_R1375_U57, new_P1_R1375_U58, new_P1_R1375_U59, new_P1_R1375_U60,
    new_P1_R1375_U61, new_P1_R1375_U62, new_P1_R1375_U63, new_P1_R1375_U64,
    new_P1_R1375_U65, new_P1_R1375_U66, new_P1_R1375_U67, new_P1_R1375_U68,
    new_P1_R1375_U69, new_P1_R1375_U70, new_P1_R1375_U71, new_P1_R1375_U72,
    new_P1_R1375_U73, new_P1_R1375_U74, new_P1_R1375_U75, new_P1_R1375_U76,
    new_P1_R1375_U77, new_P1_R1375_U78, new_P1_R1375_U79, new_P1_R1375_U80,
    new_P1_R1375_U81, new_P1_R1375_U82, new_P1_R1375_U83, new_P1_R1375_U84,
    new_P1_R1375_U85, new_P1_R1375_U86, new_P1_R1375_U87, new_P1_R1375_U88,
    new_P1_R1375_U89, new_P1_R1375_U90, new_P1_R1375_U91, new_P1_R1375_U92,
    new_P1_R1375_U93, new_P1_R1375_U94, new_P1_R1375_U95, new_P1_R1375_U96,
    new_P1_R1375_U97, new_P1_R1375_U98, new_P1_R1375_U99,
    new_P1_R1375_U100, new_P1_R1375_U101, new_P1_R1375_U102,
    new_P1_R1375_U103, new_P1_R1375_U104, new_P1_R1375_U105,
    new_P1_R1375_U106, new_P1_R1375_U107, new_P1_R1375_U108,
    new_P1_R1375_U109, new_P1_R1375_U110, new_P1_R1375_U111,
    new_P1_R1375_U112, new_P1_R1375_U113, new_P1_R1375_U114,
    new_P1_R1375_U115, new_P1_R1375_U116, new_P1_R1375_U117,
    new_P1_R1375_U118, new_P1_R1375_U119, new_P1_R1375_U120,
    new_P1_R1375_U121, new_P1_R1375_U122, new_P1_R1375_U123,
    new_P1_R1375_U124, new_P1_R1375_U125, new_P1_R1375_U126,
    new_P1_R1375_U127, new_P1_R1375_U128, new_P1_R1375_U129,
    new_P1_R1375_U130, new_P1_R1375_U131, new_P1_R1375_U132,
    new_P1_R1375_U133, new_P1_R1375_U134, new_P1_R1375_U135,
    new_P1_R1375_U136, new_P1_R1375_U137, new_P1_R1375_U138,
    new_P1_R1375_U139, new_P1_R1375_U140, new_P1_R1375_U141,
    new_P1_R1375_U142, new_P1_R1375_U143, new_P1_R1375_U144,
    new_P1_R1375_U145, new_P1_R1375_U146, new_P1_R1375_U147,
    new_P1_R1375_U148, new_P1_R1375_U149, new_P1_R1375_U150,
    new_P1_R1375_U151, new_P1_R1375_U152, new_P1_R1375_U153,
    new_P1_R1375_U154, new_P1_R1375_U155, new_P1_R1375_U156,
    new_P1_R1375_U157, new_P1_R1375_U158, new_P1_R1375_U159,
    new_P1_R1375_U160, new_P1_R1375_U161, new_P1_R1375_U162,
    new_P1_R1375_U163, new_P1_R1375_U164, new_P1_R1375_U165,
    new_P1_R1375_U166, new_P1_R1375_U167, new_P1_R1375_U168,
    new_P1_R1375_U169, new_P1_R1375_U170, new_P1_R1375_U171,
    new_P1_R1375_U172, new_P1_R1375_U173, new_P1_R1375_U174,
    new_P1_R1375_U175, new_P1_R1375_U176, new_P1_R1375_U177,
    new_P1_R1375_U178, new_P1_R1375_U179, new_P1_R1375_U180,
    new_P1_R1375_U181, new_P1_R1375_U182, new_P1_R1375_U183,
    new_P1_R1375_U184, new_P1_R1375_U185, new_P1_R1375_U186,
    new_P1_R1375_U187, new_P1_R1375_U188, new_P1_R1375_U189,
    new_P1_R1375_U190, new_P1_R1375_U191, new_P1_R1375_U192,
    new_P1_R1375_U193, new_P1_R1375_U194, new_P1_R1375_U195,
    new_P1_R1375_U196, new_P1_R1375_U197, new_P1_R1375_U198,
    new_P1_R1375_U199, new_P1_R1375_U200, new_P1_R1375_U201,
    new_P1_R1375_U202, new_P1_R1375_U203, new_P1_R1375_U204,
    new_P1_R1375_U205, new_P1_R1375_U206, new_P1_R1375_U207,
    new_P1_R1352_U6, new_P1_R1352_U7, new_P1_R1207_U6, new_P1_R1207_U7,
    new_P1_R1207_U8, new_P1_R1207_U9, new_P1_R1207_U10, new_P1_R1207_U11,
    new_P1_R1207_U12, new_P1_R1207_U13, new_P1_R1207_U14, new_P1_R1207_U15,
    new_P1_R1207_U16, new_P1_R1207_U17, new_P1_R1207_U18, new_P1_R1207_U19,
    new_P1_R1207_U20, new_P1_R1207_U21, new_P1_R1207_U22, new_P1_R1207_U23,
    new_P1_R1207_U24, new_P1_R1207_U25, new_P1_R1207_U26, new_P1_R1207_U27,
    new_P1_R1207_U28, new_P1_R1207_U29, new_P1_R1207_U30, new_P1_R1207_U31,
    new_P1_R1207_U32, new_P1_R1207_U33, new_P1_R1207_U34, new_P1_R1207_U35,
    new_P1_R1207_U36, new_P1_R1207_U37, new_P1_R1207_U38, new_P1_R1207_U39,
    new_P1_R1207_U40, new_P1_R1207_U41, new_P1_R1207_U42, new_P1_R1207_U43,
    new_P1_R1207_U44, new_P1_R1207_U45, new_P1_R1207_U46, new_P1_R1207_U47,
    new_P1_R1207_U48, new_P1_R1207_U49, new_P1_R1207_U50, new_P1_R1207_U51,
    new_P1_R1207_U52, new_P1_R1207_U53, new_P1_R1207_U54, new_P1_R1207_U55,
    new_P1_R1207_U56, new_P1_R1207_U57, new_P1_R1207_U58, new_P1_R1207_U59,
    new_P1_R1207_U60, new_P1_R1207_U61, new_P1_R1207_U62, new_P1_R1207_U63,
    new_P1_R1207_U64, new_P1_R1207_U65, new_P1_R1207_U66, new_P1_R1207_U67,
    new_P1_R1207_U68, new_P1_R1207_U69, new_P1_R1207_U70, new_P1_R1207_U71,
    new_P1_R1207_U72, new_P1_R1207_U73, new_P1_R1207_U74, new_P1_R1207_U75,
    new_P1_R1207_U76, new_P1_R1207_U77, new_P1_R1207_U78, new_P1_R1207_U79,
    new_P1_R1207_U80, new_P1_R1207_U81, new_P1_R1207_U82, new_P1_R1207_U83,
    new_P1_R1207_U84, new_P1_R1207_U85, new_P1_R1207_U86, new_P1_R1207_U87,
    new_P1_R1207_U88, new_P1_R1207_U89, new_P1_R1207_U90, new_P1_R1207_U91,
    new_P1_R1207_U92, new_P1_R1207_U93, new_P1_R1207_U94, new_P1_R1207_U95,
    new_P1_R1207_U96, new_P1_R1207_U97, new_P1_R1207_U98, new_P1_R1207_U99,
    new_P1_R1207_U100, new_P1_R1207_U101, new_P1_R1207_U102,
    new_P1_R1207_U103, new_P1_R1207_U104, new_P1_R1207_U105,
    new_P1_R1207_U106, new_P1_R1207_U107, new_P1_R1207_U108,
    new_P1_R1207_U109, new_P1_R1207_U110, new_P1_R1207_U111,
    new_P1_R1207_U112, new_P1_R1207_U113, new_P1_R1207_U114,
    new_P1_R1207_U115, new_P1_R1207_U116, new_P1_R1207_U117,
    new_P1_R1207_U118, new_P1_R1207_U119, new_P1_R1207_U120,
    new_P1_R1207_U121, new_P1_R1207_U122, new_P1_R1207_U123,
    new_P1_R1207_U124, new_P1_R1207_U125, new_P1_R1207_U126,
    new_P1_R1207_U127, new_P1_R1207_U128, new_P1_R1207_U129,
    new_P1_R1207_U130, new_P1_R1207_U131, new_P1_R1207_U132,
    new_P1_R1207_U133, new_P1_R1207_U134, new_P1_R1207_U135,
    new_P1_R1207_U136, new_P1_R1207_U137, new_P1_R1207_U138,
    new_P1_R1207_U139, new_P1_R1207_U140, new_P1_R1207_U141,
    new_P1_R1207_U142, new_P1_R1207_U143, new_P1_R1207_U144,
    new_P1_R1207_U145, new_P1_R1207_U146, new_P1_R1207_U147,
    new_P1_R1207_U148, new_P1_R1207_U149, new_P1_R1207_U150,
    new_P1_R1207_U151, new_P1_R1207_U152, new_P1_R1207_U153,
    new_P1_R1207_U154, new_P1_R1207_U155, new_P1_R1207_U156,
    new_P1_R1207_U157, new_P1_R1207_U158, new_P1_R1207_U159,
    new_P1_R1207_U160, new_P1_R1207_U161, new_P1_R1207_U162,
    new_P1_R1207_U163, new_P1_R1207_U164, new_P1_R1207_U165,
    new_P1_R1207_U166, new_P1_R1207_U167, new_P1_R1207_U168,
    new_P1_R1207_U169, new_P1_R1207_U170, new_P1_R1207_U171,
    new_P1_R1207_U172, new_P1_R1207_U173, new_P1_R1207_U174,
    new_P1_R1207_U175, new_P1_R1207_U176, new_P1_R1207_U177,
    new_P1_R1207_U178, new_P1_R1207_U179, new_P1_R1207_U180,
    new_P1_R1207_U181, new_P1_R1207_U182, new_P1_R1207_U183,
    new_P1_R1207_U184, new_P1_R1207_U185, new_P1_R1207_U186,
    new_P1_R1207_U187, new_P1_R1207_U188, new_P1_R1207_U189,
    new_P1_R1207_U190, new_P1_R1207_U191, new_P1_R1207_U192,
    new_P1_R1207_U193, new_P1_R1207_U194, new_P1_R1207_U195,
    new_P1_R1207_U196, new_P1_R1207_U197, new_P1_R1207_U198,
    new_P1_R1207_U199, new_P1_R1207_U200, new_P1_R1207_U201,
    new_P1_R1207_U202, new_P1_R1207_U203, new_P1_R1207_U204,
    new_P1_R1207_U205, new_P1_R1207_U206, new_P1_R1207_U207,
    new_P1_R1207_U208, new_P1_R1207_U209, new_P1_R1207_U210,
    new_P1_R1207_U211, new_P1_R1207_U212, new_P1_R1207_U213,
    new_P1_R1207_U214, new_P1_R1207_U215, new_P1_R1207_U216,
    new_P1_R1207_U217, new_P1_R1207_U218, new_P1_R1207_U219,
    new_P1_R1207_U220, new_P1_R1207_U221, new_P1_R1207_U222,
    new_P1_R1207_U223, new_P1_R1207_U224, new_P1_R1207_U225,
    new_P1_R1207_U226, new_P1_R1207_U227, new_P1_R1207_U228,
    new_P1_R1207_U229, new_P1_R1207_U230, new_P1_R1207_U231,
    new_P1_R1207_U232, new_P1_R1207_U233, new_P1_R1207_U234,
    new_P1_R1207_U235, new_P1_R1207_U236, new_P1_R1207_U237,
    new_P1_R1207_U238, new_P1_R1207_U239, new_P1_R1207_U240,
    new_P1_R1207_U241, new_P1_R1207_U242, new_P1_R1207_U243,
    new_P1_R1207_U244, new_P1_R1207_U245, new_P1_R1207_U246,
    new_P1_R1207_U247, new_P1_R1207_U248, new_P1_R1207_U249,
    new_P1_R1207_U250, new_P1_R1207_U251, new_P1_R1207_U252,
    new_P1_R1207_U253, new_P1_R1207_U254, new_P1_R1207_U255,
    new_P1_R1207_U256, new_P1_R1207_U257, new_P1_R1207_U258,
    new_P1_R1207_U259, new_P1_R1207_U260, new_P1_R1207_U261,
    new_P1_R1207_U262, new_P1_R1207_U263, new_P1_R1207_U264,
    new_P1_R1207_U265, new_P1_R1207_U266, new_P1_R1207_U267,
    new_P1_R1207_U268, new_P1_R1207_U269, new_P1_R1207_U270,
    new_P1_R1207_U271, new_P1_R1207_U272, new_P1_R1207_U273,
    new_P1_R1207_U274, new_P1_R1207_U275, new_P1_R1207_U276,
    new_P1_R1207_U277, new_P1_R1207_U278, new_P1_R1207_U279,
    new_P1_R1207_U280, new_P1_R1207_U281, new_P1_R1207_U282,
    new_P1_R1207_U283, new_P1_R1207_U284, new_P1_R1207_U285,
    new_P1_R1207_U286, new_P1_R1207_U287, new_P1_R1207_U288,
    new_P1_R1207_U289, new_P1_R1207_U290, new_P1_R1207_U291,
    new_P1_R1207_U292, new_P1_R1207_U293, new_P1_R1207_U294,
    new_P1_R1207_U295, new_P1_R1207_U296, new_P1_R1207_U297,
    new_P1_R1207_U298, new_P1_R1207_U299, new_P1_R1207_U300,
    new_P1_R1207_U301, new_P1_R1207_U302, new_P1_R1207_U303,
    new_P1_R1207_U304, new_P1_R1207_U305, new_P1_R1207_U306,
    new_P1_R1207_U307, new_P1_R1207_U308, new_P1_R1207_U309,
    new_P1_R1207_U310, new_P1_R1207_U311, new_P1_R1207_U312,
    new_P1_R1207_U313, new_P1_R1207_U314, new_P1_R1207_U315,
    new_P1_R1207_U316, new_P1_R1207_U317, new_P1_R1207_U318,
    new_P1_R1207_U319, new_P1_R1207_U320, new_P1_R1207_U321,
    new_P1_R1207_U322, new_P1_R1207_U323, new_P1_R1207_U324,
    new_P1_R1207_U325, new_P1_R1207_U326, new_P1_R1207_U327,
    new_P1_R1207_U328, new_P1_R1207_U329, new_P1_R1207_U330,
    new_P1_R1207_U331, new_P1_R1207_U332, new_P1_R1207_U333,
    new_P1_R1207_U334, new_P1_R1207_U335, new_P1_R1207_U336,
    new_P1_R1207_U337, new_P1_R1207_U338, new_P1_R1207_U339,
    new_P1_R1207_U340, new_P1_R1207_U341, new_P1_R1207_U342,
    new_P1_R1207_U343, new_P1_R1207_U344, new_P1_R1207_U345,
    new_P1_R1207_U346, new_P1_R1207_U347, new_P1_R1207_U348,
    new_P1_R1207_U349, new_P1_R1207_U350, new_P1_R1207_U351,
    new_P1_R1207_U352, new_P1_R1207_U353, new_P1_R1207_U354,
    new_P1_R1207_U355, new_P1_R1207_U356, new_P1_R1207_U357,
    new_P1_R1207_U358, new_P1_R1207_U359, new_P1_R1207_U360,
    new_P1_R1207_U361, new_P1_R1207_U362, new_P1_R1207_U363,
    new_P1_R1207_U364, new_P1_R1207_U365, new_P1_R1207_U366,
    new_P1_R1207_U367, new_P1_R1207_U368, new_P1_R1207_U369,
    new_P1_R1207_U370, new_P1_R1207_U371, new_P1_R1207_U372,
    new_P1_R1207_U373, new_P1_R1207_U374, new_P1_R1207_U375,
    new_P1_R1207_U376, new_P1_R1207_U377, new_P1_R1207_U378,
    new_P1_R1207_U379, new_P1_R1207_U380, new_P1_R1207_U381,
    new_P1_R1207_U382, new_P1_R1207_U383, new_P1_R1207_U384,
    new_P1_R1207_U385, new_P1_R1207_U386, new_P1_R1207_U387,
    new_P1_R1207_U388, new_P1_R1207_U389, new_P1_R1207_U390,
    new_P1_R1207_U391, new_P1_R1207_U392, new_P1_R1207_U393,
    new_P1_R1207_U394, new_P1_R1207_U395, new_P1_R1207_U396,
    new_P1_R1207_U397, new_P1_R1207_U398, new_P1_R1207_U399,
    new_P1_R1207_U400, new_P1_R1207_U401, new_P1_R1207_U402,
    new_P1_R1207_U403, new_P1_R1207_U404, new_P1_R1207_U405,
    new_P1_R1207_U406, new_P1_R1207_U407, new_P1_R1207_U408,
    new_P1_R1207_U409, new_P1_R1207_U410, new_P1_R1207_U411,
    new_P1_R1207_U412, new_P1_R1207_U413, new_P1_R1207_U414,
    new_P1_R1207_U415, new_P1_R1207_U416, new_P1_R1207_U417,
    new_P1_R1207_U418, new_P1_R1207_U419, new_P1_R1207_U420,
    new_P1_R1207_U421, new_P1_R1207_U422, new_P1_R1207_U423,
    new_P1_R1207_U424, new_P1_R1207_U425, new_P1_R1207_U426,
    new_P1_R1207_U427, new_P1_R1207_U428, new_P1_R1207_U429,
    new_P1_R1207_U430, new_P1_R1207_U431, new_P1_R1207_U432,
    new_P1_R1207_U433, new_P1_R1207_U434, new_P1_R1207_U435,
    new_P1_R1207_U436, new_P1_R1207_U437, new_P1_R1207_U438,
    new_P1_R1207_U439, new_P1_R1207_U440, new_P1_R1207_U441,
    new_P1_R1207_U442, new_P1_R1207_U443, new_P1_R1207_U444,
    new_P1_R1207_U445, new_P1_R1207_U446, new_P1_R1207_U447,
    new_P1_R1207_U448, new_P1_R1207_U449, new_P1_R1207_U450,
    new_P1_R1207_U451, new_P1_R1207_U452, new_P1_R1207_U453,
    new_P1_R1207_U454, new_P1_R1207_U455, new_P1_R1207_U456,
    new_P1_R1207_U457, new_P1_R1207_U458, new_P1_R1207_U459,
    new_P1_R1207_U460, new_P1_R1207_U461, new_P1_R1207_U462,
    new_P1_R1207_U463, new_P1_R1207_U464, new_P1_R1207_U465,
    new_P1_R1207_U466, new_P1_R1207_U467, new_P1_R1207_U468,
    new_P1_R1207_U469, new_P1_R1207_U470, new_P1_R1207_U471,
    new_P1_R1207_U472, new_P1_R1207_U473, new_P1_R1165_U4, new_P1_R1165_U5,
    new_P1_R1165_U6, new_P1_R1165_U7, new_P1_R1165_U8, new_P1_R1165_U9,
    new_P1_R1165_U10, new_P1_R1165_U11, new_P1_R1165_U12, new_P1_R1165_U13,
    new_P1_R1165_U14, new_P1_R1165_U15, new_P1_R1165_U16, new_P1_R1165_U17,
    new_P1_R1165_U18, new_P1_R1165_U19, new_P1_R1165_U20, new_P1_R1165_U21,
    new_P1_R1165_U22, new_P1_R1165_U23, new_P1_R1165_U24, new_P1_R1165_U25,
    new_P1_R1165_U26, new_P1_R1165_U27, new_P1_R1165_U28, new_P1_R1165_U29,
    new_P1_R1165_U30, new_P1_R1165_U31, new_P1_R1165_U32, new_P1_R1165_U33,
    new_P1_R1165_U34, new_P1_R1165_U35, new_P1_R1165_U36, new_P1_R1165_U37,
    new_P1_R1165_U38, new_P1_R1165_U39, new_P1_R1165_U40, new_P1_R1165_U41,
    new_P1_R1165_U42, new_P1_R1165_U43, new_P1_R1165_U44, new_P1_R1165_U45,
    new_P1_R1165_U46, new_P1_R1165_U47, new_P1_R1165_U48, new_P1_R1165_U49,
    new_P1_R1165_U50, new_P1_R1165_U51, new_P1_R1165_U52, new_P1_R1165_U53,
    new_P1_R1165_U54, new_P1_R1165_U55, new_P1_R1165_U56, new_P1_R1165_U57,
    new_P1_R1165_U58, new_P1_R1165_U59, new_P1_R1165_U60, new_P1_R1165_U61,
    new_P1_R1165_U62, new_P1_R1165_U63, new_P1_R1165_U64, new_P1_R1165_U65,
    new_P1_R1165_U66, new_P1_R1165_U67, new_P1_R1165_U68, new_P1_R1165_U69,
    new_P1_R1165_U70, new_P1_R1165_U71, new_P1_R1165_U72, new_P1_R1165_U73,
    new_P1_R1165_U74, new_P1_R1165_U75, new_P1_R1165_U76, new_P1_R1165_U77,
    new_P1_R1165_U78, new_P1_R1165_U79, new_P1_R1165_U80, new_P1_R1165_U81,
    new_P1_R1165_U82, new_P1_R1165_U83, new_P1_R1165_U84, new_P1_R1165_U85,
    new_P1_R1165_U86, new_P1_R1165_U87, new_P1_R1165_U88, new_P1_R1165_U89,
    new_P1_R1165_U90, new_P1_R1165_U91, new_P1_R1165_U92, new_P1_R1165_U93,
    new_P1_R1165_U94, new_P1_R1165_U95, new_P1_R1165_U96, new_P1_R1165_U97,
    new_P1_R1165_U98, new_P1_R1165_U99, new_P1_R1165_U100,
    new_P1_R1165_U101, new_P1_R1165_U102, new_P1_R1165_U103,
    new_P1_R1165_U104, new_P1_R1165_U105, new_P1_R1165_U106,
    new_P1_R1165_U107, new_P1_R1165_U108, new_P1_R1165_U109,
    new_P1_R1165_U110, new_P1_R1165_U111, new_P1_R1165_U112,
    new_P1_R1165_U113, new_P1_R1165_U114, new_P1_R1165_U115,
    new_P1_R1165_U116, new_P1_R1165_U117, new_P1_R1165_U118,
    new_P1_R1165_U119, new_P1_R1165_U120, new_P1_R1165_U121,
    new_P1_R1165_U122, new_P1_R1165_U123, new_P1_R1165_U124,
    new_P1_R1165_U125, new_P1_R1165_U126, new_P1_R1165_U127,
    new_P1_R1165_U128, new_P1_R1165_U129, new_P1_R1165_U130,
    new_P1_R1165_U131, new_P1_R1165_U132, new_P1_R1165_U133,
    new_P1_R1165_U134, new_P1_R1165_U135, new_P1_R1165_U136,
    new_P1_R1165_U137, new_P1_R1165_U138, new_P1_R1165_U139,
    new_P1_R1165_U140, new_P1_R1165_U141, new_P1_R1165_U142,
    new_P1_R1165_U143, new_P1_R1165_U144, new_P1_R1165_U145,
    new_P1_R1165_U146, new_P1_R1165_U147, new_P1_R1165_U148,
    new_P1_R1165_U149, new_P1_R1165_U150, new_P1_R1165_U151,
    new_P1_R1165_U152, new_P1_R1165_U153, new_P1_R1165_U154,
    new_P1_R1165_U155, new_P1_R1165_U156, new_P1_R1165_U157,
    new_P1_R1165_U158, new_P1_R1165_U159, new_P1_R1165_U160,
    new_P1_R1165_U161, new_P1_R1165_U162, new_P1_R1165_U163,
    new_P1_R1165_U164, new_P1_R1165_U165, new_P1_R1165_U166,
    new_P1_R1165_U167, new_P1_R1165_U168, new_P1_R1165_U169,
    new_P1_R1165_U170, new_P1_R1165_U171, new_P1_R1165_U172,
    new_P1_R1165_U173, new_P1_R1165_U174, new_P1_R1165_U175,
    new_P1_R1165_U176, new_P1_R1165_U177, new_P1_R1165_U178,
    new_P1_R1165_U179, new_P1_R1165_U180, new_P1_R1165_U181,
    new_P1_R1165_U182, new_P1_R1165_U183, new_P1_R1165_U184,
    new_P1_R1165_U185, new_P1_R1165_U186, new_P1_R1165_U187,
    new_P1_R1165_U188, new_P1_R1165_U189, new_P1_R1165_U190,
    new_P1_R1165_U191, new_P1_R1165_U192, new_P1_R1165_U193,
    new_P1_R1165_U194, new_P1_R1165_U195, new_P1_R1165_U196,
    new_P1_R1165_U197, new_P1_R1165_U198, new_P1_R1165_U199,
    new_P1_R1165_U200, new_P1_R1165_U201, new_P1_R1165_U202,
    new_P1_R1165_U203, new_P1_R1165_U204, new_P1_R1165_U205,
    new_P1_R1165_U206, new_P1_R1165_U207, new_P1_R1165_U208,
    new_P1_R1165_U209, new_P1_R1165_U210, new_P1_R1165_U211,
    new_P1_R1165_U212, new_P1_R1165_U213, new_P1_R1165_U214,
    new_P1_R1165_U215, new_P1_R1165_U216, new_P1_R1165_U217,
    new_P1_R1165_U218, new_P1_R1165_U219, new_P1_R1165_U220,
    new_P1_R1165_U221, new_P1_R1165_U222, new_P1_R1165_U223,
    new_P1_R1165_U224, new_P1_R1165_U225, new_P1_R1165_U226,
    new_P1_R1165_U227, new_P1_R1165_U228, new_P1_R1165_U229,
    new_P1_R1165_U230, new_P1_R1165_U231, new_P1_R1165_U232,
    new_P1_R1165_U233, new_P1_R1165_U234, new_P1_R1165_U235,
    new_P1_R1165_U236, new_P1_R1165_U237, new_P1_R1165_U238,
    new_P1_R1165_U239, new_P1_R1165_U240, new_P1_R1165_U241,
    new_P1_R1165_U242, new_P1_R1165_U243, new_P1_R1165_U244,
    new_P1_R1165_U245, new_P1_R1165_U246, new_P1_R1165_U247,
    new_P1_R1165_U248, new_P1_R1165_U249, new_P1_R1165_U250,
    new_P1_R1165_U251, new_P1_R1165_U252, new_P1_R1165_U253,
    new_P1_R1165_U254, new_P1_R1165_U255, new_P1_R1165_U256,
    new_P1_R1165_U257, new_P1_R1165_U258, new_P1_R1165_U259,
    new_P1_R1165_U260, new_P1_R1165_U261, new_P1_R1165_U262,
    new_P1_R1165_U263, new_P1_R1165_U264, new_P1_R1165_U265,
    new_P1_R1165_U266, new_P1_R1165_U267, new_P1_R1165_U268,
    new_P1_R1165_U269, new_P1_R1165_U270, new_P1_R1165_U271,
    new_P1_R1165_U272, new_P1_R1165_U273, new_P1_R1165_U274,
    new_P1_R1165_U275, new_P1_R1165_U276, new_P1_R1165_U277,
    new_P1_R1165_U278, new_P1_R1165_U279, new_P1_R1165_U280,
    new_P1_R1165_U281, new_P1_R1165_U282, new_P1_R1165_U283,
    new_P1_R1165_U284, new_P1_R1165_U285, new_P1_R1165_U286,
    new_P1_R1165_U287, new_P1_R1165_U288, new_P1_R1165_U289,
    new_P1_R1165_U290, new_P1_R1165_U291, new_P1_R1165_U292,
    new_P1_R1165_U293, new_P1_R1165_U294, new_P1_R1165_U295,
    new_P1_R1165_U296, new_P1_R1165_U297, new_P1_R1165_U298,
    new_P1_R1165_U299, new_P1_R1165_U300, new_P1_R1165_U301,
    new_P1_R1165_U302, new_P1_R1165_U303, new_P1_R1165_U304,
    new_P1_R1165_U305, new_P1_R1165_U306, new_P1_R1165_U307,
    new_P1_R1165_U308, new_P1_R1165_U309, new_P1_R1165_U310,
    new_P1_R1165_U311, new_P1_R1165_U312, new_P1_R1165_U313,
    new_P1_R1165_U314, new_P1_R1165_U315, new_P1_R1165_U316,
    new_P1_R1165_U317, new_P1_R1165_U318, new_P1_R1165_U319,
    new_P1_R1165_U320, new_P1_R1165_U321, new_P1_R1165_U322,
    new_P1_R1165_U323, new_P1_R1165_U324, new_P1_R1165_U325,
    new_P1_R1165_U326, new_P1_R1165_U327, new_P1_R1165_U328,
    new_P1_R1165_U329, new_P1_R1165_U330, new_P1_R1165_U331,
    new_P1_R1165_U332, new_P1_R1165_U333, new_P1_R1165_U334,
    new_P1_R1165_U335, new_P1_R1165_U336, new_P1_R1165_U337,
    new_P1_R1165_U338, new_P1_R1165_U339, new_P1_R1165_U340,
    new_P1_R1165_U341, new_P1_R1165_U342, new_P1_R1165_U343,
    new_P1_R1165_U344, new_P1_R1165_U345, new_P1_R1165_U346,
    new_P1_R1165_U347, new_P1_R1165_U348, new_P1_R1165_U349,
    new_P1_R1165_U350, new_P1_R1165_U351, new_P1_R1165_U352,
    new_P1_R1165_U353, new_P1_R1165_U354, new_P1_R1165_U355,
    new_P1_R1165_U356, new_P1_R1165_U357, new_P1_R1165_U358,
    new_P1_R1165_U359, new_P1_R1165_U360, new_P1_R1165_U361,
    new_P1_R1165_U362, new_P1_R1165_U363, new_P1_R1165_U364,
    new_P1_R1165_U365, new_P1_R1165_U366, new_P1_R1165_U367,
    new_P1_R1165_U368, new_P1_R1165_U369, new_P1_R1165_U370,
    new_P1_R1165_U371, new_P1_R1165_U372, new_P1_R1165_U373,
    new_P1_R1165_U374, new_P1_R1165_U375, new_P1_R1165_U376,
    new_P1_R1165_U377, new_P1_R1165_U378, new_P1_R1165_U379,
    new_P1_R1165_U380, new_P1_R1165_U381, new_P1_R1165_U382,
    new_P1_R1165_U383, new_P1_R1165_U384, new_P1_R1165_U385,
    new_P1_R1165_U386, new_P1_R1165_U387, new_P1_R1165_U388,
    new_P1_R1165_U389, new_P1_R1165_U390, new_P1_R1165_U391,
    new_P1_R1165_U392, new_P1_R1165_U393, new_P1_R1165_U394,
    new_P1_R1165_U395, new_P1_R1165_U396, new_P1_R1165_U397,
    new_P1_R1165_U398, new_P1_R1165_U399, new_P1_R1165_U400,
    new_P1_R1165_U401, new_P1_R1165_U402, new_P1_R1165_U403,
    new_P1_R1165_U404, new_P1_R1165_U405, new_P1_R1165_U406,
    new_P1_R1165_U407, new_P1_R1165_U408, new_P1_R1165_U409,
    new_P1_R1165_U410, new_P1_R1165_U411, new_P1_R1165_U412,
    new_P1_R1165_U413, new_P1_R1165_U414, new_P1_R1165_U415,
    new_P1_R1165_U416, new_P1_R1165_U417, new_P1_R1165_U418,
    new_P1_R1165_U419, new_P1_R1165_U420, new_P1_R1165_U421,
    new_P1_R1165_U422, new_P1_R1165_U423, new_P1_R1165_U424,
    new_P1_R1165_U425, new_P1_R1165_U426, new_P1_R1165_U427,
    new_P1_R1165_U428, new_P1_R1165_U429, new_P1_R1165_U430,
    new_P1_R1165_U431, new_P1_R1165_U432, new_P1_R1165_U433,
    new_P1_R1165_U434, new_P1_R1165_U435, new_P1_R1165_U436,
    new_P1_R1165_U437, new_P1_R1165_U438, new_P1_R1165_U439,
    new_P1_R1165_U440, new_P1_R1165_U441, new_P1_R1165_U442,
    new_P1_R1165_U443, new_P1_R1165_U444, new_P1_R1165_U445,
    new_P1_R1165_U446, new_P1_R1165_U447, new_P1_R1165_U448,
    new_P1_R1165_U449, new_P1_R1165_U450, new_P1_R1165_U451,
    new_P1_R1165_U452, new_P1_R1165_U453, new_P1_R1165_U454,
    new_P1_R1165_U455, new_P1_R1165_U456, new_P1_R1165_U457,
    new_P1_R1165_U458, new_P1_R1165_U459, new_P1_R1165_U460,
    new_P1_R1165_U461, new_P1_R1165_U462, new_P1_R1165_U463,
    new_P1_R1165_U464, new_P1_R1165_U465, new_P1_R1165_U466,
    new_P1_R1165_U467, new_P1_R1165_U468, new_P1_R1165_U469,
    new_P1_R1165_U470, new_P1_R1165_U471, new_P1_R1165_U472,
    new_P1_R1165_U473, new_P1_R1165_U474, new_P1_R1165_U475,
    new_P1_R1165_U476, new_P1_R1165_U477, new_P1_R1165_U478,
    new_P1_R1165_U479, new_P1_R1165_U480, new_P1_R1165_U481,
    new_P1_R1165_U482, new_P1_R1165_U483, new_P1_R1165_U484,
    new_P1_R1165_U485, new_P1_R1165_U486, new_P1_R1165_U487,
    new_P1_R1165_U488, new_P1_R1165_U489, new_P1_R1165_U490,
    new_P1_R1165_U491, new_P1_R1165_U492, new_P1_R1165_U493,
    new_P1_R1165_U494, new_P1_R1165_U495, new_P1_R1165_U496,
    new_P1_R1165_U497, new_P1_R1165_U498, new_P1_R1165_U499,
    new_P1_R1165_U500, new_P1_R1165_U501, new_P1_R1165_U502,
    new_P1_R1165_U503, new_P1_R1165_U504, new_P1_R1165_U505,
    new_P1_R1165_U506, new_P1_R1165_U507, new_P1_R1165_U508,
    new_P1_R1165_U509, new_P1_R1165_U510, new_P1_R1165_U511,
    new_P1_R1165_U512, new_P1_R1165_U513, new_P1_R1165_U514,
    new_P1_R1165_U515, new_P1_R1165_U516, new_P1_R1165_U517,
    new_P1_R1165_U518, new_P1_R1165_U519, new_P1_R1165_U520,
    new_P1_R1165_U521, new_P1_R1165_U522, new_P1_R1165_U523,
    new_P1_R1165_U524, new_P1_R1165_U525, new_P1_R1165_U526,
    new_P1_R1165_U527, new_P1_R1165_U528, new_P1_R1165_U529,
    new_P1_R1165_U530, new_P1_R1165_U531, new_P1_R1165_U532,
    new_P1_R1165_U533, new_P1_R1165_U534, new_P1_R1165_U535,
    new_P1_R1165_U536, new_P1_R1165_U537, new_P1_R1165_U538,
    new_P1_R1165_U539, new_P1_R1165_U540, new_P1_R1165_U541,
    new_P1_R1165_U542, new_P1_R1165_U543, new_P1_R1165_U544,
    new_P1_R1165_U545, new_P1_R1165_U546, new_P1_R1165_U547,
    new_P1_R1165_U548, new_P1_R1165_U549, new_P1_R1165_U550,
    new_P1_R1165_U551, new_P1_R1165_U552, new_P1_R1165_U553,
    new_P1_R1165_U554, new_P1_R1165_U555, new_P1_R1165_U556,
    new_P1_R1165_U557, new_P1_R1165_U558, new_P1_R1165_U559,
    new_P1_R1165_U560, new_P1_R1165_U561, new_P1_R1165_U562,
    new_P1_R1165_U563, new_P1_R1165_U564, new_P1_R1165_U565,
    new_P1_R1165_U566, new_P1_R1165_U567, new_P1_R1165_U568,
    new_P1_R1165_U569, new_P1_R1165_U570, new_P1_R1165_U571,
    new_P1_R1165_U572, new_P1_R1165_U573, new_P1_R1165_U574,
    new_P1_R1165_U575, new_P1_R1165_U576, new_P1_R1165_U577,
    new_P1_R1165_U578, new_P1_R1165_U579, new_P1_R1165_U580,
    new_P1_R1165_U581, new_P1_R1165_U582, new_P1_R1165_U583,
    new_P1_R1165_U584, new_P1_R1165_U585, new_P1_R1165_U586,
    new_P1_R1165_U587, new_P1_R1165_U588, new_P1_R1165_U589,
    new_P1_R1165_U590, new_P1_R1165_U591, new_P1_R1165_U592,
    new_P1_R1165_U593, new_P1_R1165_U594, new_P1_R1165_U595,
    new_P1_R1165_U596, new_P1_R1165_U597, new_P1_R1165_U598,
    new_P1_R1165_U599, new_P1_R1165_U600, new_P1_R1165_U601,
    new_P1_R1165_U602, new_P1_R1150_U6, new_P1_R1150_U7, new_P1_R1150_U8,
    new_P1_R1150_U9, new_P1_R1150_U10, new_P1_R1150_U11, new_P1_R1150_U12,
    new_P1_R1150_U13, new_P1_R1150_U14, new_P1_R1150_U15, new_P1_R1150_U16,
    new_P1_R1150_U17, new_P1_R1150_U18, new_P1_R1150_U19, new_P1_R1150_U20,
    new_P1_R1150_U21, new_P1_R1150_U22, new_P1_R1150_U23, new_P1_R1150_U24,
    new_P1_R1150_U25, new_P1_R1150_U26, new_P1_R1150_U27, new_P1_R1150_U28,
    new_P1_R1150_U29, new_P1_R1150_U30, new_P1_R1150_U31, new_P1_R1150_U32,
    new_P1_R1150_U33, new_P1_R1150_U34, new_P1_R1150_U35, new_P1_R1150_U36,
    new_P1_R1150_U37, new_P1_R1150_U38, new_P1_R1150_U39, new_P1_R1150_U40,
    new_P1_R1150_U41, new_P1_R1150_U42, new_P1_R1150_U43, new_P1_R1150_U44,
    new_P1_R1150_U45, new_P1_R1150_U46, new_P1_R1150_U47, new_P1_R1150_U48,
    new_P1_R1150_U49, new_P1_R1150_U50, new_P1_R1150_U51, new_P1_R1150_U52,
    new_P1_R1150_U53, new_P1_R1150_U54, new_P1_R1150_U55, new_P1_R1150_U56,
    new_P1_R1150_U57, new_P1_R1150_U58, new_P1_R1150_U59, new_P1_R1150_U60,
    new_P1_R1150_U61, new_P1_R1150_U62, new_P1_R1150_U63, new_P1_R1150_U64,
    new_P1_R1150_U65, new_P1_R1150_U66, new_P1_R1150_U67, new_P1_R1150_U68,
    new_P1_R1150_U69, new_P1_R1150_U70, new_P1_R1150_U71, new_P1_R1150_U72,
    new_P1_R1150_U73, new_P1_R1150_U74, new_P1_R1150_U75, new_P1_R1150_U76,
    new_P1_R1150_U77, new_P1_R1150_U78, new_P1_R1150_U79, new_P1_R1150_U80,
    new_P1_R1150_U81, new_P1_R1150_U82, new_P1_R1150_U83, new_P1_R1150_U84,
    new_P1_R1150_U85, new_P1_R1150_U86, new_P1_R1150_U87, new_P1_R1150_U88,
    new_P1_R1150_U89, new_P1_R1150_U90, new_P1_R1150_U91, new_P1_R1150_U92,
    new_P1_R1150_U93, new_P1_R1150_U94, new_P1_R1150_U95, new_P1_R1150_U96,
    new_P1_R1150_U97, new_P1_R1150_U98, new_P1_R1150_U99,
    new_P1_R1150_U100, new_P1_R1150_U101, new_P1_R1150_U102,
    new_P1_R1150_U103, new_P1_R1150_U104, new_P1_R1150_U105,
    new_P1_R1150_U106, new_P1_R1150_U107, new_P1_R1150_U108,
    new_P1_R1150_U109, new_P1_R1150_U110, new_P1_R1150_U111,
    new_P1_R1150_U112, new_P1_R1150_U113, new_P1_R1150_U114,
    new_P1_R1150_U115, new_P1_R1150_U116, new_P1_R1150_U117,
    new_P1_R1150_U118, new_P1_R1150_U119, new_P1_R1150_U120,
    new_P1_R1150_U121, new_P1_R1150_U122, new_P1_R1150_U123,
    new_P1_R1150_U124, new_P1_R1150_U125, new_P1_R1150_U126,
    new_P1_R1150_U127, new_P1_R1150_U128, new_P1_R1150_U129,
    new_P1_R1150_U130, new_P1_R1150_U131, new_P1_R1150_U132,
    new_P1_R1150_U133, new_P1_R1150_U134, new_P1_R1150_U135,
    new_P1_R1150_U136, new_P1_R1150_U137, new_P1_R1150_U138,
    new_P1_R1150_U139, new_P1_R1150_U140, new_P1_R1150_U141,
    new_P1_R1150_U142, new_P1_R1150_U143, new_P1_R1150_U144,
    new_P1_R1150_U145, new_P1_R1150_U146, new_P1_R1150_U147,
    new_P1_R1150_U148, new_P1_R1150_U149, new_P1_R1150_U150,
    new_P1_R1150_U151, new_P1_R1150_U152, new_P1_R1150_U153,
    new_P1_R1150_U154, new_P1_R1150_U155, new_P1_R1150_U156,
    new_P1_R1150_U157, new_P1_R1150_U158, new_P1_R1150_U159,
    new_P1_R1150_U160, new_P1_R1150_U161, new_P1_R1150_U162,
    new_P1_R1150_U163, new_P1_R1150_U164, new_P1_R1150_U165,
    new_P1_R1150_U166, new_P1_R1150_U167, new_P1_R1150_U168,
    new_P1_R1150_U169, new_P1_R1150_U170, new_P1_R1150_U171,
    new_P1_R1150_U172, new_P1_R1150_U173, new_P1_R1150_U174,
    new_P1_R1150_U175, new_P1_R1150_U176, new_P1_R1150_U177,
    new_P1_R1150_U178, new_P1_R1150_U179, new_P1_R1150_U180,
    new_P1_R1150_U181, new_P1_R1150_U182, new_P1_R1150_U183,
    new_P1_R1150_U184, new_P1_R1150_U185, new_P1_R1150_U186,
    new_P1_R1150_U187, new_P1_R1150_U188, new_P1_R1150_U189,
    new_P1_R1150_U190, new_P1_R1150_U191, new_P1_R1150_U192,
    new_P1_R1150_U193, new_P1_R1150_U194, new_P1_R1150_U195,
    new_P1_R1150_U196, new_P1_R1150_U197, new_P1_R1150_U198,
    new_P1_R1150_U199, new_P1_R1150_U200, new_P1_R1150_U201,
    new_P1_R1150_U202, new_P1_R1150_U203, new_P1_R1150_U204,
    new_P1_R1150_U205, new_P1_R1150_U206, new_P1_R1150_U207,
    new_P1_R1150_U208, new_P1_R1150_U209, new_P1_R1150_U210,
    new_P1_R1150_U211, new_P1_R1150_U212, new_P1_R1150_U213,
    new_P1_R1150_U214, new_P1_R1150_U215, new_P1_R1150_U216,
    new_P1_R1150_U217, new_P1_R1150_U218, new_P1_R1150_U219,
    new_P1_R1150_U220, new_P1_R1150_U221, new_P1_R1150_U222,
    new_P1_R1150_U223, new_P1_R1150_U224, new_P1_R1150_U225,
    new_P1_R1150_U226, new_P1_R1150_U227, new_P1_R1150_U228,
    new_P1_R1150_U229, new_P1_R1150_U230, new_P1_R1150_U231,
    new_P1_R1150_U232, new_P1_R1150_U233, new_P1_R1150_U234,
    new_P1_R1150_U235, new_P1_R1150_U236, new_P1_R1150_U237,
    new_P1_R1150_U238, new_P1_R1150_U239, new_P1_R1150_U240,
    new_P1_R1150_U241, new_P1_R1150_U242, new_P1_R1150_U243,
    new_P1_R1150_U244, new_P1_R1150_U245, new_P1_R1150_U246,
    new_P1_R1150_U247, new_P1_R1150_U248, new_P1_R1150_U249,
    new_P1_R1150_U250, new_P1_R1150_U251, new_P1_R1150_U252,
    new_P1_R1150_U253, new_P1_R1150_U254, new_P1_R1150_U255,
    new_P1_R1150_U256, new_P1_R1150_U257, new_P1_R1150_U258,
    new_P1_R1150_U259, new_P1_R1150_U260, new_P1_R1150_U261,
    new_P1_R1150_U262, new_P1_R1150_U263, new_P1_R1150_U264,
    new_P1_R1150_U265, new_P1_R1150_U266, new_P1_R1150_U267,
    new_P1_R1150_U268, new_P1_R1150_U269, new_P1_R1150_U270,
    new_P1_R1150_U271, new_P1_R1150_U272, new_P1_R1150_U273,
    new_P1_R1150_U274, new_P1_R1150_U275, new_P1_R1150_U276,
    new_P1_R1150_U277, new_P1_R1150_U278, new_P1_R1150_U279,
    new_P1_R1150_U280, new_P1_R1150_U281, new_P1_R1150_U282,
    new_P1_R1150_U283, new_P1_R1150_U284, new_P1_R1150_U285,
    new_P1_R1150_U286, new_P1_R1150_U287, new_P1_R1150_U288,
    new_P1_R1150_U289, new_P1_R1150_U290, new_P1_R1150_U291,
    new_P1_R1150_U292, new_P1_R1150_U293, new_P1_R1150_U294,
    new_P1_R1150_U295, new_P1_R1150_U296, new_P1_R1150_U297,
    new_P1_R1150_U298, new_P1_R1150_U299, new_P1_R1150_U300,
    new_P1_R1150_U301, new_P1_R1150_U302, new_P1_R1150_U303,
    new_P1_R1150_U304, new_P1_R1150_U305, new_P1_R1150_U306,
    new_P1_R1150_U307, new_P1_R1150_U308, new_P1_R1150_U309,
    new_P1_R1150_U310, new_P1_R1150_U311, new_P1_R1150_U312,
    new_P1_R1150_U313, new_P1_R1150_U314, new_P1_R1150_U315,
    new_P1_R1150_U316, new_P1_R1150_U317, new_P1_R1150_U318,
    new_P1_R1150_U319, new_P1_R1150_U320, new_P1_R1150_U321,
    new_P1_R1150_U322, new_P1_R1150_U323, new_P1_R1150_U324,
    new_P1_R1150_U325, new_P1_R1150_U326, new_P1_R1150_U327,
    new_P1_R1150_U328, new_P1_R1150_U329, new_P1_R1150_U330,
    new_P1_R1150_U331, new_P1_R1150_U332, new_P1_R1150_U333,
    new_P1_R1150_U334, new_P1_R1150_U335, new_P1_R1150_U336,
    new_P1_R1150_U337, new_P1_R1150_U338, new_P1_R1150_U339,
    new_P1_R1150_U340, new_P1_R1150_U341, new_P1_R1150_U342,
    new_P1_R1150_U343, new_P1_R1150_U344, new_P1_R1150_U345,
    new_P1_R1150_U346, new_P1_R1150_U347, new_P1_R1150_U348,
    new_P1_R1150_U349, new_P1_R1150_U350, new_P1_R1150_U351,
    new_P1_R1150_U352, new_P1_R1150_U353, new_P1_R1150_U354,
    new_P1_R1150_U355, new_P1_R1150_U356, new_P1_R1150_U357,
    new_P1_R1150_U358, new_P1_R1150_U359, new_P1_R1150_U360,
    new_P1_R1150_U361, new_P1_R1150_U362, new_P1_R1150_U363,
    new_P1_R1150_U364, new_P1_R1150_U365, new_P1_R1150_U366,
    new_P1_R1150_U367, new_P1_R1150_U368, new_P1_R1150_U369,
    new_P1_R1150_U370, new_P1_R1150_U371, new_P1_R1150_U372,
    new_P1_R1150_U373, new_P1_R1150_U374, new_P1_R1150_U375,
    new_P1_R1150_U376, new_P1_R1150_U377, new_P1_R1150_U378,
    new_P1_R1150_U379, new_P1_R1150_U380, new_P1_R1150_U381,
    new_P1_R1150_U382, new_P1_R1150_U383, new_P1_R1150_U384,
    new_P1_R1150_U385, new_P1_R1150_U386, new_P1_R1150_U387,
    new_P1_R1150_U388, new_P1_R1150_U389, new_P1_R1150_U390,
    new_P1_R1150_U391, new_P1_R1150_U392, new_P1_R1150_U393,
    new_P1_R1150_U394, new_P1_R1150_U395, new_P1_R1150_U396,
    new_P1_R1150_U397, new_P1_R1150_U398, new_P1_R1150_U399,
    new_P1_R1150_U400, new_P1_R1150_U401, new_P1_R1150_U402,
    new_P1_R1150_U403, new_P1_R1150_U404, new_P1_R1150_U405,
    new_P1_R1150_U406, new_P1_R1150_U407, new_P1_R1150_U408,
    new_P1_R1150_U409, new_P1_R1150_U410, new_P1_R1150_U411,
    new_P1_R1150_U412, new_P1_R1150_U413, new_P1_R1150_U414,
    new_P1_R1150_U415, new_P1_R1150_U416, new_P1_R1150_U417,
    new_P1_R1150_U418, new_P1_R1150_U419, new_P1_R1150_U420,
    new_P1_R1150_U421, new_P1_R1150_U422, new_P1_R1150_U423,
    new_P1_R1150_U424, new_P1_R1150_U425, new_P1_R1150_U426,
    new_P1_R1150_U427, new_P1_R1150_U428, new_P1_R1150_U429,
    new_P1_R1150_U430, new_P1_R1150_U431, new_P1_R1150_U432,
    new_P1_R1150_U433, new_P1_R1150_U434, new_P1_R1150_U435,
    new_P1_R1150_U436, new_P1_R1150_U437, new_P1_R1150_U438,
    new_P1_R1150_U439, new_P1_R1150_U440, new_P1_R1150_U441,
    new_P1_R1150_U442, new_P1_R1150_U443, new_P1_R1150_U444,
    new_P1_R1150_U445, new_P1_R1150_U446, new_P1_R1150_U447,
    new_P1_R1150_U448, new_P1_R1150_U449, new_P1_R1150_U450,
    new_P1_R1150_U451, new_P1_R1150_U452, new_P1_R1150_U453,
    new_P1_R1150_U454, new_P1_R1150_U455, new_P1_R1150_U456,
    new_P1_R1150_U457, new_P1_R1150_U458, new_P1_R1150_U459,
    new_P1_R1150_U460, new_P1_R1150_U461, new_P1_R1150_U462,
    new_P1_R1150_U463, new_P1_R1150_U464, new_P1_R1150_U465,
    new_P1_R1150_U466, new_P1_R1150_U467, new_P1_R1150_U468,
    new_P1_R1150_U469, new_P1_R1150_U470, new_P1_R1150_U471,
    new_P1_R1150_U472, new_P1_R1150_U473, new_P1_R1192_U6, new_P1_R1192_U7,
    new_P1_R1192_U8, new_P1_R1192_U9, new_P1_R1192_U10, new_P1_R1192_U11,
    new_P1_R1192_U12, new_P1_R1192_U13, new_P1_R1192_U14, new_P1_R1192_U15,
    new_P1_R1192_U16, new_P1_R1192_U17, new_P1_R1192_U18, new_P1_R1192_U19,
    new_P1_R1192_U20, new_P1_R1192_U21, new_P1_R1192_U22, new_P1_R1192_U23,
    new_P1_R1192_U24, new_P1_R1192_U25, new_P1_R1192_U26, new_P1_R1192_U27,
    new_P1_R1192_U28, new_P1_R1192_U29, new_P1_R1192_U30, new_P1_R1192_U31,
    new_P1_R1192_U32, new_P1_R1192_U33, new_P1_R1192_U34, new_P1_R1192_U35,
    new_P1_R1192_U36, new_P1_R1192_U37, new_P1_R1192_U38, new_P1_R1192_U39,
    new_P1_R1192_U40, new_P1_R1192_U41, new_P1_R1192_U42, new_P1_R1192_U43,
    new_P1_R1192_U44, new_P1_R1192_U45, new_P1_R1192_U46, new_P1_R1192_U47,
    new_P1_R1192_U48, new_P1_R1192_U49, new_P1_R1192_U50, new_P1_R1192_U51,
    new_P1_R1192_U52, new_P1_R1192_U53, new_P1_R1192_U54, new_P1_R1192_U55,
    new_P1_R1192_U56, new_P1_R1192_U57, new_P1_R1192_U58, new_P1_R1192_U59,
    new_P1_R1192_U60, new_P1_R1192_U61, new_P1_R1192_U62, new_P1_R1192_U63,
    new_P1_R1192_U64, new_P1_R1192_U65, new_P1_R1192_U66, new_P1_R1192_U67,
    new_P1_R1192_U68, new_P1_R1192_U69, new_P1_R1192_U70, new_P1_R1192_U71,
    new_P1_R1192_U72, new_P1_R1192_U73, new_P1_R1192_U74, new_P1_R1192_U75,
    new_P1_R1192_U76, new_P1_R1192_U77, new_P1_R1192_U78, new_P1_R1192_U79,
    new_P1_R1192_U80, new_P1_R1192_U81, new_P1_R1192_U82, new_P1_R1192_U83,
    new_P1_R1192_U84, new_P1_R1192_U85, new_P1_R1192_U86, new_P1_R1192_U87,
    new_P1_R1192_U88, new_P1_R1192_U89, new_P1_R1192_U90, new_P1_R1192_U91,
    new_P1_R1192_U92, new_P1_R1192_U93, new_P1_R1192_U94, new_P1_R1192_U95,
    new_P1_R1192_U96, new_P1_R1192_U97, new_P1_R1192_U98, new_P1_R1192_U99,
    new_P1_R1192_U100, new_P1_R1192_U101, new_P1_R1192_U102,
    new_P1_R1192_U103, new_P1_R1192_U104, new_P1_R1192_U105,
    new_P1_R1192_U106, new_P1_R1192_U107, new_P1_R1192_U108,
    new_P1_R1192_U109, new_P1_R1192_U110, new_P1_R1192_U111,
    new_P1_R1192_U112, new_P1_R1192_U113, new_P1_R1192_U114,
    new_P1_R1192_U115, new_P1_R1192_U116, new_P1_R1192_U117,
    new_P1_R1192_U118, new_P1_R1192_U119, new_P1_R1192_U120,
    new_P1_R1192_U121, new_P1_R1192_U122, new_P1_R1192_U123,
    new_P1_R1192_U124, new_P1_R1192_U125, new_P1_R1192_U126,
    new_P1_R1192_U127, new_P1_R1192_U128, new_P1_R1192_U129,
    new_P1_R1192_U130, new_P1_R1192_U131, new_P1_R1192_U132,
    new_P1_R1192_U133, new_P1_R1192_U134, new_P1_R1192_U135,
    new_P1_R1192_U136, new_P1_R1192_U137, new_P1_R1192_U138,
    new_P1_R1192_U139, new_P1_R1192_U140, new_P1_R1192_U141,
    new_P1_R1192_U142, new_P1_R1192_U143, new_P1_R1192_U144,
    new_P1_R1192_U145, new_P1_R1192_U146, new_P1_R1192_U147,
    new_P1_R1192_U148, new_P1_R1192_U149, new_P1_R1192_U150,
    new_P1_R1192_U151, new_P1_R1192_U152, new_P1_R1192_U153,
    new_P1_R1192_U154, new_P1_R1192_U155, new_P1_R1192_U156,
    new_P1_R1192_U157, new_P1_R1192_U158, new_P1_R1192_U159,
    new_P1_R1192_U160, new_P1_R1192_U161, new_P1_R1192_U162,
    new_P1_R1192_U163, new_P1_R1192_U164, new_P1_R1192_U165,
    new_P1_R1192_U166, new_P1_R1192_U167, new_P1_R1192_U168,
    new_P1_R1192_U169, new_P1_R1192_U170, new_P1_R1192_U171,
    new_P1_R1192_U172, new_P1_R1192_U173, new_P1_R1192_U174,
    new_P1_R1192_U175, new_P1_R1192_U176, new_P1_R1192_U177,
    new_P1_R1192_U178, new_P1_R1192_U179, new_P1_R1192_U180,
    new_P1_R1192_U181, new_P1_R1192_U182, new_P1_R1192_U183,
    new_P1_R1192_U184, new_P1_R1192_U185, new_P1_R1192_U186,
    new_P1_R1192_U187, new_P1_R1192_U188, new_P1_R1192_U189,
    new_P1_R1192_U190, new_P1_R1192_U191, new_P1_R1192_U192,
    new_P1_R1192_U193, new_P1_R1192_U194, new_P1_R1192_U195,
    new_P1_R1192_U196, new_P1_R1192_U197, new_P1_R1192_U198,
    new_P1_R1192_U199, new_P1_R1192_U200, new_P1_R1192_U201,
    new_P1_R1192_U202, new_P1_R1192_U203, new_P1_R1192_U204,
    new_P1_R1192_U205, new_P1_R1192_U206, new_P1_R1192_U207,
    new_P1_R1192_U208, new_P1_R1192_U209, new_P1_R1192_U210,
    new_P1_R1192_U211, new_P1_R1192_U212, new_P1_R1192_U213,
    new_P1_R1192_U214, new_P1_R1192_U215, new_P1_R1192_U216,
    new_P1_R1192_U217, new_P1_R1192_U218, new_P1_R1192_U219,
    new_P1_R1192_U220, new_P1_R1192_U221, new_P1_R1192_U222,
    new_P1_R1192_U223, new_P1_R1192_U224, new_P1_R1192_U225,
    new_P1_R1192_U226, new_P1_R1192_U227, new_P1_R1192_U228,
    new_P1_R1192_U229, new_P1_R1192_U230, new_P1_R1192_U231,
    new_P1_R1192_U232, new_P1_R1192_U233, new_P1_R1192_U234,
    new_P1_R1192_U235, new_P1_R1192_U236, new_P1_R1192_U237,
    new_P1_R1192_U238, new_P1_R1192_U239, new_P1_R1192_U240,
    new_P1_R1192_U241, new_P1_R1192_U242, new_P1_R1192_U243,
    new_P1_R1192_U244, new_P1_R1192_U245, new_P1_R1192_U246,
    new_P1_R1192_U247, new_P1_R1192_U248, new_P1_R1192_U249,
    new_P1_R1192_U250, new_P1_R1192_U251, new_P1_R1192_U252,
    new_P1_R1192_U253, new_P1_R1192_U254, new_P1_R1192_U255,
    new_P1_R1192_U256, new_P1_R1192_U257, new_P1_R1192_U258,
    new_P1_R1192_U259, new_P1_R1192_U260, new_P1_R1192_U261,
    new_P1_R1192_U262, new_P1_R1192_U263, new_P1_R1192_U264,
    new_P1_R1192_U265, new_P1_R1192_U266, new_P1_R1192_U267,
    new_P1_R1192_U268, new_P1_R1192_U269, new_P1_R1192_U270,
    new_P1_R1192_U271, new_P1_R1192_U272, new_P1_R1192_U273,
    new_P1_R1192_U274, new_P1_R1192_U275, new_P1_R1192_U276,
    new_P1_R1192_U277, new_P1_R1192_U278, new_P1_R1192_U279,
    new_P1_R1192_U280, new_P1_R1192_U281, new_P1_R1192_U282,
    new_P1_R1192_U283, new_P1_R1192_U284, new_P1_R1192_U285,
    new_P1_R1192_U286, new_P1_R1192_U287, new_P1_R1192_U288,
    new_P1_R1192_U289, new_P1_R1192_U290, new_P1_R1192_U291,
    new_P1_R1192_U292, new_P1_R1192_U293, new_P1_R1192_U294,
    new_P1_R1192_U295, new_P1_R1192_U296, new_P1_R1192_U297,
    new_P1_R1192_U298, new_P1_R1192_U299, new_P1_R1192_U300,
    new_P1_R1192_U301, new_P1_R1192_U302, new_P1_R1192_U303,
    new_P1_R1192_U304, new_P1_R1192_U305, new_P1_R1192_U306,
    new_P1_R1192_U307, new_P1_R1192_U308, new_P1_R1192_U309,
    new_P1_R1192_U310, new_P1_R1192_U311, new_P1_R1192_U312,
    new_P1_R1192_U313, new_P1_R1192_U314, new_P1_R1192_U315,
    new_P1_R1192_U316, new_P1_R1192_U317, new_P1_R1192_U318,
    new_P1_R1192_U319, new_P1_R1192_U320, new_P1_R1192_U321,
    new_P1_R1192_U322, new_P1_R1192_U323, new_P1_R1192_U324,
    new_P1_R1192_U325, new_P1_R1192_U326, new_P1_R1192_U327,
    new_P1_R1192_U328, new_P1_R1192_U329, new_P1_R1192_U330,
    new_P1_R1192_U331, new_P1_R1192_U332, new_P1_R1192_U333,
    new_P1_R1192_U334, new_P1_R1192_U335, new_P1_R1192_U336,
    new_P1_R1192_U337, new_P1_R1192_U338, new_P1_R1192_U339,
    new_P1_R1192_U340, new_P1_R1192_U341, new_P1_R1192_U342,
    new_P1_R1192_U343, new_P1_R1192_U344, new_P1_R1192_U345,
    new_P1_R1192_U346, new_P1_R1192_U347, new_P1_R1192_U348,
    new_P1_R1192_U349, new_P1_R1192_U350, new_P1_R1192_U351,
    new_P1_R1192_U352, new_P1_R1192_U353, new_P1_R1192_U354,
    new_P1_R1192_U355, new_P1_R1192_U356, new_P1_R1192_U357,
    new_P1_R1192_U358, new_P1_R1192_U359, new_P1_R1192_U360,
    new_P1_R1192_U361, new_P1_R1192_U362, new_P1_R1192_U363,
    new_P1_R1192_U364, new_P1_R1192_U365, new_P1_R1192_U366,
    new_P1_R1192_U367, new_P1_R1192_U368, new_P1_R1192_U369,
    new_P1_R1192_U370, new_P1_R1192_U371, new_P1_R1192_U372,
    new_P1_R1192_U373, new_P1_R1192_U374, new_P1_R1192_U375,
    new_P1_R1192_U376, new_P1_R1192_U377, new_P1_R1192_U378,
    new_P1_R1192_U379, new_P1_R1192_U380, new_P1_R1192_U381,
    new_P1_R1192_U382, new_P1_R1192_U383, new_P1_R1192_U384,
    new_P1_R1192_U385, new_P1_R1192_U386, new_P1_R1192_U387,
    new_P1_R1192_U388, new_P1_R1192_U389, new_P1_R1192_U390,
    new_P1_R1192_U391, new_P1_R1192_U392, new_P1_R1192_U393,
    new_P1_R1192_U394, new_P1_R1192_U395, new_P1_R1192_U396,
    new_P1_R1192_U397, new_P1_R1192_U398, new_P1_R1192_U399,
    new_P1_R1192_U400, new_P1_R1192_U401, new_P1_R1192_U402,
    new_P1_R1192_U403, new_P1_R1192_U404, new_P1_R1192_U405,
    new_P1_R1192_U406, new_P1_R1192_U407, new_P1_R1192_U408,
    new_P1_R1192_U409, new_P1_R1192_U410, new_P1_R1192_U411,
    new_P1_R1192_U412, new_P1_R1192_U413, new_P1_R1192_U414,
    new_P1_R1192_U415, new_P1_R1192_U416, new_P1_R1192_U417,
    new_P1_R1192_U418, new_P1_R1192_U419, new_P1_R1192_U420,
    new_P1_R1192_U421, new_P1_R1192_U422, new_P1_R1192_U423,
    new_P1_R1192_U424, new_P1_R1192_U425, new_P1_R1192_U426,
    new_P1_R1192_U427, new_P1_R1192_U428, new_P1_R1192_U429,
    new_P1_R1192_U430, new_P1_R1192_U431, new_P1_R1192_U432,
    new_P1_R1192_U433, new_P1_R1192_U434, new_P1_R1192_U435,
    new_P1_R1192_U436, new_P1_R1192_U437, new_P1_R1192_U438,
    new_P1_R1192_U439, new_P1_R1192_U440, new_P1_R1192_U441,
    new_P1_R1192_U442, new_P1_R1192_U443, new_P1_R1192_U444,
    new_P1_R1192_U445, new_P1_R1192_U446, new_P1_R1192_U447,
    new_P1_R1192_U448, new_P1_R1192_U449, new_P1_R1192_U450,
    new_P1_R1192_U451, new_P1_R1192_U452, new_P1_R1192_U453,
    new_P1_R1192_U454, new_P1_R1192_U455, new_P1_R1192_U456,
    new_P1_R1192_U457, new_P1_R1192_U458, new_P1_R1192_U459,
    new_P1_R1192_U460, new_P1_R1192_U461, new_P1_R1192_U462,
    new_P1_R1192_U463, new_P1_R1192_U464, new_P1_R1192_U465,
    new_P1_R1192_U466, new_P1_R1192_U467, new_P1_R1192_U468,
    new_P1_R1192_U469, new_P1_R1192_U470, new_P1_R1192_U471,
    new_P1_R1192_U472, new_P1_R1192_U473, new_P1_LT_197_U6,
    new_P1_LT_197_U7, new_P1_LT_197_U8, new_P1_LT_197_U9,
    new_P1_LT_197_U10, new_P1_LT_197_U11, new_P1_LT_197_U12,
    new_P1_LT_197_U13, new_P1_LT_197_U14, new_P1_LT_197_U15,
    new_P1_LT_197_U16, new_P1_LT_197_U17, new_P1_LT_197_U18,
    new_P1_LT_197_U19, new_P1_LT_197_U20, new_P1_LT_197_U21,
    new_P1_LT_197_U22, new_P1_LT_197_U23, new_P1_LT_197_U24,
    new_P1_LT_197_U25, new_P1_LT_197_U26, new_P1_LT_197_U27,
    new_P1_LT_197_U28, new_P1_LT_197_U29, new_P1_LT_197_U30,
    new_P1_LT_197_U31, new_P1_LT_197_U32, new_P1_LT_197_U33,
    new_P1_LT_197_U34, new_P1_LT_197_U35, new_P1_LT_197_U36,
    new_P1_LT_197_U37, new_P1_LT_197_U38, new_P1_LT_197_U39,
    new_P1_LT_197_U40, new_P1_LT_197_U41, new_P1_LT_197_U42,
    new_P1_LT_197_U43, new_P1_LT_197_U44, new_P1_LT_197_U45,
    new_P1_LT_197_U46, new_P1_LT_197_U47, new_P1_LT_197_U48,
    new_P1_LT_197_U49, new_P1_LT_197_U50, new_P1_LT_197_U51,
    new_P1_LT_197_U52, new_P1_LT_197_U53, new_P1_LT_197_U54,
    new_P1_LT_197_U55, new_P1_LT_197_U56, new_P1_LT_197_U57,
    new_P1_LT_197_U58, new_P1_LT_197_U59, new_P1_LT_197_U60,
    new_P1_LT_197_U61, new_P1_LT_197_U62, new_P1_LT_197_U63,
    new_P1_LT_197_U64, new_P1_LT_197_U65, new_P1_LT_197_U66,
    new_P1_LT_197_U67, new_P1_LT_197_U68, new_P1_LT_197_U69,
    new_P1_LT_197_U70, new_P1_LT_197_U71, new_P1_LT_197_U72,
    new_P1_LT_197_U73, new_P1_LT_197_U74, new_P1_LT_197_U75,
    new_P1_LT_197_U76, new_P1_LT_197_U77, new_P1_LT_197_U78,
    new_P1_LT_197_U79, new_P1_LT_197_U80, new_P1_LT_197_U81,
    new_P1_LT_197_U82, new_P1_LT_197_U83, new_P1_LT_197_U84,
    new_P1_LT_197_U85, new_P1_LT_197_U86, new_P1_LT_197_U87,
    new_P1_LT_197_U88, new_P1_LT_197_U89, new_P1_LT_197_U90,
    new_P1_LT_197_U91, new_P1_LT_197_U92, new_P1_LT_197_U93,
    new_P1_LT_197_U94, new_P1_LT_197_U95, new_P1_LT_197_U96,
    new_P1_LT_197_U97, new_P1_LT_197_U98, new_P1_LT_197_U99,
    new_P1_LT_197_U100, new_P1_LT_197_U101, new_P1_LT_197_U102,
    new_P1_LT_197_U103, new_P1_LT_197_U104, new_P1_LT_197_U105,
    new_P1_LT_197_U106, new_P1_LT_197_U107, new_P1_LT_197_U108,
    new_P1_LT_197_U109, new_P1_LT_197_U110, new_P1_LT_197_U111,
    new_P1_LT_197_U112, new_P1_LT_197_U113, new_P1_LT_197_U114,
    new_P1_LT_197_U115, new_P1_LT_197_U116, new_P1_LT_197_U117,
    new_P1_LT_197_U118, new_P1_LT_197_U119, new_P1_LT_197_U120,
    new_P1_LT_197_U121, new_P1_LT_197_U122, new_P1_LT_197_U123,
    new_P1_LT_197_U124, new_P1_LT_197_U125, new_P1_LT_197_U126,
    new_P1_LT_197_U127, new_P1_LT_197_U128, new_P1_LT_197_U129,
    new_P1_LT_197_U130, new_P1_LT_197_U131, new_P1_LT_197_U132,
    new_P1_LT_197_U133, new_P1_LT_197_U134, new_P1_LT_197_U135,
    new_P1_LT_197_U136, new_P1_LT_197_U137, new_P1_LT_197_U138,
    new_P1_LT_197_U139, new_P1_LT_197_U140, new_P1_LT_197_U141,
    new_P1_LT_197_U142, new_P1_LT_197_U143, new_P1_LT_197_U144,
    new_P1_LT_197_U145, new_P1_LT_197_U146, new_P1_LT_197_U147,
    new_P1_LT_197_U148, new_P1_LT_197_U149, new_P1_LT_197_U150,
    new_P1_LT_197_U151, new_P1_LT_197_U152, new_P1_LT_197_U153,
    new_P1_LT_197_U154, new_P1_LT_197_U155, new_P1_LT_197_U156,
    new_P1_LT_197_U157, new_P1_LT_197_U158, new_P1_LT_197_U159,
    new_P1_LT_197_U160, new_P1_LT_197_U161, new_P1_LT_197_U162,
    new_P1_LT_197_U163, new_P1_LT_197_U164, new_P1_LT_197_U165,
    new_P1_LT_197_U166, new_P1_LT_197_U167, new_P1_LT_197_U168,
    new_P1_LT_197_U169, new_P1_LT_197_U170, new_P1_LT_197_U171,
    new_P1_LT_197_U172, new_P1_LT_197_U173, new_P1_LT_197_U174,
    new_P1_LT_197_U175, new_P1_LT_197_U176, new_P1_LT_197_U177,
    new_P1_LT_197_U178, new_P1_LT_197_U179, new_P1_LT_197_U180,
    new_P1_LT_197_U181, new_P1_LT_197_U182, new_P1_LT_197_U183,
    new_P1_LT_197_U184, new_P1_LT_197_U185, new_P1_LT_197_U186,
    new_P1_LT_197_U187, new_P1_LT_197_U188, new_P1_LT_197_U189,
    new_P1_LT_197_U190, new_P1_LT_197_U191, new_P1_LT_197_U192,
    new_P1_LT_197_U193, new_P1_LT_197_U194, new_P1_LT_197_U195,
    new_P1_LT_197_U196, new_P1_LT_197_U197, new_P1_LT_197_U198,
    new_P1_LT_197_U199, new_P1_LT_197_U200, new_P1_R1360_U6,
    new_P1_R1360_U7, new_P1_R1360_U8, new_P1_R1360_U9, new_P1_R1360_U10,
    new_P1_R1360_U11, new_P1_R1360_U12, new_P1_R1360_U13, new_P1_R1360_U14,
    new_P1_R1360_U15, new_P1_R1360_U16, new_P1_R1360_U17, new_P1_R1360_U18,
    new_P1_R1360_U19, new_P1_R1360_U20, new_P1_R1360_U21, new_P1_R1360_U22,
    new_P1_R1360_U23, new_P1_R1360_U24, new_P1_R1360_U25, new_P1_R1360_U26,
    new_P1_R1360_U27, new_P1_R1360_U28, new_P1_R1360_U29, new_P1_R1360_U30,
    new_P1_R1360_U31, new_P1_R1360_U32, new_P1_R1360_U33, new_P1_R1360_U34,
    new_P1_R1360_U35, new_P1_R1360_U36, new_P1_R1360_U37, new_P1_R1360_U38,
    new_P1_R1360_U39, new_P1_R1360_U40, new_P1_R1360_U41, new_P1_R1360_U42,
    new_P1_R1360_U43, new_P1_R1360_U44, new_P1_R1360_U45, new_P1_R1360_U46,
    new_P1_R1360_U47, new_P1_R1360_U48, new_P1_R1360_U49, new_P1_R1360_U50,
    new_P1_R1360_U51, new_P1_R1360_U52, new_P1_R1360_U53, new_P1_R1360_U54,
    new_P1_R1360_U55, new_P1_R1360_U56, new_P1_R1360_U57, new_P1_R1360_U58,
    new_P1_R1360_U59, new_P1_R1360_U60, new_P1_R1360_U61, new_P1_R1360_U62,
    new_P1_R1360_U63, new_P1_R1360_U64, new_P1_R1360_U65, new_P1_R1360_U66,
    new_P1_R1360_U67, new_P1_R1360_U68, new_P1_R1360_U69, new_P1_R1360_U70,
    new_P1_R1360_U71, new_P1_R1360_U72, new_P1_R1360_U73, new_P1_R1360_U74,
    new_P1_R1360_U75, new_P1_R1360_U76, new_P1_R1360_U77, new_P1_R1360_U78,
    new_P1_R1360_U79, new_P1_R1360_U80, new_P1_R1360_U81, new_P1_R1360_U82,
    new_P1_R1360_U83, new_P1_R1360_U84, new_P1_R1360_U85, new_P1_R1360_U86,
    new_P1_R1360_U87, new_P1_R1360_U88, new_P1_R1360_U89, new_P1_R1360_U90,
    new_P1_R1360_U91, new_P1_R1360_U92, new_P1_R1360_U93, new_P1_R1360_U94,
    new_P1_R1360_U95, new_P1_R1360_U96, new_P1_R1360_U97, new_P1_R1360_U98,
    new_P1_R1360_U99, new_P1_R1360_U100, new_P1_R1360_U101,
    new_P1_R1360_U102, new_P1_R1360_U103, new_P1_R1360_U104,
    new_P1_R1360_U105, new_P1_R1360_U106, new_P1_R1360_U107,
    new_P1_R1360_U108, new_P1_R1360_U109, new_P1_R1360_U110,
    new_P1_R1360_U111, new_P1_R1360_U112, new_P1_R1360_U113,
    new_P1_R1360_U114, new_P1_R1360_U115, new_P1_R1360_U116,
    new_P1_R1360_U117, new_P1_R1360_U118, new_P1_R1360_U119,
    new_P1_R1360_U120, new_P1_R1360_U121, new_P1_R1360_U122,
    new_P1_R1360_U123, new_P1_R1360_U124, new_P1_R1360_U125,
    new_P1_R1360_U126, new_P1_R1360_U127, new_P1_R1360_U128,
    new_P1_R1360_U129, new_P1_R1360_U130, new_P1_R1360_U131,
    new_P1_R1360_U132, new_P1_R1360_U133, new_P1_R1360_U134,
    new_P1_R1360_U135, new_P1_R1360_U136, new_P1_R1360_U137,
    new_P1_R1360_U138, new_P1_R1360_U139, new_P1_R1360_U140,
    new_P1_R1360_U141, new_P1_R1360_U142, new_P1_R1360_U143,
    new_P1_R1360_U144, new_P1_R1360_U145, new_P1_R1360_U146,
    new_P1_R1360_U147, new_P1_R1360_U148, new_P1_R1360_U149,
    new_P1_R1360_U150, new_P1_R1360_U151, new_P1_R1360_U152,
    new_P1_R1360_U153, new_P1_R1360_U154, new_P1_R1360_U155,
    new_P1_R1360_U156, new_P1_R1360_U157, new_P1_R1360_U158,
    new_P1_R1360_U159, new_P1_R1360_U160, new_P1_R1360_U161,
    new_P1_R1360_U162, new_P1_R1360_U163, new_P1_R1360_U164,
    new_P1_R1360_U165, new_P1_R1360_U166, new_P1_R1360_U167,
    new_P1_R1360_U168, new_P1_R1360_U169, new_P1_R1360_U170,
    new_P1_R1360_U171, new_P1_R1360_U172, new_P1_R1360_U173,
    new_P1_R1360_U174, new_P1_R1360_U175, new_P1_R1360_U176,
    new_P1_R1360_U177, new_P1_R1360_U178, new_P1_R1360_U179,
    new_P1_R1360_U180, new_P1_R1360_U181, new_P1_R1360_U182,
    new_P1_R1360_U183, new_P1_R1360_U184, new_P1_R1360_U185,
    new_P1_R1360_U186, new_P1_R1360_U187, new_P1_R1360_U188,
    new_P1_R1360_U189, new_P1_R1360_U190, new_P1_R1360_U191,
    new_P1_R1360_U192, new_P1_R1360_U193, new_P1_R1360_U194,
    new_P1_R1360_U195, new_P1_R1360_U196, new_P1_R1360_U197,
    new_P1_R1360_U198, new_P1_R1360_U199, new_P1_R1360_U200,
    new_P1_R1360_U201, new_P1_R1360_U202, new_P1_R1360_U203,
    new_P1_R1360_U204, new_P1_R1360_U205, new_P1_R1171_U4, new_P1_R1171_U5,
    new_P1_R1171_U6, new_P1_R1171_U7, new_P1_R1171_U8, new_P1_R1171_U9,
    new_P1_R1171_U10, new_P1_R1171_U11, new_P1_R1171_U12, new_P1_R1171_U13,
    new_P1_R1171_U14, new_P1_R1171_U15, new_P1_R1171_U16, new_P1_R1171_U17,
    new_P1_R1171_U18, new_P1_R1171_U19, new_P1_R1171_U20, new_P1_R1171_U21,
    new_P1_R1171_U22, new_P1_R1171_U23, new_P1_R1171_U24, new_P1_R1171_U25,
    new_P1_R1171_U26, new_P1_R1171_U27, new_P1_R1171_U28, new_P1_R1171_U29,
    new_P1_R1171_U30, new_P1_R1171_U31, new_P1_R1171_U32, new_P1_R1171_U33,
    new_P1_R1171_U34, new_P1_R1171_U35, new_P1_R1171_U36, new_P1_R1171_U37,
    new_P1_R1171_U38, new_P1_R1171_U39, new_P1_R1171_U40, new_P1_R1171_U41,
    new_P1_R1171_U42, new_P1_R1171_U43, new_P1_R1171_U44, new_P1_R1171_U45,
    new_P1_R1171_U46, new_P1_R1171_U47, new_P1_R1171_U48, new_P1_R1171_U49,
    new_P1_R1171_U50, new_P1_R1171_U51, new_P1_R1171_U52, new_P1_R1171_U53,
    new_P1_R1171_U54, new_P1_R1171_U55, new_P1_R1171_U56, new_P1_R1171_U57,
    new_P1_R1171_U58, new_P1_R1171_U59, new_P1_R1171_U60, new_P1_R1171_U61,
    new_P1_R1171_U62, new_P1_R1171_U63, new_P1_R1171_U64, new_P1_R1171_U65,
    new_P1_R1171_U66, new_P1_R1171_U67, new_P1_R1171_U68, new_P1_R1171_U69,
    new_P1_R1171_U70, new_P1_R1171_U71, new_P1_R1171_U72, new_P1_R1171_U73,
    new_P1_R1171_U74, new_P1_R1171_U75, new_P1_R1171_U76, new_P1_R1171_U77,
    new_P1_R1171_U78, new_P1_R1171_U79, new_P1_R1171_U80, new_P1_R1171_U81,
    new_P1_R1171_U82, new_P1_R1171_U83, new_P1_R1171_U84, new_P1_R1171_U85,
    new_P1_R1171_U86, new_P1_R1171_U87, new_P1_R1171_U88, new_P1_R1171_U89,
    new_P1_R1171_U90, new_P1_R1171_U91, new_P1_R1171_U92, new_P1_R1171_U93,
    new_P1_R1171_U94, new_P1_R1171_U95, new_P1_R1171_U96, new_P1_R1171_U97,
    new_P1_R1171_U98, new_P1_R1171_U99, new_P1_R1171_U100,
    new_P1_R1171_U101, new_P1_R1171_U102, new_P1_R1171_U103,
    new_P1_R1171_U104, new_P1_R1171_U105, new_P1_R1171_U106,
    new_P1_R1171_U107, new_P1_R1171_U108, new_P1_R1171_U109,
    new_P1_R1171_U110, new_P1_R1171_U111, new_P1_R1171_U112,
    new_P1_R1171_U113, new_P1_R1171_U114, new_P1_R1171_U115,
    new_P1_R1171_U116, new_P1_R1171_U117, new_P1_R1171_U118,
    new_P1_R1171_U119, new_P1_R1171_U120, new_P1_R1171_U121,
    new_P1_R1171_U122, new_P1_R1171_U123, new_P1_R1171_U124,
    new_P1_R1171_U125, new_P1_R1171_U126, new_P1_R1171_U127,
    new_P1_R1171_U128, new_P1_R1171_U129, new_P1_R1171_U130,
    new_P1_R1171_U131, new_P1_R1171_U132, new_P1_R1171_U133,
    new_P1_R1171_U134, new_P1_R1171_U135, new_P1_R1171_U136,
    new_P1_R1171_U137, new_P1_R1171_U138, new_P1_R1171_U139,
    new_P1_R1171_U140, new_P1_R1171_U141, new_P1_R1171_U142,
    new_P1_R1171_U143, new_P1_R1171_U144, new_P1_R1171_U145,
    new_P1_R1171_U146, new_P1_R1171_U147, new_P1_R1171_U148,
    new_P1_R1171_U149, new_P1_R1171_U150, new_P1_R1171_U151,
    new_P1_R1171_U152, new_P1_R1171_U153, new_P1_R1171_U154,
    new_P1_R1171_U155, new_P1_R1171_U156, new_P1_R1171_U157,
    new_P1_R1171_U158, new_P1_R1171_U159, new_P1_R1171_U160,
    new_P1_R1171_U161, new_P1_R1171_U162, new_P1_R1171_U163,
    new_P1_R1171_U164, new_P1_R1171_U165, new_P1_R1171_U166,
    new_P1_R1171_U167, new_P1_R1171_U168, new_P1_R1171_U169,
    new_P1_R1171_U170, new_P1_R1171_U171, new_P1_R1171_U172,
    new_P1_R1171_U173, new_P1_R1171_U174, new_P1_R1171_U175,
    new_P1_R1171_U176, new_P1_R1171_U177, new_P1_R1171_U178,
    new_P1_R1171_U179, new_P1_R1171_U180, new_P1_R1171_U181,
    new_P1_R1171_U182, new_P1_R1171_U183, new_P1_R1171_U184,
    new_P1_R1171_U185, new_P1_R1171_U186, new_P1_R1171_U187,
    new_P1_R1171_U188, new_P1_R1171_U189, new_P1_R1171_U190,
    new_P1_R1171_U191, new_P1_R1171_U192, new_P1_R1171_U193,
    new_P1_R1171_U194, new_P1_R1171_U195, new_P1_R1171_U196,
    new_P1_R1171_U197, new_P1_R1171_U198, new_P1_R1171_U199,
    new_P1_R1171_U200, new_P1_R1171_U201, new_P1_R1171_U202,
    new_P1_R1171_U203, new_P1_R1171_U204, new_P1_R1171_U205,
    new_P1_R1171_U206, new_P1_R1171_U207, new_P1_R1171_U208,
    new_P1_R1171_U209, new_P1_R1171_U210, new_P1_R1171_U211,
    new_P1_R1171_U212, new_P1_R1171_U213, new_P1_R1171_U214,
    new_P1_R1171_U215, new_P1_R1171_U216, new_P1_R1171_U217,
    new_P1_R1171_U218, new_P1_R1171_U219, new_P1_R1171_U220,
    new_P1_R1171_U221, new_P1_R1171_U222, new_P1_R1171_U223,
    new_P1_R1171_U224, new_P1_R1171_U225, new_P1_R1171_U226,
    new_P1_R1171_U227, new_P1_R1171_U228, new_P1_R1171_U229,
    new_P1_R1171_U230, new_P1_R1171_U231, new_P1_R1171_U232,
    new_P1_R1171_U233, new_P1_R1171_U234, new_P1_R1171_U235,
    new_P1_R1171_U236, new_P1_R1171_U237, new_P1_R1171_U238,
    new_P1_R1171_U239, new_P1_R1171_U240, new_P1_R1171_U241,
    new_P1_R1171_U242, new_P1_R1171_U243, new_P1_R1171_U244,
    new_P1_R1171_U245, new_P1_R1171_U246, new_P1_R1171_U247,
    new_P1_R1171_U248, new_P1_R1171_U249, new_P1_R1171_U250,
    new_P1_R1171_U251, new_P1_R1171_U252, new_P1_R1171_U253,
    new_P1_R1171_U254, new_P1_R1171_U255, new_P1_R1171_U256,
    new_P1_R1171_U257, new_P1_R1171_U258, new_P1_R1171_U259,
    new_P1_R1171_U260, new_P1_R1171_U261, new_P1_R1171_U262,
    new_P1_R1171_U263, new_P1_R1171_U264, new_P1_R1171_U265,
    new_P1_R1171_U266, new_P1_R1171_U267, new_P1_R1171_U268,
    new_P1_R1171_U269, new_P1_R1171_U270, new_P1_R1171_U271,
    new_P1_R1171_U272, new_P1_R1171_U273, new_P1_R1171_U274,
    new_P1_R1171_U275, new_P1_R1171_U276, new_P1_R1171_U277,
    new_P1_R1171_U278, new_P1_R1171_U279, new_P1_R1171_U280,
    new_P1_R1171_U281, new_P1_R1171_U282, new_P1_R1171_U283,
    new_P1_R1171_U284, new_P1_R1171_U285, new_P1_R1171_U286,
    new_P1_R1171_U287, new_P1_R1171_U288, new_P1_R1171_U289,
    new_P1_R1171_U290, new_P1_R1171_U291, new_P1_R1171_U292,
    new_P1_R1171_U293, new_P1_R1171_U294, new_P1_R1171_U295,
    new_P1_R1171_U296, new_P1_R1171_U297, new_P1_R1171_U298,
    new_P1_R1171_U299, new_P1_R1171_U300, new_P1_R1171_U301,
    new_P1_R1171_U302, new_P1_R1171_U303, new_P1_R1171_U304,
    new_P1_R1171_U305, new_P1_R1171_U306, new_P1_R1171_U307,
    new_P1_R1171_U308, new_P1_R1171_U309, new_P1_R1171_U310,
    new_P1_R1171_U311, new_P1_R1171_U312, new_P1_R1171_U313,
    new_P1_R1171_U314, new_P1_R1171_U315, new_P1_R1171_U316,
    new_P1_R1171_U317, new_P1_R1171_U318, new_P1_R1171_U319,
    new_P1_R1171_U320, new_P1_R1171_U321, new_P1_R1171_U322,
    new_P1_R1171_U323, new_P1_R1171_U324, new_P1_R1171_U325,
    new_P1_R1171_U326, new_P1_R1171_U327, new_P1_R1171_U328,
    new_P1_R1171_U329, new_P1_R1171_U330, new_P1_R1171_U331,
    new_P1_R1171_U332, new_P1_R1171_U333, new_P1_R1171_U334,
    new_P1_R1171_U335, new_P1_R1171_U336, new_P1_R1171_U337,
    new_P1_R1171_U338, new_P1_R1171_U339, new_P1_R1171_U340,
    new_P1_R1171_U341, new_P1_R1171_U342, new_P1_R1171_U343,
    new_P1_R1171_U344, new_P1_R1171_U345, new_P1_R1171_U346,
    new_P1_R1171_U347, new_P1_R1171_U348, new_P1_R1171_U349,
    new_P1_R1171_U350, new_P1_R1171_U351, new_P1_R1171_U352,
    new_P1_R1171_U353, new_P1_R1171_U354, new_P1_R1171_U355,
    new_P1_R1171_U356, new_P1_R1171_U357, new_P1_R1171_U358,
    new_P1_R1171_U359, new_P1_R1171_U360, new_P1_R1171_U361,
    new_P1_R1171_U362, new_P1_R1171_U363, new_P1_R1171_U364,
    new_P1_R1171_U365, new_P1_R1171_U366, new_P1_R1171_U367,
    new_P1_R1171_U368, new_P1_R1171_U369, new_P1_R1171_U370,
    new_P1_R1171_U371, new_P1_R1171_U372, new_P1_R1171_U373,
    new_P1_R1171_U374, new_P1_R1171_U375, new_P1_R1171_U376,
    new_P1_R1171_U377, new_P1_R1171_U378, new_P1_R1171_U379,
    new_P1_R1171_U380, new_P1_R1171_U381, new_P1_R1171_U382,
    new_P1_R1171_U383, new_P1_R1171_U384, new_P1_R1171_U385,
    new_P1_R1171_U386, new_P1_R1171_U387, new_P1_R1171_U388,
    new_P1_R1171_U389, new_P1_R1171_U390, new_P1_R1171_U391,
    new_P1_R1171_U392, new_P1_R1171_U393, new_P1_R1171_U394,
    new_P1_R1171_U395, new_P1_R1171_U396, new_P1_R1171_U397,
    new_P1_R1171_U398, new_P1_R1171_U399, new_P1_R1171_U400,
    new_P1_R1171_U401, new_P1_R1171_U402, new_P1_R1171_U403,
    new_P1_R1171_U404, new_P1_R1171_U405, new_P1_R1171_U406,
    new_P1_R1171_U407, new_P1_R1171_U408, new_P1_R1171_U409,
    new_P1_R1171_U410, new_P1_R1171_U411, new_P1_R1171_U412,
    new_P1_R1171_U413, new_P1_R1171_U414, new_P1_R1171_U415,
    new_P1_R1171_U416, new_P1_R1171_U417, new_P1_R1171_U418,
    new_P1_R1171_U419, new_P1_R1171_U420, new_P1_R1171_U421,
    new_P1_R1171_U422, new_P1_R1171_U423, new_P1_R1171_U424,
    new_P1_R1171_U425, new_P1_R1171_U426, new_P1_R1171_U427,
    new_P1_R1171_U428, new_P1_R1171_U429, new_P1_R1171_U430,
    new_P1_R1171_U431, new_P1_R1171_U432, new_P1_R1171_U433,
    new_P1_R1171_U434, new_P1_R1171_U435, new_P1_R1171_U436,
    new_P1_R1171_U437, new_P1_R1171_U438, new_P1_R1171_U439,
    new_P1_R1171_U440, new_P1_R1171_U441, new_P1_R1171_U442,
    new_P1_R1171_U443, new_P1_R1171_U444, new_P1_R1171_U445,
    new_P1_R1171_U446, new_P1_R1171_U447, new_P1_R1171_U448,
    new_P1_R1171_U449, new_P1_R1171_U450, new_P1_R1171_U451,
    new_P1_R1171_U452, new_P1_R1171_U453, new_P1_R1171_U454,
    new_P1_R1171_U455, new_P1_R1171_U456, new_P1_R1171_U457,
    new_P1_R1171_U458, new_P1_R1171_U459, new_P1_R1171_U460,
    new_P1_R1171_U461, new_P1_R1171_U462, new_P1_R1171_U463,
    new_P1_R1171_U464, new_P1_R1171_U465, new_P1_R1171_U466,
    new_P1_R1171_U467, new_P1_R1171_U468, new_P1_R1171_U469,
    new_P1_R1171_U470, new_P1_R1171_U471, new_P1_R1171_U472,
    new_P1_R1171_U473, new_P1_R1171_U474, new_P1_R1171_U475,
    new_P1_R1171_U476, new_P1_R1171_U477, new_P1_R1171_U478,
    new_P1_R1171_U479, new_P1_R1171_U480, new_P1_R1171_U481,
    new_P1_R1171_U482, new_P1_R1171_U483, new_P1_R1171_U484,
    new_P1_R1171_U485, new_P1_R1171_U486, new_P1_R1171_U487,
    new_P1_R1171_U488, new_P1_R1171_U489, new_P1_R1171_U490,
    new_P1_R1171_U491, new_P1_R1171_U492, new_P1_R1171_U493,
    new_P1_R1171_U494, new_P1_R1171_U495, new_P1_R1171_U496,
    new_P1_R1171_U497, new_P1_R1171_U498, new_P1_R1171_U499,
    new_P1_R1171_U500, new_P1_R1171_U501, new_P1_R1171_U502,
    new_P1_R1171_U503, new_P1_R1138_U4, new_P1_R1138_U5, new_P1_R1138_U6,
    new_P1_R1138_U7, new_P1_R1138_U8, new_P1_R1138_U9, new_P1_R1138_U10,
    new_P1_R1138_U11, new_P1_R1138_U12, new_P1_R1138_U13, new_P1_R1138_U14,
    new_P1_R1138_U15, new_P1_R1138_U16, new_P1_R1138_U17, new_P1_R1138_U18,
    new_P1_R1138_U19, new_P1_R1138_U20, new_P1_R1138_U21, new_P1_R1138_U22,
    new_P1_R1138_U23, new_P1_R1138_U24, new_P1_R1138_U25, new_P1_R1138_U26,
    new_P1_R1138_U27, new_P1_R1138_U28, new_P1_R1138_U29, new_P1_R1138_U30,
    new_P1_R1138_U31, new_P1_R1138_U32, new_P1_R1138_U33, new_P1_R1138_U34,
    new_P1_R1138_U35, new_P1_R1138_U36, new_P1_R1138_U37, new_P1_R1138_U38,
    new_P1_R1138_U39, new_P1_R1138_U40, new_P1_R1138_U41, new_P1_R1138_U42,
    new_P1_R1138_U43, new_P1_R1138_U44, new_P1_R1138_U45, new_P1_R1138_U46,
    new_P1_R1138_U47, new_P1_R1138_U48, new_P1_R1138_U49, new_P1_R1138_U50,
    new_P1_R1138_U51, new_P1_R1138_U52, new_P1_R1138_U53, new_P1_R1138_U54,
    new_P1_R1138_U55, new_P1_R1138_U56, new_P1_R1138_U57, new_P1_R1138_U58,
    new_P1_R1138_U59, new_P1_R1138_U60, new_P1_R1138_U61, new_P1_R1138_U62,
    new_P1_R1138_U63, new_P1_R1138_U64, new_P1_R1138_U65, new_P1_R1138_U66,
    new_P1_R1138_U67, new_P1_R1138_U68, new_P1_R1138_U69, new_P1_R1138_U70,
    new_P1_R1138_U71, new_P1_R1138_U72, new_P1_R1138_U73, new_P1_R1138_U74,
    new_P1_R1138_U75, new_P1_R1138_U76, new_P1_R1138_U77, new_P1_R1138_U78,
    new_P1_R1138_U79, new_P1_R1138_U80, new_P1_R1138_U81, new_P1_R1138_U82,
    new_P1_R1138_U83, new_P1_R1138_U84, new_P1_R1138_U85, new_P1_R1138_U86,
    new_P1_R1138_U87, new_P1_R1138_U88, new_P1_R1138_U89, new_P1_R1138_U90,
    new_P1_R1138_U91, new_P1_R1138_U92, new_P1_R1138_U93, new_P1_R1138_U94,
    new_P1_R1138_U95, new_P1_R1138_U96, new_P1_R1138_U97, new_P1_R1138_U98,
    new_P1_R1138_U99, new_P1_R1138_U100, new_P1_R1138_U101,
    new_P1_R1138_U102, new_P1_R1138_U103, new_P1_R1138_U104,
    new_P1_R1138_U105, new_P1_R1138_U106, new_P1_R1138_U107,
    new_P1_R1138_U108, new_P1_R1138_U109, new_P1_R1138_U110,
    new_P1_R1138_U111, new_P1_R1138_U112, new_P1_R1138_U113,
    new_P1_R1138_U114, new_P1_R1138_U115, new_P1_R1138_U116,
    new_P1_R1138_U117, new_P1_R1138_U118, new_P1_R1138_U119,
    new_P1_R1138_U120, new_P1_R1138_U121, new_P1_R1138_U122,
    new_P1_R1138_U123, new_P1_R1138_U124, new_P1_R1138_U125,
    new_P1_R1138_U126, new_P1_R1138_U127, new_P1_R1138_U128,
    new_P1_R1138_U129, new_P1_R1138_U130, new_P1_R1138_U131,
    new_P1_R1138_U132, new_P1_R1138_U133, new_P1_R1138_U134,
    new_P1_R1138_U135, new_P1_R1138_U136, new_P1_R1138_U137,
    new_P1_R1138_U138, new_P1_R1138_U139, new_P1_R1138_U140,
    new_P1_R1138_U141, new_P1_R1138_U142, new_P1_R1138_U143,
    new_P1_R1138_U144, new_P1_R1138_U145, new_P1_R1138_U146,
    new_P1_R1138_U147, new_P1_R1138_U148, new_P1_R1138_U149,
    new_P1_R1138_U150, new_P1_R1138_U151, new_P1_R1138_U152,
    new_P1_R1138_U153, new_P1_R1138_U154, new_P1_R1138_U155,
    new_P1_R1138_U156, new_P1_R1138_U157, new_P1_R1138_U158,
    new_P1_R1138_U159, new_P1_R1138_U160, new_P1_R1138_U161,
    new_P1_R1138_U162, new_P1_R1138_U163, new_P1_R1138_U164,
    new_P1_R1138_U165, new_P1_R1138_U166, new_P1_R1138_U167,
    new_P1_R1138_U168, new_P1_R1138_U169, new_P1_R1138_U170,
    new_P1_R1138_U171, new_P1_R1138_U172, new_P1_R1138_U173,
    new_P1_R1138_U174, new_P1_R1138_U175, new_P1_R1138_U176,
    new_P1_R1138_U177, new_P1_R1138_U178, new_P1_R1138_U179,
    new_P1_R1138_U180, new_P1_R1138_U181, new_P1_R1138_U182,
    new_P1_R1138_U183, new_P1_R1138_U184, new_P1_R1138_U185,
    new_P1_R1138_U186, new_P1_R1138_U187, new_P1_R1138_U188,
    new_P1_R1138_U189, new_P1_R1138_U190, new_P1_R1138_U191,
    new_P1_R1138_U192, new_P1_R1138_U193, new_P1_R1138_U194,
    new_P1_R1138_U195, new_P1_R1138_U196, new_P1_R1138_U197,
    new_P1_R1138_U198, new_P1_R1138_U199, new_P1_R1138_U200,
    new_P1_R1138_U201, new_P1_R1138_U202, new_P1_R1138_U203,
    new_P1_R1138_U204, new_P1_R1138_U205, new_P1_R1138_U206,
    new_P1_R1138_U207, new_P1_R1138_U208, new_P1_R1138_U209,
    new_P1_R1138_U210, new_P1_R1138_U211, new_P1_R1138_U212,
    new_P1_R1138_U213, new_P1_R1138_U214, new_P1_R1138_U215,
    new_P1_R1138_U216, new_P1_R1138_U217, new_P1_R1138_U218,
    new_P1_R1138_U219, new_P1_R1138_U220, new_P1_R1138_U221,
    new_P1_R1138_U222, new_P1_R1138_U223, new_P1_R1138_U224,
    new_P1_R1138_U225, new_P1_R1138_U226, new_P1_R1138_U227,
    new_P1_R1138_U228, new_P1_R1138_U229, new_P1_R1138_U230,
    new_P1_R1138_U231, new_P1_R1138_U232, new_P1_R1138_U233,
    new_P1_R1138_U234, new_P1_R1138_U235, new_P1_R1138_U236,
    new_P1_R1138_U237, new_P1_R1138_U238, new_P1_R1138_U239,
    new_P1_R1138_U240, new_P1_R1138_U241, new_P1_R1138_U242,
    new_P1_R1138_U243, new_P1_R1138_U244, new_P1_R1138_U245,
    new_P1_R1138_U246, new_P1_R1138_U247, new_P1_R1138_U248,
    new_P1_R1138_U249, new_P1_R1138_U250, new_P1_R1138_U251,
    new_P1_R1138_U252, new_P1_R1138_U253, new_P1_R1138_U254,
    new_P1_R1138_U255, new_P1_R1138_U256, new_P1_R1138_U257,
    new_P1_R1138_U258, new_P1_R1138_U259, new_P1_R1138_U260,
    new_P1_R1138_U261, new_P1_R1138_U262, new_P1_R1138_U263,
    new_P1_R1138_U264, new_P1_R1138_U265, new_P1_R1138_U266,
    new_P1_R1138_U267, new_P1_R1138_U268, new_P1_R1138_U269,
    new_P1_R1138_U270, new_P1_R1138_U271, new_P1_R1138_U272,
    new_P1_R1138_U273, new_P1_R1138_U274, new_P1_R1138_U275,
    new_P1_R1138_U276, new_P1_R1138_U277, new_P1_R1138_U278,
    new_P1_R1138_U279, new_P1_R1138_U280, new_P1_R1138_U281,
    new_P1_R1138_U282, new_P1_R1138_U283, new_P1_R1138_U284,
    new_P1_R1138_U285, new_P1_R1138_U286, new_P1_R1138_U287,
    new_P1_R1138_U288, new_P1_R1138_U289, new_P1_R1138_U290,
    new_P1_R1138_U291, new_P1_R1138_U292, new_P1_R1138_U293,
    new_P1_R1138_U294, new_P1_R1138_U295, new_P1_R1138_U296,
    new_P1_R1138_U297, new_P1_R1138_U298, new_P1_R1138_U299,
    new_P1_R1138_U300, new_P1_R1138_U301, new_P1_R1138_U302,
    new_P1_R1138_U303, new_P1_R1138_U304, new_P1_R1138_U305,
    new_P1_R1138_U306, new_P1_R1138_U307, new_P1_R1138_U308,
    new_P1_R1138_U309, new_P1_R1138_U310, new_P1_R1138_U311,
    new_P1_R1138_U312, new_P1_R1138_U313, new_P1_R1138_U314,
    new_P1_R1138_U315, new_P1_R1138_U316, new_P1_R1138_U317,
    new_P1_R1138_U318, new_P1_R1138_U319, new_P1_R1138_U320,
    new_P1_R1138_U321, new_P1_R1138_U322, new_P1_R1138_U323,
    new_P1_R1138_U324, new_P1_R1138_U325, new_P1_R1138_U326,
    new_P1_R1138_U327, new_P1_R1138_U328, new_P1_R1138_U329,
    new_P1_R1138_U330, new_P1_R1138_U331, new_P1_R1138_U332,
    new_P1_R1138_U333, new_P1_R1138_U334, new_P1_R1138_U335,
    new_P1_R1138_U336, new_P1_R1138_U337, new_P1_R1138_U338,
    new_P1_R1138_U339, new_P1_R1138_U340, new_P1_R1138_U341,
    new_P1_R1138_U342, new_P1_R1138_U343, new_P1_R1138_U344,
    new_P1_R1138_U345, new_P1_R1138_U346, new_P1_R1138_U347,
    new_P1_R1138_U348, new_P1_R1138_U349, new_P1_R1138_U350,
    new_P1_R1138_U351, new_P1_R1138_U352, new_P1_R1138_U353,
    new_P1_R1138_U354, new_P1_R1138_U355, new_P1_R1138_U356,
    new_P1_R1138_U357, new_P1_R1138_U358, new_P1_R1138_U359,
    new_P1_R1138_U360, new_P1_R1138_U361, new_P1_R1138_U362,
    new_P1_R1138_U363, new_P1_R1138_U364, new_P1_R1138_U365,
    new_P1_R1138_U366, new_P1_R1138_U367, new_P1_R1138_U368,
    new_P1_R1138_U369, new_P1_R1138_U370, new_P1_R1138_U371,
    new_P1_R1138_U372, new_P1_R1138_U373, new_P1_R1138_U374,
    new_P1_R1138_U375, new_P1_R1138_U376, new_P1_R1138_U377,
    new_P1_R1138_U378, new_P1_R1138_U379, new_P1_R1138_U380,
    new_P1_R1138_U381, new_P1_R1138_U382, new_P1_R1138_U383,
    new_P1_R1138_U384, new_P1_R1138_U385, new_P1_R1138_U386,
    new_P1_R1138_U387, new_P1_R1138_U388, new_P1_R1138_U389,
    new_P1_R1138_U390, new_P1_R1138_U391, new_P1_R1138_U392,
    new_P1_R1138_U393, new_P1_R1138_U394, new_P1_R1138_U395,
    new_P1_R1138_U396, new_P1_R1138_U397, new_P1_R1138_U398,
    new_P1_R1138_U399, new_P1_R1138_U400, new_P1_R1138_U401,
    new_P1_R1138_U402, new_P1_R1138_U403, new_P1_R1138_U404,
    new_P1_R1138_U405, new_P1_R1138_U406, new_P1_R1138_U407,
    new_P1_R1138_U408, new_P1_R1138_U409, new_P1_R1138_U410,
    new_P1_R1138_U411, new_P1_R1138_U412, new_P1_R1138_U413,
    new_P1_R1138_U414, new_P1_R1138_U415, new_P1_R1138_U416,
    new_P1_R1138_U417, new_P1_R1138_U418, new_P1_R1138_U419,
    new_P1_R1138_U420, new_P1_R1138_U421, new_P1_R1138_U422,
    new_P1_R1138_U423, new_P1_R1138_U424, new_P1_R1138_U425,
    new_P1_R1138_U426, new_P1_R1138_U427, new_P1_R1138_U428,
    new_P1_R1138_U429, new_P1_R1138_U430, new_P1_R1138_U431,
    new_P1_R1138_U432, new_P1_R1138_U433, new_P1_R1138_U434,
    new_P1_R1138_U435, new_P1_R1138_U436, new_P1_R1138_U437,
    new_P1_R1138_U438, new_P1_R1138_U439, new_P1_R1138_U440,
    new_P1_R1138_U441, new_P1_R1138_U442, new_P1_R1138_U443,
    new_P1_R1138_U444, new_P1_R1138_U445, new_P1_R1138_U446,
    new_P1_R1138_U447, new_P1_R1138_U448, new_P1_R1138_U449,
    new_P1_R1138_U450, new_P1_R1138_U451, new_P1_R1138_U452,
    new_P1_R1138_U453, new_P1_R1138_U454, new_P1_R1138_U455,
    new_P1_R1138_U456, new_P1_R1138_U457, new_P1_R1138_U458,
    new_P1_R1138_U459, new_P1_R1138_U460, new_P1_R1138_U461,
    new_P1_R1138_U462, new_P1_R1138_U463, new_P1_R1138_U464,
    new_P1_R1138_U465, new_P1_R1138_U466, new_P1_R1138_U467,
    new_P1_R1138_U468, new_P1_R1138_U469, new_P1_R1138_U470,
    new_P1_R1138_U471, new_P1_R1138_U472, new_P1_R1138_U473,
    new_P1_R1138_U474, new_P1_R1138_U475, new_P1_R1138_U476,
    new_P1_R1138_U477, new_P1_R1138_U478, new_P1_R1138_U479,
    new_P1_R1138_U480, new_P1_R1138_U481, new_P1_R1138_U482,
    new_P1_R1138_U483, new_P1_R1138_U484, new_P1_R1138_U485,
    new_P1_R1138_U486, new_P1_R1138_U487, new_P1_R1138_U488,
    new_P1_R1138_U489, new_P1_R1138_U490, new_P1_R1138_U491,
    new_P1_R1138_U492, new_P1_R1138_U493, new_P1_R1138_U494,
    new_P1_R1138_U495, new_P1_R1138_U496, new_P1_R1138_U497,
    new_P1_R1138_U498, new_P1_R1138_U499, new_P1_R1138_U500,
    new_P1_R1138_U501, new_P1_R1138_U502, new_P1_R1138_U503,
    new_P1_R1222_U4, new_P1_R1222_U5, new_P1_R1222_U6, new_P1_R1222_U7,
    new_P1_R1222_U8, new_P1_R1222_U9, new_P1_R1222_U10, new_P1_R1222_U11,
    new_P1_R1222_U12, new_P1_R1222_U13, new_P1_R1222_U14, new_P1_R1222_U15,
    new_P1_R1222_U16, new_P1_R1222_U17, new_P1_R1222_U18, new_P1_R1222_U19,
    new_P1_R1222_U20, new_P1_R1222_U21, new_P1_R1222_U22, new_P1_R1222_U23,
    new_P1_R1222_U24, new_P1_R1222_U25, new_P1_R1222_U26, new_P1_R1222_U27,
    new_P1_R1222_U28, new_P1_R1222_U29, new_P1_R1222_U30, new_P1_R1222_U31,
    new_P1_R1222_U32, new_P1_R1222_U33, new_P1_R1222_U34, new_P1_R1222_U35,
    new_P1_R1222_U36, new_P1_R1222_U37, new_P1_R1222_U38, new_P1_R1222_U39,
    new_P1_R1222_U40, new_P1_R1222_U41, new_P1_R1222_U42, new_P1_R1222_U43,
    new_P1_R1222_U44, new_P1_R1222_U45, new_P1_R1222_U46, new_P1_R1222_U47,
    new_P1_R1222_U48, new_P1_R1222_U49, new_P1_R1222_U50, new_P1_R1222_U51,
    new_P1_R1222_U52, new_P1_R1222_U53, new_P1_R1222_U54, new_P1_R1222_U55,
    new_P1_R1222_U56, new_P1_R1222_U57, new_P1_R1222_U58, new_P1_R1222_U59,
    new_P1_R1222_U60, new_P1_R1222_U61, new_P1_R1222_U62, new_P1_R1222_U63,
    new_P1_R1222_U64, new_P1_R1222_U65, new_P1_R1222_U66, new_P1_R1222_U67,
    new_P1_R1222_U68, new_P1_R1222_U69, new_P1_R1222_U70, new_P1_R1222_U71,
    new_P1_R1222_U72, new_P1_R1222_U73, new_P1_R1222_U74, new_P1_R1222_U75,
    new_P1_R1222_U76, new_P1_R1222_U77, new_P1_R1222_U78, new_P1_R1222_U79,
    new_P1_R1222_U80, new_P1_R1222_U81, new_P1_R1222_U82, new_P1_R1222_U83,
    new_P1_R1222_U84, new_P1_R1222_U85, new_P1_R1222_U86, new_P1_R1222_U87,
    new_P1_R1222_U88, new_P1_R1222_U89, new_P1_R1222_U90, new_P1_R1222_U91,
    new_P1_R1222_U92, new_P1_R1222_U93, new_P1_R1222_U94, new_P1_R1222_U95,
    new_P1_R1222_U96, new_P1_R1222_U97, new_P1_R1222_U98, new_P1_R1222_U99,
    new_P1_R1222_U100, new_P1_R1222_U101, new_P1_R1222_U102,
    new_P1_R1222_U103, new_P1_R1222_U104, new_P1_R1222_U105,
    new_P1_R1222_U106, new_P1_R1222_U107, new_P1_R1222_U108,
    new_P1_R1222_U109, new_P1_R1222_U110, new_P1_R1222_U111,
    new_P1_R1222_U112, new_P1_R1222_U113, new_P1_R1222_U114,
    new_P1_R1222_U115, new_P1_R1222_U116, new_P1_R1222_U117,
    new_P1_R1222_U118, new_P1_R1222_U119, new_P1_R1222_U120,
    new_P1_R1222_U121, new_P1_R1222_U122, new_P1_R1222_U123,
    new_P1_R1222_U124, new_P1_R1222_U125, new_P1_R1222_U126,
    new_P1_R1222_U127, new_P1_R1222_U128, new_P1_R1222_U129,
    new_P1_R1222_U130, new_P1_R1222_U131, new_P1_R1222_U132,
    new_P1_R1222_U133, new_P1_R1222_U134, new_P1_R1222_U135,
    new_P1_R1222_U136, new_P1_R1222_U137, new_P1_R1222_U138,
    new_P1_R1222_U139, new_P1_R1222_U140, new_P1_R1222_U141,
    new_P1_R1222_U142, new_P1_R1222_U143, new_P1_R1222_U144,
    new_P1_R1222_U145, new_P1_R1222_U146, new_P1_R1222_U147,
    new_P1_R1222_U148, new_P1_R1222_U149, new_P1_R1222_U150,
    new_P1_R1222_U151, new_P1_R1222_U152, new_P1_R1222_U153,
    new_P1_R1222_U154, new_P1_R1222_U155, new_P1_R1222_U156,
    new_P1_R1222_U157, new_P1_R1222_U158, new_P1_R1222_U159,
    new_P1_R1222_U160, new_P1_R1222_U161, new_P1_R1222_U162,
    new_P1_R1222_U163, new_P1_R1222_U164, new_P1_R1222_U165,
    new_P1_R1222_U166, new_P1_R1222_U167, new_P1_R1222_U168,
    new_P1_R1222_U169, new_P1_R1222_U170, new_P1_R1222_U171,
    new_P1_R1222_U172, new_P1_R1222_U173, new_P1_R1222_U174,
    new_P1_R1222_U175, new_P1_R1222_U176, new_P1_R1222_U177,
    new_P1_R1222_U178, new_P1_R1222_U179, new_P1_R1222_U180,
    new_P1_R1222_U181, new_P1_R1222_U182, new_P1_R1222_U183,
    new_P1_R1222_U184, new_P1_R1222_U185, new_P1_R1222_U186,
    new_P1_R1222_U187, new_P1_R1222_U188, new_P1_R1222_U189,
    new_P1_R1222_U190, new_P1_R1222_U191, new_P1_R1222_U192,
    new_P1_R1222_U193, new_P1_R1222_U194, new_P1_R1222_U195,
    new_P1_R1222_U196, new_P1_R1222_U197, new_P1_R1222_U198,
    new_P1_R1222_U199, new_P1_R1222_U200, new_P1_R1222_U201,
    new_P1_R1222_U202, new_P1_R1222_U203, new_P1_R1222_U204,
    new_P1_R1222_U205, new_P1_R1222_U206, new_P1_R1222_U207,
    new_P1_R1222_U208, new_P1_R1222_U209, new_P1_R1222_U210,
    new_P1_R1222_U211, new_P1_R1222_U212, new_P1_R1222_U213,
    new_P1_R1222_U214, new_P1_R1222_U215, new_P1_R1222_U216,
    new_P1_R1222_U217, new_P1_R1222_U218, new_P1_R1222_U219,
    new_P1_R1222_U220, new_P1_R1222_U221, new_P1_R1222_U222,
    new_P1_R1222_U223, new_P1_R1222_U224, new_P1_R1222_U225,
    new_P1_R1222_U226, new_P1_R1222_U227, new_P1_R1222_U228,
    new_P1_R1222_U229, new_P1_R1222_U230, new_P1_R1222_U231,
    new_P1_R1222_U232, new_P1_R1222_U233, new_P1_R1222_U234,
    new_P1_R1222_U235, new_P1_R1222_U236, new_P1_R1222_U237,
    new_P1_R1222_U238, new_P1_R1222_U239, new_P1_R1222_U240,
    new_P1_R1222_U241, new_P1_R1222_U242, new_P1_R1222_U243,
    new_P1_R1222_U244, new_P1_R1222_U245, new_P1_R1222_U246,
    new_P1_R1222_U247, new_P1_R1222_U248, new_P1_R1222_U249,
    new_P1_R1222_U250, new_P1_R1222_U251, new_P1_R1222_U252,
    new_P1_R1222_U253, new_P1_R1222_U254, new_P1_R1222_U255,
    new_P1_R1222_U256, new_P1_R1222_U257, new_P1_R1222_U258,
    new_P1_R1222_U259, new_P1_R1222_U260, new_P1_R1222_U261,
    new_P1_R1222_U262, new_P1_R1222_U263, new_P1_R1222_U264,
    new_P1_R1222_U265, new_P1_R1222_U266, new_P1_R1222_U267,
    new_P1_R1222_U268, new_P1_R1222_U269, new_P1_R1222_U270,
    new_P1_R1222_U271, new_P1_R1222_U272, new_P1_R1222_U273,
    new_P1_R1222_U274, new_P1_R1222_U275, new_P1_R1222_U276,
    new_P1_R1222_U277, new_P1_R1222_U278, new_P1_R1222_U279,
    new_P1_R1222_U280, new_P1_R1222_U281, new_P1_R1222_U282,
    new_P1_R1222_U283, new_P1_R1222_U284, new_P1_R1222_U285,
    new_P1_R1222_U286, new_P1_R1222_U287, new_P1_R1222_U288,
    new_P1_R1222_U289, new_P1_R1222_U290, new_P1_R1222_U291,
    new_P1_R1222_U292, new_P1_R1222_U293, new_P1_R1222_U294,
    new_P1_R1222_U295, new_P1_R1222_U296, new_P1_R1222_U297,
    new_P1_R1222_U298, new_P1_R1222_U299, new_P1_R1222_U300,
    new_P1_R1222_U301, new_P1_R1222_U302, new_P1_R1222_U303,
    new_P1_R1222_U304, new_P1_R1222_U305, new_P1_R1222_U306,
    new_P1_R1222_U307, new_P1_R1222_U308, new_P1_R1222_U309,
    new_P1_R1222_U310, new_P1_R1222_U311, new_P1_R1222_U312,
    new_P1_R1222_U313, new_P1_R1222_U314, new_P1_R1222_U315,
    new_P1_R1222_U316, new_P1_R1222_U317, new_P1_R1222_U318,
    new_P1_R1222_U319, new_P1_R1222_U320, new_P1_R1222_U321,
    new_P1_R1222_U322, new_P1_R1222_U323, new_P1_R1222_U324,
    new_P1_R1222_U325, new_P1_R1222_U326, new_P1_R1222_U327,
    new_P1_R1222_U328, new_P1_R1222_U329, new_P1_R1222_U330,
    new_P1_R1222_U331, new_P1_R1222_U332, new_P1_R1222_U333,
    new_P1_R1222_U334, new_P1_R1222_U335, new_P1_R1222_U336,
    new_P1_R1222_U337, new_P1_R1222_U338, new_P1_R1222_U339,
    new_P1_R1222_U340, new_P1_R1222_U341, new_P1_R1222_U342,
    new_P1_R1222_U343, new_P1_R1222_U344, new_P1_R1222_U345,
    new_P1_R1222_U346, new_P1_R1222_U347, new_P1_R1222_U348,
    new_P1_R1222_U349, new_P1_R1222_U350, new_P1_R1222_U351,
    new_P1_R1222_U352, new_P1_R1222_U353, new_P1_R1222_U354,
    new_P1_R1222_U355, new_P1_R1222_U356, new_P1_R1222_U357,
    new_P1_R1222_U358, new_P1_R1222_U359, new_P1_R1222_U360,
    new_P1_R1222_U361, new_P1_R1222_U362, new_P1_R1222_U363,
    new_P1_R1222_U364, new_P1_R1222_U365, new_P1_R1222_U366,
    new_P1_R1222_U367, new_P1_R1222_U368, new_P1_R1222_U369,
    new_P1_R1222_U370, new_P1_R1222_U371, new_P1_R1222_U372,
    new_P1_R1222_U373, new_P1_R1222_U374, new_P1_R1222_U375,
    new_P1_R1222_U376, new_P1_R1222_U377, new_P1_R1222_U378,
    new_P1_R1222_U379, new_P1_R1222_U380, new_P1_R1222_U381,
    new_P1_R1222_U382, new_P1_R1222_U383, new_P1_R1222_U384,
    new_P1_R1222_U385, new_P1_R1222_U386, new_P1_R1222_U387,
    new_P1_R1222_U388, new_P1_R1222_U389, new_P1_R1222_U390,
    new_P1_R1222_U391, new_P1_R1222_U392, new_P1_R1222_U393,
    new_P1_R1222_U394, new_P1_R1222_U395, new_P1_R1222_U396,
    new_P1_R1222_U397, new_P1_R1222_U398, new_P1_R1222_U399,
    new_P1_R1222_U400, new_P1_R1222_U401, new_P1_R1222_U402,
    new_P1_R1222_U403, new_P1_R1222_U404, new_P1_R1222_U405,
    new_P1_R1222_U406, new_P1_R1222_U407, new_P1_R1222_U408,
    new_P1_R1222_U409, new_P1_R1222_U410, new_P1_R1222_U411,
    new_P1_R1222_U412, new_P1_R1222_U413, new_P1_R1222_U414,
    new_P1_R1222_U415, new_P1_R1222_U416, new_P1_R1222_U417,
    new_P1_R1222_U418, new_P1_R1222_U419, new_P1_R1222_U420,
    new_P1_R1222_U421, new_P1_R1222_U422, new_P1_R1222_U423,
    new_P1_R1222_U424, new_P1_R1222_U425, new_P1_R1222_U426,
    new_P1_R1222_U427, new_P1_R1222_U428, new_P1_R1222_U429,
    new_P1_R1222_U430, new_P1_R1222_U431, new_P1_R1222_U432,
    new_P1_R1222_U433, new_P1_R1222_U434, new_P1_R1222_U435,
    new_P1_R1222_U436, new_P1_R1222_U437, new_P1_R1222_U438,
    new_P1_R1222_U439, new_P1_R1222_U440, new_P1_R1222_U441,
    new_P1_R1222_U442, new_P1_R1222_U443, new_P1_R1222_U444,
    new_P1_R1222_U445, new_P1_R1222_U446, new_P1_R1222_U447,
    new_P1_R1222_U448, new_P1_R1222_U449, new_P1_R1222_U450,
    new_P1_R1222_U451, new_P1_R1222_U452, new_P1_R1222_U453,
    new_P1_R1222_U454, new_P1_R1222_U455, new_P1_R1222_U456,
    new_P1_R1222_U457, new_P1_R1222_U458, new_P1_R1222_U459,
    new_P1_R1222_U460, new_P1_R1222_U461, new_P1_R1222_U462,
    new_P1_R1222_U463, new_P1_R1222_U464, new_P1_R1222_U465,
    new_P1_R1222_U466, new_P1_R1222_U467, new_P1_R1222_U468,
    new_P1_R1222_U469, new_P1_R1222_U470, new_P1_R1222_U471,
    new_P1_R1222_U472, new_P1_R1222_U473, new_P1_R1222_U474,
    new_P1_R1222_U475, new_P1_R1222_U476, new_P1_R1222_U477,
    new_P1_R1222_U478, new_P1_R1222_U479, new_P1_R1222_U480,
    new_P1_R1222_U481, new_P1_R1222_U482, new_P1_R1222_U483,
    new_P1_R1222_U484, new_P1_R1222_U485, new_P1_R1222_U486,
    new_P1_R1222_U487, new_P1_R1222_U488, new_P1_R1222_U489,
    new_P1_R1222_U490, new_P1_R1222_U491, new_P1_R1222_U492,
    new_P1_R1222_U493, new_P1_R1222_U494, new_P1_R1222_U495,
    new_P1_R1222_U496, new_P1_R1222_U497, new_P1_R1222_U498,
    new_P1_R1222_U499, new_P1_R1222_U500, new_P1_R1222_U501,
    new_P1_R1222_U502, new_P1_R1222_U503, new_P2_SUB_594_U6,
    new_P2_SUB_594_U7, new_P2_SUB_594_U8, new_P2_SUB_594_U9,
    new_P2_SUB_594_U10, new_P2_SUB_594_U11, new_P2_SUB_594_U12,
    new_P2_SUB_594_U13, new_P2_SUB_594_U14, new_P2_SUB_594_U15,
    new_P2_SUB_594_U16, new_P2_SUB_594_U17, new_P2_SUB_594_U18,
    new_P2_SUB_594_U19, new_P2_SUB_594_U20, new_P2_SUB_594_U21,
    new_P2_SUB_594_U22, new_P2_SUB_594_U23, new_P2_SUB_594_U24,
    new_P2_SUB_594_U25, new_P2_SUB_594_U26, new_P2_SUB_594_U27,
    new_P2_SUB_594_U28, new_P2_SUB_594_U29, new_P2_SUB_594_U30,
    new_P2_SUB_594_U31, new_P2_SUB_594_U32, new_P2_SUB_594_U33,
    new_P2_SUB_594_U34, new_P2_SUB_594_U35, new_P2_SUB_594_U36,
    new_P2_SUB_594_U37, new_P2_SUB_594_U38, new_P2_SUB_594_U39,
    new_P2_SUB_594_U40, new_P2_SUB_594_U41, new_P2_SUB_594_U42,
    new_P2_SUB_594_U43, new_P2_SUB_594_U44, new_P2_SUB_594_U45,
    new_P2_SUB_594_U46, new_P2_SUB_594_U47, new_P2_SUB_594_U48,
    new_P2_SUB_594_U49, new_P2_SUB_594_U50, new_P2_SUB_594_U51,
    new_P2_SUB_594_U52, new_P2_SUB_594_U53, new_P2_SUB_594_U54,
    new_P2_SUB_594_U55, new_P2_SUB_594_U56, new_P2_SUB_594_U57,
    new_P2_SUB_594_U58, new_P2_SUB_594_U59, new_P2_SUB_594_U60,
    new_P2_SUB_594_U61, new_P2_SUB_594_U62, new_P2_SUB_594_U63,
    new_P2_SUB_594_U64, new_P2_SUB_594_U65, new_P2_SUB_594_U66,
    new_P2_SUB_594_U67, new_P2_SUB_594_U68, new_P2_SUB_594_U69,
    new_P2_SUB_594_U70, new_P2_SUB_594_U71, new_P2_SUB_594_U72,
    new_P2_SUB_594_U73, new_P2_SUB_594_U74, new_P2_SUB_594_U75,
    new_P2_SUB_594_U76, new_P2_SUB_594_U77, new_P2_SUB_594_U78,
    new_P2_SUB_594_U79, new_P2_SUB_594_U80, new_P2_SUB_594_U81,
    new_P2_SUB_594_U82, new_P2_SUB_594_U83, new_P2_SUB_594_U84,
    new_P2_SUB_594_U85, new_P2_SUB_594_U86, new_P2_SUB_594_U87,
    new_P2_SUB_594_U88, new_P2_SUB_594_U89, new_P2_SUB_594_U90,
    new_P2_SUB_594_U91, new_P2_SUB_594_U92, new_P2_SUB_594_U93,
    new_P2_SUB_594_U94, new_P2_SUB_594_U95, new_P2_SUB_594_U96,
    new_P2_SUB_594_U97, new_P2_SUB_594_U98, new_P2_SUB_594_U99,
    new_P2_SUB_594_U100, new_P2_SUB_594_U101, new_P2_SUB_594_U102,
    new_P2_SUB_594_U103, new_P2_SUB_594_U104, new_P2_SUB_594_U105,
    new_P2_SUB_594_U106, new_P2_SUB_594_U107, new_P2_SUB_594_U108,
    new_P2_SUB_594_U109, new_P2_SUB_594_U110, new_P2_SUB_594_U111,
    new_P2_SUB_594_U112, new_P2_SUB_594_U113, new_P2_SUB_594_U114,
    new_P2_SUB_594_U115, new_P2_SUB_594_U116, new_P2_SUB_594_U117,
    new_P2_SUB_594_U118, new_P2_SUB_594_U119, new_P2_SUB_594_U120,
    new_P2_SUB_594_U121, new_P2_SUB_594_U122, new_P2_SUB_594_U123,
    new_P2_SUB_594_U124, new_P2_SUB_594_U125, new_P2_SUB_594_U126,
    new_P2_SUB_594_U127, new_P2_SUB_594_U128, new_P2_SUB_594_U129,
    new_P2_SUB_594_U130, new_P2_SUB_594_U131, new_P2_SUB_594_U132,
    new_P2_SUB_594_U133, new_P2_SUB_594_U134, new_P2_SUB_594_U135,
    new_P2_SUB_594_U136, new_P2_SUB_594_U137, new_P2_SUB_594_U138,
    new_P2_SUB_594_U139, new_P2_SUB_594_U140, new_P2_SUB_594_U141,
    new_P2_SUB_594_U142, new_P2_SUB_594_U143, new_P2_SUB_594_U144,
    new_P2_SUB_594_U145, new_P2_SUB_594_U146, new_P2_SUB_594_U147,
    new_P2_SUB_594_U148, new_P2_SUB_594_U149, new_P2_SUB_594_U150,
    new_P2_SUB_594_U151, new_P2_SUB_594_U152, new_P2_SUB_594_U153,
    new_P2_SUB_594_U154, new_P2_SUB_594_U155, new_P2_SUB_594_U156,
    new_P2_SUB_594_U157, new_P2_SUB_594_U158, new_P2_R693_U6,
    new_P2_R693_U7, new_P2_R693_U8, new_P2_R693_U9, new_P2_R693_U10,
    new_P2_R693_U11, new_P2_R693_U12, new_P2_R693_U13, new_P2_R693_U14,
    new_P2_R693_U15, new_P2_R693_U16, new_P2_R693_U17, new_P2_R693_U18,
    new_P2_R693_U19, new_P2_R693_U20, new_P2_R693_U21, new_P2_R693_U22,
    new_P2_R693_U23, new_P2_R693_U24, new_P2_R693_U25, new_P2_R693_U26,
    new_P2_R693_U27, new_P2_R693_U28, new_P2_R693_U29, new_P2_R693_U30,
    new_P2_R693_U31, new_P2_R693_U32, new_P2_R693_U33, new_P2_R693_U34,
    new_P2_R693_U35, new_P2_R693_U36, new_P2_R693_U37, new_P2_R693_U38,
    new_P2_R693_U39, new_P2_R693_U40, new_P2_R693_U41, new_P2_R693_U42,
    new_P2_R693_U43, new_P2_R693_U44, new_P2_R693_U45, new_P2_R693_U46,
    new_P2_R693_U47, new_P2_R693_U48, new_P2_R693_U49, new_P2_R693_U50,
    new_P2_R693_U51, new_P2_R693_U52, new_P2_R693_U53, new_P2_R693_U54,
    new_P2_R693_U55, new_P2_R693_U56, new_P2_R693_U57, new_P2_R693_U58,
    new_P2_R693_U59, new_P2_R693_U60, new_P2_R693_U61, new_P2_R693_U62,
    new_P2_R693_U63, new_P2_R693_U64, new_P2_R693_U65, new_P2_R693_U66,
    new_P2_R693_U67, new_P2_R693_U68, new_P2_R693_U69, new_P2_R693_U70,
    new_P2_R693_U71, new_P2_R693_U72, new_P2_R693_U73, new_P2_R693_U74,
    new_P2_R693_U75, new_P2_R693_U76, new_P2_R693_U77, new_P2_R693_U78,
    new_P2_R693_U79, new_P2_R693_U80, new_P2_R693_U81, new_P2_R693_U82,
    new_P2_R693_U83, new_P2_R693_U84, new_P2_R693_U85, new_P2_R693_U86,
    new_P2_R693_U87, new_P2_R693_U88, new_P2_R693_U89, new_P2_R693_U90,
    new_P2_R693_U91, new_P2_R693_U92, new_P2_R693_U93, new_P2_R693_U94,
    new_P2_R693_U95, new_P2_R693_U96, new_P2_R693_U97, new_P2_R693_U98,
    new_P2_R693_U99, new_P2_R693_U100, new_P2_R693_U101, new_P2_R693_U102,
    new_P2_R693_U103, new_P2_R693_U104, new_P2_R693_U105, new_P2_R693_U106,
    new_P2_R693_U107, new_P2_R693_U108, new_P2_R693_U109, new_P2_R693_U110,
    new_P2_R693_U111, new_P2_R693_U112, new_P2_R693_U113, new_P2_R693_U114,
    new_P2_R693_U115, new_P2_R693_U116, new_P2_R693_U117, new_P2_R693_U118,
    new_P2_R693_U119, new_P2_R693_U120, new_P2_R693_U121, new_P2_R693_U122,
    new_P2_R693_U123, new_P2_R693_U124, new_P2_R693_U125, new_P2_R693_U126,
    new_P2_R693_U127, new_P2_R693_U128, new_P2_R693_U129, new_P2_R693_U130,
    new_P2_R693_U131, new_P2_R693_U132, new_P2_R693_U133, new_P2_R693_U134,
    new_P2_R693_U135, new_P2_R693_U136, new_P2_R693_U137, new_P2_R693_U138,
    new_P2_R693_U139, new_P2_R693_U140, new_P2_R693_U141, new_P2_R693_U142,
    new_P2_R693_U143, new_P2_R693_U144, new_P2_R693_U145, new_P2_R693_U146,
    new_P2_R693_U147, new_P2_R693_U148, new_P2_R693_U149, new_P2_R693_U150,
    new_P2_R693_U151, new_P2_R693_U152, new_P2_R693_U153, new_P2_R693_U154,
    new_P2_R693_U155, new_P2_R693_U156, new_P2_R693_U157, new_P2_R693_U158,
    new_P2_R693_U159, new_P2_R693_U160, new_P2_R693_U161, new_P2_R693_U162,
    new_P2_R693_U163, new_P2_R693_U164, new_P2_R693_U165, new_P2_R693_U166,
    new_P2_R693_U167, new_P2_R693_U168, new_P2_R693_U169, new_P2_R693_U170,
    new_P2_R693_U171, new_P2_R693_U172, new_P2_R693_U173, new_P2_R693_U174,
    new_P2_R693_U175, new_P2_R693_U176, new_P2_R693_U177, new_P2_R693_U178,
    new_P2_R693_U179, new_P2_R693_U180, new_P2_R693_U181, new_P2_R693_U182,
    new_P2_R693_U183, new_P2_R693_U184, new_P2_R693_U185, new_P2_R693_U186,
    new_P2_R693_U187, new_P2_R693_U188, new_P2_R693_U189, new_P2_R693_U190,
    new_P2_R693_U191, new_P2_R693_U192, new_P2_R693_U193,
    new_P2_SUB_605_U6, new_P2_SUB_605_U7, new_P2_SUB_605_U8,
    new_P2_SUB_605_U9, new_P2_SUB_605_U10, new_P2_SUB_605_U11,
    new_P2_SUB_605_U12, new_P2_SUB_605_U13, new_P2_SUB_605_U14,
    new_P2_SUB_605_U15, new_P2_SUB_605_U16, new_P2_SUB_605_U17,
    new_P2_SUB_605_U18, new_P2_SUB_605_U19, new_P2_SUB_605_U20,
    new_P2_SUB_605_U21, new_P2_SUB_605_U22, new_P2_SUB_605_U23,
    new_P2_SUB_605_U24, new_P2_SUB_605_U25, new_P2_SUB_605_U26,
    new_P2_SUB_605_U27, new_P2_SUB_605_U28, new_P2_SUB_605_U29,
    new_P2_SUB_605_U30, new_P2_SUB_605_U31, new_P2_SUB_605_U32,
    new_P2_SUB_605_U33, new_P2_SUB_605_U34, new_P2_SUB_605_U35,
    new_P2_SUB_605_U36, new_P2_SUB_605_U37, new_P2_SUB_605_U38,
    new_P2_SUB_605_U39, new_P2_SUB_605_U40, new_P2_SUB_605_U41,
    new_P2_SUB_605_U42, new_P2_SUB_605_U43, new_P2_SUB_605_U44,
    new_P2_SUB_605_U45, new_P2_SUB_605_U46, new_P2_SUB_605_U47,
    new_P2_SUB_605_U48, new_P2_SUB_605_U49, new_P2_SUB_605_U50,
    new_P2_SUB_605_U51, new_P2_SUB_605_U52, new_P2_SUB_605_U53,
    new_P2_SUB_605_U54, new_P2_SUB_605_U55, new_P2_SUB_605_U56,
    new_P2_SUB_605_U57, new_P2_SUB_605_U58, new_P2_SUB_605_U59,
    new_P2_SUB_605_U60, new_P2_SUB_605_U61, new_P2_SUB_605_U62,
    new_P2_SUB_605_U63, new_P2_SUB_605_U64, new_P2_SUB_605_U65,
    new_P2_SUB_605_U66, new_P2_SUB_605_U67, new_P2_SUB_605_U68,
    new_P2_SUB_605_U69, new_P2_SUB_605_U70, new_P2_SUB_605_U71,
    new_P2_SUB_605_U72, new_P2_SUB_605_U73, new_P2_SUB_605_U74,
    new_P2_SUB_605_U75, new_P2_SUB_605_U76, new_P2_SUB_605_U77,
    new_P2_SUB_605_U78, new_P2_SUB_605_U79, new_P2_SUB_605_U80,
    new_P2_SUB_605_U81, new_P2_SUB_605_U82, new_P2_SUB_605_U83,
    new_P2_SUB_605_U84, new_P2_SUB_605_U85, new_P2_SUB_605_U86,
    new_P2_SUB_605_U87, new_P2_SUB_605_U88, new_P2_SUB_605_U89,
    new_P2_SUB_605_U90, new_P2_SUB_605_U91, new_P2_SUB_605_U92,
    new_P2_SUB_605_U93, new_P2_SUB_605_U94, new_P2_SUB_605_U95,
    new_P2_SUB_605_U96, new_P2_SUB_605_U97, new_P2_SUB_605_U98,
    new_P2_SUB_605_U99, new_P2_SUB_605_U100, new_P2_SUB_605_U101,
    new_P2_SUB_605_U102, new_P2_SUB_605_U103, new_P2_SUB_605_U104,
    new_P2_SUB_605_U105, new_P2_SUB_605_U106, new_P2_SUB_605_U107,
    new_P2_SUB_605_U108, new_P2_SUB_605_U109, new_P2_SUB_605_U110,
    new_P2_SUB_605_U111, new_P2_SUB_605_U112, new_P2_SUB_605_U113,
    new_P2_R1095_U6, new_P2_R1095_U7, new_P2_R1095_U8, new_P2_R1095_U9,
    new_P2_R1095_U10, new_P2_R1095_U11, new_P2_R1095_U12, new_P2_R1095_U13,
    new_P2_R1095_U14, new_P2_R1095_U15, new_P2_R1095_U16, new_P2_R1095_U17,
    new_P2_R1095_U18, new_P2_R1095_U19, new_P2_R1095_U20, new_P2_R1095_U21,
    new_P2_R1095_U22, new_P2_R1095_U23, new_P2_R1095_U24, new_P2_R1095_U25,
    new_P2_R1095_U26, new_P2_R1095_U27, new_P2_R1095_U28, new_P2_R1095_U29,
    new_P2_R1095_U30, new_P2_R1095_U31, new_P2_R1095_U32, new_P2_R1095_U33,
    new_P2_R1095_U34, new_P2_R1095_U35, new_P2_R1095_U36, new_P2_R1095_U37,
    new_P2_R1095_U38, new_P2_R1095_U39, new_P2_R1095_U40, new_P2_R1095_U41,
    new_P2_R1095_U42, new_P2_R1095_U43, new_P2_R1095_U44, new_P2_R1095_U45,
    new_P2_R1095_U46, new_P2_R1095_U47, new_P2_R1095_U48, new_P2_R1095_U49,
    new_P2_R1095_U50, new_P2_R1095_U51, new_P2_R1095_U52, new_P2_R1095_U53,
    new_P2_R1095_U54, new_P2_R1095_U55, new_P2_R1095_U56, new_P2_R1095_U57,
    new_P2_R1095_U58, new_P2_R1095_U59, new_P2_R1095_U60, new_P2_R1095_U61,
    new_P2_R1095_U62, new_P2_R1095_U63, new_P2_R1095_U64, new_P2_R1095_U65,
    new_P2_R1095_U66, new_P2_R1095_U67, new_P2_R1095_U68, new_P2_R1095_U69,
    new_P2_R1095_U70, new_P2_R1095_U71, new_P2_R1095_U72, new_P2_R1095_U73,
    new_P2_R1095_U74, new_P2_R1095_U75, new_P2_R1095_U76, new_P2_R1095_U77,
    new_P2_R1095_U78, new_P2_R1095_U79, new_P2_R1095_U80, new_P2_R1095_U81,
    new_P2_R1095_U82, new_P2_R1095_U83, new_P2_R1095_U84, new_P2_R1095_U85,
    new_P2_R1095_U86, new_P2_R1095_U87, new_P2_R1095_U88, new_P2_R1095_U89,
    new_P2_R1095_U90, new_P2_R1095_U91, new_P2_R1095_U92, new_P2_R1095_U93,
    new_P2_R1095_U94, new_P2_R1095_U95, new_P2_R1095_U96, new_P2_R1095_U97,
    new_P2_R1095_U98, new_P2_R1095_U99, new_P2_R1095_U100,
    new_P2_R1095_U101, new_P2_R1095_U102, new_P2_R1095_U103,
    new_P2_R1095_U104, new_P2_R1095_U105, new_P2_R1095_U106,
    new_P2_R1095_U107, new_P2_R1095_U108, new_P2_R1095_U109,
    new_P2_R1095_U110, new_P2_R1095_U111, new_P2_R1095_U112,
    new_P2_R1095_U113, new_P2_R1095_U114, new_P2_R1095_U115,
    new_P2_R1095_U116, new_P2_R1095_U117, new_P2_R1095_U118,
    new_P2_R1095_U119, new_P2_R1095_U120, new_P2_R1095_U121,
    new_P2_R1095_U122, new_P2_R1095_U123, new_P2_R1095_U124,
    new_P2_R1095_U125, new_P2_R1095_U126, new_P2_R1095_U127,
    new_P2_R1095_U128, new_P2_R1095_U129, new_P2_R1095_U130,
    new_P2_R1095_U131, new_P2_R1095_U132, new_P2_R1095_U133,
    new_P2_R1095_U134, new_P2_R1095_U135, new_P2_R1095_U136,
    new_P2_R1095_U137, new_P2_R1095_U138, new_P2_R1095_U139,
    new_P2_R1095_U140, new_P2_R1095_U141, new_P2_R1095_U142,
    new_P2_R1095_U143, new_P2_R1095_U144, new_P2_R1095_U145,
    new_P2_R1095_U146, new_P2_R1095_U147, new_P2_R1095_U148,
    new_P2_R1095_U149, new_P2_R1095_U150, new_P2_R1095_U151,
    new_P2_R1095_U152, new_P2_R1095_U153, new_P2_R1095_U154,
    new_P2_R1095_U155, new_P2_R1095_U156, new_P2_R1095_U157,
    new_P2_R1095_U158, new_P2_R1095_U159, new_P2_R1095_U160,
    new_P2_R1095_U161, new_P2_R1095_U162, new_P2_R1095_U163,
    new_P2_R1095_U164, new_P2_R1095_U165, new_P2_R1095_U166,
    new_P2_R1095_U167, new_P2_R1095_U168, new_P2_R1095_U169,
    new_P2_R1095_U170, new_P2_R1095_U171, new_P2_R1095_U172,
    new_P2_R1095_U173, new_P2_R1095_U174, new_P2_R1095_U175,
    new_P2_R1095_U176, new_P2_R1095_U177, new_P2_R1095_U178,
    new_P2_R1095_U179, new_P2_R1095_U180, new_P2_R1095_U181,
    new_P2_R1095_U182, new_P2_R1095_U183, new_P2_R1095_U184,
    new_P2_R1095_U185, new_P2_R1095_U186, new_P2_R1095_U187,
    new_P2_R1095_U188, new_P2_R1095_U189, new_P2_R1095_U190,
    new_P2_R1095_U191, new_P2_R1095_U192, new_P2_R1095_U193,
    new_P2_R1095_U194, new_P2_R1095_U195, new_P2_R1095_U196,
    new_P2_R1095_U197, new_P2_R1095_U198, new_P2_R1095_U199,
    new_P2_R1095_U200, new_P2_R1095_U201, new_P2_R1095_U202,
    new_P2_R1095_U203, new_P2_R1095_U204, new_P2_R1095_U205,
    new_P2_R1095_U206, new_P2_R1095_U207, new_P2_R1095_U208,
    new_P2_R1095_U209, new_P2_R1095_U210, new_P2_R1095_U211,
    new_P2_R1095_U212, new_P2_R1095_U213, new_P2_R1095_U214,
    new_P2_R1095_U215, new_P2_R1095_U216, new_P2_R1095_U217,
    new_P2_R1095_U218, new_P2_R1095_U219, new_P2_R1095_U220,
    new_P2_R1095_U221, new_P2_R1095_U222, new_P2_R1095_U223,
    new_P2_R1095_U224, new_P2_R1095_U225, new_P2_R1095_U226,
    new_P2_R1095_U227, new_P2_R1095_U228, new_P2_R1095_U229,
    new_P2_R1095_U230, new_P2_R1095_U231, new_P2_R1095_U232,
    new_P2_R1095_U233, new_P2_R1095_U234, new_P2_R1095_U235,
    new_P2_R1095_U236, new_P2_R1095_U237, new_P2_R1095_U238,
    new_P2_R1095_U239, new_P2_R1095_U240, new_P2_R1095_U241,
    new_P2_R1095_U242, new_P2_R1095_U243, new_P2_R1095_U244,
    new_P2_R1095_U245, new_P2_R1095_U246, new_P2_R1095_U247,
    new_P2_R1095_U248, new_P2_R1095_U249, new_P2_R1095_U250,
    new_P2_R1095_U251, new_P2_R1095_U252, new_P2_R1095_U253,
    new_P2_R1095_U254, new_P2_R1095_U255, new_P2_R1095_U256,
    new_P2_R1095_U257, new_P2_R1095_U258, new_P2_R1095_U259,
    new_P2_R1095_U260, new_P2_R1095_U261, new_P2_R1095_U262,
    new_P2_R1095_U263, new_P2_R1095_U264, new_P2_R1095_U265,
    new_P2_R1095_U266, new_P2_R1095_U267, new_P2_R1095_U268,
    new_P2_R1095_U269, new_P2_R1095_U270, new_P2_R1095_U271,
    new_P2_R1095_U272, new_P2_R1095_U273, new_P2_R1095_U274,
    new_P2_R1095_U275, new_P2_R1095_U276, new_P2_R1095_U277,
    new_P2_R1095_U278, new_P2_R1095_U279, new_P2_R1095_U280,
    new_P2_R1095_U281, new_P2_R1095_U282, new_P2_R1095_U283,
    new_P2_R1095_U284, new_P2_R1095_U285, new_P2_R1095_U286,
    new_P2_R1095_U287, new_P2_R1095_U288, new_P2_R1095_U289,
    new_P2_R1095_U290, new_P2_R1095_U291, new_P2_R1095_U292,
    new_P2_R1095_U293, new_P2_R1095_U294, new_P2_R1095_U295,
    new_P2_R1095_U296, new_P2_R1095_U297, new_P2_R1095_U298,
    new_P2_R1095_U299, new_P2_R1095_U300, new_P2_R1095_U301,
    new_P2_R1095_U302, new_P2_R1095_U303, new_P2_R1095_U304,
    new_P2_R1095_U305, new_P2_R1095_U306, new_P2_R1095_U307,
    new_P2_R1095_U308, new_P2_R1095_U309, new_P2_R1095_U310,
    new_P2_R1095_U311, new_P2_R1095_U312, new_P2_R1095_U313,
    new_P2_R1095_U314, new_P2_R1095_U315, new_P2_R1095_U316,
    new_P2_R1095_U317, new_P2_R1095_U318, new_P2_R1095_U319,
    new_P2_R1095_U320, new_P2_R1095_U321, new_P2_R1095_U322,
    new_P2_R1095_U323, new_P2_R1095_U324, new_P2_R1095_U325,
    new_P2_R1095_U326, new_P2_R1095_U327, new_P2_R1095_U328,
    new_P2_R1095_U329, new_P2_R1095_U330, new_P2_R1095_U331,
    new_P2_R1095_U332, new_P2_R1095_U333, new_P2_R1095_U334,
    new_P2_R1095_U335, new_P2_R1095_U336, new_P2_R1095_U337,
    new_P2_R1095_U338, new_P2_R1095_U339, new_P2_R1095_U340,
    new_P2_R1095_U341, new_P2_R1095_U342, new_P2_R1095_U343,
    new_P2_R1095_U344, new_P2_R1095_U345, new_P2_R1095_U346,
    new_P2_R1095_U347, new_P2_R1095_U348, new_P2_R1095_U349,
    new_P2_R1095_U350, new_P2_R1095_U351, new_P2_R1095_U352,
    new_P2_R1095_U353, new_P2_R1095_U354, new_P2_R1095_U355,
    new_P2_R1095_U356, new_P2_R1095_U357, new_P2_R1095_U358,
    new_P2_R1095_U359, new_P2_R1095_U360, new_P2_R1095_U361,
    new_P2_R1095_U362, new_P2_R1095_U363, new_P2_R1095_U364,
    new_P2_R1095_U365, new_P2_R1095_U366, new_P2_R1095_U367,
    new_P2_R1095_U368, new_P2_R1095_U369, new_P2_R1095_U370,
    new_P2_R1095_U371, new_P2_R1095_U372, new_P2_R1095_U373,
    new_P2_R1095_U374, new_P2_R1095_U375, new_P2_R1095_U376,
    new_P2_R1095_U377, new_P2_R1095_U378, new_P2_R1095_U379,
    new_P2_R1095_U380, new_P2_R1095_U381, new_P2_R1095_U382,
    new_P2_R1095_U383, new_P2_R1095_U384, new_P2_R1095_U385,
    new_P2_R1095_U386, new_P2_R1095_U387, new_P2_R1095_U388,
    new_P2_R1095_U389, new_P2_R1095_U390, new_P2_R1095_U391,
    new_P2_R1095_U392, new_P2_R1095_U393, new_P2_R1095_U394,
    new_P2_R1095_U395, new_P2_R1095_U396, new_P2_R1095_U397,
    new_P2_R1095_U398, new_P2_R1095_U399, new_P2_R1095_U400,
    new_P2_R1095_U401, new_P2_R1095_U402, new_P2_R1095_U403,
    new_P2_R1095_U404, new_P2_R1095_U405, new_P2_R1095_U406,
    new_P2_R1095_U407, new_P2_R1095_U408, new_P2_R1095_U409,
    new_P2_R1095_U410, new_P2_R1095_U411, new_P2_R1095_U412,
    new_P2_R1095_U413, new_P2_R1095_U414, new_P2_R1095_U415,
    new_P2_R1095_U416, new_P2_R1095_U417, new_P2_R1095_U418,
    new_P2_R1095_U419, new_P2_R1095_U420, new_P2_R1095_U421,
    new_P2_R1095_U422, new_P2_R1095_U423, new_P2_R1095_U424,
    new_P2_R1095_U425, new_P2_R1095_U426, new_P2_R1095_U427,
    new_P2_R1095_U428, new_P2_R1095_U429, new_P2_R1095_U430,
    new_P2_R1095_U431, new_P2_R1095_U432, new_P2_R1095_U433,
    new_P2_R1095_U434, new_P2_R1095_U435, new_P2_R1095_U436,
    new_P2_R1095_U437, new_P2_R1095_U438, new_P2_R1095_U439,
    new_P2_R1095_U440, new_P2_R1095_U441, new_P2_R1095_U442,
    new_P2_R1095_U443, new_P2_R1095_U444, new_P2_R1095_U445,
    new_P2_R1095_U446, new_P2_R1095_U447, new_P2_R1095_U448,
    new_P2_R1095_U449, new_P2_R1095_U450, new_P2_R1095_U451,
    new_P2_R1095_U452, new_P2_R1095_U453, new_P2_R1095_U454,
    new_P2_R1095_U455, new_P2_R1095_U456, new_P2_R1095_U457,
    new_P2_R1095_U458, new_P2_R1095_U459, new_P2_R1095_U460,
    new_P2_R1095_U461, new_P2_R1095_U462, new_P2_R1095_U463,
    new_P2_R1095_U464, new_P2_R1095_U465, new_P2_R1095_U466,
    new_P2_R1095_U467, new_P2_R1095_U468, new_P2_R1095_U469,
    new_P2_R1095_U470, new_P2_R1095_U471, new_P2_R1095_U472,
    new_P2_R1095_U473, new_P2_R1095_U474, new_P2_R1095_U475,
    new_P2_R1095_U476, new_P2_R1095_U477, new_P2_R1095_U478,
    new_P2_R1095_U479, new_P2_R1095_U480, new_P2_R1095_U481,
    new_P2_R1095_U482, new_P2_R1095_U483, new_P2_R1095_U484,
    new_P2_R1095_U485, new_P2_R1095_U486, new_P2_R1095_U487,
    new_P2_R1095_U488, new_P2_R1095_U489, new_P2_R1212_U6, new_P2_R1212_U7,
    new_P2_R1212_U8, new_P2_R1212_U9, new_P2_R1212_U10, new_P2_R1212_U11,
    new_P2_R1212_U12, new_P2_R1212_U13, new_P2_R1212_U14, new_P2_R1212_U15,
    new_P2_R1212_U16, new_P2_R1212_U17, new_P2_R1212_U18, new_P2_R1212_U19,
    new_P2_R1212_U20, new_P2_R1212_U21, new_P2_R1212_U22, new_P2_R1212_U23,
    new_P2_R1212_U24, new_P2_R1212_U25, new_P2_R1212_U26, new_P2_R1212_U27,
    new_P2_R1212_U28, new_P2_R1212_U29, new_P2_R1212_U30, new_P2_R1212_U31,
    new_P2_R1212_U32, new_P2_R1212_U33, new_P2_R1212_U34, new_P2_R1212_U35,
    new_P2_R1212_U36, new_P2_R1212_U37, new_P2_R1212_U38, new_P2_R1212_U39,
    new_P2_R1212_U40, new_P2_R1212_U41, new_P2_R1212_U42, new_P2_R1212_U43,
    new_P2_R1212_U44, new_P2_R1212_U45, new_P2_R1212_U46, new_P2_R1212_U47,
    new_P2_R1212_U48, new_P2_R1212_U49, new_P2_R1212_U50, new_P2_R1212_U51,
    new_P2_R1212_U52, new_P2_R1212_U53, new_P2_R1212_U54, new_P2_R1212_U55,
    new_P2_R1212_U56, new_P2_R1212_U57, new_P2_R1212_U58, new_P2_R1212_U59,
    new_P2_R1212_U60, new_P2_R1212_U61, new_P2_R1212_U62, new_P2_R1212_U63,
    new_P2_R1212_U64, new_P2_R1212_U65, new_P2_R1212_U66, new_P2_R1212_U67,
    new_P2_R1212_U68, new_P2_R1212_U69, new_P2_R1212_U70, new_P2_R1212_U71,
    new_P2_R1212_U72, new_P2_R1212_U73, new_P2_R1212_U74, new_P2_R1212_U75,
    new_P2_R1212_U76, new_P2_R1212_U77, new_P2_R1212_U78, new_P2_R1212_U79,
    new_P2_R1212_U80, new_P2_R1212_U81, new_P2_R1212_U82, new_P2_R1212_U83,
    new_P2_R1212_U84, new_P2_R1212_U85, new_P2_R1212_U86, new_P2_R1212_U87,
    new_P2_R1212_U88, new_P2_R1212_U89, new_P2_R1212_U90, new_P2_R1212_U91,
    new_P2_R1212_U92, new_P2_R1212_U93, new_P2_R1212_U94, new_P2_R1212_U95,
    new_P2_R1212_U96, new_P2_R1212_U97, new_P2_R1212_U98, new_P2_R1212_U99,
    new_P2_R1212_U100, new_P2_R1212_U101, new_P2_R1212_U102,
    new_P2_R1212_U103, new_P2_R1212_U104, new_P2_R1212_U105,
    new_P2_R1212_U106, new_P2_R1212_U107, new_P2_R1212_U108,
    new_P2_R1212_U109, new_P2_R1212_U110, new_P2_R1212_U111,
    new_P2_R1212_U112, new_P2_R1212_U113, new_P2_R1212_U114,
    new_P2_R1212_U115, new_P2_R1212_U116, new_P2_R1212_U117,
    new_P2_R1212_U118, new_P2_R1212_U119, new_P2_R1212_U120,
    new_P2_R1212_U121, new_P2_R1212_U122, new_P2_R1212_U123,
    new_P2_R1212_U124, new_P2_R1212_U125, new_P2_R1212_U126,
    new_P2_R1212_U127, new_P2_R1212_U128, new_P2_R1212_U129,
    new_P2_R1212_U130, new_P2_R1212_U131, new_P2_R1212_U132,
    new_P2_R1212_U133, new_P2_R1212_U134, new_P2_R1212_U135,
    new_P2_R1212_U136, new_P2_R1212_U137, new_P2_R1212_U138,
    new_P2_R1212_U139, new_P2_R1212_U140, new_P2_R1212_U141,
    new_P2_R1212_U142, new_P2_R1212_U143, new_P2_R1212_U144,
    new_P2_R1212_U145, new_P2_R1212_U146, new_P2_R1212_U147,
    new_P2_R1212_U148, new_P2_R1212_U149, new_P2_R1212_U150,
    new_P2_R1212_U151, new_P2_R1212_U152, new_P2_R1212_U153,
    new_P2_R1212_U154, new_P2_R1212_U155, new_P2_R1212_U156,
    new_P2_R1212_U157, new_P2_R1212_U158, new_P2_R1212_U159,
    new_P2_R1212_U160, new_P2_R1212_U161, new_P2_R1212_U162,
    new_P2_R1212_U163, new_P2_R1212_U164, new_P2_R1212_U165,
    new_P2_R1212_U166, new_P2_R1212_U167, new_P2_R1212_U168,
    new_P2_R1212_U169, new_P2_R1212_U170, new_P2_R1212_U171,
    new_P2_R1212_U172, new_P2_R1212_U173, new_P2_R1212_U174,
    new_P2_R1212_U175, new_P2_R1212_U176, new_P2_R1212_U177,
    new_P2_R1212_U178, new_P2_R1212_U179, new_P2_R1212_U180,
    new_P2_R1212_U181, new_P2_R1212_U182, new_P2_R1212_U183,
    new_P2_R1212_U184, new_P2_R1212_U185, new_P2_R1212_U186,
    new_P2_R1212_U187, new_P2_R1212_U188, new_P2_R1212_U189,
    new_P2_R1212_U190, new_P2_R1212_U191, new_P2_R1212_U192,
    new_P2_R1212_U193, new_P2_R1212_U194, new_P2_R1212_U195,
    new_P2_R1212_U196, new_P2_R1212_U197, new_P2_R1212_U198,
    new_P2_R1212_U199, new_P2_R1212_U200, new_P2_R1212_U201,
    new_P2_R1212_U202, new_P2_R1212_U203, new_P2_R1212_U204,
    new_P2_R1212_U205, new_P2_R1212_U206, new_P2_R1212_U207,
    new_P2_R1212_U208, new_P2_R1212_U209, new_P2_R1212_U210,
    new_P2_R1212_U211, new_P2_R1212_U212, new_P2_R1212_U213,
    new_P2_R1212_U214, new_P2_R1212_U215, new_P2_R1212_U216,
    new_P2_R1212_U217, new_P2_R1212_U218, new_P2_R1212_U219,
    new_P2_R1212_U220, new_P2_R1212_U221, new_P2_R1212_U222,
    new_P2_R1212_U223, new_P2_R1212_U224, new_P2_R1212_U225,
    new_P2_R1212_U226, new_P2_R1212_U227, new_P2_R1212_U228,
    new_P2_R1212_U229, new_P2_R1212_U230, new_P2_R1212_U231,
    new_P2_R1212_U232, new_P2_R1212_U233, new_P2_R1212_U234,
    new_P2_R1212_U235, new_P2_R1212_U236, new_P2_R1212_U237,
    new_P2_R1212_U238, new_P2_R1212_U239, new_P2_R1212_U240,
    new_P2_R1212_U241, new_P2_R1212_U242, new_P2_R1212_U243,
    new_P2_R1212_U244, new_P2_R1212_U245, new_P2_R1212_U246,
    new_P2_R1212_U247, new_P2_R1212_U248, new_P2_R1212_U249,
    new_P2_R1212_U250, new_P2_R1212_U251, new_P2_R1212_U252,
    new_P2_R1212_U253, new_P2_R1212_U254, new_P2_R1212_U255,
    new_P2_R1212_U256, new_P2_R1212_U257, new_P2_R1212_U258,
    new_P2_R1212_U259, new_P2_R1212_U260, new_P2_R1212_U261,
    new_P2_R1212_U262, new_P2_R1212_U263, new_P2_R1212_U264,
    new_P2_R1212_U265, new_P2_R1212_U266, new_P2_R1212_U267,
    new_P2_R1212_U268, new_P2_R1212_U269, new_P2_R1212_U270,
    new_P2_R1212_U271, new_P2_R1212_U272, new_P2_R1212_U273,
    new_P2_R1212_U274, new_P2_R1212_U275, new_P2_R1212_U276,
    new_P2_R1209_U6, new_P2_R1209_U7, new_P2_R1209_U8, new_P2_R1209_U9,
    new_P2_R1209_U10, new_P2_R1209_U11, new_P2_R1209_U12, new_P2_R1209_U13,
    new_P2_R1209_U14, new_P2_R1209_U15, new_P2_R1209_U16, new_P2_R1209_U17,
    new_P2_R1209_U18, new_P2_R1209_U19, new_P2_R1209_U20, new_P2_R1209_U21,
    new_P2_R1209_U22, new_P2_R1209_U23, new_P2_R1209_U24, new_P2_R1209_U25,
    new_P2_R1209_U26, new_P2_R1209_U27, new_P2_R1209_U28, new_P2_R1209_U29,
    new_P2_R1209_U30, new_P2_R1209_U31, new_P2_R1209_U32, new_P2_R1209_U33,
    new_P2_R1209_U34, new_P2_R1209_U35, new_P2_R1209_U36, new_P2_R1209_U37,
    new_P2_R1209_U38, new_P2_R1209_U39, new_P2_R1209_U40, new_P2_R1209_U41,
    new_P2_R1209_U42, new_P2_R1209_U43, new_P2_R1209_U44, new_P2_R1209_U45,
    new_P2_R1209_U46, new_P2_R1209_U47, new_P2_R1209_U48, new_P2_R1209_U49,
    new_P2_R1209_U50, new_P2_R1209_U51, new_P2_R1209_U52, new_P2_R1209_U53,
    new_P2_R1209_U54, new_P2_R1209_U55, new_P2_R1209_U56, new_P2_R1209_U57,
    new_P2_R1209_U58, new_P2_R1209_U59, new_P2_R1209_U60, new_P2_R1209_U61,
    new_P2_R1209_U62, new_P2_R1209_U63, new_P2_R1209_U64, new_P2_R1209_U65,
    new_P2_R1209_U66, new_P2_R1209_U67, new_P2_R1209_U68, new_P2_R1209_U69,
    new_P2_R1209_U70, new_P2_R1209_U71, new_P2_R1209_U72, new_P2_R1209_U73,
    new_P2_R1209_U74, new_P2_R1209_U75, new_P2_R1209_U76, new_P2_R1209_U77,
    new_P2_R1209_U78, new_P2_R1209_U79, new_P2_R1209_U80, new_P2_R1209_U81,
    new_P2_R1209_U82, new_P2_R1209_U83, new_P2_R1209_U84, new_P2_R1209_U85,
    new_P2_R1209_U86, new_P2_R1209_U87, new_P2_R1209_U88, new_P2_R1209_U89,
    new_P2_R1209_U90, new_P2_R1209_U91, new_P2_R1209_U92, new_P2_R1209_U93,
    new_P2_R1209_U94, new_P2_R1209_U95, new_P2_R1209_U96, new_P2_R1209_U97,
    new_P2_R1209_U98, new_P2_R1209_U99, new_P2_R1209_U100,
    new_P2_R1209_U101, new_P2_R1209_U102, new_P2_R1209_U103,
    new_P2_R1209_U104, new_P2_R1209_U105, new_P2_R1209_U106,
    new_P2_R1209_U107, new_P2_R1209_U108, new_P2_R1209_U109,
    new_P2_R1209_U110, new_P2_R1209_U111, new_P2_R1209_U112,
    new_P2_R1209_U113, new_P2_R1209_U114, new_P2_R1209_U115,
    new_P2_R1209_U116, new_P2_R1209_U117, new_P2_R1209_U118,
    new_P2_R1209_U119, new_P2_R1209_U120, new_P2_R1209_U121,
    new_P2_R1209_U122, new_P2_R1209_U123, new_P2_R1209_U124,
    new_P2_R1209_U125, new_P2_R1209_U126, new_P2_R1209_U127,
    new_P2_R1209_U128, new_P2_R1209_U129, new_P2_R1209_U130,
    new_P2_R1209_U131, new_P2_R1209_U132, new_P2_R1209_U133,
    new_P2_R1209_U134, new_P2_R1209_U135, new_P2_R1209_U136,
    new_P2_R1209_U137, new_P2_R1209_U138, new_P2_R1209_U139,
    new_P2_R1209_U140, new_P2_R1209_U141, new_P2_R1209_U142,
    new_P2_R1209_U143, new_P2_R1209_U144, new_P2_R1209_U145,
    new_P2_R1209_U146, new_P2_R1209_U147, new_P2_R1209_U148,
    new_P2_R1209_U149, new_P2_R1209_U150, new_P2_R1209_U151,
    new_P2_R1209_U152, new_P2_R1209_U153, new_P2_R1209_U154,
    new_P2_R1209_U155, new_P2_R1209_U156, new_P2_R1209_U157,
    new_P2_R1209_U158, new_P2_R1209_U159, new_P2_R1209_U160,
    new_P2_R1209_U161, new_P2_R1209_U162, new_P2_R1209_U163,
    new_P2_R1209_U164, new_P2_R1209_U165, new_P2_R1209_U166,
    new_P2_R1209_U167, new_P2_R1209_U168, new_P2_R1209_U169,
    new_P2_R1209_U170, new_P2_R1209_U171, new_P2_R1209_U172,
    new_P2_R1209_U173, new_P2_R1209_U174, new_P2_R1209_U175,
    new_P2_R1209_U176, new_P2_R1209_U177, new_P2_R1209_U178,
    new_P2_R1209_U179, new_P2_R1209_U180, new_P2_R1209_U181,
    new_P2_R1209_U182, new_P2_R1209_U183, new_P2_R1209_U184,
    new_P2_R1209_U185, new_P2_R1209_U186, new_P2_R1209_U187,
    new_P2_R1209_U188, new_P2_R1209_U189, new_P2_R1209_U190,
    new_P2_R1209_U191, new_P2_R1209_U192, new_P2_R1209_U193,
    new_P2_R1209_U194, new_P2_R1209_U195, new_P2_R1209_U196,
    new_P2_R1209_U197, new_P2_R1209_U198, new_P2_R1209_U199,
    new_P2_R1209_U200, new_P2_R1209_U201, new_P2_R1209_U202,
    new_P2_R1209_U203, new_P2_R1209_U204, new_P2_R1209_U205,
    new_P2_R1209_U206, new_P2_R1209_U207, new_P2_R1209_U208,
    new_P2_R1209_U209, new_P2_R1209_U210, new_P2_R1209_U211,
    new_P2_R1209_U212, new_P2_R1209_U213, new_P2_R1209_U214,
    new_P2_R1209_U215, new_P2_R1209_U216, new_P2_R1209_U217,
    new_P2_R1209_U218, new_P2_R1209_U219, new_P2_R1209_U220,
    new_P2_R1209_U221, new_P2_R1209_U222, new_P2_R1209_U223,
    new_P2_R1209_U224, new_P2_R1209_U225, new_P2_R1209_U226,
    new_P2_R1209_U227, new_P2_R1209_U228, new_P2_R1209_U229,
    new_P2_R1209_U230, new_P2_R1209_U231, new_P2_R1209_U232,
    new_P2_R1209_U233, new_P2_R1209_U234, new_P2_R1209_U235,
    new_P2_R1209_U236, new_P2_R1209_U237, new_P2_R1209_U238,
    new_P2_R1209_U239, new_P2_R1209_U240, new_P2_R1209_U241,
    new_P2_R1209_U242, new_P2_R1209_U243, new_P2_R1209_U244,
    new_P2_R1209_U245, new_P2_R1209_U246, new_P2_R1209_U247,
    new_P2_R1209_U248, new_P2_R1209_U249, new_P2_R1209_U250,
    new_P2_R1209_U251, new_P2_R1209_U252, new_P2_R1209_U253,
    new_P2_R1209_U254, new_P2_R1209_U255, new_P2_R1209_U256,
    new_P2_R1209_U257, new_P2_R1209_U258, new_P2_R1209_U259,
    new_P2_R1209_U260, new_P2_R1209_U261, new_P2_R1209_U262,
    new_P2_R1209_U263, new_P2_R1209_U264, new_P2_R1209_U265,
    new_P2_R1209_U266, new_P2_R1209_U267, new_P2_R1209_U268,
    new_P2_R1209_U269, new_P2_R1209_U270, new_P2_R1209_U271,
    new_P2_R1209_U272, new_P2_R1209_U273, new_P2_R1209_U274,
    new_P2_R1209_U275, new_P2_R1209_U276, new_P2_R1300_U6, new_P2_R1300_U7,
    new_P2_R1300_U8, new_P2_R1300_U9, new_P2_R1300_U10, new_P2_R1200_U6,
    new_P2_R1200_U7, new_P2_R1200_U8, new_P2_R1200_U9, new_P2_R1200_U10,
    new_P2_R1200_U11, new_P2_R1200_U12, new_P2_R1200_U13, new_P2_R1200_U14,
    new_P2_R1200_U15, new_P2_R1200_U16, new_P2_R1200_U17, new_P2_R1200_U18,
    new_P2_R1200_U19, new_P2_R1200_U20, new_P2_R1200_U21, new_P2_R1200_U22,
    new_P2_R1200_U23, new_P2_R1200_U24, new_P2_R1200_U25, new_P2_R1200_U26,
    new_P2_R1200_U27, new_P2_R1200_U28, new_P2_R1200_U29, new_P2_R1200_U30,
    new_P2_R1200_U31, new_P2_R1200_U32, new_P2_R1200_U33, new_P2_R1200_U34,
    new_P2_R1200_U35, new_P2_R1200_U36, new_P2_R1200_U37, new_P2_R1200_U38,
    new_P2_R1200_U39, new_P2_R1200_U40, new_P2_R1200_U41, new_P2_R1200_U42,
    new_P2_R1200_U43, new_P2_R1200_U44, new_P2_R1200_U45, new_P2_R1200_U46,
    new_P2_R1200_U47, new_P2_R1200_U48, new_P2_R1200_U49, new_P2_R1200_U50,
    new_P2_R1200_U51, new_P2_R1200_U52, new_P2_R1200_U53, new_P2_R1200_U54,
    new_P2_R1200_U55, new_P2_R1200_U56, new_P2_R1200_U57, new_P2_R1200_U58,
    new_P2_R1200_U59, new_P2_R1200_U60, new_P2_R1200_U61, new_P2_R1200_U62,
    new_P2_R1200_U63, new_P2_R1200_U64, new_P2_R1200_U65, new_P2_R1200_U66,
    new_P2_R1200_U67, new_P2_R1200_U68, new_P2_R1200_U69, new_P2_R1200_U70,
    new_P2_R1200_U71, new_P2_R1200_U72, new_P2_R1200_U73, new_P2_R1200_U74,
    new_P2_R1200_U75, new_P2_R1200_U76, new_P2_R1200_U77, new_P2_R1200_U78,
    new_P2_R1200_U79, new_P2_R1200_U80, new_P2_R1200_U81, new_P2_R1200_U82,
    new_P2_R1200_U83, new_P2_R1200_U84, new_P2_R1200_U85, new_P2_R1200_U86,
    new_P2_R1200_U87, new_P2_R1200_U88, new_P2_R1200_U89, new_P2_R1200_U90,
    new_P2_R1200_U91, new_P2_R1200_U92, new_P2_R1200_U93, new_P2_R1200_U94,
    new_P2_R1200_U95, new_P2_R1200_U96, new_P2_R1200_U97, new_P2_R1200_U98,
    new_P2_R1200_U99, new_P2_R1200_U100, new_P2_R1200_U101,
    new_P2_R1200_U102, new_P2_R1200_U103, new_P2_R1200_U104,
    new_P2_R1200_U105, new_P2_R1200_U106, new_P2_R1200_U107,
    new_P2_R1200_U108, new_P2_R1200_U109, new_P2_R1200_U110,
    new_P2_R1200_U111, new_P2_R1200_U112, new_P2_R1200_U113,
    new_P2_R1200_U114, new_P2_R1200_U115, new_P2_R1200_U116,
    new_P2_R1200_U117, new_P2_R1200_U118, new_P2_R1200_U119,
    new_P2_R1200_U120, new_P2_R1200_U121, new_P2_R1200_U122,
    new_P2_R1200_U123, new_P2_R1200_U124, new_P2_R1200_U125,
    new_P2_R1200_U126, new_P2_R1200_U127, new_P2_R1200_U128,
    new_P2_R1200_U129, new_P2_R1200_U130, new_P2_R1200_U131,
    new_P2_R1200_U132, new_P2_R1200_U133, new_P2_R1200_U134,
    new_P2_R1200_U135, new_P2_R1200_U136, new_P2_R1200_U137,
    new_P2_R1200_U138, new_P2_R1200_U139, new_P2_R1200_U140,
    new_P2_R1200_U141, new_P2_R1200_U142, new_P2_R1200_U143,
    new_P2_R1200_U144, new_P2_R1200_U145, new_P2_R1200_U146,
    new_P2_R1200_U147, new_P2_R1200_U148, new_P2_R1200_U149,
    new_P2_R1200_U150, new_P2_R1200_U151, new_P2_R1200_U152,
    new_P2_R1200_U153, new_P2_R1200_U154, new_P2_R1200_U155,
    new_P2_R1200_U156, new_P2_R1200_U157, new_P2_R1200_U158,
    new_P2_R1200_U159, new_P2_R1200_U160, new_P2_R1200_U161,
    new_P2_R1200_U162, new_P2_R1200_U163, new_P2_R1200_U164,
    new_P2_R1200_U165, new_P2_R1200_U166, new_P2_R1200_U167,
    new_P2_R1200_U168, new_P2_R1200_U169, new_P2_R1200_U170,
    new_P2_R1200_U171, new_P2_R1200_U172, new_P2_R1200_U173,
    new_P2_R1200_U174, new_P2_R1200_U175, new_P2_R1200_U176,
    new_P2_R1200_U177, new_P2_R1200_U178, new_P2_R1200_U179,
    new_P2_R1200_U180, new_P2_R1200_U181, new_P2_R1200_U182,
    new_P2_R1200_U183, new_P2_R1200_U184, new_P2_R1200_U185,
    new_P2_R1200_U186, new_P2_R1200_U187, new_P2_R1200_U188,
    new_P2_R1200_U189, new_P2_R1200_U190, new_P2_R1200_U191,
    new_P2_R1200_U192, new_P2_R1200_U193, new_P2_R1200_U194,
    new_P2_R1200_U195, new_P2_R1200_U196, new_P2_R1200_U197,
    new_P2_R1200_U198, new_P2_R1200_U199, new_P2_R1200_U200,
    new_P2_R1200_U201, new_P2_R1200_U202, new_P2_R1200_U203,
    new_P2_R1200_U204, new_P2_R1200_U205, new_P2_R1200_U206,
    new_P2_R1200_U207, new_P2_R1200_U208, new_P2_R1200_U209,
    new_P2_R1200_U210, new_P2_R1200_U211, new_P2_R1200_U212,
    new_P2_R1200_U213, new_P2_R1200_U214, new_P2_R1200_U215,
    new_P2_R1200_U216, new_P2_R1200_U217, new_P2_R1200_U218,
    new_P2_R1200_U219, new_P2_R1200_U220, new_P2_R1200_U221,
    new_P2_R1200_U222, new_P2_R1200_U223, new_P2_R1200_U224,
    new_P2_R1200_U225, new_P2_R1200_U226, new_P2_R1200_U227,
    new_P2_R1200_U228, new_P2_R1200_U229, new_P2_R1200_U230,
    new_P2_R1200_U231, new_P2_R1200_U232, new_P2_R1200_U233,
    new_P2_R1200_U234, new_P2_R1200_U235, new_P2_R1200_U236,
    new_P2_R1200_U237, new_P2_R1200_U238, new_P2_R1200_U239,
    new_P2_R1200_U240, new_P2_R1200_U241, new_P2_R1200_U242,
    new_P2_R1200_U243, new_P2_R1200_U244, new_P2_R1200_U245,
    new_P2_R1200_U246, new_P2_R1200_U247, new_P2_R1200_U248,
    new_P2_R1200_U249, new_P2_R1200_U250, new_P2_R1200_U251,
    new_P2_R1200_U252, new_P2_R1200_U253, new_P2_R1200_U254,
    new_P2_R1200_U255, new_P2_R1200_U256, new_P2_R1200_U257,
    new_P2_R1200_U258, new_P2_R1200_U259, new_P2_R1200_U260,
    new_P2_R1200_U261, new_P2_R1200_U262, new_P2_R1200_U263,
    new_P2_R1200_U264, new_P2_R1200_U265, new_P2_R1200_U266,
    new_P2_R1200_U267, new_P2_R1200_U268, new_P2_R1200_U269,
    new_P2_R1200_U270, new_P2_R1200_U271, new_P2_R1200_U272,
    new_P2_R1200_U273, new_P2_R1200_U274, new_P2_R1200_U275,
    new_P2_R1200_U276, new_P2_R1200_U277, new_P2_R1200_U278,
    new_P2_R1200_U279, new_P2_R1200_U280, new_P2_R1200_U281,
    new_P2_R1200_U282, new_P2_R1200_U283, new_P2_R1200_U284,
    new_P2_R1200_U285, new_P2_R1200_U286, new_P2_R1200_U287,
    new_P2_R1200_U288, new_P2_R1200_U289, new_P2_R1200_U290,
    new_P2_R1200_U291, new_P2_R1200_U292, new_P2_R1200_U293,
    new_P2_R1200_U294, new_P2_R1200_U295, new_P2_R1200_U296,
    new_P2_R1200_U297, new_P2_R1200_U298, new_P2_R1200_U299,
    new_P2_R1200_U300, new_P2_R1200_U301, new_P2_R1200_U302,
    new_P2_R1200_U303, new_P2_R1200_U304, new_P2_R1200_U305,
    new_P2_R1200_U306, new_P2_R1200_U307, new_P2_R1200_U308,
    new_P2_R1200_U309, new_P2_R1200_U310, new_P2_R1200_U311,
    new_P2_R1200_U312, new_P2_R1200_U313, new_P2_R1200_U314,
    new_P2_R1200_U315, new_P2_R1200_U316, new_P2_R1200_U317,
    new_P2_R1200_U318, new_P2_R1200_U319, new_P2_R1200_U320,
    new_P2_R1200_U321, new_P2_R1200_U322, new_P2_R1200_U323,
    new_P2_R1200_U324, new_P2_R1200_U325, new_P2_R1200_U326,
    new_P2_R1200_U327, new_P2_R1200_U328, new_P2_R1200_U329,
    new_P2_R1200_U330, new_P2_R1200_U331, new_P2_R1200_U332,
    new_P2_R1200_U333, new_P2_R1200_U334, new_P2_R1200_U335,
    new_P2_R1200_U336, new_P2_R1200_U337, new_P2_R1200_U338,
    new_P2_R1200_U339, new_P2_R1200_U340, new_P2_R1200_U341,
    new_P2_R1200_U342, new_P2_R1200_U343, new_P2_R1200_U344,
    new_P2_R1200_U345, new_P2_R1200_U346, new_P2_R1200_U347,
    new_P2_R1200_U348, new_P2_R1200_U349, new_P2_R1200_U350,
    new_P2_R1200_U351, new_P2_R1200_U352, new_P2_R1200_U353,
    new_P2_R1200_U354, new_P2_R1200_U355, new_P2_R1200_U356,
    new_P2_R1200_U357, new_P2_R1200_U358, new_P2_R1200_U359,
    new_P2_R1200_U360, new_P2_R1200_U361, new_P2_R1200_U362,
    new_P2_R1200_U363, new_P2_R1200_U364, new_P2_R1200_U365,
    new_P2_R1200_U366, new_P2_R1200_U367, new_P2_R1200_U368,
    new_P2_R1200_U369, new_P2_R1200_U370, new_P2_R1200_U371,
    new_P2_R1200_U372, new_P2_R1200_U373, new_P2_R1200_U374,
    new_P2_R1200_U375, new_P2_R1200_U376, new_P2_R1200_U377,
    new_P2_R1200_U378, new_P2_R1200_U379, new_P2_R1200_U380,
    new_P2_R1200_U381, new_P2_R1200_U382, new_P2_R1200_U383,
    new_P2_R1200_U384, new_P2_R1200_U385, new_P2_R1200_U386,
    new_P2_R1200_U387, new_P2_R1200_U388, new_P2_R1200_U389,
    new_P2_R1200_U390, new_P2_R1200_U391, new_P2_R1200_U392,
    new_P2_R1200_U393, new_P2_R1200_U394, new_P2_R1200_U395,
    new_P2_R1200_U396, new_P2_R1200_U397, new_P2_R1200_U398,
    new_P2_R1200_U399, new_P2_R1200_U400, new_P2_R1200_U401,
    new_P2_R1200_U402, new_P2_R1200_U403, new_P2_R1200_U404,
    new_P2_R1200_U405, new_P2_R1200_U406, new_P2_R1200_U407,
    new_P2_R1200_U408, new_P2_R1200_U409, new_P2_R1200_U410,
    new_P2_R1200_U411, new_P2_R1200_U412, new_P2_R1200_U413,
    new_P2_R1200_U414, new_P2_R1200_U415, new_P2_R1200_U416,
    new_P2_R1200_U417, new_P2_R1200_U418, new_P2_R1200_U419,
    new_P2_R1200_U420, new_P2_R1200_U421, new_P2_R1200_U422,
    new_P2_R1200_U423, new_P2_R1200_U424, new_P2_R1200_U425,
    new_P2_R1200_U426, new_P2_R1200_U427, new_P2_R1200_U428,
    new_P2_R1200_U429, new_P2_R1200_U430, new_P2_R1200_U431,
    new_P2_R1200_U432, new_P2_R1200_U433, new_P2_R1200_U434,
    new_P2_R1200_U435, new_P2_R1200_U436, new_P2_R1200_U437,
    new_P2_R1200_U438, new_P2_R1200_U439, new_P2_R1200_U440,
    new_P2_R1200_U441, new_P2_R1200_U442, new_P2_R1200_U443,
    new_P2_R1200_U444, new_P2_R1200_U445, new_P2_R1200_U446,
    new_P2_R1200_U447, new_P2_R1200_U448, new_P2_R1200_U449,
    new_P2_R1200_U450, new_P2_R1200_U451, new_P2_R1200_U452,
    new_P2_R1200_U453, new_P2_R1200_U454, new_P2_R1200_U455,
    new_P2_R1200_U456, new_P2_R1200_U457, new_P2_R1200_U458,
    new_P2_R1200_U459, new_P2_R1200_U460, new_P2_R1200_U461,
    new_P2_R1200_U462, new_P2_R1200_U463, new_P2_R1200_U464,
    new_P2_R1200_U465, new_P2_R1200_U466, new_P2_R1200_U467,
    new_P2_R1200_U468, new_P2_R1200_U469, new_P2_R1200_U470,
    new_P2_R1200_U471, new_P2_R1200_U472, new_P2_R1200_U473,
    new_P2_R1200_U474, new_P2_R1200_U475, new_P2_R1200_U476,
    new_P2_R1200_U477, new_P2_R1200_U478, new_P2_R1200_U479,
    new_P2_R1200_U480, new_P2_R1200_U481, new_P2_R1200_U482,
    new_P2_R1200_U483, new_P2_R1200_U484, new_P2_R1200_U485,
    new_P2_R1200_U486, new_P2_R1200_U487, new_P2_R1200_U488,
    new_P2_R1200_U489, new_P2_R1179_U6, new_P2_R1179_U7, new_P2_R1179_U8,
    new_P2_R1179_U9, new_P2_R1179_U10, new_P2_R1179_U11, new_P2_R1179_U12,
    new_P2_R1179_U13, new_P2_R1179_U14, new_P2_R1179_U15, new_P2_R1179_U16,
    new_P2_R1179_U17, new_P2_R1179_U18, new_P2_R1179_U19, new_P2_R1179_U20,
    new_P2_R1179_U21, new_P2_R1179_U22, new_P2_R1179_U23, new_P2_R1179_U24,
    new_P2_R1179_U25, new_P2_R1179_U26, new_P2_R1179_U27, new_P2_R1179_U28,
    new_P2_R1179_U29, new_P2_R1179_U30, new_P2_R1179_U31, new_P2_R1179_U32,
    new_P2_R1179_U33, new_P2_R1179_U34, new_P2_R1179_U35, new_P2_R1179_U36,
    new_P2_R1179_U37, new_P2_R1179_U38, new_P2_R1179_U39, new_P2_R1179_U40,
    new_P2_R1179_U41, new_P2_R1179_U42, new_P2_R1179_U43, new_P2_R1179_U44,
    new_P2_R1179_U45, new_P2_R1179_U46, new_P2_R1179_U47, new_P2_R1179_U48,
    new_P2_R1179_U49, new_P2_R1179_U50, new_P2_R1179_U51, new_P2_R1179_U52,
    new_P2_R1179_U53, new_P2_R1179_U54, new_P2_R1179_U55, new_P2_R1179_U56,
    new_P2_R1179_U57, new_P2_R1179_U58, new_P2_R1179_U59, new_P2_R1179_U60,
    new_P2_R1179_U61, new_P2_R1179_U62, new_P2_R1179_U63, new_P2_R1179_U64,
    new_P2_R1179_U65, new_P2_R1179_U66, new_P2_R1179_U67, new_P2_R1179_U68,
    new_P2_R1179_U69, new_P2_R1179_U70, new_P2_R1179_U71, new_P2_R1179_U72,
    new_P2_R1179_U73, new_P2_R1179_U74, new_P2_R1179_U75, new_P2_R1179_U76,
    new_P2_R1179_U77, new_P2_R1179_U78, new_P2_R1179_U79, new_P2_R1179_U80,
    new_P2_R1179_U81, new_P2_R1179_U82, new_P2_R1179_U83, new_P2_R1179_U84,
    new_P2_R1179_U85, new_P2_R1179_U86, new_P2_R1179_U87, new_P2_R1179_U88,
    new_P2_R1179_U89, new_P2_R1179_U90, new_P2_R1179_U91, new_P2_R1179_U92,
    new_P2_R1179_U93, new_P2_R1179_U94, new_P2_R1179_U95, new_P2_R1179_U96,
    new_P2_R1179_U97, new_P2_R1179_U98, new_P2_R1179_U99,
    new_P2_R1179_U100, new_P2_R1179_U101, new_P2_R1179_U102,
    new_P2_R1179_U103, new_P2_R1179_U104, new_P2_R1179_U105,
    new_P2_R1179_U106, new_P2_R1179_U107, new_P2_R1179_U108,
    new_P2_R1179_U109, new_P2_R1179_U110, new_P2_R1179_U111,
    new_P2_R1179_U112, new_P2_R1179_U113, new_P2_R1179_U114,
    new_P2_R1179_U115, new_P2_R1179_U116, new_P2_R1179_U117,
    new_P2_R1179_U118, new_P2_R1179_U119, new_P2_R1179_U120,
    new_P2_R1179_U121, new_P2_R1179_U122, new_P2_R1179_U123,
    new_P2_R1179_U124, new_P2_R1179_U125, new_P2_R1179_U126,
    new_P2_R1179_U127, new_P2_R1179_U128, new_P2_R1179_U129,
    new_P2_R1179_U130, new_P2_R1179_U131, new_P2_R1179_U132,
    new_P2_R1179_U133, new_P2_R1179_U134, new_P2_R1179_U135,
    new_P2_R1179_U136, new_P2_R1179_U137, new_P2_R1179_U138,
    new_P2_R1179_U139, new_P2_R1179_U140, new_P2_R1179_U141,
    new_P2_R1179_U142, new_P2_R1179_U143, new_P2_R1179_U144,
    new_P2_R1179_U145, new_P2_R1179_U146, new_P2_R1179_U147,
    new_P2_R1179_U148, new_P2_R1179_U149, new_P2_R1179_U150,
    new_P2_R1179_U151, new_P2_R1179_U152, new_P2_R1179_U153,
    new_P2_R1179_U154, new_P2_R1179_U155, new_P2_R1179_U156,
    new_P2_R1179_U157, new_P2_R1179_U158, new_P2_R1179_U159,
    new_P2_R1179_U160, new_P2_R1179_U161, new_P2_R1179_U162,
    new_P2_R1179_U163, new_P2_R1179_U164, new_P2_R1179_U165,
    new_P2_R1179_U166, new_P2_R1179_U167, new_P2_R1179_U168,
    new_P2_R1179_U169, new_P2_R1179_U170, new_P2_R1179_U171,
    new_P2_R1179_U172, new_P2_R1179_U173, new_P2_R1179_U174,
    new_P2_R1179_U175, new_P2_R1179_U176, new_P2_R1179_U177,
    new_P2_R1179_U178, new_P2_R1179_U179, new_P2_R1179_U180,
    new_P2_R1179_U181, new_P2_R1179_U182, new_P2_R1179_U183,
    new_P2_R1179_U184, new_P2_R1179_U185, new_P2_R1179_U186,
    new_P2_R1179_U187, new_P2_R1179_U188, new_P2_R1179_U189,
    new_P2_R1179_U190, new_P2_R1179_U191, new_P2_R1179_U192,
    new_P2_R1179_U193, new_P2_R1179_U194, new_P2_R1179_U195,
    new_P2_R1179_U196, new_P2_R1179_U197, new_P2_R1179_U198,
    new_P2_R1179_U199, new_P2_R1179_U200, new_P2_R1179_U201,
    new_P2_R1179_U202, new_P2_R1179_U203, new_P2_R1179_U204,
    new_P2_R1179_U205, new_P2_R1179_U206, new_P2_R1179_U207,
    new_P2_R1179_U208, new_P2_R1179_U209, new_P2_R1179_U210,
    new_P2_R1179_U211, new_P2_R1179_U212, new_P2_R1179_U213,
    new_P2_R1179_U214, new_P2_R1179_U215, new_P2_R1179_U216,
    new_P2_R1179_U217, new_P2_R1179_U218, new_P2_R1179_U219,
    new_P2_R1179_U220, new_P2_R1179_U221, new_P2_R1179_U222,
    new_P2_R1179_U223, new_P2_R1179_U224, new_P2_R1179_U225,
    new_P2_R1179_U226, new_P2_R1179_U227, new_P2_R1179_U228,
    new_P2_R1179_U229, new_P2_R1179_U230, new_P2_R1179_U231,
    new_P2_R1179_U232, new_P2_R1179_U233, new_P2_R1179_U234,
    new_P2_R1179_U235, new_P2_R1179_U236, new_P2_R1179_U237,
    new_P2_R1179_U238, new_P2_R1179_U239, new_P2_R1179_U240,
    new_P2_R1179_U241, new_P2_R1179_U242, new_P2_R1179_U243,
    new_P2_R1179_U244, new_P2_R1179_U245, new_P2_R1179_U246,
    new_P2_R1179_U247, new_P2_R1179_U248, new_P2_R1179_U249,
    new_P2_R1179_U250, new_P2_R1179_U251, new_P2_R1179_U252,
    new_P2_R1179_U253, new_P2_R1179_U254, new_P2_R1179_U255,
    new_P2_R1179_U256, new_P2_R1179_U257, new_P2_R1179_U258,
    new_P2_R1179_U259, new_P2_R1179_U260, new_P2_R1179_U261,
    new_P2_R1179_U262, new_P2_R1179_U263, new_P2_R1179_U264,
    new_P2_R1179_U265, new_P2_R1179_U266, new_P2_R1179_U267,
    new_P2_R1179_U268, new_P2_R1179_U269, new_P2_R1179_U270,
    new_P2_R1179_U271, new_P2_R1179_U272, new_P2_R1179_U273,
    new_P2_R1179_U274, new_P2_R1179_U275, new_P2_R1179_U276,
    new_P2_R1179_U277, new_P2_R1179_U278, new_P2_R1179_U279,
    new_P2_R1179_U280, new_P2_R1179_U281, new_P2_R1179_U282,
    new_P2_R1179_U283, new_P2_R1179_U284, new_P2_R1179_U285,
    new_P2_R1179_U286, new_P2_R1179_U287, new_P2_R1179_U288,
    new_P2_R1179_U289, new_P2_R1179_U290, new_P2_R1179_U291,
    new_P2_R1179_U292, new_P2_R1179_U293, new_P2_R1179_U294,
    new_P2_R1179_U295, new_P2_R1179_U296, new_P2_R1179_U297,
    new_P2_R1179_U298, new_P2_R1179_U299, new_P2_R1179_U300,
    new_P2_R1179_U301, new_P2_R1179_U302, new_P2_R1179_U303,
    new_P2_R1179_U304, new_P2_R1179_U305, new_P2_R1179_U306,
    new_P2_R1179_U307, new_P2_R1179_U308, new_P2_R1179_U309,
    new_P2_R1179_U310, new_P2_R1179_U311, new_P2_R1179_U312,
    new_P2_R1179_U313, new_P2_R1179_U314, new_P2_R1179_U315,
    new_P2_R1179_U316, new_P2_R1179_U317, new_P2_R1179_U318,
    new_P2_R1179_U319, new_P2_R1179_U320, new_P2_R1179_U321,
    new_P2_R1179_U322, new_P2_R1179_U323, new_P2_R1179_U324,
    new_P2_R1179_U325, new_P2_R1179_U326, new_P2_R1179_U327,
    new_P2_R1179_U328, new_P2_R1179_U329, new_P2_R1179_U330,
    new_P2_R1179_U331, new_P2_R1179_U332, new_P2_R1179_U333,
    new_P2_R1179_U334, new_P2_R1179_U335, new_P2_R1179_U336,
    new_P2_R1179_U337, new_P2_R1179_U338, new_P2_R1179_U339,
    new_P2_R1179_U340, new_P2_R1179_U341, new_P2_R1179_U342,
    new_P2_R1179_U343, new_P2_R1179_U344, new_P2_R1179_U345,
    new_P2_R1179_U346, new_P2_R1179_U347, new_P2_R1179_U348,
    new_P2_R1179_U349, new_P2_R1179_U350, new_P2_R1179_U351,
    new_P2_R1179_U352, new_P2_R1179_U353, new_P2_R1179_U354,
    new_P2_R1179_U355, new_P2_R1179_U356, new_P2_R1179_U357,
    new_P2_R1179_U358, new_P2_R1179_U359, new_P2_R1179_U360,
    new_P2_R1179_U361, new_P2_R1179_U362, new_P2_R1179_U363,
    new_P2_R1179_U364, new_P2_R1179_U365, new_P2_R1179_U366,
    new_P2_R1179_U367, new_P2_R1179_U368, new_P2_R1179_U369,
    new_P2_R1179_U370, new_P2_R1179_U371, new_P2_R1179_U372,
    new_P2_R1179_U373, new_P2_R1179_U374, new_P2_R1179_U375,
    new_P2_R1179_U376, new_P2_R1179_U377, new_P2_R1179_U378,
    new_P2_R1179_U379, new_P2_R1179_U380, new_P2_R1179_U381,
    new_P2_R1179_U382, new_P2_R1179_U383, new_P2_R1179_U384,
    new_P2_R1179_U385, new_P2_R1179_U386, new_P2_R1179_U387,
    new_P2_R1179_U388, new_P2_R1179_U389, new_P2_R1179_U390,
    new_P2_R1179_U391, new_P2_R1179_U392, new_P2_R1179_U393,
    new_P2_R1179_U394, new_P2_R1179_U395, new_P2_R1179_U396,
    new_P2_R1179_U397, new_P2_R1179_U398, new_P2_R1179_U399,
    new_P2_R1179_U400, new_P2_R1179_U401, new_P2_R1179_U402,
    new_P2_R1179_U403, new_P2_R1179_U404, new_P2_R1179_U405,
    new_P2_R1179_U406, new_P2_R1179_U407, new_P2_R1179_U408,
    new_P2_R1179_U409, new_P2_R1179_U410, new_P2_R1179_U411,
    new_P2_R1179_U412, new_P2_R1179_U413, new_P2_R1179_U414,
    new_P2_R1179_U415, new_P2_R1179_U416, new_P2_R1179_U417,
    new_P2_R1179_U418, new_P2_R1179_U419, new_P2_R1179_U420,
    new_P2_R1179_U421, new_P2_R1179_U422, new_P2_R1179_U423,
    new_P2_R1179_U424, new_P2_R1179_U425, new_P2_R1179_U426,
    new_P2_R1179_U427, new_P2_R1179_U428, new_P2_R1179_U429,
    new_P2_R1179_U430, new_P2_R1179_U431, new_P2_R1179_U432,
    new_P2_R1179_U433, new_P2_R1179_U434, new_P2_R1179_U435,
    new_P2_R1179_U436, new_P2_R1179_U437, new_P2_R1179_U438,
    new_P2_R1179_U439, new_P2_R1179_U440, new_P2_R1179_U441,
    new_P2_R1179_U442, new_P2_R1179_U443, new_P2_R1179_U444,
    new_P2_R1179_U445, new_P2_R1179_U446, new_P2_R1179_U447,
    new_P2_R1179_U448, new_P2_R1179_U449, new_P2_R1179_U450,
    new_P2_R1179_U451, new_P2_R1179_U452, new_P2_R1179_U453,
    new_P2_R1179_U454, new_P2_R1179_U455, new_P2_R1179_U456,
    new_P2_R1179_U457, new_P2_R1179_U458, new_P2_R1179_U459,
    new_P2_R1179_U460, new_P2_R1179_U461, new_P2_R1179_U462,
    new_P2_R1179_U463, new_P2_R1179_U464, new_P2_R1179_U465,
    new_P2_R1179_U466, new_P2_R1179_U467, new_P2_R1179_U468,
    new_P2_R1179_U469, new_P2_R1179_U470, new_P2_R1179_U471,
    new_P2_R1179_U472, new_P2_R1179_U473, new_P2_R1179_U474,
    new_P2_R1179_U475, new_P2_R1179_U476, new_P2_R1179_U477,
    new_P2_R1179_U478, new_P2_R1179_U479, new_P2_R1179_U480,
    new_P2_R1179_U481, new_P2_R1179_U482, new_P2_R1179_U483,
    new_P2_R1179_U484, new_P2_R1179_U485, new_P2_R1179_U486,
    new_P2_R1179_U487, new_P2_R1179_U488, new_P2_R1179_U489,
    new_P2_R1269_U6, new_P2_R1269_U7, new_P2_R1269_U8, new_P2_R1269_U9,
    new_P2_R1269_U10, new_P2_R1269_U11, new_P2_R1269_U12, new_P2_R1269_U13,
    new_P2_R1269_U14, new_P2_R1269_U15, new_P2_R1269_U16, new_P2_R1269_U17,
    new_P2_R1269_U18, new_P2_R1269_U19, new_P2_R1269_U20, new_P2_R1269_U21,
    new_P2_R1269_U22, new_P2_R1269_U23, new_P2_R1269_U24, new_P2_R1269_U25,
    new_P2_R1269_U26, new_P2_R1269_U27, new_P2_R1269_U28, new_P2_R1269_U29,
    new_P2_R1269_U30, new_P2_R1269_U31, new_P2_R1269_U32, new_P2_R1269_U33,
    new_P2_R1269_U34, new_P2_R1269_U35, new_P2_R1269_U36, new_P2_R1269_U37,
    new_P2_R1269_U38, new_P2_R1269_U39, new_P2_R1269_U40, new_P2_R1269_U41,
    new_P2_R1269_U42, new_P2_R1269_U43, new_P2_R1269_U44, new_P2_R1269_U45,
    new_P2_R1269_U46, new_P2_R1269_U47, new_P2_R1269_U48, new_P2_R1269_U49,
    new_P2_R1269_U50, new_P2_R1269_U51, new_P2_R1269_U52, new_P2_R1269_U53,
    new_P2_R1269_U54, new_P2_R1269_U55, new_P2_R1269_U56, new_P2_R1269_U57,
    new_P2_R1269_U58, new_P2_R1269_U59, new_P2_R1269_U60, new_P2_R1269_U61,
    new_P2_R1269_U62, new_P2_R1269_U63, new_P2_R1269_U64, new_P2_R1269_U65,
    new_P2_R1269_U66, new_P2_R1269_U67, new_P2_R1269_U68, new_P2_R1269_U69,
    new_P2_R1269_U70, new_P2_R1269_U71, new_P2_R1269_U72, new_P2_R1269_U73,
    new_P2_R1269_U74, new_P2_R1269_U75, new_P2_R1269_U76, new_P2_R1269_U77,
    new_P2_R1269_U78, new_P2_R1269_U79, new_P2_R1269_U80, new_P2_R1269_U81,
    new_P2_R1269_U82, new_P2_R1269_U83, new_P2_R1269_U84, new_P2_R1269_U85,
    new_P2_R1269_U86, new_P2_R1269_U87, new_P2_R1269_U88, new_P2_R1269_U89,
    new_P2_R1269_U90, new_P2_R1269_U91, new_P2_R1269_U92, new_P2_R1269_U93,
    new_P2_R1269_U94, new_P2_R1269_U95, new_P2_R1269_U96, new_P2_R1269_U97,
    new_P2_R1269_U98, new_P2_R1269_U99, new_P2_R1269_U100,
    new_P2_R1269_U101, new_P2_R1269_U102, new_P2_R1269_U103,
    new_P2_R1269_U104, new_P2_R1269_U105, new_P2_R1269_U106,
    new_P2_R1269_U107, new_P2_R1269_U108, new_P2_R1269_U109,
    new_P2_R1269_U110, new_P2_R1269_U111, new_P2_R1269_U112,
    new_P2_R1269_U113, new_P2_R1269_U114, new_P2_R1269_U115,
    new_P2_R1269_U116, new_P2_R1269_U117, new_P2_R1269_U118,
    new_P2_R1269_U119, new_P2_R1269_U120, new_P2_R1269_U121,
    new_P2_R1269_U122, new_P2_R1269_U123, new_P2_R1269_U124,
    new_P2_R1269_U125, new_P2_R1269_U126, new_P2_R1269_U127,
    new_P2_R1269_U128, new_P2_R1269_U129, new_P2_R1269_U130,
    new_P2_R1269_U131, new_P2_R1269_U132, new_P2_R1269_U133,
    new_P2_R1269_U134, new_P2_R1269_U135, new_P2_R1269_U136,
    new_P2_R1269_U137, new_P2_R1269_U138, new_P2_R1269_U139,
    new_P2_R1269_U140, new_P2_R1269_U141, new_P2_R1269_U142,
    new_P2_R1269_U143, new_P2_R1269_U144, new_P2_R1269_U145,
    new_P2_R1269_U146, new_P2_R1269_U147, new_P2_R1269_U148,
    new_P2_R1269_U149, new_P2_R1269_U150, new_P2_R1269_U151,
    new_P2_R1269_U152, new_P2_R1269_U153, new_P2_R1269_U154,
    new_P2_R1269_U155, new_P2_R1269_U156, new_P2_R1269_U157,
    new_P2_R1269_U158, new_P2_R1269_U159, new_P2_R1269_U160,
    new_P2_R1269_U161, new_P2_R1269_U162, new_P2_R1269_U163,
    new_P2_R1269_U164, new_P2_R1269_U165, new_P2_R1269_U166,
    new_P2_R1269_U167, new_P2_R1269_U168, new_P2_R1269_U169,
    new_P2_R1269_U170, new_P2_R1269_U171, new_P2_R1269_U172,
    new_P2_R1269_U173, new_P2_R1269_U174, new_P2_R1269_U175,
    new_P2_R1269_U176, new_P2_R1269_U177, new_P2_R1269_U178,
    new_P2_R1269_U179, new_P2_R1269_U180, new_P2_R1269_U181,
    new_P2_R1269_U182, new_P2_R1269_U183, new_P2_R1269_U184,
    new_P2_R1269_U185, new_P2_R1269_U186, new_P2_R1269_U187,
    new_P2_R1269_U188, new_P2_R1269_U189, new_P2_R1269_U190,
    new_P2_R1269_U191, new_P2_R1269_U192, new_P2_R1269_U193,
    new_P2_R1269_U194, new_P2_R1269_U195, new_P2_R1269_U196,
    new_P2_R1269_U197, new_P2_R1269_U198, new_P2_R1269_U199,
    new_P2_R1269_U200, new_P2_R1269_U201, new_P2_R1269_U202,
    new_P2_R1269_U203, new_P2_R1269_U204, new_P2_R1269_U205,
    new_P2_R1269_U206, new_P2_R1269_U207, new_P2_R1269_U208,
    new_P2_R1269_U209, new_P2_R1110_U4, new_P2_R1110_U5, new_P2_R1110_U6,
    new_P2_R1110_U7, new_P2_R1110_U8, new_P2_R1110_U9, new_P2_R1110_U10,
    new_P2_R1110_U11, new_P2_R1110_U12, new_P2_R1110_U13, new_P2_R1110_U14,
    new_P2_R1110_U15, new_P2_R1110_U16, new_P2_R1110_U17, new_P2_R1110_U18,
    new_P2_R1110_U19, new_P2_R1110_U20, new_P2_R1110_U21, new_P2_R1110_U22,
    new_P2_R1110_U23, new_P2_R1110_U24, new_P2_R1110_U25, new_P2_R1110_U26,
    new_P2_R1110_U27, new_P2_R1110_U28, new_P2_R1110_U29, new_P2_R1110_U30,
    new_P2_R1110_U31, new_P2_R1110_U32, new_P2_R1110_U33, new_P2_R1110_U34,
    new_P2_R1110_U35, new_P2_R1110_U36, new_P2_R1110_U37, new_P2_R1110_U38,
    new_P2_R1110_U39, new_P2_R1110_U40, new_P2_R1110_U41, new_P2_R1110_U42,
    new_P2_R1110_U43, new_P2_R1110_U44, new_P2_R1110_U45, new_P2_R1110_U46,
    new_P2_R1110_U47, new_P2_R1110_U48, new_P2_R1110_U49, new_P2_R1110_U50,
    new_P2_R1110_U51, new_P2_R1110_U52, new_P2_R1110_U53, new_P2_R1110_U54,
    new_P2_R1110_U55, new_P2_R1110_U56, new_P2_R1110_U57, new_P2_R1110_U58,
    new_P2_R1110_U59, new_P2_R1110_U60, new_P2_R1110_U61, new_P2_R1110_U62,
    new_P2_R1110_U63, new_P2_R1110_U64, new_P2_R1110_U65, new_P2_R1110_U66,
    new_P2_R1110_U67, new_P2_R1110_U68, new_P2_R1110_U69, new_P2_R1110_U70,
    new_P2_R1110_U71, new_P2_R1110_U72, new_P2_R1110_U73, new_P2_R1110_U74,
    new_P2_R1110_U75, new_P2_R1110_U76, new_P2_R1110_U77, new_P2_R1110_U78,
    new_P2_R1110_U79, new_P2_R1110_U80, new_P2_R1110_U81, new_P2_R1110_U82,
    new_P2_R1110_U83, new_P2_R1110_U84, new_P2_R1110_U85, new_P2_R1110_U86,
    new_P2_R1110_U87, new_P2_R1110_U88, new_P2_R1110_U89, new_P2_R1110_U90,
    new_P2_R1110_U91, new_P2_R1110_U92, new_P2_R1110_U93, new_P2_R1110_U94,
    new_P2_R1110_U95, new_P2_R1110_U96, new_P2_R1110_U97, new_P2_R1110_U98,
    new_P2_R1110_U99, new_P2_R1110_U100, new_P2_R1110_U101,
    new_P2_R1110_U102, new_P2_R1110_U103, new_P2_R1110_U104,
    new_P2_R1110_U105, new_P2_R1110_U106, new_P2_R1110_U107,
    new_P2_R1110_U108, new_P2_R1110_U109, new_P2_R1110_U110,
    new_P2_R1110_U111, new_P2_R1110_U112, new_P2_R1110_U113,
    new_P2_R1110_U114, new_P2_R1110_U115, new_P2_R1110_U116,
    new_P2_R1110_U117, new_P2_R1110_U118, new_P2_R1110_U119,
    new_P2_R1110_U120, new_P2_R1110_U121, new_P2_R1110_U122,
    new_P2_R1110_U123, new_P2_R1110_U124, new_P2_R1110_U125,
    new_P2_R1110_U126, new_P2_R1110_U127, new_P2_R1110_U128,
    new_P2_R1110_U129, new_P2_R1110_U130, new_P2_R1110_U131,
    new_P2_R1110_U132, new_P2_R1110_U133, new_P2_R1110_U134,
    new_P2_R1110_U135, new_P2_R1110_U136, new_P2_R1110_U137,
    new_P2_R1110_U138, new_P2_R1110_U139, new_P2_R1110_U140,
    new_P2_R1110_U141, new_P2_R1110_U142, new_P2_R1110_U143,
    new_P2_R1110_U144, new_P2_R1110_U145, new_P2_R1110_U146,
    new_P2_R1110_U147, new_P2_R1110_U148, new_P2_R1110_U149,
    new_P2_R1110_U150, new_P2_R1110_U151, new_P2_R1110_U152,
    new_P2_R1110_U153, new_P2_R1110_U154, new_P2_R1110_U155,
    new_P2_R1110_U156, new_P2_R1110_U157, new_P2_R1110_U158,
    new_P2_R1110_U159, new_P2_R1110_U160, new_P2_R1110_U161,
    new_P2_R1110_U162, new_P2_R1110_U163, new_P2_R1110_U164,
    new_P2_R1110_U165, new_P2_R1110_U166, new_P2_R1110_U167,
    new_P2_R1110_U168, new_P2_R1110_U169, new_P2_R1110_U170,
    new_P2_R1110_U171, new_P2_R1110_U172, new_P2_R1110_U173,
    new_P2_R1110_U174, new_P2_R1110_U175, new_P2_R1110_U176,
    new_P2_R1110_U177, new_P2_R1110_U178, new_P2_R1110_U179,
    new_P2_R1110_U180, new_P2_R1110_U181, new_P2_R1110_U182,
    new_P2_R1110_U183, new_P2_R1110_U184, new_P2_R1110_U185,
    new_P2_R1110_U186, new_P2_R1110_U187, new_P2_R1110_U188,
    new_P2_R1110_U189, new_P2_R1110_U190, new_P2_R1110_U191,
    new_P2_R1110_U192, new_P2_R1110_U193, new_P2_R1110_U194,
    new_P2_R1110_U195, new_P2_R1110_U196, new_P2_R1110_U197,
    new_P2_R1110_U198, new_P2_R1110_U199, new_P2_R1110_U200,
    new_P2_R1110_U201, new_P2_R1110_U202, new_P2_R1110_U203,
    new_P2_R1110_U204, new_P2_R1110_U205, new_P2_R1110_U206,
    new_P2_R1110_U207, new_P2_R1110_U208, new_P2_R1110_U209,
    new_P2_R1110_U210, new_P2_R1110_U211, new_P2_R1110_U212,
    new_P2_R1110_U213, new_P2_R1110_U214, new_P2_R1110_U215,
    new_P2_R1110_U216, new_P2_R1110_U217, new_P2_R1110_U218,
    new_P2_R1110_U219, new_P2_R1110_U220, new_P2_R1110_U221,
    new_P2_R1110_U222, new_P2_R1110_U223, new_P2_R1110_U224,
    new_P2_R1110_U225, new_P2_R1110_U226, new_P2_R1110_U227,
    new_P2_R1110_U228, new_P2_R1110_U229, new_P2_R1110_U230,
    new_P2_R1110_U231, new_P2_R1110_U232, new_P2_R1110_U233,
    new_P2_R1110_U234, new_P2_R1110_U235, new_P2_R1110_U236,
    new_P2_R1110_U237, new_P2_R1110_U238, new_P2_R1110_U239,
    new_P2_R1110_U240, new_P2_R1110_U241, new_P2_R1110_U242,
    new_P2_R1110_U243, new_P2_R1110_U244, new_P2_R1110_U245,
    new_P2_R1110_U246, new_P2_R1110_U247, new_P2_R1110_U248,
    new_P2_R1110_U249, new_P2_R1110_U250, new_P2_R1110_U251,
    new_P2_R1110_U252, new_P2_R1110_U253, new_P2_R1110_U254,
    new_P2_R1110_U255, new_P2_R1110_U256, new_P2_R1110_U257,
    new_P2_R1110_U258, new_P2_R1110_U259, new_P2_R1110_U260,
    new_P2_R1110_U261, new_P2_R1110_U262, new_P2_R1110_U263,
    new_P2_R1110_U264, new_P2_R1110_U265, new_P2_R1110_U266,
    new_P2_R1110_U267, new_P2_R1110_U268, new_P2_R1110_U269,
    new_P2_R1110_U270, new_P2_R1110_U271, new_P2_R1110_U272,
    new_P2_R1110_U273, new_P2_R1110_U274, new_P2_R1110_U275,
    new_P2_R1110_U276, new_P2_R1110_U277, new_P2_R1110_U278,
    new_P2_R1110_U279, new_P2_R1110_U280, new_P2_R1110_U281,
    new_P2_R1110_U282, new_P2_R1110_U283, new_P2_R1110_U284,
    new_P2_R1110_U285, new_P2_R1110_U286, new_P2_R1110_U287,
    new_P2_R1110_U288, new_P2_R1110_U289, new_P2_R1110_U290,
    new_P2_R1110_U291, new_P2_R1110_U292, new_P2_R1110_U293,
    new_P2_R1110_U294, new_P2_R1110_U295, new_P2_R1110_U296,
    new_P2_R1110_U297, new_P2_R1110_U298, new_P2_R1110_U299,
    new_P2_R1110_U300, new_P2_R1110_U301, new_P2_R1110_U302,
    new_P2_R1110_U303, new_P2_R1110_U304, new_P2_R1110_U305,
    new_P2_R1110_U306, new_P2_R1110_U307, new_P2_R1110_U308,
    new_P2_R1110_U309, new_P2_R1110_U310, new_P2_R1110_U311,
    new_P2_R1110_U312, new_P2_R1110_U313, new_P2_R1110_U314,
    new_P2_R1110_U315, new_P2_R1110_U316, new_P2_R1110_U317,
    new_P2_R1110_U318, new_P2_R1110_U319, new_P2_R1110_U320,
    new_P2_R1110_U321, new_P2_R1110_U322, new_P2_R1110_U323,
    new_P2_R1110_U324, new_P2_R1110_U325, new_P2_R1110_U326,
    new_P2_R1110_U327, new_P2_R1110_U328, new_P2_R1110_U329,
    new_P2_R1110_U330, new_P2_R1110_U331, new_P2_R1110_U332,
    new_P2_R1110_U333, new_P2_R1110_U334, new_P2_R1110_U335,
    new_P2_R1110_U336, new_P2_R1110_U337, new_P2_R1110_U338,
    new_P2_R1110_U339, new_P2_R1110_U340, new_P2_R1110_U341,
    new_P2_R1110_U342, new_P2_R1110_U343, new_P2_R1110_U344,
    new_P2_R1110_U345, new_P2_R1110_U346, new_P2_R1110_U347,
    new_P2_R1110_U348, new_P2_R1110_U349, new_P2_R1110_U350,
    new_P2_R1110_U351, new_P2_R1110_U352, new_P2_R1110_U353,
    new_P2_R1110_U354, new_P2_R1110_U355, new_P2_R1110_U356,
    new_P2_R1110_U357, new_P2_R1110_U358, new_P2_R1110_U359,
    new_P2_R1110_U360, new_P2_R1110_U361, new_P2_R1110_U362,
    new_P2_R1110_U363, new_P2_R1110_U364, new_P2_R1110_U365,
    new_P2_R1110_U366, new_P2_R1110_U367, new_P2_R1110_U368,
    new_P2_R1110_U369, new_P2_R1110_U370, new_P2_R1110_U371,
    new_P2_R1110_U372, new_P2_R1110_U373, new_P2_R1110_U374,
    new_P2_R1110_U375, new_P2_R1110_U376, new_P2_R1110_U377,
    new_P2_R1110_U378, new_P2_R1110_U379, new_P2_R1110_U380,
    new_P2_R1110_U381, new_P2_R1110_U382, new_P2_R1110_U383,
    new_P2_R1110_U384, new_P2_R1110_U385, new_P2_R1110_U386,
    new_P2_R1110_U387, new_P2_R1110_U388, new_P2_R1110_U389,
    new_P2_R1110_U390, new_P2_R1110_U391, new_P2_R1110_U392,
    new_P2_R1110_U393, new_P2_R1110_U394, new_P2_R1110_U395,
    new_P2_R1110_U396, new_P2_R1110_U397, new_P2_R1110_U398,
    new_P2_R1110_U399, new_P2_R1110_U400, new_P2_R1110_U401,
    new_P2_R1110_U402, new_P2_R1110_U403, new_P2_R1110_U404,
    new_P2_R1110_U405, new_P2_R1110_U406, new_P2_R1110_U407,
    new_P2_R1110_U408, new_P2_R1110_U409, new_P2_R1110_U410,
    new_P2_R1110_U411, new_P2_R1110_U412, new_P2_R1110_U413,
    new_P2_R1110_U414, new_P2_R1110_U415, new_P2_R1110_U416,
    new_P2_R1110_U417, new_P2_R1110_U418, new_P2_R1110_U419,
    new_P2_R1110_U420, new_P2_R1110_U421, new_P2_R1110_U422,
    new_P2_R1110_U423, new_P2_R1110_U424, new_P2_R1110_U425,
    new_P2_R1110_U426, new_P2_R1110_U427, new_P2_R1110_U428,
    new_P2_R1110_U429, new_P2_R1110_U430, new_P2_R1110_U431,
    new_P2_R1110_U432, new_P2_R1110_U433, new_P2_R1110_U434,
    new_P2_R1110_U435, new_P2_R1110_U436, new_P2_R1110_U437,
    new_P2_R1110_U438, new_P2_R1110_U439, new_P2_R1110_U440,
    new_P2_R1110_U441, new_P2_R1110_U442, new_P2_R1110_U443,
    new_P2_R1110_U444, new_P2_R1110_U445, new_P2_R1110_U446,
    new_P2_R1110_U447, new_P2_R1110_U448, new_P2_R1110_U449,
    new_P2_R1110_U450, new_P2_R1110_U451, new_P2_R1110_U452,
    new_P2_R1110_U453, new_P2_R1110_U454, new_P2_R1110_U455,
    new_P2_R1110_U456, new_P2_R1110_U457, new_P2_R1110_U458,
    new_P2_R1110_U459, new_P2_R1110_U460, new_P2_R1110_U461,
    new_P2_R1110_U462, new_P2_R1110_U463, new_P2_R1110_U464,
    new_P2_R1110_U465, new_P2_R1110_U466, new_P2_R1110_U467,
    new_P2_R1110_U468, new_P2_R1110_U469, new_P2_R1110_U470,
    new_P2_R1110_U471, new_P2_R1110_U472, new_P2_R1110_U473,
    new_P2_R1110_U474, new_P2_R1110_U475, new_P2_R1110_U476,
    new_P2_R1110_U477, new_P2_R1110_U478, new_P2_R1110_U479,
    new_P2_R1110_U480, new_P2_R1110_U481, new_P2_R1110_U482,
    new_P2_R1110_U483, new_P2_R1110_U484, new_P2_R1110_U485,
    new_P2_R1110_U486, new_P2_R1110_U487, new_P2_R1110_U488,
    new_P2_R1110_U489, new_P2_R1110_U490, new_P2_R1110_U491,
    new_P2_R1110_U492, new_P2_R1110_U493, new_P2_R1110_U494,
    new_P2_R1110_U495, new_P2_R1110_U496, new_P2_R1110_U497,
    new_P2_R1110_U498, new_P2_R1110_U499, new_P2_R1110_U500,
    new_P2_R1110_U501, new_P2_R1110_U502, new_P2_R1110_U503,
    new_P2_R1110_U504, new_P2_R1297_U6, new_P2_R1297_U7, new_P2_R1077_U4,
    new_P2_R1077_U5, new_P2_R1077_U6, new_P2_R1077_U7, new_P2_R1077_U8,
    new_P2_R1077_U9, new_P2_R1077_U10, new_P2_R1077_U11, new_P2_R1077_U12,
    new_P2_R1077_U13, new_P2_R1077_U14, new_P2_R1077_U15, new_P2_R1077_U16,
    new_P2_R1077_U17, new_P2_R1077_U18, new_P2_R1077_U19, new_P2_R1077_U20,
    new_P2_R1077_U21, new_P2_R1077_U22, new_P2_R1077_U23, new_P2_R1077_U24,
    new_P2_R1077_U25, new_P2_R1077_U26, new_P2_R1077_U27, new_P2_R1077_U28,
    new_P2_R1077_U29, new_P2_R1077_U30, new_P2_R1077_U31, new_P2_R1077_U32,
    new_P2_R1077_U33, new_P2_R1077_U34, new_P2_R1077_U35, new_P2_R1077_U36,
    new_P2_R1077_U37, new_P2_R1077_U38, new_P2_R1077_U39, new_P2_R1077_U40,
    new_P2_R1077_U41, new_P2_R1077_U42, new_P2_R1077_U43, new_P2_R1077_U44,
    new_P2_R1077_U45, new_P2_R1077_U46, new_P2_R1077_U47, new_P2_R1077_U48,
    new_P2_R1077_U49, new_P2_R1077_U50, new_P2_R1077_U51, new_P2_R1077_U52,
    new_P2_R1077_U53, new_P2_R1077_U54, new_P2_R1077_U55, new_P2_R1077_U56,
    new_P2_R1077_U57, new_P2_R1077_U58, new_P2_R1077_U59, new_P2_R1077_U60,
    new_P2_R1077_U61, new_P2_R1077_U62, new_P2_R1077_U63, new_P2_R1077_U64,
    new_P2_R1077_U65, new_P2_R1077_U66, new_P2_R1077_U67, new_P2_R1077_U68,
    new_P2_R1077_U69, new_P2_R1077_U70, new_P2_R1077_U71, new_P2_R1077_U72,
    new_P2_R1077_U73, new_P2_R1077_U74, new_P2_R1077_U75, new_P2_R1077_U76,
    new_P2_R1077_U77, new_P2_R1077_U78, new_P2_R1077_U79, new_P2_R1077_U80,
    new_P2_R1077_U81, new_P2_R1077_U82, new_P2_R1077_U83, new_P2_R1077_U84,
    new_P2_R1077_U85, new_P2_R1077_U86, new_P2_R1077_U87, new_P2_R1077_U88,
    new_P2_R1077_U89, new_P2_R1077_U90, new_P2_R1077_U91, new_P2_R1077_U92,
    new_P2_R1077_U93, new_P2_R1077_U94, new_P2_R1077_U95, new_P2_R1077_U96,
    new_P2_R1077_U97, new_P2_R1077_U98, new_P2_R1077_U99,
    new_P2_R1077_U100, new_P2_R1077_U101, new_P2_R1077_U102,
    new_P2_R1077_U103, new_P2_R1077_U104, new_P2_R1077_U105,
    new_P2_R1077_U106, new_P2_R1077_U107, new_P2_R1077_U108,
    new_P2_R1077_U109, new_P2_R1077_U110, new_P2_R1077_U111,
    new_P2_R1077_U112, new_P2_R1077_U113, new_P2_R1077_U114,
    new_P2_R1077_U115, new_P2_R1077_U116, new_P2_R1077_U117,
    new_P2_R1077_U118, new_P2_R1077_U119, new_P2_R1077_U120,
    new_P2_R1077_U121, new_P2_R1077_U122, new_P2_R1077_U123,
    new_P2_R1077_U124, new_P2_R1077_U125, new_P2_R1077_U126,
    new_P2_R1077_U127, new_P2_R1077_U128, new_P2_R1077_U129,
    new_P2_R1077_U130, new_P2_R1077_U131, new_P2_R1077_U132,
    new_P2_R1077_U133, new_P2_R1077_U134, new_P2_R1077_U135,
    new_P2_R1077_U136, new_P2_R1077_U137, new_P2_R1077_U138,
    new_P2_R1077_U139, new_P2_R1077_U140, new_P2_R1077_U141,
    new_P2_R1077_U142, new_P2_R1077_U143, new_P2_R1077_U144,
    new_P2_R1077_U145, new_P2_R1077_U146, new_P2_R1077_U147,
    new_P2_R1077_U148, new_P2_R1077_U149, new_P2_R1077_U150,
    new_P2_R1077_U151, new_P2_R1077_U152, new_P2_R1077_U153,
    new_P2_R1077_U154, new_P2_R1077_U155, new_P2_R1077_U156,
    new_P2_R1077_U157, new_P2_R1077_U158, new_P2_R1077_U159,
    new_P2_R1077_U160, new_P2_R1077_U161, new_P2_R1077_U162,
    new_P2_R1077_U163, new_P2_R1077_U164, new_P2_R1077_U165,
    new_P2_R1077_U166, new_P2_R1077_U167, new_P2_R1077_U168,
    new_P2_R1077_U169, new_P2_R1077_U170, new_P2_R1077_U171,
    new_P2_R1077_U172, new_P2_R1077_U173, new_P2_R1077_U174,
    new_P2_R1077_U175, new_P2_R1077_U176, new_P2_R1077_U177,
    new_P2_R1077_U178, new_P2_R1077_U179, new_P2_R1077_U180,
    new_P2_R1077_U181, new_P2_R1077_U182, new_P2_R1077_U183,
    new_P2_R1077_U184, new_P2_R1077_U185, new_P2_R1077_U186,
    new_P2_R1077_U187, new_P2_R1077_U188, new_P2_R1077_U189,
    new_P2_R1077_U190, new_P2_R1077_U191, new_P2_R1077_U192,
    new_P2_R1077_U193, new_P2_R1077_U194, new_P2_R1077_U195,
    new_P2_R1077_U196, new_P2_R1077_U197, new_P2_R1077_U198,
    new_P2_R1077_U199, new_P2_R1077_U200, new_P2_R1077_U201,
    new_P2_R1077_U202, new_P2_R1077_U203, new_P2_R1077_U204,
    new_P2_R1077_U205, new_P2_R1077_U206, new_P2_R1077_U207,
    new_P2_R1077_U208, new_P2_R1077_U209, new_P2_R1077_U210,
    new_P2_R1077_U211, new_P2_R1077_U212, new_P2_R1077_U213,
    new_P2_R1077_U214, new_P2_R1077_U215, new_P2_R1077_U216,
    new_P2_R1077_U217, new_P2_R1077_U218, new_P2_R1077_U219,
    new_P2_R1077_U220, new_P2_R1077_U221, new_P2_R1077_U222,
    new_P2_R1077_U223, new_P2_R1077_U224, new_P2_R1077_U225,
    new_P2_R1077_U226, new_P2_R1077_U227, new_P2_R1077_U228,
    new_P2_R1077_U229, new_P2_R1077_U230, new_P2_R1077_U231,
    new_P2_R1077_U232, new_P2_R1077_U233, new_P2_R1077_U234,
    new_P2_R1077_U235, new_P2_R1077_U236, new_P2_R1077_U237,
    new_P2_R1077_U238, new_P2_R1077_U239, new_P2_R1077_U240,
    new_P2_R1077_U241, new_P2_R1077_U242, new_P2_R1077_U243,
    new_P2_R1077_U244, new_P2_R1077_U245, new_P2_R1077_U246,
    new_P2_R1077_U247, new_P2_R1077_U248, new_P2_R1077_U249,
    new_P2_R1077_U250, new_P2_R1077_U251, new_P2_R1077_U252,
    new_P2_R1077_U253, new_P2_R1077_U254, new_P2_R1077_U255,
    new_P2_R1077_U256, new_P2_R1077_U257, new_P2_R1077_U258,
    new_P2_R1077_U259, new_P2_R1077_U260, new_P2_R1077_U261,
    new_P2_R1077_U262, new_P2_R1077_U263, new_P2_R1077_U264,
    new_P2_R1077_U265, new_P2_R1077_U266, new_P2_R1077_U267,
    new_P2_R1077_U268, new_P2_R1077_U269, new_P2_R1077_U270,
    new_P2_R1077_U271, new_P2_R1077_U272, new_P2_R1077_U273,
    new_P2_R1077_U274, new_P2_R1077_U275, new_P2_R1077_U276,
    new_P2_R1077_U277, new_P2_R1077_U278, new_P2_R1077_U279,
    new_P2_R1077_U280, new_P2_R1077_U281, new_P2_R1077_U282,
    new_P2_R1077_U283, new_P2_R1077_U284, new_P2_R1077_U285,
    new_P2_R1077_U286, new_P2_R1077_U287, new_P2_R1077_U288,
    new_P2_R1077_U289, new_P2_R1077_U290, new_P2_R1077_U291,
    new_P2_R1077_U292, new_P2_R1077_U293, new_P2_R1077_U294,
    new_P2_R1077_U295, new_P2_R1077_U296, new_P2_R1077_U297,
    new_P2_R1077_U298, new_P2_R1077_U299, new_P2_R1077_U300,
    new_P2_R1077_U301, new_P2_R1077_U302, new_P2_R1077_U303,
    new_P2_R1077_U304, new_P2_R1077_U305, new_P2_R1077_U306,
    new_P2_R1077_U307, new_P2_R1077_U308, new_P2_R1077_U309,
    new_P2_R1077_U310, new_P2_R1077_U311, new_P2_R1077_U312,
    new_P2_R1077_U313, new_P2_R1077_U314, new_P2_R1077_U315,
    new_P2_R1077_U316, new_P2_R1077_U317, new_P2_R1077_U318,
    new_P2_R1077_U319, new_P2_R1077_U320, new_P2_R1077_U321,
    new_P2_R1077_U322, new_P2_R1077_U323, new_P2_R1077_U324,
    new_P2_R1077_U325, new_P2_R1077_U326, new_P2_R1077_U327,
    new_P2_R1077_U328, new_P2_R1077_U329, new_P2_R1077_U330,
    new_P2_R1077_U331, new_P2_R1077_U332, new_P2_R1077_U333,
    new_P2_R1077_U334, new_P2_R1077_U335, new_P2_R1077_U336,
    new_P2_R1077_U337, new_P2_R1077_U338, new_P2_R1077_U339,
    new_P2_R1077_U340, new_P2_R1077_U341, new_P2_R1077_U342,
    new_P2_R1077_U343, new_P2_R1077_U344, new_P2_R1077_U345,
    new_P2_R1077_U346, new_P2_R1077_U347, new_P2_R1077_U348,
    new_P2_R1077_U349, new_P2_R1077_U350, new_P2_R1077_U351,
    new_P2_R1077_U352, new_P2_R1077_U353, new_P2_R1077_U354,
    new_P2_R1077_U355, new_P2_R1077_U356, new_P2_R1077_U357,
    new_P2_R1077_U358, new_P2_R1077_U359, new_P2_R1077_U360,
    new_P2_R1077_U361, new_P2_R1077_U362, new_P2_R1077_U363,
    new_P2_R1077_U364, new_P2_R1077_U365, new_P2_R1077_U366,
    new_P2_R1077_U367, new_P2_R1077_U368, new_P2_R1077_U369,
    new_P2_R1077_U370, new_P2_R1077_U371, new_P2_R1077_U372,
    new_P2_R1077_U373, new_P2_R1077_U374, new_P2_R1077_U375,
    new_P2_R1077_U376, new_P2_R1077_U377, new_P2_R1077_U378,
    new_P2_R1077_U379, new_P2_R1077_U380, new_P2_R1077_U381,
    new_P2_R1077_U382, new_P2_R1077_U383, new_P2_R1077_U384,
    new_P2_R1077_U385, new_P2_R1077_U386, new_P2_R1077_U387,
    new_P2_R1077_U388, new_P2_R1077_U389, new_P2_R1077_U390,
    new_P2_R1077_U391, new_P2_R1077_U392, new_P2_R1077_U393,
    new_P2_R1077_U394, new_P2_R1077_U395, new_P2_R1077_U396,
    new_P2_R1077_U397, new_P2_R1077_U398, new_P2_R1077_U399,
    new_P2_R1077_U400, new_P2_R1077_U401, new_P2_R1077_U402,
    new_P2_R1077_U403, new_P2_R1077_U404, new_P2_R1077_U405,
    new_P2_R1077_U406, new_P2_R1077_U407, new_P2_R1077_U408,
    new_P2_R1077_U409, new_P2_R1077_U410, new_P2_R1077_U411,
    new_P2_R1077_U412, new_P2_R1077_U413, new_P2_R1077_U414,
    new_P2_R1077_U415, new_P2_R1077_U416, new_P2_R1077_U417,
    new_P2_R1077_U418, new_P2_R1077_U419, new_P2_R1077_U420,
    new_P2_R1077_U421, new_P2_R1077_U422, new_P2_R1077_U423,
    new_P2_R1077_U424, new_P2_R1077_U425, new_P2_R1077_U426,
    new_P2_R1077_U427, new_P2_R1077_U428, new_P2_R1077_U429,
    new_P2_R1077_U430, new_P2_R1077_U431, new_P2_R1077_U432,
    new_P2_R1077_U433, new_P2_R1077_U434, new_P2_R1077_U435,
    new_P2_R1077_U436, new_P2_R1077_U437, new_P2_R1077_U438,
    new_P2_R1077_U439, new_P2_R1077_U440, new_P2_R1077_U441,
    new_P2_R1077_U442, new_P2_R1077_U443, new_P2_R1077_U444,
    new_P2_R1077_U445, new_P2_R1077_U446, new_P2_R1077_U447,
    new_P2_R1077_U448, new_P2_R1077_U449, new_P2_R1077_U450,
    new_P2_R1077_U451, new_P2_R1077_U452, new_P2_R1077_U453,
    new_P2_R1077_U454, new_P2_R1077_U455, new_P2_R1077_U456,
    new_P2_R1077_U457, new_P2_R1077_U458, new_P2_R1077_U459,
    new_P2_R1077_U460, new_P2_R1077_U461, new_P2_R1077_U462,
    new_P2_R1077_U463, new_P2_R1077_U464, new_P2_R1077_U465,
    new_P2_R1077_U466, new_P2_R1077_U467, new_P2_R1077_U468,
    new_P2_R1077_U469, new_P2_R1077_U470, new_P2_R1077_U471,
    new_P2_R1077_U472, new_P2_R1077_U473, new_P2_R1077_U474,
    new_P2_R1077_U475, new_P2_R1077_U476, new_P2_R1077_U477,
    new_P2_R1077_U478, new_P2_R1077_U479, new_P2_R1077_U480,
    new_P2_R1077_U481, new_P2_R1077_U482, new_P2_R1077_U483,
    new_P2_R1077_U484, new_P2_R1077_U485, new_P2_R1077_U486,
    new_P2_R1077_U487, new_P2_R1077_U488, new_P2_R1077_U489,
    new_P2_R1077_U490, new_P2_R1077_U491, new_P2_R1077_U492,
    new_P2_R1077_U493, new_P2_R1077_U494, new_P2_R1077_U495,
    new_P2_R1077_U496, new_P2_R1077_U497, new_P2_R1077_U498,
    new_P2_R1077_U499, new_P2_R1077_U500, new_P2_R1077_U501,
    new_P2_R1077_U502, new_P2_R1077_U503, new_P2_R1077_U504,
    new_P2_R1143_U4, new_P2_R1143_U5, new_P2_R1143_U6, new_P2_R1143_U7,
    new_P2_R1143_U8, new_P2_R1143_U9, new_P2_R1143_U10, new_P2_R1143_U11,
    new_P2_R1143_U12, new_P2_R1143_U13, new_P2_R1143_U14, new_P2_R1143_U15,
    new_P2_R1143_U16, new_P2_R1143_U17, new_P2_R1143_U18, new_P2_R1143_U19,
    new_P2_R1143_U20, new_P2_R1143_U21, new_P2_R1143_U22, new_P2_R1143_U23,
    new_P2_R1143_U24, new_P2_R1143_U25, new_P2_R1143_U26, new_P2_R1143_U27,
    new_P2_R1143_U28, new_P2_R1143_U29, new_P2_R1143_U30, new_P2_R1143_U31,
    new_P2_R1143_U32, new_P2_R1143_U33, new_P2_R1143_U34, new_P2_R1143_U35,
    new_P2_R1143_U36, new_P2_R1143_U37, new_P2_R1143_U38, new_P2_R1143_U39,
    new_P2_R1143_U40, new_P2_R1143_U41, new_P2_R1143_U42, new_P2_R1143_U43,
    new_P2_R1143_U44, new_P2_R1143_U45, new_P2_R1143_U46, new_P2_R1143_U47,
    new_P2_R1143_U48, new_P2_R1143_U49, new_P2_R1143_U50, new_P2_R1143_U51,
    new_P2_R1143_U52, new_P2_R1143_U53, new_P2_R1143_U54, new_P2_R1143_U55,
    new_P2_R1143_U56, new_P2_R1143_U57, new_P2_R1143_U58, new_P2_R1143_U59,
    new_P2_R1143_U60, new_P2_R1143_U61, new_P2_R1143_U62, new_P2_R1143_U63,
    new_P2_R1143_U64, new_P2_R1143_U65, new_P2_R1143_U66, new_P2_R1143_U67,
    new_P2_R1143_U68, new_P2_R1143_U69, new_P2_R1143_U70, new_P2_R1143_U71,
    new_P2_R1143_U72, new_P2_R1143_U73, new_P2_R1143_U74, new_P2_R1143_U75,
    new_P2_R1143_U76, new_P2_R1143_U77, new_P2_R1143_U78, new_P2_R1143_U79,
    new_P2_R1143_U80, new_P2_R1143_U81, new_P2_R1143_U82, new_P2_R1143_U83,
    new_P2_R1143_U84, new_P2_R1143_U85, new_P2_R1143_U86, new_P2_R1143_U87,
    new_P2_R1143_U88, new_P2_R1143_U89, new_P2_R1143_U90, new_P2_R1143_U91,
    new_P2_R1143_U92, new_P2_R1143_U93, new_P2_R1143_U94, new_P2_R1143_U95,
    new_P2_R1143_U96, new_P2_R1143_U97, new_P2_R1143_U98, new_P2_R1143_U99,
    new_P2_R1143_U100, new_P2_R1143_U101, new_P2_R1143_U102,
    new_P2_R1143_U103, new_P2_R1143_U104, new_P2_R1143_U105,
    new_P2_R1143_U106, new_P2_R1143_U107, new_P2_R1143_U108,
    new_P2_R1143_U109, new_P2_R1143_U110, new_P2_R1143_U111,
    new_P2_R1143_U112, new_P2_R1143_U113, new_P2_R1143_U114,
    new_P2_R1143_U115, new_P2_R1143_U116, new_P2_R1143_U117,
    new_P2_R1143_U118, new_P2_R1143_U119, new_P2_R1143_U120,
    new_P2_R1143_U121, new_P2_R1143_U122, new_P2_R1143_U123,
    new_P2_R1143_U124, new_P2_R1143_U125, new_P2_R1143_U126,
    new_P2_R1143_U127, new_P2_R1143_U128, new_P2_R1143_U129,
    new_P2_R1143_U130, new_P2_R1143_U131, new_P2_R1143_U132,
    new_P2_R1143_U133, new_P2_R1143_U134, new_P2_R1143_U135,
    new_P2_R1143_U136, new_P2_R1143_U137, new_P2_R1143_U138,
    new_P2_R1143_U139, new_P2_R1143_U140, new_P2_R1143_U141,
    new_P2_R1143_U142, new_P2_R1143_U143, new_P2_R1143_U144,
    new_P2_R1143_U145, new_P2_R1143_U146, new_P2_R1143_U147,
    new_P2_R1143_U148, new_P2_R1143_U149, new_P2_R1143_U150,
    new_P2_R1143_U151, new_P2_R1143_U152, new_P2_R1143_U153,
    new_P2_R1143_U154, new_P2_R1143_U155, new_P2_R1143_U156,
    new_P2_R1143_U157, new_P2_R1143_U158, new_P2_R1143_U159,
    new_P2_R1143_U160, new_P2_R1143_U161, new_P2_R1143_U162,
    new_P2_R1143_U163, new_P2_R1143_U164, new_P2_R1143_U165,
    new_P2_R1143_U166, new_P2_R1143_U167, new_P2_R1143_U168,
    new_P2_R1143_U169, new_P2_R1143_U170, new_P2_R1143_U171,
    new_P2_R1143_U172, new_P2_R1143_U173, new_P2_R1143_U174,
    new_P2_R1143_U175, new_P2_R1143_U176, new_P2_R1143_U177,
    new_P2_R1143_U178, new_P2_R1143_U179, new_P2_R1143_U180,
    new_P2_R1143_U181, new_P2_R1143_U182, new_P2_R1143_U183,
    new_P2_R1143_U184, new_P2_R1143_U185, new_P2_R1143_U186,
    new_P2_R1143_U187, new_P2_R1143_U188, new_P2_R1143_U189,
    new_P2_R1143_U190, new_P2_R1143_U191, new_P2_R1143_U192,
    new_P2_R1143_U193, new_P2_R1143_U194, new_P2_R1143_U195,
    new_P2_R1143_U196, new_P2_R1143_U197, new_P2_R1143_U198,
    new_P2_R1143_U199, new_P2_R1143_U200, new_P2_R1143_U201,
    new_P2_R1143_U202, new_P2_R1143_U203, new_P2_R1143_U204,
    new_P2_R1143_U205, new_P2_R1143_U206, new_P2_R1143_U207,
    new_P2_R1143_U208, new_P2_R1143_U209, new_P2_R1143_U210,
    new_P2_R1143_U211, new_P2_R1143_U212, new_P2_R1143_U213,
    new_P2_R1143_U214, new_P2_R1143_U215, new_P2_R1143_U216,
    new_P2_R1143_U217, new_P2_R1143_U218, new_P2_R1143_U219,
    new_P2_R1143_U220, new_P2_R1143_U221, new_P2_R1143_U222,
    new_P2_R1143_U223, new_P2_R1143_U224, new_P2_R1143_U225,
    new_P2_R1143_U226, new_P2_R1143_U227, new_P2_R1143_U228,
    new_P2_R1143_U229, new_P2_R1143_U230, new_P2_R1143_U231,
    new_P2_R1143_U232, new_P2_R1143_U233, new_P2_R1143_U234,
    new_P2_R1143_U235, new_P2_R1143_U236, new_P2_R1143_U237,
    new_P2_R1143_U238, new_P2_R1143_U239, new_P2_R1143_U240,
    new_P2_R1143_U241, new_P2_R1143_U242, new_P2_R1143_U243,
    new_P2_R1143_U244, new_P2_R1143_U245, new_P2_R1143_U246,
    new_P2_R1143_U247, new_P2_R1143_U248, new_P2_R1143_U249,
    new_P2_R1143_U250, new_P2_R1143_U251, new_P2_R1143_U252,
    new_P2_R1143_U253, new_P2_R1143_U254, new_P2_R1143_U255,
    new_P2_R1143_U256, new_P2_R1143_U257, new_P2_R1143_U258,
    new_P2_R1143_U259, new_P2_R1143_U260, new_P2_R1143_U261,
    new_P2_R1143_U262, new_P2_R1143_U263, new_P2_R1143_U264,
    new_P2_R1143_U265, new_P2_R1143_U266, new_P2_R1143_U267,
    new_P2_R1143_U268, new_P2_R1143_U269, new_P2_R1143_U270,
    new_P2_R1143_U271, new_P2_R1143_U272, new_P2_R1143_U273,
    new_P2_R1143_U274, new_P2_R1143_U275, new_P2_R1143_U276,
    new_P2_R1143_U277, new_P2_R1143_U278, new_P2_R1143_U279,
    new_P2_R1143_U280, new_P2_R1143_U281, new_P2_R1143_U282,
    new_P2_R1143_U283, new_P2_R1143_U284, new_P2_R1143_U285,
    new_P2_R1143_U286, new_P2_R1143_U287, new_P2_R1143_U288,
    new_P2_R1143_U289, new_P2_R1143_U290, new_P2_R1143_U291,
    new_P2_R1143_U292, new_P2_R1143_U293, new_P2_R1143_U294,
    new_P2_R1143_U295, new_P2_R1143_U296, new_P2_R1143_U297,
    new_P2_R1143_U298, new_P2_R1143_U299, new_P2_R1143_U300,
    new_P2_R1143_U301, new_P2_R1143_U302, new_P2_R1143_U303,
    new_P2_R1143_U304, new_P2_R1143_U305, new_P2_R1143_U306,
    new_P2_R1143_U307, new_P2_R1143_U308, new_P2_R1143_U309,
    new_P2_R1143_U310, new_P2_R1143_U311, new_P2_R1143_U312,
    new_P2_R1143_U313, new_P2_R1143_U314, new_P2_R1143_U315,
    new_P2_R1143_U316, new_P2_R1143_U317, new_P2_R1143_U318,
    new_P2_R1143_U319, new_P2_R1143_U320, new_P2_R1143_U321,
    new_P2_R1143_U322, new_P2_R1143_U323, new_P2_R1143_U324,
    new_P2_R1143_U325, new_P2_R1143_U326, new_P2_R1143_U327,
    new_P2_R1143_U328, new_P2_R1143_U329, new_P2_R1143_U330,
    new_P2_R1143_U331, new_P2_R1143_U332, new_P2_R1143_U333,
    new_P2_R1143_U334, new_P2_R1143_U335, new_P2_R1143_U336,
    new_P2_R1143_U337, new_P2_R1143_U338, new_P2_R1143_U339,
    new_P2_R1143_U340, new_P2_R1143_U341, new_P2_R1143_U342,
    new_P2_R1143_U343, new_P2_R1143_U344, new_P2_R1143_U345,
    new_P2_R1143_U346, new_P2_R1143_U347, new_P2_R1143_U348,
    new_P2_R1143_U349, new_P2_R1143_U350, new_P2_R1143_U351,
    new_P2_R1143_U352, new_P2_R1143_U353, new_P2_R1143_U354,
    new_P2_R1143_U355, new_P2_R1143_U356, new_P2_R1143_U357,
    new_P2_R1143_U358, new_P2_R1143_U359, new_P2_R1143_U360,
    new_P2_R1143_U361, new_P2_R1143_U362, new_P2_R1143_U363,
    new_P2_R1143_U364, new_P2_R1143_U365, new_P2_R1143_U366,
    new_P2_R1143_U367, new_P2_R1143_U368, new_P2_R1143_U369,
    new_P2_R1143_U370, new_P2_R1143_U371, new_P2_R1143_U372,
    new_P2_R1143_U373, new_P2_R1143_U374, new_P2_R1143_U375,
    new_P2_R1143_U376, new_P2_R1143_U377, new_P2_R1143_U378,
    new_P2_R1143_U379, new_P2_R1143_U380, new_P2_R1143_U381,
    new_P2_R1143_U382, new_P2_R1143_U383, new_P2_R1143_U384,
    new_P2_R1143_U385, new_P2_R1143_U386, new_P2_R1143_U387,
    new_P2_R1143_U388, new_P2_R1143_U389, new_P2_R1143_U390,
    new_P2_R1143_U391, new_P2_R1143_U392, new_P2_R1143_U393,
    new_P2_R1143_U394, new_P2_R1143_U395, new_P2_R1143_U396,
    new_P2_R1143_U397, new_P2_R1143_U398, new_P2_R1143_U399,
    new_P2_R1143_U400, new_P2_R1143_U401, new_P2_R1143_U402,
    new_P2_R1143_U403, new_P2_R1143_U404, new_P2_R1143_U405,
    new_P2_R1143_U406, new_P2_R1143_U407, new_P2_R1143_U408,
    new_P2_R1143_U409, new_P2_R1143_U410, new_P2_R1143_U411,
    new_P2_R1143_U412, new_P2_R1143_U413, new_P2_R1143_U414,
    new_P2_R1143_U415, new_P2_R1143_U416, new_P2_R1143_U417,
    new_P2_R1143_U418, new_P2_R1143_U419, new_P2_R1143_U420,
    new_P2_R1143_U421, new_P2_R1143_U422, new_P2_R1143_U423,
    new_P2_R1143_U424, new_P2_R1143_U425, new_P2_R1143_U426,
    new_P2_R1143_U427, new_P2_R1143_U428, new_P2_R1143_U429,
    new_P2_R1143_U430, new_P2_R1143_U431, new_P2_R1143_U432,
    new_P2_R1143_U433, new_P2_R1143_U434, new_P2_R1143_U435,
    new_P2_R1143_U436, new_P2_R1143_U437, new_P2_R1143_U438,
    new_P2_R1143_U439, new_P2_R1143_U440, new_P2_R1143_U441,
    new_P2_R1143_U442, new_P2_R1143_U443, new_P2_R1143_U444,
    new_P2_R1143_U445, new_P2_R1143_U446, new_P2_R1143_U447,
    new_P2_R1143_U448, new_P2_R1143_U449, new_P2_R1143_U450,
    new_P2_R1143_U451, new_P2_R1143_U452, new_P2_R1143_U453,
    new_P2_R1143_U454, new_P2_R1143_U455, new_P2_R1143_U456,
    new_P2_R1143_U457, new_P2_R1143_U458, new_P2_R1143_U459,
    new_P2_R1143_U460, new_P2_R1143_U461, new_P2_R1143_U462,
    new_P2_R1143_U463, new_P2_R1143_U464, new_P2_R1143_U465,
    new_P2_R1143_U466, new_P2_R1143_U467, new_P2_R1143_U468,
    new_P2_R1143_U469, new_P2_R1143_U470, new_P2_R1143_U471,
    new_P2_R1143_U472, new_P2_R1143_U473, new_P2_R1143_U474,
    new_P2_R1143_U475, new_P2_R1143_U476, new_P2_R1143_U477,
    new_P2_R1143_U478, new_P2_R1143_U479, new_P2_R1143_U480,
    new_P2_R1143_U481, new_P2_R1143_U482, new_P2_R1143_U483,
    new_P2_R1143_U484, new_P2_R1143_U485, new_P2_R1143_U486,
    new_P2_R1143_U487, new_P2_R1143_U488, new_P2_R1143_U489,
    new_P2_R1143_U490, new_P2_R1143_U491, new_P2_R1143_U492,
    new_P2_R1143_U493, new_P2_R1143_U494, new_P2_R1143_U495,
    new_P2_R1143_U496, new_P2_R1143_U497, new_P2_R1143_U498,
    new_P2_R1143_U499, new_P2_R1143_U500, new_P2_R1143_U501,
    new_P2_R1143_U502, new_P2_R1143_U503, new_P2_R1143_U504,
    new_P2_R1158_U4, new_P2_R1158_U5, new_P2_R1158_U6, new_P2_R1158_U7,
    new_P2_R1158_U8, new_P2_R1158_U9, new_P2_R1158_U10, new_P2_R1158_U11,
    new_P2_R1158_U12, new_P2_R1158_U13, new_P2_R1158_U14, new_P2_R1158_U15,
    new_P2_R1158_U16, new_P2_R1158_U17, new_P2_R1158_U18, new_P2_R1158_U19,
    new_P2_R1158_U20, new_P2_R1158_U21, new_P2_R1158_U22, new_P2_R1158_U23,
    new_P2_R1158_U24, new_P2_R1158_U25, new_P2_R1158_U26, new_P2_R1158_U27,
    new_P2_R1158_U28, new_P2_R1158_U29, new_P2_R1158_U30, new_P2_R1158_U31,
    new_P2_R1158_U32, new_P2_R1158_U33, new_P2_R1158_U34, new_P2_R1158_U35,
    new_P2_R1158_U36, new_P2_R1158_U37, new_P2_R1158_U38, new_P2_R1158_U39,
    new_P2_R1158_U40, new_P2_R1158_U41, new_P2_R1158_U42, new_P2_R1158_U43,
    new_P2_R1158_U44, new_P2_R1158_U45, new_P2_R1158_U46, new_P2_R1158_U47,
    new_P2_R1158_U48, new_P2_R1158_U49, new_P2_R1158_U50, new_P2_R1158_U51,
    new_P2_R1158_U52, new_P2_R1158_U53, new_P2_R1158_U54, new_P2_R1158_U55,
    new_P2_R1158_U56, new_P2_R1158_U57, new_P2_R1158_U58, new_P2_R1158_U59,
    new_P2_R1158_U60, new_P2_R1158_U61, new_P2_R1158_U62, new_P2_R1158_U63,
    new_P2_R1158_U64, new_P2_R1158_U65, new_P2_R1158_U66, new_P2_R1158_U67,
    new_P2_R1158_U68, new_P2_R1158_U69, new_P2_R1158_U70, new_P2_R1158_U71,
    new_P2_R1158_U72, new_P2_R1158_U73, new_P2_R1158_U74, new_P2_R1158_U75,
    new_P2_R1158_U76, new_P2_R1158_U77, new_P2_R1158_U78, new_P2_R1158_U79,
    new_P2_R1158_U80, new_P2_R1158_U81, new_P2_R1158_U82, new_P2_R1158_U83,
    new_P2_R1158_U84, new_P2_R1158_U85, new_P2_R1158_U86, new_P2_R1158_U87,
    new_P2_R1158_U88, new_P2_R1158_U89, new_P2_R1158_U90, new_P2_R1158_U91,
    new_P2_R1158_U92, new_P2_R1158_U93, new_P2_R1158_U94, new_P2_R1158_U95,
    new_P2_R1158_U96, new_P2_R1158_U97, new_P2_R1158_U98, new_P2_R1158_U99,
    new_P2_R1158_U100, new_P2_R1158_U101, new_P2_R1158_U102,
    new_P2_R1158_U103, new_P2_R1158_U104, new_P2_R1158_U105,
    new_P2_R1158_U106, new_P2_R1158_U107, new_P2_R1158_U108,
    new_P2_R1158_U109, new_P2_R1158_U110, new_P2_R1158_U111,
    new_P2_R1158_U112, new_P2_R1158_U113, new_P2_R1158_U114,
    new_P2_R1158_U115, new_P2_R1158_U116, new_P2_R1158_U117,
    new_P2_R1158_U118, new_P2_R1158_U119, new_P2_R1158_U120,
    new_P2_R1158_U121, new_P2_R1158_U122, new_P2_R1158_U123,
    new_P2_R1158_U124, new_P2_R1158_U125, new_P2_R1158_U126,
    new_P2_R1158_U127, new_P2_R1158_U128, new_P2_R1158_U129,
    new_P2_R1158_U130, new_P2_R1158_U131, new_P2_R1158_U132,
    new_P2_R1158_U133, new_P2_R1158_U134, new_P2_R1158_U135,
    new_P2_R1158_U136, new_P2_R1158_U137, new_P2_R1158_U138,
    new_P2_R1158_U139, new_P2_R1158_U140, new_P2_R1158_U141,
    new_P2_R1158_U142, new_P2_R1158_U143, new_P2_R1158_U144,
    new_P2_R1158_U145, new_P2_R1158_U146, new_P2_R1158_U147,
    new_P2_R1158_U148, new_P2_R1158_U149, new_P2_R1158_U150,
    new_P2_R1158_U151, new_P2_R1158_U152, new_P2_R1158_U153,
    new_P2_R1158_U154, new_P2_R1158_U155, new_P2_R1158_U156,
    new_P2_R1158_U157, new_P2_R1158_U158, new_P2_R1158_U159,
    new_P2_R1158_U160, new_P2_R1158_U161, new_P2_R1158_U162,
    new_P2_R1158_U163, new_P2_R1158_U164, new_P2_R1158_U165,
    new_P2_R1158_U166, new_P2_R1158_U167, new_P2_R1158_U168,
    new_P2_R1158_U169, new_P2_R1158_U170, new_P2_R1158_U171,
    new_P2_R1158_U172, new_P2_R1158_U173, new_P2_R1158_U174,
    new_P2_R1158_U175, new_P2_R1158_U176, new_P2_R1158_U177,
    new_P2_R1158_U178, new_P2_R1158_U179, new_P2_R1158_U180,
    new_P2_R1158_U181, new_P2_R1158_U182, new_P2_R1158_U183,
    new_P2_R1158_U184, new_P2_R1158_U185, new_P2_R1158_U186,
    new_P2_R1158_U187, new_P2_R1158_U188, new_P2_R1158_U189,
    new_P2_R1158_U190, new_P2_R1158_U191, new_P2_R1158_U192,
    new_P2_R1158_U193, new_P2_R1158_U194, new_P2_R1158_U195,
    new_P2_R1158_U196, new_P2_R1158_U197, new_P2_R1158_U198,
    new_P2_R1158_U199, new_P2_R1158_U200, new_P2_R1158_U201,
    new_P2_R1158_U202, new_P2_R1158_U203, new_P2_R1158_U204,
    new_P2_R1158_U205, new_P2_R1158_U206, new_P2_R1158_U207,
    new_P2_R1158_U208, new_P2_R1158_U209, new_P2_R1158_U210,
    new_P2_R1158_U211, new_P2_R1158_U212, new_P2_R1158_U213,
    new_P2_R1158_U214, new_P2_R1158_U215, new_P2_R1158_U216,
    new_P2_R1158_U217, new_P2_R1158_U218, new_P2_R1158_U219,
    new_P2_R1158_U220, new_P2_R1158_U221, new_P2_R1158_U222,
    new_P2_R1158_U223, new_P2_R1158_U224, new_P2_R1158_U225,
    new_P2_R1158_U226, new_P2_R1158_U227, new_P2_R1158_U228,
    new_P2_R1158_U229, new_P2_R1158_U230, new_P2_R1158_U231,
    new_P2_R1158_U232, new_P2_R1158_U233, new_P2_R1158_U234,
    new_P2_R1158_U235, new_P2_R1158_U236, new_P2_R1158_U237,
    new_P2_R1158_U238, new_P2_R1158_U239, new_P2_R1158_U240,
    new_P2_R1158_U241, new_P2_R1158_U242, new_P2_R1158_U243,
    new_P2_R1158_U244, new_P2_R1158_U245, new_P2_R1158_U246,
    new_P2_R1158_U247, new_P2_R1158_U248, new_P2_R1158_U249,
    new_P2_R1158_U250, new_P2_R1158_U251, new_P2_R1158_U252,
    new_P2_R1158_U253, new_P2_R1158_U254, new_P2_R1158_U255,
    new_P2_R1158_U256, new_P2_R1158_U257, new_P2_R1158_U258,
    new_P2_R1158_U259, new_P2_R1158_U260, new_P2_R1158_U261,
    new_P2_R1158_U262, new_P2_R1158_U263, new_P2_R1158_U264,
    new_P2_R1158_U265, new_P2_R1158_U266, new_P2_R1158_U267,
    new_P2_R1158_U268, new_P2_R1158_U269, new_P2_R1158_U270,
    new_P2_R1158_U271, new_P2_R1158_U272, new_P2_R1158_U273,
    new_P2_R1158_U274, new_P2_R1158_U275, new_P2_R1158_U276,
    new_P2_R1158_U277, new_P2_R1158_U278, new_P2_R1158_U279,
    new_P2_R1158_U280, new_P2_R1158_U281, new_P2_R1158_U282,
    new_P2_R1158_U283, new_P2_R1158_U284, new_P2_R1158_U285,
    new_P2_R1158_U286, new_P2_R1158_U287, new_P2_R1158_U288,
    new_P2_R1158_U289, new_P2_R1158_U290, new_P2_R1158_U291,
    new_P2_R1158_U292, new_P2_R1158_U293, new_P2_R1158_U294,
    new_P2_R1158_U295, new_P2_R1158_U296, new_P2_R1158_U297,
    new_P2_R1158_U298, new_P2_R1158_U299, new_P2_R1158_U300,
    new_P2_R1158_U301, new_P2_R1158_U302, new_P2_R1158_U303,
    new_P2_R1158_U304, new_P2_R1158_U305, new_P2_R1158_U306,
    new_P2_R1158_U307, new_P2_R1158_U308, new_P2_R1158_U309,
    new_P2_R1158_U310, new_P2_R1158_U311, new_P2_R1158_U312,
    new_P2_R1158_U313, new_P2_R1158_U314, new_P2_R1158_U315,
    new_P2_R1158_U316, new_P2_R1158_U317, new_P2_R1158_U318,
    new_P2_R1158_U319, new_P2_R1158_U320, new_P2_R1158_U321,
    new_P2_R1158_U322, new_P2_R1158_U323, new_P2_R1158_U324,
    new_P2_R1158_U325, new_P2_R1158_U326, new_P2_R1158_U327,
    new_P2_R1158_U328, new_P2_R1158_U329, new_P2_R1158_U330,
    new_P2_R1158_U331, new_P2_R1158_U332, new_P2_R1158_U333,
    new_P2_R1158_U334, new_P2_R1158_U335, new_P2_R1158_U336,
    new_P2_R1158_U337, new_P2_R1158_U338, new_P2_R1158_U339,
    new_P2_R1158_U340, new_P2_R1158_U341, new_P2_R1158_U342,
    new_P2_R1158_U343, new_P2_R1158_U344, new_P2_R1158_U345,
    new_P2_R1158_U346, new_P2_R1158_U347, new_P2_R1158_U348,
    new_P2_R1158_U349, new_P2_R1158_U350, new_P2_R1158_U351,
    new_P2_R1158_U352, new_P2_R1158_U353, new_P2_R1158_U354,
    new_P2_R1158_U355, new_P2_R1158_U356, new_P2_R1158_U357,
    new_P2_R1158_U358, new_P2_R1158_U359, new_P2_R1158_U360,
    new_P2_R1158_U361, new_P2_R1158_U362, new_P2_R1158_U363,
    new_P2_R1158_U364, new_P2_R1158_U365, new_P2_R1158_U366,
    new_P2_R1158_U367, new_P2_R1158_U368, new_P2_R1158_U369,
    new_P2_R1158_U370, new_P2_R1158_U371, new_P2_R1158_U372,
    new_P2_R1158_U373, new_P2_R1158_U374, new_P2_R1158_U375,
    new_P2_R1158_U376, new_P2_R1158_U377, new_P2_R1158_U378,
    new_P2_R1158_U379, new_P2_R1158_U380, new_P2_R1158_U381,
    new_P2_R1158_U382, new_P2_R1158_U383, new_P2_R1158_U384,
    new_P2_R1158_U385, new_P2_R1158_U386, new_P2_R1158_U387,
    new_P2_R1158_U388, new_P2_R1158_U389, new_P2_R1158_U390,
    new_P2_R1158_U391, new_P2_R1158_U392, new_P2_R1158_U393,
    new_P2_R1158_U394, new_P2_R1158_U395, new_P2_R1158_U396,
    new_P2_R1158_U397, new_P2_R1158_U398, new_P2_R1158_U399,
    new_P2_R1158_U400, new_P2_R1158_U401, new_P2_R1158_U402,
    new_P2_R1158_U403, new_P2_R1158_U404, new_P2_R1158_U405,
    new_P2_R1158_U406, new_P2_R1158_U407, new_P2_R1158_U408,
    new_P2_R1158_U409, new_P2_R1158_U410, new_P2_R1158_U411,
    new_P2_R1158_U412, new_P2_R1158_U413, new_P2_R1158_U414,
    new_P2_R1158_U415, new_P2_R1158_U416, new_P2_R1158_U417,
    new_P2_R1158_U418, new_P2_R1158_U419, new_P2_R1158_U420,
    new_P2_R1158_U421, new_P2_R1158_U422, new_P2_R1158_U423,
    new_P2_R1158_U424, new_P2_R1158_U425, new_P2_R1158_U426,
    new_P2_R1158_U427, new_P2_R1158_U428, new_P2_R1158_U429,
    new_P2_R1158_U430, new_P2_R1158_U431, new_P2_R1158_U432,
    new_P2_R1158_U433, new_P2_R1158_U434, new_P2_R1158_U435,
    new_P2_R1158_U436, new_P2_R1158_U437, new_P2_R1158_U438,
    new_P2_R1158_U439, new_P2_R1158_U440, new_P2_R1158_U441,
    new_P2_R1158_U442, new_P2_R1158_U443, new_P2_R1158_U444,
    new_P2_R1158_U445, new_P2_R1158_U446, new_P2_R1158_U447,
    new_P2_R1158_U448, new_P2_R1158_U449, new_P2_R1158_U450,
    new_P2_R1158_U451, new_P2_R1158_U452, new_P2_R1158_U453,
    new_P2_R1158_U454, new_P2_R1158_U455, new_P2_R1158_U456,
    new_P2_R1158_U457, new_P2_R1158_U458, new_P2_R1158_U459,
    new_P2_R1158_U460, new_P2_R1158_U461, new_P2_R1158_U462,
    new_P2_R1158_U463, new_P2_R1158_U464, new_P2_R1158_U465,
    new_P2_R1158_U466, new_P2_R1158_U467, new_P2_R1158_U468,
    new_P2_R1158_U469, new_P2_R1158_U470, new_P2_R1158_U471,
    new_P2_R1158_U472, new_P2_R1158_U473, new_P2_R1158_U474,
    new_P2_R1158_U475, new_P2_R1158_U476, new_P2_R1158_U477,
    new_P2_R1158_U478, new_P2_R1158_U479, new_P2_R1158_U480,
    new_P2_R1158_U481, new_P2_R1158_U482, new_P2_R1158_U483,
    new_P2_R1158_U484, new_P2_R1158_U485, new_P2_R1158_U486,
    new_P2_R1158_U487, new_P2_R1158_U488, new_P2_R1158_U489,
    new_P2_R1158_U490, new_P2_R1158_U491, new_P2_R1158_U492,
    new_P2_R1158_U493, new_P2_R1158_U494, new_P2_R1158_U495,
    new_P2_R1158_U496, new_P2_R1158_U497, new_P2_R1158_U498,
    new_P2_R1158_U499, new_P2_R1158_U500, new_P2_R1158_U501,
    new_P2_R1158_U502, new_P2_R1158_U503, new_P2_R1158_U504,
    new_P2_R1158_U505, new_P2_R1158_U506, new_P2_R1158_U507,
    new_P2_R1158_U508, new_P2_R1158_U509, new_P2_R1158_U510,
    new_P2_R1158_U511, new_P2_R1158_U512, new_P2_R1158_U513,
    new_P2_R1158_U514, new_P2_R1158_U515, new_P2_R1158_U516,
    new_P2_R1158_U517, new_P2_R1158_U518, new_P2_R1158_U519,
    new_P2_R1158_U520, new_P2_R1158_U521, new_P2_R1158_U522,
    new_P2_R1158_U523, new_P2_R1158_U524, new_P2_R1158_U525,
    new_P2_R1158_U526, new_P2_R1158_U527, new_P2_R1158_U528,
    new_P2_R1158_U529, new_P2_R1158_U530, new_P2_R1158_U531,
    new_P2_R1158_U532, new_P2_R1158_U533, new_P2_R1158_U534,
    new_P2_R1158_U535, new_P2_R1158_U536, new_P2_R1158_U537,
    new_P2_R1158_U538, new_P2_R1158_U539, new_P2_R1158_U540,
    new_P2_R1158_U541, new_P2_R1158_U542, new_P2_R1158_U543,
    new_P2_R1158_U544, new_P2_R1158_U545, new_P2_R1158_U546,
    new_P2_R1158_U547, new_P2_R1158_U548, new_P2_R1158_U549,
    new_P2_R1158_U550, new_P2_R1158_U551, new_P2_R1158_U552,
    new_P2_R1158_U553, new_P2_R1158_U554, new_P2_R1158_U555,
    new_P2_R1158_U556, new_P2_R1158_U557, new_P2_R1158_U558,
    new_P2_R1158_U559, new_P2_R1158_U560, new_P2_R1158_U561,
    new_P2_R1158_U562, new_P2_R1158_U563, new_P2_R1158_U564,
    new_P2_R1158_U565, new_P2_R1158_U566, new_P2_R1158_U567,
    new_P2_R1158_U568, new_P2_R1158_U569, new_P2_R1158_U570,
    new_P2_R1158_U571, new_P2_R1158_U572, new_P2_R1158_U573,
    new_P2_R1158_U574, new_P2_R1158_U575, new_P2_R1158_U576,
    new_P2_R1158_U577, new_P2_R1158_U578, new_P2_R1158_U579,
    new_P2_R1158_U580, new_P2_R1158_U581, new_P2_R1158_U582,
    new_P2_R1158_U583, new_P2_R1158_U584, new_P2_R1158_U585,
    new_P2_R1158_U586, new_P2_R1158_U587, new_P2_R1158_U588,
    new_P2_R1158_U589, new_P2_R1158_U590, new_P2_R1158_U591,
    new_P2_R1158_U592, new_P2_R1158_U593, new_P2_R1158_U594,
    new_P2_R1158_U595, new_P2_R1158_U596, new_P2_R1158_U597,
    new_P2_R1158_U598, new_P2_R1158_U599, new_P2_R1158_U600,
    new_P2_R1158_U601, new_P2_R1158_U602, new_P2_R1158_U603,
    new_P2_R1158_U604, new_P2_R1158_U605, new_P2_R1158_U606,
    new_P2_R1158_U607, new_P2_R1158_U608, new_P2_R1158_U609,
    new_P2_R1158_U610, new_P2_R1158_U611, new_P2_R1158_U612,
    new_P2_R1158_U613, new_P2_R1158_U614, new_P2_R1158_U615,
    new_P2_R1158_U616, new_P2_R1158_U617, new_P2_R1158_U618,
    new_P2_R1158_U619, new_P2_R1158_U620, new_P2_R1158_U621,
    new_P2_R1158_U622, new_P2_R1158_U623, new_P2_R1158_U624,
    new_P2_R1158_U625, new_P2_R1158_U626, new_P2_R1158_U627,
    new_P2_R1158_U628, new_P2_R1158_U629, new_P2_R1158_U630,
    new_P2_R1158_U631, new_P2_R1158_U632, new_P2_R1158_U633,
    new_P2_R1158_U634, new_P2_R1131_U6, new_P2_R1131_U7, new_P2_R1131_U8,
    new_P2_R1131_U9, new_P2_R1131_U10, new_P2_R1131_U11, new_P2_R1131_U12,
    new_P2_R1131_U13, new_P2_R1131_U14, new_P2_R1131_U15, new_P2_R1131_U16,
    new_P2_R1131_U17, new_P2_R1131_U18, new_P2_R1131_U19, new_P2_R1131_U20,
    new_P2_R1131_U21, new_P2_R1131_U22, new_P2_R1131_U23, new_P2_R1131_U24,
    new_P2_R1131_U25, new_P2_R1131_U26, new_P2_R1131_U27, new_P2_R1131_U28,
    new_P2_R1131_U29, new_P2_R1131_U30, new_P2_R1131_U31, new_P2_R1131_U32,
    new_P2_R1131_U33, new_P2_R1131_U34, new_P2_R1131_U35, new_P2_R1131_U36,
    new_P2_R1131_U37, new_P2_R1131_U38, new_P2_R1131_U39, new_P2_R1131_U40,
    new_P2_R1131_U41, new_P2_R1131_U42, new_P2_R1131_U43, new_P2_R1131_U44,
    new_P2_R1131_U45, new_P2_R1131_U46, new_P2_R1131_U47, new_P2_R1131_U48,
    new_P2_R1131_U49, new_P2_R1131_U50, new_P2_R1131_U51, new_P2_R1131_U52,
    new_P2_R1131_U53, new_P2_R1131_U54, new_P2_R1131_U55, new_P2_R1131_U56,
    new_P2_R1131_U57, new_P2_R1131_U58, new_P2_R1131_U59, new_P2_R1131_U60,
    new_P2_R1131_U61, new_P2_R1131_U62, new_P2_R1131_U63, new_P2_R1131_U64,
    new_P2_R1131_U65, new_P2_R1131_U66, new_P2_R1131_U67, new_P2_R1131_U68,
    new_P2_R1131_U69, new_P2_R1131_U70, new_P2_R1131_U71, new_P2_R1131_U72,
    new_P2_R1131_U73, new_P2_R1131_U74, new_P2_R1131_U75, new_P2_R1131_U76,
    new_P2_R1131_U77, new_P2_R1131_U78, new_P2_R1131_U79, new_P2_R1131_U80,
    new_P2_R1131_U81, new_P2_R1131_U82, new_P2_R1131_U83, new_P2_R1131_U84,
    new_P2_R1131_U85, new_P2_R1131_U86, new_P2_R1131_U87, new_P2_R1131_U88,
    new_P2_R1131_U89, new_P2_R1131_U90, new_P2_R1131_U91, new_P2_R1131_U92,
    new_P2_R1131_U93, new_P2_R1131_U94, new_P2_R1131_U95, new_P2_R1131_U96,
    new_P2_R1131_U97, new_P2_R1131_U98, new_P2_R1131_U99,
    new_P2_R1131_U100, new_P2_R1131_U101, new_P2_R1131_U102,
    new_P2_R1131_U103, new_P2_R1131_U104, new_P2_R1131_U105,
    new_P2_R1131_U106, new_P2_R1131_U107, new_P2_R1131_U108,
    new_P2_R1131_U109, new_P2_R1131_U110, new_P2_R1131_U111,
    new_P2_R1131_U112, new_P2_R1131_U113, new_P2_R1131_U114,
    new_P2_R1131_U115, new_P2_R1131_U116, new_P2_R1131_U117,
    new_P2_R1131_U118, new_P2_R1131_U119, new_P2_R1131_U120,
    new_P2_R1131_U121, new_P2_R1131_U122, new_P2_R1131_U123,
    new_P2_R1131_U124, new_P2_R1131_U125, new_P2_R1131_U126,
    new_P2_R1131_U127, new_P2_R1131_U128, new_P2_R1131_U129,
    new_P2_R1131_U130, new_P2_R1131_U131, new_P2_R1131_U132,
    new_P2_R1131_U133, new_P2_R1131_U134, new_P2_R1131_U135,
    new_P2_R1131_U136, new_P2_R1131_U137, new_P2_R1131_U138,
    new_P2_R1131_U139, new_P2_R1131_U140, new_P2_R1131_U141,
    new_P2_R1131_U142, new_P2_R1131_U143, new_P2_R1131_U144,
    new_P2_R1131_U145, new_P2_R1131_U146, new_P2_R1131_U147,
    new_P2_R1131_U148, new_P2_R1131_U149, new_P2_R1131_U150,
    new_P2_R1131_U151, new_P2_R1131_U152, new_P2_R1131_U153,
    new_P2_R1131_U154, new_P2_R1131_U155, new_P2_R1131_U156,
    new_P2_R1131_U157, new_P2_R1131_U158, new_P2_R1131_U159,
    new_P2_R1131_U160, new_P2_R1131_U161, new_P2_R1131_U162,
    new_P2_R1131_U163, new_P2_R1131_U164, new_P2_R1131_U165,
    new_P2_R1131_U166, new_P2_R1131_U167, new_P2_R1131_U168,
    new_P2_R1131_U169, new_P2_R1131_U170, new_P2_R1131_U171,
    new_P2_R1131_U172, new_P2_R1131_U173, new_P2_R1131_U174,
    new_P2_R1131_U175, new_P2_R1131_U176, new_P2_R1131_U177,
    new_P2_R1131_U178, new_P2_R1131_U179, new_P2_R1131_U180,
    new_P2_R1131_U181, new_P2_R1131_U182, new_P2_R1131_U183,
    new_P2_R1131_U184, new_P2_R1131_U185, new_P2_R1131_U186,
    new_P2_R1131_U187, new_P2_R1131_U188, new_P2_R1131_U189,
    new_P2_R1131_U190, new_P2_R1131_U191, new_P2_R1131_U192,
    new_P2_R1131_U193, new_P2_R1131_U194, new_P2_R1131_U195,
    new_P2_R1131_U196, new_P2_R1131_U197, new_P2_R1131_U198,
    new_P2_R1131_U199, new_P2_R1131_U200, new_P2_R1131_U201,
    new_P2_R1131_U202, new_P2_R1131_U203, new_P2_R1131_U204,
    new_P2_R1131_U205, new_P2_R1131_U206, new_P2_R1131_U207,
    new_P2_R1131_U208, new_P2_R1131_U209, new_P2_R1131_U210,
    new_P2_R1131_U211, new_P2_R1131_U212, new_P2_R1131_U213,
    new_P2_R1131_U214, new_P2_R1131_U215, new_P2_R1131_U216,
    new_P2_R1131_U217, new_P2_R1131_U218, new_P2_R1131_U219,
    new_P2_R1131_U220, new_P2_R1131_U221, new_P2_R1131_U222,
    new_P2_R1131_U223, new_P2_R1131_U224, new_P2_R1131_U225,
    new_P2_R1131_U226, new_P2_R1131_U227, new_P2_R1131_U228,
    new_P2_R1131_U229, new_P2_R1131_U230, new_P2_R1131_U231,
    new_P2_R1131_U232, new_P2_R1131_U233, new_P2_R1131_U234,
    new_P2_R1131_U235, new_P2_R1131_U236, new_P2_R1131_U237,
    new_P2_R1131_U238, new_P2_R1131_U239, new_P2_R1131_U240,
    new_P2_R1131_U241, new_P2_R1131_U242, new_P2_R1131_U243,
    new_P2_R1131_U244, new_P2_R1131_U245, new_P2_R1131_U246,
    new_P2_R1131_U247, new_P2_R1131_U248, new_P2_R1131_U249,
    new_P2_R1131_U250, new_P2_R1131_U251, new_P2_R1131_U252,
    new_P2_R1131_U253, new_P2_R1131_U254, new_P2_R1131_U255,
    new_P2_R1131_U256, new_P2_R1131_U257, new_P2_R1131_U258,
    new_P2_R1131_U259, new_P2_R1131_U260, new_P2_R1131_U261,
    new_P2_R1131_U262, new_P2_R1131_U263, new_P2_R1131_U264,
    new_P2_R1131_U265, new_P2_R1131_U266, new_P2_R1131_U267,
    new_P2_R1131_U268, new_P2_R1131_U269, new_P2_R1131_U270,
    new_P2_R1131_U271, new_P2_R1131_U272, new_P2_R1131_U273,
    new_P2_R1131_U274, new_P2_R1131_U275, new_P2_R1131_U276,
    new_P2_R1131_U277, new_P2_R1131_U278, new_P2_R1131_U279,
    new_P2_R1131_U280, new_P2_R1131_U281, new_P2_R1131_U282,
    new_P2_R1131_U283, new_P2_R1131_U284, new_P2_R1131_U285,
    new_P2_R1131_U286, new_P2_R1131_U287, new_P2_R1131_U288,
    new_P2_R1131_U289, new_P2_R1131_U290, new_P2_R1131_U291,
    new_P2_R1131_U292, new_P2_R1131_U293, new_P2_R1131_U294,
    new_P2_R1131_U295, new_P2_R1131_U296, new_P2_R1131_U297,
    new_P2_R1131_U298, new_P2_R1131_U299, new_P2_R1131_U300,
    new_P2_R1131_U301, new_P2_R1131_U302, new_P2_R1131_U303,
    new_P2_R1131_U304, new_P2_R1131_U305, new_P2_R1131_U306,
    new_P2_R1131_U307, new_P2_R1131_U308, new_P2_R1131_U309,
    new_P2_R1131_U310, new_P2_R1131_U311, new_P2_R1131_U312,
    new_P2_R1131_U313, new_P2_R1131_U314, new_P2_R1131_U315,
    new_P2_R1131_U316, new_P2_R1131_U317, new_P2_R1131_U318,
    new_P2_R1131_U319, new_P2_R1131_U320, new_P2_R1131_U321,
    new_P2_R1131_U322, new_P2_R1131_U323, new_P2_R1131_U324,
    new_P2_R1131_U325, new_P2_R1131_U326, new_P2_R1131_U327,
    new_P2_R1131_U328, new_P2_R1131_U329, new_P2_R1131_U330,
    new_P2_R1131_U331, new_P2_R1131_U332, new_P2_R1131_U333,
    new_P2_R1131_U334, new_P2_R1131_U335, new_P2_R1131_U336,
    new_P2_R1131_U337, new_P2_R1131_U338, new_P2_R1131_U339,
    new_P2_R1131_U340, new_P2_R1131_U341, new_P2_R1131_U342,
    new_P2_R1131_U343, new_P2_R1131_U344, new_P2_R1131_U345,
    new_P2_R1131_U346, new_P2_R1131_U347, new_P2_R1131_U348,
    new_P2_R1131_U349, new_P2_R1131_U350, new_P2_R1131_U351,
    new_P2_R1131_U352, new_P2_R1131_U353, new_P2_R1131_U354,
    new_P2_R1131_U355, new_P2_R1131_U356, new_P2_R1131_U357,
    new_P2_R1131_U358, new_P2_R1131_U359, new_P2_R1131_U360,
    new_P2_R1131_U361, new_P2_R1131_U362, new_P2_R1131_U363,
    new_P2_R1131_U364, new_P2_R1131_U365, new_P2_R1131_U366,
    new_P2_R1131_U367, new_P2_R1131_U368, new_P2_R1131_U369,
    new_P2_R1131_U370, new_P2_R1131_U371, new_P2_R1131_U372,
    new_P2_R1131_U373, new_P2_R1131_U374, new_P2_R1131_U375,
    new_P2_R1131_U376, new_P2_R1131_U377, new_P2_R1131_U378,
    new_P2_R1131_U379, new_P2_R1131_U380, new_P2_R1131_U381,
    new_P2_R1131_U382, new_P2_R1131_U383, new_P2_R1131_U384,
    new_P2_R1131_U385, new_P2_R1131_U386, new_P2_R1131_U387,
    new_P2_R1131_U388, new_P2_R1131_U389, new_P2_R1131_U390,
    new_P2_R1131_U391, new_P2_R1131_U392, new_P2_R1131_U393,
    new_P2_R1131_U394, new_P2_R1131_U395, new_P2_R1131_U396,
    new_P2_R1131_U397, new_P2_R1131_U398, new_P2_R1131_U399,
    new_P2_R1131_U400, new_P2_R1131_U401, new_P2_R1131_U402,
    new_P2_R1131_U403, new_P2_R1131_U404, new_P2_R1131_U405,
    new_P2_R1131_U406, new_P2_R1131_U407, new_P2_R1131_U408,
    new_P2_R1131_U409, new_P2_R1131_U410, new_P2_R1131_U411,
    new_P2_R1131_U412, new_P2_R1131_U413, new_P2_R1131_U414,
    new_P2_R1131_U415, new_P2_R1131_U416, new_P2_R1131_U417,
    new_P2_R1131_U418, new_P2_R1131_U419, new_P2_R1131_U420,
    new_P2_R1131_U421, new_P2_R1131_U422, new_P2_R1131_U423,
    new_P2_R1131_U424, new_P2_R1131_U425, new_P2_R1131_U426,
    new_P2_R1131_U427, new_P2_R1131_U428, new_P2_R1131_U429,
    new_P2_R1131_U430, new_P2_R1131_U431, new_P2_R1131_U432,
    new_P2_R1131_U433, new_P2_R1131_U434, new_P2_R1131_U435,
    new_P2_R1131_U436, new_P2_R1131_U437, new_P2_R1131_U438,
    new_P2_R1131_U439, new_P2_R1131_U440, new_P2_R1131_U441,
    new_P2_R1131_U442, new_P2_R1131_U443, new_P2_R1131_U444,
    new_P2_R1131_U445, new_P2_R1131_U446, new_P2_R1131_U447,
    new_P2_R1131_U448, new_P2_R1131_U449, new_P2_R1131_U450,
    new_P2_R1131_U451, new_P2_R1131_U452, new_P2_R1131_U453,
    new_P2_R1131_U454, new_P2_R1131_U455, new_P2_R1131_U456,
    new_P2_R1131_U457, new_P2_R1131_U458, new_P2_R1131_U459,
    new_P2_R1131_U460, new_P2_R1131_U461, new_P2_R1131_U462,
    new_P2_R1131_U463, new_P2_R1131_U464, new_P2_R1131_U465,
    new_P2_R1131_U466, new_P2_R1131_U467, new_P2_R1131_U468,
    new_P2_R1131_U469, new_P2_R1131_U470, new_P2_R1131_U471,
    new_P2_R1131_U472, new_P2_R1131_U473, new_P2_R1131_U474,
    new_P2_R1131_U475, new_P2_R1131_U476, new_P2_R1131_U477,
    new_P2_R1131_U478, new_P2_R1131_U479, new_P2_R1131_U480,
    new_P2_R1131_U481, new_P2_R1131_U482, new_P2_R1131_U483,
    new_P2_R1131_U484, new_P2_R1131_U485, new_P2_R1131_U486,
    new_P2_R1131_U487, new_P2_R1131_U488, new_P2_R1131_U489,
    new_P2_R1054_U6, new_P2_R1054_U7, new_P2_R1054_U8, new_P2_R1054_U9,
    new_P2_R1054_U10, new_P2_R1054_U11, new_P2_R1054_U12, new_P2_R1054_U13,
    new_P2_R1054_U14, new_P2_R1054_U15, new_P2_R1054_U16, new_P2_R1054_U17,
    new_P2_R1054_U18, new_P2_R1054_U19, new_P2_R1054_U20, new_P2_R1054_U21,
    new_P2_R1054_U22, new_P2_R1054_U23, new_P2_R1054_U24, new_P2_R1054_U25,
    new_P2_R1054_U26, new_P2_R1054_U27, new_P2_R1054_U28, new_P2_R1054_U29,
    new_P2_R1054_U30, new_P2_R1054_U31, new_P2_R1054_U32, new_P2_R1054_U33,
    new_P2_R1054_U34, new_P2_R1054_U35, new_P2_R1054_U36, new_P2_R1054_U37,
    new_P2_R1054_U38, new_P2_R1054_U39, new_P2_R1054_U40, new_P2_R1054_U41,
    new_P2_R1054_U42, new_P2_R1054_U43, new_P2_R1054_U44, new_P2_R1054_U45,
    new_P2_R1054_U46, new_P2_R1054_U47, new_P2_R1054_U48, new_P2_R1054_U49,
    new_P2_R1054_U50, new_P2_R1054_U51, new_P2_R1054_U52, new_P2_R1054_U53,
    new_P2_R1054_U54, new_P2_R1054_U55, new_P2_R1054_U56, new_P2_R1054_U57,
    new_P2_R1054_U58, new_P2_R1054_U59, new_P2_R1054_U60, new_P2_R1054_U61,
    new_P2_R1054_U62, new_P2_R1054_U63, new_P2_R1054_U64, new_P2_R1054_U65,
    new_P2_R1054_U66, new_P2_R1054_U67, new_P2_R1054_U68, new_P2_R1054_U69,
    new_P2_R1054_U70, new_P2_R1054_U71, new_P2_R1054_U72, new_P2_R1054_U73,
    new_P2_R1054_U74, new_P2_R1054_U75, new_P2_R1054_U76, new_P2_R1054_U77,
    new_P2_R1054_U78, new_P2_R1054_U79, new_P2_R1054_U80, new_P2_R1054_U81,
    new_P2_R1054_U82, new_P2_R1054_U83, new_P2_R1054_U84, new_P2_R1054_U85,
    new_P2_R1054_U86, new_P2_R1054_U87, new_P2_R1054_U88, new_P2_R1054_U89,
    new_P2_R1054_U90, new_P2_R1054_U91, new_P2_R1054_U92, new_P2_R1054_U93,
    new_P2_R1054_U94, new_P2_R1054_U95, new_P2_R1054_U96, new_P2_R1054_U97,
    new_P2_R1054_U98, new_P2_R1054_U99, new_P2_R1054_U100,
    new_P2_R1054_U101, new_P2_R1054_U102, new_P2_R1054_U103,
    new_P2_R1054_U104, new_P2_R1054_U105, new_P2_R1054_U106,
    new_P2_R1054_U107, new_P2_R1054_U108, new_P2_R1054_U109,
    new_P2_R1054_U110, new_P2_R1054_U111, new_P2_R1054_U112,
    new_P2_R1054_U113, new_P2_R1054_U114, new_P2_R1054_U115,
    new_P2_R1054_U116, new_P2_R1054_U117, new_P2_R1054_U118,
    new_P2_R1054_U119, new_P2_R1054_U120, new_P2_R1054_U121,
    new_P2_R1054_U122, new_P2_R1054_U123, new_P2_R1054_U124,
    new_P2_R1054_U125, new_P2_R1054_U126, new_P2_R1054_U127,
    new_P2_R1054_U128, new_P2_R1054_U129, new_P2_R1054_U130,
    new_P2_R1054_U131, new_P2_R1054_U132, new_P2_R1054_U133,
    new_P2_R1054_U134, new_P2_R1054_U135, new_P2_R1054_U136,
    new_P2_R1054_U137, new_P2_R1054_U138, new_P2_R1054_U139,
    new_P2_R1054_U140, new_P2_R1054_U141, new_P2_R1054_U142,
    new_P2_R1054_U143, new_P2_R1054_U144, new_P2_R1054_U145,
    new_P2_R1054_U146, new_P2_R1054_U147, new_P2_R1054_U148,
    new_P2_R1054_U149, new_P2_R1054_U150, new_P2_R1054_U151,
    new_P2_R1054_U152, new_P2_R1054_U153, new_P2_R1054_U154,
    new_P2_R1054_U155, new_P2_R1054_U156, new_P2_R1054_U157,
    new_P2_R1054_U158, new_P2_R1054_U159, new_P2_R1054_U160,
    new_P2_R1054_U161, new_P2_R1054_U162, new_P2_R1054_U163,
    new_P2_R1054_U164, new_P2_R1054_U165, new_P2_R1054_U166,
    new_P2_R1054_U167, new_P2_R1054_U168, new_P2_R1054_U169,
    new_P2_R1054_U170, new_P2_R1054_U171, new_P2_R1054_U172,
    new_P2_R1054_U173, new_P2_R1054_U174, new_P2_R1054_U175,
    new_P2_R1054_U176, new_P2_R1054_U177, new_P2_R1054_U178,
    new_P2_R1054_U179, new_P2_R1054_U180, new_P2_R1054_U181,
    new_P2_R1054_U182, new_P2_R1054_U183, new_P2_R1054_U184,
    new_P2_R1054_U185, new_P2_R1054_U186, new_P2_R1054_U187,
    new_P2_R1054_U188, new_P2_R1054_U189, new_P2_R1054_U190,
    new_P2_R1054_U191, new_P2_R1054_U192, new_P2_R1054_U193,
    new_P2_R1054_U194, new_P2_R1054_U195, new_P2_R1054_U196,
    new_P2_R1054_U197, new_P2_R1054_U198, new_P2_R1054_U199,
    new_P2_R1054_U200, new_P2_R1054_U201, new_P2_R1054_U202,
    new_P2_R1054_U203, new_P2_R1054_U204, new_P2_R1054_U205,
    new_P2_R1054_U206, new_P2_R1054_U207, new_P2_R1054_U208,
    new_P2_R1054_U209, new_P2_R1054_U210, new_P2_R1054_U211,
    new_P2_R1054_U212, new_P2_R1054_U213, new_P2_R1054_U214,
    new_P2_R1054_U215, new_P2_R1054_U216, new_P2_R1054_U217,
    new_P2_R1054_U218, new_P2_R1054_U219, new_P2_R1054_U220,
    new_P2_R1054_U221, new_P2_R1054_U222, new_P2_R1054_U223,
    new_P2_R1054_U224, new_P2_R1054_U225, new_P2_R1054_U226,
    new_P2_R1054_U227, new_P2_R1054_U228, new_P2_R1054_U229,
    new_P2_R1054_U230, new_P2_R1054_U231, new_P2_R1054_U232,
    new_P2_R1054_U233, new_P2_R1054_U234, new_P2_R1054_U235,
    new_P2_R1054_U236, new_P2_R1054_U237, new_P2_R1054_U238,
    new_P2_R1054_U239, new_P2_R1054_U240, new_P2_R1054_U241,
    new_P2_R1054_U242, new_P2_R1054_U243, new_P2_R1054_U244,
    new_P2_R1054_U245, new_P2_R1054_U246, new_P2_R1054_U247,
    new_P2_R1054_U248, new_P2_R1054_U249, new_P2_R1054_U250,
    new_P2_R1054_U251, new_P2_R1054_U252, new_P2_R1054_U253,
    new_P2_R1054_U254, new_P2_R1054_U255, new_P2_R1054_U256,
    new_P2_R1054_U257, new_P2_R1054_U258, new_P2_R1054_U259,
    new_P2_R1054_U260, new_P2_R1054_U261, new_P2_R1054_U262,
    new_P2_R1054_U263, new_P2_R1054_U264, new_P2_R1054_U265,
    new_P2_R1054_U266, new_P2_R1054_U267, new_P2_R1054_U268,
    new_P2_R1054_U269, new_P2_R1054_U270, new_P2_R1054_U271,
    new_P2_R1054_U272, new_P2_R1054_U273, new_P2_R1054_U274,
    new_P2_R1054_U275, new_P2_R1054_U276, new_P2_R1054_U277,
    new_P2_R1054_U278, new_P2_R1054_U279, new_P2_R1054_U280,
    new_P2_R1054_U281, new_P2_R1054_U282, new_P2_R1054_U283,
    new_P2_R1054_U284, new_P2_R1054_U285, new_P2_R1054_U286,
    new_P2_R1054_U287, new_P2_R1054_U288, new_P2_R1054_U289,
    new_P2_R1054_U290, new_P2_R1054_U291, new_P2_R1054_U292,
    new_P2_R1054_U293, new_P2_R1054_U294, new_P2_R1161_U4, new_P2_R1161_U5,
    new_P2_R1161_U6, new_P2_R1161_U7, new_P2_R1161_U8, new_P2_R1161_U9,
    new_P2_R1161_U10, new_P2_R1161_U11, new_P2_R1161_U12, new_P2_R1161_U13,
    new_P2_R1161_U14, new_P2_R1161_U15, new_P2_R1161_U16, new_P2_R1161_U17,
    new_P2_R1161_U18, new_P2_R1161_U19, new_P2_R1161_U20, new_P2_R1161_U21,
    new_P2_R1161_U22, new_P2_R1161_U23, new_P2_R1161_U24, new_P2_R1161_U25,
    new_P2_R1161_U26, new_P2_R1161_U27, new_P2_R1161_U28, new_P2_R1161_U29,
    new_P2_R1161_U30, new_P2_R1161_U31, new_P2_R1161_U32, new_P2_R1161_U33,
    new_P2_R1161_U34, new_P2_R1161_U35, new_P2_R1161_U36, new_P2_R1161_U37,
    new_P2_R1161_U38, new_P2_R1161_U39, new_P2_R1161_U40, new_P2_R1161_U41,
    new_P2_R1161_U42, new_P2_R1161_U43, new_P2_R1161_U44, new_P2_R1161_U45,
    new_P2_R1161_U46, new_P2_R1161_U47, new_P2_R1161_U48, new_P2_R1161_U49,
    new_P2_R1161_U50, new_P2_R1161_U51, new_P2_R1161_U52, new_P2_R1161_U53,
    new_P2_R1161_U54, new_P2_R1161_U55, new_P2_R1161_U56, new_P2_R1161_U57,
    new_P2_R1161_U58, new_P2_R1161_U59, new_P2_R1161_U60, new_P2_R1161_U61,
    new_P2_R1161_U62, new_P2_R1161_U63, new_P2_R1161_U64, new_P2_R1161_U65,
    new_P2_R1161_U66, new_P2_R1161_U67, new_P2_R1161_U68, new_P2_R1161_U69,
    new_P2_R1161_U70, new_P2_R1161_U71, new_P2_R1161_U72, new_P2_R1161_U73,
    new_P2_R1161_U74, new_P2_R1161_U75, new_P2_R1161_U76, new_P2_R1161_U77,
    new_P2_R1161_U78, new_P2_R1161_U79, new_P2_R1161_U80, new_P2_R1161_U81,
    new_P2_R1161_U82, new_P2_R1161_U83, new_P2_R1161_U84, new_P2_R1161_U85,
    new_P2_R1161_U86, new_P2_R1161_U87, new_P2_R1161_U88, new_P2_R1161_U89,
    new_P2_R1161_U90, new_P2_R1161_U91, new_P2_R1161_U92, new_P2_R1161_U93,
    new_P2_R1161_U94, new_P2_R1161_U95, new_P2_R1161_U96, new_P2_R1161_U97,
    new_P2_R1161_U98, new_P2_R1161_U99, new_P2_R1161_U100,
    new_P2_R1161_U101, new_P2_R1161_U102, new_P2_R1161_U103,
    new_P2_R1161_U104, new_P2_R1161_U105, new_P2_R1161_U106,
    new_P2_R1161_U107, new_P2_R1161_U108, new_P2_R1161_U109,
    new_P2_R1161_U110, new_P2_R1161_U111, new_P2_R1161_U112,
    new_P2_R1161_U113, new_P2_R1161_U114, new_P2_R1161_U115,
    new_P2_R1161_U116, new_P2_R1161_U117, new_P2_R1161_U118,
    new_P2_R1161_U119, new_P2_R1161_U120, new_P2_R1161_U121,
    new_P2_R1161_U122, new_P2_R1161_U123, new_P2_R1161_U124,
    new_P2_R1161_U125, new_P2_R1161_U126, new_P2_R1161_U127,
    new_P2_R1161_U128, new_P2_R1161_U129, new_P2_R1161_U130,
    new_P2_R1161_U131, new_P2_R1161_U132, new_P2_R1161_U133,
    new_P2_R1161_U134, new_P2_R1161_U135, new_P2_R1161_U136,
    new_P2_R1161_U137, new_P2_R1161_U138, new_P2_R1161_U139,
    new_P2_R1161_U140, new_P2_R1161_U141, new_P2_R1161_U142,
    new_P2_R1161_U143, new_P2_R1161_U144, new_P2_R1161_U145,
    new_P2_R1161_U146, new_P2_R1161_U147, new_P2_R1161_U148,
    new_P2_R1161_U149, new_P2_R1161_U150, new_P2_R1161_U151,
    new_P2_R1161_U152, new_P2_R1161_U153, new_P2_R1161_U154,
    new_P2_R1161_U155, new_P2_R1161_U156, new_P2_R1161_U157,
    new_P2_R1161_U158, new_P2_R1161_U159, new_P2_R1161_U160,
    new_P2_R1161_U161, new_P2_R1161_U162, new_P2_R1161_U163,
    new_P2_R1161_U164, new_P2_R1161_U165, new_P2_R1161_U166,
    new_P2_R1161_U167, new_P2_R1161_U168, new_P2_R1161_U169,
    new_P2_R1161_U170, new_P2_R1161_U171, new_P2_R1161_U172,
    new_P2_R1161_U173, new_P2_R1161_U174, new_P2_R1161_U175,
    new_P2_R1161_U176, new_P2_R1161_U177, new_P2_R1161_U178,
    new_P2_R1161_U179, new_P2_R1161_U180, new_P2_R1161_U181,
    new_P2_R1161_U182, new_P2_R1161_U183, new_P2_R1161_U184,
    new_P2_R1161_U185, new_P2_R1161_U186, new_P2_R1161_U187,
    new_P2_R1161_U188, new_P2_R1161_U189, new_P2_R1161_U190,
    new_P2_R1161_U191, new_P2_R1161_U192, new_P2_R1161_U193,
    new_P2_R1161_U194, new_P2_R1161_U195, new_P2_R1161_U196,
    new_P2_R1161_U197, new_P2_R1161_U198, new_P2_R1161_U199,
    new_P2_R1161_U200, new_P2_R1161_U201, new_P2_R1161_U202,
    new_P2_R1161_U203, new_P2_R1161_U204, new_P2_R1161_U205,
    new_P2_R1161_U206, new_P2_R1161_U207, new_P2_R1161_U208,
    new_P2_R1161_U209, new_P2_R1161_U210, new_P2_R1161_U211,
    new_P2_R1161_U212, new_P2_R1161_U213, new_P2_R1161_U214,
    new_P2_R1161_U215, new_P2_R1161_U216, new_P2_R1161_U217,
    new_P2_R1161_U218, new_P2_R1161_U219, new_P2_R1161_U220,
    new_P2_R1161_U221, new_P2_R1161_U222, new_P2_R1161_U223,
    new_P2_R1161_U224, new_P2_R1161_U225, new_P2_R1161_U226,
    new_P2_R1161_U227, new_P2_R1161_U228, new_P2_R1161_U229,
    new_P2_R1161_U230, new_P2_R1161_U231, new_P2_R1161_U232,
    new_P2_R1161_U233, new_P2_R1161_U234, new_P2_R1161_U235,
    new_P2_R1161_U236, new_P2_R1161_U237, new_P2_R1161_U238,
    new_P2_R1161_U239, new_P2_R1161_U240, new_P2_R1161_U241,
    new_P2_R1161_U242, new_P2_R1161_U243, new_P2_R1161_U244,
    new_P2_R1161_U245, new_P2_R1161_U246, new_P2_R1161_U247,
    new_P2_R1161_U248, new_P2_R1161_U249, new_P2_R1161_U250,
    new_P2_R1161_U251, new_P2_R1161_U252, new_P2_R1161_U253,
    new_P2_R1161_U254, new_P2_R1161_U255, new_P2_R1161_U256,
    new_P2_R1161_U257, new_P2_R1161_U258, new_P2_R1161_U259,
    new_P2_R1161_U260, new_P2_R1161_U261, new_P2_R1161_U262,
    new_P2_R1161_U263, new_P2_R1161_U264, new_P2_R1161_U265,
    new_P2_R1161_U266, new_P2_R1161_U267, new_P2_R1161_U268,
    new_P2_R1161_U269, new_P2_R1161_U270, new_P2_R1161_U271,
    new_P2_R1161_U272, new_P2_R1161_U273, new_P2_R1161_U274,
    new_P2_R1161_U275, new_P2_R1161_U276, new_P2_R1161_U277,
    new_P2_R1161_U278, new_P2_R1161_U279, new_P2_R1161_U280,
    new_P2_R1161_U281, new_P2_R1161_U282, new_P2_R1161_U283,
    new_P2_R1161_U284, new_P2_R1161_U285, new_P2_R1161_U286,
    new_P2_R1161_U287, new_P2_R1161_U288, new_P2_R1161_U289,
    new_P2_R1161_U290, new_P2_R1161_U291, new_P2_R1161_U292,
    new_P2_R1161_U293, new_P2_R1161_U294, new_P2_R1161_U295,
    new_P2_R1161_U296, new_P2_R1161_U297, new_P2_R1161_U298,
    new_P2_R1161_U299, new_P2_R1161_U300, new_P2_R1161_U301,
    new_P2_R1161_U302, new_P2_R1161_U303, new_P2_R1161_U304,
    new_P2_R1161_U305, new_P2_R1161_U306, new_P2_R1161_U307,
    new_P2_R1161_U308, new_P2_R1161_U309, new_P2_R1161_U310,
    new_P2_R1161_U311, new_P2_R1161_U312, new_P2_R1161_U313,
    new_P2_R1161_U314, new_P2_R1161_U315, new_P2_R1161_U316,
    new_P2_R1161_U317, new_P2_R1161_U318, new_P2_R1161_U319,
    new_P2_R1161_U320, new_P2_R1161_U321, new_P2_R1161_U322,
    new_P2_R1161_U323, new_P2_R1161_U324, new_P2_R1161_U325,
    new_P2_R1161_U326, new_P2_R1161_U327, new_P2_R1161_U328,
    new_P2_R1161_U329, new_P2_R1161_U330, new_P2_R1161_U331,
    new_P2_R1161_U332, new_P2_R1161_U333, new_P2_R1161_U334,
    new_P2_R1161_U335, new_P2_R1161_U336, new_P2_R1161_U337,
    new_P2_R1161_U338, new_P2_R1161_U339, new_P2_R1161_U340,
    new_P2_R1161_U341, new_P2_R1161_U342, new_P2_R1161_U343,
    new_P2_R1161_U344, new_P2_R1161_U345, new_P2_R1161_U346,
    new_P2_R1161_U347, new_P2_R1161_U348, new_P2_R1161_U349,
    new_P2_R1161_U350, new_P2_R1161_U351, new_P2_R1161_U352,
    new_P2_R1161_U353, new_P2_R1161_U354, new_P2_R1161_U355,
    new_P2_R1161_U356, new_P2_R1161_U357, new_P2_R1161_U358,
    new_P2_R1161_U359, new_P2_R1161_U360, new_P2_R1161_U361,
    new_P2_R1161_U362, new_P2_R1161_U363, new_P2_R1161_U364,
    new_P2_R1161_U365, new_P2_R1161_U366, new_P2_R1161_U367,
    new_P2_R1161_U368, new_P2_R1161_U369, new_P2_R1161_U370,
    new_P2_R1161_U371, new_P2_R1161_U372, new_P2_R1161_U373,
    new_P2_R1161_U374, new_P2_R1161_U375, new_P2_R1161_U376,
    new_P2_R1161_U377, new_P2_R1161_U378, new_P2_R1161_U379,
    new_P2_R1161_U380, new_P2_R1161_U381, new_P2_R1161_U382,
    new_P2_R1161_U383, new_P2_R1161_U384, new_P2_R1161_U385,
    new_P2_R1161_U386, new_P2_R1161_U387, new_P2_R1161_U388,
    new_P2_R1161_U389, new_P2_R1161_U390, new_P2_R1161_U391,
    new_P2_R1161_U392, new_P2_R1161_U393, new_P2_R1161_U394,
    new_P2_R1161_U395, new_P2_R1161_U396, new_P2_R1161_U397,
    new_P2_R1161_U398, new_P2_R1161_U399, new_P2_R1161_U400,
    new_P2_R1161_U401, new_P2_R1161_U402, new_P2_R1161_U403,
    new_P2_R1161_U404, new_P2_R1161_U405, new_P2_R1161_U406,
    new_P2_R1161_U407, new_P2_R1161_U408, new_P2_R1161_U409,
    new_P2_R1161_U410, new_P2_R1161_U411, new_P2_R1161_U412,
    new_P2_R1161_U413, new_P2_R1161_U414, new_P2_R1161_U415,
    new_P2_R1161_U416, new_P2_R1161_U417, new_P2_R1161_U418,
    new_P2_R1161_U419, new_P2_R1161_U420, new_P2_R1161_U421,
    new_P2_R1161_U422, new_P2_R1161_U423, new_P2_R1161_U424,
    new_P2_R1161_U425, new_P2_R1161_U426, new_P2_R1161_U427,
    new_P2_R1161_U428, new_P2_R1161_U429, new_P2_R1161_U430,
    new_P2_R1161_U431, new_P2_R1161_U432, new_P2_R1161_U433,
    new_P2_R1161_U434, new_P2_R1161_U435, new_P2_R1161_U436,
    new_P2_R1161_U437, new_P2_R1161_U438, new_P2_R1161_U439,
    new_P2_R1161_U440, new_P2_R1161_U441, new_P2_R1161_U442,
    new_P2_R1161_U443, new_P2_R1161_U444, new_P2_R1161_U445,
    new_P2_R1161_U446, new_not_keyinput0, new_not_keyinput1,
    new_not_keyinput2, new_not_keyinput3, new_not_keyinput4, new_not_0,
    new_and_1, new_not_2, new_and_3, new_not_4, new_and_5, new_not_6,
    new_and_7, new_not_9, new_and_10, new_not_11, new_and_12, new_not_13,
    new_and_14, new_not_16, new_and_17, new_not_18, new_and_19,
    new_not_Q_0, new_not_Q_1, new_not_Q_2, new_not_Q_3, new_count_state_1,
    new_count_state_2, new_count_state_3, new_count_state_4,
    new_count_state_5, new_count_state_6, new_count_state_7,
    new_count_state_8, new_count_state_9, new_count_state_10,
    new_count_state_11, new_count_state_12, new_count_state_13,
    new_count_state_14, new_count_state_15, new_y_mux_key0_and_0,
    new_y_mux_key0_and_1, new_y_mux_key0, new_y_mux_key1_and_0,
    new_y_mux_key1_and_1, new_y_mux_key1, new_y_mux_key2_and_0,
    new_y_mux_key2_and_1, new_y_mux_key2, new_y_mux_key3_and_0,
    new_y_mux_key3_and_1, new_y_mux_key3, new_y_mux_key4_and_0,
    new_y_mux_key4_and_1, new_y_mux_key4, new_y_mux_key5_and_0,
    new_y_mux_key5_and_1, new_y_mux_key5, new_y_mux_key6_and_0,
    new_y_mux_key6_and_1, new_y_mux_key6, new_y_mux_key7_and_0,
    new_y_mux_key7_and_1, new_y_mux_key7, new_y_mux_key8_and_0,
    new_y_mux_key8_and_1, new_y_mux_key8, new_y_mux_key9_and_0,
    new_y_mux_key9_and_1, new_y_mux_key9, new_y_mux_key10_and_0,
    new_y_mux_key10_and_1, new_y_mux_key10, new_y_mux_key11_and_0,
    new_y_mux_key11_and_1, new_y_mux_key11, new_y_mux_key12_and_0,
    new_y_mux_key12_and_1, new_y_mux_key12, new_y_mux_key13_and_0,
    new_y_mux_key13_and_1, new_y_mux_key13, new_y_mux_key14_and_0,
    new_y_mux_key14_and_1, new_y_mux_key14, new_y_mux_key15_and_0,
    new_y_mux_key15_and_1, new_y_mux_key15, new__state_1, new__state_2,
    new__state_3, new__state_4, new__state_5, new__state_6, new__state_7,
    new__state_8, new__state_9, new__state_10, new__state_11,
    new__state_12, new__state_13, new__state_14, new__state_15,
    new__state_17, new__state_18, new__state_19, new__state_20,
    new__state_21, new__state_22, new__state_23, new__state_25,
    new__state_26, new__state_27, new__state_29, new_s__state_1,
    new_not_s__state_1, new_I0__state_1, new_I1__state_1,
    new_and_mux__state_1, new_and_mux__state_1_2, new_y_mux_16,
    new_s__state_3, new_not_s__state_3, new_I0__state_3, new_I1__state_3,
    new_and_mux__state_3, new_and_mux__state_3_2, new_y_mux_17,
    new_s__state_5, new_not_s__state_5, new_I0__state_5, new_I1__state_5,
    new_and_mux__state_5, new_and_mux__state_5_2, new_y_mux_18,
    new_s__state_7, new_not_s__state_7, new_I0__state_7, new_I1__state_7,
    new_and_mux__state_7, new_and_mux__state_7_2, new_y_mux_19,
    new_s__state_9, new_not_s__state_9, new_I0__state_9, new_I1__state_9,
    new_and_mux__state_9, new_and_mux__state_9_2, new_y_mux_20,
    new_s__state_11, new_not_s__state_11, new_I0__state_11,
    new_I1__state_11, new_and_mux__state_11, new_and_mux__state_11_2,
    new_y_mux_21, new_s__state_13, new_not_s__state_13, new_I0__state_13,
    new_I1__state_13, new_and_mux__state_13, new_and_mux__state_13_2,
    new_y_mux_22, new_s__state_15, new_not_s__state_15, new_I0__state_15,
    new_I1__state_15, new_and_mux__state_15, new_and_mux__state_15_2,
    new_y_mux_23, new_s__state_17, new_not_s__state_17, new_I0__state_17,
    new_I1__state_17, new_and_mux__state_17, new_and_mux__state_17_2,
    new_y_mux_24, new_s__state_19, new_not_s__state_19, new_I0__state_19,
    new_I1__state_19, new_and_mux__state_19, new_and_mux__state_19_2,
    new_y_mux_25, new_s__state_21, new_not_s__state_21, new_I0__state_21,
    new_I1__state_21, new_and_mux__state_21, new_and_mux__state_21_2,
    new_y_mux_26, new_s__state_23, new_not_s__state_23, new_I0__state_23,
    new_I1__state_23, new_and_mux__state_23, new_and_mux__state_23_2,
    new_y_mux_27, new_s__state_25, new_not_s__state_25, new_I0__state_25,
    new_I1__state_25, new_and_mux__state_25, new_and_mux__state_25_2,
    new_y_mux_28, new_s__state_27, new_not_s__state_27, new_I0__state_27,
    new_I1__state_27, new_and_mux__state_27, new_and_mux__state_27_2,
    new_y_mux_29, new_s__state_29, new_not_s__state_29, new_I0__state_29,
    new_I1__state_29, new_and_mux__state_29, new_and_mux__state_29_2, n120,
    n125, n130, n135, n140, n145, n150, n155, n160, n165, n170, n175, n180,
    n185, n190, n195, n200, n205, n210, n215, n220, n225, n230, n235, n240,
    n245, n250, n255, n260, n265, n270, n275, n280, n285, n290, n295, n300,
    n305, n310, n315, n320, n325, n330, n335, n340, n345, n350, n355, n360,
    n365, n370, n375, n380, n385, n390, n395, n400, n405, n410, n415, n420,
    n425, n430, n435, n440, n445, n450, n455, n460, n465, n470, n475, n480,
    n485, n490, n495, n500, n505, n510, n515, n520, n525, n530, n535, n540,
    n545, n550, n555, n560, n565, n570, n575, n580, n585, n590, n595, n600,
    n605, n610, n615, n620, n625, n630, n635, n640, n645, n650, n655, n660,
    n665, n670, n675, n680, n685, n690, n695, n700, n705, n710, n715, n720,
    n725, n730, n735, n740, n745, n750, n755, n760, n765, n770, n775, n780,
    n785, n790, n795, n800, n805, n810, n815, n820, n825, n830, n835, n840,
    n845, n850, n855, n860, n865, n870, n875, n880, n885, n890, n895, n900,
    n905, n910, n915, n920, n925, n930, n935, n940, n945, n950, n955, n960,
    n965, n970, n975, n980, n985, n990, n995, n1000, n1005, n1010, n1015,
    n1020, n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065,
    n1070, n1075, n1080, n1085, n1090, n1095, n1100, n1105, n1110, n1115,
    n1120, n1125, n1130, n1135, n1140, n1145, n1150, n1155, n1160, n1165,
    n1170, n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215,
    n1220, n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265,
    n1270, n1275, n1280, n1285, n1290, n1295, n1300, n1305, n1310, n1315,
    n1320, n1325, n1330, n1335, n1340, n1345, n1350, n1355, n1360, n1365,
    n1370, n1375, n1380, n1385, n1390, n1395, n1400, n1405, n1410, n1415,
    n1420, n1425, n1430, n1435, n1440, n1445, n1450, n1455, n1460, n1465,
    n1470, n1475, n1480, n1485, n1490, n1495, n1500, n1505, n1510, n1515,
    n1520, n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565,
    n1570, n1575, n1580, n1585, n1590, n1595, n1600, n1605, n1610, n1615,
    n1620, n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665,
    n1670, n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715,
    n1720, n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765,
    n1770, n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815,
    n1820, n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865,
    n1870, n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1910, n1915,
    n1920, n1925, n1930, n1935, n1940, n1945, n1950, n1955, n1960, n1965,
    n1970, n1975, n1980, n1985, n1990, n1995, n2000, n2005, n2010, n2015,
    n2020, n2025, n2030, n2035, n2040, n2045, n2050, n2055, n2060, n2065,
    n2070, n2075, n2080, n2085, n2090, n2095, n2100, n2105, n2110, n2115,
    n2120, n2125, n2130, n2135, n2140, n2145, n2150, n2155, n2160, n2165,
    n2170, n2175, n2180, n2185, n2190, n2195, n2200, n2205, n2210, n2215,
    n2220, n2225, n2230, n2235, n2240, n2245, n2250, n2255, n2260, n2265,
    n2270, n2275, n2280, n2285, n2290, n2295, n2300, n2305, n2310, n2315,
    n2320, n2325, n2330, n2335, n2340, n2345, n2350, n2355, n2360, n2365,
    n2370, n2375, n2380, n2385, n2390, n2395, n2400, n2405, n2410, n2415,
    n2420, n2425, n2430, n2435, n2440, n2445, n2450, n2455, n2460, n2465,
    n2470, n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510, n2515,
    n2520, n2525, n2530, n2535, n2540, n2545, n2550, n2555, n2560, n2565,
    n41480, n41483, n41486, n41489;
  assign new_P2_R1161_U504 = ~new_P2_U3387 | ~new_P2_R1161_U30;
  assign new_P2_R1161_U503 = ~new_P2_U3076 | ~new_P2_R1161_U29;
  assign new_P2_R1161_U502 = ~new_P2_U3419 | ~new_P2_R1161_U64;
  assign new_U25 = ~new_U136 | ~new_U135;
  assign new_U26 = ~new_U138 | ~new_U137;
  assign new_U27 = ~new_U140 | ~new_U139;
  assign new_U28 = ~new_U142 | ~new_U141;
  assign new_U29 = ~new_U144 | ~new_U143;
  assign new_U30 = ~new_U146 | ~new_U145;
  assign new_U31 = ~new_U148 | ~new_U147;
  assign new_U32 = ~new_U150 | ~new_U149;
  assign new_U33 = ~new_U152 | ~new_U151;
  assign new_U34 = ~new_U154 | ~new_U153;
  assign new_U35 = ~new_U156 | ~new_U155;
  assign new_U36 = ~new_U158 | ~new_U157;
  assign new_U37 = ~new_U160 | ~new_U159;
  assign new_U38 = ~new_U162 | ~new_U161;
  assign new_U39 = ~new_U164 | ~new_U163;
  assign new_U40 = ~new_U166 | ~new_U165;
  assign new_U41 = ~new_U168 | ~new_U167;
  assign new_U42 = ~new_U170 | ~new_U169;
  assign new_U43 = ~new_U172 | ~new_U171;
  assign new_U44 = ~new_U174 | ~new_U173;
  assign new_U45 = ~new_U176 | ~new_U175;
  assign new_U46 = ~new_U178 | ~new_U177;
  assign new_U47 = ~new_U180 | ~new_U179;
  assign new_U48 = ~new_U182 | ~new_U181;
  assign new_U49 = ~new_U184 | ~new_U183;
  assign new_U50 = ~new_U186 | ~new_U185;
  assign new_U51 = ~new_U188 | ~new_U187;
  assign new_U52 = ~new_U190 | ~new_U189;
  assign new_U53 = ~new_U192 | ~new_U191;
  assign new_U54 = ~new_U194 | ~new_U193;
  assign new_U55 = ~new_U196 | ~new_U195;
  assign new_U56 = ~new_U198 | ~new_U197;
  assign new_U57 = ~new_U200 | ~new_U199;
  assign new_U58 = ~new_U202 | ~new_U201;
  assign new_U59 = ~new_U204 | ~new_U203;
  assign new_U60 = ~new_U206 | ~new_U205;
  assign new_U61 = ~new_U208 | ~new_U207;
  assign new_U62 = ~new_U210 | ~new_U209;
  assign new_U63 = ~new_U212 | ~new_U211;
  assign new_U64 = ~new_U214 | ~new_U213;
  assign new_U65 = ~new_U216 | ~new_U215;
  assign new_U66 = ~new_U218 | ~new_U217;
  assign new_U67 = ~new_U220 | ~new_U219;
  assign new_U68 = ~new_U222 | ~new_U221;
  assign new_U69 = ~new_U224 | ~new_U223;
  assign new_U70 = ~new_U226 | ~new_U225;
  assign new_U71 = ~new_U228 | ~new_U227;
  assign new_U72 = ~new_U230 | ~new_U229;
  assign new_U73 = ~new_U232 | ~new_U231;
  assign new_U74 = ~new_U234 | ~new_U233;
  assign new_U75 = ~new_U236 | ~new_U235;
  assign new_U76 = ~new_U238 | ~new_U237;
  assign new_U77 = ~new_U240 | ~new_U239;
  assign new_U78 = ~new_U242 | ~new_U241;
  assign new_U79 = ~new_U244 | ~new_U243;
  assign new_U80 = ~new_U246 | ~new_U245;
  assign new_U81 = ~new_U248 | ~new_U247;
  assign new_U82 = ~new_U250 | ~new_U249;
  assign new_U83 = ~new_U252 | ~new_U251;
  assign new_U84 = ~new_U254 | ~new_U253;
  assign new_U85 = ~new_U256 | ~new_U255;
  assign new_U86 = ~new_U258 | ~new_U257;
  assign new_U87 = ~new_U260 | ~new_U259;
  assign new_U88 = ~new_U262 | ~new_U261;
  assign new_U89 = ~new_U264 | ~new_U263;
  assign new_U90 = ~new_U266 | ~new_U265;
  assign new_U91 = ~new_U268 | ~new_U267;
  assign new_U92 = ~new_U270 | ~new_U269;
  assign new_U93 = ~new_U272 | ~new_U271;
  assign new_U94 = ~new_U274 | ~new_U273;
  assign new_U95 = ~new_U276 | ~new_U275;
  assign new_U96 = ~new_U278 | ~new_U277;
  assign new_U97 = ~new_U280 | ~new_U279;
  assign new_U98 = ~new_U282 | ~new_U281;
  assign new_U99 = ~new_U284 | ~new_U283;
  assign new_U100 = ~new_U286 | ~new_U285;
  assign new_U101 = ~new_U288 | ~new_U287;
  assign new_U102 = ~new_U290 | ~new_U289;
  assign new_U103 = ~new_U292 | ~new_U291;
  assign new_U104 = ~new_U294 | ~new_U293;
  assign new_U105 = ~new_U296 | ~new_U295;
  assign new_U106 = ~new_U298 | ~new_U297;
  assign new_U107 = ~new_U300 | ~new_U299;
  assign new_U108 = ~new_U302 | ~new_U301;
  assign new_U109 = ~new_U304 | ~new_U303;
  assign new_U110 = ~new_U306 | ~new_U305;
  assign new_U111 = ~new_U308 | ~new_U307;
  assign new_U112 = ~new_U310 | ~new_U309;
  assign new_U113 = ~new_U312 | ~new_U311;
  assign new_U114 = ~new_U314 | ~new_U313;
  assign new_U115 = ~new_U316 | ~new_U315;
  assign new_U116 = ~new_U318 | ~new_U317;
  assign new_U117 = ~new_U320 | ~new_U319;
  assign new_U118 = ~new_U322 | ~new_U321;
  assign new_U119 = ~new_U324 | ~new_U323;
  assign new_U120 = ~new_U326 | ~new_U325;
  assign new_U121 = ~P2_WR_REG;
  assign new_U122 = ~P1_WR_REG;
  assign U123 = new_U132 & new_U131;
  assign new_U124 = ~P2_RD_REG;
  assign new_U125 = ~P1_RD_REG;
  assign U126 = new_U134 & new_U133;
  assign new_U127 = ~new_U129 | ~new_U128;
  assign new_U128 = ~new_LT_1075_19_U6 | ~new_LT_1075_U6 | ~new_U125;
  assign new_U129 = ~P2_ADDR_REG_19_ | ~P1_ADDR_REG_19_ | ~new_U124;
  assign new_U130 = ~new_U127;
  assign new_U131 = ~P2_WR_REG | ~new_U122;
  assign new_U132 = ~P1_WR_REG | ~new_U121;
  assign new_U133 = ~P2_RD_REG | ~new_U125;
  assign new_U134 = ~P1_RD_REG | ~new_U124;
  assign new_U135 = ~P1_DATAO_REG_9_ | ~new_U127;
  assign new_U136 = ~new_R140_U84 | ~new_U130;
  assign new_U137 = ~P1_DATAO_REG_8_ | ~new_U127;
  assign new_U138 = ~new_R140_U85 | ~new_U130;
  assign new_U139 = ~P1_DATAO_REG_7_ | ~new_U127;
  assign new_U140 = ~new_R140_U86 | ~new_U130;
  assign new_U141 = ~P1_DATAO_REG_6_ | ~new_U127;
  assign new_U142 = ~new_R140_U87 | ~new_U130;
  assign new_U143 = ~P1_DATAO_REG_5_ | ~new_U127;
  assign new_U144 = ~new_R140_U88 | ~new_U130;
  assign new_U145 = ~P1_DATAO_REG_4_ | ~new_U127;
  assign new_U146 = ~new_R140_U89 | ~new_U130;
  assign new_U147 = ~P1_DATAO_REG_3_ | ~new_U127;
  assign new_U148 = ~new_R140_U90 | ~new_U130;
  assign new_U149 = ~P1_DATAO_REG_31_ | ~new_U127;
  assign new_U150 = ~new_R140_U11 | ~new_U130;
  assign new_U151 = ~P1_DATAO_REG_30_ | ~new_U127;
  assign new_U152 = ~new_R140_U91 | ~new_U130;
  assign new_U153 = ~P1_DATAO_REG_2_ | ~new_U127;
  assign new_U154 = ~new_R140_U92 | ~new_U130;
  assign new_U155 = ~P1_DATAO_REG_29_ | ~new_U127;
  assign new_U156 = ~new_R140_U93 | ~new_U130;
  assign new_U157 = ~P1_DATAO_REG_28_ | ~new_U127;
  assign new_U158 = ~new_R140_U94 | ~new_U130;
  assign new_U159 = ~P1_DATAO_REG_27_ | ~new_U127;
  assign new_U160 = ~new_R140_U95 | ~new_U130;
  assign new_U161 = ~P1_DATAO_REG_26_ | ~new_U127;
  assign new_U162 = ~new_R140_U96 | ~new_U130;
  assign new_U163 = ~P1_DATAO_REG_25_ | ~new_U127;
  assign new_U164 = ~new_R140_U97 | ~new_U130;
  assign new_U165 = ~P1_DATAO_REG_24_ | ~new_U127;
  assign new_U166 = ~new_R140_U98 | ~new_U130;
  assign new_U167 = ~P1_DATAO_REG_23_ | ~new_U127;
  assign new_U168 = ~new_R140_U99 | ~new_U130;
  assign new_U169 = ~P1_DATAO_REG_22_ | ~new_U127;
  assign new_U170 = ~new_R140_U100 | ~new_U130;
  assign new_U171 = ~P1_DATAO_REG_21_ | ~new_U127;
  assign new_U172 = ~new_R140_U101 | ~new_U130;
  assign new_U173 = ~P1_DATAO_REG_20_ | ~new_U127;
  assign new_U174 = ~new_R140_U102 | ~new_U130;
  assign new_U175 = ~P1_DATAO_REG_1_ | ~new_U127;
  assign new_U176 = ~new_R140_U10 | ~new_U130;
  assign new_U177 = ~P1_DATAO_REG_19_ | ~new_U127;
  assign new_U178 = ~new_R140_U103 | ~new_U130;
  assign new_U179 = ~P1_DATAO_REG_18_ | ~new_U127;
  assign new_U180 = ~new_R140_U104 | ~new_U130;
  assign new_U181 = ~P1_DATAO_REG_17_ | ~new_U127;
  assign new_U182 = ~new_R140_U105 | ~new_U130;
  assign new_U183 = ~P1_DATAO_REG_16_ | ~new_U127;
  assign new_U184 = ~new_R140_U106 | ~new_U130;
  assign new_U185 = ~P1_DATAO_REG_15_ | ~new_U127;
  assign new_U186 = ~new_R140_U107 | ~new_U130;
  assign new_U187 = ~P1_DATAO_REG_14_ | ~new_U127;
  assign new_U188 = ~new_R140_U108 | ~new_U130;
  assign new_U189 = ~P1_DATAO_REG_13_ | ~new_U127;
  assign new_U190 = ~new_R140_U109 | ~new_U130;
  assign new_U191 = ~P1_DATAO_REG_12_ | ~new_U127;
  assign new_U192 = ~new_R140_U110 | ~new_U130;
  assign new_U193 = ~P1_DATAO_REG_11_ | ~new_U127;
  assign new_U194 = ~new_R140_U111 | ~new_U130;
  assign new_U195 = ~P1_DATAO_REG_10_ | ~new_U127;
  assign new_U196 = ~new_R140_U112 | ~new_U130;
  assign new_U197 = ~P1_DATAO_REG_0_ | ~new_U127;
  assign new_U198 = ~new_R140_U83 | ~new_U130;
  assign new_U199 = ~new_R140_U84 | ~new_U127;
  assign new_U200 = ~P2_DATAO_REG_9_ | ~new_U130;
  assign new_U201 = ~new_R140_U85 | ~new_U127;
  assign new_U202 = ~P2_DATAO_REG_8_ | ~new_U130;
  assign new_U203 = ~new_R140_U86 | ~new_U127;
  assign new_U204 = ~P2_DATAO_REG_7_ | ~new_U130;
  assign new_U205 = ~new_R140_U87 | ~new_U127;
  assign new_U206 = ~P2_DATAO_REG_6_ | ~new_U130;
  assign new_U207 = ~new_R140_U88 | ~new_U127;
  assign new_U208 = ~P2_DATAO_REG_5_ | ~new_U130;
  assign new_U209 = ~new_R140_U89 | ~new_U127;
  assign new_U210 = ~P2_DATAO_REG_4_ | ~new_U130;
  assign new_U211 = ~new_R140_U90 | ~new_U127;
  assign new_U212 = ~P2_DATAO_REG_3_ | ~new_U130;
  assign new_U213 = ~new_R140_U11 | ~new_U127;
  assign new_U214 = ~P2_DATAO_REG_31_ | ~new_U130;
  assign new_U215 = ~new_R140_U91 | ~new_U127;
  assign new_U216 = ~P2_DATAO_REG_30_ | ~new_U130;
  assign new_U217 = ~new_R140_U92 | ~new_U127;
  assign new_U218 = ~P2_DATAO_REG_2_ | ~new_U130;
  assign new_U219 = ~new_R140_U93 | ~new_U127;
  assign new_U220 = ~P2_DATAO_REG_29_ | ~new_U130;
  assign new_U221 = ~new_R140_U94 | ~new_U127;
  assign new_U222 = ~P2_DATAO_REG_28_ | ~new_U130;
  assign new_U223 = ~new_R140_U95 | ~new_U127;
  assign new_U224 = ~P2_DATAO_REG_27_ | ~new_U130;
  assign new_U225 = ~new_R140_U96 | ~new_U127;
  assign new_U226 = ~P2_DATAO_REG_26_ | ~new_U130;
  assign new_U227 = ~new_R140_U97 | ~new_U127;
  assign new_U228 = ~P2_DATAO_REG_25_ | ~new_U130;
  assign new_U229 = ~new_R140_U98 | ~new_U127;
  assign new_U230 = ~P2_DATAO_REG_24_ | ~new_U130;
  assign new_U231 = ~new_R140_U99 | ~new_U127;
  assign new_U232 = ~P2_DATAO_REG_23_ | ~new_U130;
  assign new_U233 = ~new_R140_U100 | ~new_U127;
  assign new_U234 = ~P2_DATAO_REG_22_ | ~new_U130;
  assign new_U235 = ~new_R140_U101 | ~new_U127;
  assign new_U236 = ~P2_DATAO_REG_21_ | ~new_U130;
  assign new_U237 = ~new_R140_U102 | ~new_U127;
  assign new_U238 = ~P2_DATAO_REG_20_ | ~new_U130;
  assign new_U239 = ~new_R140_U10 | ~new_U127;
  assign new_U240 = ~P2_DATAO_REG_1_ | ~new_U130;
  assign new_U241 = ~new_R140_U103 | ~new_U127;
  assign new_U242 = ~P2_DATAO_REG_19_ | ~new_U130;
  assign new_U243 = ~new_R140_U104 | ~new_U127;
  assign new_U244 = ~P2_DATAO_REG_18_ | ~new_U130;
  assign new_U245 = ~new_R140_U105 | ~new_U127;
  assign new_U246 = ~P2_DATAO_REG_17_ | ~new_U130;
  assign new_U247 = ~new_R140_U106 | ~new_U127;
  assign new_U248 = ~P2_DATAO_REG_16_ | ~new_U130;
  assign new_U249 = ~new_R140_U107 | ~new_U127;
  assign new_U250 = ~P2_DATAO_REG_15_ | ~new_U130;
  assign new_U251 = ~new_R140_U108 | ~new_U127;
  assign new_U252 = ~P2_DATAO_REG_14_ | ~new_U130;
  assign new_U253 = ~new_R140_U109 | ~new_U127;
  assign new_U254 = ~P2_DATAO_REG_13_ | ~new_U130;
  assign new_U255 = ~new_R140_U110 | ~new_U127;
  assign new_U256 = ~P2_DATAO_REG_12_ | ~new_U130;
  assign new_U257 = ~new_R140_U111 | ~new_U127;
  assign new_U258 = ~P2_DATAO_REG_11_ | ~new_U130;
  assign new_U259 = ~new_R140_U112 | ~new_U127;
  assign new_U260 = ~P2_DATAO_REG_10_ | ~new_U130;
  assign new_U261 = ~new_R140_U83 | ~new_U127;
  assign new_U262 = ~P2_DATAO_REG_0_ | ~new_U130;
  assign new_U263 = ~P2_DATAO_REG_9_ | ~new_U127;
  assign new_U264 = ~new_U130 | ~P1_DATAO_REG_9_;
  assign new_U265 = ~P2_DATAO_REG_8_ | ~new_U127;
  assign new_U266 = ~P1_DATAO_REG_8_ | ~new_U130;
  assign new_U267 = ~P2_DATAO_REG_7_ | ~new_U127;
  assign new_U268 = ~P1_DATAO_REG_7_ | ~new_U130;
  assign new_U269 = ~P2_DATAO_REG_6_ | ~new_U127;
  assign new_U270 = ~P1_DATAO_REG_6_ | ~new_U130;
  assign new_U271 = ~P2_DATAO_REG_5_ | ~new_U127;
  assign new_U272 = ~P1_DATAO_REG_5_ | ~new_U130;
  assign new_U273 = ~P2_DATAO_REG_4_ | ~new_U127;
  assign new_U274 = ~P1_DATAO_REG_4_ | ~new_U130;
  assign new_U275 = ~P2_DATAO_REG_31_ | ~new_U127;
  assign new_U276 = ~P1_DATAO_REG_31_ | ~new_U130;
  assign new_U277 = ~P2_DATAO_REG_30_ | ~new_U127;
  assign new_U278 = ~P1_DATAO_REG_30_ | ~new_U130;
  assign new_U279 = ~P2_DATAO_REG_3_ | ~new_U127;
  assign new_U280 = ~P1_DATAO_REG_3_ | ~new_U130;
  assign new_U281 = ~P2_DATAO_REG_29_ | ~new_U127;
  assign new_U282 = ~P1_DATAO_REG_29_ | ~new_U130;
  assign new_U283 = ~P2_DATAO_REG_28_ | ~new_U127;
  assign new_U284 = ~P1_DATAO_REG_28_ | ~new_U130;
  assign new_U285 = ~P2_DATAO_REG_27_ | ~new_U127;
  assign new_U286 = ~P1_DATAO_REG_27_ | ~new_U130;
  assign new_U287 = ~P2_DATAO_REG_26_ | ~new_U127;
  assign new_U288 = ~P1_DATAO_REG_26_ | ~new_U130;
  assign new_U289 = ~P2_DATAO_REG_25_ | ~new_U127;
  assign new_U290 = ~P1_DATAO_REG_25_ | ~new_U130;
  assign new_U291 = ~P2_DATAO_REG_24_ | ~new_U127;
  assign new_U292 = ~P1_DATAO_REG_24_ | ~new_U130;
  assign new_U293 = ~P2_DATAO_REG_23_ | ~new_U127;
  assign new_U294 = ~P1_DATAO_REG_23_ | ~new_U130;
  assign new_U295 = ~P2_DATAO_REG_22_ | ~new_U127;
  assign new_U296 = ~P1_DATAO_REG_22_ | ~new_U130;
  assign new_U297 = ~P2_DATAO_REG_21_ | ~new_U127;
  assign new_U298 = ~P1_DATAO_REG_21_ | ~new_U130;
  assign new_U299 = ~P2_DATAO_REG_20_ | ~new_U127;
  assign new_U300 = ~P1_DATAO_REG_20_ | ~new_U130;
  assign new_U301 = ~P2_DATAO_REG_2_ | ~new_U127;
  assign new_U302 = ~P1_DATAO_REG_2_ | ~new_U130;
  assign new_U303 = ~P2_DATAO_REG_19_ | ~new_U127;
  assign new_U304 = ~P1_DATAO_REG_19_ | ~new_U130;
  assign new_U305 = ~P2_DATAO_REG_18_ | ~new_U127;
  assign new_U306 = ~P1_DATAO_REG_18_ | ~new_U130;
  assign new_U307 = ~P2_DATAO_REG_17_ | ~new_U127;
  assign new_U308 = ~P1_DATAO_REG_17_ | ~new_U130;
  assign new_U309 = ~P2_DATAO_REG_16_ | ~new_U127;
  assign new_U310 = ~P1_DATAO_REG_16_ | ~new_U130;
  assign new_U311 = ~P2_DATAO_REG_15_ | ~new_U127;
  assign new_U312 = ~P1_DATAO_REG_15_ | ~new_U130;
  assign new_U313 = ~P2_DATAO_REG_14_ | ~new_U127;
  assign new_U314 = ~P1_DATAO_REG_14_ | ~new_U130;
  assign new_U315 = ~P2_DATAO_REG_13_ | ~new_U127;
  assign new_U316 = ~P1_DATAO_REG_13_ | ~new_U130;
  assign new_U317 = ~P2_DATAO_REG_12_ | ~new_U127;
  assign new_U318 = ~P1_DATAO_REG_12_ | ~new_U130;
  assign new_U319 = ~P2_DATAO_REG_11_ | ~new_U127;
  assign new_U320 = ~P1_DATAO_REG_11_ | ~new_U130;
  assign new_U321 = ~P2_DATAO_REG_10_ | ~new_U127;
  assign new_U322 = ~P1_DATAO_REG_10_ | ~new_U130;
  assign new_U323 = ~P2_DATAO_REG_1_ | ~new_U127;
  assign new_U324 = ~P1_DATAO_REG_1_ | ~new_U130;
  assign new_U325 = ~P2_DATAO_REG_0_ | ~new_U127;
  assign new_U326 = ~P1_DATAO_REG_0_ | ~new_U130;
  assign new_P2_R1161_U501 = ~new_P2_U3061 | ~new_P2_R1161_U63;
  assign new_P2_R1161_U500 = ~new_P2_R1161_U244 | ~new_P2_R1161_U498;
  assign new_P2_R1161_U499 = ~new_P2_R1161_U363 | ~new_P2_R1161_U167;
  assign new_P2_R1161_U498 = ~new_P2_R1161_U497 | ~new_P2_R1161_U496;
  assign new_P2_R1161_U497 = ~new_P2_U3422 | ~new_P2_R1161_U67;
  assign new_P2_R1161_U496 = ~new_P2_U3062 | ~new_P2_R1161_U66;
  assign new_P2_R1161_U495 = ~new_P2_R1161_U493 | ~new_P2_R1161_U338;
  assign new_P2_R1161_U494 = ~new_P2_R1161_U362 | ~new_P2_R1161_U93;
  assign new_P2_R1161_U493 = ~new_P2_R1161_U492 | ~new_P2_R1161_U491;
  assign new_P2_R1161_U492 = ~new_P2_U3425 | ~new_P2_R1161_U70;
  assign new_P2_R1161_U491 = ~new_P2_U3071 | ~new_P2_R1161_U69;
  assign new_P2_R1161_U490 = ~new_P2_U3428 | ~new_P2_R1161_U62;
  assign new_P1_U3014 = new_P1_U3956 & new_P1_U3443;
  assign new_P1_U3015 = new_P1_U3449 & new_P1_U3446;
  assign new_P1_U3016 = new_P1_U3630 & new_P1_U3625;
  assign new_P1_U3017 = new_P1_U3444 & new_P1_U3445;
  assign new_P1_U3018 = new_P1_U5711 & new_P1_U3444;
  assign new_P1_U3019 = new_P1_U5708 & new_P1_U3445;
  assign new_P1_U3020 = new_P1_U5708 & new_P1_U5711;
  assign new_P1_U3021 = new_P1_U5368 & new_P1_U3421;
  assign new_P1_U3022 = new_P1_U3046 & P1_STATE_REG;
  assign new_P1_U3023 = new_P1_U3049 & new_P1_U5690;
  assign new_P1_U3024 = new_P1_U3807 & new_P1_U3423;
  assign new_P1_U3025 = new_P1_U3987 & new_P1_U5699;
  assign new_P1_U3026 = new_P1_U3953 & new_P1_U5690;
  assign new_P1_U3027 = new_P1_U3871 & new_P1_U3972;
  assign new_P1_U3028 = new_P1_U3357 & P1_STATE_REG;
  assign new_P1_U3029 = new_P1_U3964 & new_P1_U3989;
  assign new_P1_U3030 = new_P1_U3989 & new_P1_U3422;
  assign new_P1_U3031 = new_P1_U3957 & new_P1_U3989;
  assign new_P1_U3032 = new_P1_U3965 & new_P1_U3989;
  assign new_P1_U3033 = new_P1_U3987 & new_P1_U3446;
  assign new_P1_U3034 = new_P1_U3972 & new_P1_U5699;
  assign new_P1_U3035 = new_P1_U3989 & new_P1_U3025;
  assign new_P1_U3036 = new_P1_U3972 & new_P1_U3446;
  assign new_P1_U3037 = new_P1_U5702 & new_P1_U4880;
  assign new_P1_U3038 = new_P1_U3024 & new_P1_U5702;
  assign new_P1_U3039 = new_P1_U5699 & new_P1_U4880;
  assign new_P1_U3040 = new_P1_U3024 & new_P1_U5699;
  assign new_P1_U3041 = new_P1_U3015 & new_P1_U4880;
  assign new_P1_U3042 = new_P1_U3024 & new_P1_U3015;
  assign new_P1_U3043 = new_P1_U3022 & new_P1_U3423;
  assign new_P1_U3044 = new_P1_U5113 & P1_STATE_REG;
  assign new_P1_U3045 = new_P1_U3022 & new_P1_U5115;
  assign new_P1_U3046 = new_P1_U5677 & new_P1_U3421;
  assign new_P1_U3047 = new_P1_U3631 & new_P1_U3016;
  assign new_P1_U3048 = new_P1_U5690 & new_P1_U3442;
  assign new_P1_U3049 = new_P1_U5684 & new_P1_U5693;
  assign new_P1_U3050 = new_P1_U3435 & new_P1_U3437;
  assign new_P1_U3051 = new_P1_U4699 & new_P1_U4700 & new_P1_U4706 & new_P1_U4703;
  assign new_P1_U3052 = new_P1_U6070 & new_P1_U6069;
  assign new_P1_U3053 = ~new_P1_U4639 | ~new_P1_U4636 | ~new_P1_U4637 | ~new_P1_U4638;
  assign new_P1_U3054 = ~new_P1_U4658 | ~new_P1_U4655 | ~new_P1_U4656 | ~new_P1_U4657;
  assign new_P1_U3055 = ~new_P1_U4674 | ~new_P1_U4675 | ~new_P1_U4677 | ~new_P1_U4676;
  assign new_P1_U3056 = ~new_P1_U4713 | ~new_P1_U4714 | ~new_P1_U4715;
  assign new_P1_U3057 = ~new_P1_U4620 | ~new_P1_U4617 | ~new_P1_U4618 | ~new_P1_U4619;
  assign new_P1_U3058 = ~new_P1_U4601 | ~new_P1_U4598 | ~new_P1_U4599 | ~new_P1_U4600;
  assign new_P1_U3059 = ~new_P1_U4693 | ~new_P1_U4694 | ~new_P1_U4695;
  assign new_P1_U3060 = ~new_P1_U4199 | ~new_P1_U4200 | ~new_P1_U4202 | ~new_P1_U4201;
  assign new_P1_U3061 = ~new_P1_U4544 | ~new_P1_U4541 | ~new_P1_U4542 | ~new_P1_U4543;
  assign new_P1_U3062 = ~new_P1_U4316 | ~new_P1_U4313 | ~new_P1_U4314 | ~new_P1_U4315;
  assign new_P1_U3063 = ~new_P1_U4335 | ~new_P1_U4332 | ~new_P1_U4333 | ~new_P1_U4334;
  assign new_P1_U3064 = ~new_P1_U4180 | ~new_P1_U4181 | ~new_P1_U4183 | ~new_P1_U4182;
  assign new_P1_U3065 = ~new_P1_U4582 | ~new_P1_U4579 | ~new_P1_U4580 | ~new_P1_U4581;
  assign new_P1_U3066 = ~new_P1_U4563 | ~new_P1_U4560 | ~new_P1_U4561 | ~new_P1_U4562;
  assign new_P1_U3067 = ~new_P1_U4218 | ~new_P1_U4219 | ~new_P1_U4221 | ~new_P1_U4220;
  assign new_P1_U3068 = ~new_P1_U4156 | ~new_P1_U4157 | ~new_P1_U4159 | ~new_P1_U4158;
  assign new_P1_U3069 = ~new_P1_U4449 | ~new_P1_U4446 | ~new_P1_U4447 | ~new_P1_U4448;
  assign new_P1_U3070 = ~new_P1_U4256 | ~new_P1_U4257 | ~new_P1_U4259 | ~new_P1_U4258;
  assign new_P1_U3071 = ~new_P1_U4237 | ~new_P1_U4238 | ~new_P1_U4240 | ~new_P1_U4239;
  assign new_P1_U3072 = ~new_P1_U4354 | ~new_P1_U4351 | ~new_P1_U4352 | ~new_P1_U4353;
  assign new_P1_U3073 = ~new_P1_U4430 | ~new_P1_U4427 | ~new_P1_U4428 | ~new_P1_U4429;
  assign new_P1_U3074 = ~new_P1_U4411 | ~new_P1_U4408 | ~new_P1_U4409 | ~new_P1_U4410;
  assign new_P1_U3075 = ~new_P1_U4525 | ~new_P1_U4522 | ~new_P1_U4523 | ~new_P1_U4524;
  assign new_P1_U3076 = ~new_P1_U4506 | ~new_P1_U4503 | ~new_P1_U4504 | ~new_P1_U4505;
  assign new_P1_U3077 = ~new_P1_U4161 | ~new_P1_U4162 | ~new_P1_U4164 | ~new_P1_U4163;
  assign new_P1_U3078 = ~new_P1_U4137 | ~new_P1_U4138 | ~new_P1_U4140 | ~new_P1_U4139;
  assign new_P1_U3079 = ~new_P1_U4392 | ~new_P1_U4389 | ~new_P1_U4390 | ~new_P1_U4391;
  assign new_P1_U3080 = ~new_P1_U4373 | ~new_P1_U4370 | ~new_P1_U4371 | ~new_P1_U4372;
  assign new_P1_U3081 = ~new_P1_U4487 | ~new_P1_U4484 | ~new_P1_U4485 | ~new_P1_U4486;
  assign new_P1_U3082 = ~new_P1_U4468 | ~new_P1_U4465 | ~new_P1_U4466 | ~new_P1_U4467;
  assign new_P1_U3083 = ~new_P1_U4297 | ~new_P1_U4294 | ~new_P1_U4295 | ~new_P1_U4296;
  assign new_P1_U3084 = ~new_P1_U4275 | ~new_P1_U4276 | ~new_P1_U4278 | ~new_P1_U4277;
  assign n1335 = ~new_P1_U4887 | ~P1_STATE_REG;
  assign n1330 = ~P1_STATE_REG;
  assign new_P1_U3087 = ~new_P1_U5576 | ~new_P1_U5575;
  assign new_P1_U3088 = ~new_P1_U5578 | ~new_P1_U5577;
  assign new_P1_U3089 = ~new_P1_U5582 | ~new_P1_U5583 | ~new_P1_U5584;
  assign new_P1_U3090 = ~new_P1_U3895 | ~new_P1_U5586;
  assign new_P1_U3091 = ~new_P1_U3896 | ~new_P1_U5589;
  assign new_P1_U3092 = ~new_P1_U3897 | ~new_P1_U5592;
  assign new_P1_U3093 = ~new_P1_U3898 | ~new_P1_U5595;
  assign new_P1_U3094 = ~new_P1_U3899 | ~new_P1_U5598;
  assign new_P1_U3095 = ~new_P1_U3900 | ~new_P1_U5601;
  assign new_P1_U3096 = ~new_P1_U3901 | ~new_P1_U5604;
  assign new_P1_U3097 = ~new_P1_U3902 | ~new_P1_U5607;
  assign new_P1_U3098 = ~new_P1_U3903 | ~new_P1_U5610;
  assign new_P1_U3099 = ~new_P1_U3904 | ~new_P1_U5616;
  assign new_P1_U3100 = ~new_P1_U3905 | ~new_P1_U5619;
  assign new_P1_U3101 = ~new_P1_U3906 | ~new_P1_U5622;
  assign new_P1_U3102 = ~new_P1_U3907 | ~new_P1_U5625;
  assign new_P1_U3103 = ~new_P1_U3908 | ~new_P1_U5628;
  assign new_P1_U3104 = ~new_P1_U3909 | ~new_P1_U5631;
  assign new_P1_U3105 = ~new_P1_U5633 | ~new_P1_U5634 | ~new_P1_U5635;
  assign new_P1_U3106 = ~new_P1_U5636 | ~new_P1_U5637 | ~new_P1_U5638;
  assign new_P1_U3107 = ~new_P1_U5639 | ~new_P1_U5640 | ~new_P1_U5641;
  assign new_P1_U3108 = ~new_P1_U5642 | ~new_P1_U5643 | ~new_P1_U5644;
  assign new_P1_U3109 = ~new_P1_U5557 | ~new_P1_U5558 | ~new_P1_U5559;
  assign new_P1_U3110 = ~new_P1_U5560 | ~new_P1_U5561 | ~new_P1_U5562;
  assign new_P1_U3111 = ~new_P1_U5563 | ~new_P1_U5564 | ~new_P1_U5565;
  assign new_P1_U3112 = ~new_P1_U5566 | ~new_P1_U5567 | ~new_P1_U5568;
  assign new_P1_U3113 = ~new_P1_U5569 | ~new_P1_U5570 | ~new_P1_U5571;
  assign new_P1_U3114 = ~new_P1_U5572 | ~new_P1_U5573 | ~new_P1_U5574;
  assign new_P1_U3115 = ~new_P1_U5579 | ~new_P1_U5580 | ~new_P1_U5581;
  assign new_P1_U3116 = ~new_P1_U5612 | ~new_P1_U5613 | ~new_P1_U5614;
  assign new_P1_U3117 = ~new_P1_U5645 | ~new_P1_U5646 | ~new_P1_U5647;
  assign new_P1_U3118 = ~new_P1_U5649 | ~new_P1_U5648;
  assign new_P1_U3119 = ~new_P1_U5506 | ~new_P1_U5505;
  assign new_P1_U3120 = ~new_P1_U5508 | ~new_P1_U5507;
  assign new_P1_U3121 = ~new_P1_U5512 | ~new_P1_U3438 | ~new_P1_U5511;
  assign new_P1_U3122 = ~new_P1_U3879 | ~new_P1_U5513;
  assign new_P1_U3123 = ~new_P1_U3880 | ~new_P1_U5515;
  assign new_P1_U3124 = ~new_P1_U3881 | ~new_P1_U5517;
  assign new_P1_U3125 = ~new_P1_U3882 | ~new_P1_U5519;
  assign new_P1_U3126 = ~new_P1_U3883 | ~new_P1_U5521;
  assign new_P1_U3127 = ~new_P1_U3884 | ~new_P1_U5523;
  assign new_P1_U3128 = ~new_P1_U3885 | ~new_P1_U5525;
  assign new_P1_U3129 = ~new_P1_U3886 | ~new_P1_U5527;
  assign new_P1_U3130 = ~new_P1_U3887 | ~new_P1_U5529;
  assign new_P1_U3131 = ~new_P1_U3888 | ~new_P1_U5534;
  assign new_P1_U3132 = ~new_P1_U3889 | ~new_P1_U5536;
  assign new_P1_U3133 = ~new_P1_U3890 | ~new_P1_U5538;
  assign new_P1_U3134 = ~new_P1_U3891 | ~new_P1_U5540;
  assign new_P1_U3135 = ~new_P1_U3892 | ~new_P1_U5542;
  assign new_P1_U3136 = ~new_P1_U3893 | ~new_P1_U5544;
  assign new_P1_U3137 = ~new_P1_U5545 | ~new_P1_U5546 | ~new_P1_U3438;
  assign new_P1_U3138 = ~new_P1_U5547 | ~new_P1_U5548 | ~new_P1_U3438;
  assign new_P1_U3139 = ~new_P1_U5549 | ~new_P1_U5550 | ~new_P1_U3438;
  assign new_P1_U3140 = ~new_P1_U5551 | ~new_P1_U5552 | ~new_P1_U3438;
  assign new_P1_U3141 = ~new_P1_U5493 | ~new_P1_U5494 | ~new_P1_U3438;
  assign new_P1_U3142 = ~new_P1_U5495 | ~new_P1_U5496 | ~new_P1_U3438;
  assign new_P1_U3143 = ~new_P1_U5497 | ~new_P1_U5498 | ~new_P1_U3438;
  assign new_P1_U3144 = ~new_P1_U5499 | ~new_P1_U5500 | ~new_P1_U3438;
  assign new_P1_U3145 = ~new_P1_U5501 | ~new_P1_U5502 | ~new_P1_U3438;
  assign new_P1_U3146 = ~new_P1_U5503 | ~new_P1_U5504 | ~new_P1_U3438;
  assign new_P1_U3147 = ~new_P1_U5509 | ~new_P1_U5510 | ~new_P1_U3438;
  assign new_P1_U3148 = ~new_P1_U5531 | ~new_P1_U5532 | ~new_P1_U3438;
  assign new_P1_U3149 = ~new_P1_U5553 | ~new_P1_U5554 | ~new_P1_U3438;
  assign new_P1_U3150 = ~new_P1_U3894 | ~new_P1_U5556;
  assign new_P1_U3151 = ~new_P1_U3953 | ~new_P1_U3438;
  assign new_P1_U3152 = ~new_P1_U5677 | ~new_P1_U3372;
  assign new_P1_U3153 = ~new_P1_U5448 | ~new_P1_U5447;
  assign new_P1_U3154 = ~new_P1_U5450 | ~new_P1_U5449;
  assign new_P1_U3155 = ~new_P1_U5452 | ~new_P1_U5451;
  assign new_P1_U3156 = ~new_P1_U5454 | ~new_P1_U5453;
  assign new_P1_U3157 = ~new_P1_U5456 | ~new_P1_U5455;
  assign new_P1_U3158 = ~new_P1_U5458 | ~new_P1_U5457;
  assign new_P1_U3159 = ~new_P1_U5460 | ~new_P1_U5459;
  assign new_P1_U3160 = ~new_P1_U5462 | ~new_P1_U5461;
  assign new_P1_U3161 = ~new_P1_U5464 | ~new_P1_U5463;
  assign new_P1_U3162 = ~new_P1_U5468 | ~new_P1_U5467;
  assign new_P1_U3163 = ~new_P1_U5470 | ~new_P1_U5469;
  assign new_P1_U3164 = ~new_P1_U5472 | ~new_P1_U5471;
  assign new_P1_U3165 = ~new_P1_U5474 | ~new_P1_U5473;
  assign new_P1_U3166 = ~new_P1_U5476 | ~new_P1_U5475;
  assign new_P1_U3167 = ~new_P1_U5478 | ~new_P1_U5477;
  assign new_P1_U3168 = ~new_P1_U5480 | ~new_P1_U5479;
  assign new_P1_U3169 = ~new_P1_U5482 | ~new_P1_U5481;
  assign new_P1_U3170 = ~new_P1_U5484 | ~new_P1_U5483;
  assign new_P1_U3171 = ~new_P1_U5486 | ~new_P1_U5485;
  assign new_P1_U3172 = ~new_P1_U5434 | ~new_P1_U5433;
  assign new_P1_U3173 = ~new_P1_U5436 | ~new_P1_U5435;
  assign new_P1_U3174 = ~new_P1_U5438 | ~new_P1_U5437;
  assign new_P1_U3175 = ~new_P1_U5440 | ~new_P1_U5439;
  assign new_P1_U3176 = ~new_P1_U5442 | ~new_P1_U5441;
  assign new_P1_U3177 = ~new_P1_U5444 | ~new_P1_U5443;
  assign new_P1_U3178 = ~new_P1_U5446 | ~new_P1_U5445;
  assign new_P1_U3179 = ~new_P1_U5466 | ~new_P1_U5465;
  assign new_P1_U3180 = ~new_P1_U5488 | ~new_P1_U5487;
  assign new_P1_U3181 = ~new_P1_U5489 | ~new_P1_U5490 | ~new_P1_U5491;
  assign new_P1_U3182 = ~new_P1_U5389 | ~new_P1_U5388;
  assign new_P1_U3183 = ~new_P1_U5391 | ~new_P1_U5390;
  assign new_P1_U3184 = ~new_P1_U5393 | ~new_P1_U5392;
  assign new_P1_U3185 = ~new_P1_U5395 | ~new_P1_U5394;
  assign new_P1_U3186 = ~new_P1_U5397 | ~new_P1_U5396;
  assign new_P1_U3187 = ~new_P1_U5399 | ~new_P1_U5398;
  assign new_P1_U3188 = ~new_P1_U5401 | ~new_P1_U5400;
  assign new_P1_U3189 = ~new_P1_U5403 | ~new_P1_U5402;
  assign new_P1_U3190 = ~new_P1_U5405 | ~new_P1_U5404;
  assign new_P1_U3191 = ~new_P1_U5409 | ~new_P1_U5408;
  assign new_P1_U3192 = ~new_P1_U5411 | ~new_P1_U5410;
  assign new_P1_U3193 = ~new_P1_U5413 | ~new_P1_U5412;
  assign new_P1_U3194 = ~new_P1_U5415 | ~new_P1_U5414;
  assign new_P1_U3195 = ~new_P1_U5417 | ~new_P1_U5416;
  assign new_P1_U3196 = ~new_P1_U5419 | ~new_P1_U5418;
  assign new_P1_U3197 = ~new_P1_U5421 | ~new_P1_U5420;
  assign new_P1_U3198 = ~new_P1_U5423 | ~new_P1_U5422;
  assign new_P1_U3199 = ~new_P1_U5425 | ~new_P1_U5424;
  assign new_P1_U3200 = ~new_P1_U5427 | ~new_P1_U5426;
  assign new_P1_U3201 = ~new_P1_U5375 | ~new_P1_U5374;
  assign new_P1_U3202 = ~new_P1_U5377 | ~new_P1_U5376;
  assign new_P1_U3203 = ~new_P1_U5379 | ~new_P1_U5378;
  assign new_P1_U3204 = ~new_P1_U5381 | ~new_P1_U5380;
  assign new_P1_U3205 = ~new_P1_U5383 | ~new_P1_U5382;
  assign new_P1_U3206 = ~new_P1_U5385 | ~new_P1_U5384;
  assign new_P1_U3207 = ~new_P1_U5387 | ~new_P1_U5386;
  assign new_P1_U3208 = ~new_P1_U5407 | ~new_P1_U5406;
  assign new_P1_U3209 = ~new_P1_U5429 | ~new_P1_U5428;
  assign new_P1_U3210 = ~new_P1_U3878 | ~new_P1_U5430;
  assign new_P1_U3211 = new_P1_U5367 & new_P1_U3421;
  assign new_P1_U3212 = ~new_P1_U5365 | ~new_P1_U6236 | ~new_P1_U6235;
  assign n1325 = ~new_P1_U5361 | ~new_P1_U5360 | ~new_P1_U5362 | ~new_P1_U5359 | ~new_P1_U5358;
  assign n1320 = ~new_P1_U5352 | ~new_P1_U5351 | ~new_P1_U5353 | ~new_P1_U5350 | ~new_P1_U5349;
  assign n1315 = ~new_P1_U5343 | ~new_P1_U5342 | ~new_P1_U5344 | ~new_P1_U5341 | ~new_P1_U5340;
  assign n1310 = ~new_P1_U5334 | ~new_P1_U5333 | ~new_P1_U5335 | ~new_P1_U5332 | ~new_P1_U5331;
  assign n1305 = ~new_P1_U5325 | ~new_P1_U5324 | ~new_P1_U5326 | ~new_P1_U5323 | ~new_P1_U5322;
  assign n1300 = ~new_P1_U5316 | ~new_P1_U5315 | ~new_P1_U5317 | ~new_P1_U5314 | ~new_P1_U5313;
  assign n1295 = ~new_P1_U5307 | ~new_P1_U5306 | ~new_P1_U5308 | ~new_P1_U5305 | ~new_P1_U5304;
  assign n1290 = ~new_P1_U5298 | ~new_P1_U5297 | ~new_P1_U5299 | ~new_P1_U5296 | ~new_P1_U5295;
  assign n1285 = ~new_P1_U5289 | ~new_P1_U5288 | ~new_P1_U5290 | ~new_P1_U5287 | ~new_P1_U5286;
  assign n1280 = ~new_P1_U5279 | ~new_P1_U3876 | ~new_P1_U5278 | ~new_P1_U5277;
  assign n1275 = ~new_P1_U5271 | ~new_P1_U5270 | ~new_P1_U5272 | ~new_P1_U5269 | ~new_P1_U5268;
  assign n1270 = ~new_P1_U5262 | ~new_P1_U5261 | ~new_P1_U5263 | ~new_P1_U5260 | ~new_P1_U5259;
  assign n1265 = ~new_P1_U5253 | ~new_P1_U5252 | ~new_P1_U5254 | ~new_P1_U5251 | ~new_P1_U5250;
  assign n1260 = ~new_P1_U5244 | ~new_P1_U5243 | ~new_P1_U5245 | ~new_P1_U5242 | ~new_P1_U5241;
  assign n1255 = ~new_P1_U5235 | ~new_P1_U5234 | ~new_P1_U5236 | ~new_P1_U5233 | ~new_P1_U5232;
  assign n1250 = ~new_P1_U5226 | ~new_P1_U5225 | ~new_P1_U5227 | ~new_P1_U5224 | ~new_P1_U5223;
  assign n1245 = ~new_P1_U5217 | ~new_P1_U5216 | ~new_P1_U5218 | ~new_P1_U5215 | ~new_P1_U5214;
  assign n1240 = ~new_P1_U5208 | ~new_P1_U5207 | ~new_P1_U5209 | ~new_P1_U5206 | ~new_P1_U5205;
  assign n1235 = ~new_P1_U5199 | ~new_P1_U5198 | ~new_P1_U5200 | ~new_P1_U5197 | ~new_P1_U5196;
  assign n1230 = ~new_P1_U3874 | ~new_P1_U3875 | ~new_P1_U5189;
  assign n1225 = ~new_P1_U5182 | ~new_P1_U5181 | ~new_P1_U5183 | ~new_P1_U5180 | ~new_P1_U5179;
  assign n1220 = ~new_P1_U5173 | ~new_P1_U5172 | ~new_P1_U5174 | ~new_P1_U5171 | ~new_P1_U5170;
  assign n1215 = ~new_P1_U5164 | ~new_P1_U5163 | ~new_P1_U5165 | ~new_P1_U5162 | ~new_P1_U5161;
  assign n1210 = ~new_P1_U5155 | ~new_P1_U5154 | ~new_P1_U5156 | ~new_P1_U5153 | ~new_P1_U5152;
  assign n1205 = ~new_P1_U3872 | ~new_P1_U5145 | ~new_P1_U5144 | ~new_P1_U5143;
  assign n1200 = ~new_P1_U5137 | ~new_P1_U5136 | ~new_P1_U5138 | ~new_P1_U5135 | ~new_P1_U5134;
  assign n1195 = ~new_P1_U5128 | ~new_P1_U5127 | ~new_P1_U5129 | ~new_P1_U5126 | ~new_P1_U5125;
  assign n1190 = ~new_P1_U5119 | ~new_P1_U5118 | ~new_P1_U5120 | ~new_P1_U5117 | ~new_P1_U5116;
  assign n1185 = ~new_P1_U5106 | ~new_P1_U5105 | ~new_P1_U5107 | ~new_P1_U5104 | ~new_P1_U5103;
  assign n1180 = new_P1_U3866 & new_P1_U5650;
  assign n1015 = ~new_P1_U3849 | ~new_P1_U3848;
  assign n1010 = ~new_P1_U3847 | ~new_P1_U3846;
  assign n1005 = ~new_P1_U3845 | ~new_P1_U3844;
  assign n1000 = ~new_P1_U3842 | ~new_P1_U3841;
  assign n995 = ~new_P1_U3840 | ~new_P1_U3839;
  assign n990 = ~new_P1_U3837 | ~new_P1_U3836;
  assign n985 = ~new_P1_U3835 | ~new_P1_U3834;
  assign n980 = ~new_P1_U5010 | ~new_P1_U3832 | ~new_P1_U3833;
  assign n975 = ~new_P1_U5000 | ~new_P1_U3830 | ~new_P1_U3831;
  assign n970 = ~new_P1_U4990 | ~new_P1_U3828 | ~new_P1_U3829;
  assign n965 = ~new_P1_U4980 | ~new_P1_U3826 | ~new_P1_U3827;
  assign n960 = ~new_P1_U4970 | ~new_P1_U3824 | ~new_P1_U3825;
  assign n955 = ~new_P1_U4960 | ~new_P1_U3822 | ~new_P1_U3823;
  assign n950 = ~new_P1_U4950 | ~new_P1_U3820 | ~new_P1_U3821;
  assign n945 = ~new_P1_U4940 | ~new_P1_U3818 | ~new_P1_U3819;
  assign n940 = ~new_P1_U4930 | ~new_P1_U3816 | ~new_P1_U3817;
  assign n935 = ~new_P1_U4920 | ~new_P1_U3814 | ~new_P1_U3815;
  assign n930 = ~new_P1_U4910 | ~new_P1_U3812 | ~new_P1_U3813;
  assign n925 = ~new_P1_U4900 | ~new_P1_U3810 | ~new_P1_U3811;
  assign n920 = ~new_P1_U4890 | ~new_P1_U3808 | ~new_P1_U3809;
  assign n915 = ~new_P1_U4879 | ~new_P1_U3947 | ~new_P1_U4878;
  assign n910 = ~new_P1_U4877 | ~new_P1_U3946 | ~new_P1_U4876;
  assign n900 = ~new_P1_U3943 | ~new_P1_U4869 | ~new_P1_U3799 | ~new_P1_U3800;
  assign n895 = ~new_P1_U3942 | ~new_P1_U4864 | ~new_P1_U3797 | ~new_P1_U3798;
  assign n890 = ~new_P1_U3941 | ~new_P1_U4859 | ~new_P1_U3795 | ~new_P1_U3796;
  assign n885 = ~new_P1_U3940 | ~new_P1_U4854 | ~new_P1_U3793 | ~new_P1_U3794;
  assign n880 = ~new_P1_U3939 | ~new_P1_U4849 | ~new_P1_U3791 | ~new_P1_U3792;
  assign n875 = ~new_P1_U3938 | ~new_P1_U3790 | ~new_P1_U3789;
  assign n870 = ~new_P1_U3937 | ~new_P1_U3788 | ~new_P1_U3787;
  assign n865 = ~new_P1_U3786 | ~new_P1_U3936;
  assign n860 = ~new_P1_U3935 | ~new_P1_U3785 | ~new_P1_U3784;
  assign n855 = ~new_P1_U3783 | ~new_P1_U3934;
  assign n850 = ~new_P1_U3782 | ~new_P1_U3933;
  assign n845 = ~new_P1_U3781 | ~new_P1_U3932;
  assign n840 = ~new_P1_U3780 | ~new_P1_U3931;
  assign n835 = ~new_P1_U3779 | ~new_P1_U3930;
  assign n830 = ~new_P1_U3778 | ~new_P1_U3929;
  assign n825 = ~new_P1_U3928 | ~new_P1_U3777 | ~new_P1_U3776;
  assign n820 = ~new_P1_U3927 | ~new_P1_U3775 | ~new_P1_U3774;
  assign n815 = ~new_P1_U3926 | ~new_P1_U3773 | ~new_P1_U3772;
  assign n810 = ~new_P1_U3925 | ~new_P1_U4779 | ~new_P1_U3770 | ~new_P1_U3771;
  assign n805 = ~new_P1_U3924 | ~new_P1_U4774 | ~new_P1_U3768 | ~new_P1_U3769;
  assign n800 = ~new_P1_U3923 | ~new_P1_U4769 | ~new_P1_U3766 | ~new_P1_U3767;
  assign n795 = ~new_P1_U3922 | ~new_P1_U4764 | ~new_P1_U3764 | ~new_P1_U3765;
  assign n790 = ~new_P1_U3921 | ~new_P1_U4759 | ~new_P1_U3762 | ~new_P1_U3763;
  assign n785 = ~new_P1_U3920 | ~new_P1_U4754 | ~new_P1_U3760 | ~new_P1_U3761;
  assign n780 = ~new_P1_U3919 | ~new_P1_U4749 | ~new_P1_U3758 | ~new_P1_U3759;
  assign n775 = ~new_P1_U3918 | ~new_P1_U3757 | ~new_P1_U3756;
  assign n770 = ~new_P1_U3755 | ~new_P1_U3754;
  assign n765 = ~new_P1_U3753 | ~new_P1_U3752;
  assign n760 = ~new_P1_U3751 | ~new_P1_U3750;
  assign n435 = P1_D_REG_31_ & new_P1_U3911;
  assign n430 = P1_D_REG_30_ & new_P1_U3911;
  assign n425 = P1_D_REG_29_ & new_P1_U3911;
  assign n420 = P1_D_REG_28_ & new_P1_U3911;
  assign n415 = P1_D_REG_27_ & new_P1_U3911;
  assign n410 = P1_D_REG_26_ & new_P1_U3911;
  assign n405 = P1_D_REG_25_ & new_P1_U3911;
  assign n400 = P1_D_REG_24_ & new_P1_U3911;
  assign n395 = P1_D_REG_23_ & new_P1_U3911;
  assign n390 = P1_D_REG_22_ & new_P1_U3911;
  assign n385 = P1_D_REG_21_ & new_P1_U3911;
  assign n380 = P1_D_REG_20_ & new_P1_U3911;
  assign n375 = P1_D_REG_19_ & new_P1_U3911;
  assign n370 = P1_D_REG_18_ & new_P1_U3911;
  assign n365 = P1_D_REG_17_ & new_P1_U3911;
  assign n360 = P1_D_REG_16_ & new_P1_U3911;
  assign n355 = P1_D_REG_15_ & new_P1_U3911;
  assign n350 = P1_D_REG_14_ & new_P1_U3911;
  assign n345 = P1_D_REG_13_ & new_P1_U3911;
  assign n340 = P1_D_REG_12_ & new_P1_U3911;
  assign n335 = P1_D_REG_11_ & new_P1_U3911;
  assign n330 = P1_D_REG_10_ & new_P1_U3911;
  assign n325 = P1_D_REG_9_ & new_P1_U3911;
  assign n320 = P1_D_REG_8_ & new_P1_U3911;
  assign n315 = P1_D_REG_7_ & new_P1_U3911;
  assign n310 = P1_D_REG_6_ & new_P1_U3911;
  assign n305 = P1_D_REG_5_ & new_P1_U3911;
  assign n300 = P1_D_REG_4_ & new_P1_U3911;
  assign n295 = P1_D_REG_3_ & new_P1_U3911;
  assign n290 = P1_D_REG_2_ & new_P1_U3911;
  assign n275 = ~new_P1_U4098 | ~new_P1_U4099 | ~new_P1_U4100;
  assign n270 = ~new_P1_U4095 | ~new_P1_U4096 | ~new_P1_U4097;
  assign n265 = ~new_P1_U4092 | ~new_P1_U4093 | ~new_P1_U4094;
  assign n260 = ~new_P1_U4089 | ~new_P1_U4090 | ~new_P1_U4091;
  assign n255 = ~new_P1_U4086 | ~new_P1_U4087 | ~new_P1_U4088;
  assign n250 = ~new_P1_U4083 | ~new_P1_U4084 | ~new_P1_U4085;
  assign n245 = ~new_P1_U4080 | ~new_P1_U4081 | ~new_P1_U4082;
  assign n240 = ~new_P1_U4077 | ~new_P1_U4078 | ~new_P1_U4079;
  assign n235 = ~new_P1_U4074 | ~new_P1_U4075 | ~new_P1_U4076;
  assign n230 = ~new_P1_U4071 | ~new_P1_U4072 | ~new_P1_U4073;
  assign n225 = ~new_P1_U4068 | ~new_P1_U4069 | ~new_P1_U4070;
  assign n220 = ~new_P1_U4065 | ~new_P1_U4066 | ~new_P1_U4067;
  assign n215 = ~new_P1_U4062 | ~new_P1_U4063 | ~new_P1_U4064;
  assign n210 = ~new_P1_U4059 | ~new_P1_U4060 | ~new_P1_U4061;
  assign n205 = ~new_P1_U4056 | ~new_P1_U4057 | ~new_P1_U4058;
  assign n200 = ~new_P1_U4053 | ~new_P1_U4054 | ~new_P1_U4055;
  assign n195 = ~new_P1_U4050 | ~new_P1_U4051 | ~new_P1_U4052;
  assign n190 = ~new_P1_U4047 | ~new_P1_U4048 | ~new_P1_U4049;
  assign n185 = ~new_P1_U4044 | ~new_P1_U4045 | ~new_P1_U4046;
  assign n180 = ~new_P1_U4041 | ~new_P1_U4042 | ~new_P1_U4043;
  assign n175 = ~new_P1_U4038 | ~new_P1_U4039 | ~new_P1_U4040;
  assign n170 = ~new_P1_U4035 | ~new_P1_U4036 | ~new_P1_U4037;
  assign n165 = ~new_P1_U4032 | ~new_P1_U4033 | ~new_P1_U4034;
  assign n160 = ~new_P1_U4029 | ~new_P1_U4030 | ~new_P1_U4031;
  assign n155 = ~new_P1_U4026 | ~new_P1_U4027 | ~new_P1_U4028;
  assign n150 = ~new_P1_U4023 | ~new_P1_U4024 | ~new_P1_U4025;
  assign n145 = ~new_P1_U4020 | ~new_P1_U4021 | ~new_P1_U4022;
  assign n140 = ~new_P1_U4017 | ~new_P1_U4018 | ~new_P1_U4019;
  assign n135 = ~new_P1_U4014 | ~new_P1_U4015 | ~new_P1_U4016;
  assign n130 = ~new_P1_U4011 | ~new_P1_U4012 | ~new_P1_U4013;
  assign n125 = ~new_P1_U4008 | ~new_P1_U4009 | ~new_P1_U4010;
  assign new_P1_U3355 = ~new_P1_U4005 | ~new_P1_U4006 | ~new_P1_U4007;
  assign n905 = ~new_P1_U3944 | ~new_P1_U4873 | ~new_P1_U4875 | ~new_P1_U4874 | ~new_P1_U4872;
  assign new_P1_U3357 = ~P1_STATE_REG | ~new_P1_U3910;
  assign new_P1_U3358 = ~new_P1_U3437 | ~new_P1_U5669;
  assign new_P1_U3359 = ~P1_B_REG;
  assign new_P1_U3360 = ~new_P1_U3437 | ~new_P1_U5674 | ~new_P1_U5673;
  assign new_P1_U3361 = ~new_P1_U3048 | ~new_P1_U3443;
  assign new_P1_U3362 = ~new_P1_U3443 | ~new_P1_U3441 | ~new_P1_U3442;
  assign new_P1_U3363 = ~new_P1_U3441 | ~new_P1_U5687;
  assign new_P1_U3364 = ~new_P1_U4001 | ~new_P1_U3443;
  assign new_P1_U3365 = ~new_P1_U3447 | ~new_P1_U3441 | ~new_P1_U3442;
  assign new_P1_U3366 = ~new_P1_U4001 | ~new_P1_U3447;
  assign new_P1_U3367 = ~new_P1_U5690 | ~new_P1_U5687;
  assign new_P1_U3368 = ~new_P1_U4002 | ~new_P1_U3443;
  assign new_P1_U3369 = ~new_P1_U3960 | ~new_P1_U5693;
  assign new_P1_U3370 = ~new_P1_U4002 | ~new_P1_U3447;
  assign new_P1_U3371 = ~new_P1_U3956 | ~new_P1_U5684;
  assign new_P1_U3372 = ~new_P1_U5684 | ~new_P1_U3442;
  assign new_P1_U3373 = ~new_P1_U3443 | ~new_P1_U3447;
  assign new_P1_U3374 = ~new_P1_U3618 | ~new_P1_U3619 | ~new_P1_U4149 | ~new_P1_U4148 | ~new_P1_U4147;
  assign new_P1_U3375 = ~P1_REG2_REG_0_;
  assign new_P1_U3376 = ~new_P1_U3635 | ~new_P1_U3633 | ~new_P1_U4167 | ~new_P1_U4166;
  assign new_P1_U3377 = ~new_P1_U3639 | ~new_P1_U3637 | ~new_P1_U4186 | ~new_P1_U4185;
  assign new_P1_U3378 = ~new_P1_U3642 | ~new_P1_U4207 | ~new_P1_U4206 | ~new_P1_U4205 | ~new_P1_U4204;
  assign new_P1_U3379 = ~new_P1_U3645 | ~new_P1_U4226 | ~new_P1_U4225 | ~new_P1_U4224 | ~new_P1_U4223;
  assign new_P1_U3380 = ~new_P1_U3649 | ~new_P1_U3647 | ~new_P1_U4243 | ~new_P1_U4242;
  assign new_P1_U3381 = ~new_P1_U3653 | ~new_P1_U3651 | ~new_P1_U4262 | ~new_P1_U4261;
  assign new_P1_U3382 = ~new_P1_U3657 | ~new_P1_U3655 | ~new_P1_U4281 | ~new_P1_U4280;
  assign new_P1_U3383 = ~new_P1_U3661 | ~new_P1_U3659 | ~new_P1_U4300 | ~new_P1_U4299;
  assign new_P1_U3384 = ~new_P1_U3665 | ~new_P1_U3663 | ~new_P1_U4319 | ~new_P1_U4318;
  assign new_P1_U3385 = ~new_P1_U3669 | ~new_P1_U3667 | ~new_P1_U4338 | ~new_P1_U4337;
  assign new_P1_U3386 = ~new_P1_U3673 | ~new_P1_U3671 | ~new_P1_U4357 | ~new_P1_U4356;
  assign new_P1_U3387 = ~new_P1_U3677 | ~new_P1_U3675 | ~new_P1_U4376 | ~new_P1_U4375;
  assign new_P1_U3388 = ~new_P1_U3681 | ~new_P1_U3679 | ~new_P1_U4395 | ~new_P1_U4394;
  assign new_P1_U3389 = ~new_P1_U3685 | ~new_P1_U3683 | ~new_P1_U4414 | ~new_P1_U4413;
  assign new_P1_U3390 = ~new_P1_U3689 | ~new_P1_U3687 | ~new_P1_U4433 | ~new_P1_U4432;
  assign new_P1_U3391 = ~new_P1_U3693 | ~new_P1_U3691 | ~new_P1_U4452 | ~new_P1_U4451;
  assign new_P1_U3392 = ~new_P1_U3697 | ~new_P1_U3695 | ~new_P1_U4471 | ~new_P1_U4470;
  assign new_P1_U3393 = ~new_P1_U3701 | ~new_P1_U3699 | ~new_P1_U4490 | ~new_P1_U4489;
  assign new_P1_U3394 = ~new_P1_U3705 | ~new_P1_U3703 | ~new_P1_U4509 | ~new_P1_U4508;
  assign new_P1_U3395 = ~new_U76 | ~new_P1_U3912;
  assign new_P1_U3396 = ~new_P1_U3709 | ~new_P1_U3707 | ~new_P1_U4528 | ~new_P1_U4527;
  assign new_P1_U3397 = ~new_U75 | ~new_P1_U3912;
  assign new_P1_U3398 = ~new_P1_U3713 | ~new_P1_U3711 | ~new_P1_U4547 | ~new_P1_U4546;
  assign new_P1_U3399 = ~new_U74 | ~new_P1_U3912;
  assign new_P1_U3400 = ~new_P1_U3717 | ~new_P1_U3715 | ~new_P1_U4566 | ~new_P1_U4565;
  assign new_P1_U3401 = ~new_U73 | ~new_P1_U3912;
  assign new_P1_U3402 = ~new_P1_U3721 | ~new_P1_U3719 | ~new_P1_U4585 | ~new_P1_U4584;
  assign new_P1_U3403 = ~new_U72 | ~new_P1_U3912;
  assign new_P1_U3404 = ~new_P1_U3725 | ~new_P1_U3723 | ~new_P1_U4604 | ~new_P1_U4603;
  assign new_P1_U3405 = ~new_U71 | ~new_P1_U3912;
  assign new_P1_U3406 = ~new_P1_U3729 | ~new_P1_U3727 | ~new_P1_U4623 | ~new_P1_U4622;
  assign new_P1_U3407 = ~new_U70 | ~new_P1_U3912;
  assign new_P1_U3408 = ~new_P1_U3733 | ~new_P1_U3731 | ~new_P1_U4642 | ~new_P1_U4641;
  assign new_P1_U3409 = ~new_U69 | ~new_P1_U3912;
  assign new_P1_U3410 = ~new_P1_U3737 | ~new_P1_U3735 | ~new_P1_U4661 | ~new_P1_U4660;
  assign new_P1_U3411 = ~new_U68 | ~new_P1_U3912;
  assign new_P1_U3412 = ~new_P1_U3741 | ~new_P1_U3739 | ~new_P1_U4680 | ~new_P1_U4679;
  assign new_P1_U3413 = ~new_U67 | ~new_P1_U3912;
  assign new_P1_U3414 = ~new_U65 | ~new_P1_U3912;
  assign new_P1_U3415 = ~new_U64 | ~new_P1_U3912;
  assign new_P1_U3416 = ~new_P1_U3953 | ~new_P1_U5693;
  assign new_P1_U3417 = ~new_P1_U3022 | ~new_P1_U4724;
  assign new_P1_U3418 = ~new_P1_U3988 | ~new_P1_U5690;
  assign new_P1_U3419 = ~new_P1_U3048 | ~new_P1_U3447;
  assign new_P1_U3420 = ~new_P1_U3023 | ~new_P1_U5687;
  assign new_P1_U3421 = ~new_P1_U3050 | ~new_P1_U3436;
  assign new_P1_U3422 = ~new_P1_U3966 | ~new_P1_U4725;
  assign new_P1_U3423 = ~new_P1_U3424 | ~new_P1_U4888;
  assign new_P1_U3424 = ~new_P1_U4102 | ~new_P1_U5677;
  assign new_P1_U3425 = ~new_P1_U3999 | ~P1_STATE_REG;
  assign new_P1_U3426 = ~new_P1_U3438 | ~new_P1_U5687;
  assign new_P1_U3427 = ~new_P1_U3014 | ~new_P1_U3015;
  assign new_P1_U3428 = ~new_P1_U3443 | ~new_P1_U3438;
  assign new_P1_U3429 = ~new_P1_U3022 | ~new_P1_U3422;
  assign new_P1_U3430 = ~new_P1_U3867 | ~new_P1_U3016;
  assign new_P1_U3431 = ~new_P1_U3014 | ~new_P1_U3022;
  assign new_P1_U3432 = ~new_P1_U3870 | ~new_P1_U5101;
  assign new_P1_U3433 = ~new_P1_U3442 | ~new_P1_U5693;
  assign new_P1_U3434 = ~new_P1_U5371 | ~new_P1_U5370;
  assign new_P1_U3435 = ~new_P1_U5665 | ~new_P1_U5664;
  assign new_P1_U3436 = ~new_P1_U5668 | ~new_P1_U5667;
  assign new_P1_U3437 = ~new_P1_U5671 | ~new_P1_U5670;
  assign new_P1_U3438 = ~new_P1_U5676 | ~new_P1_U5675;
  assign n280 = ~new_P1_U5679 | ~new_P1_U5678;
  assign n285 = ~new_P1_U5681 | ~new_P1_U5680;
  assign new_P1_U3441 = ~new_P1_U5689 | ~new_P1_U5688;
  assign new_P1_U3442 = ~new_P1_U5686 | ~new_P1_U5685;
  assign new_P1_U3443 = ~new_P1_U5683 | ~new_P1_U5682;
  assign new_P1_U3444 = ~new_P1_U5707 | ~new_P1_U5706;
  assign new_P1_U3445 = ~new_P1_U5710 | ~new_P1_U5709;
  assign new_P1_U3446 = ~new_P1_U5698 | ~new_P1_U5697;
  assign new_P1_U3447 = ~new_P1_U5692 | ~new_P1_U5691;
  assign new_P1_U3448 = ~new_P1_U5695 | ~new_P1_U5694;
  assign new_P1_U3449 = ~new_P1_U5701 | ~new_P1_U5700;
  assign new_P1_U3450 = ~new_P1_U5704 | ~new_P1_U5703;
  assign new_P1_U3451 = ~new_P1_U5718 | ~new_P1_U5717;
  assign new_P1_U3452 = ~new_P1_U5715 | ~new_P1_U5714;
  assign n440 = ~new_P1_U5721 | ~new_P1_U5720;
  assign new_P1_U3454 = ~new_P1_U5723 | ~new_P1_U5722;
  assign new_P1_U3455 = ~new_P1_U5725 | ~new_P1_U5724;
  assign n445 = ~new_P1_U5728 | ~new_P1_U5727;
  assign new_P1_U3457 = ~new_P1_U5730 | ~new_P1_U5729;
  assign new_P1_U3458 = ~new_P1_U5732 | ~new_P1_U5731;
  assign n450 = ~new_P1_U5735 | ~new_P1_U5734;
  assign new_P1_U3460 = ~new_P1_U5737 | ~new_P1_U5736;
  assign new_P1_U3461 = ~new_P1_U5739 | ~new_P1_U5738;
  assign n455 = ~new_P1_U5742 | ~new_P1_U5741;
  assign new_P1_U3463 = ~new_P1_U5744 | ~new_P1_U5743;
  assign new_P1_U3464 = ~new_P1_U5746 | ~new_P1_U5745;
  assign n460 = ~new_P1_U5749 | ~new_P1_U5748;
  assign new_P1_U3466 = ~new_P1_U5751 | ~new_P1_U5750;
  assign new_P1_U3467 = ~new_P1_U5753 | ~new_P1_U5752;
  assign n465 = ~new_P1_U5756 | ~new_P1_U5755;
  assign new_P1_U3469 = ~new_P1_U5758 | ~new_P1_U5757;
  assign new_P1_U3470 = ~new_P1_U5760 | ~new_P1_U5759;
  assign n470 = ~new_P1_U5763 | ~new_P1_U5762;
  assign new_P1_U3472 = ~new_P1_U5765 | ~new_P1_U5764;
  assign new_P1_U3473 = ~new_P1_U5767 | ~new_P1_U5766;
  assign n475 = ~new_P1_U5770 | ~new_P1_U5769;
  assign new_P1_U3475 = ~new_P1_U5772 | ~new_P1_U5771;
  assign new_P1_U3476 = ~new_P1_U5774 | ~new_P1_U5773;
  assign n480 = ~new_P1_U5777 | ~new_P1_U5776;
  assign new_P1_U3478 = ~new_P1_U5779 | ~new_P1_U5778;
  assign new_P1_U3479 = ~new_P1_U5781 | ~new_P1_U5780;
  assign n485 = ~new_P1_U5784 | ~new_P1_U5783;
  assign new_P1_U3481 = ~new_P1_U5786 | ~new_P1_U5785;
  assign new_P1_U3482 = ~new_P1_U5788 | ~new_P1_U5787;
  assign n490 = ~new_P1_U5791 | ~new_P1_U5790;
  assign new_P1_U3484 = ~new_P1_U5793 | ~new_P1_U5792;
  assign new_P1_U3485 = ~new_P1_U5795 | ~new_P1_U5794;
  assign n495 = ~new_P1_U5798 | ~new_P1_U5797;
  assign new_P1_U3487 = ~new_P1_U5800 | ~new_P1_U5799;
  assign new_P1_U3488 = ~new_P1_U5802 | ~new_P1_U5801;
  assign n500 = ~new_P1_U5805 | ~new_P1_U5804;
  assign new_P1_U3490 = ~new_P1_U5807 | ~new_P1_U5806;
  assign new_P1_U3491 = ~new_P1_U5809 | ~new_P1_U5808;
  assign n505 = ~new_P1_U5812 | ~new_P1_U5811;
  assign new_P1_U3493 = ~new_P1_U5814 | ~new_P1_U5813;
  assign new_P1_U3494 = ~new_P1_U5816 | ~new_P1_U5815;
  assign n510 = ~new_P1_U5819 | ~new_P1_U5818;
  assign new_P1_U3496 = ~new_P1_U5821 | ~new_P1_U5820;
  assign new_P1_U3497 = ~new_P1_U5823 | ~new_P1_U5822;
  assign n515 = ~new_P1_U5826 | ~new_P1_U5825;
  assign new_P1_U3499 = ~new_P1_U5828 | ~new_P1_U5827;
  assign new_P1_U3500 = ~new_P1_U5830 | ~new_P1_U5829;
  assign n520 = ~new_P1_U5833 | ~new_P1_U5832;
  assign new_P1_U3502 = ~new_P1_U5835 | ~new_P1_U5834;
  assign new_P1_U3503 = ~new_P1_U5837 | ~new_P1_U5836;
  assign n525 = ~new_P1_U5840 | ~new_P1_U5839;
  assign new_P1_U3505 = ~new_P1_U5842 | ~new_P1_U5841;
  assign new_P1_U3506 = ~new_P1_U5844 | ~new_P1_U5843;
  assign n530 = ~new_P1_U5847 | ~new_P1_U5846;
  assign new_P1_U3508 = ~new_P1_U5849 | ~new_P1_U5848;
  assign n535 = ~new_P1_U5852 | ~new_P1_U5851;
  assign n540 = ~new_P1_U5854 | ~new_P1_U5853;
  assign n545 = ~new_P1_U5856 | ~new_P1_U5855;
  assign n550 = ~new_P1_U5858 | ~new_P1_U5857;
  assign n555 = ~new_P1_U5860 | ~new_P1_U5859;
  assign n560 = ~new_P1_U5862 | ~new_P1_U5861;
  assign n565 = ~new_P1_U5864 | ~new_P1_U5863;
  assign n570 = ~new_P1_U5866 | ~new_P1_U5865;
  assign n575 = ~new_P1_U5868 | ~new_P1_U5867;
  assign n580 = ~new_P1_U5870 | ~new_P1_U5869;
  assign n585 = ~new_P1_U5872 | ~new_P1_U5871;
  assign n590 = ~new_P1_U5874 | ~new_P1_U5873;
  assign n595 = ~new_P1_U5876 | ~new_P1_U5875;
  assign n600 = ~new_P1_U5878 | ~new_P1_U5877;
  assign n605 = ~new_P1_U5880 | ~new_P1_U5879;
  assign n610 = ~new_P1_U5882 | ~new_P1_U5881;
  assign n615 = ~new_P1_U5884 | ~new_P1_U5883;
  assign n620 = ~new_P1_U5886 | ~new_P1_U5885;
  assign n625 = ~new_P1_U5888 | ~new_P1_U5887;
  assign n630 = ~new_P1_U5890 | ~new_P1_U5889;
  assign n635 = ~new_P1_U5892 | ~new_P1_U5891;
  assign n640 = ~new_P1_U5894 | ~new_P1_U5893;
  assign n645 = ~new_P1_U5896 | ~new_P1_U5895;
  assign n650 = ~new_P1_U5898 | ~new_P1_U5897;
  assign n655 = ~new_P1_U5900 | ~new_P1_U5899;
  assign n660 = ~new_P1_U5902 | ~new_P1_U5901;
  assign n665 = ~new_P1_U5904 | ~new_P1_U5903;
  assign n670 = ~new_P1_U5906 | ~new_P1_U5905;
  assign n675 = ~new_P1_U5908 | ~new_P1_U5907;
  assign n680 = ~new_P1_U5910 | ~new_P1_U5909;
  assign n685 = ~new_P1_U5912 | ~new_P1_U5911;
  assign n690 = ~new_P1_U5914 | ~new_P1_U5913;
  assign n695 = ~new_P1_U5916 | ~new_P1_U5915;
  assign n700 = ~new_P1_U5918 | ~new_P1_U5917;
  assign n705 = ~new_P1_U5920 | ~new_P1_U5919;
  assign n710 = ~new_P1_U5922 | ~new_P1_U5921;
  assign n715 = ~new_P1_U5924 | ~new_P1_U5923;
  assign n720 = ~new_P1_U5926 | ~new_P1_U5925;
  assign n725 = ~new_P1_U5928 | ~new_P1_U5927;
  assign n730 = ~new_P1_U5930 | ~new_P1_U5929;
  assign n735 = ~new_P1_U5932 | ~new_P1_U5931;
  assign n740 = ~new_P1_U5934 | ~new_P1_U5933;
  assign n745 = ~new_P1_U5936 | ~new_P1_U5935;
  assign n750 = ~new_P1_U5938 | ~new_P1_U5937;
  assign n755 = ~new_P1_U5940 | ~new_P1_U5939;
  assign n1020 = ~new_P1_U6006 | ~new_P1_U6005;
  assign n1025 = ~new_P1_U6008 | ~new_P1_U6007;
  assign n1030 = ~new_P1_U6010 | ~new_P1_U6009;
  assign n1035 = ~new_P1_U6012 | ~new_P1_U6011;
  assign n1040 = ~new_P1_U6014 | ~new_P1_U6013;
  assign n1045 = ~new_P1_U6016 | ~new_P1_U6015;
  assign n1050 = ~new_P1_U6018 | ~new_P1_U6017;
  assign n1055 = ~new_P1_U6020 | ~new_P1_U6019;
  assign n1060 = ~new_P1_U6022 | ~new_P1_U6021;
  assign n1065 = ~new_P1_U6024 | ~new_P1_U6023;
  assign n1070 = ~new_P1_U6026 | ~new_P1_U6025;
  assign n1075 = ~new_P1_U6028 | ~new_P1_U6027;
  assign n1080 = ~new_P1_U6030 | ~new_P1_U6029;
  assign n1085 = ~new_P1_U6032 | ~new_P1_U6031;
  assign n1090 = ~new_P1_U6034 | ~new_P1_U6033;
  assign n1095 = ~new_P1_U6036 | ~new_P1_U6035;
  assign n1100 = ~new_P1_U6038 | ~new_P1_U6037;
  assign n1105 = ~new_P1_U6040 | ~new_P1_U6039;
  assign n1110 = ~new_P1_U6042 | ~new_P1_U6041;
  assign n1115 = ~new_P1_U6044 | ~new_P1_U6043;
  assign n1120 = ~new_P1_U6046 | ~new_P1_U6045;
  assign n1125 = ~new_P1_U6048 | ~new_P1_U6047;
  assign n1130 = ~new_P1_U6050 | ~new_P1_U6049;
  assign n1135 = ~new_P1_U6052 | ~new_P1_U6051;
  assign n1140 = ~new_P1_U6054 | ~new_P1_U6053;
  assign n1145 = ~new_P1_U6056 | ~new_P1_U6055;
  assign n1150 = ~new_P1_U6058 | ~new_P1_U6057;
  assign n1155 = ~new_P1_U6060 | ~new_P1_U6059;
  assign n1160 = ~new_P1_U6062 | ~new_P1_U6061;
  assign n1165 = ~new_P1_U6064 | ~new_P1_U6063;
  assign n1170 = ~new_P1_U6066 | ~new_P1_U6065;
  assign n1175 = ~new_P1_U6068 | ~new_P1_U6067;
  assign new_P1_U3586 = ~new_P1_U6172 | ~new_P1_U6171;
  assign new_P1_U3587 = ~new_P1_U6174 | ~new_P1_U6173;
  assign new_P1_U3588 = ~new_P1_U6176 | ~new_P1_U6175;
  assign new_P1_U3589 = ~new_P1_U6178 | ~new_P1_U6177;
  assign new_P1_U3590 = ~new_P1_U6180 | ~new_P1_U6179;
  assign new_P1_U3591 = ~new_P1_U6182 | ~new_P1_U6181;
  assign new_P1_U3592 = ~new_P1_U6184 | ~new_P1_U6183;
  assign new_P1_U3593 = ~new_P1_U6186 | ~new_P1_U6185;
  assign new_P1_U3594 = ~new_P1_U6188 | ~new_P1_U6187;
  assign new_P1_U3595 = ~new_P1_U6190 | ~new_P1_U6189;
  assign new_P1_U3596 = ~new_P1_U6192 | ~new_P1_U6191;
  assign new_P1_U3597 = ~new_P1_U6194 | ~new_P1_U6193;
  assign new_P1_U3598 = ~new_P1_U6196 | ~new_P1_U6195;
  assign new_P1_U3599 = ~new_P1_U6198 | ~new_P1_U6197;
  assign new_P1_U3600 = ~new_P1_U6200 | ~new_P1_U6199;
  assign new_P1_U3601 = ~new_P1_U6202 | ~new_P1_U6201;
  assign new_P1_U3602 = ~new_P1_U6204 | ~new_P1_U6203;
  assign new_P1_U3603 = ~new_P1_U6206 | ~new_P1_U6205;
  assign new_P1_U3604 = ~new_P1_U6208 | ~new_P1_U6207;
  assign new_P1_U3605 = ~new_P1_U6210 | ~new_P1_U6209;
  assign new_P1_U3606 = ~new_P1_U6212 | ~new_P1_U6211;
  assign new_P1_U3607 = ~new_P1_U6214 | ~new_P1_U6213;
  assign new_P1_U3608 = ~new_P1_U6216 | ~new_P1_U6215;
  assign new_P1_U3609 = ~new_P1_U6218 | ~new_P1_U6217;
  assign new_P1_U3610 = ~new_P1_U6220 | ~new_P1_U6219;
  assign new_P1_U3611 = ~new_P1_U6222 | ~new_P1_U6221;
  assign new_P1_U3612 = ~new_P1_U6224 | ~new_P1_U6223;
  assign new_P1_U3613 = ~new_P1_U6226 | ~new_P1_U6225;
  assign new_P1_U3614 = ~new_P1_U6228 | ~new_P1_U6227;
  assign new_P1_U3615 = ~new_P1_U6230 | ~new_P1_U6229;
  assign new_P1_U3616 = ~new_P1_U6232 | ~new_P1_U6231;
  assign new_P1_U3617 = ~new_P1_U6234 | ~new_P1_U6233;
  assign new_P1_U3618 = new_P1_U4144 & new_P1_U4143;
  assign new_P1_U3619 = new_P1_U4146 & new_P1_U4145;
  assign new_P1_U3620 = new_P1_U4151 & new_P1_U4154 & new_P1_U4152 & new_P1_U4153;
  assign new_P1_U3621 = new_P1_U4105 & new_P1_U4106 & new_P1_U4108 & new_P1_U4107;
  assign new_P1_U3622 = new_P1_U4109 & new_P1_U4110 & new_P1_U4112 & new_P1_U4111;
  assign new_P1_U3623 = new_P1_U4113 & new_P1_U4114 & new_P1_U4116 & new_P1_U4115;
  assign new_P1_U3624 = new_P1_U4119 & new_P1_U4118 & new_P1_U4117;
  assign new_P1_U3625 = new_P1_U3621 & new_P1_U3622 & new_P1_U3624 & new_P1_U3623;
  assign new_P1_U3626 = new_P1_U4120 & new_P1_U4121 & new_P1_U4123 & new_P1_U4122;
  assign new_P1_U3627 = new_P1_U4124 & new_P1_U4125 & new_P1_U4127 & new_P1_U4126;
  assign new_P1_U3628 = new_P1_U4128 & new_P1_U4129 & new_P1_U4131 & new_P1_U4130;
  assign new_P1_U3629 = new_P1_U4134 & new_P1_U4133 & new_P1_U4132;
  assign new_P1_U3630 = new_P1_U3626 & new_P1_U3627 & new_P1_U3629 & new_P1_U3628;
  assign new_P1_U3631 = new_P1_U5716 & new_P1_U4136;
  assign new_P1_U3632 = new_P1_U5719 & new_P1_U3022;
  assign new_P1_U3633 = new_P1_U4169 & new_P1_U4168;
  assign new_P1_U3634 = new_P1_U4171 & new_P1_U4170;
  assign new_P1_U3635 = new_P1_U3634 & new_P1_U4173 & new_P1_U4172;
  assign new_P1_U3636 = new_P1_U4175 & new_P1_U4178 & new_P1_U4176 & new_P1_U4177;
  assign new_P1_U3637 = new_P1_U4188 & new_P1_U4187;
  assign new_P1_U3638 = new_P1_U4190 & new_P1_U4189;
  assign new_P1_U3639 = new_P1_U3638 & new_P1_U4192 & new_P1_U4191;
  assign new_P1_U3640 = new_P1_U4194 & new_P1_U4197 & new_P1_U4195 & new_P1_U4196;
  assign new_P1_U3641 = new_P1_U4209 & new_P1_U4208;
  assign new_P1_U3642 = new_P1_U3641 & new_P1_U4211 & new_P1_U4210;
  assign new_P1_U3643 = new_P1_U4213 & new_P1_U4216 & new_P1_U4214 & new_P1_U4215;
  assign new_P1_U3644 = new_P1_U4228 & new_P1_U4227;
  assign new_P1_U3645 = new_P1_U3644 & new_P1_U4230 & new_P1_U4229;
  assign new_P1_U3646 = new_P1_U4232 & new_P1_U4235 & new_P1_U4233 & new_P1_U4234;
  assign new_P1_U3647 = new_P1_U4245 & new_P1_U4244;
  assign new_P1_U3648 = new_P1_U4247 & new_P1_U4246;
  assign new_P1_U3649 = new_P1_U3648 & new_P1_U4249 & new_P1_U4248;
  assign new_P1_U3650 = new_P1_U4251 & new_P1_U4254 & new_P1_U4252 & new_P1_U4253;
  assign new_P1_U3651 = new_P1_U4264 & new_P1_U4263;
  assign new_P1_U3652 = new_P1_U4266 & new_P1_U4265;
  assign new_P1_U3653 = new_P1_U3652 & new_P1_U4268 & new_P1_U4267;
  assign new_P1_U3654 = new_P1_U4270 & new_P1_U4273 & new_P1_U4271 & new_P1_U4272;
  assign new_P1_U3655 = new_P1_U4283 & new_P1_U4282;
  assign new_P1_U3656 = new_P1_U4285 & new_P1_U4284;
  assign new_P1_U3657 = new_P1_U3656 & new_P1_U4287 & new_P1_U4286;
  assign new_P1_U3658 = new_P1_U4289 & new_P1_U4292 & new_P1_U4290 & new_P1_U4291;
  assign new_P1_U3659 = new_P1_U4302 & new_P1_U4301;
  assign new_P1_U3660 = new_P1_U4304 & new_P1_U4303;
  assign new_P1_U3661 = new_P1_U3660 & new_P1_U4306 & new_P1_U4305;
  assign new_P1_U3662 = new_P1_U4308 & new_P1_U4311 & new_P1_U4309 & new_P1_U4310;
  assign new_P1_U3663 = new_P1_U4321 & new_P1_U4320;
  assign new_P1_U3664 = new_P1_U4323 & new_P1_U4322;
  assign new_P1_U3665 = new_P1_U3664 & new_P1_U4325 & new_P1_U4324;
  assign new_P1_U3666 = new_P1_U4327 & new_P1_U4330 & new_P1_U4328 & new_P1_U4329;
  assign new_P1_U3667 = new_P1_U4340 & new_P1_U4339;
  assign new_P1_U3668 = new_P1_U4342 & new_P1_U4341;
  assign new_P1_U3669 = new_P1_U3668 & new_P1_U4344 & new_P1_U4343;
  assign new_P1_U3670 = new_P1_U4346 & new_P1_U4349 & new_P1_U4347 & new_P1_U4348;
  assign new_P1_U3671 = new_P1_U4359 & new_P1_U4358;
  assign new_P1_U3672 = new_P1_U4361 & new_P1_U4360;
  assign new_P1_U3673 = new_P1_U3672 & new_P1_U4363 & new_P1_U4362;
  assign new_P1_U3674 = new_P1_U4367 & new_P1_U4366 & new_P1_U4368 & new_P1_U4365;
  assign new_P1_U3675 = new_P1_U4378 & new_P1_U4377;
  assign new_P1_U3676 = new_P1_U4380 & new_P1_U4379;
  assign new_P1_U3677 = new_P1_U3676 & new_P1_U4382 & new_P1_U4381;
  assign new_P1_U3678 = new_P1_U4386 & new_P1_U4385 & new_P1_U4387 & new_P1_U4384;
  assign new_P1_U3679 = new_P1_U4397 & new_P1_U4396;
  assign new_P1_U3680 = new_P1_U4399 & new_P1_U4398;
  assign new_P1_U3681 = new_P1_U3680 & new_P1_U4401 & new_P1_U4400;
  assign new_P1_U3682 = new_P1_U4403 & new_P1_U4404 & new_P1_U4406 & new_P1_U4405;
  assign new_P1_U3683 = new_P1_U4416 & new_P1_U4415;
  assign new_P1_U3684 = new_P1_U4418 & new_P1_U4417;
  assign new_P1_U3685 = new_P1_U3684 & new_P1_U4420 & new_P1_U4419;
  assign new_P1_U3686 = new_P1_U4424 & new_P1_U4425 & new_P1_U4423 & new_P1_U4422;
  assign new_P1_U3687 = new_P1_U4435 & new_P1_U4434;
  assign new_P1_U3688 = new_P1_U4437 & new_P1_U4436;
  assign new_P1_U3689 = new_P1_U3688 & new_P1_U4439 & new_P1_U4438;
  assign new_P1_U3690 = new_P1_U4443 & new_P1_U4444 & new_P1_U4442 & new_P1_U4441;
  assign new_P1_U3691 = new_P1_U4454 & new_P1_U4453;
  assign new_P1_U3692 = new_P1_U4456 & new_P1_U4455;
  assign new_P1_U3693 = new_P1_U3692 & new_P1_U4458 & new_P1_U4457;
  assign new_P1_U3694 = new_P1_U4462 & new_P1_U4463 & new_P1_U4461 & new_P1_U4460;
  assign new_P1_U3695 = new_P1_U4473 & new_P1_U4472;
  assign new_P1_U3696 = new_P1_U4475 & new_P1_U4474;
  assign new_P1_U3697 = new_P1_U3696 & new_P1_U4477 & new_P1_U4476;
  assign new_P1_U3698 = new_P1_U4481 & new_P1_U4482 & new_P1_U4480 & new_P1_U4479;
  assign new_P1_U3699 = new_P1_U4492 & new_P1_U4491;
  assign new_P1_U3700 = new_P1_U4494 & new_P1_U4493;
  assign new_P1_U3701 = new_P1_U3700 & new_P1_U4496 & new_P1_U4495;
  assign new_P1_U3702 = new_P1_U4500 & new_P1_U4501 & new_P1_U4499 & new_P1_U4498;
  assign new_P1_U3703 = new_P1_U4511 & new_P1_U4510;
  assign new_P1_U3704 = new_P1_U4513 & new_P1_U4512;
  assign new_P1_U3705 = new_P1_U3704 & new_P1_U4515 & new_P1_U4514;
  assign new_P1_U3706 = new_P1_U4519 & new_P1_U4520 & new_P1_U4518 & new_P1_U4517;
  assign new_P1_U3707 = new_P1_U4530 & new_P1_U4529;
  assign new_P1_U3708 = new_P1_U4532 & new_P1_U4531;
  assign new_P1_U3709 = new_P1_U3708 & new_P1_U4534 & new_P1_U4533;
  assign new_P1_U3710 = new_P1_U4536 & new_P1_U4537 & new_P1_U4539 & new_P1_U4538;
  assign new_P1_U3711 = new_P1_U4549 & new_P1_U4548;
  assign new_P1_U3712 = new_P1_U4551 & new_P1_U4550;
  assign new_P1_U3713 = new_P1_U3712 & new_P1_U4553 & new_P1_U4552;
  assign new_P1_U3714 = new_P1_U4557 & new_P1_U4558 & new_P1_U4556 & new_P1_U4555;
  assign new_P1_U3715 = new_P1_U4568 & new_P1_U4567;
  assign new_P1_U3716 = new_P1_U4570 & new_P1_U4569;
  assign new_P1_U3717 = new_P1_U3716 & new_P1_U4572 & new_P1_U4571;
  assign new_P1_U3718 = new_P1_U4574 & new_P1_U4575 & new_P1_U4577 & new_P1_U4576;
  assign new_P1_U3719 = new_P1_U4587 & new_P1_U4586;
  assign new_P1_U3720 = new_P1_U4589 & new_P1_U4588;
  assign new_P1_U3721 = new_P1_U3720 & new_P1_U4591 & new_P1_U4590;
  assign new_P1_U3722 = new_P1_U4595 & new_P1_U4594 & new_P1_U4596 & new_P1_U4593;
  assign new_P1_U3723 = new_P1_U4606 & new_P1_U4605;
  assign new_P1_U3724 = new_P1_U4608 & new_P1_U4607;
  assign new_P1_U3725 = new_P1_U3724 & new_P1_U4610 & new_P1_U4609;
  assign new_P1_U3726 = new_P1_U4612 & new_P1_U4615 & new_P1_U4613 & new_P1_U4614;
  assign new_P1_U3727 = new_P1_U4625 & new_P1_U4624;
  assign new_P1_U3728 = new_P1_U4627 & new_P1_U4626;
  assign new_P1_U3729 = new_P1_U3728 & new_P1_U4629 & new_P1_U4628;
  assign new_P1_U3730 = new_P1_U4631 & new_P1_U4634 & new_P1_U4632 & new_P1_U4633;
  assign new_P1_U3731 = new_P1_U4644 & new_P1_U4643;
  assign new_P1_U3732 = new_P1_U4646 & new_P1_U4645;
  assign new_P1_U3733 = new_P1_U3732 & new_P1_U4648 & new_P1_U4647;
  assign new_P1_U3734 = new_P1_U4650 & new_P1_U4653 & new_P1_U4651 & new_P1_U4652;
  assign new_P1_U3735 = new_P1_U4663 & new_P1_U4662;
  assign new_P1_U3736 = new_P1_U4665 & new_P1_U4664;
  assign new_P1_U3737 = new_P1_U3736 & new_P1_U4667 & new_P1_U4666;
  assign new_P1_U3738 = new_P1_U4669 & new_P1_U4672 & new_P1_U4670 & new_P1_U4671;
  assign new_P1_U3739 = new_P1_U4682 & new_P1_U4681;
  assign new_P1_U3740 = new_P1_U4684 & new_P1_U4683;
  assign new_P1_U3741 = new_P1_U3740 & new_P1_U4686 & new_P1_U4685;
  assign new_P1_U3742 = new_P1_U4688 & new_P1_U4691 & new_P1_U4689 & new_P1_U4690;
  assign new_P1_U3743 = new_P1_U4698 & new_P1_U3987;
  assign new_P1_U3744 = new_P1_U4704 & new_P1_U4702 & new_P1_U4701;
  assign new_P1_U3745 = new_P1_U4707 & new_P1_U4705;
  assign new_P1_U3746 = new_P1_U4709 & new_P1_U4710 & new_P1_U4711;
  assign new_P1_U3747 = new_P1_U3987 & new_P1_U4698;
  assign new_P1_U3748 = new_P1_U3022 & new_P1_U3451;
  assign new_P1_U3749 = new_P1_U3452 & new_P1_U5719 & new_P1_U3969;
  assign new_P1_U3750 = new_P1_U4729 & new_P1_U4728 & new_P1_U4727;
  assign new_P1_U3751 = new_P1_U3915 & new_P1_U4731 & new_P1_U4730;
  assign new_P1_U3752 = new_P1_U4734 & new_P1_U4733 & new_P1_U4732;
  assign new_P1_U3753 = new_P1_U3916 & new_P1_U4736 & new_P1_U4735;
  assign new_P1_U3754 = new_P1_U4739 & new_P1_U4738 & new_P1_U4737;
  assign new_P1_U3755 = new_P1_U3917 & new_P1_U4741 & new_P1_U4740;
  assign new_P1_U3756 = new_P1_U4744 & new_P1_U4743 & new_P1_U4742;
  assign new_P1_U3757 = new_P1_U4746 & new_P1_U4745;
  assign new_P1_U3758 = new_P1_U4748 & new_P1_U4747;
  assign new_P1_U3759 = new_P1_U4751 & new_P1_U4750;
  assign new_P1_U3760 = new_P1_U4753 & new_P1_U4752;
  assign new_P1_U3761 = new_P1_U4756 & new_P1_U4755;
  assign new_P1_U3762 = new_P1_U4758 & new_P1_U4757;
  assign new_P1_U3763 = new_P1_U4761 & new_P1_U4760;
  assign new_P1_U3764 = new_P1_U4763 & new_P1_U4762;
  assign new_P1_U3765 = new_P1_U4766 & new_P1_U4765;
  assign new_P1_U3766 = new_P1_U4768 & new_P1_U4767;
  assign new_P1_U3767 = new_P1_U4771 & new_P1_U4770;
  assign new_P1_U3768 = new_P1_U4773 & new_P1_U4772;
  assign new_P1_U3769 = new_P1_U4776 & new_P1_U4775;
  assign new_P1_U3770 = new_P1_U4778 & new_P1_U4777;
  assign new_P1_U3771 = new_P1_U4781 & new_P1_U4780;
  assign new_P1_U3772 = new_P1_U4784 & new_P1_U4783 & new_P1_U4782;
  assign new_P1_U3773 = new_P1_U4786 & new_P1_U4785;
  assign new_P1_U3774 = new_P1_U4789 & new_P1_U4788 & new_P1_U4787;
  assign new_P1_U3775 = new_P1_U4791 & new_P1_U4790;
  assign new_P1_U3776 = new_P1_U4794 & new_P1_U4793 & new_P1_U4792;
  assign new_P1_U3777 = new_P1_U4796 & new_P1_U4795;
  assign new_P1_U3778 = new_P1_U4801 & new_P1_U4800 & new_P1_U4799 & new_P1_U4798 & new_P1_U4797;
  assign new_P1_U3779 = new_P1_U4806 & new_P1_U4805 & new_P1_U4804 & new_P1_U4803 & new_P1_U4802;
  assign new_P1_U3780 = new_P1_U4811 & new_P1_U4810 & new_P1_U4809 & new_P1_U4808 & new_P1_U4807;
  assign new_P1_U3781 = new_P1_U4816 & new_P1_U4815 & new_P1_U4814 & new_P1_U4813 & new_P1_U4812;
  assign new_P1_U3782 = new_P1_U4821 & new_P1_U4820 & new_P1_U4819 & new_P1_U4818 & new_P1_U4817;
  assign new_P1_U3783 = new_P1_U4826 & new_P1_U4825 & new_P1_U4824 & new_P1_U4823 & new_P1_U4822;
  assign new_P1_U3784 = new_P1_U4829 & new_P1_U4828 & new_P1_U4827;
  assign new_P1_U3785 = new_P1_U4831 & new_P1_U4830;
  assign new_P1_U3786 = new_P1_U4836 & new_P1_U4835 & new_P1_U4834 & new_P1_U4833 & new_P1_U4832;
  assign new_P1_U3787 = new_P1_U4839 & new_P1_U4838 & new_P1_U4837;
  assign new_P1_U3788 = new_P1_U4841 & new_P1_U4840;
  assign new_P1_U3789 = new_P1_U4844 & new_P1_U4843 & new_P1_U4842;
  assign new_P1_U3790 = new_P1_U4846 & new_P1_U4845;
  assign new_P1_U3791 = new_P1_U4848 & new_P1_U4847;
  assign new_P1_U3792 = new_P1_U4851 & new_P1_U4850;
  assign new_P1_U3793 = new_P1_U4853 & new_P1_U4852;
  assign new_P1_U3794 = new_P1_U4856 & new_P1_U4855;
  assign new_P1_U3795 = new_P1_U4858 & new_P1_U4857;
  assign new_P1_U3796 = new_P1_U4861 & new_P1_U4860;
  assign new_P1_U3797 = new_P1_U4863 & new_P1_U4862;
  assign new_P1_U3798 = new_P1_U4866 & new_P1_U4865;
  assign new_P1_U3799 = new_P1_U4868 & new_P1_U4867;
  assign new_P1_U3800 = new_P1_U4871 & new_P1_U4870;
  assign new_P1_U3801 = new_P1_U5658 & new_P1_U5657 & new_P1_U4707;
  assign new_P1_U3802 = new_P1_U5660 & new_P1_U5659;
  assign new_P1_U3803 = new_P1_U3366 & new_P1_U3419 & new_P1_U3370;
  assign new_P1_U3804 = new_P1_U3361 & new_P1_U3368 & new_P1_U3365;
  assign new_P1_U3805 = new_P1_U3362 & new_P1_U3364;
  assign new_P1_U3806 = new_P1_U3805 & new_P1_U3420;
  assign new_P1_U3807 = new_P1_U3438 & P1_STATE_REG;
  assign new_P1_U3808 = new_P1_U4891 & new_P1_U4892;
  assign new_P1_U3809 = new_P1_U4894 & new_P1_U4895 & new_P1_U4893;
  assign new_P1_U3810 = new_P1_U4901 & new_P1_U4902;
  assign new_P1_U3811 = new_P1_U4904 & new_P1_U4905 & new_P1_U4903;
  assign new_P1_U3812 = new_P1_U4911 & new_P1_U4912;
  assign new_P1_U3813 = new_P1_U4914 & new_P1_U4915 & new_P1_U4913;
  assign new_P1_U3814 = new_P1_U4921 & new_P1_U4922;
  assign new_P1_U3815 = new_P1_U4924 & new_P1_U4925 & new_P1_U4923;
  assign new_P1_U3816 = new_P1_U4931 & new_P1_U4932;
  assign new_P1_U3817 = new_P1_U4934 & new_P1_U4935 & new_P1_U4933;
  assign new_P1_U3818 = new_P1_U4941 & new_P1_U4942;
  assign new_P1_U3819 = new_P1_U4944 & new_P1_U4945 & new_P1_U4943;
  assign new_P1_U3820 = new_P1_U4951 & new_P1_U4952;
  assign new_P1_U3821 = new_P1_U4954 & new_P1_U4955 & new_P1_U4953;
  assign new_P1_U3822 = new_P1_U4961 & new_P1_U4962;
  assign new_P1_U3823 = new_P1_U4964 & new_P1_U4965 & new_P1_U4963;
  assign new_P1_U3824 = new_P1_U4971 & new_P1_U4972;
  assign new_P1_U3825 = new_P1_U4974 & new_P1_U4975 & new_P1_U4973;
  assign new_P1_U3826 = new_P1_U4981 & new_P1_U4982;
  assign new_P1_U3827 = new_P1_U4984 & new_P1_U4985 & new_P1_U4983;
  assign new_P1_U3828 = new_P1_U4991 & new_P1_U4992;
  assign new_P1_U3829 = new_P1_U4994 & new_P1_U4995 & new_P1_U4993;
  assign new_P1_U3830 = new_P1_U5001 & new_P1_U5002;
  assign new_P1_U3831 = new_P1_U5004 & new_P1_U5005 & new_P1_U5003;
  assign new_P1_U3832 = new_P1_U5011 & new_P1_U5012;
  assign new_P1_U3833 = new_P1_U5015 & new_P1_U5014 & new_P1_U5013;
  assign new_P1_U3834 = new_P1_U5020 & new_P1_U5021 & new_P1_U5022;
  assign new_P1_U3835 = new_P1_U5025 & new_P1_U5024 & new_P1_U5023;
  assign new_P1_U3836 = new_P1_U5030 & new_P1_U5031 & new_P1_U5032;
  assign new_P1_U3837 = new_P1_U5035 & new_P1_U5034 & new_P1_U5033;
  assign new_P1_U3838 = new_P1_U5040 & new_P1_U3998;
  assign new_P1_U3839 = new_P1_U3838 & new_P1_U5042 & new_P1_U5041;
  assign new_P1_U3840 = new_P1_U5045 & new_P1_U5044 & new_P1_U5043;
  assign new_P1_U3841 = new_P1_U5050 & new_P1_U5051 & new_P1_U5052;
  assign new_P1_U3842 = new_P1_U5055 & new_P1_U5054 & new_P1_U5053;
  assign new_P1_U3843 = new_P1_U5060 & new_P1_U3998;
  assign new_P1_U3844 = new_P1_U3843 & new_P1_U5062 & new_P1_U5061;
  assign new_P1_U3845 = new_P1_U5065 & new_P1_U5064 & new_P1_U5063;
  assign new_P1_U3846 = new_P1_U5070 & new_P1_U5071 & new_P1_U5072;
  assign new_P1_U3847 = new_P1_U5075 & new_P1_U5074 & new_P1_U5073;
  assign new_P1_U3848 = new_P1_U5080 & new_P1_U5081 & new_P1_U5082;
  assign new_P1_U3849 = new_P1_U5085 & new_P1_U5084 & new_P1_U5083;
  assign new_P1_U3850 = P1_STATE_REG & new_P1_U3428;
  assign new_P1_U3851 = new_P1_U3850 & new_P1_U3424;
  assign new_P1_U3852 = new_P1_U6117 & new_P1_U6114 & new_P1_U6111;
  assign new_P1_U3853 = new_P1_U6129 & new_P1_U3854 & new_P1_U3852;
  assign new_P1_U3854 = new_P1_U6120 & new_P1_U6126 & new_P1_U6123;
  assign new_P1_U3855 = new_P1_U6141 & new_P1_U6138 & new_P1_U6135;
  assign new_P1_U3856 = new_P1_U6150 & new_P1_U6147 & new_P1_U6144;
  assign new_P1_U3857 = new_P1_U6132 & new_P1_U3856 & new_P1_U3855;
  assign new_P1_U3858 = new_P1_U6075 & new_P1_U6078 & new_P1_U6081 & new_P1_U3863 & new_P1_U3862;
  assign new_P1_U3859 = new_P1_U6168 & new_P1_U6156 & new_P1_U6159 & new_P1_U6165 & new_P1_U6162;
  assign new_P1_U3860 = new_P1_U3859 & new_P1_U6153 & new_P1_U6108 & new_P1_U3857 & new_P1_U3853;
  assign new_P1_U3861 = new_P1_U6102 & new_P1_U3858;
  assign new_P1_U3862 = new_P1_U6084 & new_P1_U6087 & new_P1_U6093 & new_P1_U6090;
  assign new_P1_U3863 = new_P1_U6099 & new_P1_U6096;
  assign new_P1_U3864 = new_P1_U5087 & new_P1_U5090 & new_P1_U5091;
  assign new_P1_U3865 = new_P1_U3052 & new_P1_U5690;
  assign new_P1_U3866 = new_P1_U5651 & new_P1_U5652;
  assign new_P1_U3867 = new_P1_U3451 & new_P1_U3452;
  assign new_P1_U3868 = new_P1_U3420 & new_P1_U3371 & new_P1_U3369;
  assign new_P1_U3869 = new_P1_U5677 & new_P1_U3969;
  assign new_P1_U3870 = new_P1_U3424 & new_P1_U3869;
  assign new_P1_U3871 = new_P1_U3022 & new_P1_U5100;
  assign new_P1_U3872 = new_P1_U5147 & new_P1_U5146;
  assign new_P1_U3873 = new_P1_U3994 & new_P1_U3078;
  assign new_P1_U3874 = new_P1_U5188 & new_P1_U5187;
  assign new_P1_U3875 = new_P1_U5191 & new_P1_U5190;
  assign new_P1_U3876 = new_P1_U5281 & new_P1_U5280;
  assign new_P1_U3877 = new_P1_U3433 & new_P1_U5366;
  assign new_P1_U3878 = new_P1_U5431 & new_P1_U5432;
  assign new_P1_U3879 = new_P1_U5514 & new_P1_U3438;
  assign new_P1_U3880 = new_P1_U5516 & new_P1_U3438;
  assign new_P1_U3881 = new_P1_U5518 & new_P1_U3438;
  assign new_P1_U3882 = new_P1_U5520 & new_P1_U3438;
  assign new_P1_U3883 = new_P1_U5522 & new_P1_U3438;
  assign new_P1_U3884 = new_P1_U5524 & new_P1_U3438;
  assign new_P1_U3885 = new_P1_U5526 & new_P1_U3438;
  assign new_P1_U3886 = new_P1_U5528 & new_P1_U3438;
  assign new_P1_U3887 = new_P1_U5530 & new_P1_U3438;
  assign new_P1_U3888 = new_P1_U3438 & new_P1_U5533;
  assign new_P1_U3889 = new_P1_U3438 & new_P1_U5535;
  assign new_P1_U3890 = new_P1_U3438 & new_P1_U5537;
  assign new_P1_U3891 = new_P1_U3438 & new_P1_U5539;
  assign new_P1_U3892 = new_P1_U3438 & new_P1_U5541;
  assign new_P1_U3893 = new_P1_U3438 & new_P1_U5543;
  assign new_P1_U3894 = new_P1_U3438 & new_P1_U5555;
  assign new_P1_U3895 = new_P1_U5587 & new_P1_U5585;
  assign new_P1_U3896 = new_P1_U5590 & new_P1_U5588;
  assign new_P1_U3897 = new_P1_U5593 & new_P1_U5591;
  assign new_P1_U3898 = new_P1_U5596 & new_P1_U5594;
  assign new_P1_U3899 = new_P1_U5599 & new_P1_U5597;
  assign new_P1_U3900 = new_P1_U5602 & new_P1_U5600;
  assign new_P1_U3901 = new_P1_U5605 & new_P1_U5603;
  assign new_P1_U3902 = new_P1_U5608 & new_P1_U5606;
  assign new_P1_U3903 = new_P1_U5611 & new_P1_U5609;
  assign new_P1_U3904 = new_P1_U5617 & new_P1_U5615;
  assign new_P1_U3905 = new_P1_U5620 & new_P1_U5618;
  assign new_P1_U3906 = new_P1_U5623 & new_P1_U5621;
  assign new_P1_U3907 = new_P1_U5626 & new_P1_U5624;
  assign new_P1_U3908 = new_P1_U5629 & new_P1_U5627;
  assign new_P1_U3909 = new_P1_U5632 & new_P1_U5630;
  assign new_P1_U3910 = ~P1_IR_REG_31_;
  assign new_P1_U3911 = ~new_P1_U3022 | ~new_P1_U3360;
  assign new_P1_U3912 = ~new_P1_U5702 | ~new_P1_U5699;
  assign new_P1_U3913 = ~new_P1_U3632 | ~new_P1_U3047;
  assign new_P1_U3914 = ~new_P1_U3748 | ~new_P1_U3047;
  assign new_P1_U3915 = new_P1_U5942 & new_P1_U5941;
  assign new_P1_U3916 = new_P1_U5944 & new_P1_U5943;
  assign new_P1_U3917 = new_P1_U5946 & new_P1_U5945;
  assign new_P1_U3918 = new_P1_U5948 & new_P1_U5947;
  assign new_P1_U3919 = new_P1_U5950 & new_P1_U5949;
  assign new_P1_U3920 = new_P1_U5952 & new_P1_U5951;
  assign new_P1_U3921 = new_P1_U5954 & new_P1_U5953;
  assign new_P1_U3922 = new_P1_U5956 & new_P1_U5955;
  assign new_P1_U3923 = new_P1_U5958 & new_P1_U5957;
  assign new_P1_U3924 = new_P1_U5960 & new_P1_U5959;
  assign new_P1_U3925 = new_P1_U5962 & new_P1_U5961;
  assign new_P1_U3926 = new_P1_U5964 & new_P1_U5963;
  assign new_P1_U3927 = new_P1_U5966 & new_P1_U5965;
  assign new_P1_U3928 = new_P1_U5968 & new_P1_U5967;
  assign new_P1_U3929 = new_P1_U5970 & new_P1_U5969;
  assign new_P1_U3930 = new_P1_U5972 & new_P1_U5971;
  assign new_P1_U3931 = new_P1_U5974 & new_P1_U5973;
  assign new_P1_U3932 = new_P1_U5976 & new_P1_U5975;
  assign new_P1_U3933 = new_P1_U5978 & new_P1_U5977;
  assign new_P1_U3934 = new_P1_U5980 & new_P1_U5979;
  assign new_P1_U3935 = new_P1_U5982 & new_P1_U5981;
  assign new_P1_U3936 = new_P1_U5984 & new_P1_U5983;
  assign new_P1_U3937 = new_P1_U5986 & new_P1_U5985;
  assign new_P1_U3938 = new_P1_U5988 & new_P1_U5987;
  assign new_P1_U3939 = new_P1_U5990 & new_P1_U5989;
  assign new_P1_U3940 = new_P1_U5992 & new_P1_U5991;
  assign new_P1_U3941 = new_P1_U5994 & new_P1_U5993;
  assign new_P1_U3942 = new_P1_U5996 & new_P1_U5995;
  assign new_P1_U3943 = new_P1_U5998 & new_P1_U5997;
  assign new_P1_U3944 = new_P1_U6000 & new_P1_U5999;
  assign new_P1_U3945 = ~new_P1_U3747 | ~new_P1_U3056;
  assign new_P1_U3946 = new_P1_U6002 & new_P1_U6001;
  assign new_P1_U3947 = new_P1_U6004 & new_P1_U6003;
  assign new_P1_U3948 = ~new_P1_R1375_U14;
  assign new_P1_U3949 = ~new_P1_R1360_U14;
  assign new_P1_U3950 = new_P1_U6072 & new_P1_U6071;
  assign new_P1_U3951 = ~new_P1_U3861 | ~new_P1_U3860 | ~new_P1_U6105;
  assign new_P1_U3952 = ~new_P1_R1352_U6;
  assign new_P1_U3953 = ~new_P1_U3372;
  assign new_P1_U3954 = ~new_P1_U3426;
  assign new_P1_U3955 = ~new_P1_U3428;
  assign new_P1_U3956 = ~new_P1_U3370;
  assign new_P1_U3957 = ~new_P1_U3419;
  assign new_P1_U3958 = ~new_P1_U3366;
  assign new_P1_U3959 = ~new_P1_U3365;
  assign new_P1_U3960 = ~new_P1_U3368;
  assign new_P1_U3961 = ~new_P1_U3361;
  assign new_P1_U3962 = ~new_P1_U3364;
  assign new_P1_U3963 = ~new_P1_U3362;
  assign new_P1_U3964 = ~new_P1_U3420;
  assign new_P1_U3965 = ~new_P1_U3418;
  assign new_P1_U3966 = ~new_P1_U3049 | ~new_P1_U4001;
  assign new_P1_U3967 = ~new_P1_U3371;
  assign new_P1_U3968 = ~new_P1_U3369;
  assign new_P1_U3969 = ~new_P1_U3987 | ~new_P1_U3367;
  assign new_P1_U3970 = ~new_P1_U3049 | ~new_P1_U3421;
  assign new_P1_U3971 = ~new_P1_U3912;
  assign new_P1_U3972 = ~new_P1_U3430;
  assign n1340 = ~new_P1_U3425;
  assign new_P1_U3974 = ~new_P1_U3411;
  assign new_P1_U3975 = ~new_P1_U3409;
  assign new_P1_U3976 = ~new_P1_U3407;
  assign new_P1_U3977 = ~new_P1_U3405;
  assign new_P1_U3978 = ~new_P1_U3403;
  assign new_P1_U3979 = ~new_P1_U3401;
  assign new_P1_U3980 = ~new_P1_U3399;
  assign new_P1_U3981 = ~new_P1_U3397;
  assign new_P1_U3982 = ~new_P1_U3395;
  assign new_P1_U3983 = ~new_P1_U3415;
  assign new_P1_U3984 = ~new_P1_U3414;
  assign new_P1_U3985 = ~new_P1_U3413;
  assign new_P1_U3986 = ~new_P1_U3427;
  assign new_P1_U3987 = ~new_P1_U3373;
  assign new_P1_U3988 = ~new_P1_U3416;
  assign new_P1_U3989 = ~new_P1_U3417;
  assign new_P1_U3990 = ~new_P1_U3914;
  assign new_P1_U3991 = ~new_P1_U3913;
  assign new_P1_U3992 = ~new_P1_U3911;
  assign new_P1_U3993 = ~new_P1_U3945;
  assign new_P1_U3994 = ~new_P1_U3431;
  assign new_P1_U3995 = ~new_P1_U3432 | ~P1_STATE_REG;
  assign new_P1_U3996 = ~new_P1_U3965 | ~new_P1_U3022;
  assign new_P1_U3997 = ~new_P1_U3429;
  assign new_P1_U3998 = ~n1340 | ~new_P1_U3212;
  assign new_P1_U3999 = ~new_P1_U3424;
  assign new_P1_U4000 = ~new_P1_U3433;
  assign new_P1_U4001 = ~new_P1_U3363;
  assign new_P1_U4002 = ~new_P1_U3367;
  assign new_P1_U4003 = ~new_P1_U3358;
  assign new_P1_U4004 = ~new_P1_U3357;
  assign new_P1_U4005 = ~new_U88 | ~n1330;
  assign new_P1_U4006 = ~P1_IR_REG_0_ | ~new_P1_U3028;
  assign new_P1_U4007 = ~P1_IR_REG_0_ | ~new_P1_U4004;
  assign new_P1_U4008 = ~new_U77 | ~n1330;
  assign new_P1_U4009 = ~new_P1_SUB_84_U40 | ~new_P1_U3028;
  assign new_P1_U4010 = ~P1_IR_REG_1_ | ~new_P1_U4004;
  assign new_P1_U4011 = ~new_U66 | ~n1330;
  assign new_P1_U4012 = ~new_P1_SUB_84_U21 | ~new_P1_U3028;
  assign new_P1_U4013 = ~P1_IR_REG_2_ | ~new_P1_U4004;
  assign new_P1_U4014 = ~new_U63 | ~n1330;
  assign new_P1_U4015 = ~new_P1_SUB_84_U22 | ~new_P1_U3028;
  assign new_P1_U4016 = ~P1_IR_REG_3_ | ~new_P1_U4004;
  assign new_P1_U4017 = ~new_U62 | ~n1330;
  assign new_P1_U4018 = ~new_P1_SUB_84_U23 | ~new_P1_U3028;
  assign new_P1_U4019 = ~P1_IR_REG_4_ | ~new_P1_U4004;
  assign new_P1_U4020 = ~new_U61 | ~n1330;
  assign new_P1_U4021 = ~new_P1_SUB_84_U162 | ~new_P1_U3028;
  assign new_P1_U4022 = ~P1_IR_REG_5_ | ~new_P1_U4004;
  assign new_P1_U4023 = ~new_U60 | ~n1330;
  assign new_P1_U4024 = ~new_P1_SUB_84_U24 | ~new_P1_U3028;
  assign new_P1_U4025 = ~P1_IR_REG_6_ | ~new_P1_U4004;
  assign new_P1_U4026 = ~new_U59 | ~n1330;
  assign new_P1_U4027 = ~new_P1_SUB_84_U25 | ~new_P1_U3028;
  assign new_P1_U4028 = ~P1_IR_REG_7_ | ~new_P1_U4004;
  assign new_P1_U4029 = ~new_U58 | ~n1330;
  assign new_P1_U4030 = ~new_P1_SUB_84_U26 | ~new_P1_U3028;
  assign new_P1_U4031 = ~P1_IR_REG_8_ | ~new_P1_U4004;
  assign new_P1_U4032 = ~new_U57 | ~n1330;
  assign new_P1_U4033 = ~new_P1_SUB_84_U160 | ~new_P1_U3028;
  assign new_P1_U4034 = ~P1_IR_REG_9_ | ~new_P1_U4004;
  assign new_P1_U4035 = ~new_U87 | ~n1330;
  assign new_P1_U4036 = ~new_P1_SUB_84_U6 | ~new_P1_U3028;
  assign new_P1_U4037 = ~P1_IR_REG_10_ | ~new_P1_U4004;
  assign new_P1_U4038 = ~new_U86 | ~n1330;
  assign new_P1_U4039 = ~new_P1_SUB_84_U7 | ~new_P1_U3028;
  assign new_P1_U4040 = ~P1_IR_REG_11_ | ~new_P1_U4004;
  assign new_P1_U4041 = ~new_U85 | ~n1330;
  assign new_P1_U4042 = ~new_P1_SUB_84_U8 | ~new_P1_U3028;
  assign new_P1_U4043 = ~P1_IR_REG_12_ | ~new_P1_U4004;
  assign new_P1_U4044 = ~new_U84 | ~n1330;
  assign new_P1_U4045 = ~new_P1_SUB_84_U179 | ~new_P1_U3028;
  assign new_P1_U4046 = ~P1_IR_REG_13_ | ~new_P1_U4004;
  assign new_P1_U4047 = ~new_U83 | ~n1330;
  assign new_P1_U4048 = ~new_P1_SUB_84_U9 | ~new_P1_U3028;
  assign new_P1_U4049 = ~P1_IR_REG_14_ | ~new_P1_U4004;
  assign new_P1_U4050 = ~new_U82 | ~n1330;
  assign new_P1_U4051 = ~new_P1_SUB_84_U10 | ~new_P1_U3028;
  assign new_P1_U4052 = ~P1_IR_REG_15_ | ~new_P1_U4004;
  assign new_P1_U4053 = ~new_U81 | ~n1330;
  assign new_P1_U4054 = ~new_P1_SUB_84_U11 | ~new_P1_U3028;
  assign new_P1_U4055 = ~P1_IR_REG_16_ | ~new_P1_U4004;
  assign new_P1_U4056 = ~new_U80 | ~n1330;
  assign new_P1_U4057 = ~new_P1_SUB_84_U177 | ~new_P1_U3028;
  assign new_P1_U4058 = ~P1_IR_REG_17_ | ~new_P1_U4004;
  assign new_P1_U4059 = ~new_U79 | ~n1330;
  assign new_P1_U4060 = ~new_P1_SUB_84_U12 | ~new_P1_U3028;
  assign new_P1_U4061 = ~P1_IR_REG_18_ | ~new_P1_U4004;
  assign new_P1_U4062 = ~new_U78 | ~n1330;
  assign new_P1_U4063 = ~new_P1_SUB_84_U13 | ~new_P1_U3028;
  assign new_P1_U4064 = ~P1_IR_REG_19_ | ~new_P1_U4004;
  assign new_P1_U4065 = ~new_U76 | ~n1330;
  assign new_P1_U4066 = ~new_P1_SUB_84_U14 | ~new_P1_U3028;
  assign new_P1_U4067 = ~P1_IR_REG_20_ | ~new_P1_U4004;
  assign new_P1_U4068 = ~new_U75 | ~n1330;
  assign new_P1_U4069 = ~new_P1_SUB_84_U173 | ~new_P1_U3028;
  assign new_P1_U4070 = ~P1_IR_REG_21_ | ~new_P1_U4004;
  assign new_P1_U4071 = ~new_U74 | ~n1330;
  assign new_P1_U4072 = ~new_P1_SUB_84_U15 | ~new_P1_U3028;
  assign new_P1_U4073 = ~P1_IR_REG_22_ | ~new_P1_U4004;
  assign new_P1_U4074 = ~new_U73 | ~n1330;
  assign new_P1_U4075 = ~new_P1_SUB_84_U16 | ~new_P1_U3028;
  assign new_P1_U4076 = ~P1_IR_REG_23_ | ~new_P1_U4004;
  assign new_P1_U4077 = ~new_U72 | ~n1330;
  assign new_P1_U4078 = ~new_P1_SUB_84_U17 | ~new_P1_U3028;
  assign new_P1_U4079 = ~P1_IR_REG_24_ | ~new_P1_U4004;
  assign new_P1_U4080 = ~new_U71 | ~n1330;
  assign new_P1_U4081 = ~new_P1_SUB_84_U170 | ~new_P1_U3028;
  assign new_P1_U4082 = ~P1_IR_REG_25_ | ~new_P1_U4004;
  assign new_P1_U4083 = ~new_U70 | ~n1330;
  assign new_P1_U4084 = ~new_P1_SUB_84_U18 | ~new_P1_U3028;
  assign new_P1_U4085 = ~P1_IR_REG_26_ | ~new_P1_U4004;
  assign new_P1_U4086 = ~new_U69 | ~n1330;
  assign new_P1_U4087 = ~new_P1_SUB_84_U42 | ~new_P1_U3028;
  assign new_P1_U4088 = ~P1_IR_REG_27_ | ~new_P1_U4004;
  assign new_P1_U4089 = ~new_U68 | ~n1330;
  assign new_P1_U4090 = ~new_P1_SUB_84_U19 | ~new_P1_U3028;
  assign new_P1_U4091 = ~P1_IR_REG_28_ | ~new_P1_U4004;
  assign new_P1_U4092 = ~new_U67 | ~n1330;
  assign new_P1_U4093 = ~new_P1_SUB_84_U20 | ~new_P1_U3028;
  assign new_P1_U4094 = ~P1_IR_REG_29_ | ~new_P1_U4004;
  assign new_P1_U4095 = ~new_U65 | ~n1330;
  assign new_P1_U4096 = ~new_P1_SUB_84_U165 | ~new_P1_U3028;
  assign new_P1_U4097 = ~P1_IR_REG_30_ | ~new_P1_U4004;
  assign new_P1_U4098 = ~new_U64 | ~n1330;
  assign new_P1_U4099 = ~new_P1_SUB_84_U41 | ~new_P1_U3028;
  assign new_P1_U4100 = ~P1_IR_REG_31_ | ~new_P1_U4004;
  assign new_P1_U4101 = ~new_P1_U3360;
  assign new_P1_U4102 = ~new_P1_U3421;
  assign new_P1_U4103 = ~new_P1_U3358 | ~new_P1_U5666;
  assign new_P1_U4104 = ~new_P1_U3358 | ~new_P1_U5669;
  assign new_P1_U4105 = ~new_P1_U4101 | ~P1_D_REG_10_;
  assign new_P1_U4106 = ~new_P1_U4101 | ~P1_D_REG_11_;
  assign new_P1_U4107 = ~new_P1_U4101 | ~P1_D_REG_12_;
  assign new_P1_U4108 = ~new_P1_U4101 | ~P1_D_REG_13_;
  assign new_P1_U4109 = ~new_P1_U4101 | ~P1_D_REG_14_;
  assign new_P1_U4110 = ~new_P1_U4101 | ~P1_D_REG_15_;
  assign new_P1_U4111 = ~new_P1_U4101 | ~P1_D_REG_16_;
  assign new_P1_U4112 = ~new_P1_U4101 | ~P1_D_REG_17_;
  assign new_P1_U4113 = ~new_P1_U4101 | ~P1_D_REG_18_;
  assign new_P1_U4114 = ~new_P1_U4101 | ~P1_D_REG_19_;
  assign new_P1_U4115 = ~new_P1_U4101 | ~P1_D_REG_20_;
  assign new_P1_U4116 = ~new_P1_U4101 | ~P1_D_REG_21_;
  assign new_P1_U4117 = ~new_P1_U4101 | ~P1_D_REG_22_;
  assign new_P1_U4118 = ~new_P1_U4101 | ~P1_D_REG_23_;
  assign new_P1_U4119 = ~new_P1_U4101 | ~P1_D_REG_24_;
  assign new_P1_U4120 = ~new_P1_U4101 | ~P1_D_REG_25_;
  assign new_P1_U4121 = ~new_P1_U4101 | ~P1_D_REG_26_;
  assign new_P1_U4122 = ~new_P1_U4101 | ~P1_D_REG_27_;
  assign new_P1_U4123 = ~new_P1_U4101 | ~P1_D_REG_28_;
  assign new_P1_U4124 = ~new_P1_U4101 | ~P1_D_REG_29_;
  assign new_P1_U4125 = ~new_P1_U4101 | ~P1_D_REG_2_;
  assign new_P1_U4126 = ~new_P1_U4101 | ~P1_D_REG_30_;
  assign new_P1_U4127 = ~new_P1_U4101 | ~P1_D_REG_31_;
  assign new_P1_U4128 = ~new_P1_U4101 | ~P1_D_REG_3_;
  assign new_P1_U4129 = ~new_P1_U4101 | ~P1_D_REG_4_;
  assign new_P1_U4130 = ~new_P1_U4101 | ~P1_D_REG_5_;
  assign new_P1_U4131 = ~new_P1_U4101 | ~P1_D_REG_6_;
  assign new_P1_U4132 = ~new_P1_U4101 | ~P1_D_REG_7_;
  assign new_P1_U4133 = ~new_P1_U4101 | ~P1_D_REG_8_;
  assign new_P1_U4134 = ~new_P1_U4101 | ~P1_D_REG_9_;
  assign new_P1_U4135 = ~new_P1_U5690 | ~new_P1_U5693;
  assign new_P1_U4136 = ~new_P1_U3367 | ~new_P1_U5713 | ~new_P1_U5712;
  assign new_P1_U4137 = ~new_P1_U3018 | ~P1_REG2_REG_1_;
  assign new_P1_U4138 = ~new_P1_U3019 | ~P1_REG1_REG_1_;
  assign new_P1_U4139 = ~new_P1_U3020 | ~P1_REG0_REG_1_;
  assign new_P1_U4140 = ~P1_REG3_REG_1_ | ~new_P1_U3017;
  assign new_P1_U4141 = ~new_P1_U3078;
  assign new_P1_U4142 = ~new_P1_U3966 | ~new_P1_U3416;
  assign new_P1_U4143 = ~new_P1_U3961 | ~new_P1_R1150_U18;
  assign new_P1_U4144 = ~new_P1_U3963 | ~new_P1_R1117_U18;
  assign new_P1_U4145 = ~new_P1_U3962 | ~new_P1_R1138_U96;
  assign new_P1_U4146 = ~new_P1_U3959 | ~new_P1_R1192_U18;
  assign new_P1_U4147 = ~new_P1_U3958 | ~new_P1_R1207_U18;
  assign new_P1_U4148 = ~new_P1_U3968 | ~new_P1_R1171_U96;
  assign new_P1_U4149 = ~new_P1_U3967 | ~new_P1_R1240_U96;
  assign new_P1_U4150 = ~new_P1_U3374;
  assign new_P1_U4151 = ~new_P1_R1222_U96 | ~new_P1_U3026;
  assign new_P1_U4152 = ~new_P1_U3025 | ~new_P1_U3078;
  assign new_P1_U4153 = ~new_P1_U3450 | ~new_P1_U3023;
  assign new_P1_U4154 = ~new_P1_U3450 | ~new_P1_U4142;
  assign new_P1_U4155 = ~new_P1_U3620 | ~new_P1_U4150;
  assign new_P1_U4156 = ~P1_REG2_REG_2_ | ~new_P1_U3018;
  assign new_P1_U4157 = ~P1_REG1_REG_2_ | ~new_P1_U3019;
  assign new_P1_U4158 = ~P1_REG0_REG_2_ | ~new_P1_U3020;
  assign new_P1_U4159 = ~P1_REG3_REG_2_ | ~new_P1_U3017;
  assign new_P1_U4160 = ~new_P1_U3068;
  assign new_P1_U4161 = ~P1_REG0_REG_0_ | ~new_P1_U3020;
  assign new_P1_U4162 = ~P1_REG1_REG_0_ | ~new_P1_U3019;
  assign new_P1_U4163 = ~P1_REG2_REG_0_ | ~new_P1_U3018;
  assign new_P1_U4164 = ~P1_REG3_REG_0_ | ~new_P1_U3017;
  assign new_P1_U4165 = ~new_P1_U3077;
  assign new_P1_U4166 = ~new_P1_U3033 | ~new_P1_U3077;
  assign new_P1_U4167 = ~new_P1_R1150_U96 | ~new_P1_U3961;
  assign new_P1_U4168 = ~new_P1_R1117_U96 | ~new_P1_U3963;
  assign new_P1_U4169 = ~new_P1_R1138_U95 | ~new_P1_U3962;
  assign new_P1_U4170 = ~new_P1_R1192_U96 | ~new_P1_U3959;
  assign new_P1_U4171 = ~new_P1_R1207_U96 | ~new_P1_U3958;
  assign new_P1_U4172 = ~new_P1_R1171_U95 | ~new_P1_U3968;
  assign new_P1_U4173 = ~new_P1_R1240_U95 | ~new_P1_U3967;
  assign new_P1_U4174 = ~new_P1_U3376;
  assign new_P1_U4175 = ~new_P1_R1222_U95 | ~new_P1_U3026;
  assign new_P1_U4176 = ~new_P1_U3025 | ~new_P1_U3068;
  assign new_P1_U4177 = ~new_P1_R1282_U57 | ~new_P1_U3023;
  assign new_P1_U4178 = ~new_P1_U3455 | ~new_P1_U4142;
  assign new_P1_U4179 = ~new_P1_U3636 | ~new_P1_U4174;
  assign new_P1_U4180 = ~P1_REG2_REG_3_ | ~new_P1_U3018;
  assign new_P1_U4181 = ~P1_REG1_REG_3_ | ~new_P1_U3019;
  assign new_P1_U4182 = ~P1_REG0_REG_3_ | ~new_P1_U3020;
  assign new_P1_U4183 = ~new_P1_ADD_95_U4 | ~new_P1_U3017;
  assign new_P1_U4184 = ~new_P1_U3064;
  assign new_P1_U4185 = ~new_P1_U3033 | ~new_P1_U3078;
  assign new_P1_U4186 = ~new_P1_R1150_U106 | ~new_P1_U3961;
  assign new_P1_U4187 = ~new_P1_R1117_U106 | ~new_P1_U3963;
  assign new_P1_U4188 = ~new_P1_R1138_U17 | ~new_P1_U3962;
  assign new_P1_U4189 = ~new_P1_R1192_U106 | ~new_P1_U3959;
  assign new_P1_U4190 = ~new_P1_R1207_U106 | ~new_P1_U3958;
  assign new_P1_U4191 = ~new_P1_R1171_U17 | ~new_P1_U3968;
  assign new_P1_U4192 = ~new_P1_R1240_U17 | ~new_P1_U3967;
  assign new_P1_U4193 = ~new_P1_U3377;
  assign new_P1_U4194 = ~new_P1_R1222_U17 | ~new_P1_U3026;
  assign new_P1_U4195 = ~new_P1_U3025 | ~new_P1_U3064;
  assign new_P1_U4196 = ~new_P1_R1282_U18 | ~new_P1_U3023;
  assign new_P1_U4197 = ~new_P1_U3458 | ~new_P1_U4142;
  assign new_P1_U4198 = ~new_P1_U3640 | ~new_P1_U4193;
  assign new_P1_U4199 = ~P1_REG2_REG_4_ | ~new_P1_U3018;
  assign new_P1_U4200 = ~P1_REG1_REG_4_ | ~new_P1_U3019;
  assign new_P1_U4201 = ~P1_REG0_REG_4_ | ~new_P1_U3020;
  assign new_P1_U4202 = ~new_P1_ADD_95_U59 | ~new_P1_U3017;
  assign new_P1_U4203 = ~new_P1_U3060;
  assign new_P1_U4204 = ~new_P1_U3033 | ~new_P1_U3068;
  assign new_P1_U4205 = ~new_P1_R1150_U15 | ~new_P1_U3961;
  assign new_P1_U4206 = ~new_P1_R1117_U15 | ~new_P1_U3963;
  assign new_P1_U4207 = ~new_P1_R1138_U101 | ~new_P1_U3962;
  assign new_P1_U4208 = ~new_P1_R1192_U15 | ~new_P1_U3959;
  assign new_P1_U4209 = ~new_P1_R1207_U15 | ~new_P1_U3958;
  assign new_P1_U4210 = ~new_P1_R1171_U101 | ~new_P1_U3968;
  assign new_P1_U4211 = ~new_P1_R1240_U101 | ~new_P1_U3967;
  assign new_P1_U4212 = ~new_P1_U3378;
  assign new_P1_U4213 = ~new_P1_R1222_U101 | ~new_P1_U3026;
  assign new_P1_U4214 = ~new_P1_U3025 | ~new_P1_U3060;
  assign new_P1_U4215 = ~new_P1_R1282_U20 | ~new_P1_U3023;
  assign new_P1_U4216 = ~new_P1_U3461 | ~new_P1_U4142;
  assign new_P1_U4217 = ~new_P1_U3643 | ~new_P1_U4212;
  assign new_P1_U4218 = ~P1_REG2_REG_5_ | ~new_P1_U3018;
  assign new_P1_U4219 = ~P1_REG1_REG_5_ | ~new_P1_U3019;
  assign new_P1_U4220 = ~P1_REG0_REG_5_ | ~new_P1_U3020;
  assign new_P1_U4221 = ~new_P1_ADD_95_U58 | ~new_P1_U3017;
  assign new_P1_U4222 = ~new_P1_U3067;
  assign new_P1_U4223 = ~new_P1_U3033 | ~new_P1_U3064;
  assign new_P1_U4224 = ~new_P1_R1150_U105 | ~new_P1_U3961;
  assign new_P1_U4225 = ~new_P1_R1117_U105 | ~new_P1_U3963;
  assign new_P1_U4226 = ~new_P1_R1138_U100 | ~new_P1_U3962;
  assign new_P1_U4227 = ~new_P1_R1192_U105 | ~new_P1_U3959;
  assign new_P1_U4228 = ~new_P1_R1207_U105 | ~new_P1_U3958;
  assign new_P1_U4229 = ~new_P1_R1171_U100 | ~new_P1_U3968;
  assign new_P1_U4230 = ~new_P1_R1240_U100 | ~new_P1_U3967;
  assign new_P1_U4231 = ~new_P1_U3379;
  assign new_P1_U4232 = ~new_P1_R1222_U100 | ~new_P1_U3026;
  assign new_P1_U4233 = ~new_P1_U3025 | ~new_P1_U3067;
  assign new_P1_U4234 = ~new_P1_R1282_U21 | ~new_P1_U3023;
  assign new_P1_U4235 = ~new_P1_U3464 | ~new_P1_U4142;
  assign new_P1_U4236 = ~new_P1_U3646 | ~new_P1_U4231;
  assign new_P1_U4237 = ~P1_REG2_REG_6_ | ~new_P1_U3018;
  assign new_P1_U4238 = ~P1_REG1_REG_6_ | ~new_P1_U3019;
  assign new_P1_U4239 = ~P1_REG0_REG_6_ | ~new_P1_U3020;
  assign new_P1_U4240 = ~new_P1_ADD_95_U57 | ~new_P1_U3017;
  assign new_P1_U4241 = ~new_P1_U3071;
  assign new_P1_U4242 = ~new_P1_U3033 | ~new_P1_U3060;
  assign new_P1_U4243 = ~new_P1_R1150_U104 | ~new_P1_U3961;
  assign new_P1_U4244 = ~new_P1_R1117_U104 | ~new_P1_U3963;
  assign new_P1_U4245 = ~new_P1_R1138_U18 | ~new_P1_U3962;
  assign new_P1_U4246 = ~new_P1_R1192_U104 | ~new_P1_U3959;
  assign new_P1_U4247 = ~new_P1_R1207_U104 | ~new_P1_U3958;
  assign new_P1_U4248 = ~new_P1_R1171_U18 | ~new_P1_U3968;
  assign new_P1_U4249 = ~new_P1_R1240_U18 | ~new_P1_U3967;
  assign new_P1_U4250 = ~new_P1_U3380;
  assign new_P1_U4251 = ~new_P1_R1222_U18 | ~new_P1_U3026;
  assign new_P1_U4252 = ~new_P1_U3025 | ~new_P1_U3071;
  assign new_P1_U4253 = ~new_P1_R1282_U65 | ~new_P1_U3023;
  assign new_P1_U4254 = ~new_P1_U3467 | ~new_P1_U4142;
  assign new_P1_U4255 = ~new_P1_U3650 | ~new_P1_U4250;
  assign new_P1_U4256 = ~P1_REG2_REG_7_ | ~new_P1_U3018;
  assign new_P1_U4257 = ~P1_REG1_REG_7_ | ~new_P1_U3019;
  assign new_P1_U4258 = ~P1_REG0_REG_7_ | ~new_P1_U3020;
  assign new_P1_U4259 = ~new_P1_ADD_95_U56 | ~new_P1_U3017;
  assign new_P1_U4260 = ~new_P1_U3070;
  assign new_P1_U4261 = ~new_P1_U3033 | ~new_P1_U3067;
  assign new_P1_U4262 = ~new_P1_R1150_U16 | ~new_P1_U3961;
  assign new_P1_U4263 = ~new_P1_R1117_U16 | ~new_P1_U3963;
  assign new_P1_U4264 = ~new_P1_R1138_U99 | ~new_P1_U3962;
  assign new_P1_U4265 = ~new_P1_R1192_U16 | ~new_P1_U3959;
  assign new_P1_U4266 = ~new_P1_R1207_U16 | ~new_P1_U3958;
  assign new_P1_U4267 = ~new_P1_R1171_U99 | ~new_P1_U3968;
  assign new_P1_U4268 = ~new_P1_R1240_U99 | ~new_P1_U3967;
  assign new_P1_U4269 = ~new_P1_U3381;
  assign new_P1_U4270 = ~new_P1_R1222_U99 | ~new_P1_U3026;
  assign new_P1_U4271 = ~new_P1_U3025 | ~new_P1_U3070;
  assign new_P1_U4272 = ~new_P1_R1282_U22 | ~new_P1_U3023;
  assign new_P1_U4273 = ~new_P1_U3470 | ~new_P1_U4142;
  assign new_P1_U4274 = ~new_P1_U3654 | ~new_P1_U4269;
  assign new_P1_U4275 = ~P1_REG2_REG_8_ | ~new_P1_U3018;
  assign new_P1_U4276 = ~P1_REG1_REG_8_ | ~new_P1_U3019;
  assign new_P1_U4277 = ~P1_REG0_REG_8_ | ~new_P1_U3020;
  assign new_P1_U4278 = ~new_P1_ADD_95_U55 | ~new_P1_U3017;
  assign new_P1_U4279 = ~new_P1_U3084;
  assign new_P1_U4280 = ~new_P1_U3033 | ~new_P1_U3071;
  assign new_P1_U4281 = ~new_P1_R1150_U103 | ~new_P1_U3961;
  assign new_P1_U4282 = ~new_P1_R1117_U103 | ~new_P1_U3963;
  assign new_P1_U4283 = ~new_P1_R1138_U19 | ~new_P1_U3962;
  assign new_P1_U4284 = ~new_P1_R1192_U103 | ~new_P1_U3959;
  assign new_P1_U4285 = ~new_P1_R1207_U103 | ~new_P1_U3958;
  assign new_P1_U4286 = ~new_P1_R1171_U19 | ~new_P1_U3968;
  assign new_P1_U4287 = ~new_P1_R1240_U19 | ~new_P1_U3967;
  assign new_P1_U4288 = ~new_P1_U3382;
  assign new_P1_U4289 = ~new_P1_R1222_U19 | ~new_P1_U3026;
  assign new_P1_U4290 = ~new_P1_U3025 | ~new_P1_U3084;
  assign new_P1_U4291 = ~new_P1_R1282_U23 | ~new_P1_U3023;
  assign new_P1_U4292 = ~new_P1_U3473 | ~new_P1_U4142;
  assign new_P1_U4293 = ~new_P1_U3658 | ~new_P1_U4288;
  assign new_P1_U4294 = ~P1_REG2_REG_9_ | ~new_P1_U3018;
  assign new_P1_U4295 = ~P1_REG1_REG_9_ | ~new_P1_U3019;
  assign new_P1_U4296 = ~P1_REG0_REG_9_ | ~new_P1_U3020;
  assign new_P1_U4297 = ~new_P1_ADD_95_U54 | ~new_P1_U3017;
  assign new_P1_U4298 = ~new_P1_U3083;
  assign new_P1_U4299 = ~new_P1_U3033 | ~new_P1_U3070;
  assign new_P1_U4300 = ~new_P1_R1150_U17 | ~new_P1_U3961;
  assign new_P1_U4301 = ~new_P1_R1117_U17 | ~new_P1_U3963;
  assign new_P1_U4302 = ~new_P1_R1138_U98 | ~new_P1_U3962;
  assign new_P1_U4303 = ~new_P1_R1192_U17 | ~new_P1_U3959;
  assign new_P1_U4304 = ~new_P1_R1207_U17 | ~new_P1_U3958;
  assign new_P1_U4305 = ~new_P1_R1171_U98 | ~new_P1_U3968;
  assign new_P1_U4306 = ~new_P1_R1240_U98 | ~new_P1_U3967;
  assign new_P1_U4307 = ~new_P1_U3383;
  assign new_P1_U4308 = ~new_P1_R1222_U98 | ~new_P1_U3026;
  assign new_P1_U4309 = ~new_P1_U3025 | ~new_P1_U3083;
  assign new_P1_U4310 = ~new_P1_R1282_U24 | ~new_P1_U3023;
  assign new_P1_U4311 = ~new_P1_U3476 | ~new_P1_U4142;
  assign new_P1_U4312 = ~new_P1_U3662 | ~new_P1_U4307;
  assign new_P1_U4313 = ~P1_REG2_REG_10_ | ~new_P1_U3018;
  assign new_P1_U4314 = ~P1_REG1_REG_10_ | ~new_P1_U3019;
  assign new_P1_U4315 = ~P1_REG0_REG_10_ | ~new_P1_U3020;
  assign new_P1_U4316 = ~new_P1_ADD_95_U78 | ~new_P1_U3017;
  assign new_P1_U4317 = ~new_P1_U3062;
  assign new_P1_U4318 = ~new_P1_U3033 | ~new_P1_U3084;
  assign new_P1_U4319 = ~new_P1_R1150_U102 | ~new_P1_U3961;
  assign new_P1_U4320 = ~new_P1_R1117_U102 | ~new_P1_U3963;
  assign new_P1_U4321 = ~new_P1_R1138_U97 | ~new_P1_U3962;
  assign new_P1_U4322 = ~new_P1_R1192_U102 | ~new_P1_U3959;
  assign new_P1_U4323 = ~new_P1_R1207_U102 | ~new_P1_U3958;
  assign new_P1_U4324 = ~new_P1_R1171_U97 | ~new_P1_U3968;
  assign new_P1_U4325 = ~new_P1_R1240_U97 | ~new_P1_U3967;
  assign new_P1_U4326 = ~new_P1_U3384;
  assign new_P1_U4327 = ~new_P1_R1222_U97 | ~new_P1_U3026;
  assign new_P1_U4328 = ~new_P1_U3025 | ~new_P1_U3062;
  assign new_P1_U4329 = ~new_P1_R1282_U63 | ~new_P1_U3023;
  assign new_P1_U4330 = ~new_P1_U3479 | ~new_P1_U4142;
  assign new_P1_U4331 = ~new_P1_U3666 | ~new_P1_U4326;
  assign new_P1_U4332 = ~P1_REG2_REG_11_ | ~new_P1_U3018;
  assign new_P1_U4333 = ~P1_REG1_REG_11_ | ~new_P1_U3019;
  assign new_P1_U4334 = ~P1_REG0_REG_11_ | ~new_P1_U3020;
  assign new_P1_U4335 = ~new_P1_ADD_95_U77 | ~new_P1_U3017;
  assign new_P1_U4336 = ~new_P1_U3063;
  assign new_P1_U4337 = ~new_P1_U3033 | ~new_P1_U3083;
  assign new_P1_U4338 = ~new_P1_R1150_U112 | ~new_P1_U3961;
  assign new_P1_U4339 = ~new_P1_R1117_U112 | ~new_P1_U3963;
  assign new_P1_U4340 = ~new_P1_R1138_U11 | ~new_P1_U3962;
  assign new_P1_U4341 = ~new_P1_R1192_U112 | ~new_P1_U3959;
  assign new_P1_U4342 = ~new_P1_R1207_U112 | ~new_P1_U3958;
  assign new_P1_U4343 = ~new_P1_R1171_U11 | ~new_P1_U3968;
  assign new_P1_U4344 = ~new_P1_R1240_U11 | ~new_P1_U3967;
  assign new_P1_U4345 = ~new_P1_U3385;
  assign new_P1_U4346 = ~new_P1_R1222_U11 | ~new_P1_U3026;
  assign new_P1_U4347 = ~new_P1_U3025 | ~new_P1_U3063;
  assign new_P1_U4348 = ~new_P1_R1282_U6 | ~new_P1_U3023;
  assign new_P1_U4349 = ~new_P1_U3482 | ~new_P1_U4142;
  assign new_P1_U4350 = ~new_P1_U3670 | ~new_P1_U4345;
  assign new_P1_U4351 = ~P1_REG2_REG_12_ | ~new_P1_U3018;
  assign new_P1_U4352 = ~P1_REG1_REG_12_ | ~new_P1_U3019;
  assign new_P1_U4353 = ~P1_REG0_REG_12_ | ~new_P1_U3020;
  assign new_P1_U4354 = ~new_P1_ADD_95_U76 | ~new_P1_U3017;
  assign new_P1_U4355 = ~new_P1_U3072;
  assign new_P1_U4356 = ~new_P1_U3033 | ~new_P1_U3062;
  assign new_P1_U4357 = ~new_P1_R1150_U10 | ~new_P1_U3961;
  assign new_P1_U4358 = ~new_P1_R1117_U10 | ~new_P1_U3963;
  assign new_P1_U4359 = ~new_P1_R1138_U115 | ~new_P1_U3962;
  assign new_P1_U4360 = ~new_P1_R1192_U10 | ~new_P1_U3959;
  assign new_P1_U4361 = ~new_P1_R1207_U10 | ~new_P1_U3958;
  assign new_P1_U4362 = ~new_P1_R1171_U115 | ~new_P1_U3968;
  assign new_P1_U4363 = ~new_P1_R1240_U115 | ~new_P1_U3967;
  assign new_P1_U4364 = ~new_P1_U3386;
  assign new_P1_U4365 = ~new_P1_R1222_U115 | ~new_P1_U3026;
  assign new_P1_U4366 = ~new_P1_U3025 | ~new_P1_U3072;
  assign new_P1_U4367 = ~new_P1_R1282_U7 | ~new_P1_U3023;
  assign new_P1_U4368 = ~new_P1_U3485 | ~new_P1_U4142;
  assign new_P1_U4369 = ~new_P1_U3674 | ~new_P1_U4364;
  assign new_P1_U4370 = ~P1_REG2_REG_13_ | ~new_P1_U3018;
  assign new_P1_U4371 = ~P1_REG1_REG_13_ | ~new_P1_U3019;
  assign new_P1_U4372 = ~P1_REG0_REG_13_ | ~new_P1_U3020;
  assign new_P1_U4373 = ~new_P1_ADD_95_U75 | ~new_P1_U3017;
  assign new_P1_U4374 = ~new_P1_U3080;
  assign new_P1_U4375 = ~new_P1_U3033 | ~new_P1_U3063;
  assign new_P1_U4376 = ~new_P1_R1150_U101 | ~new_P1_U3961;
  assign new_P1_U4377 = ~new_P1_R1117_U101 | ~new_P1_U3963;
  assign new_P1_U4378 = ~new_P1_R1138_U114 | ~new_P1_U3962;
  assign new_P1_U4379 = ~new_P1_R1192_U101 | ~new_P1_U3959;
  assign new_P1_U4380 = ~new_P1_R1207_U101 | ~new_P1_U3958;
  assign new_P1_U4381 = ~new_P1_R1171_U114 | ~new_P1_U3968;
  assign new_P1_U4382 = ~new_P1_R1240_U114 | ~new_P1_U3967;
  assign new_P1_U4383 = ~new_P1_U3387;
  assign new_P1_U4384 = ~new_P1_R1222_U114 | ~new_P1_U3026;
  assign new_P1_U4385 = ~new_P1_U3025 | ~new_P1_U3080;
  assign new_P1_U4386 = ~new_P1_R1282_U8 | ~new_P1_U3023;
  assign new_P1_U4387 = ~new_P1_U3488 | ~new_P1_U4142;
  assign new_P1_U4388 = ~new_P1_U3678 | ~new_P1_U4383;
  assign new_P1_U4389 = ~P1_REG2_REG_14_ | ~new_P1_U3018;
  assign new_P1_U4390 = ~P1_REG1_REG_14_ | ~new_P1_U3019;
  assign new_P1_U4391 = ~P1_REG0_REG_14_ | ~new_P1_U3020;
  assign new_P1_U4392 = ~new_P1_ADD_95_U74 | ~new_P1_U3017;
  assign new_P1_U4393 = ~new_P1_U3079;
  assign new_P1_U4394 = ~new_P1_U3033 | ~new_P1_U3072;
  assign new_P1_U4395 = ~new_P1_R1150_U100 | ~new_P1_U3961;
  assign new_P1_U4396 = ~new_P1_R1117_U100 | ~new_P1_U3963;
  assign new_P1_U4397 = ~new_P1_R1138_U12 | ~new_P1_U3962;
  assign new_P1_U4398 = ~new_P1_R1192_U100 | ~new_P1_U3959;
  assign new_P1_U4399 = ~new_P1_R1207_U100 | ~new_P1_U3958;
  assign new_P1_U4400 = ~new_P1_R1171_U12 | ~new_P1_U3968;
  assign new_P1_U4401 = ~new_P1_R1240_U12 | ~new_P1_U3967;
  assign new_P1_U4402 = ~new_P1_U3388;
  assign new_P1_U4403 = ~new_P1_R1222_U12 | ~new_P1_U3026;
  assign new_P1_U4404 = ~new_P1_U3025 | ~new_P1_U3079;
  assign new_P1_U4405 = ~new_P1_R1282_U86 | ~new_P1_U3023;
  assign new_P1_U4406 = ~new_P1_U3491 | ~new_P1_U4142;
  assign new_P1_U4407 = ~new_P1_U3682 | ~new_P1_U4402;
  assign new_P1_U4408 = ~P1_REG2_REG_15_ | ~new_P1_U3018;
  assign new_P1_U4409 = ~P1_REG1_REG_15_ | ~new_P1_U3019;
  assign new_P1_U4410 = ~P1_REG0_REG_15_ | ~new_P1_U3020;
  assign new_P1_U4411 = ~new_P1_ADD_95_U73 | ~new_P1_U3017;
  assign new_P1_U4412 = ~new_P1_U3074;
  assign new_P1_U4413 = ~new_P1_U3033 | ~new_P1_U3080;
  assign new_P1_U4414 = ~new_P1_R1150_U111 | ~new_P1_U3961;
  assign new_P1_U4415 = ~new_P1_R1117_U111 | ~new_P1_U3963;
  assign new_P1_U4416 = ~new_P1_R1138_U113 | ~new_P1_U3962;
  assign new_P1_U4417 = ~new_P1_R1192_U111 | ~new_P1_U3959;
  assign new_P1_U4418 = ~new_P1_R1207_U111 | ~new_P1_U3958;
  assign new_P1_U4419 = ~new_P1_R1171_U113 | ~new_P1_U3968;
  assign new_P1_U4420 = ~new_P1_R1240_U113 | ~new_P1_U3967;
  assign new_P1_U4421 = ~new_P1_U3389;
  assign new_P1_U4422 = ~new_P1_R1222_U113 | ~new_P1_U3026;
  assign new_P1_U4423 = ~new_P1_U3025 | ~new_P1_U3074;
  assign new_P1_U4424 = ~new_P1_R1282_U9 | ~new_P1_U3023;
  assign new_P1_U4425 = ~new_P1_U3494 | ~new_P1_U4142;
  assign new_P1_U4426 = ~new_P1_U3686 | ~new_P1_U4421;
  assign new_P1_U4427 = ~P1_REG2_REG_16_ | ~new_P1_U3018;
  assign new_P1_U4428 = ~P1_REG1_REG_16_ | ~new_P1_U3019;
  assign new_P1_U4429 = ~P1_REG0_REG_16_ | ~new_P1_U3020;
  assign new_P1_U4430 = ~new_P1_ADD_95_U72 | ~new_P1_U3017;
  assign new_P1_U4431 = ~new_P1_U3073;
  assign new_P1_U4432 = ~new_P1_U3033 | ~new_P1_U3079;
  assign new_P1_U4433 = ~new_P1_R1150_U110 | ~new_P1_U3961;
  assign new_P1_U4434 = ~new_P1_R1117_U110 | ~new_P1_U3963;
  assign new_P1_U4435 = ~new_P1_R1138_U112 | ~new_P1_U3962;
  assign new_P1_U4436 = ~new_P1_R1192_U110 | ~new_P1_U3959;
  assign new_P1_U4437 = ~new_P1_R1207_U110 | ~new_P1_U3958;
  assign new_P1_U4438 = ~new_P1_R1171_U112 | ~new_P1_U3968;
  assign new_P1_U4439 = ~new_P1_R1240_U112 | ~new_P1_U3967;
  assign new_P1_U4440 = ~new_P1_U3390;
  assign new_P1_U4441 = ~new_P1_R1222_U112 | ~new_P1_U3026;
  assign new_P1_U4442 = ~new_P1_U3025 | ~new_P1_U3073;
  assign new_P1_U4443 = ~new_P1_R1282_U10 | ~new_P1_U3023;
  assign new_P1_U4444 = ~new_P1_U3497 | ~new_P1_U4142;
  assign new_P1_U4445 = ~new_P1_U3690 | ~new_P1_U4440;
  assign new_P1_U4446 = ~P1_REG2_REG_17_ | ~new_P1_U3018;
  assign new_P1_U4447 = ~P1_REG1_REG_17_ | ~new_P1_U3019;
  assign new_P1_U4448 = ~P1_REG0_REG_17_ | ~new_P1_U3020;
  assign new_P1_U4449 = ~new_P1_ADD_95_U71 | ~new_P1_U3017;
  assign new_P1_U4450 = ~new_P1_U3069;
  assign new_P1_U4451 = ~new_P1_U3033 | ~new_P1_U3074;
  assign new_P1_U4452 = ~new_P1_R1150_U11 | ~new_P1_U3961;
  assign new_P1_U4453 = ~new_P1_R1117_U11 | ~new_P1_U3963;
  assign new_P1_U4454 = ~new_P1_R1138_U111 | ~new_P1_U3962;
  assign new_P1_U4455 = ~new_P1_R1192_U11 | ~new_P1_U3959;
  assign new_P1_U4456 = ~new_P1_R1207_U11 | ~new_P1_U3958;
  assign new_P1_U4457 = ~new_P1_R1171_U111 | ~new_P1_U3968;
  assign new_P1_U4458 = ~new_P1_R1240_U111 | ~new_P1_U3967;
  assign new_P1_U4459 = ~new_P1_U3391;
  assign new_P1_U4460 = ~new_P1_R1222_U111 | ~new_P1_U3026;
  assign new_P1_U4461 = ~new_P1_U3025 | ~new_P1_U3069;
  assign new_P1_U4462 = ~new_P1_R1282_U11 | ~new_P1_U3023;
  assign new_P1_U4463 = ~new_P1_U3500 | ~new_P1_U4142;
  assign new_P1_U4464 = ~new_P1_U3694 | ~new_P1_U4459;
  assign new_P1_U4465 = ~P1_REG2_REG_18_ | ~new_P1_U3018;
  assign new_P1_U4466 = ~P1_REG1_REG_18_ | ~new_P1_U3019;
  assign new_P1_U4467 = ~P1_REG0_REG_18_ | ~new_P1_U3020;
  assign new_P1_U4468 = ~new_P1_ADD_95_U70 | ~new_P1_U3017;
  assign new_P1_U4469 = ~new_P1_U3082;
  assign new_P1_U4470 = ~new_P1_U3033 | ~new_P1_U3073;
  assign new_P1_U4471 = ~new_P1_R1150_U99 | ~new_P1_U3961;
  assign new_P1_U4472 = ~new_P1_R1117_U99 | ~new_P1_U3963;
  assign new_P1_U4473 = ~new_P1_R1138_U13 | ~new_P1_U3962;
  assign new_P1_U4474 = ~new_P1_R1192_U99 | ~new_P1_U3959;
  assign new_P1_U4475 = ~new_P1_R1207_U99 | ~new_P1_U3958;
  assign new_P1_U4476 = ~new_P1_R1171_U13 | ~new_P1_U3968;
  assign new_P1_U4477 = ~new_P1_R1240_U13 | ~new_P1_U3967;
  assign new_P1_U4478 = ~new_P1_U3392;
  assign new_P1_U4479 = ~new_P1_R1222_U13 | ~new_P1_U3026;
  assign new_P1_U4480 = ~new_P1_U3025 | ~new_P1_U3082;
  assign new_P1_U4481 = ~new_P1_R1282_U84 | ~new_P1_U3023;
  assign new_P1_U4482 = ~new_P1_U3503 | ~new_P1_U4142;
  assign new_P1_U4483 = ~new_P1_U3698 | ~new_P1_U4478;
  assign new_P1_U4484 = ~P1_REG2_REG_19_ | ~new_P1_U3018;
  assign new_P1_U4485 = ~P1_REG1_REG_19_ | ~new_P1_U3019;
  assign new_P1_U4486 = ~P1_REG0_REG_19_ | ~new_P1_U3020;
  assign new_P1_U4487 = ~new_P1_ADD_95_U69 | ~new_P1_U3017;
  assign new_P1_U4488 = ~new_P1_U3081;
  assign new_P1_U4489 = ~new_P1_U3033 | ~new_P1_U3069;
  assign new_P1_U4490 = ~new_P1_R1150_U98 | ~new_P1_U3961;
  assign new_P1_U4491 = ~new_P1_R1117_U98 | ~new_P1_U3963;
  assign new_P1_U4492 = ~new_P1_R1138_U110 | ~new_P1_U3962;
  assign new_P1_U4493 = ~new_P1_R1192_U98 | ~new_P1_U3959;
  assign new_P1_U4494 = ~new_P1_R1207_U98 | ~new_P1_U3958;
  assign new_P1_U4495 = ~new_P1_R1171_U110 | ~new_P1_U3968;
  assign new_P1_U4496 = ~new_P1_R1240_U110 | ~new_P1_U3967;
  assign new_P1_U4497 = ~new_P1_U3393;
  assign new_P1_U4498 = ~new_P1_R1222_U110 | ~new_P1_U3026;
  assign new_P1_U4499 = ~new_P1_U3025 | ~new_P1_U3081;
  assign new_P1_U4500 = ~new_P1_R1282_U12 | ~new_P1_U3023;
  assign new_P1_U4501 = ~new_P1_U3506 | ~new_P1_U4142;
  assign new_P1_U4502 = ~new_P1_U3702 | ~new_P1_U4497;
  assign new_P1_U4503 = ~P1_REG2_REG_20_ | ~new_P1_U3018;
  assign new_P1_U4504 = ~P1_REG1_REG_20_ | ~new_P1_U3019;
  assign new_P1_U4505 = ~P1_REG0_REG_20_ | ~new_P1_U3020;
  assign new_P1_U4506 = ~new_P1_ADD_95_U68 | ~new_P1_U3017;
  assign new_P1_U4507 = ~new_P1_U3076;
  assign new_P1_U4508 = ~new_P1_U3033 | ~new_P1_U3082;
  assign new_P1_U4509 = ~new_P1_R1150_U97 | ~new_P1_U3961;
  assign new_P1_U4510 = ~new_P1_R1117_U97 | ~new_P1_U3963;
  assign new_P1_U4511 = ~new_P1_R1138_U109 | ~new_P1_U3962;
  assign new_P1_U4512 = ~new_P1_R1192_U97 | ~new_P1_U3959;
  assign new_P1_U4513 = ~new_P1_R1207_U97 | ~new_P1_U3958;
  assign new_P1_U4514 = ~new_P1_R1171_U109 | ~new_P1_U3968;
  assign new_P1_U4515 = ~new_P1_R1240_U109 | ~new_P1_U3967;
  assign new_P1_U4516 = ~new_P1_U3394;
  assign new_P1_U4517 = ~new_P1_R1222_U109 | ~new_P1_U3026;
  assign new_P1_U4518 = ~new_P1_U3025 | ~new_P1_U3076;
  assign new_P1_U4519 = ~new_P1_R1282_U82 | ~new_P1_U3023;
  assign new_P1_U4520 = ~new_P1_U3508 | ~new_P1_U4142;
  assign new_P1_U4521 = ~new_P1_U3706 | ~new_P1_U4516;
  assign new_P1_U4522 = ~P1_REG2_REG_21_ | ~new_P1_U3018;
  assign new_P1_U4523 = ~P1_REG1_REG_21_ | ~new_P1_U3019;
  assign new_P1_U4524 = ~P1_REG0_REG_21_ | ~new_P1_U3020;
  assign new_P1_U4525 = ~new_P1_ADD_95_U67 | ~new_P1_U3017;
  assign new_P1_U4526 = ~new_P1_U3075;
  assign new_P1_U4527 = ~new_P1_U3033 | ~new_P1_U3081;
  assign new_P1_U4528 = ~new_P1_R1150_U95 | ~new_P1_U3961;
  assign new_P1_U4529 = ~new_P1_R1117_U95 | ~new_P1_U3963;
  assign new_P1_U4530 = ~new_P1_R1138_U14 | ~new_P1_U3962;
  assign new_P1_U4531 = ~new_P1_R1192_U95 | ~new_P1_U3959;
  assign new_P1_U4532 = ~new_P1_R1207_U95 | ~new_P1_U3958;
  assign new_P1_U4533 = ~new_P1_R1171_U14 | ~new_P1_U3968;
  assign new_P1_U4534 = ~new_P1_R1240_U14 | ~new_P1_U3967;
  assign new_P1_U4535 = ~new_P1_U3396;
  assign new_P1_U4536 = ~new_P1_R1222_U14 | ~new_P1_U3026;
  assign new_P1_U4537 = ~new_P1_U3025 | ~new_P1_U3075;
  assign new_P1_U4538 = ~new_P1_R1282_U13 | ~new_P1_U3023;
  assign new_P1_U4539 = ~new_P1_U3982 | ~new_P1_U4142;
  assign new_P1_U4540 = ~new_P1_U3710 | ~new_P1_U4535;
  assign new_P1_U4541 = ~P1_REG2_REG_22_ | ~new_P1_U3018;
  assign new_P1_U4542 = ~P1_REG1_REG_22_ | ~new_P1_U3019;
  assign new_P1_U4543 = ~P1_REG0_REG_22_ | ~new_P1_U3020;
  assign new_P1_U4544 = ~new_P1_ADD_95_U66 | ~new_P1_U3017;
  assign new_P1_U4545 = ~new_P1_U3061;
  assign new_P1_U4546 = ~new_P1_U3033 | ~new_P1_U3076;
  assign new_P1_U4547 = ~new_P1_R1150_U109 | ~new_P1_U3961;
  assign new_P1_U4548 = ~new_P1_R1117_U109 | ~new_P1_U3963;
  assign new_P1_U4549 = ~new_P1_R1138_U15 | ~new_P1_U3962;
  assign new_P1_U4550 = ~new_P1_R1192_U109 | ~new_P1_U3959;
  assign new_P1_U4551 = ~new_P1_R1207_U109 | ~new_P1_U3958;
  assign new_P1_U4552 = ~new_P1_R1171_U15 | ~new_P1_U3968;
  assign new_P1_U4553 = ~new_P1_R1240_U15 | ~new_P1_U3967;
  assign new_P1_U4554 = ~new_P1_U3398;
  assign new_P1_U4555 = ~new_P1_R1222_U15 | ~new_P1_U3026;
  assign new_P1_U4556 = ~new_P1_U3025 | ~new_P1_U3061;
  assign new_P1_U4557 = ~new_P1_R1282_U78 | ~new_P1_U3023;
  assign new_P1_U4558 = ~new_P1_U3981 | ~new_P1_U4142;
  assign new_P1_U4559 = ~new_P1_U3714 | ~new_P1_U4554;
  assign new_P1_U4560 = ~P1_REG2_REG_23_ | ~new_P1_U3018;
  assign new_P1_U4561 = ~P1_REG1_REG_23_ | ~new_P1_U3019;
  assign new_P1_U4562 = ~P1_REG0_REG_23_ | ~new_P1_U3020;
  assign new_P1_U4563 = ~new_P1_ADD_95_U65 | ~new_P1_U3017;
  assign new_P1_U4564 = ~new_P1_U3066;
  assign new_P1_U4565 = ~new_P1_U3033 | ~new_P1_U3075;
  assign new_P1_U4566 = ~new_P1_R1150_U108 | ~new_P1_U3961;
  assign new_P1_U4567 = ~new_P1_R1117_U108 | ~new_P1_U3963;
  assign new_P1_U4568 = ~new_P1_R1138_U108 | ~new_P1_U3962;
  assign new_P1_U4569 = ~new_P1_R1192_U108 | ~new_P1_U3959;
  assign new_P1_U4570 = ~new_P1_R1207_U108 | ~new_P1_U3958;
  assign new_P1_U4571 = ~new_P1_R1171_U108 | ~new_P1_U3968;
  assign new_P1_U4572 = ~new_P1_R1240_U108 | ~new_P1_U3967;
  assign new_P1_U4573 = ~new_P1_U3400;
  assign new_P1_U4574 = ~new_P1_R1222_U108 | ~new_P1_U3026;
  assign new_P1_U4575 = ~new_P1_U3025 | ~new_P1_U3066;
  assign new_P1_U4576 = ~new_P1_R1282_U14 | ~new_P1_U3023;
  assign new_P1_U4577 = ~new_P1_U3980 | ~new_P1_U4142;
  assign new_P1_U4578 = ~new_P1_U3718 | ~new_P1_U4573;
  assign new_P1_U4579 = ~P1_REG2_REG_24_ | ~new_P1_U3018;
  assign new_P1_U4580 = ~P1_REG1_REG_24_ | ~new_P1_U3019;
  assign new_P1_U4581 = ~P1_REG0_REG_24_ | ~new_P1_U3020;
  assign new_P1_U4582 = ~new_P1_ADD_95_U64 | ~new_P1_U3017;
  assign new_P1_U4583 = ~new_P1_U3065;
  assign new_P1_U4584 = ~new_P1_U3033 | ~new_P1_U3061;
  assign new_P1_U4585 = ~new_P1_R1150_U12 | ~new_P1_U3961;
  assign new_P1_U4586 = ~new_P1_R1117_U12 | ~new_P1_U3963;
  assign new_P1_U4587 = ~new_P1_R1138_U107 | ~new_P1_U3962;
  assign new_P1_U4588 = ~new_P1_R1192_U12 | ~new_P1_U3959;
  assign new_P1_U4589 = ~new_P1_R1207_U12 | ~new_P1_U3958;
  assign new_P1_U4590 = ~new_P1_R1171_U107 | ~new_P1_U3968;
  assign new_P1_U4591 = ~new_P1_R1240_U107 | ~new_P1_U3967;
  assign new_P1_U4592 = ~new_P1_U3402;
  assign new_P1_U4593 = ~new_P1_R1222_U107 | ~new_P1_U3026;
  assign new_P1_U4594 = ~new_P1_U3025 | ~new_P1_U3065;
  assign new_P1_U4595 = ~new_P1_R1282_U76 | ~new_P1_U3023;
  assign new_P1_U4596 = ~new_P1_U3979 | ~new_P1_U4142;
  assign new_P1_U4597 = ~new_P1_U3722 | ~new_P1_U4592;
  assign new_P1_U4598 = ~P1_REG2_REG_25_ | ~new_P1_U3018;
  assign new_P1_U4599 = ~P1_REG1_REG_25_ | ~new_P1_U3019;
  assign new_P1_U4600 = ~P1_REG0_REG_25_ | ~new_P1_U3020;
  assign new_P1_U4601 = ~new_P1_ADD_95_U63 | ~new_P1_U3017;
  assign new_P1_U4602 = ~new_P1_U3058;
  assign new_P1_U4603 = ~new_P1_U3033 | ~new_P1_U3066;
  assign new_P1_U4604 = ~new_P1_R1150_U94 | ~new_P1_U3961;
  assign new_P1_U4605 = ~new_P1_R1117_U94 | ~new_P1_U3963;
  assign new_P1_U4606 = ~new_P1_R1138_U106 | ~new_P1_U3962;
  assign new_P1_U4607 = ~new_P1_R1192_U94 | ~new_P1_U3959;
  assign new_P1_U4608 = ~new_P1_R1207_U94 | ~new_P1_U3958;
  assign new_P1_U4609 = ~new_P1_R1171_U106 | ~new_P1_U3968;
  assign new_P1_U4610 = ~new_P1_R1240_U106 | ~new_P1_U3967;
  assign new_P1_U4611 = ~new_P1_U3404;
  assign new_P1_U4612 = ~new_P1_R1222_U106 | ~new_P1_U3026;
  assign new_P1_U4613 = ~new_P1_U3025 | ~new_P1_U3058;
  assign new_P1_U4614 = ~new_P1_R1282_U15 | ~new_P1_U3023;
  assign new_P1_U4615 = ~new_P1_U3978 | ~new_P1_U4142;
  assign new_P1_U4616 = ~new_P1_U3726 | ~new_P1_U4611;
  assign new_P1_U4617 = ~P1_REG2_REG_26_ | ~new_P1_U3018;
  assign new_P1_U4618 = ~P1_REG1_REG_26_ | ~new_P1_U3019;
  assign new_P1_U4619 = ~P1_REG0_REG_26_ | ~new_P1_U3020;
  assign new_P1_U4620 = ~new_P1_ADD_95_U62 | ~new_P1_U3017;
  assign new_P1_U4621 = ~new_P1_U3057;
  assign new_P1_U4622 = ~new_P1_U3033 | ~new_P1_U3065;
  assign new_P1_U4623 = ~new_P1_R1150_U93 | ~new_P1_U3961;
  assign new_P1_U4624 = ~new_P1_R1117_U93 | ~new_P1_U3963;
  assign new_P1_U4625 = ~new_P1_R1138_U105 | ~new_P1_U3962;
  assign new_P1_U4626 = ~new_P1_R1192_U93 | ~new_P1_U3959;
  assign new_P1_U4627 = ~new_P1_R1207_U93 | ~new_P1_U3958;
  assign new_P1_U4628 = ~new_P1_R1171_U105 | ~new_P1_U3968;
  assign new_P1_U4629 = ~new_P1_R1240_U105 | ~new_P1_U3967;
  assign new_P1_U4630 = ~new_P1_U3406;
  assign new_P1_U4631 = ~new_P1_R1222_U105 | ~new_P1_U3026;
  assign new_P1_U4632 = ~new_P1_U3025 | ~new_P1_U3057;
  assign new_P1_U4633 = ~new_P1_R1282_U74 | ~new_P1_U3023;
  assign new_P1_U4634 = ~new_P1_U3977 | ~new_P1_U4142;
  assign new_P1_U4635 = ~new_P1_U3730 | ~new_P1_U4630;
  assign new_P1_U4636 = ~P1_REG2_REG_27_ | ~new_P1_U3018;
  assign new_P1_U4637 = ~P1_REG1_REG_27_ | ~new_P1_U3019;
  assign new_P1_U4638 = ~P1_REG0_REG_27_ | ~new_P1_U3020;
  assign new_P1_U4639 = ~new_P1_ADD_95_U61 | ~new_P1_U3017;
  assign new_P1_U4640 = ~new_P1_U3053;
  assign new_P1_U4641 = ~new_P1_U3033 | ~new_P1_U3058;
  assign new_P1_U4642 = ~new_P1_R1150_U107 | ~new_P1_U3961;
  assign new_P1_U4643 = ~new_P1_R1117_U107 | ~new_P1_U3963;
  assign new_P1_U4644 = ~new_P1_R1138_U16 | ~new_P1_U3962;
  assign new_P1_U4645 = ~new_P1_R1192_U107 | ~new_P1_U3959;
  assign new_P1_U4646 = ~new_P1_R1207_U107 | ~new_P1_U3958;
  assign new_P1_U4647 = ~new_P1_R1171_U16 | ~new_P1_U3968;
  assign new_P1_U4648 = ~new_P1_R1240_U16 | ~new_P1_U3967;
  assign new_P1_U4649 = ~new_P1_U3408;
  assign new_P1_U4650 = ~new_P1_R1222_U16 | ~new_P1_U3026;
  assign new_P1_U4651 = ~new_P1_U3025 | ~new_P1_U3053;
  assign new_P1_U4652 = ~new_P1_R1282_U16 | ~new_P1_U3023;
  assign new_P1_U4653 = ~new_P1_U3976 | ~new_P1_U4142;
  assign new_P1_U4654 = ~new_P1_U3734 | ~new_P1_U4649;
  assign new_P1_U4655 = ~P1_REG2_REG_28_ | ~new_P1_U3018;
  assign new_P1_U4656 = ~P1_REG1_REG_28_ | ~new_P1_U3019;
  assign new_P1_U4657 = ~P1_REG0_REG_28_ | ~new_P1_U3020;
  assign new_P1_U4658 = ~new_P1_ADD_95_U60 | ~new_P1_U3017;
  assign new_P1_U4659 = ~new_P1_U3054;
  assign new_P1_U4660 = ~new_P1_U3033 | ~new_P1_U3057;
  assign new_P1_U4661 = ~new_P1_R1150_U13 | ~new_P1_U3961;
  assign new_P1_U4662 = ~new_P1_R1117_U13 | ~new_P1_U3963;
  assign new_P1_U4663 = ~new_P1_R1138_U104 | ~new_P1_U3962;
  assign new_P1_U4664 = ~new_P1_R1192_U13 | ~new_P1_U3959;
  assign new_P1_U4665 = ~new_P1_R1207_U13 | ~new_P1_U3958;
  assign new_P1_U4666 = ~new_P1_R1171_U104 | ~new_P1_U3968;
  assign new_P1_U4667 = ~new_P1_R1240_U104 | ~new_P1_U3967;
  assign new_P1_U4668 = ~new_P1_U3410;
  assign new_P1_U4669 = ~new_P1_R1222_U104 | ~new_P1_U3026;
  assign new_P1_U4670 = ~new_P1_U3025 | ~new_P1_U3054;
  assign new_P1_U4671 = ~new_P1_R1282_U72 | ~new_P1_U3023;
  assign new_P1_U4672 = ~new_P1_U3975 | ~new_P1_U4142;
  assign new_P1_U4673 = ~new_P1_U3738 | ~new_P1_U4668;
  assign new_P1_U4674 = ~new_P1_ADD_95_U5 | ~new_P1_U3017;
  assign new_P1_U4675 = ~P1_REG2_REG_29_ | ~new_P1_U3018;
  assign new_P1_U4676 = ~P1_REG1_REG_29_ | ~new_P1_U3019;
  assign new_P1_U4677 = ~P1_REG0_REG_29_ | ~new_P1_U3020;
  assign new_P1_U4678 = ~new_P1_U3055;
  assign new_P1_U4679 = ~new_P1_U3033 | ~new_P1_U3053;
  assign new_P1_U4680 = ~new_P1_R1150_U92 | ~new_P1_U3961;
  assign new_P1_U4681 = ~new_P1_R1117_U92 | ~new_P1_U3963;
  assign new_P1_U4682 = ~new_P1_R1138_U103 | ~new_P1_U3962;
  assign new_P1_U4683 = ~new_P1_R1192_U92 | ~new_P1_U3959;
  assign new_P1_U4684 = ~new_P1_R1207_U92 | ~new_P1_U3958;
  assign new_P1_U4685 = ~new_P1_R1171_U103 | ~new_P1_U3968;
  assign new_P1_U4686 = ~new_P1_R1240_U103 | ~new_P1_U3967;
  assign new_P1_U4687 = ~new_P1_U3412;
  assign new_P1_U4688 = ~new_P1_R1222_U103 | ~new_P1_U3026;
  assign new_P1_U4689 = ~new_P1_U3025 | ~new_P1_U3055;
  assign new_P1_U4690 = ~new_P1_R1282_U17 | ~new_P1_U3023;
  assign new_P1_U4691 = ~new_P1_U3974 | ~new_P1_U4142;
  assign new_P1_U4692 = ~new_P1_U3742 | ~new_P1_U4687;
  assign new_P1_U4693 = ~P1_REG2_REG_30_ | ~new_P1_U3018;
  assign new_P1_U4694 = ~P1_REG1_REG_30_ | ~new_P1_U3019;
  assign new_P1_U4695 = ~P1_REG0_REG_30_ | ~new_P1_U3020;
  assign new_P1_U4696 = ~new_P1_U3059;
  assign new_P1_U4697 = ~new_P1_U5699 | ~new_P1_U3359;
  assign new_P1_U4698 = ~new_P1_U3912 | ~new_P1_U4697;
  assign new_P1_U4699 = ~new_P1_U3743 | ~new_P1_U3059;
  assign new_P1_U4700 = ~new_P1_U3033 | ~new_P1_U3054;
  assign new_P1_U4701 = ~new_P1_R1150_U14 | ~new_P1_U3961;
  assign new_P1_U4702 = ~new_P1_R1117_U14 | ~new_P1_U3963;
  assign new_P1_U4703 = ~new_P1_R1138_U102 | ~new_P1_U3962;
  assign new_P1_U4704 = ~new_P1_R1192_U14 | ~new_P1_U3959;
  assign new_P1_U4705 = ~new_P1_R1207_U14 | ~new_P1_U3958;
  assign new_P1_U4706 = ~new_P1_R1171_U102 | ~new_P1_U3968;
  assign new_P1_U4707 = ~new_P1_R1240_U102 | ~new_P1_U3967;
  assign new_P1_U4708 = ~new_P1_U3801 | ~new_P1_U3802 | ~new_P1_U3051;
  assign new_P1_U4709 = ~new_P1_R1222_U102 | ~new_P1_U3026;
  assign new_P1_U4710 = ~new_P1_R1282_U70 | ~new_P1_U3023;
  assign new_P1_U4711 = ~new_P1_U3985 | ~new_P1_U4142;
  assign new_P1_U4712 = ~new_P1_U3744 | ~new_P1_U3745 | ~new_P1_U3746 | ~new_P1_U3051;
  assign new_P1_U4713 = ~P1_REG2_REG_31_ | ~new_P1_U3018;
  assign new_P1_U4714 = ~P1_REG1_REG_31_ | ~new_P1_U3019;
  assign new_P1_U4715 = ~P1_REG0_REG_31_ | ~new_P1_U3020;
  assign new_P1_U4716 = ~new_P1_U3056;
  assign new_P1_U4717 = ~new_P1_R1282_U19 | ~new_P1_U3023;
  assign new_P1_U4718 = ~new_P1_U3984 | ~new_P1_U4142;
  assign new_P1_U4719 = ~new_P1_U4717 | ~new_P1_U4718 | ~new_P1_U3945;
  assign new_P1_U4720 = ~new_P1_R1282_U68 | ~new_P1_U3023;
  assign new_P1_U4721 = ~new_P1_U3983 | ~new_P1_U4142;
  assign new_P1_U4722 = ~new_P1_U4720 | ~new_P1_U4721 | ~new_P1_U3945;
  assign new_P1_U4723 = ~new_P1_U3749 | ~new_P1_U3016;
  assign new_P1_U4724 = ~new_P1_U3418 | ~new_P1_U4723;
  assign new_P1_U4725 = ~new_P1_U3988 | ~new_P1_U3441;
  assign new_P1_U4726 = ~new_P1_U3422;
  assign new_P1_U4727 = ~new_P1_U3035 | ~new_P1_U3078;
  assign new_P1_U4728 = ~new_P1_U3032 | ~P1_REG3_REG_0_;
  assign new_P1_U4729 = ~new_P1_U3031 | ~new_P1_R1222_U96;
  assign new_P1_U4730 = ~new_P1_U3030 | ~new_P1_U3450;
  assign new_P1_U4731 = ~new_P1_U3029 | ~new_P1_U3450;
  assign new_P1_U4732 = ~new_P1_U3035 | ~new_P1_U3068;
  assign new_P1_U4733 = ~new_P1_U3032 | ~P1_REG3_REG_1_;
  assign new_P1_U4734 = ~new_P1_U3031 | ~new_P1_R1222_U95;
  assign new_P1_U4735 = ~new_P1_U3030 | ~new_P1_U3455;
  assign new_P1_U4736 = ~new_P1_U3029 | ~new_P1_R1282_U57;
  assign new_P1_U4737 = ~new_P1_U3035 | ~new_P1_U3064;
  assign new_P1_U4738 = ~new_P1_U3032 | ~P1_REG3_REG_2_;
  assign new_P1_U4739 = ~new_P1_U3031 | ~new_P1_R1222_U17;
  assign new_P1_U4740 = ~new_P1_U3030 | ~new_P1_U3458;
  assign new_P1_U4741 = ~new_P1_U3029 | ~new_P1_R1282_U18;
  assign new_P1_U4742 = ~new_P1_U3035 | ~new_P1_U3060;
  assign new_P1_U4743 = ~new_P1_U3032 | ~new_P1_ADD_95_U4;
  assign new_P1_U4744 = ~new_P1_U3031 | ~new_P1_R1222_U101;
  assign new_P1_U4745 = ~new_P1_U3030 | ~new_P1_U3461;
  assign new_P1_U4746 = ~new_P1_U3029 | ~new_P1_R1282_U20;
  assign new_P1_U4747 = ~new_P1_U3035 | ~new_P1_U3067;
  assign new_P1_U4748 = ~new_P1_U3032 | ~new_P1_ADD_95_U59;
  assign new_P1_U4749 = ~new_P1_U3031 | ~new_P1_R1222_U100;
  assign new_P1_U4750 = ~new_P1_U3030 | ~new_P1_U3464;
  assign new_P1_U4751 = ~new_P1_U3029 | ~new_P1_R1282_U21;
  assign new_P1_U4752 = ~new_P1_U3035 | ~new_P1_U3071;
  assign new_P1_U4753 = ~new_P1_U3032 | ~new_P1_ADD_95_U58;
  assign new_P1_U4754 = ~new_P1_U3031 | ~new_P1_R1222_U18;
  assign new_P1_U4755 = ~new_P1_U3030 | ~new_P1_U3467;
  assign new_P1_U4756 = ~new_P1_U3029 | ~new_P1_R1282_U65;
  assign new_P1_U4757 = ~new_P1_U3035 | ~new_P1_U3070;
  assign new_P1_U4758 = ~new_P1_U3032 | ~new_P1_ADD_95_U57;
  assign new_P1_U4759 = ~new_P1_U3031 | ~new_P1_R1222_U99;
  assign new_P1_U4760 = ~new_P1_U3030 | ~new_P1_U3470;
  assign new_P1_U4761 = ~new_P1_U3029 | ~new_P1_R1282_U22;
  assign new_P1_U4762 = ~new_P1_U3035 | ~new_P1_U3084;
  assign new_P1_U4763 = ~new_P1_U3032 | ~new_P1_ADD_95_U56;
  assign new_P1_U4764 = ~new_P1_U3031 | ~new_P1_R1222_U19;
  assign new_P1_U4765 = ~new_P1_U3030 | ~new_P1_U3473;
  assign new_P1_U4766 = ~new_P1_U3029 | ~new_P1_R1282_U23;
  assign new_P1_U4767 = ~new_P1_U3035 | ~new_P1_U3083;
  assign new_P1_U4768 = ~new_P1_U3032 | ~new_P1_ADD_95_U55;
  assign new_P1_U4769 = ~new_P1_U3031 | ~new_P1_R1222_U98;
  assign new_P1_U4770 = ~new_P1_U3030 | ~new_P1_U3476;
  assign new_P1_U4771 = ~new_P1_U3029 | ~new_P1_R1282_U24;
  assign new_P1_U4772 = ~new_P1_U3035 | ~new_P1_U3062;
  assign new_P1_U4773 = ~new_P1_U3032 | ~new_P1_ADD_95_U54;
  assign new_P1_U4774 = ~new_P1_U3031 | ~new_P1_R1222_U97;
  assign new_P1_U4775 = ~new_P1_U3030 | ~new_P1_U3479;
  assign new_P1_U4776 = ~new_P1_U3029 | ~new_P1_R1282_U63;
  assign new_P1_U4777 = ~new_P1_U3035 | ~new_P1_U3063;
  assign new_P1_U4778 = ~new_P1_U3032 | ~new_P1_ADD_95_U78;
  assign new_P1_U4779 = ~new_P1_U3031 | ~new_P1_R1222_U11;
  assign new_P1_U4780 = ~new_P1_U3030 | ~new_P1_U3482;
  assign new_P1_U4781 = ~new_P1_U3029 | ~new_P1_R1282_U6;
  assign new_P1_U4782 = ~new_P1_U3035 | ~new_P1_U3072;
  assign new_P1_U4783 = ~new_P1_U3032 | ~new_P1_ADD_95_U77;
  assign new_P1_U4784 = ~new_P1_U3031 | ~new_P1_R1222_U115;
  assign new_P1_U4785 = ~new_P1_U3030 | ~new_P1_U3485;
  assign new_P1_U4786 = ~new_P1_U3029 | ~new_P1_R1282_U7;
  assign new_P1_U4787 = ~new_P1_U3035 | ~new_P1_U3080;
  assign new_P1_U4788 = ~new_P1_U3032 | ~new_P1_ADD_95_U76;
  assign new_P1_U4789 = ~new_P1_U3031 | ~new_P1_R1222_U114;
  assign new_P1_U4790 = ~new_P1_U3030 | ~new_P1_U3488;
  assign new_P1_U4791 = ~new_P1_U3029 | ~new_P1_R1282_U8;
  assign new_P1_U4792 = ~new_P1_U3035 | ~new_P1_U3079;
  assign new_P1_U4793 = ~new_P1_U3032 | ~new_P1_ADD_95_U75;
  assign new_P1_U4794 = ~new_P1_U3031 | ~new_P1_R1222_U12;
  assign new_P1_U4795 = ~new_P1_U3030 | ~new_P1_U3491;
  assign new_P1_U4796 = ~new_P1_U3029 | ~new_P1_R1282_U86;
  assign new_P1_U4797 = ~new_P1_U3035 | ~new_P1_U3074;
  assign new_P1_U4798 = ~new_P1_U3032 | ~new_P1_ADD_95_U74;
  assign new_P1_U4799 = ~new_P1_U3031 | ~new_P1_R1222_U113;
  assign new_P1_U4800 = ~new_P1_U3030 | ~new_P1_U3494;
  assign new_P1_U4801 = ~new_P1_U3029 | ~new_P1_R1282_U9;
  assign new_P1_U4802 = ~new_P1_U3035 | ~new_P1_U3073;
  assign new_P1_U4803 = ~new_P1_U3032 | ~new_P1_ADD_95_U73;
  assign new_P1_U4804 = ~new_P1_U3031 | ~new_P1_R1222_U112;
  assign new_P1_U4805 = ~new_P1_U3030 | ~new_P1_U3497;
  assign new_P1_U4806 = ~new_P1_U3029 | ~new_P1_R1282_U10;
  assign new_P1_U4807 = ~new_P1_U3035 | ~new_P1_U3069;
  assign new_P1_U4808 = ~new_P1_U3032 | ~new_P1_ADD_95_U72;
  assign new_P1_U4809 = ~new_P1_U3031 | ~new_P1_R1222_U111;
  assign new_P1_U4810 = ~new_P1_U3030 | ~new_P1_U3500;
  assign new_P1_U4811 = ~new_P1_U3029 | ~new_P1_R1282_U11;
  assign new_P1_U4812 = ~new_P1_U3035 | ~new_P1_U3082;
  assign new_P1_U4813 = ~new_P1_U3032 | ~new_P1_ADD_95_U71;
  assign new_P1_U4814 = ~new_P1_U3031 | ~new_P1_R1222_U13;
  assign new_P1_U4815 = ~new_P1_U3030 | ~new_P1_U3503;
  assign new_P1_U4816 = ~new_P1_U3029 | ~new_P1_R1282_U84;
  assign new_P1_U4817 = ~new_P1_U3035 | ~new_P1_U3081;
  assign new_P1_U4818 = ~new_P1_U3032 | ~new_P1_ADD_95_U70;
  assign new_P1_U4819 = ~new_P1_U3031 | ~new_P1_R1222_U110;
  assign new_P1_U4820 = ~new_P1_U3030 | ~new_P1_U3506;
  assign new_P1_U4821 = ~new_P1_U3029 | ~new_P1_R1282_U12;
  assign new_P1_U4822 = ~new_P1_U3035 | ~new_P1_U3076;
  assign new_P1_U4823 = ~new_P1_U3032 | ~new_P1_ADD_95_U69;
  assign new_P1_U4824 = ~new_P1_U3031 | ~new_P1_R1222_U109;
  assign new_P1_U4825 = ~new_P1_U3030 | ~new_P1_U3508;
  assign new_P1_U4826 = ~new_P1_U3029 | ~new_P1_R1282_U82;
  assign new_P1_U4827 = ~new_P1_U3035 | ~new_P1_U3075;
  assign new_P1_U4828 = ~new_P1_U3032 | ~new_P1_ADD_95_U68;
  assign new_P1_U4829 = ~new_P1_U3031 | ~new_P1_R1222_U14;
  assign new_P1_U4830 = ~new_P1_U3030 | ~new_P1_U3982;
  assign new_P1_U4831 = ~new_P1_U3029 | ~new_P1_R1282_U13;
  assign new_P1_U4832 = ~new_P1_U3035 | ~new_P1_U3061;
  assign new_P1_U4833 = ~new_P1_U3032 | ~new_P1_ADD_95_U67;
  assign new_P1_U4834 = ~new_P1_U3031 | ~new_P1_R1222_U15;
  assign new_P1_U4835 = ~new_P1_U3030 | ~new_P1_U3981;
  assign new_P1_U4836 = ~new_P1_U3029 | ~new_P1_R1282_U78;
  assign new_P1_U4837 = ~new_P1_U3035 | ~new_P1_U3066;
  assign new_P1_U4838 = ~new_P1_U3032 | ~new_P1_ADD_95_U66;
  assign new_P1_U4839 = ~new_P1_U3031 | ~new_P1_R1222_U108;
  assign new_P1_U4840 = ~new_P1_U3030 | ~new_P1_U3980;
  assign new_P1_U4841 = ~new_P1_U3029 | ~new_P1_R1282_U14;
  assign new_P1_U4842 = ~new_P1_U3035 | ~new_P1_U3065;
  assign new_P1_U4843 = ~new_P1_U3032 | ~new_P1_ADD_95_U65;
  assign new_P1_U4844 = ~new_P1_U3031 | ~new_P1_R1222_U107;
  assign new_P1_U4845 = ~new_P1_U3030 | ~new_P1_U3979;
  assign new_P1_U4846 = ~new_P1_U3029 | ~new_P1_R1282_U76;
  assign new_P1_U4847 = ~new_P1_U3035 | ~new_P1_U3058;
  assign new_P1_U4848 = ~new_P1_U3032 | ~new_P1_ADD_95_U64;
  assign new_P1_U4849 = ~new_P1_U3031 | ~new_P1_R1222_U106;
  assign new_P1_U4850 = ~new_P1_U3030 | ~new_P1_U3978;
  assign new_P1_U4851 = ~new_P1_U3029 | ~new_P1_R1282_U15;
  assign new_P1_U4852 = ~new_P1_U3035 | ~new_P1_U3057;
  assign new_P1_U4853 = ~new_P1_U3032 | ~new_P1_ADD_95_U63;
  assign new_P1_U4854 = ~new_P1_U3031 | ~new_P1_R1222_U105;
  assign new_P1_U4855 = ~new_P1_U3030 | ~new_P1_U3977;
  assign new_P1_U4856 = ~new_P1_U3029 | ~new_P1_R1282_U74;
  assign new_P1_U4857 = ~new_P1_U3035 | ~new_P1_U3053;
  assign new_P1_U4858 = ~new_P1_U3032 | ~new_P1_ADD_95_U62;
  assign new_P1_U4859 = ~new_P1_U3031 | ~new_P1_R1222_U16;
  assign new_P1_U4860 = ~new_P1_U3030 | ~new_P1_U3976;
  assign new_P1_U4861 = ~new_P1_U3029 | ~new_P1_R1282_U16;
  assign new_P1_U4862 = ~new_P1_U3035 | ~new_P1_U3054;
  assign new_P1_U4863 = ~new_P1_U3032 | ~new_P1_ADD_95_U61;
  assign new_P1_U4864 = ~new_P1_U3031 | ~new_P1_R1222_U104;
  assign new_P1_U4865 = ~new_P1_U3030 | ~new_P1_U3975;
  assign new_P1_U4866 = ~new_P1_U3029 | ~new_P1_R1282_U72;
  assign new_P1_U4867 = ~new_P1_U3035 | ~new_P1_U3055;
  assign new_P1_U4868 = ~new_P1_U3032 | ~new_P1_ADD_95_U60;
  assign new_P1_U4869 = ~new_P1_U3031 | ~new_P1_R1222_U103;
  assign new_P1_U4870 = ~new_P1_U3030 | ~new_P1_U3974;
  assign new_P1_U4871 = ~new_P1_U3029 | ~new_P1_R1282_U17;
  assign new_P1_U4872 = ~new_P1_U3032 | ~new_P1_ADD_95_U5;
  assign new_P1_U4873 = ~new_P1_U3031 | ~new_P1_R1222_U102;
  assign new_P1_U4874 = ~new_P1_U3030 | ~new_P1_U3985;
  assign new_P1_U4875 = ~new_P1_U3029 | ~new_P1_R1282_U70;
  assign new_P1_U4876 = ~new_P1_U3030 | ~new_P1_U3984;
  assign new_P1_U4877 = ~new_P1_U3029 | ~new_P1_R1282_U19;
  assign new_P1_U4878 = ~new_P1_U3030 | ~new_P1_U3983;
  assign new_P1_U4879 = ~new_P1_U3029 | ~new_P1_R1282_U68;
  assign new_P1_U4880 = ~new_P1_U3418 | ~new_P1_U4726 | ~new_P1_U3806 | ~new_P1_U3804 | ~new_P1_U3803;
  assign new_P1_U4881 = ~new_P1_R1105_U13 | ~new_P1_U3041;
  assign new_P1_U4882 = ~new_P1_U3039 | ~new_P1_U3442;
  assign new_P1_U4883 = ~new_P1_R1162_U13 | ~new_P1_U3037;
  assign new_P1_U4884 = ~new_P1_U4883 | ~new_P1_U4882 | ~new_P1_U4881;
  assign new_P1_U4885 = ~new_P1_U3046 | ~new_P1_U3373;
  assign new_P1_U4886 = ~new_P1_U5677 | ~new_P1_U4885;
  assign new_P1_U4887 = ~new_P1_U4886 | ~new_P1_U3912;
  assign new_P1_U4888 = ~n1335;
  assign new_P1_U4889 = ~new_P1_U3423;
  assign new_P1_U4890 = ~new_P1_U3043 | ~new_P1_U4884;
  assign new_P1_U4891 = ~new_P1_U3042 | ~new_P1_R1105_U13;
  assign new_P1_U4892 = ~P1_REG3_REG_19_ | ~n1330;
  assign new_P1_U4893 = ~new_P1_U3040 | ~new_P1_U3442;
  assign new_P1_U4894 = ~new_P1_U3038 | ~new_P1_R1162_U13;
  assign new_P1_U4895 = ~P1_ADDR_REG_19_ | ~new_P1_U4889;
  assign new_P1_U4896 = ~new_P1_R1105_U75 | ~new_P1_U3041;
  assign new_P1_U4897 = ~new_P1_U3039 | ~new_P1_U3505;
  assign new_P1_U4898 = ~new_P1_R1162_U75 | ~new_P1_U3037;
  assign new_P1_U4899 = ~new_P1_U4898 | ~new_P1_U4897 | ~new_P1_U4896;
  assign new_P1_U4900 = ~new_P1_U3043 | ~new_P1_U4899;
  assign new_P1_U4901 = ~new_P1_R1105_U75 | ~new_P1_U3042;
  assign new_P1_U4902 = ~P1_REG3_REG_18_ | ~n1330;
  assign new_P1_U4903 = ~new_P1_U3040 | ~new_P1_U3505;
  assign new_P1_U4904 = ~new_P1_R1162_U75 | ~new_P1_U3038;
  assign new_P1_U4905 = ~P1_ADDR_REG_18_ | ~new_P1_U4889;
  assign new_P1_U4906 = ~new_P1_R1105_U12 | ~new_P1_U3041;
  assign new_P1_U4907 = ~new_P1_U3039 | ~new_P1_U3502;
  assign new_P1_U4908 = ~new_P1_R1162_U12 | ~new_P1_U3037;
  assign new_P1_U4909 = ~new_P1_U4908 | ~new_P1_U4907 | ~new_P1_U4906;
  assign new_P1_U4910 = ~new_P1_U3043 | ~new_P1_U4909;
  assign new_P1_U4911 = ~new_P1_R1105_U12 | ~new_P1_U3042;
  assign new_P1_U4912 = ~P1_REG3_REG_17_ | ~n1330;
  assign new_P1_U4913 = ~new_P1_U3040 | ~new_P1_U3502;
  assign new_P1_U4914 = ~new_P1_R1162_U12 | ~new_P1_U3038;
  assign new_P1_U4915 = ~P1_ADDR_REG_17_ | ~new_P1_U4889;
  assign new_P1_U4916 = ~new_P1_R1105_U76 | ~new_P1_U3041;
  assign new_P1_U4917 = ~new_P1_U3039 | ~new_P1_U3499;
  assign new_P1_U4918 = ~new_P1_R1162_U76 | ~new_P1_U3037;
  assign new_P1_U4919 = ~new_P1_U4918 | ~new_P1_U4917 | ~new_P1_U4916;
  assign new_P1_U4920 = ~new_P1_U3043 | ~new_P1_U4919;
  assign new_P1_U4921 = ~new_P1_R1105_U76 | ~new_P1_U3042;
  assign new_P1_U4922 = ~P1_REG3_REG_16_ | ~n1330;
  assign new_P1_U4923 = ~new_P1_U3040 | ~new_P1_U3499;
  assign new_P1_U4924 = ~new_P1_R1162_U76 | ~new_P1_U3038;
  assign new_P1_U4925 = ~P1_ADDR_REG_16_ | ~new_P1_U4889;
  assign new_P1_U4926 = ~new_P1_R1105_U77 | ~new_P1_U3041;
  assign new_P1_U4927 = ~new_P1_U3039 | ~new_P1_U3496;
  assign new_P1_U4928 = ~new_P1_R1162_U77 | ~new_P1_U3037;
  assign new_P1_U4929 = ~new_P1_U4928 | ~new_P1_U4927 | ~new_P1_U4926;
  assign new_P1_U4930 = ~new_P1_U3043 | ~new_P1_U4929;
  assign new_P1_U4931 = ~new_P1_R1105_U77 | ~new_P1_U3042;
  assign new_P1_U4932 = ~P1_REG3_REG_15_ | ~n1330;
  assign new_P1_U4933 = ~new_P1_U3040 | ~new_P1_U3496;
  assign new_P1_U4934 = ~new_P1_R1162_U77 | ~new_P1_U3038;
  assign new_P1_U4935 = ~P1_ADDR_REG_15_ | ~new_P1_U4889;
  assign new_P1_U4936 = ~new_P1_R1105_U78 | ~new_P1_U3041;
  assign new_P1_U4937 = ~new_P1_U3039 | ~new_P1_U3493;
  assign new_P1_U4938 = ~new_P1_R1162_U78 | ~new_P1_U3037;
  assign new_P1_U4939 = ~new_P1_U4938 | ~new_P1_U4937 | ~new_P1_U4936;
  assign new_P1_U4940 = ~new_P1_U3043 | ~new_P1_U4939;
  assign new_P1_U4941 = ~new_P1_R1105_U78 | ~new_P1_U3042;
  assign new_P1_U4942 = ~P1_REG3_REG_14_ | ~n1330;
  assign new_P1_U4943 = ~new_P1_U3040 | ~new_P1_U3493;
  assign new_P1_U4944 = ~new_P1_R1162_U78 | ~new_P1_U3038;
  assign new_P1_U4945 = ~P1_ADDR_REG_14_ | ~new_P1_U4889;
  assign new_P1_U4946 = ~new_P1_R1105_U11 | ~new_P1_U3041;
  assign new_P1_U4947 = ~new_P1_U3039 | ~new_P1_U3490;
  assign new_P1_U4948 = ~new_P1_R1162_U11 | ~new_P1_U3037;
  assign new_P1_U4949 = ~new_P1_U4948 | ~new_P1_U4947 | ~new_P1_U4946;
  assign new_P1_U4950 = ~new_P1_U3043 | ~new_P1_U4949;
  assign new_P1_U4951 = ~new_P1_R1105_U11 | ~new_P1_U3042;
  assign new_P1_U4952 = ~P1_REG3_REG_13_ | ~n1330;
  assign new_P1_U4953 = ~new_P1_U3040 | ~new_P1_U3490;
  assign new_P1_U4954 = ~new_P1_R1162_U11 | ~new_P1_U3038;
  assign new_P1_U4955 = ~P1_ADDR_REG_13_ | ~new_P1_U4889;
  assign new_P1_U4956 = ~new_P1_R1105_U79 | ~new_P1_U3041;
  assign new_P1_U4957 = ~new_P1_U3039 | ~new_P1_U3487;
  assign new_P1_U4958 = ~new_P1_R1162_U79 | ~new_P1_U3037;
  assign new_P1_U4959 = ~new_P1_U4958 | ~new_P1_U4957 | ~new_P1_U4956;
  assign new_P1_U4960 = ~new_P1_U3043 | ~new_P1_U4959;
  assign new_P1_U4961 = ~new_P1_R1105_U79 | ~new_P1_U3042;
  assign new_P1_U4962 = ~P1_REG3_REG_12_ | ~n1330;
  assign new_P1_U4963 = ~new_P1_U3040 | ~new_P1_U3487;
  assign new_P1_U4964 = ~new_P1_R1162_U79 | ~new_P1_U3038;
  assign new_P1_U4965 = ~P1_ADDR_REG_12_ | ~new_P1_U4889;
  assign new_P1_U4966 = ~new_P1_R1105_U80 | ~new_P1_U3041;
  assign new_P1_U4967 = ~new_P1_U3039 | ~new_P1_U3484;
  assign new_P1_U4968 = ~new_P1_R1162_U80 | ~new_P1_U3037;
  assign new_P1_U4969 = ~new_P1_U4968 | ~new_P1_U4967 | ~new_P1_U4966;
  assign new_P1_U4970 = ~new_P1_U3043 | ~new_P1_U4969;
  assign new_P1_U4971 = ~new_P1_R1105_U80 | ~new_P1_U3042;
  assign new_P1_U4972 = ~P1_REG3_REG_11_ | ~n1330;
  assign new_P1_U4973 = ~new_P1_U3040 | ~new_P1_U3484;
  assign new_P1_U4974 = ~new_P1_R1162_U80 | ~new_P1_U3038;
  assign new_P1_U4975 = ~P1_ADDR_REG_11_ | ~new_P1_U4889;
  assign new_P1_U4976 = ~new_P1_R1105_U10 | ~new_P1_U3041;
  assign new_P1_U4977 = ~new_P1_U3039 | ~new_P1_U3481;
  assign new_P1_U4978 = ~new_P1_R1162_U10 | ~new_P1_U3037;
  assign new_P1_U4979 = ~new_P1_U4978 | ~new_P1_U4977 | ~new_P1_U4976;
  assign new_P1_U4980 = ~new_P1_U3043 | ~new_P1_U4979;
  assign new_P1_U4981 = ~new_P1_R1105_U10 | ~new_P1_U3042;
  assign new_P1_U4982 = ~P1_REG3_REG_10_ | ~n1330;
  assign new_P1_U4983 = ~new_P1_U3040 | ~new_P1_U3481;
  assign new_P1_U4984 = ~new_P1_R1162_U10 | ~new_P1_U3038;
  assign new_P1_U4985 = ~P1_ADDR_REG_10_ | ~new_P1_U4889;
  assign new_P1_U4986 = ~new_P1_R1105_U70 | ~new_P1_U3041;
  assign new_P1_U4987 = ~new_P1_U3039 | ~new_P1_U3478;
  assign new_P1_U4988 = ~new_P1_R1162_U70 | ~new_P1_U3037;
  assign new_P1_U4989 = ~new_P1_U4988 | ~new_P1_U4987 | ~new_P1_U4986;
  assign new_P1_U4990 = ~new_P1_U3043 | ~new_P1_U4989;
  assign new_P1_U4991 = ~new_P1_R1105_U70 | ~new_P1_U3042;
  assign new_P1_U4992 = ~P1_REG3_REG_9_ | ~n1330;
  assign new_P1_U4993 = ~new_P1_U3040 | ~new_P1_U3478;
  assign new_P1_U4994 = ~new_P1_R1162_U70 | ~new_P1_U3038;
  assign new_P1_U4995 = ~P1_ADDR_REG_9_ | ~new_P1_U4889;
  assign new_P1_U4996 = ~new_P1_R1105_U71 | ~new_P1_U3041;
  assign new_P1_U4997 = ~new_P1_U3039 | ~new_P1_U3475;
  assign new_P1_U4998 = ~new_P1_R1162_U71 | ~new_P1_U3037;
  assign new_P1_U4999 = ~new_P1_U4998 | ~new_P1_U4997 | ~new_P1_U4996;
  assign new_P1_U5000 = ~new_P1_U3043 | ~new_P1_U4999;
  assign new_P1_U5001 = ~new_P1_R1105_U71 | ~new_P1_U3042;
  assign new_P1_U5002 = ~P1_REG3_REG_8_ | ~n1330;
  assign new_P1_U5003 = ~new_P1_U3040 | ~new_P1_U3475;
  assign new_P1_U5004 = ~new_P1_R1162_U71 | ~new_P1_U3038;
  assign new_P1_U5005 = ~P1_ADDR_REG_8_ | ~new_P1_U4889;
  assign new_P1_U5006 = ~new_P1_R1105_U16 | ~new_P1_U3041;
  assign new_P1_U5007 = ~new_P1_U3039 | ~new_P1_U3472;
  assign new_P1_U5008 = ~new_P1_R1162_U16 | ~new_P1_U3037;
  assign new_P1_U5009 = ~new_P1_U5008 | ~new_P1_U5007 | ~new_P1_U5006;
  assign new_P1_U5010 = ~new_P1_U3043 | ~new_P1_U5009;
  assign new_P1_U5011 = ~new_P1_R1105_U16 | ~new_P1_U3042;
  assign new_P1_U5012 = ~P1_REG3_REG_7_ | ~n1330;
  assign new_P1_U5013 = ~new_P1_U3040 | ~new_P1_U3472;
  assign new_P1_U5014 = ~new_P1_R1162_U16 | ~new_P1_U3038;
  assign new_P1_U5015 = ~P1_ADDR_REG_7_ | ~new_P1_U4889;
  assign new_P1_U5016 = ~new_P1_R1105_U72 | ~new_P1_U3041;
  assign new_P1_U5017 = ~new_P1_U3039 | ~new_P1_U3469;
  assign new_P1_U5018 = ~new_P1_R1162_U72 | ~new_P1_U3037;
  assign new_P1_U5019 = ~new_P1_U5018 | ~new_P1_U5017 | ~new_P1_U5016;
  assign new_P1_U5020 = ~new_P1_U3043 | ~new_P1_U5019;
  assign new_P1_U5021 = ~new_P1_R1105_U72 | ~new_P1_U3042;
  assign new_P1_U5022 = ~P1_REG3_REG_6_ | ~n1330;
  assign new_P1_U5023 = ~new_P1_U3040 | ~new_P1_U3469;
  assign new_P1_U5024 = ~new_P1_R1162_U72 | ~new_P1_U3038;
  assign new_P1_U5025 = ~P1_ADDR_REG_6_ | ~new_P1_U4889;
  assign new_P1_U5026 = ~new_P1_R1105_U15 | ~new_P1_U3041;
  assign new_P1_U5027 = ~new_P1_U3039 | ~new_P1_U3466;
  assign new_P1_U5028 = ~new_P1_R1162_U15 | ~new_P1_U3037;
  assign new_P1_U5029 = ~new_P1_U5028 | ~new_P1_U5027 | ~new_P1_U5026;
  assign new_P1_U5030 = ~new_P1_U3043 | ~new_P1_U5029;
  assign new_P1_U5031 = ~new_P1_R1105_U15 | ~new_P1_U3042;
  assign new_P1_U5032 = ~P1_REG3_REG_5_ | ~n1330;
  assign new_P1_U5033 = ~new_P1_U3040 | ~new_P1_U3466;
  assign new_P1_U5034 = ~new_P1_R1162_U15 | ~new_P1_U3038;
  assign new_P1_U5035 = ~P1_ADDR_REG_5_ | ~new_P1_U4889;
  assign new_P1_U5036 = ~new_P1_R1105_U73 | ~new_P1_U3041;
  assign new_P1_U5037 = ~new_P1_U3039 | ~new_P1_U3463;
  assign new_P1_U5038 = ~new_P1_R1162_U73 | ~new_P1_U3037;
  assign new_P1_U5039 = ~new_P1_U5038 | ~new_P1_U5037 | ~new_P1_U5036;
  assign new_P1_U5040 = ~new_P1_U3043 | ~new_P1_U5039;
  assign new_P1_U5041 = ~new_P1_R1105_U73 | ~new_P1_U3042;
  assign new_P1_U5042 = ~P1_REG3_REG_4_ | ~n1330;
  assign new_P1_U5043 = ~new_P1_U3040 | ~new_P1_U3463;
  assign new_P1_U5044 = ~new_P1_R1162_U73 | ~new_P1_U3038;
  assign new_P1_U5045 = ~P1_ADDR_REG_4_ | ~new_P1_U4889;
  assign new_P1_U5046 = ~new_P1_R1105_U74 | ~new_P1_U3041;
  assign new_P1_U5047 = ~new_P1_U3039 | ~new_P1_U3460;
  assign new_P1_U5048 = ~new_P1_R1162_U74 | ~new_P1_U3037;
  assign new_P1_U5049 = ~new_P1_U5048 | ~new_P1_U5047 | ~new_P1_U5046;
  assign new_P1_U5050 = ~new_P1_U3043 | ~new_P1_U5049;
  assign new_P1_U5051 = ~new_P1_R1105_U74 | ~new_P1_U3042;
  assign new_P1_U5052 = ~P1_REG3_REG_3_ | ~n1330;
  assign new_P1_U5053 = ~new_P1_U3040 | ~new_P1_U3460;
  assign new_P1_U5054 = ~new_P1_R1162_U74 | ~new_P1_U3038;
  assign new_P1_U5055 = ~P1_ADDR_REG_3_ | ~new_P1_U4889;
  assign new_P1_U5056 = ~new_P1_R1105_U14 | ~new_P1_U3041;
  assign new_P1_U5057 = ~new_P1_U3039 | ~new_P1_U3457;
  assign new_P1_U5058 = ~new_P1_R1162_U14 | ~new_P1_U3037;
  assign new_P1_U5059 = ~new_P1_U5058 | ~new_P1_U5057 | ~new_P1_U5056;
  assign new_P1_U5060 = ~new_P1_U3043 | ~new_P1_U5059;
  assign new_P1_U5061 = ~new_P1_R1105_U14 | ~new_P1_U3042;
  assign new_P1_U5062 = ~P1_REG3_REG_2_ | ~n1330;
  assign new_P1_U5063 = ~new_P1_U3040 | ~new_P1_U3457;
  assign new_P1_U5064 = ~new_P1_R1162_U14 | ~new_P1_U3038;
  assign new_P1_U5065 = ~P1_ADDR_REG_2_ | ~new_P1_U4889;
  assign new_P1_U5066 = ~new_P1_R1105_U68 | ~new_P1_U3041;
  assign new_P1_U5067 = ~new_P1_U3039 | ~new_P1_U3454;
  assign new_P1_U5068 = ~new_P1_R1162_U68 | ~new_P1_U3037;
  assign new_P1_U5069 = ~new_P1_U5068 | ~new_P1_U5067 | ~new_P1_U5066;
  assign new_P1_U5070 = ~new_P1_U3043 | ~new_P1_U5069;
  assign new_P1_U5071 = ~new_P1_R1105_U68 | ~new_P1_U3042;
  assign new_P1_U5072 = ~P1_REG3_REG_1_ | ~n1330;
  assign new_P1_U5073 = ~new_P1_U3040 | ~new_P1_U3454;
  assign new_P1_U5074 = ~new_P1_R1162_U68 | ~new_P1_U3038;
  assign new_P1_U5075 = ~P1_ADDR_REG_1_ | ~new_P1_U4889;
  assign new_P1_U5076 = ~new_P1_R1105_U69 | ~new_P1_U3041;
  assign new_P1_U5077 = ~new_P1_U3039 | ~new_P1_U3448;
  assign new_P1_U5078 = ~new_P1_R1162_U69 | ~new_P1_U3037;
  assign new_P1_U5079 = ~new_P1_U5078 | ~new_P1_U5077 | ~new_P1_U5076;
  assign new_P1_U5080 = ~new_P1_U3043 | ~new_P1_U5079;
  assign new_P1_U5081 = ~new_P1_R1105_U69 | ~new_P1_U3042;
  assign new_P1_U5082 = ~P1_REG3_REG_0_ | ~n1330;
  assign new_P1_U5083 = ~new_P1_U3040 | ~new_P1_U3448;
  assign new_P1_U5084 = ~new_P1_R1162_U69 | ~new_P1_U3038;
  assign new_P1_U5085 = ~P1_ADDR_REG_0_ | ~new_P1_U4889;
  assign new_P1_U5086 = ~new_P1_U3951;
  assign new_P1_U5087 = ~new_P1_LT_197_U13 | ~new_P1_U3954 | ~new_P1_U3987;
  assign new_P1_U5088 = ~new_P1_U5677 | ~new_P1_U3427;
  assign new_P1_U5089 = ~new_P1_U3851 | ~new_P1_U5088;
  assign new_P1_U5090 = ~new_P1_U3949 | ~new_P1_U3022 | ~new_P1_U3986;
  assign new_P1_U5091 = ~P1_B_REG | ~new_P1_U5089;
  assign new_P1_U5092 = ~new_P1_U3036 | ~new_P1_U3079;
  assign new_P1_U5093 = ~new_P1_U3034 | ~new_P1_U3073;
  assign new_P1_U5094 = ~new_P1_ADD_95_U73 | ~new_P1_U3430;
  assign new_P1_U5095 = ~new_P1_U5093 | ~new_P1_U5094 | ~new_P1_U5092;
  assign new_P1_U5096 = ~new_P1_U3362 | ~new_P1_U3364 | ~new_P1_U3361;
  assign new_P1_U5097 = ~new_P1_U3365 | ~new_P1_U3366 | ~new_P1_U3419;
  assign new_P1_U5098 = ~new_P1_U5684 | ~new_P1_U5097;
  assign new_P1_U5099 = ~new_P1_U5693 | ~new_P1_U5096;
  assign new_P1_U5100 = ~new_P1_U3868 | ~new_P1_U5099 | ~new_P1_U5098;
  assign new_P1_U5101 = ~new_P1_U5100 | ~new_P1_U3430;
  assign new_P1_U5102 = ~new_P1_U3432;
  assign new_P1_U5103 = ~new_P1_U3497 | ~new_P1_U5656;
  assign new_P1_U5104 = ~new_P1_ADD_95_U73 | ~new_P1_U5655;
  assign new_P1_U5105 = ~new_P1_U3994 | ~new_P1_U5095;
  assign new_P1_U5106 = ~new_P1_R1165_U104 | ~new_P1_U3027;
  assign new_P1_U5107 = ~P1_REG3_REG_15_ | ~n1330;
  assign new_P1_U5108 = ~new_P1_U3036 | ~new_P1_U3058;
  assign new_P1_U5109 = ~new_P1_U3034 | ~new_P1_U3053;
  assign new_P1_U5110 = ~new_P1_ADD_95_U62 | ~new_P1_U3430;
  assign new_P1_U5111 = ~new_P1_U5109 | ~new_P1_U5110 | ~new_P1_U5108;
  assign new_P1_U5112 = ~new_P1_U3422 | ~new_P1_U3430;
  assign new_P1_U5113 = ~new_P1_U5102 | ~new_P1_U5112;
  assign new_P1_U5114 = ~new_P1_U3972 | ~new_P1_U3422;
  assign new_P1_U5115 = ~new_P1_U3418 | ~new_P1_U5114;
  assign new_P1_U5116 = ~new_P1_U3045 | ~new_P1_U3976;
  assign new_P1_U5117 = ~new_P1_U3044 | ~new_P1_ADD_95_U62;
  assign new_P1_U5118 = ~new_P1_U3994 | ~new_P1_U5111;
  assign new_P1_U5119 = ~new_P1_R1165_U13 | ~new_P1_U3027;
  assign new_P1_U5120 = ~P1_REG3_REG_26_ | ~n1330;
  assign new_P1_U5121 = ~new_P1_U3036 | ~new_P1_U3067;
  assign new_P1_U5122 = ~new_P1_U3034 | ~new_P1_U3070;
  assign new_P1_U5123 = ~new_P1_ADD_95_U57 | ~new_P1_U3430;
  assign new_P1_U5124 = ~new_P1_U5123 | ~new_P1_U5122 | ~new_P1_U5121;
  assign new_P1_U5125 = ~new_P1_U3470 | ~new_P1_U5656;
  assign new_P1_U5126 = ~new_P1_ADD_95_U57 | ~new_P1_U5655;
  assign new_P1_U5127 = ~new_P1_U3994 | ~new_P1_U5124;
  assign new_P1_U5128 = ~new_P1_R1165_U89 | ~new_P1_U3027;
  assign new_P1_U5129 = ~P1_REG3_REG_6_ | ~n1330;
  assign new_P1_U5130 = ~new_P1_U3036 | ~new_P1_U3069;
  assign new_P1_U5131 = ~new_P1_U3034 | ~new_P1_U3081;
  assign new_P1_U5132 = ~new_P1_ADD_95_U70 | ~new_P1_U3430;
  assign new_P1_U5133 = ~new_P1_U5131 | ~new_P1_U5132 | ~new_P1_U5130;
  assign new_P1_U5134 = ~new_P1_U3506 | ~new_P1_U5656;
  assign new_P1_U5135 = ~new_P1_ADD_95_U70 | ~new_P1_U5655;
  assign new_P1_U5136 = ~new_P1_U3994 | ~new_P1_U5133;
  assign new_P1_U5137 = ~new_P1_R1165_U102 | ~new_P1_U3027;
  assign new_P1_U5138 = ~P1_REG3_REG_18_ | ~n1330;
  assign new_P1_U5139 = ~new_P1_U3036 | ~new_P1_U3078;
  assign new_P1_U5140 = ~new_P1_U3034 | ~new_P1_U3064;
  assign new_P1_U5141 = ~P1_REG3_REG_2_ | ~new_P1_U3430;
  assign new_P1_U5142 = ~new_P1_U5141 | ~new_P1_U5140 | ~new_P1_U5139;
  assign new_P1_U5143 = ~new_P1_U3458 | ~new_P1_U5656;
  assign new_P1_U5144 = ~P1_REG3_REG_2_ | ~new_P1_U5655;
  assign new_P1_U5145 = ~new_P1_U3994 | ~new_P1_U5142;
  assign new_P1_U5146 = ~new_P1_R1165_U92 | ~new_P1_U3027;
  assign new_P1_U5147 = ~P1_REG3_REG_2_ | ~n1330;
  assign new_P1_U5148 = ~new_P1_U3036 | ~new_P1_U3062;
  assign new_P1_U5149 = ~new_P1_U3034 | ~new_P1_U3072;
  assign new_P1_U5150 = ~new_P1_ADD_95_U77 | ~new_P1_U3430;
  assign new_P1_U5151 = ~new_P1_U5150 | ~new_P1_U5149 | ~new_P1_U5148;
  assign new_P1_U5152 = ~new_P1_U3485 | ~new_P1_U5656;
  assign new_P1_U5153 = ~new_P1_ADD_95_U77 | ~new_P1_U5655;
  assign new_P1_U5154 = ~new_P1_U3994 | ~new_P1_U5151;
  assign new_P1_U5155 = ~new_P1_R1165_U107 | ~new_P1_U3027;
  assign new_P1_U5156 = ~P1_REG3_REG_11_ | ~n1330;
  assign new_P1_U5157 = ~new_P1_U3036 | ~new_P1_U3075;
  assign new_P1_U5158 = ~new_P1_U3034 | ~new_P1_U3066;
  assign new_P1_U5159 = ~new_P1_ADD_95_U66 | ~new_P1_U3430;
  assign new_P1_U5160 = ~new_P1_U5158 | ~new_P1_U5159 | ~new_P1_U5157;
  assign new_P1_U5161 = ~new_P1_U3045 | ~new_P1_U3980;
  assign new_P1_U5162 = ~new_P1_U3044 | ~new_P1_ADD_95_U66;
  assign new_P1_U5163 = ~new_P1_U3994 | ~new_P1_U5160;
  assign new_P1_U5164 = ~new_P1_R1165_U98 | ~new_P1_U3027;
  assign new_P1_U5165 = ~P1_REG3_REG_22_ | ~n1330;
  assign new_P1_U5166 = ~new_P1_U3036 | ~new_P1_U3072;
  assign new_P1_U5167 = ~new_P1_U3034 | ~new_P1_U3079;
  assign new_P1_U5168 = ~new_P1_ADD_95_U75 | ~new_P1_U3430;
  assign new_P1_U5169 = ~new_P1_U5167 | ~new_P1_U5168 | ~new_P1_U5166;
  assign new_P1_U5170 = ~new_P1_U3491 | ~new_P1_U5656;
  assign new_P1_U5171 = ~new_P1_ADD_95_U75 | ~new_P1_U5655;
  assign new_P1_U5172 = ~new_P1_U3994 | ~new_P1_U5169;
  assign new_P1_U5173 = ~new_P1_R1165_U10 | ~new_P1_U3027;
  assign new_P1_U5174 = ~P1_REG3_REG_13_ | ~n1330;
  assign new_P1_U5175 = ~new_P1_U3036 | ~new_P1_U3081;
  assign new_P1_U5176 = ~new_P1_U3034 | ~new_P1_U3075;
  assign new_P1_U5177 = ~new_P1_ADD_95_U68 | ~new_P1_U3430;
  assign new_P1_U5178 = ~new_P1_U5176 | ~new_P1_U5177 | ~new_P1_U5175;
  assign new_P1_U5179 = ~new_P1_U3045 | ~new_P1_U3982;
  assign new_P1_U5180 = ~new_P1_U3044 | ~new_P1_ADD_95_U68;
  assign new_P1_U5181 = ~new_P1_U3994 | ~new_P1_U5178;
  assign new_P1_U5182 = ~new_P1_R1165_U99 | ~new_P1_U3027;
  assign new_P1_U5183 = ~P1_REG3_REG_20_ | ~n1330;
  assign new_P1_U5184 = ~new_P1_U3431 | ~new_P1_U3429;
  assign new_P1_U5185 = ~new_P1_U5184 | ~new_P1_U3430;
  assign new_P1_U5186 = ~new_P1_U3995 | ~new_P1_U5185;
  assign new_P1_U5187 = ~new_P1_U3873 | ~new_P1_U3034;
  assign new_P1_U5188 = ~new_P1_U3450 | ~new_P1_U5656;
  assign new_P1_U5189 = ~P1_REG3_REG_0_ | ~new_P1_U5186;
  assign new_P1_U5190 = ~new_P1_R1165_U86 | ~new_P1_U3027;
  assign new_P1_U5191 = ~P1_REG3_REG_0_ | ~n1330;
  assign new_P1_U5192 = ~new_P1_U3036 | ~new_P1_U3084;
  assign new_P1_U5193 = ~new_P1_U3034 | ~new_P1_U3062;
  assign new_P1_U5194 = ~new_P1_ADD_95_U54 | ~new_P1_U3430;
  assign new_P1_U5195 = ~new_P1_U5194 | ~new_P1_U5193 | ~new_P1_U5192;
  assign new_P1_U5196 = ~new_P1_U3479 | ~new_P1_U5656;
  assign new_P1_U5197 = ~new_P1_ADD_95_U54 | ~new_P1_U5655;
  assign new_P1_U5198 = ~new_P1_U3994 | ~new_P1_U5195;
  assign new_P1_U5199 = ~new_P1_R1165_U87 | ~new_P1_U3027;
  assign new_P1_U5200 = ~P1_REG3_REG_9_ | ~n1330;
  assign new_P1_U5201 = ~new_P1_U3036 | ~new_P1_U3064;
  assign new_P1_U5202 = ~new_P1_U3034 | ~new_P1_U3067;
  assign new_P1_U5203 = ~new_P1_ADD_95_U59 | ~new_P1_U3430;
  assign new_P1_U5204 = ~new_P1_U5203 | ~new_P1_U5202 | ~new_P1_U5201;
  assign new_P1_U5205 = ~new_P1_U3464 | ~new_P1_U5656;
  assign new_P1_U5206 = ~new_P1_ADD_95_U59 | ~new_P1_U5655;
  assign new_P1_U5207 = ~new_P1_U3994 | ~new_P1_U5204;
  assign new_P1_U5208 = ~new_P1_R1165_U91 | ~new_P1_U3027;
  assign new_P1_U5209 = ~P1_REG3_REG_4_ | ~n1330;
  assign new_P1_U5210 = ~new_P1_U3036 | ~new_P1_U3066;
  assign new_P1_U5211 = ~new_P1_U3034 | ~new_P1_U3058;
  assign new_P1_U5212 = ~new_P1_ADD_95_U64 | ~new_P1_U3430;
  assign new_P1_U5213 = ~new_P1_U5211 | ~new_P1_U5212 | ~new_P1_U5210;
  assign new_P1_U5214 = ~new_P1_U3045 | ~new_P1_U3978;
  assign new_P1_U5215 = ~new_P1_U3044 | ~new_P1_ADD_95_U64;
  assign new_P1_U5216 = ~new_P1_U3994 | ~new_P1_U5213;
  assign new_P1_U5217 = ~new_P1_R1165_U96 | ~new_P1_U3027;
  assign new_P1_U5218 = ~P1_REG3_REG_24_ | ~n1330;
  assign new_P1_U5219 = ~new_P1_U3036 | ~new_P1_U3073;
  assign new_P1_U5220 = ~new_P1_U3034 | ~new_P1_U3082;
  assign new_P1_U5221 = ~new_P1_ADD_95_U71 | ~new_P1_U3430;
  assign new_P1_U5222 = ~new_P1_U5220 | ~new_P1_U5221 | ~new_P1_U5219;
  assign new_P1_U5223 = ~new_P1_U3503 | ~new_P1_U5656;
  assign new_P1_U5224 = ~new_P1_ADD_95_U71 | ~new_P1_U5655;
  assign new_P1_U5225 = ~new_P1_U3994 | ~new_P1_U5222;
  assign new_P1_U5226 = ~new_P1_R1165_U11 | ~new_P1_U3027;
  assign new_P1_U5227 = ~P1_REG3_REG_17_ | ~n1330;
  assign new_P1_U5228 = ~new_P1_U3036 | ~new_P1_U3060;
  assign new_P1_U5229 = ~new_P1_U3034 | ~new_P1_U3071;
  assign new_P1_U5230 = ~new_P1_ADD_95_U58 | ~new_P1_U3430;
  assign new_P1_U5231 = ~new_P1_U5230 | ~new_P1_U5229 | ~new_P1_U5228;
  assign new_P1_U5232 = ~new_P1_U3467 | ~new_P1_U5656;
  assign new_P1_U5233 = ~new_P1_ADD_95_U58 | ~new_P1_U5655;
  assign new_P1_U5234 = ~new_P1_U3994 | ~new_P1_U5231;
  assign new_P1_U5235 = ~new_P1_R1165_U90 | ~new_P1_U3027;
  assign new_P1_U5236 = ~P1_REG3_REG_5_ | ~n1330;
  assign new_P1_U5237 = ~new_P1_U3036 | ~new_P1_U3074;
  assign new_P1_U5238 = ~new_P1_U3034 | ~new_P1_U3069;
  assign new_P1_U5239 = ~new_P1_ADD_95_U72 | ~new_P1_U3430;
  assign new_P1_U5240 = ~new_P1_U5238 | ~new_P1_U5239 | ~new_P1_U5237;
  assign new_P1_U5241 = ~new_P1_U3500 | ~new_P1_U5656;
  assign new_P1_U5242 = ~new_P1_ADD_95_U72 | ~new_P1_U5655;
  assign new_P1_U5243 = ~new_P1_U3994 | ~new_P1_U5240;
  assign new_P1_U5244 = ~new_P1_R1165_U103 | ~new_P1_U3027;
  assign new_P1_U5245 = ~P1_REG3_REG_16_ | ~n1330;
  assign new_P1_U5246 = ~new_P1_U3036 | ~new_P1_U3065;
  assign new_P1_U5247 = ~new_P1_U3034 | ~new_P1_U3057;
  assign new_P1_U5248 = ~new_P1_ADD_95_U63 | ~new_P1_U3430;
  assign new_P1_U5249 = ~new_P1_U5247 | ~new_P1_U5248 | ~new_P1_U5246;
  assign new_P1_U5250 = ~new_P1_U3045 | ~new_P1_U3977;
  assign new_P1_U5251 = ~new_P1_U3044 | ~new_P1_ADD_95_U63;
  assign new_P1_U5252 = ~new_P1_U3994 | ~new_P1_U5249;
  assign new_P1_U5253 = ~new_P1_R1165_U95 | ~new_P1_U3027;
  assign new_P1_U5254 = ~P1_REG3_REG_25_ | ~n1330;
  assign new_P1_U5255 = ~new_P1_U3036 | ~new_P1_U3063;
  assign new_P1_U5256 = ~new_P1_U3034 | ~new_P1_U3080;
  assign new_P1_U5257 = ~new_P1_ADD_95_U76 | ~new_P1_U3430;
  assign new_P1_U5258 = ~new_P1_U5256 | ~new_P1_U5257 | ~new_P1_U5255;
  assign new_P1_U5259 = ~new_P1_U3488 | ~new_P1_U5656;
  assign new_P1_U5260 = ~new_P1_ADD_95_U76 | ~new_P1_U5655;
  assign new_P1_U5261 = ~new_P1_U3994 | ~new_P1_U5258;
  assign new_P1_U5262 = ~new_P1_R1165_U106 | ~new_P1_U3027;
  assign new_P1_U5263 = ~P1_REG3_REG_12_ | ~n1330;
  assign new_P1_U5264 = ~new_P1_U3036 | ~new_P1_U3076;
  assign new_P1_U5265 = ~new_P1_U3034 | ~new_P1_U3061;
  assign new_P1_U5266 = ~new_P1_ADD_95_U67 | ~new_P1_U3430;
  assign new_P1_U5267 = ~new_P1_U5265 | ~new_P1_U5266 | ~new_P1_U5264;
  assign new_P1_U5268 = ~new_P1_U3045 | ~new_P1_U3981;
  assign new_P1_U5269 = ~new_P1_U3044 | ~new_P1_ADD_95_U67;
  assign new_P1_U5270 = ~new_P1_U3994 | ~new_P1_U5267;
  assign new_P1_U5271 = ~new_P1_R1165_U12 | ~new_P1_U3027;
  assign new_P1_U5272 = ~P1_REG3_REG_21_ | ~n1330;
  assign new_P1_U5273 = ~new_P1_U3036 | ~new_P1_U3077;
  assign new_P1_U5274 = ~new_P1_U3034 | ~new_P1_U3068;
  assign new_P1_U5275 = ~P1_REG3_REG_1_ | ~new_P1_U3430;
  assign new_P1_U5276 = ~new_P1_U5275 | ~new_P1_U5274 | ~new_P1_U5273;
  assign new_P1_U5277 = ~new_P1_U3455 | ~new_P1_U5656;
  assign new_P1_U5278 = ~P1_REG3_REG_1_ | ~new_P1_U5655;
  assign new_P1_U5279 = ~new_P1_U3994 | ~new_P1_U5276;
  assign new_P1_U5280 = ~new_P1_R1165_U100 | ~new_P1_U3027;
  assign new_P1_U5281 = ~P1_REG3_REG_1_ | ~n1330;
  assign new_P1_U5282 = ~new_P1_U3036 | ~new_P1_U3070;
  assign new_P1_U5283 = ~new_P1_U3034 | ~new_P1_U3083;
  assign new_P1_U5284 = ~new_P1_ADD_95_U55 | ~new_P1_U3430;
  assign new_P1_U5285 = ~new_P1_U5284 | ~new_P1_U5283 | ~new_P1_U5282;
  assign new_P1_U5286 = ~new_P1_U3476 | ~new_P1_U5656;
  assign new_P1_U5287 = ~new_P1_ADD_95_U55 | ~new_P1_U5655;
  assign new_P1_U5288 = ~new_P1_U3994 | ~new_P1_U5285;
  assign new_P1_U5289 = ~new_P1_R1165_U88 | ~new_P1_U3027;
  assign new_P1_U5290 = ~P1_REG3_REG_8_ | ~n1330;
  assign new_P1_U5291 = ~new_P1_U3036 | ~new_P1_U3053;
  assign new_P1_U5292 = ~new_P1_U3034 | ~new_P1_U3055;
  assign new_P1_U5293 = ~new_P1_ADD_95_U60 | ~new_P1_U3430;
  assign new_P1_U5294 = ~new_P1_U5293 | ~new_P1_U5292 | ~new_P1_U5291;
  assign new_P1_U5295 = ~new_P1_U3045 | ~new_P1_U3974;
  assign new_P1_U5296 = ~new_P1_U3044 | ~new_P1_ADD_95_U60;
  assign new_P1_U5297 = ~new_P1_U3994 | ~new_P1_U5294;
  assign new_P1_U5298 = ~new_P1_R1165_U93 | ~new_P1_U3027;
  assign new_P1_U5299 = ~P1_REG3_REG_28_ | ~n1330;
  assign new_P1_U5300 = ~new_P1_U3036 | ~new_P1_U3082;
  assign new_P1_U5301 = ~new_P1_U3034 | ~new_P1_U3076;
  assign new_P1_U5302 = ~new_P1_ADD_95_U69 | ~new_P1_U3430;
  assign new_P1_U5303 = ~new_P1_U5301 | ~new_P1_U5302 | ~new_P1_U5300;
  assign new_P1_U5304 = ~new_P1_U3508 | ~new_P1_U5656;
  assign new_P1_U5305 = ~new_P1_ADD_95_U69 | ~new_P1_U5655;
  assign new_P1_U5306 = ~new_P1_U3994 | ~new_P1_U5303;
  assign new_P1_U5307 = ~new_P1_R1165_U101 | ~new_P1_U3027;
  assign new_P1_U5308 = ~P1_REG3_REG_19_ | ~n1330;
  assign new_P1_U5309 = ~new_P1_U3036 | ~new_P1_U3068;
  assign new_P1_U5310 = ~new_P1_U3034 | ~new_P1_U3060;
  assign new_P1_U5311 = ~new_P1_ADD_95_U4 | ~new_P1_U3430;
  assign new_P1_U5312 = ~new_P1_U5311 | ~new_P1_U5310 | ~new_P1_U5309;
  assign new_P1_U5313 = ~new_P1_U3461 | ~new_P1_U5656;
  assign new_P1_U5314 = ~new_P1_ADD_95_U4 | ~new_P1_U5655;
  assign new_P1_U5315 = ~new_P1_U3994 | ~new_P1_U5312;
  assign new_P1_U5316 = ~new_P1_R1165_U14 | ~new_P1_U3027;
  assign new_P1_U5317 = ~P1_REG3_REG_3_ | ~n1330;
  assign new_P1_U5318 = ~new_P1_U3036 | ~new_P1_U3083;
  assign new_P1_U5319 = ~new_P1_U3034 | ~new_P1_U3063;
  assign new_P1_U5320 = ~new_P1_ADD_95_U78 | ~new_P1_U3430;
  assign new_P1_U5321 = ~new_P1_U5320 | ~new_P1_U5319 | ~new_P1_U5318;
  assign new_P1_U5322 = ~new_P1_U3482 | ~new_P1_U5656;
  assign new_P1_U5323 = ~new_P1_ADD_95_U78 | ~new_P1_U5655;
  assign new_P1_U5324 = ~new_P1_U3994 | ~new_P1_U5321;
  assign new_P1_U5325 = ~new_P1_R1165_U108 | ~new_P1_U3027;
  assign new_P1_U5326 = ~P1_REG3_REG_10_ | ~n1330;
  assign new_P1_U5327 = ~new_P1_U3036 | ~new_P1_U3061;
  assign new_P1_U5328 = ~new_P1_U3034 | ~new_P1_U3065;
  assign new_P1_U5329 = ~new_P1_ADD_95_U65 | ~new_P1_U3430;
  assign new_P1_U5330 = ~new_P1_U5328 | ~new_P1_U5329 | ~new_P1_U5327;
  assign new_P1_U5331 = ~new_P1_U3045 | ~new_P1_U3979;
  assign new_P1_U5332 = ~new_P1_U3044 | ~new_P1_ADD_95_U65;
  assign new_P1_U5333 = ~new_P1_U3994 | ~new_P1_U5330;
  assign new_P1_U5334 = ~new_P1_R1165_U97 | ~new_P1_U3027;
  assign new_P1_U5335 = ~P1_REG3_REG_23_ | ~n1330;
  assign new_P1_U5336 = ~new_P1_U3036 | ~new_P1_U3080;
  assign new_P1_U5337 = ~new_P1_U3034 | ~new_P1_U3074;
  assign new_P1_U5338 = ~new_P1_ADD_95_U74 | ~new_P1_U3430;
  assign new_P1_U5339 = ~new_P1_U5337 | ~new_P1_U5338 | ~new_P1_U5336;
  assign new_P1_U5340 = ~new_P1_U3494 | ~new_P1_U5656;
  assign new_P1_U5341 = ~new_P1_ADD_95_U74 | ~new_P1_U5655;
  assign new_P1_U5342 = ~new_P1_U3994 | ~new_P1_U5339;
  assign new_P1_U5343 = ~new_P1_R1165_U105 | ~new_P1_U3027;
  assign new_P1_U5344 = ~P1_REG3_REG_14_ | ~n1330;
  assign new_P1_U5345 = ~new_P1_U3036 | ~new_P1_U3057;
  assign new_P1_U5346 = ~new_P1_U3034 | ~new_P1_U3054;
  assign new_P1_U5347 = ~new_P1_ADD_95_U61 | ~new_P1_U3430;
  assign new_P1_U5348 = ~new_P1_U5346 | ~new_P1_U5347 | ~new_P1_U5345;
  assign new_P1_U5349 = ~new_P1_U3045 | ~new_P1_U3975;
  assign new_P1_U5350 = ~new_P1_U3044 | ~new_P1_ADD_95_U61;
  assign new_P1_U5351 = ~new_P1_U3994 | ~new_P1_U5348;
  assign new_P1_U5352 = ~new_P1_R1165_U94 | ~new_P1_U3027;
  assign new_P1_U5353 = ~P1_REG3_REG_27_ | ~n1330;
  assign new_P1_U5354 = ~new_P1_U3036 | ~new_P1_U3071;
  assign new_P1_U5355 = ~new_P1_U3034 | ~new_P1_U3084;
  assign new_P1_U5356 = ~new_P1_ADD_95_U56 | ~new_P1_U3430;
  assign new_P1_U5357 = ~new_P1_U5356 | ~new_P1_U5355 | ~new_P1_U5354;
  assign new_P1_U5358 = ~new_P1_U3473 | ~new_P1_U5656;
  assign new_P1_U5359 = ~new_P1_ADD_95_U56 | ~new_P1_U5655;
  assign new_P1_U5360 = ~new_P1_U3994 | ~new_P1_U5357;
  assign new_P1_U5361 = ~new_P1_R1165_U15 | ~new_P1_U3027;
  assign new_P1_U5362 = ~P1_REG3_REG_7_ | ~n1330;
  assign new_P1_U5363 = ~new_P1_U3449 | ~new_P1_U3375;
  assign new_P1_U5364 = ~new_P1_U3446 | ~new_P1_U5363;
  assign new_P1_U5365 = ~new_P1_R1165_U86 | ~new_P1_U5702 | ~new_P1_U3446;
  assign new_P1_U5366 = ~new_P1_U3447 | ~new_P1_U3441;
  assign new_P1_U5367 = ~new_P1_U3877 | ~new_P1_U3970;
  assign new_P1_U5368 = ~new_P1_U3370 | ~new_P1_U3419;
  assign new_P1_U5369 = ~new_P1_U3365 | ~new_P1_U3368 | ~new_P1_U3363;
  assign new_P1_U5370 = ~new_P1_U4000 | ~new_P1_U3421;
  assign new_P1_U5371 = ~new_P1_U5369 | ~new_P1_U3421;
  assign new_P1_U5372 = ~new_P1_U3434;
  assign new_P1_U5373 = ~new_P1_U5372 | ~new_P1_U3970;
  assign new_P1_U5374 = ~new_P1_U3479 | ~new_P1_U5373;
  assign new_P1_U5375 = ~new_P1_U3021 | ~new_P1_U3083;
  assign new_P1_U5376 = ~new_P1_U3476 | ~new_P1_U5373;
  assign new_P1_U5377 = ~new_P1_U3021 | ~new_P1_U3084;
  assign new_P1_U5378 = ~new_P1_U3473 | ~new_P1_U5373;
  assign new_P1_U5379 = ~new_P1_U3021 | ~new_P1_U3070;
  assign new_P1_U5380 = ~new_P1_U3470 | ~new_P1_U5373;
  assign new_P1_U5381 = ~new_P1_U3021 | ~new_P1_U3071;
  assign new_P1_U5382 = ~new_P1_U3467 | ~new_P1_U5373;
  assign new_P1_U5383 = ~new_P1_U3021 | ~new_P1_U3067;
  assign new_P1_U5384 = ~new_P1_U3464 | ~new_P1_U5373;
  assign new_P1_U5385 = ~new_P1_U3021 | ~new_P1_U3060;
  assign new_P1_U5386 = ~new_P1_U3461 | ~new_P1_U5373;
  assign new_P1_U5387 = ~new_P1_U3021 | ~new_P1_U3064;
  assign new_P1_U5388 = ~new_P1_U3974 | ~new_P1_U5373;
  assign new_P1_U5389 = ~new_P1_U3021 | ~new_P1_U3054;
  assign new_P1_U5390 = ~new_P1_U3975 | ~new_P1_U5373;
  assign new_P1_U5391 = ~new_P1_U3021 | ~new_P1_U3053;
  assign new_P1_U5392 = ~new_P1_U3976 | ~new_P1_U5373;
  assign new_P1_U5393 = ~new_P1_U3021 | ~new_P1_U3057;
  assign new_P1_U5394 = ~new_P1_U3977 | ~new_P1_U5373;
  assign new_P1_U5395 = ~new_P1_U3021 | ~new_P1_U3058;
  assign new_P1_U5396 = ~new_P1_U3978 | ~new_P1_U5373;
  assign new_P1_U5397 = ~new_P1_U3021 | ~new_P1_U3065;
  assign new_P1_U5398 = ~new_P1_U3979 | ~new_P1_U5373;
  assign new_P1_U5399 = ~new_P1_U3021 | ~new_P1_U3066;
  assign new_P1_U5400 = ~new_P1_U3980 | ~new_P1_U5373;
  assign new_P1_U5401 = ~new_P1_U3021 | ~new_P1_U3061;
  assign new_P1_U5402 = ~new_P1_U3981 | ~new_P1_U5373;
  assign new_P1_U5403 = ~new_P1_U3021 | ~new_P1_U3075;
  assign new_P1_U5404 = ~new_P1_U3982 | ~new_P1_U5373;
  assign new_P1_U5405 = ~new_P1_U3021 | ~new_P1_U3076;
  assign new_P1_U5406 = ~new_P1_U3458 | ~new_P1_U5373;
  assign new_P1_U5407 = ~new_P1_U3021 | ~new_P1_U3068;
  assign new_P1_U5408 = ~new_P1_U3508 | ~new_P1_U5373;
  assign new_P1_U5409 = ~new_P1_U3021 | ~new_P1_U3081;
  assign new_P1_U5410 = ~new_P1_U3506 | ~new_P1_U5373;
  assign new_P1_U5411 = ~new_P1_U3021 | ~new_P1_U3082;
  assign new_P1_U5412 = ~new_P1_U3503 | ~new_P1_U5373;
  assign new_P1_U5413 = ~new_P1_U3021 | ~new_P1_U3069;
  assign new_P1_U5414 = ~new_P1_U3500 | ~new_P1_U5373;
  assign new_P1_U5415 = ~new_P1_U3021 | ~new_P1_U3073;
  assign new_P1_U5416 = ~new_P1_U3497 | ~new_P1_U5373;
  assign new_P1_U5417 = ~new_P1_U3021 | ~new_P1_U3074;
  assign new_P1_U5418 = ~new_P1_U3494 | ~new_P1_U5373;
  assign new_P1_U5419 = ~new_P1_U3021 | ~new_P1_U3079;
  assign new_P1_U5420 = ~new_P1_U3491 | ~new_P1_U5373;
  assign new_P1_U5421 = ~new_P1_U3021 | ~new_P1_U3080;
  assign new_P1_U5422 = ~new_P1_U3488 | ~new_P1_U5373;
  assign new_P1_U5423 = ~new_P1_U3021 | ~new_P1_U3072;
  assign new_P1_U5424 = ~new_P1_U3485 | ~new_P1_U5373;
  assign new_P1_U5425 = ~new_P1_U3021 | ~new_P1_U3063;
  assign new_P1_U5426 = ~new_P1_U3482 | ~new_P1_U5373;
  assign new_P1_U5427 = ~new_P1_U3021 | ~new_P1_U3062;
  assign new_P1_U5428 = ~new_P1_U3455 | ~new_P1_U5373;
  assign new_P1_U5429 = ~new_P1_U3021 | ~new_P1_U3078;
  assign new_P1_U5430 = ~new_P1_U3450 | ~new_P1_U5373;
  assign new_P1_U5431 = ~new_P1_U3021 | ~new_P1_U3077;
  assign new_P1_U5432 = ~new_P1_U4102 | ~P1_REG1_REG_0_;
  assign new_P1_U5433 = ~new_P1_U3021 | ~new_P1_U3479;
  assign new_P1_U5434 = ~new_P1_U3434 | ~new_P1_U3083;
  assign new_P1_U5435 = ~new_P1_U3021 | ~new_P1_U3476;
  assign new_P1_U5436 = ~new_P1_U3434 | ~new_P1_U3084;
  assign new_P1_U5437 = ~new_P1_U3021 | ~new_P1_U3473;
  assign new_P1_U5438 = ~new_P1_U3434 | ~new_P1_U3070;
  assign new_P1_U5439 = ~new_P1_U3021 | ~new_P1_U3470;
  assign new_P1_U5440 = ~new_P1_U3434 | ~new_P1_U3071;
  assign new_P1_U5441 = ~new_P1_U3021 | ~new_P1_U3467;
  assign new_P1_U5442 = ~new_P1_U3434 | ~new_P1_U3067;
  assign new_P1_U5443 = ~new_P1_U3021 | ~new_P1_U3464;
  assign new_P1_U5444 = ~new_P1_U3434 | ~new_P1_U3060;
  assign new_P1_U5445 = ~new_P1_U3021 | ~new_P1_U3461;
  assign new_P1_U5446 = ~new_P1_U3434 | ~new_P1_U3064;
  assign new_P1_U5447 = ~new_P1_U3021 | ~new_P1_U3974;
  assign new_P1_U5448 = ~new_P1_U3434 | ~new_P1_U3054;
  assign new_P1_U5449 = ~new_P1_U3021 | ~new_P1_U3975;
  assign new_P1_U5450 = ~new_P1_U3434 | ~new_P1_U3053;
  assign new_P1_U5451 = ~new_P1_U3021 | ~new_P1_U3976;
  assign new_P1_U5452 = ~new_P1_U3434 | ~new_P1_U3057;
  assign new_P1_U5453 = ~new_P1_U3021 | ~new_P1_U3977;
  assign new_P1_U5454 = ~new_P1_U3434 | ~new_P1_U3058;
  assign new_P1_U5455 = ~new_P1_U3021 | ~new_P1_U3978;
  assign new_P1_U5456 = ~new_P1_U3434 | ~new_P1_U3065;
  assign new_P1_U5457 = ~new_P1_U3021 | ~new_P1_U3979;
  assign new_P1_U5458 = ~new_P1_U3434 | ~new_P1_U3066;
  assign new_P1_U5459 = ~new_P1_U3021 | ~new_P1_U3980;
  assign new_P1_U5460 = ~new_P1_U3434 | ~new_P1_U3061;
  assign new_P1_U5461 = ~new_P1_U3021 | ~new_P1_U3981;
  assign new_P1_U5462 = ~new_P1_U3434 | ~new_P1_U3075;
  assign new_P1_U5463 = ~new_P1_U3021 | ~new_P1_U3982;
  assign new_P1_U5464 = ~new_P1_U3434 | ~new_P1_U3076;
  assign new_P1_U5465 = ~new_P1_U3021 | ~new_P1_U3458;
  assign new_P1_U5466 = ~new_P1_U3434 | ~new_P1_U3068;
  assign new_P1_U5467 = ~new_P1_U3021 | ~new_P1_U3508;
  assign new_P1_U5468 = ~new_P1_U3434 | ~new_P1_U3081;
  assign new_P1_U5469 = ~new_P1_U3021 | ~new_P1_U3506;
  assign new_P1_U5470 = ~new_P1_U3434 | ~new_P1_U3082;
  assign new_P1_U5471 = ~new_P1_U3021 | ~new_P1_U3503;
  assign new_P1_U5472 = ~new_P1_U3434 | ~new_P1_U3069;
  assign new_P1_U5473 = ~new_P1_U3021 | ~new_P1_U3500;
  assign new_P1_U5474 = ~new_P1_U3434 | ~new_P1_U3073;
  assign new_P1_U5475 = ~new_P1_U3021 | ~new_P1_U3497;
  assign new_P1_U5476 = ~new_P1_U3434 | ~new_P1_U3074;
  assign new_P1_U5477 = ~new_P1_U3021 | ~new_P1_U3494;
  assign new_P1_U5478 = ~new_P1_U3434 | ~new_P1_U3079;
  assign new_P1_U5479 = ~new_P1_U3021 | ~new_P1_U3491;
  assign new_P1_U5480 = ~new_P1_U3434 | ~new_P1_U3080;
  assign new_P1_U5481 = ~new_P1_U3021 | ~new_P1_U3488;
  assign new_P1_U5482 = ~new_P1_U3434 | ~new_P1_U3072;
  assign new_P1_U5483 = ~new_P1_U3021 | ~new_P1_U3485;
  assign new_P1_U5484 = ~new_P1_U3434 | ~new_P1_U3063;
  assign new_P1_U5485 = ~new_P1_U3021 | ~new_P1_U3482;
  assign new_P1_U5486 = ~new_P1_U3434 | ~new_P1_U3062;
  assign new_P1_U5487 = ~new_P1_U3021 | ~new_P1_U3455;
  assign new_P1_U5488 = ~new_P1_U3434 | ~new_P1_U3078;
  assign new_P1_U5489 = ~new_P1_U3021 | ~new_P1_U3450;
  assign new_P1_U5490 = ~new_P1_U3434 | ~new_P1_U3077;
  assign new_P1_U5491 = ~new_P1_U4102 | ~new_P1_U3448;
  assign new_P1_U5492 = ~new_P1_U3426 | ~new_P1_U3428;
  assign new_P1_U5493 = ~new_P1_U3953 | ~new_P1_U3479;
  assign new_P1_U5494 = ~new_P1_U3586 | ~new_P1_U5492;
  assign new_P1_U5495 = ~new_P1_U3953 | ~new_P1_U3476;
  assign new_P1_U5496 = ~new_P1_U3587 | ~new_P1_U5492;
  assign new_P1_U5497 = ~new_P1_U3953 | ~new_P1_U3473;
  assign new_P1_U5498 = ~new_P1_U3588 | ~new_P1_U5492;
  assign new_P1_U5499 = ~new_P1_U3953 | ~new_P1_U3470;
  assign new_P1_U5500 = ~new_P1_U3589 | ~new_P1_U5492;
  assign new_P1_U5501 = ~new_P1_U3953 | ~new_P1_U3467;
  assign new_P1_U5502 = ~new_P1_U3590 | ~new_P1_U5492;
  assign new_P1_U5503 = ~new_P1_U3953 | ~new_P1_U3464;
  assign new_P1_U5504 = ~new_P1_U3591 | ~new_P1_U5492;
  assign new_P1_U5505 = ~new_P1_U3593 | ~new_P1_U5492;
  assign new_P1_U5506 = ~new_P1_U3983 | ~new_P1_U3953;
  assign new_P1_U5507 = ~new_P1_U3594 | ~new_P1_U5492;
  assign new_P1_U5508 = ~new_P1_U3984 | ~new_P1_U3953;
  assign new_P1_U5509 = ~new_P1_U3953 | ~new_P1_U3461;
  assign new_P1_U5510 = ~new_P1_U3592 | ~new_P1_U5492;
  assign new_P1_U5511 = ~new_P1_U3596 | ~new_P1_U5492;
  assign new_P1_U5512 = ~new_P1_U3985 | ~new_P1_U3953;
  assign new_P1_U5513 = ~new_P1_U3597 | ~new_P1_U5492;
  assign new_P1_U5514 = ~new_P1_U3974 | ~new_P1_U3953;
  assign new_P1_U5515 = ~new_P1_U3598 | ~new_P1_U5492;
  assign new_P1_U5516 = ~new_P1_U3975 | ~new_P1_U3953;
  assign new_P1_U5517 = ~new_P1_U3599 | ~new_P1_U5492;
  assign new_P1_U5518 = ~new_P1_U3976 | ~new_P1_U3953;
  assign new_P1_U5519 = ~new_P1_U3600 | ~new_P1_U5492;
  assign new_P1_U5520 = ~new_P1_U3977 | ~new_P1_U3953;
  assign new_P1_U5521 = ~new_P1_U3601 | ~new_P1_U5492;
  assign new_P1_U5522 = ~new_P1_U3978 | ~new_P1_U3953;
  assign new_P1_U5523 = ~new_P1_U3602 | ~new_P1_U5492;
  assign new_P1_U5524 = ~new_P1_U3979 | ~new_P1_U3953;
  assign new_P1_U5525 = ~new_P1_U3603 | ~new_P1_U5492;
  assign new_P1_U5526 = ~new_P1_U3980 | ~new_P1_U3953;
  assign new_P1_U5527 = ~new_P1_U3604 | ~new_P1_U5492;
  assign new_P1_U5528 = ~new_P1_U3981 | ~new_P1_U3953;
  assign new_P1_U5529 = ~new_P1_U3605 | ~new_P1_U5492;
  assign new_P1_U5530 = ~new_P1_U3982 | ~new_P1_U3953;
  assign new_P1_U5531 = ~new_P1_U3953 | ~new_P1_U3458;
  assign new_P1_U5532 = ~new_P1_U3595 | ~new_P1_U5492;
  assign new_P1_U5533 = ~new_P1_U3953 | ~new_P1_U3508;
  assign new_P1_U5534 = ~new_P1_U3607 | ~new_P1_U5492;
  assign new_P1_U5535 = ~new_P1_U3953 | ~new_P1_U3506;
  assign new_P1_U5536 = ~new_P1_U3608 | ~new_P1_U5492;
  assign new_P1_U5537 = ~new_P1_U3953 | ~new_P1_U3503;
  assign new_P1_U5538 = ~new_P1_U3609 | ~new_P1_U5492;
  assign new_P1_U5539 = ~new_P1_U3953 | ~new_P1_U3500;
  assign new_P1_U5540 = ~new_P1_U3610 | ~new_P1_U5492;
  assign new_P1_U5541 = ~new_P1_U3953 | ~new_P1_U3497;
  assign new_P1_U5542 = ~new_P1_U3611 | ~new_P1_U5492;
  assign new_P1_U5543 = ~new_P1_U3953 | ~new_P1_U3494;
  assign new_P1_U5544 = ~new_P1_U3612 | ~new_P1_U5492;
  assign new_P1_U5545 = ~new_P1_U3953 | ~new_P1_U3491;
  assign new_P1_U5546 = ~new_P1_U3613 | ~new_P1_U5492;
  assign new_P1_U5547 = ~new_P1_U3953 | ~new_P1_U3488;
  assign new_P1_U5548 = ~new_P1_U3614 | ~new_P1_U5492;
  assign new_P1_U5549 = ~new_P1_U3953 | ~new_P1_U3485;
  assign new_P1_U5550 = ~new_P1_U3615 | ~new_P1_U5492;
  assign new_P1_U5551 = ~new_P1_U3953 | ~new_P1_U3482;
  assign new_P1_U5552 = ~new_P1_U3616 | ~new_P1_U5492;
  assign new_P1_U5553 = ~new_P1_U3953 | ~new_P1_U3455;
  assign new_P1_U5554 = ~new_P1_U3606 | ~new_P1_U5492;
  assign new_P1_U5555 = ~new_P1_U3953 | ~new_P1_U3450;
  assign new_P1_U5556 = ~new_P1_U3617 | ~new_P1_U5492;
  assign new_P1_U5557 = ~new_P1_U3479 | ~new_P1_U5492;
  assign new_P1_U5558 = ~new_P1_U3953 | ~new_P1_U3586;
  assign new_P1_U5559 = ~new_P1_U5677 | ~new_P1_U3084;
  assign new_P1_U5560 = ~new_P1_U3476 | ~new_P1_U5492;
  assign new_P1_U5561 = ~new_P1_U3953 | ~new_P1_U3587;
  assign new_P1_U5562 = ~new_P1_U5677 | ~new_P1_U3070;
  assign new_P1_U5563 = ~new_P1_U3473 | ~new_P1_U5492;
  assign new_P1_U5564 = ~new_P1_U3953 | ~new_P1_U3588;
  assign new_P1_U5565 = ~new_P1_U5677 | ~new_P1_U3071;
  assign new_P1_U5566 = ~new_P1_U3470 | ~new_P1_U5492;
  assign new_P1_U5567 = ~new_P1_U3953 | ~new_P1_U3589;
  assign new_P1_U5568 = ~new_P1_U5677 | ~new_P1_U3067;
  assign new_P1_U5569 = ~new_P1_U3467 | ~new_P1_U5492;
  assign new_P1_U5570 = ~new_P1_U3953 | ~new_P1_U3590;
  assign new_P1_U5571 = ~new_P1_U5677 | ~new_P1_U3060;
  assign new_P1_U5572 = ~new_P1_U3464 | ~new_P1_U5492;
  assign new_P1_U5573 = ~new_P1_U3953 | ~new_P1_U3591;
  assign new_P1_U5574 = ~new_P1_U5677 | ~new_P1_U3064;
  assign new_P1_U5575 = ~new_P1_U3983 | ~new_P1_U5492;
  assign new_P1_U5576 = ~new_P1_U3953 | ~new_P1_U3593;
  assign new_P1_U5577 = ~new_P1_U3984 | ~new_P1_U5492;
  assign new_P1_U5578 = ~new_P1_U3953 | ~new_P1_U3594;
  assign new_P1_U5579 = ~new_P1_U3461 | ~new_P1_U5492;
  assign new_P1_U5580 = ~new_P1_U3953 | ~new_P1_U3592;
  assign new_P1_U5581 = ~new_P1_U5677 | ~new_P1_U3068;
  assign new_P1_U5582 = ~new_P1_U3985 | ~new_P1_U5492;
  assign new_P1_U5583 = ~new_P1_U3953 | ~new_P1_U3596;
  assign new_P1_U5584 = ~new_P1_U5677 | ~new_P1_U3054;
  assign new_P1_U5585 = ~new_P1_U3974 | ~new_P1_U5492;
  assign new_P1_U5586 = ~new_P1_U3953 | ~new_P1_U3597;
  assign new_P1_U5587 = ~new_P1_U5677 | ~new_P1_U3053;
  assign new_P1_U5588 = ~new_P1_U3975 | ~new_P1_U5492;
  assign new_P1_U5589 = ~new_P1_U3953 | ~new_P1_U3598;
  assign new_P1_U5590 = ~new_P1_U5677 | ~new_P1_U3057;
  assign new_P1_U5591 = ~new_P1_U3976 | ~new_P1_U5492;
  assign new_P1_U5592 = ~new_P1_U3953 | ~new_P1_U3599;
  assign new_P1_U5593 = ~new_P1_U5677 | ~new_P1_U3058;
  assign new_P1_U5594 = ~new_P1_U3977 | ~new_P1_U5492;
  assign new_P1_U5595 = ~new_P1_U3953 | ~new_P1_U3600;
  assign new_P1_U5596 = ~new_P1_U5677 | ~new_P1_U3065;
  assign new_P1_U5597 = ~new_P1_U3978 | ~new_P1_U5492;
  assign new_P1_U5598 = ~new_P1_U3953 | ~new_P1_U3601;
  assign new_P1_U5599 = ~new_P1_U5677 | ~new_P1_U3066;
  assign new_P1_U5600 = ~new_P1_U3979 | ~new_P1_U5492;
  assign new_P1_U5601 = ~new_P1_U3953 | ~new_P1_U3602;
  assign new_P1_U5602 = ~new_P1_U5677 | ~new_P1_U3061;
  assign new_P1_U5603 = ~new_P1_U3980 | ~new_P1_U5492;
  assign new_P1_U5604 = ~new_P1_U3953 | ~new_P1_U3603;
  assign new_P1_U5605 = ~new_P1_U5677 | ~new_P1_U3075;
  assign new_P1_U5606 = ~new_P1_U3981 | ~new_P1_U5492;
  assign new_P1_U5607 = ~new_P1_U3953 | ~new_P1_U3604;
  assign new_P1_U5608 = ~new_P1_U5677 | ~new_P1_U3076;
  assign new_P1_U5609 = ~new_P1_U3982 | ~new_P1_U5492;
  assign new_P1_U5610 = ~new_P1_U3953 | ~new_P1_U3605;
  assign new_P1_U5611 = ~new_P1_U5677 | ~new_P1_U3081;
  assign new_P1_U5612 = ~new_P1_U3458 | ~new_P1_U5492;
  assign new_P1_U5613 = ~new_P1_U3953 | ~new_P1_U3595;
  assign new_P1_U5614 = ~new_P1_U5677 | ~new_P1_U3078;
  assign new_P1_U5615 = ~new_P1_U3508 | ~new_P1_U5492;
  assign new_P1_U5616 = ~new_P1_U3953 | ~new_P1_U3607;
  assign new_P1_U5617 = ~new_P1_U5677 | ~new_P1_U3082;
  assign new_P1_U5618 = ~new_P1_U3506 | ~new_P1_U5492;
  assign new_P1_U5619 = ~new_P1_U3953 | ~new_P1_U3608;
  assign new_P1_U5620 = ~new_P1_U5677 | ~new_P1_U3069;
  assign new_P1_U5621 = ~new_P1_U3503 | ~new_P1_U5492;
  assign new_P1_U5622 = ~new_P1_U3953 | ~new_P1_U3609;
  assign new_P1_U5623 = ~new_P1_U5677 | ~new_P1_U3073;
  assign new_P1_U5624 = ~new_P1_U3500 | ~new_P1_U5492;
  assign new_P1_U5625 = ~new_P1_U3953 | ~new_P1_U3610;
  assign new_P1_U5626 = ~new_P1_U5677 | ~new_P1_U3074;
  assign new_P1_U5627 = ~new_P1_U3497 | ~new_P1_U5492;
  assign new_P1_U5628 = ~new_P1_U3953 | ~new_P1_U3611;
  assign new_P1_U5629 = ~new_P1_U5677 | ~new_P1_U3079;
  assign new_P1_U5630 = ~new_P1_U3494 | ~new_P1_U5492;
  assign new_P1_U5631 = ~new_P1_U3953 | ~new_P1_U3612;
  assign new_P1_U5632 = ~new_P1_U5677 | ~new_P1_U3080;
  assign new_P1_U5633 = ~new_P1_U3491 | ~new_P1_U5492;
  assign new_P1_U5634 = ~new_P1_U3953 | ~new_P1_U3613;
  assign new_P1_U5635 = ~new_P1_U5677 | ~new_P1_U3072;
  assign new_P1_U5636 = ~new_P1_U3488 | ~new_P1_U5492;
  assign new_P1_U5637 = ~new_P1_U3953 | ~new_P1_U3614;
  assign new_P1_U5638 = ~new_P1_U5677 | ~new_P1_U3063;
  assign new_P1_U5639 = ~new_P1_U3485 | ~new_P1_U5492;
  assign new_P1_U5640 = ~new_P1_U3953 | ~new_P1_U3615;
  assign new_P1_U5641 = ~new_P1_U5677 | ~new_P1_U3062;
  assign new_P1_U5642 = ~new_P1_U3482 | ~new_P1_U5492;
  assign new_P1_U5643 = ~new_P1_U3953 | ~new_P1_U3616;
  assign new_P1_U5644 = ~new_P1_U5677 | ~new_P1_U3083;
  assign new_P1_U5645 = ~new_P1_U3455 | ~new_P1_U5492;
  assign new_P1_U5646 = ~new_P1_U3953 | ~new_P1_U3606;
  assign new_P1_U5647 = ~new_P1_U5677 | ~new_P1_U3077;
  assign new_P1_U5648 = ~new_P1_U3450 | ~new_P1_U5492;
  assign new_P1_U5649 = ~new_P1_U3953 | ~new_P1_U3617;
  assign new_P1_U5650 = ~new_P1_U3864 | ~new_P1_U3052 | ~new_P1_U5662 | ~new_P1_U3950;
  assign new_P1_U5651 = ~n1330 | ~new_P1_U5091;
  assign new_P1_U5652 = ~new_P1_U3865 | ~new_P1_U5091 | ~new_P1_U5090;
  assign new_P1_U5653 = ~new_P1_U3997 | ~new_P1_U3430;
  assign new_P1_U5654 = ~new_P1_U3972 | ~new_P1_U3997;
  assign new_P1_U5655 = ~new_P1_U5653 | ~new_P1_U3995;
  assign new_P1_U5656 = ~new_P1_U5654 | ~new_P1_U3996;
  assign new_P1_U5657 = ~new_P1_R1207_U14 | ~new_P1_U3958;
  assign new_P1_U5658 = ~new_P1_R1192_U14 | ~new_P1_U3959;
  assign new_P1_U5659 = ~new_P1_R1150_U14 | ~new_P1_U3961;
  assign new_P1_U5660 = ~new_P1_R1117_U14 | ~new_P1_U3963;
  assign new_P1_U5661 = ~new_P1_U5666 | ~new_P1_U5672;
  assign new_P1_U5662 = ~new_P1_U5693 | ~new_P1_U6170 | ~new_P1_U6169;
  assign new_P1_U5663 = ~new_P1_U3442 | ~new_P1_U3438;
  assign new_P1_U5664 = ~P1_IR_REG_24_ | ~new_P1_U3910;
  assign new_P1_U5665 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U17;
  assign new_P1_U5666 = ~new_P1_U3435;
  assign new_P1_U5667 = ~P1_IR_REG_25_ | ~new_P1_U3910;
  assign new_P1_U5668 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U170;
  assign new_P1_U5669 = ~new_P1_U3436;
  assign new_P1_U5670 = ~P1_IR_REG_26_ | ~new_P1_U3910;
  assign new_P1_U5671 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U18;
  assign new_P1_U5672 = ~new_P1_U3437;
  assign new_P1_U5673 = ~new_P1_U3050 | ~new_P1_U3359;
  assign new_P1_U5674 = ~P1_B_REG | ~new_P1_U4003 | ~new_P1_U5666;
  assign new_P1_U5675 = ~P1_IR_REG_23_ | ~new_P1_U3910;
  assign new_P1_U5676 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U16;
  assign new_P1_U5677 = ~new_P1_U3438;
  assign new_P1_U5678 = ~P1_D_REG_0_ | ~new_P1_U3911;
  assign new_P1_U5679 = ~new_P1_U3992 | ~new_P1_U4103;
  assign new_P1_U5680 = ~P1_D_REG_1_ | ~new_P1_U3911;
  assign new_P1_U5681 = ~new_P1_U3992 | ~new_P1_U4104;
  assign new_P1_U5682 = ~P1_IR_REG_22_ | ~new_P1_U3910;
  assign new_P1_U5683 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U15;
  assign new_P1_U5684 = ~new_P1_U3443;
  assign new_P1_U5685 = ~P1_IR_REG_19_ | ~new_P1_U3910;
  assign new_P1_U5686 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U13;
  assign new_P1_U5687 = ~new_P1_U3442;
  assign new_P1_U5688 = ~P1_IR_REG_20_ | ~new_P1_U3910;
  assign new_P1_U5689 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U14;
  assign new_P1_U5690 = ~new_P1_U3441;
  assign new_P1_U5691 = ~P1_IR_REG_21_ | ~new_P1_U3910;
  assign new_P1_U5692 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U173;
  assign new_P1_U5693 = ~new_P1_U3447;
  assign new_P1_U5694 = ~P1_IR_REG_0_ | ~new_P1_U3910;
  assign new_P1_U5695 = ~P1_IR_REG_31_ | ~P1_IR_REG_0_;
  assign new_P1_U5696 = ~new_P1_U3448;
  assign new_P1_U5697 = ~P1_IR_REG_28_ | ~new_P1_U3910;
  assign new_P1_U5698 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U19;
  assign new_P1_U5699 = ~new_P1_U3446;
  assign new_P1_U5700 = ~P1_IR_REG_27_ | ~new_P1_U3910;
  assign new_P1_U5701 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U42;
  assign new_P1_U5702 = ~new_P1_U3449;
  assign new_P1_U5703 = ~new_U88 | ~new_P1_U3912;
  assign new_P1_U5704 = ~new_P1_U3971 | ~new_P1_U3448;
  assign new_P1_U5705 = ~new_P1_U3450;
  assign new_P1_U5706 = ~P1_IR_REG_30_ | ~new_P1_U3910;
  assign new_P1_U5707 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U165;
  assign new_P1_U5708 = ~new_P1_U3444;
  assign new_P1_U5709 = ~P1_IR_REG_29_ | ~new_P1_U3910;
  assign new_P1_U5710 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U20;
  assign new_P1_U5711 = ~new_P1_U3445;
  assign new_P1_U5712 = ~new_P1_U3443 | ~new_P1_U5693;
  assign new_P1_U5713 = ~new_P1_U5684 | ~new_P1_U4135;
  assign new_P1_U5714 = ~P1_D_REG_1_ | ~new_P1_U4101;
  assign new_P1_U5715 = ~new_P1_U4104 | ~new_P1_U3360;
  assign new_P1_U5716 = ~new_P1_U3452;
  assign new_P1_U5717 = ~new_P1_U5661 | ~new_P1_U3360;
  assign new_P1_U5718 = ~P1_D_REG_0_ | ~new_P1_U4101;
  assign new_P1_U5719 = ~new_P1_U3451;
  assign new_P1_U5720 = ~P1_REG0_REG_0_ | ~new_P1_U3913;
  assign new_P1_U5721 = ~new_P1_U3991 | ~new_P1_U4155;
  assign new_P1_U5722 = ~P1_IR_REG_1_ | ~new_P1_U3910;
  assign new_P1_U5723 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U40;
  assign new_P1_U5724 = ~new_U77 | ~new_P1_U3912;
  assign new_P1_U5725 = ~new_P1_U3454 | ~new_P1_U3971;
  assign new_P1_U5726 = ~new_P1_U3455;
  assign new_P1_U5727 = ~P1_REG0_REG_1_ | ~new_P1_U3913;
  assign new_P1_U5728 = ~new_P1_U3991 | ~new_P1_U4179;
  assign new_P1_U5729 = ~P1_IR_REG_2_ | ~new_P1_U3910;
  assign new_P1_U5730 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U21;
  assign new_P1_U5731 = ~new_U66 | ~new_P1_U3912;
  assign new_P1_U5732 = ~new_P1_U3457 | ~new_P1_U3971;
  assign new_P1_U5733 = ~new_P1_U3458;
  assign new_P1_U5734 = ~P1_REG0_REG_2_ | ~new_P1_U3913;
  assign new_P1_U5735 = ~new_P1_U3991 | ~new_P1_U4198;
  assign new_P1_U5736 = ~P1_IR_REG_3_ | ~new_P1_U3910;
  assign new_P1_U5737 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U22;
  assign new_P1_U5738 = ~new_U63 | ~new_P1_U3912;
  assign new_P1_U5739 = ~new_P1_U3460 | ~new_P1_U3971;
  assign new_P1_U5740 = ~new_P1_U3461;
  assign new_P1_U5741 = ~P1_REG0_REG_3_ | ~new_P1_U3913;
  assign new_P1_U5742 = ~new_P1_U3991 | ~new_P1_U4217;
  assign new_P1_U5743 = ~P1_IR_REG_4_ | ~new_P1_U3910;
  assign new_P1_U5744 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U23;
  assign new_P1_U5745 = ~new_U62 | ~new_P1_U3912;
  assign new_P1_U5746 = ~new_P1_U3463 | ~new_P1_U3971;
  assign new_P1_U5747 = ~new_P1_U3464;
  assign new_P1_U5748 = ~P1_REG0_REG_4_ | ~new_P1_U3913;
  assign new_P1_U5749 = ~new_P1_U3991 | ~new_P1_U4236;
  assign new_P1_U5750 = ~P1_IR_REG_5_ | ~new_P1_U3910;
  assign new_P1_U5751 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U162;
  assign new_P1_U5752 = ~new_U61 | ~new_P1_U3912;
  assign new_P1_U5753 = ~new_P1_U3466 | ~new_P1_U3971;
  assign new_P1_U5754 = ~new_P1_U3467;
  assign new_P1_U5755 = ~P1_REG0_REG_5_ | ~new_P1_U3913;
  assign new_P1_U5756 = ~new_P1_U3991 | ~new_P1_U4255;
  assign new_P1_U5757 = ~P1_IR_REG_6_ | ~new_P1_U3910;
  assign new_P1_U5758 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U24;
  assign new_P1_U5759 = ~new_U60 | ~new_P1_U3912;
  assign new_P1_U5760 = ~new_P1_U3469 | ~new_P1_U3971;
  assign new_P1_U5761 = ~new_P1_U3470;
  assign new_P1_U5762 = ~P1_REG0_REG_6_ | ~new_P1_U3913;
  assign new_P1_U5763 = ~new_P1_U3991 | ~new_P1_U4274;
  assign new_P1_U5764 = ~P1_IR_REG_7_ | ~new_P1_U3910;
  assign new_P1_U5765 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U25;
  assign new_P1_U5766 = ~new_U59 | ~new_P1_U3912;
  assign new_P1_U5767 = ~new_P1_U3472 | ~new_P1_U3971;
  assign new_P1_U5768 = ~new_P1_U3473;
  assign new_P1_U5769 = ~P1_REG0_REG_7_ | ~new_P1_U3913;
  assign new_P1_U5770 = ~new_P1_U3991 | ~new_P1_U4293;
  assign new_P1_U5771 = ~P1_IR_REG_8_ | ~new_P1_U3910;
  assign new_P1_U5772 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U26;
  assign new_P1_U5773 = ~new_U58 | ~new_P1_U3912;
  assign new_P1_U5774 = ~new_P1_U3475 | ~new_P1_U3971;
  assign new_P1_U5775 = ~new_P1_U3476;
  assign new_P1_U5776 = ~P1_REG0_REG_8_ | ~new_P1_U3913;
  assign new_P1_U5777 = ~new_P1_U3991 | ~new_P1_U4312;
  assign new_P1_U5778 = ~P1_IR_REG_9_ | ~new_P1_U3910;
  assign new_P1_U5779 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U160;
  assign new_P1_U5780 = ~new_U57 | ~new_P1_U3912;
  assign new_P1_U5781 = ~new_P1_U3478 | ~new_P1_U3971;
  assign new_P1_U5782 = ~new_P1_U3479;
  assign new_P1_U5783 = ~P1_REG0_REG_9_ | ~new_P1_U3913;
  assign new_P1_U5784 = ~new_P1_U3991 | ~new_P1_U4331;
  assign new_P1_U5785 = ~P1_IR_REG_10_ | ~new_P1_U3910;
  assign new_P1_U5786 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U6;
  assign new_P1_U5787 = ~new_U87 | ~new_P1_U3912;
  assign new_P1_U5788 = ~new_P1_U3481 | ~new_P1_U3971;
  assign new_P1_U5789 = ~new_P1_U3482;
  assign new_P1_U5790 = ~P1_REG0_REG_10_ | ~new_P1_U3913;
  assign new_P1_U5791 = ~new_P1_U3991 | ~new_P1_U4350;
  assign new_P1_U5792 = ~P1_IR_REG_11_ | ~new_P1_U3910;
  assign new_P1_U5793 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U7;
  assign new_P1_U5794 = ~new_U86 | ~new_P1_U3912;
  assign new_P1_U5795 = ~new_P1_U3484 | ~new_P1_U3971;
  assign new_P1_U5796 = ~new_P1_U3485;
  assign new_P1_U5797 = ~P1_REG0_REG_11_ | ~new_P1_U3913;
  assign new_P1_U5798 = ~new_P1_U3991 | ~new_P1_U4369;
  assign new_P1_U5799 = ~P1_IR_REG_12_ | ~new_P1_U3910;
  assign new_P1_U5800 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U8;
  assign new_P1_U5801 = ~new_U85 | ~new_P1_U3912;
  assign new_P1_U5802 = ~new_P1_U3487 | ~new_P1_U3971;
  assign new_P1_U5803 = ~new_P1_U3488;
  assign new_P1_U5804 = ~P1_REG0_REG_12_ | ~new_P1_U3913;
  assign new_P1_U5805 = ~new_P1_U3991 | ~new_P1_U4388;
  assign new_P1_U5806 = ~P1_IR_REG_13_ | ~new_P1_U3910;
  assign new_P1_U5807 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U179;
  assign new_P1_U5808 = ~new_U84 | ~new_P1_U3912;
  assign new_P1_U5809 = ~new_P1_U3490 | ~new_P1_U3971;
  assign new_P1_U5810 = ~new_P1_U3491;
  assign new_P1_U5811 = ~P1_REG0_REG_13_ | ~new_P1_U3913;
  assign new_P1_U5812 = ~new_P1_U3991 | ~new_P1_U4407;
  assign new_P1_U5813 = ~P1_IR_REG_14_ | ~new_P1_U3910;
  assign new_P1_U5814 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U9;
  assign new_P1_U5815 = ~new_U83 | ~new_P1_U3912;
  assign new_P1_U5816 = ~new_P1_U3493 | ~new_P1_U3971;
  assign new_P1_U5817 = ~new_P1_U3494;
  assign new_P1_U5818 = ~P1_REG0_REG_14_ | ~new_P1_U3913;
  assign new_P1_U5819 = ~new_P1_U3991 | ~new_P1_U4426;
  assign new_P1_U5820 = ~P1_IR_REG_15_ | ~new_P1_U3910;
  assign new_P1_U5821 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U10;
  assign new_P1_U5822 = ~new_U82 | ~new_P1_U3912;
  assign new_P1_U5823 = ~new_P1_U3496 | ~new_P1_U3971;
  assign new_P1_U5824 = ~new_P1_U3497;
  assign new_P1_U5825 = ~P1_REG0_REG_15_ | ~new_P1_U3913;
  assign new_P1_U5826 = ~new_P1_U3991 | ~new_P1_U4445;
  assign new_P1_U5827 = ~P1_IR_REG_16_ | ~new_P1_U3910;
  assign new_P1_U5828 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U11;
  assign new_P1_U5829 = ~new_U81 | ~new_P1_U3912;
  assign new_P1_U5830 = ~new_P1_U3499 | ~new_P1_U3971;
  assign new_P1_U5831 = ~new_P1_U3500;
  assign new_P1_U5832 = ~P1_REG0_REG_16_ | ~new_P1_U3913;
  assign new_P1_U5833 = ~new_P1_U3991 | ~new_P1_U4464;
  assign new_P1_U5834 = ~P1_IR_REG_17_ | ~new_P1_U3910;
  assign new_P1_U5835 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U177;
  assign new_P1_U5836 = ~new_U80 | ~new_P1_U3912;
  assign new_P1_U5837 = ~new_P1_U3502 | ~new_P1_U3971;
  assign new_P1_U5838 = ~new_P1_U3503;
  assign new_P1_U5839 = ~P1_REG0_REG_17_ | ~new_P1_U3913;
  assign new_P1_U5840 = ~new_P1_U3991 | ~new_P1_U4483;
  assign new_P1_U5841 = ~P1_IR_REG_18_ | ~new_P1_U3910;
  assign new_P1_U5842 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U12;
  assign new_P1_U5843 = ~new_U79 | ~new_P1_U3912;
  assign new_P1_U5844 = ~new_P1_U3505 | ~new_P1_U3971;
  assign new_P1_U5845 = ~new_P1_U3506;
  assign new_P1_U5846 = ~P1_REG0_REG_18_ | ~new_P1_U3913;
  assign new_P1_U5847 = ~new_P1_U3991 | ~new_P1_U4502;
  assign new_P1_U5848 = ~new_U78 | ~new_P1_U3912;
  assign new_P1_U5849 = ~new_P1_U3971 | ~new_P1_U3442;
  assign new_P1_U5850 = ~new_P1_U3508;
  assign new_P1_U5851 = ~P1_REG0_REG_19_ | ~new_P1_U3913;
  assign new_P1_U5852 = ~new_P1_U3991 | ~new_P1_U4521;
  assign new_P1_U5853 = ~P1_REG0_REG_20_ | ~new_P1_U3913;
  assign new_P1_U5854 = ~new_P1_U3991 | ~new_P1_U4540;
  assign new_P1_U5855 = ~P1_REG0_REG_21_ | ~new_P1_U3913;
  assign new_P1_U5856 = ~new_P1_U3991 | ~new_P1_U4559;
  assign new_P1_U5857 = ~P1_REG0_REG_22_ | ~new_P1_U3913;
  assign new_P1_U5858 = ~new_P1_U3991 | ~new_P1_U4578;
  assign new_P1_U5859 = ~P1_REG0_REG_23_ | ~new_P1_U3913;
  assign new_P1_U5860 = ~new_P1_U3991 | ~new_P1_U4597;
  assign new_P1_U5861 = ~P1_REG0_REG_24_ | ~new_P1_U3913;
  assign new_P1_U5862 = ~new_P1_U3991 | ~new_P1_U4616;
  assign new_P1_U5863 = ~P1_REG0_REG_25_ | ~new_P1_U3913;
  assign new_P1_U5864 = ~new_P1_U3991 | ~new_P1_U4635;
  assign new_P1_U5865 = ~P1_REG0_REG_26_ | ~new_P1_U3913;
  assign new_P1_U5866 = ~new_P1_U3991 | ~new_P1_U4654;
  assign new_P1_U5867 = ~P1_REG0_REG_27_ | ~new_P1_U3913;
  assign new_P1_U5868 = ~new_P1_U3991 | ~new_P1_U4673;
  assign new_P1_U5869 = ~P1_REG0_REG_28_ | ~new_P1_U3913;
  assign new_P1_U5870 = ~new_P1_U3991 | ~new_P1_U4692;
  assign new_P1_U5871 = ~P1_REG0_REG_29_ | ~new_P1_U3913;
  assign new_P1_U5872 = ~new_P1_U3991 | ~new_P1_U4712;
  assign new_P1_U5873 = ~P1_REG0_REG_30_ | ~new_P1_U3913;
  assign new_P1_U5874 = ~new_P1_U3991 | ~new_P1_U4719;
  assign new_P1_U5875 = ~P1_REG0_REG_31_ | ~new_P1_U3913;
  assign new_P1_U5876 = ~new_P1_U3991 | ~new_P1_U4722;
  assign new_P1_U5877 = ~P1_REG1_REG_0_ | ~new_P1_U3914;
  assign new_P1_U5878 = ~new_P1_U3990 | ~new_P1_U4155;
  assign new_P1_U5879 = ~P1_REG1_REG_1_ | ~new_P1_U3914;
  assign new_P1_U5880 = ~new_P1_U3990 | ~new_P1_U4179;
  assign new_P1_U5881 = ~P1_REG1_REG_2_ | ~new_P1_U3914;
  assign new_P1_U5882 = ~new_P1_U3990 | ~new_P1_U4198;
  assign new_P1_U5883 = ~P1_REG1_REG_3_ | ~new_P1_U3914;
  assign new_P1_U5884 = ~new_P1_U3990 | ~new_P1_U4217;
  assign new_P1_U5885 = ~P1_REG1_REG_4_ | ~new_P1_U3914;
  assign new_P1_U5886 = ~new_P1_U3990 | ~new_P1_U4236;
  assign new_P1_U5887 = ~P1_REG1_REG_5_ | ~new_P1_U3914;
  assign new_P1_U5888 = ~new_P1_U3990 | ~new_P1_U4255;
  assign new_P1_U5889 = ~P1_REG1_REG_6_ | ~new_P1_U3914;
  assign new_P1_U5890 = ~new_P1_U3990 | ~new_P1_U4274;
  assign new_P1_U5891 = ~P1_REG1_REG_7_ | ~new_P1_U3914;
  assign new_P1_U5892 = ~new_P1_U3990 | ~new_P1_U4293;
  assign new_P1_U5893 = ~P1_REG1_REG_8_ | ~new_P1_U3914;
  assign new_P1_U5894 = ~new_P1_U3990 | ~new_P1_U4312;
  assign new_P1_U5895 = ~P1_REG1_REG_9_ | ~new_P1_U3914;
  assign new_P1_U5896 = ~new_P1_U3990 | ~new_P1_U4331;
  assign new_P1_U5897 = ~P1_REG1_REG_10_ | ~new_P1_U3914;
  assign new_P1_U5898 = ~new_P1_U3990 | ~new_P1_U4350;
  assign new_P1_U5899 = ~P1_REG1_REG_11_ | ~new_P1_U3914;
  assign new_P1_U5900 = ~new_P1_U3990 | ~new_P1_U4369;
  assign new_P1_U5901 = ~P1_REG1_REG_12_ | ~new_P1_U3914;
  assign new_P1_U5902 = ~new_P1_U3990 | ~new_P1_U4388;
  assign new_P1_U5903 = ~P1_REG1_REG_13_ | ~new_P1_U3914;
  assign new_P1_U5904 = ~new_P1_U3990 | ~new_P1_U4407;
  assign new_P1_U5905 = ~P1_REG1_REG_14_ | ~new_P1_U3914;
  assign new_P1_U5906 = ~new_P1_U3990 | ~new_P1_U4426;
  assign new_P1_U5907 = ~P1_REG1_REG_15_ | ~new_P1_U3914;
  assign new_P1_U5908 = ~new_P1_U3990 | ~new_P1_U4445;
  assign new_P1_U5909 = ~P1_REG1_REG_16_ | ~new_P1_U3914;
  assign new_P1_U5910 = ~new_P1_U3990 | ~new_P1_U4464;
  assign new_P1_U5911 = ~P1_REG1_REG_17_ | ~new_P1_U3914;
  assign new_P1_U5912 = ~new_P1_U3990 | ~new_P1_U4483;
  assign new_P1_U5913 = ~P1_REG1_REG_18_ | ~new_P1_U3914;
  assign new_P1_U5914 = ~new_P1_U3990 | ~new_P1_U4502;
  assign new_P1_U5915 = ~P1_REG1_REG_19_ | ~new_P1_U3914;
  assign new_P1_U5916 = ~new_P1_U3990 | ~new_P1_U4521;
  assign new_P1_U5917 = ~P1_REG1_REG_20_ | ~new_P1_U3914;
  assign new_P1_U5918 = ~new_P1_U3990 | ~new_P1_U4540;
  assign new_P1_U5919 = ~P1_REG1_REG_21_ | ~new_P1_U3914;
  assign new_P1_U5920 = ~new_P1_U3990 | ~new_P1_U4559;
  assign new_P1_U5921 = ~P1_REG1_REG_22_ | ~new_P1_U3914;
  assign new_P1_U5922 = ~new_P1_U3990 | ~new_P1_U4578;
  assign new_P1_U5923 = ~P1_REG1_REG_23_ | ~new_P1_U3914;
  assign new_P1_U5924 = ~new_P1_U3990 | ~new_P1_U4597;
  assign new_P1_U5925 = ~P1_REG1_REG_24_ | ~new_P1_U3914;
  assign new_P1_U5926 = ~new_P1_U3990 | ~new_P1_U4616;
  assign new_P1_U5927 = ~P1_REG1_REG_25_ | ~new_P1_U3914;
  assign new_P1_U5928 = ~new_P1_U3990 | ~new_P1_U4635;
  assign new_P1_U5929 = ~P1_REG1_REG_26_ | ~new_P1_U3914;
  assign new_P1_U5930 = ~new_P1_U3990 | ~new_P1_U4654;
  assign new_P1_U5931 = ~P1_REG1_REG_27_ | ~new_P1_U3914;
  assign new_P1_U5932 = ~new_P1_U3990 | ~new_P1_U4673;
  assign new_P1_U5933 = ~P1_REG1_REG_28_ | ~new_P1_U3914;
  assign new_P1_U5934 = ~new_P1_U3990 | ~new_P1_U4692;
  assign new_P1_U5935 = ~P1_REG1_REG_29_ | ~new_P1_U3914;
  assign new_P1_U5936 = ~new_P1_U3990 | ~new_P1_U4712;
  assign new_P1_U5937 = ~P1_REG1_REG_30_ | ~new_P1_U3914;
  assign new_P1_U5938 = ~new_P1_U3990 | ~new_P1_U4719;
  assign new_P1_U5939 = ~P1_REG1_REG_31_ | ~new_P1_U3914;
  assign new_P1_U5940 = ~new_P1_U3990 | ~new_P1_U4722;
  assign new_P1_U5941 = ~P1_REG2_REG_0_ | ~new_P1_U3417;
  assign new_P1_U5942 = ~new_P1_U3989 | ~new_P1_U3374;
  assign new_P1_U5943 = ~P1_REG2_REG_1_ | ~new_P1_U3417;
  assign new_P1_U5944 = ~new_P1_U3989 | ~new_P1_U3376;
  assign new_P1_U5945 = ~P1_REG2_REG_2_ | ~new_P1_U3417;
  assign new_P1_U5946 = ~new_P1_U3989 | ~new_P1_U3377;
  assign new_P1_U5947 = ~P1_REG2_REG_3_ | ~new_P1_U3417;
  assign new_P1_U5948 = ~new_P1_U3989 | ~new_P1_U3378;
  assign new_P1_U5949 = ~P1_REG2_REG_4_ | ~new_P1_U3417;
  assign new_P1_U5950 = ~new_P1_U3989 | ~new_P1_U3379;
  assign new_P1_U5951 = ~P1_REG2_REG_5_ | ~new_P1_U3417;
  assign new_P1_U5952 = ~new_P1_U3989 | ~new_P1_U3380;
  assign new_P1_U5953 = ~P1_REG2_REG_6_ | ~new_P1_U3417;
  assign new_P1_U5954 = ~new_P1_U3989 | ~new_P1_U3381;
  assign new_P1_U5955 = ~P1_REG2_REG_7_ | ~new_P1_U3417;
  assign new_P1_U5956 = ~new_P1_U3989 | ~new_P1_U3382;
  assign new_P1_U5957 = ~P1_REG2_REG_8_ | ~new_P1_U3417;
  assign new_P1_U5958 = ~new_P1_U3989 | ~new_P1_U3383;
  assign new_P1_U5959 = ~P1_REG2_REG_9_ | ~new_P1_U3417;
  assign new_P1_U5960 = ~new_P1_U3989 | ~new_P1_U3384;
  assign new_P1_U5961 = ~P1_REG2_REG_10_ | ~new_P1_U3417;
  assign new_P1_U5962 = ~new_P1_U3989 | ~new_P1_U3385;
  assign new_P1_U5963 = ~P1_REG2_REG_11_ | ~new_P1_U3417;
  assign new_P1_U5964 = ~new_P1_U3989 | ~new_P1_U3386;
  assign new_P1_U5965 = ~P1_REG2_REG_12_ | ~new_P1_U3417;
  assign new_P1_U5966 = ~new_P1_U3989 | ~new_P1_U3387;
  assign new_P1_U5967 = ~P1_REG2_REG_13_ | ~new_P1_U3417;
  assign new_P1_U5968 = ~new_P1_U3989 | ~new_P1_U3388;
  assign new_P1_U5969 = ~P1_REG2_REG_14_ | ~new_P1_U3417;
  assign new_P1_U5970 = ~new_P1_U3989 | ~new_P1_U3389;
  assign new_P1_U5971 = ~P1_REG2_REG_15_ | ~new_P1_U3417;
  assign new_P1_U5972 = ~new_P1_U3989 | ~new_P1_U3390;
  assign new_P1_U5973 = ~P1_REG2_REG_16_ | ~new_P1_U3417;
  assign new_P1_U5974 = ~new_P1_U3989 | ~new_P1_U3391;
  assign new_P1_U5975 = ~P1_REG2_REG_17_ | ~new_P1_U3417;
  assign new_P1_U5976 = ~new_P1_U3989 | ~new_P1_U3392;
  assign new_P1_U5977 = ~P1_REG2_REG_18_ | ~new_P1_U3417;
  assign new_P1_U5978 = ~new_P1_U3989 | ~new_P1_U3393;
  assign new_P1_U5979 = ~P1_REG2_REG_19_ | ~new_P1_U3417;
  assign new_P1_U5980 = ~new_P1_U3989 | ~new_P1_U3394;
  assign new_P1_U5981 = ~P1_REG2_REG_20_ | ~new_P1_U3417;
  assign new_P1_U5982 = ~new_P1_U3989 | ~new_P1_U3396;
  assign new_P1_U5983 = ~P1_REG2_REG_21_ | ~new_P1_U3417;
  assign new_P1_U5984 = ~new_P1_U3989 | ~new_P1_U3398;
  assign new_P1_U5985 = ~P1_REG2_REG_22_ | ~new_P1_U3417;
  assign new_P1_U5986 = ~new_P1_U3989 | ~new_P1_U3400;
  assign new_P1_U5987 = ~P1_REG2_REG_23_ | ~new_P1_U3417;
  assign new_P1_U5988 = ~new_P1_U3989 | ~new_P1_U3402;
  assign new_P1_U5989 = ~P1_REG2_REG_24_ | ~new_P1_U3417;
  assign new_P1_U5990 = ~new_P1_U3989 | ~new_P1_U3404;
  assign new_P1_U5991 = ~P1_REG2_REG_25_ | ~new_P1_U3417;
  assign new_P1_U5992 = ~new_P1_U3989 | ~new_P1_U3406;
  assign new_P1_U5993 = ~P1_REG2_REG_26_ | ~new_P1_U3417;
  assign new_P1_U5994 = ~new_P1_U3989 | ~new_P1_U3408;
  assign new_P1_U5995 = ~P1_REG2_REG_27_ | ~new_P1_U3417;
  assign new_P1_U5996 = ~new_P1_U3989 | ~new_P1_U3410;
  assign new_P1_U5997 = ~P1_REG2_REG_28_ | ~new_P1_U3417;
  assign new_P1_U5998 = ~new_P1_U3989 | ~new_P1_U3412;
  assign new_P1_U5999 = ~P1_REG2_REG_29_ | ~new_P1_U3417;
  assign new_P1_U6000 = ~new_P1_U3989 | ~new_P1_U4708;
  assign new_P1_U6001 = ~P1_REG2_REG_30_ | ~new_P1_U3417;
  assign new_P1_U6002 = ~new_P1_U3993 | ~new_P1_U3989;
  assign new_P1_U6003 = ~P1_REG2_REG_31_ | ~new_P1_U3417;
  assign new_P1_U6004 = ~new_P1_U3993 | ~new_P1_U3989;
  assign new_P1_U6005 = ~P1_DATAO_REG_0_ | ~new_P1_U3425;
  assign new_P1_U6006 = ~n1340 | ~new_P1_U3077;
  assign new_P1_U6007 = ~P1_DATAO_REG_1_ | ~new_P1_U3425;
  assign new_P1_U6008 = ~n1340 | ~new_P1_U3078;
  assign new_P1_U6009 = ~P1_DATAO_REG_2_ | ~new_P1_U3425;
  assign new_P1_U6010 = ~n1340 | ~new_P1_U3068;
  assign new_P1_U6011 = ~P1_DATAO_REG_3_ | ~new_P1_U3425;
  assign new_P1_U6012 = ~n1340 | ~new_P1_U3064;
  assign new_P1_U6013 = ~P1_DATAO_REG_4_ | ~new_P1_U3425;
  assign new_P1_U6014 = ~n1340 | ~new_P1_U3060;
  assign new_P1_U6015 = ~P1_DATAO_REG_5_ | ~new_P1_U3425;
  assign new_P1_U6016 = ~n1340 | ~new_P1_U3067;
  assign new_P1_U6017 = ~P1_DATAO_REG_6_ | ~new_P1_U3425;
  assign new_P1_U6018 = ~n1340 | ~new_P1_U3071;
  assign new_P1_U6019 = ~P1_DATAO_REG_7_ | ~new_P1_U3425;
  assign new_P1_U6020 = ~n1340 | ~new_P1_U3070;
  assign new_P1_U6021 = ~P1_DATAO_REG_8_ | ~new_P1_U3425;
  assign new_P1_U6022 = ~n1340 | ~new_P1_U3084;
  assign new_P1_U6023 = ~P1_DATAO_REG_9_ | ~new_P1_U3425;
  assign new_P1_U6024 = ~n1340 | ~new_P1_U3083;
  assign new_P1_U6025 = ~P1_DATAO_REG_10_ | ~new_P1_U3425;
  assign new_P1_U6026 = ~n1340 | ~new_P1_U3062;
  assign new_P1_U6027 = ~P1_DATAO_REG_11_ | ~new_P1_U3425;
  assign new_P1_U6028 = ~n1340 | ~new_P1_U3063;
  assign new_P1_U6029 = ~P1_DATAO_REG_12_ | ~new_P1_U3425;
  assign new_P1_U6030 = ~n1340 | ~new_P1_U3072;
  assign new_P1_U6031 = ~P1_DATAO_REG_13_ | ~new_P1_U3425;
  assign new_P1_U6032 = ~n1340 | ~new_P1_U3080;
  assign new_P1_U6033 = ~P1_DATAO_REG_14_ | ~new_P1_U3425;
  assign new_P1_U6034 = ~n1340 | ~new_P1_U3079;
  assign new_P1_U6035 = ~P1_DATAO_REG_15_ | ~new_P1_U3425;
  assign new_P1_U6036 = ~n1340 | ~new_P1_U3074;
  assign new_P1_U6037 = ~P1_DATAO_REG_16_ | ~new_P1_U3425;
  assign new_P1_U6038 = ~n1340 | ~new_P1_U3073;
  assign new_P1_U6039 = ~P1_DATAO_REG_17_ | ~new_P1_U3425;
  assign new_P1_U6040 = ~n1340 | ~new_P1_U3069;
  assign new_P1_U6041 = ~P1_DATAO_REG_18_ | ~new_P1_U3425;
  assign new_P1_U6042 = ~n1340 | ~new_P1_U3082;
  assign new_P1_U6043 = ~P1_DATAO_REG_19_ | ~new_P1_U3425;
  assign new_P1_U6044 = ~n1340 | ~new_P1_U3081;
  assign new_P1_U6045 = ~P1_DATAO_REG_20_ | ~new_P1_U3425;
  assign new_P1_U6046 = ~n1340 | ~new_P1_U3076;
  assign new_P1_U6047 = ~P1_DATAO_REG_21_ | ~new_P1_U3425;
  assign new_P1_U6048 = ~n1340 | ~new_P1_U3075;
  assign new_P1_U6049 = ~P1_DATAO_REG_22_ | ~new_P1_U3425;
  assign new_P1_U6050 = ~n1340 | ~new_P1_U3061;
  assign new_P1_U6051 = ~P1_DATAO_REG_23_ | ~new_P1_U3425;
  assign new_P1_U6052 = ~n1340 | ~new_P1_U3066;
  assign new_P1_U6053 = ~P1_DATAO_REG_24_ | ~new_P1_U3425;
  assign new_P1_U6054 = ~n1340 | ~new_P1_U3065;
  assign new_P1_U6055 = ~P1_DATAO_REG_25_ | ~new_P1_U3425;
  assign new_P1_U6056 = ~n1340 | ~new_P1_U3058;
  assign new_P1_U6057 = ~P1_DATAO_REG_26_ | ~new_P1_U3425;
  assign new_P1_U6058 = ~n1340 | ~new_P1_U3057;
  assign new_P1_U6059 = ~P1_DATAO_REG_27_ | ~new_P1_U3425;
  assign new_P1_U6060 = ~n1340 | ~new_P1_U3053;
  assign new_P1_U6061 = ~P1_DATAO_REG_28_ | ~new_P1_U3425;
  assign new_P1_U6062 = ~n1340 | ~new_P1_U3054;
  assign new_P1_U6063 = ~P1_DATAO_REG_29_ | ~new_P1_U3425;
  assign new_P1_U6064 = ~n1340 | ~new_P1_U3055;
  assign new_P1_U6065 = ~P1_DATAO_REG_30_ | ~new_P1_U3425;
  assign new_P1_U6066 = ~n1340 | ~new_P1_U3059;
  assign new_P1_U6067 = ~P1_DATAO_REG_31_ | ~new_P1_U3425;
  assign new_P1_U6068 = ~n1340 | ~new_P1_U3056;
  assign new_P1_U6069 = ~new_P1_U3948 | ~new_P1_U3048 | ~new_P1_U3438;
  assign new_P1_U6070 = ~new_P1_R1375_U14 | ~new_P1_U3954 | ~new_P1_U5690;
  assign new_P1_U6071 = ~new_P1_U3949 | ~new_P1_U3438 | ~new_P1_U5684 | ~new_P1_U3447;
  assign new_P1_U6072 = ~new_P1_R1360_U14 | ~new_P1_U3955 | ~new_P1_U3959;
  assign new_P1_U6073 = ~new_P1_U3985 | ~new_P1_U3055;
  assign new_P1_U6074 = ~new_P1_U3413 | ~new_P1_U4678;
  assign new_P1_U6075 = ~new_P1_U6074 | ~new_P1_U6073;
  assign new_P1_U6076 = ~new_P1_U3974 | ~new_P1_U3054;
  assign new_P1_U6077 = ~new_P1_U3411 | ~new_P1_U4659;
  assign new_P1_U6078 = ~new_P1_U6077 | ~new_P1_U6076;
  assign new_P1_U6079 = ~new_P1_U3975 | ~new_P1_U3053;
  assign new_P1_U6080 = ~new_P1_U3409 | ~new_P1_U4640;
  assign new_P1_U6081 = ~new_P1_U6080 | ~new_P1_U6079;
  assign new_P1_U6082 = ~new_P1_U3978 | ~new_P1_U3065;
  assign new_P1_U6083 = ~new_P1_U3403 | ~new_P1_U4583;
  assign new_P1_U6084 = ~new_P1_U6083 | ~new_P1_U6082;
  assign new_P1_U6085 = ~new_P1_U3979 | ~new_P1_U3066;
  assign new_P1_U6086 = ~new_P1_U3401 | ~new_P1_U4564;
  assign new_P1_U6087 = ~new_P1_U6086 | ~new_P1_U6085;
  assign new_P1_U6088 = ~new_P1_U3981 | ~new_P1_U3075;
  assign new_P1_U6089 = ~new_P1_U3397 | ~new_P1_U4526;
  assign new_P1_U6090 = ~new_P1_U6089 | ~new_P1_U6088;
  assign new_P1_U6091 = ~new_P1_U3980 | ~new_P1_U3061;
  assign new_P1_U6092 = ~new_P1_U3399 | ~new_P1_U4545;
  assign new_P1_U6093 = ~new_P1_U6092 | ~new_P1_U6091;
  assign new_P1_U6094 = ~new_P1_U3977 | ~new_P1_U3058;
  assign new_P1_U6095 = ~new_P1_U3405 | ~new_P1_U4602;
  assign new_P1_U6096 = ~new_P1_U6095 | ~new_P1_U6094;
  assign new_P1_U6097 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_U6098 = ~new_P1_U3407 | ~new_P1_U4621;
  assign new_P1_U6099 = ~new_P1_U6098 | ~new_P1_U6097;
  assign new_P1_U6100 = ~new_P1_U3984 | ~new_P1_U3059;
  assign new_P1_U6101 = ~new_P1_U3414 | ~new_P1_U4696;
  assign new_P1_U6102 = ~new_P1_U6101 | ~new_P1_U6100;
  assign new_P1_U6103 = ~new_P1_U3983 | ~new_P1_U3056;
  assign new_P1_U6104 = ~new_P1_U3415 | ~new_P1_U4716;
  assign new_P1_U6105 = ~new_P1_U6104 | ~new_P1_U6103;
  assign new_P1_U6106 = ~new_P1_U5838 | ~new_P1_U4450;
  assign new_P1_U6107 = ~new_P1_U3503 | ~new_P1_U3069;
  assign new_P1_U6108 = ~new_P1_U6107 | ~new_P1_U6106;
  assign new_P1_U6109 = ~new_P1_U5775 | ~new_P1_U4279;
  assign new_P1_U6110 = ~new_P1_U3476 | ~new_P1_U3084;
  assign new_P1_U6111 = ~new_P1_U6110 | ~new_P1_U6109;
  assign new_P1_U6112 = ~new_P1_U5782 | ~new_P1_U4298;
  assign new_P1_U6113 = ~new_P1_U3479 | ~new_P1_U3083;
  assign new_P1_U6114 = ~new_P1_U6113 | ~new_P1_U6112;
  assign new_P1_U6115 = ~new_P1_U5810 | ~new_P1_U4374;
  assign new_P1_U6116 = ~new_P1_U3491 | ~new_P1_U3080;
  assign new_P1_U6117 = ~new_P1_U6116 | ~new_P1_U6115;
  assign new_P1_U6118 = ~new_P1_U5817 | ~new_P1_U4393;
  assign new_P1_U6119 = ~new_P1_U3494 | ~new_P1_U3079;
  assign new_P1_U6120 = ~new_P1_U6119 | ~new_P1_U6118;
  assign new_P1_U6121 = ~new_P1_U5705 | ~new_P1_U4165;
  assign new_P1_U6122 = ~new_P1_U3450 | ~new_P1_U3077;
  assign new_P1_U6123 = ~new_P1_U6122 | ~new_P1_U6121;
  assign new_P1_U6124 = ~new_P1_U5726 | ~new_P1_U4141;
  assign new_P1_U6125 = ~new_P1_U3455 | ~new_P1_U3078;
  assign new_P1_U6126 = ~new_P1_U6125 | ~new_P1_U6124;
  assign new_P1_U6127 = ~new_P1_U5824 | ~new_P1_U4412;
  assign new_P1_U6128 = ~new_P1_U3497 | ~new_P1_U3074;
  assign new_P1_U6129 = ~new_P1_U6128 | ~new_P1_U6127;
  assign new_P1_U6130 = ~new_P1_U5831 | ~new_P1_U4431;
  assign new_P1_U6131 = ~new_P1_U3500 | ~new_P1_U3073;
  assign new_P1_U6132 = ~new_P1_U6131 | ~new_P1_U6130;
  assign new_P1_U6133 = ~new_P1_U5761 | ~new_P1_U4241;
  assign new_P1_U6134 = ~new_P1_U3470 | ~new_P1_U3071;
  assign new_P1_U6135 = ~new_P1_U6134 | ~new_P1_U6133;
  assign new_P1_U6136 = ~new_P1_U5768 | ~new_P1_U4260;
  assign new_P1_U6137 = ~new_P1_U3473 | ~new_P1_U3070;
  assign new_P1_U6138 = ~new_P1_U6137 | ~new_P1_U6136;
  assign new_P1_U6139 = ~new_P1_U5803 | ~new_P1_U4355;
  assign new_P1_U6140 = ~new_P1_U3488 | ~new_P1_U3072;
  assign new_P1_U6141 = ~new_P1_U6140 | ~new_P1_U6139;
  assign new_P1_U6142 = ~new_P1_U5733 | ~new_P1_U4160;
  assign new_P1_U6143 = ~new_P1_U3458 | ~new_P1_U3068;
  assign new_P1_U6144 = ~new_P1_U6143 | ~new_P1_U6142;
  assign new_P1_U6145 = ~new_P1_U5740 | ~new_P1_U4184;
  assign new_P1_U6146 = ~new_P1_U3461 | ~new_P1_U3064;
  assign new_P1_U6147 = ~new_P1_U6146 | ~new_P1_U6145;
  assign new_P1_U6148 = ~new_P1_U5754 | ~new_P1_U4222;
  assign new_P1_U6149 = ~new_P1_U3467 | ~new_P1_U3067;
  assign new_P1_U6150 = ~new_P1_U6149 | ~new_P1_U6148;
  assign new_P1_U6151 = ~new_P1_U5845 | ~new_P1_U4469;
  assign new_P1_U6152 = ~new_P1_U3506 | ~new_P1_U3082;
  assign new_P1_U6153 = ~new_P1_U6152 | ~new_P1_U6151;
  assign new_P1_U6154 = ~new_P1_U5850 | ~new_P1_U4488;
  assign new_P1_U6155 = ~new_P1_U3508 | ~new_P1_U3081;
  assign new_P1_U6156 = ~new_P1_U6155 | ~new_P1_U6154;
  assign new_P1_U6157 = ~new_P1_U5747 | ~new_P1_U4203;
  assign new_P1_U6158 = ~new_P1_U3464 | ~new_P1_U3060;
  assign new_P1_U6159 = ~new_P1_U6158 | ~new_P1_U6157;
  assign new_P1_U6160 = ~new_P1_U5796 | ~new_P1_U4336;
  assign new_P1_U6161 = ~new_P1_U3485 | ~new_P1_U3063;
  assign new_P1_U6162 = ~new_P1_U6161 | ~new_P1_U6160;
  assign new_P1_U6163 = ~new_P1_U5789 | ~new_P1_U4317;
  assign new_P1_U6164 = ~new_P1_U3482 | ~new_P1_U3062;
  assign new_P1_U6165 = ~new_P1_U6164 | ~new_P1_U6163;
  assign new_P1_U6166 = ~new_P1_U3982 | ~new_P1_U3076;
  assign new_P1_U6167 = ~new_P1_U3395 | ~new_P1_U4507;
  assign new_P1_U6168 = ~new_P1_U6167 | ~new_P1_U6166;
  assign new_P1_U6169 = ~new_P1_U5663 | ~new_P1_U3951;
  assign new_P1_U6170 = ~new_P1_U5086 | ~new_P1_U3426;
  assign new_P1_U6171 = ~new_P1_U3083 | ~new_P1_R1352_U6;
  assign new_P1_U6172 = ~new_P1_U3083 | ~new_P1_U3952;
  assign new_P1_U6173 = ~new_P1_U3084 | ~new_P1_R1352_U6;
  assign new_P1_U6174 = ~new_P1_U3084 | ~new_P1_U3952;
  assign new_P1_U6175 = ~new_P1_U3070 | ~new_P1_R1352_U6;
  assign new_P1_U6176 = ~new_P1_U3070 | ~new_P1_U3952;
  assign new_P1_U6177 = ~new_P1_U3071 | ~new_P1_R1352_U6;
  assign new_P1_U6178 = ~new_P1_U3071 | ~new_P1_U3952;
  assign new_P1_U6179 = ~new_P1_U3067 | ~new_P1_R1352_U6;
  assign new_P1_U6180 = ~new_P1_U3067 | ~new_P1_U3952;
  assign new_P1_U6181 = ~new_P1_U3060 | ~new_P1_R1352_U6;
  assign new_P1_U6182 = ~new_P1_U3060 | ~new_P1_U3952;
  assign new_P1_U6183 = ~new_P1_U3064 | ~new_P1_R1352_U6;
  assign new_P1_U6184 = ~new_P1_U3064 | ~new_P1_U3952;
  assign new_P1_U6185 = ~new_P1_R1309_U8 | ~new_P1_R1352_U6;
  assign new_P1_U6186 = ~new_P1_U3056 | ~new_P1_U3952;
  assign new_P1_U6187 = ~new_P1_R1309_U6 | ~new_P1_R1352_U6;
  assign new_P1_U6188 = ~new_P1_U3059 | ~new_P1_U3952;
  assign new_P1_U6189 = ~new_P1_U3068 | ~new_P1_R1352_U6;
  assign new_P1_U6190 = ~new_P1_U3068 | ~new_P1_U3952;
  assign new_P1_U6191 = ~new_P1_U3055 | ~new_P1_R1352_U6;
  assign new_P1_U6192 = ~new_P1_U3055 | ~new_P1_U3952;
  assign new_P1_U6193 = ~new_P1_U3054 | ~new_P1_R1352_U6;
  assign new_P1_U6194 = ~new_P1_U3054 | ~new_P1_U3952;
  assign new_P1_U6195 = ~new_P1_U3053 | ~new_P1_R1352_U6;
  assign new_P1_U6196 = ~new_P1_U3053 | ~new_P1_U3952;
  assign new_P1_U6197 = ~new_P1_U3057 | ~new_P1_R1352_U6;
  assign new_P1_U6198 = ~new_P1_U3057 | ~new_P1_U3952;
  assign new_P1_U6199 = ~new_P1_U3058 | ~new_P1_R1352_U6;
  assign new_P1_U6200 = ~new_P1_U3058 | ~new_P1_U3952;
  assign new_P1_U6201 = ~new_P1_U3065 | ~new_P1_R1352_U6;
  assign new_P1_U6202 = ~new_P1_U3065 | ~new_P1_U3952;
  assign new_P1_U6203 = ~new_P1_U3066 | ~new_P1_R1352_U6;
  assign new_P1_U6204 = ~new_P1_U3066 | ~new_P1_U3952;
  assign new_P1_U6205 = ~new_P1_U3061 | ~new_P1_R1352_U6;
  assign new_P1_U6206 = ~new_P1_U3061 | ~new_P1_U3952;
  assign new_P1_U6207 = ~new_P1_U3075 | ~new_P1_R1352_U6;
  assign new_P1_U6208 = ~new_P1_U3075 | ~new_P1_U3952;
  assign new_P1_U6209 = ~new_P1_U3076 | ~new_P1_R1352_U6;
  assign new_P1_U6210 = ~new_P1_U3076 | ~new_P1_U3952;
  assign new_P1_U6211 = ~new_P1_U3078 | ~new_P1_R1352_U6;
  assign new_P1_U6212 = ~new_P1_U3078 | ~new_P1_U3952;
  assign new_P1_U6213 = ~new_P1_U3081 | ~new_P1_R1352_U6;
  assign new_P1_U6214 = ~new_P1_U3081 | ~new_P1_U3952;
  assign new_P1_U6215 = ~new_P1_U3082 | ~new_P1_R1352_U6;
  assign new_P1_U6216 = ~new_P1_U3082 | ~new_P1_U3952;
  assign new_P1_U6217 = ~new_P1_U3069 | ~new_P1_R1352_U6;
  assign new_P1_U6218 = ~new_P1_U3069 | ~new_P1_U3952;
  assign new_P1_U6219 = ~new_P1_U3073 | ~new_P1_R1352_U6;
  assign new_P1_U6220 = ~new_P1_U3073 | ~new_P1_U3952;
  assign new_P1_U6221 = ~new_P1_U3074 | ~new_P1_R1352_U6;
  assign new_P1_U6222 = ~new_P1_U3074 | ~new_P1_U3952;
  assign new_P1_U6223 = ~new_P1_U3079 | ~new_P1_R1352_U6;
  assign new_P1_U6224 = ~new_P1_U3079 | ~new_P1_U3952;
  assign new_P1_U6225 = ~new_P1_U3080 | ~new_P1_R1352_U6;
  assign new_P1_U6226 = ~new_P1_U3080 | ~new_P1_U3952;
  assign new_P1_U6227 = ~new_P1_U3072 | ~new_P1_R1352_U6;
  assign new_P1_U6228 = ~new_P1_U3072 | ~new_P1_U3952;
  assign new_P1_U6229 = ~new_P1_U3063 | ~new_P1_R1352_U6;
  assign new_P1_U6230 = ~new_P1_U3063 | ~new_P1_U3952;
  assign new_P1_U6231 = ~new_P1_U3062 | ~new_P1_R1352_U6;
  assign new_P1_U6232 = ~new_P1_U3062 | ~new_P1_U3952;
  assign new_P1_U6233 = ~new_P1_U3077 | ~new_P1_R1352_U6;
  assign new_P1_U6234 = ~new_P1_U3077 | ~new_P1_U3952;
  assign new_P1_U6235 = ~new_P1_U3448 | ~new_P1_U5364;
  assign new_P1_U6236 = ~new_P1_U5696 | ~new_P1_U3015 | ~P1_REG2_REG_0_;
  assign new_P2_R1161_U489 = ~new_P2_U3079 | ~new_P2_R1161_U61;
  assign new_P2_R1161_U488 = ~new_P2_R1161_U254 | ~new_P2_R1161_U486;
  assign new_P2_R1161_U487 = ~new_P2_R1161_U165 | ~new_P2_R1161_U166;
  assign new_P2_R1161_U486 = ~new_P2_R1161_U485 | ~new_P2_R1161_U484;
  assign new_P2_R1161_U485 = ~new_P2_U3431 | ~new_P2_R1161_U72;
  assign new_P2_R1161_U484 = ~new_P2_U3078 | ~new_P2_R1161_U71;
  assign new_P2_R1161_U483 = ~new_P2_U3431 | ~new_P2_R1161_U72;
  assign new_P2_R1161_U482 = ~new_P2_U3078 | ~new_P2_R1161_U71;
  assign new_P2_R1161_U481 = ~new_P2_R1161_U258 | ~new_P2_R1161_U479;
  assign new_P2_R1161_U480 = ~new_P2_R1161_U163 | ~new_P2_R1161_U164;
  assign new_P2_R1161_U479 = ~new_P2_R1161_U478 | ~new_P2_R1161_U477;
  assign new_P2_R1161_U478 = ~new_P2_U3434 | ~new_P2_R1161_U74;
  assign new_P2_R1161_U477 = ~new_P2_U3073 | ~new_P2_R1161_U73;
  assign new_P2_R1161_U476 = ~new_P2_U3434 | ~new_P2_R1161_U74;
  assign new_P2_R1161_U475 = ~new_P2_U3073 | ~new_P2_R1161_U73;
  assign new_P2_R1161_U474 = ~new_P2_R1161_U472 | ~new_P2_R1161_U262;
  assign new_P2_R1161_U473 = ~new_P2_R1161_U361 | ~new_P2_R1161_U92;
  assign new_P2_R1161_U472 = ~new_P2_R1161_U471 | ~new_P2_R1161_U470;
  assign new_P2_R1161_U471 = ~new_P2_U3437 | ~new_P2_R1161_U57;
  assign new_P2_R1161_U470 = ~new_P2_U3072 | ~new_P2_R1161_U56;
  assign new_P2_R1161_U469 = ~new_P2_U3440 | ~new_P2_R1161_U58;
  assign new_P2_R1161_U468 = ~new_P2_U3068 | ~new_P2_R1161_U60;
  assign new_P2_R1161_U467 = ~new_P2_R1161_U270 | ~new_P2_R1161_U465;
  assign new_P2_R1161_U466 = ~new_P2_R1161_U360 | ~new_P2_R1161_U162;
  assign new_P2_U3013 = new_P2_U3380 & new_P2_U5446;
  assign new_P2_U3014 = new_P2_U3380 & new_P2_U3379;
  assign new_P2_U3015 = new_P2_U5449 & new_P2_U3379;
  assign new_P2_U3016 = new_P2_U5449 & new_P2_U5446;
  assign new_P2_U3017 = new_P2_U3870 & new_P2_U5443;
  assign new_P2_U3018 = new_P2_U3587 & new_P2_U3582;
  assign new_P2_U3019 = new_P2_U3381 & new_P2_U3382;
  assign new_P2_U3020 = new_P2_U5458 & new_P2_U3381;
  assign new_P2_U3021 = new_P2_U5455 & new_P2_U3382;
  assign new_P2_U3022 = new_P2_U5458 & new_P2_U5455;
  assign new_P2_U3023 = new_P2_U3046 & P2_STATE_REG;
  assign new_P2_U3024 = new_P2_U3701 & new_P2_U3366;
  assign new_P2_U3025 = new_P2_U3907 & new_P2_U4069;
  assign new_P2_U3026 = new_P2_U3015 & new_P2_U5443;
  assign new_P2_U3027 = new_P2_U3297 & P2_STATE_REG;
  assign new_P2_U3028 = new_P2_U3882 & new_P2_U3908;
  assign new_P2_U3029 = new_P2_U3908 & new_P2_U3365;
  assign new_P2_U3030 = new_P2_U3698 & new_P2_U3908;
  assign new_P2_U3031 = new_P2_U3886 & new_P2_U3023;
  assign new_P2_U3032 = new_P2_U3891 & new_P2_U4069;
  assign new_P2_U3033 = new_P2_U3907 & new_P2_U4085;
  assign new_P2_U3034 = new_P2_U3908 & new_P2_U3025;
  assign new_P2_U3035 = new_P2_U3023 & new_P2_U4985;
  assign new_P2_U3036 = new_P2_U3891 & new_P2_U4085;
  assign new_P2_U3037 = new_P2_U5464 & new_P2_U4750;
  assign new_P2_U3038 = new_P2_U3024 & new_P2_U5464;
  assign new_P2_U3039 = new_P2_U5461 & new_P2_U4750;
  assign new_P2_U3040 = new_P2_U3888 & new_P2_U4750;
  assign new_P2_U3041 = new_P2_U3024 & new_P2_U3888;
  assign new_P2_U3042 = new_P2_U3023 & new_P2_U3366;
  assign new_P2_U3043 = new_P2_U3023 & new_P2_U3365;
  assign new_P2_U3044 = new_P2_U5000 & P2_STATE_REG;
  assign new_P2_U3045 = new_P2_U3023 & new_P2_U5002;
  assign new_P2_U3046 = new_P2_U5436 & new_P2_U3362;
  assign new_P2_U3047 = new_P2_U3697 & new_P2_U3018;
  assign new_P2_U3048 = new_P2_U3696 & new_P2_U3018;
  assign new_P2_U3049 = new_P2_U4745 & new_P2_U4744;
  assign new_P2_U3050 = new_P2_U4755 & P2_STATE_REG;
  assign new_P2_U3051 = n2565 & new_P2_U4757;
  assign new_P2_U3052 = ~new_P2_U4531 | ~new_P2_U4532 | ~new_P2_U4534 | ~new_P2_U4533;
  assign new_P2_U3053 = ~new_P2_U4549 | ~new_P2_U4550 | ~new_P2_U4552 | ~new_P2_U4551;
  assign new_P2_U3054 = ~new_P2_U4567 | ~new_P2_U4568 | ~new_P2_U4570 | ~new_P2_U4569;
  assign new_P2_U3055 = ~new_P2_U4605 | ~new_P2_U4606 | ~new_P2_U4608 | ~new_P2_U4607;
  assign new_P2_U3056 = ~new_P2_U4513 | ~new_P2_U4514 | ~new_P2_U4516 | ~new_P2_U4515;
  assign new_P2_U3057 = ~new_P2_U4495 | ~new_P2_U4496 | ~new_P2_U4498 | ~new_P2_U4497;
  assign new_P2_U3058 = ~new_P2_U4585 | ~new_P2_U4586 | ~new_P2_U4588 | ~new_P2_U4587;
  assign new_P2_U3059 = ~new_P2_U4117 | ~new_P2_U4118 | ~new_P2_U4120 | ~new_P2_U4119;
  assign new_P2_U3060 = ~new_P2_U4441 | ~new_P2_U4442 | ~new_P2_U4444 | ~new_P2_U4443;
  assign new_P2_U3061 = ~new_P2_U4225 | ~new_P2_U4226 | ~new_P2_U4228 | ~new_P2_U4227;
  assign new_P2_U3062 = ~new_P2_U4243 | ~new_P2_U4244 | ~new_P2_U4246 | ~new_P2_U4245;
  assign new_P2_U3063 = ~new_P2_U4099 | ~new_P2_U4100 | ~new_P2_U4102 | ~new_P2_U4101;
  assign new_P2_U3064 = ~new_P2_U4477 | ~new_P2_U4478 | ~new_P2_U4480 | ~new_P2_U4479;
  assign new_P2_U3065 = ~new_P2_U4459 | ~new_P2_U4460 | ~new_P2_U4462 | ~new_P2_U4461;
  assign new_P2_U3066 = ~new_P2_U4135 | ~new_P2_U4136 | ~new_P2_U4138 | ~new_P2_U4137;
  assign new_P2_U3067 = ~new_P2_U4074 | ~new_P2_U4075 | ~new_P2_U4077 | ~new_P2_U4076;
  assign new_P2_U3068 = ~new_P2_U4351 | ~new_P2_U4352 | ~new_P2_U4354 | ~new_P2_U4353;
  assign new_P2_U3069 = ~new_P2_U4171 | ~new_P2_U4172 | ~new_P2_U4174 | ~new_P2_U4173;
  assign new_P2_U3070 = ~new_P2_U4153 | ~new_P2_U4154 | ~new_P2_U4156 | ~new_P2_U4155;
  assign new_P2_U3071 = ~new_P2_U4261 | ~new_P2_U4262 | ~new_P2_U4264 | ~new_P2_U4263;
  assign new_P2_U3072 = ~new_P2_U4333 | ~new_P2_U4334 | ~new_P2_U4336 | ~new_P2_U4335;
  assign new_P2_U3073 = ~new_P2_U4315 | ~new_P2_U4316 | ~new_P2_U4318 | ~new_P2_U4317;
  assign new_P2_U3074 = ~new_P2_U4423 | ~new_P2_U4424 | ~new_P2_U4426 | ~new_P2_U4425;
  assign new_P2_U3075 = ~new_P2_U4405 | ~new_P2_U4406 | ~new_P2_U4408 | ~new_P2_U4407;
  assign new_P2_U3076 = ~new_P2_U4079 | ~new_P2_U4080 | ~new_P2_U4082 | ~new_P2_U4081;
  assign new_P2_U3077 = ~new_P2_U4055 | ~new_P2_U4056 | ~new_P2_U4058 | ~new_P2_U4057;
  assign new_P2_U3078 = ~new_P2_U4297 | ~new_P2_U4298 | ~new_P2_U4300 | ~new_P2_U4299;
  assign new_P2_U3079 = ~new_P2_U4279 | ~new_P2_U4280 | ~new_P2_U4282 | ~new_P2_U4281;
  assign new_P2_U3080 = ~new_P2_U4387 | ~new_P2_U4388 | ~new_P2_U4390 | ~new_P2_U4389;
  assign new_P2_U3081 = ~new_P2_U4369 | ~new_P2_U4370 | ~new_P2_U4372 | ~new_P2_U4371;
  assign new_P2_U3082 = ~new_P2_U4207 | ~new_P2_U4208 | ~new_P2_U4210 | ~new_P2_U4209;
  assign new_P2_U3083 = ~new_P2_U4189 | ~new_P2_U4190 | ~new_P2_U4192 | ~new_P2_U4191;
  assign new_P2_U3084 = ~new_P2_U5337 | ~new_P2_U5336;
  assign new_P2_U3085 = ~new_P2_U5339 | ~new_P2_U5338;
  assign new_P2_U3086 = ~new_P2_U5344 | ~new_P2_U5345 | ~new_P2_U5343;
  assign new_P2_U3087 = ~new_P2_U5347 | ~new_P2_U5348 | ~new_P2_U5346;
  assign new_P2_U3088 = ~new_P2_U5350 | ~new_P2_U5351 | ~new_P2_U5349;
  assign new_P2_U3089 = ~new_P2_U5353 | ~new_P2_U5354 | ~new_P2_U5352;
  assign new_P2_U3090 = ~new_P2_U5356 | ~new_P2_U5357 | ~new_P2_U5355;
  assign new_P2_U3091 = ~new_P2_U5359 | ~new_P2_U5360 | ~new_P2_U5358;
  assign new_P2_U3092 = ~new_P2_U5362 | ~new_P2_U5363 | ~new_P2_U5361;
  assign new_P2_U3093 = ~new_P2_U5365 | ~new_P2_U5366 | ~new_P2_U5364;
  assign new_P2_U3094 = ~new_P2_U5368 | ~new_P2_U5369 | ~new_P2_U5367;
  assign new_P2_U3095 = ~new_P2_U5371 | ~new_P2_U5372 | ~new_P2_U5370;
  assign new_P2_U3096 = ~new_P2_U5376 | ~new_P2_U5377 | ~new_P2_U5378;
  assign new_P2_U3097 = ~new_P2_U5379 | ~new_P2_U5380 | ~new_P2_U5381;
  assign new_P2_U3098 = ~new_P2_U5382 | ~new_P2_U5383 | ~new_P2_U5384;
  assign new_P2_U3099 = ~new_P2_U5385 | ~new_P2_U5386 | ~new_P2_U5387;
  assign new_P2_U3100 = ~new_P2_U5388 | ~new_P2_U5389 | ~new_P2_U5390;
  assign new_P2_U3101 = ~new_P2_U5391 | ~new_P2_U5392 | ~new_P2_U5393;
  assign new_P2_U3102 = ~new_P2_U5394 | ~new_P2_U5395 | ~new_P2_U5396;
  assign new_P2_U3103 = ~new_P2_U5397 | ~new_P2_U5398 | ~new_P2_U5399;
  assign new_P2_U3104 = ~new_P2_U5400 | ~new_P2_U5401 | ~new_P2_U5402;
  assign new_P2_U3105 = ~new_P2_U5403 | ~new_P2_U5404 | ~new_P2_U5405;
  assign new_P2_U3106 = ~new_P2_U5318 | ~new_P2_U5319 | ~new_P2_U5320;
  assign new_P2_U3107 = ~new_P2_U5321 | ~new_P2_U5322 | ~new_P2_U5323;
  assign new_P2_U3108 = ~new_P2_U5324 | ~new_P2_U5325 | ~new_P2_U5326;
  assign new_P2_U3109 = ~new_P2_U5327 | ~new_P2_U5328 | ~new_P2_U5329;
  assign new_P2_U3110 = ~new_P2_U5330 | ~new_P2_U5331 | ~new_P2_U5332;
  assign new_P2_U3111 = ~new_P2_U5335 | ~new_P2_U5334 | ~new_P2_U5333;
  assign new_P2_U3112 = ~new_P2_U5342 | ~new_P2_U5341 | ~new_P2_U5340;
  assign new_P2_U3113 = ~new_P2_U5375 | ~new_P2_U5374 | ~new_P2_U5373;
  assign new_P2_U3114 = ~new_P2_U5408 | ~new_P2_U5407 | ~new_P2_U5406;
  assign new_P2_U3115 = ~new_P2_U5410 | ~new_P2_U5409;
  assign new_P2_U3116 = ~new_P2_U5267 | ~new_P2_U5266;
  assign new_P2_U3117 = ~new_P2_U5269 | ~new_P2_U5268;
  assign new_P2_U3118 = ~new_P2_U5272 | ~new_P2_U5273 | ~new_P2_U3375;
  assign new_P2_U3119 = ~new_P2_U5274 | ~new_P2_U5275 | ~new_P2_U3375;
  assign new_P2_U3120 = ~new_P2_U5276 | ~new_P2_U5277 | ~new_P2_U3375;
  assign new_P2_U3121 = ~new_P2_U5278 | ~new_P2_U5279 | ~new_P2_U3375;
  assign new_P2_U3122 = ~new_P2_U5280 | ~new_P2_U5281 | ~new_P2_U3375;
  assign new_P2_U3123 = ~new_P2_U5282 | ~new_P2_U5283 | ~new_P2_U3375;
  assign new_P2_U3124 = ~new_P2_U5284 | ~new_P2_U5285 | ~new_P2_U3375;
  assign new_P2_U3125 = ~new_P2_U5286 | ~new_P2_U5287 | ~new_P2_U3375;
  assign new_P2_U3126 = ~new_P2_U5288 | ~new_P2_U5289 | ~new_P2_U3375;
  assign new_P2_U3127 = ~new_P2_U5290 | ~new_P2_U5291 | ~new_P2_U3375;
  assign new_P2_U3128 = ~new_P2_U5294 | ~new_P2_U5295 | ~new_P2_U3375;
  assign new_P2_U3129 = ~new_P2_U5296 | ~new_P2_U5297 | ~new_P2_U3375;
  assign new_P2_U3130 = ~new_P2_U5298 | ~new_P2_U5299 | ~new_P2_U3375;
  assign new_P2_U3131 = ~new_P2_U5300 | ~new_P2_U5301 | ~new_P2_U3375;
  assign new_P2_U3132 = ~new_P2_U5302 | ~new_P2_U5303 | ~new_P2_U3375;
  assign new_P2_U3133 = ~new_P2_U5304 | ~new_P2_U5305 | ~new_P2_U3375;
  assign new_P2_U3134 = ~new_P2_U5306 | ~new_P2_U5307 | ~new_P2_U3375;
  assign new_P2_U3135 = ~new_P2_U5308 | ~new_P2_U5309 | ~new_P2_U3375;
  assign new_P2_U3136 = ~new_P2_U5310 | ~new_P2_U5311 | ~new_P2_U3375;
  assign new_P2_U3137 = ~new_P2_U5312 | ~new_P2_U5313 | ~new_P2_U3375;
  assign new_P2_U3138 = ~new_P2_U5254 | ~new_P2_U5255 | ~new_P2_U3375;
  assign new_P2_U3139 = ~new_P2_U5256 | ~new_P2_U5257 | ~new_P2_U3375;
  assign new_P2_U3140 = ~new_P2_U5258 | ~new_P2_U5259 | ~new_P2_U3375;
  assign new_P2_U3141 = ~new_P2_U5260 | ~new_P2_U5261 | ~new_P2_U3375;
  assign new_P2_U3142 = ~new_P2_U5262 | ~new_P2_U5263 | ~new_P2_U3375;
  assign new_P2_U3143 = ~new_P2_U3822 | ~new_P2_U5265;
  assign new_P2_U3144 = ~new_P2_U3823 | ~new_P2_U5271;
  assign new_P2_U3145 = ~new_P2_U3824 | ~new_P2_U5293;
  assign new_P2_U3146 = ~new_P2_U3825 | ~new_P2_U5315;
  assign new_P2_U3147 = ~new_P2_U3826 | ~new_P2_U5317;
  assign new_P2_U3148 = ~new_P2_U3375 | ~new_P2_U3385 | ~new_P2_U5449;
  assign new_P2_U3149 = ~new_P2_U3818 | ~new_P2_U3013;
  assign n2560 = ~new_P2_U3817 | ~new_P2_U5249;
  assign n2555 = ~P2_STATE_REG;
  assign new_P2_U3152 = ~new_P2_U3359 | ~new_P2_U5940 | ~new_P2_U5939;
  assign n2550 = ~new_P2_U5246 | ~new_P2_U3816 | ~new_P2_U5245 | ~new_P2_U5244;
  assign n2545 = ~new_P2_U5237 | ~new_P2_U5235 | ~new_P2_U5236 | ~new_P2_U3815;
  assign n2540 = ~new_P2_U5228 | ~new_P2_U3814 | ~new_P2_U5227 | ~new_P2_U5226;
  assign n2535 = ~new_P2_U5219 | ~new_P2_U5217 | ~new_P2_U5218 | ~new_P2_U3813;
  assign n2530 = ~new_P2_U5210 | ~new_P2_U3812 | ~new_P2_U5209 | ~new_P2_U5208;
  assign n2525 = ~new_P2_U3811 | ~new_P2_U3810 | ~new_P2_U5200;
  assign n2520 = ~new_P2_U5192 | ~new_P2_U5190 | ~new_P2_U5191 | ~new_P2_U3809;
  assign n2515 = ~new_P2_U5183 | ~new_P2_U5181 | ~new_P2_U5182 | ~new_P2_U3808;
  assign n2510 = ~new_P2_U5174 | ~new_P2_U3807 | ~new_P2_U5173 | ~new_P2_U5172;
  assign n2505 = ~new_P2_U3806 | ~new_P2_U3805 | ~new_P2_U5164;
  assign n2500 = ~new_P2_U5156 | ~new_P2_U5154 | ~new_P2_U5155 | ~new_P2_U3804;
  assign n2495 = ~new_P2_U5147 | ~new_P2_U3803 | ~new_P2_U5146 | ~new_P2_U5145;
  assign n2490 = ~new_P2_U5138 | ~new_P2_U5136 | ~new_P2_U5137 | ~new_P2_U3802;
  assign n2485 = ~new_P2_U5129 | ~new_P2_U3801 | ~new_P2_U5128 | ~new_P2_U5127;
  assign n2480 = ~new_P2_U5120 | ~new_P2_U3800 | ~new_P2_U5119 | ~new_P2_U5118;
  assign n2475 = ~new_P2_U5111 | ~new_P2_U3799 | ~new_P2_U5110 | ~new_P2_U5109;
  assign n2470 = ~new_P2_U5102 | ~new_P2_U5100 | ~new_P2_U5101 | ~new_P2_U3798;
  assign n2465 = ~new_P2_U3797 | ~new_P2_U3796 | ~new_P2_U5092;
  assign n2460 = ~new_P2_U5084 | ~new_P2_U3795 | ~new_P2_U5083 | ~new_P2_U5082;
  assign n2455 = ~new_P2_U5075 | ~new_P2_U3794;
  assign n2450 = ~new_P2_U5068 | ~new_P2_U5066 | ~new_P2_U5067 | ~new_P2_U3791;
  assign n2445 = ~new_P2_U5059 | ~new_P2_U3790 | ~new_P2_U5058 | ~new_P2_U5057;
  assign n2440 = ~new_P2_U5050 | ~new_P2_U5048 | ~new_P2_U5049 | ~new_P2_U3789;
  assign n2435 = ~new_P2_U5041 | ~new_P2_U3788 | ~new_P2_U5040 | ~new_P2_U5039;
  assign n2430 = ~new_P2_U3787 | ~new_P2_U3786 | ~new_P2_U5031;
  assign n2425 = ~new_P2_U5023 | ~new_P2_U3785 | ~new_P2_U5022 | ~new_P2_U5021;
  assign n2420 = ~new_P2_U5014 | ~new_P2_U3784 | ~new_P2_U5013 | ~new_P2_U5012;
  assign n2415 = ~new_P2_U5005 | ~new_P2_U5003 | ~new_P2_U5004 | ~new_P2_U3783;
  assign n2410 = ~new_P2_U4992 | ~new_P2_U3782 | ~new_P2_U4991 | ~new_P2_U4990;
  assign n2240 = ~new_P2_U4969 | ~new_P2_U3761;
  assign n2235 = ~new_P2_U4958 | ~new_P2_U3758;
  assign n2230 = ~new_P2_U4947 | ~new_P2_U3755;
  assign n2225 = ~new_P2_U3752 | ~new_P2_U4937 | ~new_P2_U4936;
  assign n2220 = ~new_P2_U3749 | ~new_P2_U4926 | ~new_P2_U4925;
  assign n2215 = ~new_P2_U4912 | ~new_P2_U3748 | ~new_P2_U4914 | ~new_P2_U3746;
  assign n2210 = ~new_P2_U4901 | ~new_P2_U4903 | ~new_P2_U3743;
  assign n2205 = ~new_P2_U3740 | ~new_P2_U3741 | ~new_P2_U4892;
  assign n2200 = ~new_P2_U3737 | ~new_P2_U3738 | ~new_P2_U4881;
  assign n2195 = ~new_P2_U4870 | ~new_P2_U3734;
  assign n2190 = ~new_P2_U4859 | ~new_P2_U3731;
  assign n2185 = ~new_P2_U4848 | ~new_P2_U3728;
  assign n2180 = ~new_P2_U4837 | ~new_P2_U3725;
  assign n2175 = ~new_P2_U4826 | ~new_P2_U3722;
  assign n2170 = ~new_P2_U4815 | ~new_P2_U3719;
  assign n2165 = ~new_P2_U4804 | ~new_P2_U3716;
  assign n2160 = ~new_P2_U4793 | ~new_P2_U3713;
  assign n2155 = ~new_P2_U4782 | ~new_P2_U3710;
  assign n2150 = ~new_P2_U4771 | ~new_P2_U3707;
  assign n2145 = ~new_P2_U4760 | ~new_P2_U3704;
  assign n2140 = ~new_P2_U4748 | ~new_P2_U4749 | ~new_P2_U3049;
  assign n2135 = ~new_P2_U4746 | ~new_P2_U4747 | ~new_P2_U3049;
  assign n2130 = ~new_P2_U3862 | ~new_P2_U4741 | ~new_P2_U4742 | ~new_P2_U4743;
  assign n2125 = ~new_P2_U3861 | ~new_P2_U4738 | ~new_P2_U4740 | ~new_P2_U4739 | ~new_P2_U4737;
  assign n2120 = ~new_P2_U3860 | ~new_P2_U4734 | ~new_P2_U4736 | ~new_P2_U4735 | ~new_P2_U4733;
  assign n2115 = ~new_P2_U3859 | ~new_P2_U4730 | ~new_P2_U4732 | ~new_P2_U4731 | ~new_P2_U4729;
  assign n2110 = ~new_P2_U3858 | ~new_P2_U4726 | ~new_P2_U4728 | ~new_P2_U4727 | ~new_P2_U4725;
  assign n2105 = ~new_P2_U3857 | ~new_P2_U4722 | ~new_P2_U4724 | ~new_P2_U4723 | ~new_P2_U4721;
  assign n2100 = ~new_P2_U3856 | ~new_P2_U4718 | ~new_P2_U4720 | ~new_P2_U4719 | ~new_P2_U4717;
  assign n2095 = ~new_P2_U3855 | ~new_P2_U4714 | ~new_P2_U4716 | ~new_P2_U4715 | ~new_P2_U4713;
  assign n2090 = ~new_P2_U3854 | ~new_P2_U4710 | ~new_P2_U4712 | ~new_P2_U4711 | ~new_P2_U4709;
  assign n2085 = ~new_P2_U3853 | ~new_P2_U4706 | ~new_P2_U4708 | ~new_P2_U4707 | ~new_P2_U4705;
  assign n2080 = ~new_P2_U3852 | ~new_P2_U4702 | ~new_P2_U4704 | ~new_P2_U4703 | ~new_P2_U4701;
  assign n2075 = ~new_P2_U3851 | ~new_P2_U4698 | ~new_P2_U4700 | ~new_P2_U4699 | ~new_P2_U4697;
  assign n2070 = ~new_P2_U3850 | ~new_P2_U4694 | ~new_P2_U4696 | ~new_P2_U4695 | ~new_P2_U4693;
  assign n2065 = ~new_P2_U3849 | ~new_P2_U4690 | ~new_P2_U4692 | ~new_P2_U4691 | ~new_P2_U4689;
  assign n2060 = ~new_P2_U3848 | ~new_P2_U4686 | ~new_P2_U4688 | ~new_P2_U4687 | ~new_P2_U4685;
  assign n2055 = ~new_P2_U3847 | ~new_P2_U4682 | ~new_P2_U4684 | ~new_P2_U4683 | ~new_P2_U4681;
  assign n2050 = ~new_P2_U3846 | ~new_P2_U4678 | ~new_P2_U4680 | ~new_P2_U4679 | ~new_P2_U4677;
  assign n2045 = ~new_P2_U3845 | ~new_P2_U4674 | ~new_P2_U4676 | ~new_P2_U4675 | ~new_P2_U4673;
  assign n2040 = ~new_P2_U3844 | ~new_P2_U4670 | ~new_P2_U4672 | ~new_P2_U4671 | ~new_P2_U4669;
  assign n2035 = ~new_P2_U3843 | ~new_P2_U4666 | ~new_P2_U4668 | ~new_P2_U4667 | ~new_P2_U4665;
  assign n2030 = ~new_P2_U3842 | ~new_P2_U4662 | ~new_P2_U4664 | ~new_P2_U4663 | ~new_P2_U4661;
  assign n2025 = ~new_P2_U3841 | ~new_P2_U4657 | ~new_P2_U4658 | ~new_P2_U4660 | ~new_P2_U4659;
  assign n2020 = ~new_P2_U3840 | ~new_P2_U4653 | ~new_P2_U4654 | ~new_P2_U4656 | ~new_P2_U4655;
  assign n2015 = ~new_P2_U4652 | ~new_P2_U3839 | ~new_P2_U4651 | ~new_P2_U4650 | ~new_P2_U4649;
  assign n2010 = ~new_P2_U4648 | ~new_P2_U3838 | ~new_P2_U4647 | ~new_P2_U4646 | ~new_P2_U4645;
  assign n2005 = ~new_P2_U4644 | ~new_P2_U3837 | ~new_P2_U4643 | ~new_P2_U4642 | ~new_P2_U4641;
  assign n2000 = ~new_P2_U4640 | ~new_P2_U3836 | ~new_P2_U4639 | ~new_P2_U4638 | ~new_P2_U4637;
  assign n1995 = ~new_P2_U4636 | ~new_P2_U3835 | ~new_P2_U4635 | ~new_P2_U4634 | ~new_P2_U4633;
  assign n1990 = ~new_P2_U4632 | ~new_P2_U3834 | ~new_P2_U4631 | ~new_P2_U4630 | ~new_P2_U4629;
  assign n1985 = ~new_P2_U4628 | ~new_P2_U3833 | ~new_P2_U4627 | ~new_P2_U4626 | ~new_P2_U4625;
  assign n1660 = P2_D_REG_31_ & new_P2_U3828;
  assign n1655 = P2_D_REG_30_ & new_P2_U3828;
  assign n1650 = P2_D_REG_29_ & new_P2_U3828;
  assign n1645 = P2_D_REG_28_ & new_P2_U3828;
  assign n1640 = P2_D_REG_27_ & new_P2_U3828;
  assign n1635 = P2_D_REG_26_ & new_P2_U3828;
  assign n1630 = P2_D_REG_25_ & new_P2_U3828;
  assign n1625 = P2_D_REG_24_ & new_P2_U3828;
  assign n1620 = P2_D_REG_23_ & new_P2_U3828;
  assign n1615 = P2_D_REG_22_ & new_P2_U3828;
  assign n1610 = P2_D_REG_21_ & new_P2_U3828;
  assign n1605 = P2_D_REG_20_ & new_P2_U3828;
  assign n1600 = P2_D_REG_19_ & new_P2_U3828;
  assign n1595 = P2_D_REG_18_ & new_P2_U3828;
  assign n1590 = P2_D_REG_17_ & new_P2_U3828;
  assign n1585 = P2_D_REG_16_ & new_P2_U3828;
  assign n1580 = P2_D_REG_15_ & new_P2_U3828;
  assign n1575 = P2_D_REG_14_ & new_P2_U3828;
  assign n1570 = P2_D_REG_13_ & new_P2_U3828;
  assign n1565 = P2_D_REG_12_ & new_P2_U3828;
  assign n1560 = P2_D_REG_11_ & new_P2_U3828;
  assign n1555 = P2_D_REG_10_ & new_P2_U3828;
  assign n1550 = P2_D_REG_9_ & new_P2_U3828;
  assign n1545 = P2_D_REG_8_ & new_P2_U3828;
  assign n1540 = P2_D_REG_7_ & new_P2_U3828;
  assign n1535 = P2_D_REG_6_ & new_P2_U3828;
  assign n1530 = P2_D_REG_5_ & new_P2_U3828;
  assign n1525 = P2_D_REG_4_ & new_P2_U3828;
  assign n1520 = P2_D_REG_3_ & new_P2_U3828;
  assign n1515 = P2_D_REG_2_ & new_P2_U3828;
  assign n1500 = ~new_P2_U4011 | ~new_P2_U4012 | ~new_P2_U4013;
  assign n1495 = ~new_P2_U4008 | ~new_P2_U4009 | ~new_P2_U4010;
  assign n1490 = ~new_P2_U4005 | ~new_P2_U4006 | ~new_P2_U4007;
  assign n1485 = ~new_P2_U4002 | ~new_P2_U4003 | ~new_P2_U4004;
  assign n1480 = ~new_P2_U3999 | ~new_P2_U4000 | ~new_P2_U4001;
  assign n1475 = ~new_P2_U3996 | ~new_P2_U3997 | ~new_P2_U3998;
  assign n1470 = ~new_P2_U3993 | ~new_P2_U3994 | ~new_P2_U3995;
  assign n1465 = ~new_P2_U3990 | ~new_P2_U3991 | ~new_P2_U3992;
  assign n1460 = ~new_P2_U3987 | ~new_P2_U3988 | ~new_P2_U3989;
  assign n1455 = ~new_P2_U3984 | ~new_P2_U3985 | ~new_P2_U3986;
  assign n1450 = ~new_P2_U3981 | ~new_P2_U3982 | ~new_P2_U3983;
  assign n1445 = ~new_P2_U3978 | ~new_P2_U3979 | ~new_P2_U3980;
  assign n1440 = ~new_P2_U3975 | ~new_P2_U3976 | ~new_P2_U3977;
  assign n1435 = ~new_P2_U3972 | ~new_P2_U3973 | ~new_P2_U3974;
  assign n1430 = ~new_P2_U3969 | ~new_P2_U3970 | ~new_P2_U3971;
  assign n1425 = ~new_P2_U3966 | ~new_P2_U3967 | ~new_P2_U3968;
  assign n1420 = ~new_P2_U3963 | ~new_P2_U3964 | ~new_P2_U3965;
  assign n1415 = ~new_P2_U3960 | ~new_P2_U3961 | ~new_P2_U3962;
  assign n1410 = ~new_P2_U3957 | ~new_P2_U3958 | ~new_P2_U3959;
  assign n1405 = ~new_P2_U3954 | ~new_P2_U3955 | ~new_P2_U3956;
  assign n1400 = ~new_P2_U3951 | ~new_P2_U3952 | ~new_P2_U3953;
  assign n1395 = ~new_P2_U3948 | ~new_P2_U3949 | ~new_P2_U3950;
  assign n1390 = ~new_P2_U3945 | ~new_P2_U3946 | ~new_P2_U3947;
  assign n1385 = ~new_P2_U3942 | ~new_P2_U3943 | ~new_P2_U3944;
  assign n1380 = ~new_P2_U3939 | ~new_P2_U3940 | ~new_P2_U3941;
  assign n1375 = ~new_P2_U3936 | ~new_P2_U3937 | ~new_P2_U3938;
  assign n1370 = ~new_P2_U3933 | ~new_P2_U3934 | ~new_P2_U3935;
  assign n1365 = ~new_P2_U3930 | ~new_P2_U3931 | ~new_P2_U3932;
  assign n1360 = ~new_P2_U3927 | ~new_P2_U3928 | ~new_P2_U3929;
  assign n1355 = ~new_P2_U3924 | ~new_P2_U3925 | ~new_P2_U3926;
  assign n1350 = ~new_P2_U3921 | ~new_P2_U3922 | ~new_P2_U3923;
  assign n1345 = ~new_P2_U3918 | ~new_P2_U3919 | ~new_P2_U3920;
  assign n2405 = new_P2_U3780 & new_P2_U5417;
  assign new_P2_U3297 = ~P2_STATE_REG | ~new_P2_U3827;
  assign new_P2_U3298 = ~P2_B_REG;
  assign new_P2_U3299 = ~new_P2_U3374 | ~new_P2_U5427;
  assign new_P2_U3300 = ~new_P2_U3374 | ~new_P2_U4014;
  assign new_P2_U3301 = ~new_P2_U3013 | ~new_P2_U5443;
  assign new_P2_U3302 = ~new_P2_U3014 | ~new_P2_U5452;
  assign new_P2_U3303 = ~new_P2_U3588 | ~new_P2_U3018;
  assign new_P2_U3304 = ~new_P2_U3589 | ~new_P2_U3018;
  assign new_P2_U3305 = ~new_P2_U3014 | ~new_P2_U5443;
  assign new_P2_U3306 = ~new_P2_U3014 | ~new_P2_U3378;
  assign new_P2_U3307 = ~new_P2_U3013 | ~new_P2_U3378;
  assign new_P2_U3308 = ~new_P2_U3378 | ~new_P2_U3385 | ~new_P2_U3379;
  assign new_P2_U3309 = ~new_P2_U3378 | ~new_P2_U5446 | ~new_P2_U3385;
  assign new_P2_U3310 = ~new_P2_U5452 | ~new_P2_U3013;
  assign new_P2_U3311 = ~new_P2_U3874 | ~new_P2_U5443;
  assign new_P2_U3312 = ~new_P2_U3016 | ~new_P2_U3385;
  assign new_P2_U3313 = ~new_P2_U3385 | ~new_P2_U3380;
  assign new_P2_U3314 = ~new_P2_U3575 | ~new_P2_U3576 | ~new_P2_U4067 | ~new_P2_U4066 | ~new_P2_U4065;
  assign new_P2_U3315 = ~new_P2_U3592 | ~new_P2_U3590 | ~new_P2_U4087 | ~new_P2_U4086;
  assign new_P2_U3316 = ~new_P2_U3596 | ~new_P2_U3594 | ~new_P2_U4105 | ~new_P2_U4104;
  assign new_P2_U3317 = ~new_P2_U3600 | ~new_P2_U3598 | ~new_P2_U4123 | ~new_P2_U4122;
  assign new_P2_U3318 = ~new_P2_U3604 | ~new_P2_U3602 | ~new_P2_U4141 | ~new_P2_U4140;
  assign new_P2_U3319 = ~new_P2_U3608 | ~new_P2_U3606 | ~new_P2_U4159 | ~new_P2_U4158;
  assign new_P2_U3320 = ~new_P2_U3612 | ~new_P2_U3610 | ~new_P2_U4177 | ~new_P2_U4176;
  assign new_P2_U3321 = ~new_P2_U3616 | ~new_P2_U3614 | ~new_P2_U4195 | ~new_P2_U4194;
  assign new_P2_U3322 = ~new_P2_U3619 | ~new_P2_U4215 | ~new_P2_U4214 | ~new_P2_U4213 | ~new_P2_U4212;
  assign new_P2_U3323 = ~new_P2_U3622 | ~new_P2_U4233 | ~new_P2_U4232 | ~new_P2_U4231 | ~new_P2_U4230;
  assign new_P2_U3324 = ~new_P2_U3625 | ~new_P2_U4251 | ~new_P2_U4250 | ~new_P2_U4249 | ~new_P2_U4248;
  assign new_P2_U3325 = ~new_P2_U3628 | ~new_P2_U4269 | ~new_P2_U4268 | ~new_P2_U4267 | ~new_P2_U4266;
  assign new_P2_U3326 = ~new_P2_U3632 | ~new_P2_U3630 | ~new_P2_U4285 | ~new_P2_U4284;
  assign new_P2_U3327 = ~new_P2_U3636 | ~new_P2_U3634 | ~new_P2_U4303 | ~new_P2_U4302;
  assign new_P2_U3328 = ~new_P2_U3639 | ~new_P2_U4323 | ~new_P2_U4322 | ~new_P2_U4321 | ~new_P2_U4320;
  assign new_P2_U3329 = ~new_P2_U3642 | ~new_P2_U4341 | ~new_P2_U4340 | ~new_P2_U4339 | ~new_P2_U4338;
  assign new_P2_U3330 = ~new_P2_U3645 | ~new_P2_U4359 | ~new_P2_U4358 | ~new_P2_U4357 | ~new_P2_U4356;
  assign new_P2_U3331 = ~new_P2_U3649 | ~new_P2_U3647 | ~new_P2_U4375 | ~new_P2_U4374;
  assign new_P2_U3332 = ~new_P2_U3653 | ~new_P2_U3651 | ~new_P2_U4393 | ~new_P2_U4392;
  assign new_P2_U3333 = ~new_P2_U3657 | ~new_P2_U3655 | ~new_P2_U4411 | ~new_P2_U4410;
  assign new_P2_U3334 = ~new_U44 | ~new_P2_U3829;
  assign new_P2_U3335 = ~new_P2_U3661 | ~new_P2_U3659 | ~new_P2_U4429 | ~new_P2_U4428;
  assign new_P2_U3336 = ~new_U43 | ~new_P2_U3829;
  assign new_P2_U3337 = ~new_P2_U3664 | ~new_P2_U4449 | ~new_P2_U4448 | ~new_P2_U4447 | ~new_P2_U4446;
  assign new_P2_U3338 = ~new_U42 | ~new_P2_U3829;
  assign new_P2_U3339 = ~new_P2_U3667 | ~new_P2_U4467 | ~new_P2_U4466 | ~new_P2_U4465 | ~new_P2_U4464;
  assign new_P2_U3340 = ~new_U41 | ~new_P2_U3829;
  assign new_P2_U3341 = ~new_P2_U3670 | ~new_P2_U4485 | ~new_P2_U4484 | ~new_P2_U4483 | ~new_P2_U4482;
  assign new_P2_U3342 = ~new_U40 | ~new_P2_U3829;
  assign new_P2_U3343 = ~new_P2_U3674 | ~new_P2_U3672 | ~new_P2_U4501 | ~new_P2_U4500;
  assign new_P2_U3344 = ~new_U39 | ~new_P2_U3829;
  assign new_P2_U3345 = ~new_P2_U3678 | ~new_P2_U3676 | ~new_P2_U4519 | ~new_P2_U4518;
  assign new_P2_U3346 = ~new_U38 | ~new_P2_U3829;
  assign new_P2_U3347 = ~new_P2_U3682 | ~new_P2_U3680 | ~new_P2_U4537 | ~new_P2_U4536;
  assign new_P2_U3348 = ~new_U37 | ~new_P2_U3829;
  assign new_P2_U3349 = ~new_P2_U3686 | ~new_P2_U3684 | ~new_P2_U4555 | ~new_P2_U4554;
  assign new_P2_U3350 = ~new_U36 | ~new_P2_U3829;
  assign new_P2_U3351 = ~new_P2_U3690 | ~new_P2_U3688 | ~new_P2_U4573 | ~new_P2_U4572;
  assign new_P2_U3352 = ~new_P2_U3383 | ~new_P2_U3384;
  assign new_P2_U3353 = ~new_U35 | ~new_P2_U3829;
  assign new_P2_U3354 = ~new_P2_U3694 | ~new_P2_U3692;
  assign new_P2_U3355 = ~new_U33 | ~new_P2_U3829;
  assign new_P2_U3356 = ~new_U32 | ~new_P2_U3829;
  assign new_P2_U3357 = ~new_P2_U3015 | ~new_P2_U5452;
  assign new_P2_U3358 = ~new_P2_U3023 | ~new_P2_U4623;
  assign new_P2_U3359 = ~new_P2_U5443 | ~new_P2_U3385;
  assign new_P2_U3360 = ~new_P2_U3875 | ~new_P2_U5443;
  assign new_P2_U3361 = ~new_P2_U3055 | ~new_P2_U3907 | ~new_P2_U4591;
  assign new_P2_U3362 = ~new_P2_U3372 | ~new_P2_U3373 | ~new_P2_U3374;
  assign new_P2_U3363 = ~new_P2_U3699 | ~new_P2_U3906;
  assign new_P2_U3364 = ~new_P2_U3313 | ~new_P2_U3829;
  assign new_P2_U3365 = ~new_P2_U3873 | ~new_P2_U5419;
  assign new_P2_U3366 = ~new_P2_U3700 | ~new_P2_U3050;
  assign new_P2_U3367 = ~new_P2_U3878 | ~new_P2_U3385;
  assign new_P2_U3368 = ~new_P2_U3764 | ~new_P2_U3886;
  assign new_P2_U3369 = ~new_P2_U3872 | ~new_P2_U3378;
  assign new_P2_U3370 = ~new_P2_U3781 | ~new_P2_U4988 | ~new_P2_U4987;
  assign new_P2_U3371 = ~new_P2_U5413 | ~new_P2_U3913;
  assign new_P2_U3372 = ~new_P2_U5423 | ~new_P2_U5422;
  assign new_P2_U3373 = ~new_P2_U5426 | ~new_P2_U5425;
  assign new_P2_U3374 = ~new_P2_U5429 | ~new_P2_U5428;
  assign new_P2_U3375 = ~new_P2_U5435 | ~new_P2_U5434;
  assign n1505 = ~new_P2_U5438 | ~new_P2_U5437;
  assign n1510 = ~new_P2_U5440 | ~new_P2_U5439;
  assign new_P2_U3378 = ~new_P2_U5442 | ~new_P2_U5441;
  assign new_P2_U3379 = ~new_P2_U5445 | ~new_P2_U5444;
  assign new_P2_U3380 = ~new_P2_U5448 | ~new_P2_U5447;
  assign new_P2_U3381 = ~new_P2_U5454 | ~new_P2_U5453;
  assign new_P2_U3382 = ~new_P2_U5457 | ~new_P2_U5456;
  assign new_P2_U3383 = ~new_P2_U5460 | ~new_P2_U5459;
  assign new_P2_U3384 = ~new_P2_U5463 | ~new_P2_U5462;
  assign new_P2_U3385 = ~new_P2_U5451 | ~new_P2_U5450;
  assign new_P2_U3386 = ~new_P2_U5466 | ~new_P2_U5465;
  assign new_P2_U3387 = ~new_P2_U5468 | ~new_P2_U5467;
  assign new_P2_U3388 = ~new_P2_U5471 | ~new_P2_U5470;
  assign new_P2_U3389 = ~new_P2_U5474 | ~new_P2_U5473;
  assign n1665 = ~new_P2_U5480 | ~new_P2_U5479;
  assign new_P2_U3391 = ~new_P2_U5482 | ~new_P2_U5481;
  assign new_P2_U3392 = ~new_P2_U5484 | ~new_P2_U5483;
  assign n1670 = ~new_P2_U5487 | ~new_P2_U5486;
  assign new_P2_U3394 = ~new_P2_U5489 | ~new_P2_U5488;
  assign new_P2_U3395 = ~new_P2_U5491 | ~new_P2_U5490;
  assign n1675 = ~new_P2_U5494 | ~new_P2_U5493;
  assign new_P2_U3397 = ~new_P2_U5496 | ~new_P2_U5495;
  assign new_P2_U3398 = ~new_P2_U5498 | ~new_P2_U5497;
  assign n1680 = ~new_P2_U5501 | ~new_P2_U5500;
  assign new_P2_U3400 = ~new_P2_U5503 | ~new_P2_U5502;
  assign new_P2_U3401 = ~new_P2_U5505 | ~new_P2_U5504;
  assign n1685 = ~new_P2_U5508 | ~new_P2_U5507;
  assign new_P2_U3403 = ~new_P2_U5510 | ~new_P2_U5509;
  assign new_P2_U3404 = ~new_P2_U5512 | ~new_P2_U5511;
  assign n1690 = ~new_P2_U5515 | ~new_P2_U5514;
  assign new_P2_U3406 = ~new_P2_U5517 | ~new_P2_U5516;
  assign new_P2_U3407 = ~new_P2_U5519 | ~new_P2_U5518;
  assign n1695 = ~new_P2_U5522 | ~new_P2_U5521;
  assign new_P2_U3409 = ~new_P2_U5524 | ~new_P2_U5523;
  assign new_P2_U3410 = ~new_P2_U5526 | ~new_P2_U5525;
  assign n1700 = ~new_P2_U5529 | ~new_P2_U5528;
  assign new_P2_U3412 = ~new_P2_U5531 | ~new_P2_U5530;
  assign new_P2_U3413 = ~new_P2_U5533 | ~new_P2_U5532;
  assign n1705 = ~new_P2_U5536 | ~new_P2_U5535;
  assign new_P2_U3415 = ~new_P2_U5538 | ~new_P2_U5537;
  assign new_P2_U3416 = ~new_P2_U5540 | ~new_P2_U5539;
  assign n1710 = ~new_P2_U5543 | ~new_P2_U5542;
  assign new_P2_U3418 = ~new_P2_U5545 | ~new_P2_U5544;
  assign new_P2_U3419 = ~new_P2_U5547 | ~new_P2_U5546;
  assign n1715 = ~new_P2_U5550 | ~new_P2_U5549;
  assign new_P2_U3421 = ~new_P2_U5552 | ~new_P2_U5551;
  assign new_P2_U3422 = ~new_P2_U5554 | ~new_P2_U5553;
  assign n1720 = ~new_P2_U5557 | ~new_P2_U5556;
  assign new_P2_U3424 = ~new_P2_U5559 | ~new_P2_U5558;
  assign new_P2_U3425 = ~new_P2_U5561 | ~new_P2_U5560;
  assign n1725 = ~new_P2_U5564 | ~new_P2_U5563;
  assign new_P2_U3427 = ~new_P2_U5566 | ~new_P2_U5565;
  assign new_P2_U3428 = ~new_P2_U5568 | ~new_P2_U5567;
  assign n1730 = ~new_P2_U5571 | ~new_P2_U5570;
  assign new_P2_U3430 = ~new_P2_U5573 | ~new_P2_U5572;
  assign new_P2_U3431 = ~new_P2_U5575 | ~new_P2_U5574;
  assign n1735 = ~new_P2_U5578 | ~new_P2_U5577;
  assign new_P2_U3433 = ~new_P2_U5580 | ~new_P2_U5579;
  assign new_P2_U3434 = ~new_P2_U5582 | ~new_P2_U5581;
  assign n1740 = ~new_P2_U5585 | ~new_P2_U5584;
  assign new_P2_U3436 = ~new_P2_U5587 | ~new_P2_U5586;
  assign new_P2_U3437 = ~new_P2_U5589 | ~new_P2_U5588;
  assign n1745 = ~new_P2_U5592 | ~new_P2_U5591;
  assign new_P2_U3439 = ~new_P2_U5594 | ~new_P2_U5593;
  assign new_P2_U3440 = ~new_P2_U5596 | ~new_P2_U5595;
  assign n1750 = ~new_P2_U5599 | ~new_P2_U5598;
  assign new_P2_U3442 = ~new_P2_U5601 | ~new_P2_U5600;
  assign new_P2_U3443 = ~new_P2_U5603 | ~new_P2_U5602;
  assign n1755 = ~new_P2_U5606 | ~new_P2_U5605;
  assign new_P2_U3445 = ~new_P2_U5608 | ~new_P2_U5607;
  assign n1760 = ~new_P2_U5611 | ~new_P2_U5610;
  assign n1765 = ~new_P2_U5613 | ~new_P2_U5612;
  assign n1770 = ~new_P2_U5615 | ~new_P2_U5614;
  assign n1775 = ~new_P2_U5617 | ~new_P2_U5616;
  assign n1780 = ~new_P2_U5619 | ~new_P2_U5618;
  assign n1785 = ~new_P2_U5621 | ~new_P2_U5620;
  assign n1790 = ~new_P2_U5623 | ~new_P2_U5622;
  assign n1795 = ~new_P2_U5625 | ~new_P2_U5624;
  assign n1800 = ~new_P2_U5627 | ~new_P2_U5626;
  assign n1805 = ~new_P2_U5629 | ~new_P2_U5628;
  assign n1810 = ~new_P2_U5631 | ~new_P2_U5630;
  assign n1815 = ~new_P2_U5633 | ~new_P2_U5632;
  assign n1820 = ~new_P2_U5635 | ~new_P2_U5634;
  assign n1825 = ~new_P2_U5639 | ~new_P2_U5638;
  assign n1830 = ~new_P2_U5641 | ~new_P2_U5640;
  assign n1835 = ~new_P2_U5643 | ~new_P2_U5642;
  assign n1840 = ~new_P2_U5645 | ~new_P2_U5644;
  assign n1845 = ~new_P2_U5647 | ~new_P2_U5646;
  assign n1850 = ~new_P2_U5649 | ~new_P2_U5648;
  assign n1855 = ~new_P2_U5651 | ~new_P2_U5650;
  assign n1860 = ~new_P2_U5653 | ~new_P2_U5652;
  assign n1865 = ~new_P2_U5655 | ~new_P2_U5654;
  assign n1870 = ~new_P2_U5657 | ~new_P2_U5656;
  assign n1875 = ~new_P2_U5659 | ~new_P2_U5658;
  assign n1880 = ~new_P2_U5661 | ~new_P2_U5660;
  assign n1885 = ~new_P2_U5663 | ~new_P2_U5662;
  assign n1890 = ~new_P2_U5665 | ~new_P2_U5664;
  assign n1895 = ~new_P2_U5667 | ~new_P2_U5666;
  assign n1900 = ~new_P2_U5669 | ~new_P2_U5668;
  assign n1905 = ~new_P2_U5671 | ~new_P2_U5670;
  assign n1910 = ~new_P2_U5673 | ~new_P2_U5672;
  assign n1915 = ~new_P2_U5675 | ~new_P2_U5674;
  assign n1920 = ~new_P2_U5677 | ~new_P2_U5676;
  assign n1925 = ~new_P2_U5679 | ~new_P2_U5678;
  assign n1930 = ~new_P2_U5681 | ~new_P2_U5680;
  assign n1935 = ~new_P2_U5683 | ~new_P2_U5682;
  assign n1940 = ~new_P2_U5685 | ~new_P2_U5684;
  assign n1945 = ~new_P2_U5687 | ~new_P2_U5686;
  assign n1950 = ~new_P2_U5689 | ~new_P2_U5688;
  assign n1955 = ~new_P2_U5691 | ~new_P2_U5690;
  assign n1960 = ~new_P2_U5693 | ~new_P2_U5692;
  assign n1965 = ~new_P2_U5695 | ~new_P2_U5694;
  assign n1970 = ~new_P2_U5697 | ~new_P2_U5696;
  assign n1975 = ~new_P2_U5699 | ~new_P2_U5698;
  assign n1980 = ~new_P2_U5701 | ~new_P2_U5700;
  assign n2245 = ~new_P2_U5766 | ~new_P2_U5765;
  assign n2250 = ~new_P2_U5768 | ~new_P2_U5767;
  assign n2255 = ~new_P2_U5770 | ~new_P2_U5769;
  assign n2260 = ~new_P2_U5772 | ~new_P2_U5771;
  assign n2265 = ~new_P2_U5774 | ~new_P2_U5773;
  assign n2270 = ~new_P2_U5776 | ~new_P2_U5775;
  assign n2275 = ~new_P2_U5778 | ~new_P2_U5777;
  assign n2280 = ~new_P2_U5780 | ~new_P2_U5779;
  assign n2285 = ~new_P2_U5782 | ~new_P2_U5781;
  assign n2290 = ~new_P2_U5784 | ~new_P2_U5783;
  assign n2295 = ~new_P2_U5786 | ~new_P2_U5785;
  assign n2300 = ~new_P2_U5788 | ~new_P2_U5787;
  assign n2305 = ~new_P2_U5790 | ~new_P2_U5789;
  assign n2310 = ~new_P2_U5792 | ~new_P2_U5791;
  assign n2315 = ~new_P2_U5794 | ~new_P2_U5793;
  assign n2320 = ~new_P2_U5796 | ~new_P2_U5795;
  assign n2325 = ~new_P2_U5798 | ~new_P2_U5797;
  assign n2330 = ~new_P2_U5800 | ~new_P2_U5799;
  assign n2335 = ~new_P2_U5802 | ~new_P2_U5801;
  assign n2340 = ~new_P2_U5804 | ~new_P2_U5803;
  assign n2345 = ~new_P2_U5806 | ~new_P2_U5805;
  assign n2350 = ~new_P2_U5808 | ~new_P2_U5807;
  assign n2355 = ~new_P2_U5810 | ~new_P2_U5809;
  assign n2360 = ~new_P2_U5812 | ~new_P2_U5811;
  assign n2365 = ~new_P2_U5814 | ~new_P2_U5813;
  assign n2370 = ~new_P2_U5816 | ~new_P2_U5815;
  assign n2375 = ~new_P2_U5818 | ~new_P2_U5817;
  assign n2380 = ~new_P2_U5820 | ~new_P2_U5819;
  assign n2385 = ~new_P2_U5822 | ~new_P2_U5821;
  assign n2390 = ~new_P2_U5824 | ~new_P2_U5823;
  assign n2395 = ~new_P2_U5826 | ~new_P2_U5825;
  assign n2400 = ~new_P2_U5828 | ~new_P2_U5827;
  assign new_P2_U3523 = ~new_P2_U5942 | ~new_P2_U5941;
  assign new_P2_U3524 = ~new_P2_U5944 | ~new_P2_U5943;
  assign new_P2_U3525 = ~new_P2_U5946 | ~new_P2_U5945;
  assign new_P2_U3526 = ~new_P2_U5948 | ~new_P2_U5947;
  assign new_P2_U3527 = ~new_P2_U5950 | ~new_P2_U5949;
  assign new_P2_U3528 = ~new_P2_U5952 | ~new_P2_U5951;
  assign new_P2_U3529 = ~new_P2_U5954 | ~new_P2_U5953;
  assign new_P2_U3530 = ~new_P2_U5956 | ~new_P2_U5955;
  assign new_P2_U3531 = ~new_P2_U5958 | ~new_P2_U5957;
  assign new_P2_U3532 = ~new_P2_U5960 | ~new_P2_U5959;
  assign new_P2_U3533 = ~new_P2_U5962 | ~new_P2_U5961;
  assign new_P2_U3534 = ~new_P2_U5964 | ~new_P2_U5963;
  assign new_P2_U3535 = ~new_P2_U5966 | ~new_P2_U5965;
  assign new_P2_U3536 = ~new_P2_U5968 | ~new_P2_U5967;
  assign new_P2_U3537 = ~new_P2_U5970 | ~new_P2_U5969;
  assign new_P2_U3538 = ~new_P2_U5972 | ~new_P2_U5971;
  assign new_P2_U3539 = ~new_P2_U5974 | ~new_P2_U5973;
  assign new_P2_U3540 = ~new_P2_U5976 | ~new_P2_U5975;
  assign new_P2_U3541 = ~new_P2_U5978 | ~new_P2_U5977;
  assign new_P2_U3542 = ~new_P2_U5980 | ~new_P2_U5979;
  assign new_P2_U3543 = ~new_P2_U5982 | ~new_P2_U5981;
  assign new_P2_U3544 = ~new_P2_U5984 | ~new_P2_U5983;
  assign new_P2_U3545 = ~new_P2_U5986 | ~new_P2_U5985;
  assign new_P2_U3546 = ~new_P2_U5988 | ~new_P2_U5987;
  assign new_P2_U3547 = ~new_P2_U5990 | ~new_P2_U5989;
  assign new_P2_U3548 = ~new_P2_U5992 | ~new_P2_U5991;
  assign new_P2_U3549 = ~new_P2_U5994 | ~new_P2_U5993;
  assign new_P2_U3550 = ~new_P2_U5996 | ~new_P2_U5995;
  assign new_P2_U3551 = ~new_P2_U5998 | ~new_P2_U5997;
  assign new_P2_U3552 = ~new_P2_U6000 | ~new_P2_U5999;
  assign new_P2_U3553 = ~new_P2_U6002 | ~new_P2_U6001;
  assign new_P2_U3554 = ~new_P2_U6004 | ~new_P2_U6003;
  assign new_P2_U3555 = ~new_P2_U6006 | ~new_P2_U6005;
  assign new_P2_U3556 = ~new_P2_U6008 | ~new_P2_U6007;
  assign new_P2_U3557 = ~new_P2_U6010 | ~new_P2_U6009;
  assign new_P2_U3558 = ~new_P2_U6012 | ~new_P2_U6011;
  assign new_P2_U3559 = ~new_P2_U6014 | ~new_P2_U6013;
  assign new_P2_U3560 = ~new_P2_U6016 | ~new_P2_U6015;
  assign new_P2_U3561 = ~new_P2_U6018 | ~new_P2_U6017;
  assign new_P2_U3562 = ~new_P2_U6020 | ~new_P2_U6019;
  assign new_P2_U3563 = ~new_P2_U6022 | ~new_P2_U6021;
  assign new_P2_U3564 = ~new_P2_U6024 | ~new_P2_U6023;
  assign new_P2_U3565 = ~new_P2_U6026 | ~new_P2_U6025;
  assign new_P2_U3566 = ~new_P2_U6028 | ~new_P2_U6027;
  assign new_P2_U3567 = ~new_P2_U6030 | ~new_P2_U6029;
  assign new_P2_U3568 = ~new_P2_U6032 | ~new_P2_U6031;
  assign new_P2_U3569 = ~new_P2_U6034 | ~new_P2_U6033;
  assign new_P2_U3570 = ~new_P2_U6036 | ~new_P2_U6035;
  assign new_P2_U3571 = ~new_P2_U6038 | ~new_P2_U6037;
  assign new_P2_U3572 = ~new_P2_U6040 | ~new_P2_U6039;
  assign new_P2_U3573 = ~new_P2_U6042 | ~new_P2_U6041;
  assign new_P2_U3574 = ~new_P2_U6044 | ~new_P2_U6043;
  assign new_P2_U3575 = new_P2_U4062 & new_P2_U4061;
  assign new_P2_U3576 = new_P2_U4064 & new_P2_U4063;
  assign new_P2_U3577 = new_P2_U4071 & new_P2_U4072 & new_P2_U4070;
  assign new_P2_U3578 = new_P2_U4018 & new_P2_U4019 & new_P2_U4021 & new_P2_U4020;
  assign new_P2_U3579 = new_P2_U4022 & new_P2_U4023 & new_P2_U4025 & new_P2_U4024;
  assign new_P2_U3580 = new_P2_U4026 & new_P2_U4027 & new_P2_U4029 & new_P2_U4028;
  assign new_P2_U3581 = new_P2_U4032 & new_P2_U4031 & new_P2_U4030;
  assign new_P2_U3582 = new_P2_U3578 & new_P2_U3579 & new_P2_U3581 & new_P2_U3580;
  assign new_P2_U3583 = new_P2_U4033 & new_P2_U4034 & new_P2_U4036 & new_P2_U4035;
  assign new_P2_U3584 = new_P2_U4037 & new_P2_U4038 & new_P2_U4040 & new_P2_U4039;
  assign new_P2_U3585 = new_P2_U4041 & new_P2_U4042 & new_P2_U4044 & new_P2_U4043;
  assign new_P2_U3586 = new_P2_U4047 & new_P2_U4046 & new_P2_U4045;
  assign new_P2_U3587 = new_P2_U3583 & new_P2_U3584 & new_P2_U3586 & new_P2_U3585;
  assign new_P2_U3588 = new_P2_U3389 & new_P2_U3388;
  assign new_P2_U3589 = new_P2_U5475 & new_P2_U5472;
  assign new_P2_U3590 = new_P2_U4089 & new_P2_U4088;
  assign new_P2_U3591 = new_P2_U4091 & new_P2_U4090;
  assign new_P2_U3592 = new_P2_U3591 & new_P2_U4093 & new_P2_U4092;
  assign new_P2_U3593 = new_P2_U4095 & new_P2_U4096 & new_P2_U4097;
  assign new_P2_U3594 = new_P2_U4107 & new_P2_U4106;
  assign new_P2_U3595 = new_P2_U4109 & new_P2_U4108;
  assign new_P2_U3596 = new_P2_U3595 & new_P2_U4111 & new_P2_U4110;
  assign new_P2_U3597 = new_P2_U4113 & new_P2_U4114 & new_P2_U4115;
  assign new_P2_U3598 = new_P2_U4125 & new_P2_U4124;
  assign new_P2_U3599 = new_P2_U4127 & new_P2_U4126;
  assign new_P2_U3600 = new_P2_U3599 & new_P2_U4129 & new_P2_U4128;
  assign new_P2_U3601 = new_P2_U4131 & new_P2_U4132 & new_P2_U4133;
  assign new_P2_U3602 = new_P2_U4143 & new_P2_U4142;
  assign new_P2_U3603 = new_P2_U4145 & new_P2_U4144;
  assign new_P2_U3604 = new_P2_U3603 & new_P2_U4147 & new_P2_U4146;
  assign new_P2_U3605 = new_P2_U4149 & new_P2_U4150 & new_P2_U4151;
  assign new_P2_U3606 = new_P2_U4161 & new_P2_U4160;
  assign new_P2_U3607 = new_P2_U4163 & new_P2_U4162;
  assign new_P2_U3608 = new_P2_U3607 & new_P2_U4165 & new_P2_U4164;
  assign new_P2_U3609 = new_P2_U4167 & new_P2_U4168 & new_P2_U4169;
  assign new_P2_U3610 = new_P2_U4179 & new_P2_U4178;
  assign new_P2_U3611 = new_P2_U4181 & new_P2_U4180;
  assign new_P2_U3612 = new_P2_U3611 & new_P2_U4183 & new_P2_U4182;
  assign new_P2_U3613 = new_P2_U4185 & new_P2_U4186 & new_P2_U4187;
  assign new_P2_U3614 = new_P2_U4197 & new_P2_U4196;
  assign new_P2_U3615 = new_P2_U4199 & new_P2_U4198;
  assign new_P2_U3616 = new_P2_U3615 & new_P2_U4201 & new_P2_U4200;
  assign new_P2_U3617 = new_P2_U4203 & new_P2_U4204 & new_P2_U4205;
  assign new_P2_U3618 = new_P2_U4217 & new_P2_U4216;
  assign new_P2_U3619 = new_P2_U3618 & new_P2_U4219 & new_P2_U4218;
  assign new_P2_U3620 = new_P2_U4221 & new_P2_U4222 & new_P2_U4223;
  assign new_P2_U3621 = new_P2_U4235 & new_P2_U4234;
  assign new_P2_U3622 = new_P2_U3621 & new_P2_U4237 & new_P2_U4236;
  assign new_P2_U3623 = new_P2_U4239 & new_P2_U4240 & new_P2_U4241;
  assign new_P2_U3624 = new_P2_U4253 & new_P2_U4252;
  assign new_P2_U3625 = new_P2_U3624 & new_P2_U4255 & new_P2_U4254;
  assign new_P2_U3626 = new_P2_U4257 & new_P2_U4258 & new_P2_U4259;
  assign new_P2_U3627 = new_P2_U4271 & new_P2_U4270;
  assign new_P2_U3628 = new_P2_U3627 & new_P2_U4273 & new_P2_U4272;
  assign new_P2_U3629 = new_P2_U4275 & new_P2_U4276 & new_P2_U4277;
  assign new_P2_U3630 = new_P2_U4287 & new_P2_U4286;
  assign new_P2_U3631 = new_P2_U4289 & new_P2_U4288;
  assign new_P2_U3632 = new_P2_U3631 & new_P2_U4291 & new_P2_U4290;
  assign new_P2_U3633 = new_P2_U4293 & new_P2_U4294 & new_P2_U4295;
  assign new_P2_U3634 = new_P2_U4305 & new_P2_U4304;
  assign new_P2_U3635 = new_P2_U4307 & new_P2_U4306;
  assign new_P2_U3636 = new_P2_U3635 & new_P2_U4309 & new_P2_U4308;
  assign new_P2_U3637 = new_P2_U4311 & new_P2_U4312 & new_P2_U4313;
  assign new_P2_U3638 = new_P2_U4325 & new_P2_U4324;
  assign new_P2_U3639 = new_P2_U3638 & new_P2_U4327 & new_P2_U4326;
  assign new_P2_U3640 = new_P2_U4329 & new_P2_U4330 & new_P2_U4331;
  assign new_P2_U3641 = new_P2_U4343 & new_P2_U4342;
  assign new_P2_U3642 = new_P2_U3641 & new_P2_U4345 & new_P2_U4344;
  assign new_P2_U3643 = new_P2_U4347 & new_P2_U4348 & new_P2_U4349;
  assign new_P2_U3644 = new_P2_U4361 & new_P2_U4360;
  assign new_P2_U3645 = new_P2_U3644 & new_P2_U4363 & new_P2_U4362;
  assign new_P2_U3646 = new_P2_U4365 & new_P2_U4366 & new_P2_U4367;
  assign new_P2_U3647 = new_P2_U4377 & new_P2_U4376;
  assign new_P2_U3648 = new_P2_U4379 & new_P2_U4378;
  assign new_P2_U3649 = new_P2_U3648 & new_P2_U4381 & new_P2_U4380;
  assign new_P2_U3650 = new_P2_U4383 & new_P2_U4384 & new_P2_U4385;
  assign new_P2_U3651 = new_P2_U4395 & new_P2_U4394;
  assign new_P2_U3652 = new_P2_U4397 & new_P2_U4396;
  assign new_P2_U3653 = new_P2_U3652 & new_P2_U4399 & new_P2_U4398;
  assign new_P2_U3654 = new_P2_U4401 & new_P2_U4402 & new_P2_U4403;
  assign new_P2_U3655 = new_P2_U4413 & new_P2_U4412;
  assign new_P2_U3656 = new_P2_U4415 & new_P2_U4414;
  assign new_P2_U3657 = new_P2_U3656 & new_P2_U4417 & new_P2_U4416;
  assign new_P2_U3658 = new_P2_U4419 & new_P2_U4420 & new_P2_U4421;
  assign new_P2_U3659 = new_P2_U4431 & new_P2_U4430;
  assign new_P2_U3660 = new_P2_U4433 & new_P2_U4432;
  assign new_P2_U3661 = new_P2_U3660 & new_P2_U4435 & new_P2_U4434;
  assign new_P2_U3662 = new_P2_U4437 & new_P2_U4438 & new_P2_U4439;
  assign new_P2_U3663 = new_P2_U4451 & new_P2_U4450;
  assign new_P2_U3664 = new_P2_U3663 & new_P2_U4453 & new_P2_U4452;
  assign new_P2_U3665 = new_P2_U4455 & new_P2_U4456 & new_P2_U4457;
  assign new_P2_U3666 = new_P2_U4469 & new_P2_U4468;
  assign new_P2_U3667 = new_P2_U3666 & new_P2_U4471 & new_P2_U4470;
  assign new_P2_U3668 = new_P2_U4473 & new_P2_U4474 & new_P2_U4475;
  assign new_P2_U3669 = new_P2_U4487 & new_P2_U4486;
  assign new_P2_U3670 = new_P2_U3669 & new_P2_U4489 & new_P2_U4488;
  assign new_P2_U3671 = new_P2_U4491 & new_P2_U4492 & new_P2_U4493;
  assign new_P2_U3672 = new_P2_U4503 & new_P2_U4502;
  assign new_P2_U3673 = new_P2_U4505 & new_P2_U4504;
  assign new_P2_U3674 = new_P2_U3673 & new_P2_U4507 & new_P2_U4506;
  assign new_P2_U3675 = new_P2_U4509 & new_P2_U4510 & new_P2_U4511;
  assign new_P2_U3676 = new_P2_U4521 & new_P2_U4520;
  assign new_P2_U3677 = new_P2_U4523 & new_P2_U4522;
  assign new_P2_U3678 = new_P2_U3677 & new_P2_U4525 & new_P2_U4524;
  assign new_P2_U3679 = new_P2_U4527 & new_P2_U4528 & new_P2_U4529;
  assign new_P2_U3680 = new_P2_U4539 & new_P2_U4538;
  assign new_P2_U3681 = new_P2_U4541 & new_P2_U4540;
  assign new_P2_U3682 = new_P2_U3681 & new_P2_U4543 & new_P2_U4542;
  assign new_P2_U3683 = new_P2_U4545 & new_P2_U4546 & new_P2_U4547;
  assign new_P2_U3684 = new_P2_U4557 & new_P2_U4556;
  assign new_P2_U3685 = new_P2_U4559 & new_P2_U4558;
  assign new_P2_U3686 = new_P2_U3685 & new_P2_U4561 & new_P2_U4560;
  assign new_P2_U3687 = new_P2_U4563 & new_P2_U4564 & new_P2_U4565;
  assign new_P2_U3688 = new_P2_U4575 & new_P2_U4574;
  assign new_P2_U3689 = new_P2_U4577 & new_P2_U4576;
  assign new_P2_U3690 = new_P2_U3689 & new_P2_U4579 & new_P2_U4578;
  assign new_P2_U3691 = new_P2_U4581 & new_P2_U4582 & new_P2_U4583;
  assign new_P2_U3692 = new_P2_U4596 & new_P2_U4595 & new_P2_U4594 & new_P2_U4593 & new_P2_U4592;
  assign new_P2_U3693 = new_P2_U4598 & new_P2_U4597;
  assign new_P2_U3694 = new_P2_U3693 & new_P2_U4600 & new_P2_U4599;
  assign new_P2_U3695 = new_P2_U4603 & new_P2_U4602;
  assign new_P2_U3696 = new_P2_U5472 & new_P2_U3389;
  assign new_P2_U3697 = new_P2_U5475 & new_P2_U3388;
  assign new_P2_U3698 = new_P2_U3916 & new_P2_U3379;
  assign new_P2_U3699 = new_P2_U5436 & P2_STATE_REG;
  assign new_P2_U3700 = new_P2_U5420 & new_P2_U3364;
  assign new_P2_U3701 = new_P2_U3375 & P2_STATE_REG;
  assign new_P2_U3702 = new_P2_U3307 & new_P2_U3306 & new_P2_U3305 & new_P2_U3301 & new_P2_U3308;
  assign new_P2_U3703 = new_P2_U3309 & new_P2_U3360;
  assign new_P2_U3704 = new_P2_U3706 & new_P2_U4761 & new_P2_U4759 & new_P2_U4758;
  assign new_P2_U3705 = new_P2_U4764 & new_P2_U4762;
  assign new_P2_U3706 = new_P2_U3705 & new_P2_U4763;
  assign new_P2_U3707 = new_P2_U3709 & new_P2_U4772 & new_P2_U4770 & new_P2_U4769;
  assign new_P2_U3708 = new_P2_U4775 & new_P2_U4773;
  assign new_P2_U3709 = new_P2_U3708 & new_P2_U4774;
  assign new_P2_U3710 = new_P2_U3712 & new_P2_U4783 & new_P2_U4781 & new_P2_U4780;
  assign new_P2_U3711 = new_P2_U4786 & new_P2_U4784;
  assign new_P2_U3712 = new_P2_U3711 & new_P2_U4785;
  assign new_P2_U3713 = new_P2_U3715 & new_P2_U4794 & new_P2_U4792 & new_P2_U4791;
  assign new_P2_U3714 = new_P2_U4797 & new_P2_U4795;
  assign new_P2_U3715 = new_P2_U3714 & new_P2_U4796;
  assign new_P2_U3716 = new_P2_U3718 & new_P2_U4805 & new_P2_U4803 & new_P2_U4802;
  assign new_P2_U3717 = new_P2_U4808 & new_P2_U4806;
  assign new_P2_U3718 = new_P2_U3717 & new_P2_U4807;
  assign new_P2_U3719 = new_P2_U3721 & new_P2_U4816 & new_P2_U4814 & new_P2_U4813;
  assign new_P2_U3720 = new_P2_U4819 & new_P2_U4817;
  assign new_P2_U3721 = new_P2_U3720 & new_P2_U4818;
  assign new_P2_U3722 = new_P2_U3724 & new_P2_U4827 & new_P2_U4825 & new_P2_U4824;
  assign new_P2_U3723 = new_P2_U4830 & new_P2_U4828;
  assign new_P2_U3724 = new_P2_U3723 & new_P2_U4829;
  assign new_P2_U3725 = new_P2_U3727 & new_P2_U4838 & new_P2_U4836 & new_P2_U4835;
  assign new_P2_U3726 = new_P2_U4841 & new_P2_U4839;
  assign new_P2_U3727 = new_P2_U3726 & new_P2_U4840;
  assign new_P2_U3728 = new_P2_U3730 & new_P2_U4846 & new_P2_U4847 & new_P2_U4849;
  assign new_P2_U3729 = new_P2_U4852 & new_P2_U4850;
  assign new_P2_U3730 = new_P2_U3729 & new_P2_U4851;
  assign new_P2_U3731 = new_P2_U3733 & new_P2_U4857 & new_P2_U4858 & new_P2_U4860;
  assign new_P2_U3732 = new_P2_U4863 & new_P2_U4861;
  assign new_P2_U3733 = new_P2_U3732 & new_P2_U4862;
  assign new_P2_U3734 = new_P2_U3736 & new_P2_U4868 & new_P2_U4869 & new_P2_U4871;
  assign new_P2_U3735 = new_P2_U4874 & new_P2_U4872;
  assign new_P2_U3736 = new_P2_U3735 & new_P2_U4873;
  assign new_P2_U3737 = new_P2_U4880 & new_P2_U4879;
  assign new_P2_U3738 = new_P2_U4882 & new_P2_U3739 & new_P2_U4884;
  assign new_P2_U3739 = new_P2_U4885 & new_P2_U4883;
  assign new_P2_U3740 = new_P2_U4891 & new_P2_U4890;
  assign new_P2_U3741 = new_P2_U4893 & new_P2_U3742 & new_P2_U4895;
  assign new_P2_U3742 = new_P2_U4896 & new_P2_U4894;
  assign new_P2_U3743 = new_P2_U3745 & new_P2_U4904 & new_P2_U4902;
  assign new_P2_U3744 = new_P2_U4907 & new_P2_U4905;
  assign new_P2_U3745 = new_P2_U3744 & new_P2_U4906;
  assign new_P2_U3746 = new_P2_U4915 & new_P2_U4913;
  assign new_P2_U3747 = new_P2_U4918 & new_P2_U4916;
  assign new_P2_U3748 = new_P2_U3747 & new_P2_U4917;
  assign new_P2_U3749 = new_P2_U4923 & new_P2_U4924 & new_P2_U3751;
  assign new_P2_U3750 = new_P2_U4929 & new_P2_U4927;
  assign new_P2_U3751 = new_P2_U3750 & new_P2_U4928;
  assign new_P2_U3752 = new_P2_U4934 & new_P2_U4935 & new_P2_U3754;
  assign new_P2_U3753 = new_P2_U4940 & new_P2_U4938;
  assign new_P2_U3754 = new_P2_U3753 & new_P2_U4939;
  assign new_P2_U3755 = new_P2_U3757 & new_P2_U4945 & new_P2_U4946 & new_P2_U4948;
  assign new_P2_U3756 = new_P2_U4951 & new_P2_U4949;
  assign new_P2_U3757 = new_P2_U3756 & new_P2_U4950;
  assign new_P2_U3758 = new_P2_U3760 & new_P2_U4959 & new_P2_U4957 & new_P2_U4956;
  assign new_P2_U3759 = new_P2_U4962 & new_P2_U4960;
  assign new_P2_U3760 = new_P2_U3759 & new_P2_U4961;
  assign new_P2_U3761 = new_P2_U3763 & new_P2_U4970 & new_P2_U4968 & new_P2_U4967;
  assign new_P2_U3762 = new_P2_U4973 & new_P2_U4971;
  assign new_P2_U3763 = new_P2_U3762 & new_P2_U4972;
  assign new_P2_U3764 = new_P2_U5464 & new_P2_U3383;
  assign new_P2_U3765 = ~new_P2_U5830 | ~new_P2_U5829;
  assign new_P2_U3766 = new_P2_U5911 & new_P2_U5908;
  assign new_P2_U3767 = new_P2_U5893 & new_P2_U3766 & new_P2_U3769 & new_P2_U3768;
  assign new_P2_U3768 = new_P2_U5899 & new_P2_U5896;
  assign new_P2_U3769 = new_P2_U5905 & new_P2_U5902;
  assign new_P2_U3770 = new_P2_U5872 & new_P2_U5878 & new_P2_U5875;
  assign new_P2_U3771 = new_P2_U5890 & new_P2_U5881 & new_P2_U5887 & new_P2_U5884;
  assign new_P2_U3772 = new_P2_U5869 & new_P2_U3771 & new_P2_U3770;
  assign new_P2_U3773 = new_P2_U5854 & new_P2_U5857 & new_P2_U5863 & new_P2_U5860;
  assign new_P2_U3774 = new_P2_U5851 & new_P2_U5848;
  assign new_P2_U3775 = new_P2_U5917 & new_P2_U5920 & new_P2_U5926 & new_P2_U5923;
  assign new_P2_U3776 = new_P2_U5842 & new_P2_U5839 & new_P2_U5836;
  assign new_P2_U3777 = new_P2_U3776 & new_P2_U5845 & new_P2_U5866 & new_P2_U3773 & new_P2_U3774;
  assign new_P2_U3778 = new_P2_U5929 & new_P2_U3775 & new_P2_U5914 & new_P2_U3767 & new_P2_U3772;
  assign new_P2_U3779 = new_P2_U4976 & new_P2_U4977 & new_P2_U3866;
  assign new_P2_U3780 = new_P2_U5412 & new_P2_U5411;
  assign new_P2_U3781 = new_P2_U3876 & new_P2_U4986 & new_P2_U5436 & new_P2_U3362;
  assign new_P2_U3782 = new_P2_U4994 & new_P2_U4993;
  assign new_P2_U3783 = new_P2_U5007 & new_P2_U5006;
  assign new_P2_U3784 = new_P2_U5016 & new_P2_U5015;
  assign new_P2_U3785 = new_P2_U5025 & new_P2_U5024;
  assign new_P2_U3786 = new_P2_U5032 & new_P2_U5030;
  assign new_P2_U3787 = new_P2_U5034 & new_P2_U5033;
  assign new_P2_U3788 = new_P2_U5043 & new_P2_U5042;
  assign new_P2_U3789 = new_P2_U5052 & new_P2_U5051;
  assign new_P2_U3790 = new_P2_U5061 & new_P2_U5060;
  assign new_P2_U3791 = new_P2_U5070 & new_P2_U5069;
  assign new_P2_U3792 = new_P2_U3031 & new_P2_U3077;
  assign new_P2_U3793 = new_P2_U5074 & new_P2_U5073;
  assign new_P2_U3794 = new_P2_U3793 & new_P2_U5077 & new_P2_U5076;
  assign new_P2_U3795 = new_P2_U5086 & new_P2_U5085;
  assign new_P2_U3796 = new_P2_U5093 & new_P2_U5091;
  assign new_P2_U3797 = new_P2_U5095 & new_P2_U5094;
  assign new_P2_U3798 = new_P2_U5104 & new_P2_U5103;
  assign new_P2_U3799 = new_P2_U5113 & new_P2_U5112;
  assign new_P2_U3800 = new_P2_U5122 & new_P2_U5121;
  assign new_P2_U3801 = new_P2_U5131 & new_P2_U5130;
  assign new_P2_U3802 = new_P2_U5140 & new_P2_U5139;
  assign new_P2_U3803 = new_P2_U5149 & new_P2_U5148;
  assign new_P2_U3804 = new_P2_U5158 & new_P2_U5157;
  assign new_P2_U3805 = new_P2_U5165 & new_P2_U5163;
  assign new_P2_U3806 = new_P2_U5167 & new_P2_U5166;
  assign new_P2_U3807 = new_P2_U5176 & new_P2_U5175;
  assign new_P2_U3808 = new_P2_U5185 & new_P2_U5184;
  assign new_P2_U3809 = new_P2_U5194 & new_P2_U5193;
  assign new_P2_U3810 = new_P2_U5201 & new_P2_U5199;
  assign new_P2_U3811 = new_P2_U5203 & new_P2_U5202;
  assign new_P2_U3812 = new_P2_U5212 & new_P2_U5211;
  assign new_P2_U3813 = new_P2_U5221 & new_P2_U5220;
  assign new_P2_U3814 = new_P2_U5230 & new_P2_U5229;
  assign new_P2_U3815 = new_P2_U5239 & new_P2_U5238;
  assign new_P2_U3816 = new_P2_U5248 & new_P2_U5247;
  assign new_P2_U3817 = new_P2_U5250 & P2_STATE_REG;
  assign new_P2_U3818 = new_P2_U5436 & new_P2_U3385;
  assign new_P2_U3819 = new_P2_U3385 & new_P2_U3375;
  assign new_P2_U3820 = new_P2_U3302 & new_P2_U3871 & new_P2_U3312;
  assign new_P2_U3821 = new_P2_U3310 & new_P2_U3357 & new_P2_U3873;
  assign new_P2_U3822 = new_P2_U3375 & new_P2_U5264;
  assign new_P2_U3823 = new_P2_U3375 & new_P2_U5270;
  assign new_P2_U3824 = new_P2_U3375 & new_P2_U5292;
  assign new_P2_U3825 = new_P2_U3375 & new_P2_U5314;
  assign new_P2_U3826 = new_P2_U3375 & new_P2_U5316;
  assign new_P2_U3827 = ~P2_IR_REG_31_;
  assign new_P2_U3828 = ~new_P2_U3023 | ~new_P2_U3300;
  assign new_P2_U3829 = ~new_P2_U5464 | ~new_P2_U5461;
  assign new_P2_U3830 = ~new_P2_U5452 | ~new_P2_U5443;
  assign new_P2_U3831 = ~new_P2_U3023 | ~new_P2_U4054;
  assign new_P2_U3832 = ~new_P2_U3023 | ~new_P2_U4618;
  assign new_P2_U3833 = new_P2_U5703 & new_P2_U5702;
  assign new_P2_U3834 = new_P2_U5705 & new_P2_U5704;
  assign new_P2_U3835 = new_P2_U5707 & new_P2_U5706;
  assign new_P2_U3836 = new_P2_U5709 & new_P2_U5708;
  assign new_P2_U3837 = new_P2_U5711 & new_P2_U5710;
  assign new_P2_U3838 = new_P2_U5713 & new_P2_U5712;
  assign new_P2_U3839 = new_P2_U5715 & new_P2_U5714;
  assign new_P2_U3840 = new_P2_U5717 & new_P2_U5716;
  assign new_P2_U3841 = new_P2_U5719 & new_P2_U5718;
  assign new_P2_U3842 = new_P2_U5721 & new_P2_U5720;
  assign new_P2_U3843 = new_P2_U5723 & new_P2_U5722;
  assign new_P2_U3844 = new_P2_U5725 & new_P2_U5724;
  assign new_P2_U3845 = new_P2_U5727 & new_P2_U5726;
  assign new_P2_U3846 = new_P2_U5729 & new_P2_U5728;
  assign new_P2_U3847 = new_P2_U5731 & new_P2_U5730;
  assign new_P2_U3848 = new_P2_U5733 & new_P2_U5732;
  assign new_P2_U3849 = new_P2_U5735 & new_P2_U5734;
  assign new_P2_U3850 = new_P2_U5737 & new_P2_U5736;
  assign new_P2_U3851 = new_P2_U5739 & new_P2_U5738;
  assign new_P2_U3852 = new_P2_U5741 & new_P2_U5740;
  assign new_P2_U3853 = new_P2_U5743 & new_P2_U5742;
  assign new_P2_U3854 = new_P2_U5745 & new_P2_U5744;
  assign new_P2_U3855 = new_P2_U5747 & new_P2_U5746;
  assign new_P2_U3856 = new_P2_U5749 & new_P2_U5748;
  assign new_P2_U3857 = new_P2_U5751 & new_P2_U5750;
  assign new_P2_U3858 = new_P2_U5753 & new_P2_U5752;
  assign new_P2_U3859 = new_P2_U5755 & new_P2_U5754;
  assign new_P2_U3860 = new_P2_U5757 & new_P2_U5756;
  assign new_P2_U3861 = new_P2_U5759 & new_P2_U5758;
  assign new_P2_U3862 = new_P2_U5761 & new_P2_U5760;
  assign new_P2_U3863 = ~new_P2_R1269_U22;
  assign new_P2_U3864 = ~new_P2_U3778 | ~new_P2_U3777;
  assign new_P2_U3865 = ~new_P2_R693_U14;
  assign new_P2_U3866 = new_P2_U5936 & new_P2_U5935;
  assign new_P2_U3867 = ~new_P2_R1297_U6;
  assign new_P2_U3868 = ~new_P2_U3356;
  assign new_P2_U3869 = ~new_P2_U3355;
  assign new_P2_U3870 = ~new_P2_U3312;
  assign new_P2_U3871 = ~new_P2_U3015 | ~new_P2_U3385;
  assign new_P2_U3872 = ~new_P2_U3302;
  assign new_P2_U3873 = ~new_P2_U3016 | ~new_P2_U5452;
  assign new_P2_U3874 = ~new_P2_U3310;
  assign new_P2_U3875 = ~new_P2_U3357;
  assign new_P2_U3876 = ~new_P2_U3014 | ~new_P2_U3385;
  assign new_P2_U3877 = ~new_P2_U3308;
  assign new_P2_U3878 = ~new_P2_U3301;
  assign new_P2_U3879 = ~new_P2_U3305;
  assign new_P2_U3880 = ~new_P2_U3307;
  assign new_P2_U3881 = ~new_P2_U3306;
  assign new_P2_U3882 = ~new_P2_U3360;
  assign new_P2_U3883 = ~new_P2_U3311;
  assign new_P2_U3884 = ~new_P2_U3874 | ~new_P2_U3378;
  assign new_P2_U3885 = ~new_P2_U3369;
  assign new_P2_U3886 = ~new_P2_U3367;
  assign new_P2_U3887 = ~new_P2_U3309;
  assign new_P2_U3888 = ~new_P2_U3352;
  assign new_P2_U3889 = ~new_P2_U3829;
  assign new_P2_U3890 = ~new_P2_U3303;
  assign new_P2_U3891 = ~new_P2_U3304;
  assign new_P2_U3892 = ~new_P2_U5461 | ~new_P2_U3384;
  assign n2565 = ~new_P2_U3363;
  assign new_P2_U3894 = ~new_P2_U3364;
  assign new_P2_U3895 = ~new_P2_U3350;
  assign new_P2_U3896 = ~new_P2_U3348;
  assign new_P2_U3897 = ~new_P2_U3346;
  assign new_P2_U3898 = ~new_P2_U3344;
  assign new_P2_U3899 = ~new_P2_U3342;
  assign new_P2_U3900 = ~new_P2_U3340;
  assign new_P2_U3901 = ~new_P2_U3338;
  assign new_P2_U3902 = ~new_P2_U3336;
  assign new_P2_U3903 = ~new_P2_U3334;
  assign new_P2_U3904 = ~new_P2_U3353;
  assign new_P2_U3905 = ~new_P2_U3368;
  assign new_P2_U3906 = ~new_P2_U3362;
  assign new_P2_U3907 = ~new_P2_U3313;
  assign new_P2_U3908 = ~new_P2_U3358;
  assign new_P2_U3909 = ~new_P2_U3832;
  assign new_P2_U3910 = ~new_P2_U3831;
  assign new_P2_U3911 = ~new_P2_U3828;
  assign new_P2_U3912 = ~new_P2_U3361;
  assign new_P2_U3913 = ~new_P2_U3370 | ~P2_STATE_REG;
  assign new_P2_U3914 = ~new_P2_U3882 | ~new_P2_U3023;
  assign new_P2_U3915 = ~new_P2_U3299;
  assign new_P2_U3916 = ~new_P2_U3359;
  assign new_P2_U3917 = ~new_P2_U3297;
  assign new_P2_U3918 = ~new_U56 | ~n2555;
  assign new_P2_U3919 = ~P2_IR_REG_0_ | ~new_P2_U3027;
  assign new_P2_U3920 = ~P2_IR_REG_0_ | ~new_P2_U3917;
  assign new_P2_U3921 = ~new_U45 | ~n2555;
  assign new_P2_U3922 = ~new_P2_SUB_594_U53 | ~new_P2_U3027;
  assign new_P2_U3923 = ~P2_IR_REG_1_ | ~new_P2_U3917;
  assign new_P2_U3924 = ~new_U34 | ~n2555;
  assign new_P2_U3925 = ~new_P2_SUB_594_U23 | ~new_P2_U3027;
  assign new_P2_U3926 = ~P2_IR_REG_2_ | ~new_P2_U3917;
  assign new_P2_U3927 = ~new_U31 | ~n2555;
  assign new_P2_U3928 = ~new_P2_SUB_594_U24 | ~new_P2_U3027;
  assign new_P2_U3929 = ~P2_IR_REG_3_ | ~new_P2_U3917;
  assign new_P2_U3930 = ~new_U30 | ~n2555;
  assign new_P2_U3931 = ~new_P2_SUB_594_U25 | ~new_P2_U3027;
  assign new_P2_U3932 = ~P2_IR_REG_4_ | ~new_P2_U3917;
  assign new_P2_U3933 = ~new_U29 | ~n2555;
  assign new_P2_U3934 = ~new_P2_SUB_594_U72 | ~new_P2_U3027;
  assign new_P2_U3935 = ~P2_IR_REG_5_ | ~new_P2_U3917;
  assign new_P2_U3936 = ~new_U28 | ~n2555;
  assign new_P2_U3937 = ~new_P2_SUB_594_U26 | ~new_P2_U3027;
  assign new_P2_U3938 = ~P2_IR_REG_6_ | ~new_P2_U3917;
  assign new_P2_U3939 = ~new_U27 | ~n2555;
  assign new_P2_U3940 = ~new_P2_SUB_594_U27 | ~new_P2_U3027;
  assign new_P2_U3941 = ~P2_IR_REG_7_ | ~new_P2_U3917;
  assign new_P2_U3942 = ~new_U26 | ~n2555;
  assign new_P2_U3943 = ~new_P2_SUB_594_U28 | ~new_P2_U3027;
  assign new_P2_U3944 = ~P2_IR_REG_8_ | ~new_P2_U3917;
  assign new_P2_U3945 = ~new_U25 | ~n2555;
  assign new_P2_U3946 = ~new_P2_SUB_594_U70 | ~new_P2_U3027;
  assign new_P2_U3947 = ~P2_IR_REG_9_ | ~new_P2_U3917;
  assign new_P2_U3948 = ~new_U55 | ~n2555;
  assign new_P2_U3949 = ~new_P2_SUB_594_U8 | ~new_P2_U3027;
  assign new_P2_U3950 = ~P2_IR_REG_10_ | ~new_P2_U3917;
  assign new_P2_U3951 = ~new_U54 | ~n2555;
  assign new_P2_U3952 = ~new_P2_SUB_594_U9 | ~new_P2_U3027;
  assign new_P2_U3953 = ~P2_IR_REG_11_ | ~new_P2_U3917;
  assign new_P2_U3954 = ~new_U53 | ~n2555;
  assign new_P2_U3955 = ~new_P2_SUB_594_U10 | ~new_P2_U3027;
  assign new_P2_U3956 = ~P2_IR_REG_12_ | ~new_P2_U3917;
  assign new_P2_U3957 = ~new_U52 | ~n2555;
  assign new_P2_U3958 = ~new_P2_SUB_594_U87 | ~new_P2_U3027;
  assign new_P2_U3959 = ~P2_IR_REG_13_ | ~new_P2_U3917;
  assign new_P2_U3960 = ~new_U51 | ~n2555;
  assign new_P2_U3961 = ~new_P2_SUB_594_U11 | ~new_P2_U3027;
  assign new_P2_U3962 = ~P2_IR_REG_14_ | ~new_P2_U3917;
  assign new_P2_U3963 = ~new_U50 | ~n2555;
  assign new_P2_U3964 = ~new_P2_SUB_594_U12 | ~new_P2_U3027;
  assign new_P2_U3965 = ~P2_IR_REG_15_ | ~new_P2_U3917;
  assign new_P2_U3966 = ~new_U49 | ~n2555;
  assign new_P2_U3967 = ~new_P2_SUB_594_U13 | ~new_P2_U3027;
  assign new_P2_U3968 = ~P2_IR_REG_16_ | ~new_P2_U3917;
  assign new_P2_U3969 = ~new_U48 | ~n2555;
  assign new_P2_U3970 = ~new_P2_SUB_594_U85 | ~new_P2_U3027;
  assign new_P2_U3971 = ~P2_IR_REG_17_ | ~new_P2_U3917;
  assign new_P2_U3972 = ~new_U47 | ~n2555;
  assign new_P2_U3973 = ~new_P2_SUB_594_U14 | ~new_P2_U3027;
  assign new_P2_U3974 = ~P2_IR_REG_18_ | ~new_P2_U3917;
  assign new_P2_U3975 = ~new_U46 | ~n2555;
  assign new_P2_U3976 = ~new_P2_SUB_594_U15 | ~new_P2_U3027;
  assign new_P2_U3977 = ~P2_IR_REG_19_ | ~new_P2_U3917;
  assign new_P2_U3978 = ~new_U44 | ~n2555;
  assign new_P2_U3979 = ~new_P2_SUB_594_U16 | ~new_P2_U3027;
  assign new_P2_U3980 = ~P2_IR_REG_20_ | ~new_P2_U3917;
  assign new_P2_U3981 = ~new_U43 | ~n2555;
  assign new_P2_U3982 = ~new_P2_SUB_594_U81 | ~new_P2_U3027;
  assign new_P2_U3983 = ~P2_IR_REG_21_ | ~new_P2_U3917;
  assign new_P2_U3984 = ~new_U42 | ~n2555;
  assign new_P2_U3985 = ~new_P2_SUB_594_U17 | ~new_P2_U3027;
  assign new_P2_U3986 = ~P2_IR_REG_22_ | ~new_P2_U3917;
  assign new_P2_U3987 = ~new_U41 | ~n2555;
  assign new_P2_U3988 = ~new_P2_SUB_594_U18 | ~new_P2_U3027;
  assign new_P2_U3989 = ~P2_IR_REG_23_ | ~new_P2_U3917;
  assign new_P2_U3990 = ~new_U40 | ~n2555;
  assign new_P2_U3991 = ~new_P2_SUB_594_U19 | ~new_P2_U3027;
  assign new_P2_U3992 = ~P2_IR_REG_24_ | ~new_P2_U3917;
  assign new_P2_U3993 = ~new_U39 | ~n2555;
  assign new_P2_U3994 = ~new_P2_SUB_594_U79 | ~new_P2_U3027;
  assign new_P2_U3995 = ~P2_IR_REG_25_ | ~new_P2_U3917;
  assign new_P2_U3996 = ~new_U38 | ~n2555;
  assign new_P2_U3997 = ~new_P2_SUB_594_U20 | ~new_P2_U3027;
  assign new_P2_U3998 = ~P2_IR_REG_26_ | ~new_P2_U3917;
  assign new_P2_U3999 = ~new_U37 | ~n2555;
  assign new_P2_U4000 = ~new_P2_SUB_594_U77 | ~new_P2_U3027;
  assign new_P2_U4001 = ~P2_IR_REG_27_ | ~new_P2_U3917;
  assign new_P2_U4002 = ~new_U36 | ~n2555;
  assign new_P2_U4003 = ~new_P2_SUB_594_U21 | ~new_P2_U3027;
  assign new_P2_U4004 = ~P2_IR_REG_28_ | ~new_P2_U3917;
  assign new_P2_U4005 = ~new_U35 | ~n2555;
  assign new_P2_U4006 = ~new_P2_SUB_594_U22 | ~new_P2_U3027;
  assign new_P2_U4007 = ~P2_IR_REG_29_ | ~new_P2_U3917;
  assign new_P2_U4008 = ~new_U33 | ~n2555;
  assign new_P2_U4009 = ~new_P2_SUB_594_U75 | ~new_P2_U3027;
  assign new_P2_U4010 = ~P2_IR_REG_30_ | ~new_P2_U3917;
  assign new_P2_U4011 = ~new_U32 | ~n2555;
  assign new_P2_U4012 = ~new_P2_SUB_594_U54 | ~new_P2_U3027;
  assign new_P2_U4013 = ~P2_IR_REG_31_ | ~new_P2_U3917;
  assign new_P2_U4014 = ~new_P2_U3915 | ~new_P2_U5433;
  assign new_P2_U4015 = ~new_P2_U3300;
  assign new_P2_U4016 = ~new_P2_U3299 | ~new_P2_U5424;
  assign new_P2_U4017 = ~new_P2_U3299 | ~new_P2_U5427;
  assign new_P2_U4018 = ~new_P2_U4015 | ~P2_D_REG_10_;
  assign new_P2_U4019 = ~new_P2_U4015 | ~P2_D_REG_11_;
  assign new_P2_U4020 = ~new_P2_U4015 | ~P2_D_REG_12_;
  assign new_P2_U4021 = ~new_P2_U4015 | ~P2_D_REG_13_;
  assign new_P2_U4022 = ~new_P2_U4015 | ~P2_D_REG_14_;
  assign new_P2_U4023 = ~new_P2_U4015 | ~P2_D_REG_15_;
  assign new_P2_U4024 = ~new_P2_U4015 | ~P2_D_REG_16_;
  assign new_P2_U4025 = ~new_P2_U4015 | ~P2_D_REG_17_;
  assign new_P2_U4026 = ~new_P2_U4015 | ~P2_D_REG_18_;
  assign new_P2_U4027 = ~new_P2_U4015 | ~P2_D_REG_19_;
  assign new_P2_U4028 = ~new_P2_U4015 | ~P2_D_REG_20_;
  assign new_P2_U4029 = ~new_P2_U4015 | ~P2_D_REG_21_;
  assign new_P2_U4030 = ~new_P2_U4015 | ~P2_D_REG_22_;
  assign new_P2_U4031 = ~new_P2_U4015 | ~P2_D_REG_23_;
  assign new_P2_U4032 = ~new_P2_U4015 | ~P2_D_REG_24_;
  assign new_P2_U4033 = ~new_P2_U4015 | ~P2_D_REG_25_;
  assign new_P2_U4034 = ~new_P2_U4015 | ~P2_D_REG_26_;
  assign new_P2_U4035 = ~new_P2_U4015 | ~P2_D_REG_27_;
  assign new_P2_U4036 = ~new_P2_U4015 | ~P2_D_REG_28_;
  assign new_P2_U4037 = ~new_P2_U4015 | ~P2_D_REG_29_;
  assign new_P2_U4038 = ~new_P2_U4015 | ~P2_D_REG_2_;
  assign new_P2_U4039 = ~new_P2_U4015 | ~P2_D_REG_30_;
  assign new_P2_U4040 = ~new_P2_U4015 | ~P2_D_REG_31_;
  assign new_P2_U4041 = ~new_P2_U4015 | ~P2_D_REG_3_;
  assign new_P2_U4042 = ~new_P2_U4015 | ~P2_D_REG_4_;
  assign new_P2_U4043 = ~new_P2_U4015 | ~P2_D_REG_5_;
  assign new_P2_U4044 = ~new_P2_U4015 | ~P2_D_REG_6_;
  assign new_P2_U4045 = ~new_P2_U4015 | ~P2_D_REG_7_;
  assign new_P2_U4046 = ~new_P2_U4015 | ~P2_D_REG_8_;
  assign new_P2_U4047 = ~new_P2_U4015 | ~P2_D_REG_9_;
  assign new_P2_U4048 = ~new_P2_U3830;
  assign new_P2_U4049 = ~new_P2_U5452 | ~new_P2_U5446;
  assign new_P2_U4050 = ~new_P2_U5478 | ~new_P2_U4049;
  assign new_P2_U4051 = ~new_P2_U3369 | ~new_P2_U3367;
  assign new_P2_U4052 = ~new_P2_U3890 | ~new_P2_U4051;
  assign new_P2_U4053 = ~new_P2_U3891 | ~new_P2_U4050;
  assign new_P2_U4054 = ~new_P2_U4053 | ~new_P2_U4052;
  assign new_P2_U4055 = ~new_P2_U3022 | ~P2_REG0_REG_1_;
  assign new_P2_U4056 = ~P2_REG1_REG_1_ | ~new_P2_U3021;
  assign new_P2_U4057 = ~P2_REG2_REG_1_ | ~new_P2_U3020;
  assign new_P2_U4058 = ~P2_REG3_REG_1_ | ~new_P2_U3019;
  assign new_P2_U4059 = ~new_P2_U3077;
  assign new_P2_U4060 = ~new_P2_U3873 | ~new_P2_U3357;
  assign new_P2_U4061 = ~new_P2_U3879 | ~new_P2_R1110_U95;
  assign new_P2_U4062 = ~new_P2_U3881 | ~new_P2_R1077_U95;
  assign new_P2_U4063 = ~new_P2_U3880 | ~new_P2_R1095_U25;
  assign new_P2_U4064 = ~new_P2_U3877 | ~new_P2_R1143_U95;
  assign new_P2_U4065 = ~new_P2_U3887 | ~new_P2_R1161_U95;
  assign new_P2_U4066 = ~new_P2_U3883 | ~new_P2_R1131_U25;
  assign new_P2_U4067 = ~new_P2_U3017 | ~new_P2_R1200_U25;
  assign new_P2_U4068 = ~new_P2_U3314;
  assign new_P2_U4069 = ~new_P2_U3352 | ~new_P2_U3829;
  assign new_P2_U4070 = ~new_P2_R1179_U25 | ~new_P2_U3026;
  assign new_P2_U4071 = ~new_P2_U3025 | ~new_P2_U3077;
  assign new_P2_U4072 = ~new_P2_U3387 | ~new_P2_U4060;
  assign new_P2_U4073 = ~new_P2_U3577 | ~new_P2_U4068;
  assign new_P2_U4074 = ~P2_REG0_REG_2_ | ~new_P2_U3022;
  assign new_P2_U4075 = ~P2_REG1_REG_2_ | ~new_P2_U3021;
  assign new_P2_U4076 = ~P2_REG2_REG_2_ | ~new_P2_U3020;
  assign new_P2_U4077 = ~P2_REG3_REG_2_ | ~new_P2_U3019;
  assign new_P2_U4078 = ~new_P2_U3067;
  assign new_P2_U4079 = ~P2_REG0_REG_0_ | ~new_P2_U3022;
  assign new_P2_U4080 = ~P2_REG1_REG_0_ | ~new_P2_U3021;
  assign new_P2_U4081 = ~P2_REG2_REG_0_ | ~new_P2_U3020;
  assign new_P2_U4082 = ~P2_REG3_REG_0_ | ~new_P2_U3019;
  assign new_P2_U4083 = ~new_P2_U3076;
  assign new_P2_U4084 = ~new_P2_U5464 | ~new_P2_U3383;
  assign new_P2_U4085 = ~new_P2_U3892 | ~new_P2_U4084;
  assign new_P2_U4086 = ~new_P2_U3033 | ~new_P2_U3076;
  assign new_P2_U4087 = ~new_P2_R1110_U94 | ~new_P2_U3879;
  assign new_P2_U4088 = ~new_P2_R1077_U94 | ~new_P2_U3881;
  assign new_P2_U4089 = ~new_P2_R1095_U102 | ~new_P2_U3880;
  assign new_P2_U4090 = ~new_P2_R1143_U94 | ~new_P2_U3877;
  assign new_P2_U4091 = ~new_P2_R1161_U94 | ~new_P2_U3887;
  assign new_P2_U4092 = ~new_P2_R1131_U102 | ~new_P2_U3883;
  assign new_P2_U4093 = ~new_P2_R1200_U102 | ~new_P2_U3017;
  assign new_P2_U4094 = ~new_P2_U3315;
  assign new_P2_U4095 = ~new_P2_R1179_U102 | ~new_P2_U3026;
  assign new_P2_U4096 = ~new_P2_U3025 | ~new_P2_U3067;
  assign new_P2_U4097 = ~new_P2_U3392 | ~new_P2_U4060;
  assign new_P2_U4098 = ~new_P2_U3593 | ~new_P2_U4094;
  assign new_P2_U4099 = ~P2_REG0_REG_3_ | ~new_P2_U3022;
  assign new_P2_U4100 = ~P2_REG1_REG_3_ | ~new_P2_U3021;
  assign new_P2_U4101 = ~P2_REG2_REG_3_ | ~new_P2_U3020;
  assign new_P2_U4102 = ~new_P2_SUB_605_U26 | ~new_P2_U3019;
  assign new_P2_U4103 = ~new_P2_U3063;
  assign new_P2_U4104 = ~new_P2_U3033 | ~new_P2_U3077;
  assign new_P2_U4105 = ~new_P2_R1110_U16 | ~new_P2_U3879;
  assign new_P2_U4106 = ~new_P2_R1077_U16 | ~new_P2_U3881;
  assign new_P2_U4107 = ~new_P2_R1095_U112 | ~new_P2_U3880;
  assign new_P2_U4108 = ~new_P2_R1143_U16 | ~new_P2_U3877;
  assign new_P2_U4109 = ~new_P2_R1161_U16 | ~new_P2_U3887;
  assign new_P2_U4110 = ~new_P2_R1131_U112 | ~new_P2_U3883;
  assign new_P2_U4111 = ~new_P2_R1200_U112 | ~new_P2_U3017;
  assign new_P2_U4112 = ~new_P2_U3316;
  assign new_P2_U4113 = ~new_P2_R1179_U112 | ~new_P2_U3026;
  assign new_P2_U4114 = ~new_P2_U3025 | ~new_P2_U3063;
  assign new_P2_U4115 = ~new_P2_U3395 | ~new_P2_U4060;
  assign new_P2_U4116 = ~new_P2_U3597 | ~new_P2_U4112;
  assign new_P2_U4117 = ~P2_REG0_REG_4_ | ~new_P2_U3022;
  assign new_P2_U4118 = ~P2_REG1_REG_4_ | ~new_P2_U3021;
  assign new_P2_U4119 = ~P2_REG2_REG_4_ | ~new_P2_U3020;
  assign new_P2_U4120 = ~new_P2_SUB_605_U30 | ~new_P2_U3019;
  assign new_P2_U4121 = ~new_P2_U3059;
  assign new_P2_U4122 = ~new_P2_U3033 | ~new_P2_U3067;
  assign new_P2_U4123 = ~new_P2_R1110_U100 | ~new_P2_U3879;
  assign new_P2_U4124 = ~new_P2_R1077_U100 | ~new_P2_U3881;
  assign new_P2_U4125 = ~new_P2_R1095_U22 | ~new_P2_U3880;
  assign new_P2_U4126 = ~new_P2_R1143_U100 | ~new_P2_U3877;
  assign new_P2_U4127 = ~new_P2_R1161_U100 | ~new_P2_U3887;
  assign new_P2_U4128 = ~new_P2_R1131_U22 | ~new_P2_U3883;
  assign new_P2_U4129 = ~new_P2_R1200_U22 | ~new_P2_U3017;
  assign new_P2_U4130 = ~new_P2_U3317;
  assign new_P2_U4131 = ~new_P2_R1179_U22 | ~new_P2_U3026;
  assign new_P2_U4132 = ~new_P2_U3025 | ~new_P2_U3059;
  assign new_P2_U4133 = ~new_P2_U3398 | ~new_P2_U4060;
  assign new_P2_U4134 = ~new_P2_U3601 | ~new_P2_U4130;
  assign new_P2_U4135 = ~P2_REG0_REG_5_ | ~new_P2_U3022;
  assign new_P2_U4136 = ~P2_REG1_REG_5_ | ~new_P2_U3021;
  assign new_P2_U4137 = ~P2_REG2_REG_5_ | ~new_P2_U3020;
  assign new_P2_U4138 = ~new_P2_SUB_605_U22 | ~new_P2_U3019;
  assign new_P2_U4139 = ~new_P2_U3066;
  assign new_P2_U4140 = ~new_P2_U3033 | ~new_P2_U3063;
  assign new_P2_U4141 = ~new_P2_R1110_U99 | ~new_P2_U3879;
  assign new_P2_U4142 = ~new_P2_R1077_U99 | ~new_P2_U3881;
  assign new_P2_U4143 = ~new_P2_R1095_U111 | ~new_P2_U3880;
  assign new_P2_U4144 = ~new_P2_R1143_U99 | ~new_P2_U3877;
  assign new_P2_U4145 = ~new_P2_R1161_U99 | ~new_P2_U3887;
  assign new_P2_U4146 = ~new_P2_R1131_U111 | ~new_P2_U3883;
  assign new_P2_U4147 = ~new_P2_R1200_U111 | ~new_P2_U3017;
  assign new_P2_U4148 = ~new_P2_U3318;
  assign new_P2_U4149 = ~new_P2_R1179_U111 | ~new_P2_U3026;
  assign new_P2_U4150 = ~new_P2_U3025 | ~new_P2_U3066;
  assign new_P2_U4151 = ~new_P2_U3401 | ~new_P2_U4060;
  assign new_P2_U4152 = ~new_P2_U3605 | ~new_P2_U4148;
  assign new_P2_U4153 = ~P2_REG0_REG_6_ | ~new_P2_U3022;
  assign new_P2_U4154 = ~P2_REG1_REG_6_ | ~new_P2_U3021;
  assign new_P2_U4155 = ~P2_REG2_REG_6_ | ~new_P2_U3020;
  assign new_P2_U4156 = ~new_P2_SUB_605_U8 | ~new_P2_U3019;
  assign new_P2_U4157 = ~new_P2_U3070;
  assign new_P2_U4158 = ~new_P2_U3033 | ~new_P2_U3059;
  assign new_P2_U4159 = ~new_P2_R1110_U17 | ~new_P2_U3879;
  assign new_P2_U4160 = ~new_P2_R1077_U17 | ~new_P2_U3881;
  assign new_P2_U4161 = ~new_P2_R1095_U110 | ~new_P2_U3880;
  assign new_P2_U4162 = ~new_P2_R1143_U17 | ~new_P2_U3877;
  assign new_P2_U4163 = ~new_P2_R1161_U17 | ~new_P2_U3887;
  assign new_P2_U4164 = ~new_P2_R1131_U110 | ~new_P2_U3883;
  assign new_P2_U4165 = ~new_P2_R1200_U110 | ~new_P2_U3017;
  assign new_P2_U4166 = ~new_P2_U3319;
  assign new_P2_U4167 = ~new_P2_R1179_U110 | ~new_P2_U3026;
  assign new_P2_U4168 = ~new_P2_U3025 | ~new_P2_U3070;
  assign new_P2_U4169 = ~new_P2_U3404 | ~new_P2_U4060;
  assign new_P2_U4170 = ~new_P2_U3609 | ~new_P2_U4166;
  assign new_P2_U4171 = ~P2_REG0_REG_7_ | ~new_P2_U3022;
  assign new_P2_U4172 = ~P2_REG1_REG_7_ | ~new_P2_U3021;
  assign new_P2_U4173 = ~P2_REG2_REG_7_ | ~new_P2_U3020;
  assign new_P2_U4174 = ~new_P2_SUB_605_U18 | ~new_P2_U3019;
  assign new_P2_U4175 = ~new_P2_U3069;
  assign new_P2_U4176 = ~new_P2_U3033 | ~new_P2_U3066;
  assign new_P2_U4177 = ~new_P2_R1110_U98 | ~new_P2_U3879;
  assign new_P2_U4178 = ~new_P2_R1077_U98 | ~new_P2_U3881;
  assign new_P2_U4179 = ~new_P2_R1095_U23 | ~new_P2_U3880;
  assign new_P2_U4180 = ~new_P2_R1143_U98 | ~new_P2_U3877;
  assign new_P2_U4181 = ~new_P2_R1161_U98 | ~new_P2_U3887;
  assign new_P2_U4182 = ~new_P2_R1131_U23 | ~new_P2_U3883;
  assign new_P2_U4183 = ~new_P2_R1200_U23 | ~new_P2_U3017;
  assign new_P2_U4184 = ~new_P2_U3320;
  assign new_P2_U4185 = ~new_P2_R1179_U23 | ~new_P2_U3026;
  assign new_P2_U4186 = ~new_P2_U3025 | ~new_P2_U3069;
  assign new_P2_U4187 = ~new_P2_U3407 | ~new_P2_U4060;
  assign new_P2_U4188 = ~new_P2_U3613 | ~new_P2_U4184;
  assign new_P2_U4189 = ~P2_REG0_REG_8_ | ~new_P2_U3022;
  assign new_P2_U4190 = ~P2_REG1_REG_8_ | ~new_P2_U3021;
  assign new_P2_U4191 = ~P2_REG2_REG_8_ | ~new_P2_U3020;
  assign new_P2_U4192 = ~new_P2_SUB_605_U12 | ~new_P2_U3019;
  assign new_P2_U4193 = ~new_P2_U3083;
  assign new_P2_U4194 = ~new_P2_U3033 | ~new_P2_U3070;
  assign new_P2_U4195 = ~new_P2_R1110_U18 | ~new_P2_U3879;
  assign new_P2_U4196 = ~new_P2_R1077_U18 | ~new_P2_U3881;
  assign new_P2_U4197 = ~new_P2_R1095_U109 | ~new_P2_U3880;
  assign new_P2_U4198 = ~new_P2_R1143_U18 | ~new_P2_U3877;
  assign new_P2_U4199 = ~new_P2_R1161_U18 | ~new_P2_U3887;
  assign new_P2_U4200 = ~new_P2_R1131_U109 | ~new_P2_U3883;
  assign new_P2_U4201 = ~new_P2_R1200_U109 | ~new_P2_U3017;
  assign new_P2_U4202 = ~new_P2_U3321;
  assign new_P2_U4203 = ~new_P2_R1179_U109 | ~new_P2_U3026;
  assign new_P2_U4204 = ~new_P2_U3025 | ~new_P2_U3083;
  assign new_P2_U4205 = ~new_P2_U3410 | ~new_P2_U4060;
  assign new_P2_U4206 = ~new_P2_U3617 | ~new_P2_U4202;
  assign new_P2_U4207 = ~P2_REG0_REG_9_ | ~new_P2_U3022;
  assign new_P2_U4208 = ~P2_REG1_REG_9_ | ~new_P2_U3021;
  assign new_P2_U4209 = ~P2_REG2_REG_9_ | ~new_P2_U3020;
  assign new_P2_U4210 = ~new_P2_SUB_605_U14 | ~new_P2_U3019;
  assign new_P2_U4211 = ~new_P2_U3082;
  assign new_P2_U4212 = ~new_P2_U3033 | ~new_P2_U3069;
  assign new_P2_U4213 = ~new_P2_R1110_U97 | ~new_P2_U3879;
  assign new_P2_U4214 = ~new_P2_R1077_U97 | ~new_P2_U3881;
  assign new_P2_U4215 = ~new_P2_R1095_U24 | ~new_P2_U3880;
  assign new_P2_U4216 = ~new_P2_R1143_U97 | ~new_P2_U3877;
  assign new_P2_U4217 = ~new_P2_R1161_U97 | ~new_P2_U3887;
  assign new_P2_U4218 = ~new_P2_R1131_U24 | ~new_P2_U3883;
  assign new_P2_U4219 = ~new_P2_R1200_U24 | ~new_P2_U3017;
  assign new_P2_U4220 = ~new_P2_U3322;
  assign new_P2_U4221 = ~new_P2_R1179_U24 | ~new_P2_U3026;
  assign new_P2_U4222 = ~new_P2_U3025 | ~new_P2_U3082;
  assign new_P2_U4223 = ~new_P2_U3413 | ~new_P2_U4060;
  assign new_P2_U4224 = ~new_P2_U3620 | ~new_P2_U4220;
  assign new_P2_U4225 = ~P2_REG0_REG_10_ | ~new_P2_U3022;
  assign new_P2_U4226 = ~P2_REG1_REG_10_ | ~new_P2_U3021;
  assign new_P2_U4227 = ~P2_REG2_REG_10_ | ~new_P2_U3020;
  assign new_P2_U4228 = ~new_P2_SUB_605_U13 | ~new_P2_U3019;
  assign new_P2_U4229 = ~new_P2_U3061;
  assign new_P2_U4230 = ~new_P2_U3033 | ~new_P2_U3083;
  assign new_P2_U4231 = ~new_P2_R1110_U96 | ~new_P2_U3879;
  assign new_P2_U4232 = ~new_P2_R1077_U96 | ~new_P2_U3881;
  assign new_P2_U4233 = ~new_P2_R1095_U108 | ~new_P2_U3880;
  assign new_P2_U4234 = ~new_P2_R1143_U96 | ~new_P2_U3877;
  assign new_P2_U4235 = ~new_P2_R1161_U96 | ~new_P2_U3887;
  assign new_P2_U4236 = ~new_P2_R1131_U108 | ~new_P2_U3883;
  assign new_P2_U4237 = ~new_P2_R1200_U108 | ~new_P2_U3017;
  assign new_P2_U4238 = ~new_P2_U3323;
  assign new_P2_U4239 = ~new_P2_R1179_U108 | ~new_P2_U3026;
  assign new_P2_U4240 = ~new_P2_U3025 | ~new_P2_U3061;
  assign new_P2_U4241 = ~new_P2_U3416 | ~new_P2_U4060;
  assign new_P2_U4242 = ~new_P2_U3623 | ~new_P2_U4238;
  assign new_P2_U4243 = ~P2_REG0_REG_11_ | ~new_P2_U3022;
  assign new_P2_U4244 = ~P2_REG1_REG_11_ | ~new_P2_U3021;
  assign new_P2_U4245 = ~P2_REG2_REG_11_ | ~new_P2_U3020;
  assign new_P2_U4246 = ~new_P2_SUB_605_U9 | ~new_P2_U3019;
  assign new_P2_U4247 = ~new_P2_U3062;
  assign new_P2_U4248 = ~new_P2_U3033 | ~new_P2_U3082;
  assign new_P2_U4249 = ~new_P2_R1110_U10 | ~new_P2_U3879;
  assign new_P2_U4250 = ~new_P2_R1077_U10 | ~new_P2_U3881;
  assign new_P2_U4251 = ~new_P2_R1095_U118 | ~new_P2_U3880;
  assign new_P2_U4252 = ~new_P2_R1143_U10 | ~new_P2_U3877;
  assign new_P2_U4253 = ~new_P2_R1161_U10 | ~new_P2_U3887;
  assign new_P2_U4254 = ~new_P2_R1131_U118 | ~new_P2_U3883;
  assign new_P2_U4255 = ~new_P2_R1200_U118 | ~new_P2_U3017;
  assign new_P2_U4256 = ~new_P2_U3324;
  assign new_P2_U4257 = ~new_P2_R1179_U118 | ~new_P2_U3026;
  assign new_P2_U4258 = ~new_P2_U3025 | ~new_P2_U3062;
  assign new_P2_U4259 = ~new_P2_U3419 | ~new_P2_U4060;
  assign new_P2_U4260 = ~new_P2_U3626 | ~new_P2_U4256;
  assign new_P2_U4261 = ~P2_REG0_REG_12_ | ~new_P2_U3022;
  assign new_P2_U4262 = ~P2_REG1_REG_12_ | ~new_P2_U3021;
  assign new_P2_U4263 = ~P2_REG2_REG_12_ | ~new_P2_U3020;
  assign new_P2_U4264 = ~new_P2_SUB_605_U24 | ~new_P2_U3019;
  assign new_P2_U4265 = ~new_P2_U3071;
  assign new_P2_U4266 = ~new_P2_U3033 | ~new_P2_U3061;
  assign new_P2_U4267 = ~new_P2_R1110_U114 | ~new_P2_U3879;
  assign new_P2_U4268 = ~new_P2_R1077_U114 | ~new_P2_U3881;
  assign new_P2_U4269 = ~new_P2_R1095_U17 | ~new_P2_U3880;
  assign new_P2_U4270 = ~new_P2_R1143_U114 | ~new_P2_U3877;
  assign new_P2_U4271 = ~new_P2_R1161_U114 | ~new_P2_U3887;
  assign new_P2_U4272 = ~new_P2_R1131_U17 | ~new_P2_U3883;
  assign new_P2_U4273 = ~new_P2_R1200_U17 | ~new_P2_U3017;
  assign new_P2_U4274 = ~new_P2_U3325;
  assign new_P2_U4275 = ~new_P2_R1179_U17 | ~new_P2_U3026;
  assign new_P2_U4276 = ~new_P2_U3025 | ~new_P2_U3071;
  assign new_P2_U4277 = ~new_P2_U3422 | ~new_P2_U4060;
  assign new_P2_U4278 = ~new_P2_U3629 | ~new_P2_U4274;
  assign new_P2_U4279 = ~P2_REG0_REG_13_ | ~new_P2_U3022;
  assign new_P2_U4280 = ~P2_REG1_REG_13_ | ~new_P2_U3021;
  assign new_P2_U4281 = ~P2_REG2_REG_13_ | ~new_P2_U3020;
  assign new_P2_U4282 = ~new_P2_SUB_605_U25 | ~new_P2_U3019;
  assign new_P2_U4283 = ~new_P2_U3079;
  assign new_P2_U4284 = ~new_P2_U3033 | ~new_P2_U3062;
  assign new_P2_U4285 = ~new_P2_R1110_U113 | ~new_P2_U3879;
  assign new_P2_U4286 = ~new_P2_R1077_U113 | ~new_P2_U3881;
  assign new_P2_U4287 = ~new_P2_R1095_U107 | ~new_P2_U3880;
  assign new_P2_U4288 = ~new_P2_R1143_U113 | ~new_P2_U3877;
  assign new_P2_U4289 = ~new_P2_R1161_U113 | ~new_P2_U3887;
  assign new_P2_U4290 = ~new_P2_R1131_U107 | ~new_P2_U3883;
  assign new_P2_U4291 = ~new_P2_R1200_U107 | ~new_P2_U3017;
  assign new_P2_U4292 = ~new_P2_U3326;
  assign new_P2_U4293 = ~new_P2_R1179_U107 | ~new_P2_U3026;
  assign new_P2_U4294 = ~new_P2_U3025 | ~new_P2_U3079;
  assign new_P2_U4295 = ~new_P2_U3425 | ~new_P2_U4060;
  assign new_P2_U4296 = ~new_P2_U3633 | ~new_P2_U4292;
  assign new_P2_U4297 = ~P2_REG0_REG_14_ | ~new_P2_U3022;
  assign new_P2_U4298 = ~P2_REG1_REG_14_ | ~new_P2_U3021;
  assign new_P2_U4299 = ~P2_REG2_REG_14_ | ~new_P2_U3020;
  assign new_P2_U4300 = ~new_P2_SUB_605_U31 | ~new_P2_U3019;
  assign new_P2_U4301 = ~new_P2_U3078;
  assign new_P2_U4302 = ~new_P2_U3033 | ~new_P2_U3071;
  assign new_P2_U4303 = ~new_P2_R1110_U11 | ~new_P2_U3879;
  assign new_P2_U4304 = ~new_P2_R1077_U11 | ~new_P2_U3881;
  assign new_P2_U4305 = ~new_P2_R1095_U106 | ~new_P2_U3880;
  assign new_P2_U4306 = ~new_P2_R1143_U11 | ~new_P2_U3877;
  assign new_P2_U4307 = ~new_P2_R1161_U11 | ~new_P2_U3887;
  assign new_P2_U4308 = ~new_P2_R1131_U106 | ~new_P2_U3883;
  assign new_P2_U4309 = ~new_P2_R1200_U106 | ~new_P2_U3017;
  assign new_P2_U4310 = ~new_P2_U3327;
  assign new_P2_U4311 = ~new_P2_R1179_U106 | ~new_P2_U3026;
  assign new_P2_U4312 = ~new_P2_U3025 | ~new_P2_U3078;
  assign new_P2_U4313 = ~new_P2_U3428 | ~new_P2_U4060;
  assign new_P2_U4314 = ~new_P2_U3637 | ~new_P2_U4310;
  assign new_P2_U4315 = ~P2_REG0_REG_15_ | ~new_P2_U3022;
  assign new_P2_U4316 = ~P2_REG1_REG_15_ | ~new_P2_U3021;
  assign new_P2_U4317 = ~P2_REG2_REG_15_ | ~new_P2_U3020;
  assign new_P2_U4318 = ~new_P2_SUB_605_U21 | ~new_P2_U3019;
  assign new_P2_U4319 = ~new_P2_U3073;
  assign new_P2_U4320 = ~new_P2_U3033 | ~new_P2_U3079;
  assign new_P2_U4321 = ~new_P2_R1110_U112 | ~new_P2_U3879;
  assign new_P2_U4322 = ~new_P2_R1077_U112 | ~new_P2_U3881;
  assign new_P2_U4323 = ~new_P2_R1095_U117 | ~new_P2_U3880;
  assign new_P2_U4324 = ~new_P2_R1143_U112 | ~new_P2_U3877;
  assign new_P2_U4325 = ~new_P2_R1161_U112 | ~new_P2_U3887;
  assign new_P2_U4326 = ~new_P2_R1131_U117 | ~new_P2_U3883;
  assign new_P2_U4327 = ~new_P2_R1200_U117 | ~new_P2_U3017;
  assign new_P2_U4328 = ~new_P2_U3328;
  assign new_P2_U4329 = ~new_P2_R1179_U117 | ~new_P2_U3026;
  assign new_P2_U4330 = ~new_P2_U3025 | ~new_P2_U3073;
  assign new_P2_U4331 = ~new_P2_U3431 | ~new_P2_U4060;
  assign new_P2_U4332 = ~new_P2_U3640 | ~new_P2_U4328;
  assign new_P2_U4333 = ~P2_REG0_REG_16_ | ~new_P2_U3022;
  assign new_P2_U4334 = ~P2_REG1_REG_16_ | ~new_P2_U3021;
  assign new_P2_U4335 = ~P2_REG2_REG_16_ | ~new_P2_U3020;
  assign new_P2_U4336 = ~new_P2_SUB_605_U7 | ~new_P2_U3019;
  assign new_P2_U4337 = ~new_P2_U3072;
  assign new_P2_U4338 = ~new_P2_U3033 | ~new_P2_U3078;
  assign new_P2_U4339 = ~new_P2_R1110_U111 | ~new_P2_U3879;
  assign new_P2_U4340 = ~new_P2_R1077_U111 | ~new_P2_U3881;
  assign new_P2_U4341 = ~new_P2_R1095_U116 | ~new_P2_U3880;
  assign new_P2_U4342 = ~new_P2_R1143_U111 | ~new_P2_U3877;
  assign new_P2_U4343 = ~new_P2_R1161_U111 | ~new_P2_U3887;
  assign new_P2_U4344 = ~new_P2_R1131_U116 | ~new_P2_U3883;
  assign new_P2_U4345 = ~new_P2_R1200_U116 | ~new_P2_U3017;
  assign new_P2_U4346 = ~new_P2_U3329;
  assign new_P2_U4347 = ~new_P2_R1179_U116 | ~new_P2_U3026;
  assign new_P2_U4348 = ~new_P2_U3025 | ~new_P2_U3072;
  assign new_P2_U4349 = ~new_P2_U3434 | ~new_P2_U4060;
  assign new_P2_U4350 = ~new_P2_U3643 | ~new_P2_U4346;
  assign new_P2_U4351 = ~P2_REG0_REG_17_ | ~new_P2_U3022;
  assign new_P2_U4352 = ~P2_REG1_REG_17_ | ~new_P2_U3021;
  assign new_P2_U4353 = ~P2_REG2_REG_17_ | ~new_P2_U3020;
  assign new_P2_U4354 = ~new_P2_SUB_605_U19 | ~new_P2_U3019;
  assign new_P2_U4355 = ~new_P2_U3068;
  assign new_P2_U4356 = ~new_P2_U3033 | ~new_P2_U3073;
  assign new_P2_U4357 = ~new_P2_R1110_U110 | ~new_P2_U3879;
  assign new_P2_U4358 = ~new_P2_R1077_U110 | ~new_P2_U3881;
  assign new_P2_U4359 = ~new_P2_R1095_U18 | ~new_P2_U3880;
  assign new_P2_U4360 = ~new_P2_R1143_U110 | ~new_P2_U3877;
  assign new_P2_U4361 = ~new_P2_R1161_U110 | ~new_P2_U3887;
  assign new_P2_U4362 = ~new_P2_R1131_U18 | ~new_P2_U3883;
  assign new_P2_U4363 = ~new_P2_R1200_U18 | ~new_P2_U3017;
  assign new_P2_U4364 = ~new_P2_U3330;
  assign new_P2_U4365 = ~new_P2_R1179_U18 | ~new_P2_U3026;
  assign new_P2_U4366 = ~new_P2_U3025 | ~new_P2_U3068;
  assign new_P2_U4367 = ~new_P2_U3437 | ~new_P2_U4060;
  assign new_P2_U4368 = ~new_P2_U3646 | ~new_P2_U4364;
  assign new_P2_U4369 = ~P2_REG0_REG_18_ | ~new_P2_U3022;
  assign new_P2_U4370 = ~P2_REG1_REG_18_ | ~new_P2_U3021;
  assign new_P2_U4371 = ~P2_REG2_REG_18_ | ~new_P2_U3020;
  assign new_P2_U4372 = ~new_P2_SUB_605_U11 | ~new_P2_U3019;
  assign new_P2_U4373 = ~new_P2_U3081;
  assign new_P2_U4374 = ~new_P2_U3033 | ~new_P2_U3072;
  assign new_P2_U4375 = ~new_P2_R1110_U12 | ~new_P2_U3879;
  assign new_P2_U4376 = ~new_P2_R1077_U12 | ~new_P2_U3881;
  assign new_P2_U4377 = ~new_P2_R1095_U105 | ~new_P2_U3880;
  assign new_P2_U4378 = ~new_P2_R1143_U12 | ~new_P2_U3877;
  assign new_P2_U4379 = ~new_P2_R1161_U12 | ~new_P2_U3887;
  assign new_P2_U4380 = ~new_P2_R1131_U105 | ~new_P2_U3883;
  assign new_P2_U4381 = ~new_P2_R1200_U105 | ~new_P2_U3017;
  assign new_P2_U4382 = ~new_P2_U3331;
  assign new_P2_U4383 = ~new_P2_R1179_U105 | ~new_P2_U3026;
  assign new_P2_U4384 = ~new_P2_U3025 | ~new_P2_U3081;
  assign new_P2_U4385 = ~new_P2_U3440 | ~new_P2_U4060;
  assign new_P2_U4386 = ~new_P2_U3650 | ~new_P2_U4382;
  assign new_P2_U4387 = ~P2_REG0_REG_19_ | ~new_P2_U3022;
  assign new_P2_U4388 = ~P2_REG1_REG_19_ | ~new_P2_U3021;
  assign new_P2_U4389 = ~P2_REG2_REG_19_ | ~new_P2_U3020;
  assign new_P2_U4390 = ~new_P2_SUB_605_U15 | ~new_P2_U3019;
  assign new_P2_U4391 = ~new_P2_U3080;
  assign new_P2_U4392 = ~new_P2_U3033 | ~new_P2_U3068;
  assign new_P2_U4393 = ~new_P2_R1110_U109 | ~new_P2_U3879;
  assign new_P2_U4394 = ~new_P2_R1077_U109 | ~new_P2_U3881;
  assign new_P2_U4395 = ~new_P2_R1095_U104 | ~new_P2_U3880;
  assign new_P2_U4396 = ~new_P2_R1143_U109 | ~new_P2_U3877;
  assign new_P2_U4397 = ~new_P2_R1161_U109 | ~new_P2_U3887;
  assign new_P2_U4398 = ~new_P2_R1131_U104 | ~new_P2_U3883;
  assign new_P2_U4399 = ~new_P2_R1200_U104 | ~new_P2_U3017;
  assign new_P2_U4400 = ~new_P2_U3332;
  assign new_P2_U4401 = ~new_P2_R1179_U104 | ~new_P2_U3026;
  assign new_P2_U4402 = ~new_P2_U3025 | ~new_P2_U3080;
  assign new_P2_U4403 = ~new_P2_U3443 | ~new_P2_U4060;
  assign new_P2_U4404 = ~new_P2_U3654 | ~new_P2_U4400;
  assign new_P2_U4405 = ~P2_REG2_REG_20_ | ~new_P2_U3020;
  assign new_P2_U4406 = ~P2_REG1_REG_20_ | ~new_P2_U3021;
  assign new_P2_U4407 = ~P2_REG0_REG_20_ | ~new_P2_U3022;
  assign new_P2_U4408 = ~new_P2_SUB_605_U20 | ~new_P2_U3019;
  assign new_P2_U4409 = ~new_P2_U3075;
  assign new_P2_U4410 = ~new_P2_U3033 | ~new_P2_U3081;
  assign new_P2_U4411 = ~new_P2_R1110_U108 | ~new_P2_U3879;
  assign new_P2_U4412 = ~new_P2_R1077_U108 | ~new_P2_U3881;
  assign new_P2_U4413 = ~new_P2_R1095_U103 | ~new_P2_U3880;
  assign new_P2_U4414 = ~new_P2_R1143_U108 | ~new_P2_U3877;
  assign new_P2_U4415 = ~new_P2_R1161_U108 | ~new_P2_U3887;
  assign new_P2_U4416 = ~new_P2_R1131_U103 | ~new_P2_U3883;
  assign new_P2_U4417 = ~new_P2_R1200_U103 | ~new_P2_U3017;
  assign new_P2_U4418 = ~new_P2_U3333;
  assign new_P2_U4419 = ~new_P2_R1179_U103 | ~new_P2_U3026;
  assign new_P2_U4420 = ~new_P2_U3025 | ~new_P2_U3075;
  assign new_P2_U4421 = ~new_P2_U3445 | ~new_P2_U4060;
  assign new_P2_U4422 = ~new_P2_U3658 | ~new_P2_U4418;
  assign new_P2_U4423 = ~P2_REG2_REG_21_ | ~new_P2_U3020;
  assign new_P2_U4424 = ~P2_REG1_REG_21_ | ~new_P2_U3021;
  assign new_P2_U4425 = ~P2_REG0_REG_21_ | ~new_P2_U3022;
  assign new_P2_U4426 = ~new_P2_SUB_605_U28 | ~new_P2_U3019;
  assign new_P2_U4427 = ~new_P2_U3074;
  assign new_P2_U4428 = ~new_P2_U3033 | ~new_P2_U3080;
  assign new_P2_U4429 = ~new_P2_R1110_U13 | ~new_P2_U3879;
  assign new_P2_U4430 = ~new_P2_R1077_U13 | ~new_P2_U3881;
  assign new_P2_U4431 = ~new_P2_R1095_U101 | ~new_P2_U3880;
  assign new_P2_U4432 = ~new_P2_R1143_U13 | ~new_P2_U3877;
  assign new_P2_U4433 = ~new_P2_R1161_U13 | ~new_P2_U3887;
  assign new_P2_U4434 = ~new_P2_R1131_U101 | ~new_P2_U3883;
  assign new_P2_U4435 = ~new_P2_R1200_U101 | ~new_P2_U3017;
  assign new_P2_U4436 = ~new_P2_U3335;
  assign new_P2_U4437 = ~new_P2_R1179_U101 | ~new_P2_U3026;
  assign new_P2_U4438 = ~new_P2_U3025 | ~new_P2_U3074;
  assign new_P2_U4439 = ~new_P2_U3903 | ~new_P2_U4060;
  assign new_P2_U4440 = ~new_P2_U3662 | ~new_P2_U4436;
  assign new_P2_U4441 = ~P2_REG2_REG_22_ | ~new_P2_U3020;
  assign new_P2_U4442 = ~P2_REG1_REG_22_ | ~new_P2_U3021;
  assign new_P2_U4443 = ~P2_REG0_REG_22_ | ~new_P2_U3022;
  assign new_P2_U4444 = ~new_P2_SUB_605_U17 | ~new_P2_U3019;
  assign new_P2_U4445 = ~new_P2_U3060;
  assign new_P2_U4446 = ~new_P2_U3033 | ~new_P2_U3075;
  assign new_P2_U4447 = ~new_P2_R1110_U14 | ~new_P2_U3879;
  assign new_P2_U4448 = ~new_P2_R1077_U14 | ~new_P2_U3881;
  assign new_P2_U4449 = ~new_P2_R1095_U115 | ~new_P2_U3880;
  assign new_P2_U4450 = ~new_P2_R1143_U14 | ~new_P2_U3877;
  assign new_P2_U4451 = ~new_P2_R1161_U14 | ~new_P2_U3887;
  assign new_P2_U4452 = ~new_P2_R1131_U115 | ~new_P2_U3883;
  assign new_P2_U4453 = ~new_P2_R1200_U115 | ~new_P2_U3017;
  assign new_P2_U4454 = ~new_P2_U3337;
  assign new_P2_U4455 = ~new_P2_R1179_U115 | ~new_P2_U3026;
  assign new_P2_U4456 = ~new_P2_U3025 | ~new_P2_U3060;
  assign new_P2_U4457 = ~new_P2_U3902 | ~new_P2_U4060;
  assign new_P2_U4458 = ~new_P2_U3665 | ~new_P2_U4454;
  assign new_P2_U4459 = ~P2_REG2_REG_23_ | ~new_P2_U3020;
  assign new_P2_U4460 = ~P2_REG1_REG_23_ | ~new_P2_U3021;
  assign new_P2_U4461 = ~P2_REG0_REG_23_ | ~new_P2_U3022;
  assign new_P2_U4462 = ~new_P2_SUB_605_U6 | ~new_P2_U3019;
  assign new_P2_U4463 = ~new_P2_U3065;
  assign new_P2_U4464 = ~new_P2_U3033 | ~new_P2_U3074;
  assign new_P2_U4465 = ~new_P2_R1110_U107 | ~new_P2_U3879;
  assign new_P2_U4466 = ~new_P2_R1077_U107 | ~new_P2_U3881;
  assign new_P2_U4467 = ~new_P2_R1095_U114 | ~new_P2_U3880;
  assign new_P2_U4468 = ~new_P2_R1143_U107 | ~new_P2_U3877;
  assign new_P2_U4469 = ~new_P2_R1161_U107 | ~new_P2_U3887;
  assign new_P2_U4470 = ~new_P2_R1131_U114 | ~new_P2_U3883;
  assign new_P2_U4471 = ~new_P2_R1200_U114 | ~new_P2_U3017;
  assign new_P2_U4472 = ~new_P2_U3339;
  assign new_P2_U4473 = ~new_P2_R1179_U114 | ~new_P2_U3026;
  assign new_P2_U4474 = ~new_P2_U3025 | ~new_P2_U3065;
  assign new_P2_U4475 = ~new_P2_U3901 | ~new_P2_U4060;
  assign new_P2_U4476 = ~new_P2_U3668 | ~new_P2_U4472;
  assign new_P2_U4477 = ~P2_REG2_REG_24_ | ~new_P2_U3020;
  assign new_P2_U4478 = ~P2_REG1_REG_24_ | ~new_P2_U3021;
  assign new_P2_U4479 = ~P2_REG0_REG_24_ | ~new_P2_U3022;
  assign new_P2_U4480 = ~new_P2_SUB_605_U10 | ~new_P2_U3019;
  assign new_P2_U4481 = ~new_P2_U3064;
  assign new_P2_U4482 = ~new_P2_U3033 | ~new_P2_U3060;
  assign new_P2_U4483 = ~new_P2_R1110_U106 | ~new_P2_U3879;
  assign new_P2_U4484 = ~new_P2_R1077_U106 | ~new_P2_U3881;
  assign new_P2_U4485 = ~new_P2_R1095_U19 | ~new_P2_U3880;
  assign new_P2_U4486 = ~new_P2_R1143_U106 | ~new_P2_U3877;
  assign new_P2_U4487 = ~new_P2_R1161_U106 | ~new_P2_U3887;
  assign new_P2_U4488 = ~new_P2_R1131_U19 | ~new_P2_U3883;
  assign new_P2_U4489 = ~new_P2_R1200_U19 | ~new_P2_U3017;
  assign new_P2_U4490 = ~new_P2_U3341;
  assign new_P2_U4491 = ~new_P2_R1179_U19 | ~new_P2_U3026;
  assign new_P2_U4492 = ~new_P2_U3025 | ~new_P2_U3064;
  assign new_P2_U4493 = ~new_P2_U3900 | ~new_P2_U4060;
  assign new_P2_U4494 = ~new_P2_U3671 | ~new_P2_U4490;
  assign new_P2_U4495 = ~P2_REG2_REG_25_ | ~new_P2_U3020;
  assign new_P2_U4496 = ~P2_REG1_REG_25_ | ~new_P2_U3021;
  assign new_P2_U4497 = ~P2_REG0_REG_25_ | ~new_P2_U3022;
  assign new_P2_U4498 = ~new_P2_SUB_605_U16 | ~new_P2_U3019;
  assign new_P2_U4499 = ~new_P2_U3057;
  assign new_P2_U4500 = ~new_P2_U3033 | ~new_P2_U3065;
  assign new_P2_U4501 = ~new_P2_R1110_U105 | ~new_P2_U3879;
  assign new_P2_U4502 = ~new_P2_R1077_U105 | ~new_P2_U3881;
  assign new_P2_U4503 = ~new_P2_R1095_U100 | ~new_P2_U3880;
  assign new_P2_U4504 = ~new_P2_R1143_U105 | ~new_P2_U3877;
  assign new_P2_U4505 = ~new_P2_R1161_U105 | ~new_P2_U3887;
  assign new_P2_U4506 = ~new_P2_R1131_U100 | ~new_P2_U3883;
  assign new_P2_U4507 = ~new_P2_R1200_U100 | ~new_P2_U3017;
  assign new_P2_U4508 = ~new_P2_U3343;
  assign new_P2_U4509 = ~new_P2_R1179_U100 | ~new_P2_U3026;
  assign new_P2_U4510 = ~new_P2_U3025 | ~new_P2_U3057;
  assign new_P2_U4511 = ~new_P2_U3899 | ~new_P2_U4060;
  assign new_P2_U4512 = ~new_P2_U3675 | ~new_P2_U4508;
  assign new_P2_U4513 = ~P2_REG2_REG_26_ | ~new_P2_U3020;
  assign new_P2_U4514 = ~P2_REG1_REG_26_ | ~new_P2_U3021;
  assign new_P2_U4515 = ~P2_REG0_REG_26_ | ~new_P2_U3022;
  assign new_P2_U4516 = ~new_P2_SUB_605_U27 | ~new_P2_U3019;
  assign new_P2_U4517 = ~new_P2_U3056;
  assign new_P2_U4518 = ~new_P2_U3033 | ~new_P2_U3064;
  assign new_P2_U4519 = ~new_P2_R1110_U104 | ~new_P2_U3879;
  assign new_P2_U4520 = ~new_P2_R1077_U104 | ~new_P2_U3881;
  assign new_P2_U4521 = ~new_P2_R1095_U99 | ~new_P2_U3880;
  assign new_P2_U4522 = ~new_P2_R1143_U104 | ~new_P2_U3877;
  assign new_P2_U4523 = ~new_P2_R1161_U104 | ~new_P2_U3887;
  assign new_P2_U4524 = ~new_P2_R1131_U99 | ~new_P2_U3883;
  assign new_P2_U4525 = ~new_P2_R1200_U99 | ~new_P2_U3017;
  assign new_P2_U4526 = ~new_P2_U3345;
  assign new_P2_U4527 = ~new_P2_R1179_U99 | ~new_P2_U3026;
  assign new_P2_U4528 = ~new_P2_U3025 | ~new_P2_U3056;
  assign new_P2_U4529 = ~new_P2_U3898 | ~new_P2_U4060;
  assign new_P2_U4530 = ~new_P2_U3679 | ~new_P2_U4526;
  assign new_P2_U4531 = ~P2_REG2_REG_27_ | ~new_P2_U3020;
  assign new_P2_U4532 = ~P2_REG1_REG_27_ | ~new_P2_U3021;
  assign new_P2_U4533 = ~P2_REG0_REG_27_ | ~new_P2_U3022;
  assign new_P2_U4534 = ~new_P2_SUB_605_U23 | ~new_P2_U3019;
  assign new_P2_U4535 = ~new_P2_U3052;
  assign new_P2_U4536 = ~new_P2_U3033 | ~new_P2_U3057;
  assign new_P2_U4537 = ~new_P2_R1110_U15 | ~new_P2_U3879;
  assign new_P2_U4538 = ~new_P2_R1077_U15 | ~new_P2_U3881;
  assign new_P2_U4539 = ~new_P2_R1095_U113 | ~new_P2_U3880;
  assign new_P2_U4540 = ~new_P2_R1143_U15 | ~new_P2_U3877;
  assign new_P2_U4541 = ~new_P2_R1161_U15 | ~new_P2_U3887;
  assign new_P2_U4542 = ~new_P2_R1131_U113 | ~new_P2_U3883;
  assign new_P2_U4543 = ~new_P2_R1200_U113 | ~new_P2_U3017;
  assign new_P2_U4544 = ~new_P2_U3347;
  assign new_P2_U4545 = ~new_P2_R1179_U113 | ~new_P2_U3026;
  assign new_P2_U4546 = ~new_P2_U3025 | ~new_P2_U3052;
  assign new_P2_U4547 = ~new_P2_U3897 | ~new_P2_U4060;
  assign new_P2_U4548 = ~new_P2_U3683 | ~new_P2_U4544;
  assign new_P2_U4549 = ~P2_REG2_REG_28_ | ~new_P2_U3020;
  assign new_P2_U4550 = ~P2_REG1_REG_28_ | ~new_P2_U3021;
  assign new_P2_U4551 = ~P2_REG0_REG_28_ | ~new_P2_U3022;
  assign new_P2_U4552 = ~new_P2_SUB_605_U29 | ~new_P2_U3019;
  assign new_P2_U4553 = ~new_P2_U3053;
  assign new_P2_U4554 = ~new_P2_U3033 | ~new_P2_U3056;
  assign new_P2_U4555 = ~new_P2_R1110_U103 | ~new_P2_U3879;
  assign new_P2_U4556 = ~new_P2_R1077_U103 | ~new_P2_U3881;
  assign new_P2_U4557 = ~new_P2_R1095_U20 | ~new_P2_U3880;
  assign new_P2_U4558 = ~new_P2_R1143_U103 | ~new_P2_U3877;
  assign new_P2_U4559 = ~new_P2_R1161_U103 | ~new_P2_U3887;
  assign new_P2_U4560 = ~new_P2_R1131_U20 | ~new_P2_U3883;
  assign new_P2_U4561 = ~new_P2_R1200_U20 | ~new_P2_U3017;
  assign new_P2_U4562 = ~new_P2_U3349;
  assign new_P2_U4563 = ~new_P2_R1179_U20 | ~new_P2_U3026;
  assign new_P2_U4564 = ~new_P2_U3025 | ~new_P2_U3053;
  assign new_P2_U4565 = ~new_P2_U3896 | ~new_P2_U4060;
  assign new_P2_U4566 = ~new_P2_U3687 | ~new_P2_U4562;
  assign new_P2_U4567 = ~new_P2_SUB_605_U94 | ~new_P2_U3019;
  assign new_P2_U4568 = ~P2_REG2_REG_29_ | ~new_P2_U3020;
  assign new_P2_U4569 = ~P2_REG1_REG_29_ | ~new_P2_U3021;
  assign new_P2_U4570 = ~P2_REG0_REG_29_ | ~new_P2_U3022;
  assign new_P2_U4571 = ~new_P2_U3054;
  assign new_P2_U4572 = ~new_P2_U3033 | ~new_P2_U3052;
  assign new_P2_U4573 = ~new_P2_R1110_U102 | ~new_P2_U3879;
  assign new_P2_U4574 = ~new_P2_R1077_U102 | ~new_P2_U3881;
  assign new_P2_U4575 = ~new_P2_R1095_U98 | ~new_P2_U3880;
  assign new_P2_U4576 = ~new_P2_R1143_U102 | ~new_P2_U3877;
  assign new_P2_U4577 = ~new_P2_R1161_U102 | ~new_P2_U3887;
  assign new_P2_U4578 = ~new_P2_R1131_U98 | ~new_P2_U3883;
  assign new_P2_U4579 = ~new_P2_R1200_U98 | ~new_P2_U3017;
  assign new_P2_U4580 = ~new_P2_U3351;
  assign new_P2_U4581 = ~new_P2_R1179_U98 | ~new_P2_U3026;
  assign new_P2_U4582 = ~new_P2_U3025 | ~new_P2_U3054;
  assign new_P2_U4583 = ~new_P2_U3895 | ~new_P2_U4060;
  assign new_P2_U4584 = ~new_P2_U3691 | ~new_P2_U4580;
  assign new_P2_U4585 = ~P2_REG2_REG_30_ | ~new_P2_U3020;
  assign new_P2_U4586 = ~P2_REG1_REG_30_ | ~new_P2_U3021;
  assign new_P2_U4587 = ~P2_REG0_REG_30_ | ~new_P2_U3022;
  assign new_P2_U4588 = ~new_P2_SUB_605_U94 | ~new_P2_U3019;
  assign new_P2_U4589 = ~new_P2_U3058;
  assign new_P2_U4590 = ~new_P2_U3888 | ~new_P2_U3298;
  assign new_P2_U4591 = ~new_P2_U3829 | ~new_P2_U4590;
  assign new_P2_U4592 = ~new_P2_U3058 | ~new_P2_U4591 | ~new_P2_U3907;
  assign new_P2_U4593 = ~new_P2_U3033 | ~new_P2_U3053;
  assign new_P2_U4594 = ~new_P2_R1110_U101 | ~new_P2_U3879;
  assign new_P2_U4595 = ~new_P2_R1077_U101 | ~new_P2_U3881;
  assign new_P2_U4596 = ~new_P2_R1095_U21 | ~new_P2_U3880;
  assign new_P2_U4597 = ~new_P2_R1143_U101 | ~new_P2_U3877;
  assign new_P2_U4598 = ~new_P2_R1161_U101 | ~new_P2_U3887;
  assign new_P2_U4599 = ~new_P2_R1131_U21 | ~new_P2_U3883;
  assign new_P2_U4600 = ~new_P2_R1200_U21 | ~new_P2_U3017;
  assign new_P2_U4601 = ~new_P2_U3354;
  assign new_P2_U4602 = ~new_P2_R1179_U21 | ~new_P2_U3026;
  assign new_P2_U4603 = ~new_P2_U3904 | ~new_P2_U4060;
  assign new_P2_U4604 = ~new_P2_U3695 | ~new_P2_U4601;
  assign new_P2_U4605 = ~new_P2_SUB_605_U94 | ~new_P2_U3019;
  assign new_P2_U4606 = ~P2_REG2_REG_31_ | ~new_P2_U3020;
  assign new_P2_U4607 = ~P2_REG1_REG_31_ | ~new_P2_U3021;
  assign new_P2_U4608 = ~P2_REG0_REG_31_ | ~new_P2_U3022;
  assign new_P2_U4609 = ~new_P2_U3055;
  assign new_P2_U4610 = ~new_P2_U3869 | ~new_P2_U4060;
  assign new_P2_U4611 = ~new_P2_U3361 | ~new_P2_U4610;
  assign new_P2_U4612 = ~new_P2_U3868 | ~new_P2_U4060;
  assign new_P2_U4613 = ~new_P2_U3361 | ~new_P2_U4612;
  assign new_P2_U4614 = ~new_P2_U3302 | ~new_P2_U5637 | ~new_P2_U5636;
  assign new_P2_U4615 = ~new_P2_U3884 | ~new_P2_U3367;
  assign new_P2_U4616 = ~new_P2_U3048 | ~new_P2_U4615;
  assign new_P2_U4617 = ~new_P2_U3047 | ~new_P2_U4614;
  assign new_P2_U4618 = ~new_P2_U4617 | ~new_P2_U4616;
  assign new_P2_U4619 = ~new_P2_U5452 | ~new_P2_U3379;
  assign new_P2_U4620 = ~new_P2_U3830 | ~new_P2_U4619 | ~new_P2_U3380;
  assign new_P2_U4621 = ~new_P2_U3048 | ~new_P2_U4620;
  assign new_P2_U4622 = ~new_P2_U3047 | ~new_P2_U4615;
  assign new_P2_U4623 = ~new_P2_U4622 | ~new_P2_U4621 | ~new_P2_U3360;
  assign new_P2_U4624 = ~new_P2_U3365;
  assign new_P2_U4625 = ~new_P2_U3034 | ~new_P2_U3077;
  assign new_P2_U4626 = ~new_P2_U3030 | ~new_P2_R1179_U25;
  assign new_P2_U4627 = ~new_P2_U3029 | ~new_P2_U3387;
  assign new_P2_U4628 = ~new_P2_U3028 | ~P2_REG3_REG_0_;
  assign new_P2_U4629 = ~new_P2_U3034 | ~new_P2_U3067;
  assign new_P2_U4630 = ~new_P2_U3030 | ~new_P2_R1179_U102;
  assign new_P2_U4631 = ~new_P2_U3029 | ~new_P2_U3392;
  assign new_P2_U4632 = ~new_P2_U3028 | ~P2_REG3_REG_1_;
  assign new_P2_U4633 = ~new_P2_U3034 | ~new_P2_U3063;
  assign new_P2_U4634 = ~new_P2_U3030 | ~new_P2_R1179_U112;
  assign new_P2_U4635 = ~new_P2_U3029 | ~new_P2_U3395;
  assign new_P2_U4636 = ~new_P2_U3028 | ~P2_REG3_REG_2_;
  assign new_P2_U4637 = ~new_P2_U3034 | ~new_P2_U3059;
  assign new_P2_U4638 = ~new_P2_U3030 | ~new_P2_R1179_U22;
  assign new_P2_U4639 = ~new_P2_U3029 | ~new_P2_U3398;
  assign new_P2_U4640 = ~new_P2_U3028 | ~new_P2_SUB_605_U26;
  assign new_P2_U4641 = ~new_P2_U3034 | ~new_P2_U3066;
  assign new_P2_U4642 = ~new_P2_U3030 | ~new_P2_R1179_U111;
  assign new_P2_U4643 = ~new_P2_U3029 | ~new_P2_U3401;
  assign new_P2_U4644 = ~new_P2_U3028 | ~new_P2_SUB_605_U30;
  assign new_P2_U4645 = ~new_P2_U3034 | ~new_P2_U3070;
  assign new_P2_U4646 = ~new_P2_U3030 | ~new_P2_R1179_U110;
  assign new_P2_U4647 = ~new_P2_U3029 | ~new_P2_U3404;
  assign new_P2_U4648 = ~new_P2_U3028 | ~new_P2_SUB_605_U22;
  assign new_P2_U4649 = ~new_P2_U3034 | ~new_P2_U3069;
  assign new_P2_U4650 = ~new_P2_U3030 | ~new_P2_R1179_U23;
  assign new_P2_U4651 = ~new_P2_U3029 | ~new_P2_U3407;
  assign new_P2_U4652 = ~new_P2_U3028 | ~new_P2_SUB_605_U8;
  assign new_P2_U4653 = ~new_P2_U3034 | ~new_P2_U3083;
  assign new_P2_U4654 = ~new_P2_U3030 | ~new_P2_R1179_U109;
  assign new_P2_U4655 = ~new_P2_U3029 | ~new_P2_U3410;
  assign new_P2_U4656 = ~new_P2_U3028 | ~new_P2_SUB_605_U18;
  assign new_P2_U4657 = ~new_P2_U3034 | ~new_P2_U3082;
  assign new_P2_U4658 = ~new_P2_U3030 | ~new_P2_R1179_U24;
  assign new_P2_U4659 = ~new_P2_U3029 | ~new_P2_U3413;
  assign new_P2_U4660 = ~new_P2_U3028 | ~new_P2_SUB_605_U12;
  assign new_P2_U4661 = ~new_P2_U3034 | ~new_P2_U3061;
  assign new_P2_U4662 = ~new_P2_U3030 | ~new_P2_R1179_U108;
  assign new_P2_U4663 = ~new_P2_U3029 | ~new_P2_U3416;
  assign new_P2_U4664 = ~new_P2_U3028 | ~new_P2_SUB_605_U14;
  assign new_P2_U4665 = ~new_P2_U3034 | ~new_P2_U3062;
  assign new_P2_U4666 = ~new_P2_U3030 | ~new_P2_R1179_U118;
  assign new_P2_U4667 = ~new_P2_U3029 | ~new_P2_U3419;
  assign new_P2_U4668 = ~new_P2_U3028 | ~new_P2_SUB_605_U13;
  assign new_P2_U4669 = ~new_P2_U3034 | ~new_P2_U3071;
  assign new_P2_U4670 = ~new_P2_U3030 | ~new_P2_R1179_U17;
  assign new_P2_U4671 = ~new_P2_U3029 | ~new_P2_U3422;
  assign new_P2_U4672 = ~new_P2_U3028 | ~new_P2_SUB_605_U9;
  assign new_P2_U4673 = ~new_P2_U3034 | ~new_P2_U3079;
  assign new_P2_U4674 = ~new_P2_U3030 | ~new_P2_R1179_U107;
  assign new_P2_U4675 = ~new_P2_U3029 | ~new_P2_U3425;
  assign new_P2_U4676 = ~new_P2_U3028 | ~new_P2_SUB_605_U24;
  assign new_P2_U4677 = ~new_P2_U3034 | ~new_P2_U3078;
  assign new_P2_U4678 = ~new_P2_U3030 | ~new_P2_R1179_U106;
  assign new_P2_U4679 = ~new_P2_U3029 | ~new_P2_U3428;
  assign new_P2_U4680 = ~new_P2_U3028 | ~new_P2_SUB_605_U25;
  assign new_P2_U4681 = ~new_P2_U3034 | ~new_P2_U3073;
  assign new_P2_U4682 = ~new_P2_U3030 | ~new_P2_R1179_U117;
  assign new_P2_U4683 = ~new_P2_U3029 | ~new_P2_U3431;
  assign new_P2_U4684 = ~new_P2_U3028 | ~new_P2_SUB_605_U31;
  assign new_P2_U4685 = ~new_P2_U3034 | ~new_P2_U3072;
  assign new_P2_U4686 = ~new_P2_U3030 | ~new_P2_R1179_U116;
  assign new_P2_U4687 = ~new_P2_U3029 | ~new_P2_U3434;
  assign new_P2_U4688 = ~new_P2_U3028 | ~new_P2_SUB_605_U21;
  assign new_P2_U4689 = ~new_P2_U3034 | ~new_P2_U3068;
  assign new_P2_U4690 = ~new_P2_U3030 | ~new_P2_R1179_U18;
  assign new_P2_U4691 = ~new_P2_U3029 | ~new_P2_U3437;
  assign new_P2_U4692 = ~new_P2_U3028 | ~new_P2_SUB_605_U7;
  assign new_P2_U4693 = ~new_P2_U3034 | ~new_P2_U3081;
  assign new_P2_U4694 = ~new_P2_U3030 | ~new_P2_R1179_U105;
  assign new_P2_U4695 = ~new_P2_U3029 | ~new_P2_U3440;
  assign new_P2_U4696 = ~new_P2_U3028 | ~new_P2_SUB_605_U19;
  assign new_P2_U4697 = ~new_P2_U3034 | ~new_P2_U3080;
  assign new_P2_U4698 = ~new_P2_U3030 | ~new_P2_R1179_U104;
  assign new_P2_U4699 = ~new_P2_U3029 | ~new_P2_U3443;
  assign new_P2_U4700 = ~new_P2_U3028 | ~new_P2_SUB_605_U11;
  assign new_P2_U4701 = ~new_P2_U3034 | ~new_P2_U3075;
  assign new_P2_U4702 = ~new_P2_U3030 | ~new_P2_R1179_U103;
  assign new_P2_U4703 = ~new_P2_U3029 | ~new_P2_U3445;
  assign new_P2_U4704 = ~new_P2_U3028 | ~new_P2_SUB_605_U15;
  assign new_P2_U4705 = ~new_P2_U3034 | ~new_P2_U3074;
  assign new_P2_U4706 = ~new_P2_U3030 | ~new_P2_R1179_U101;
  assign new_P2_U4707 = ~new_P2_U3029 | ~new_P2_U3903;
  assign new_P2_U4708 = ~new_P2_U3028 | ~new_P2_SUB_605_U20;
  assign new_P2_U4709 = ~new_P2_U3034 | ~new_P2_U3060;
  assign new_P2_U4710 = ~new_P2_U3030 | ~new_P2_R1179_U115;
  assign new_P2_U4711 = ~new_P2_U3029 | ~new_P2_U3902;
  assign new_P2_U4712 = ~new_P2_U3028 | ~new_P2_SUB_605_U28;
  assign new_P2_U4713 = ~new_P2_U3034 | ~new_P2_U3065;
  assign new_P2_U4714 = ~new_P2_U3030 | ~new_P2_R1179_U114;
  assign new_P2_U4715 = ~new_P2_U3029 | ~new_P2_U3901;
  assign new_P2_U4716 = ~new_P2_U3028 | ~new_P2_SUB_605_U17;
  assign new_P2_U4717 = ~new_P2_U3034 | ~new_P2_U3064;
  assign new_P2_U4718 = ~new_P2_U3030 | ~new_P2_R1179_U19;
  assign new_P2_U4719 = ~new_P2_U3029 | ~new_P2_U3900;
  assign new_P2_U4720 = ~new_P2_U3028 | ~new_P2_SUB_605_U6;
  assign new_P2_U4721 = ~new_P2_U3034 | ~new_P2_U3057;
  assign new_P2_U4722 = ~new_P2_U3030 | ~new_P2_R1179_U100;
  assign new_P2_U4723 = ~new_P2_U3029 | ~new_P2_U3899;
  assign new_P2_U4724 = ~new_P2_U3028 | ~new_P2_SUB_605_U10;
  assign new_P2_U4725 = ~new_P2_U3034 | ~new_P2_U3056;
  assign new_P2_U4726 = ~new_P2_U3030 | ~new_P2_R1179_U99;
  assign new_P2_U4727 = ~new_P2_U3029 | ~new_P2_U3898;
  assign new_P2_U4728 = ~new_P2_U3028 | ~new_P2_SUB_605_U16;
  assign new_P2_U4729 = ~new_P2_U3034 | ~new_P2_U3052;
  assign new_P2_U4730 = ~new_P2_U3030 | ~new_P2_R1179_U113;
  assign new_P2_U4731 = ~new_P2_U3029 | ~new_P2_U3897;
  assign new_P2_U4732 = ~new_P2_U3028 | ~new_P2_SUB_605_U27;
  assign new_P2_U4733 = ~new_P2_U3034 | ~new_P2_U3053;
  assign new_P2_U4734 = ~new_P2_U3030 | ~new_P2_R1179_U20;
  assign new_P2_U4735 = ~new_P2_U3029 | ~new_P2_U3896;
  assign new_P2_U4736 = ~new_P2_U3028 | ~new_P2_SUB_605_U23;
  assign new_P2_U4737 = ~new_P2_U3034 | ~new_P2_U3054;
  assign new_P2_U4738 = ~new_P2_U3030 | ~new_P2_R1179_U98;
  assign new_P2_U4739 = ~new_P2_U3029 | ~new_P2_U3895;
  assign new_P2_U4740 = ~new_P2_U3028 | ~new_P2_SUB_605_U29;
  assign new_P2_U4741 = ~new_P2_U3030 | ~new_P2_R1179_U21;
  assign new_P2_U4742 = ~new_P2_U3029 | ~new_P2_U3904;
  assign new_P2_U4743 = ~new_P2_U3028 | ~new_P2_SUB_605_U94;
  assign new_P2_U4744 = ~new_P2_U3028 | ~new_P2_SUB_605_U94;
  assign new_P2_U4745 = ~new_P2_U3912 | ~new_P2_U3908;
  assign new_P2_U4746 = ~new_P2_U3029 | ~new_P2_U3869;
  assign new_P2_U4747 = ~P2_REG2_REG_30_ | ~new_P2_U3358;
  assign new_P2_U4748 = ~new_P2_U3029 | ~new_P2_U3868;
  assign new_P2_U4749 = ~P2_REG2_REG_31_ | ~new_P2_U3358;
  assign new_P2_U4750 = ~new_P2_U3702 | ~new_P2_U3703 | ~new_P2_U4624 | ~new_P2_U3359;
  assign new_P2_U4751 = ~new_P2_R1212_U6 | ~new_P2_U3040;
  assign new_P2_U4752 = ~new_P2_U3039 | ~new_P2_U3379;
  assign new_P2_U4753 = ~new_P2_R1209_U6 | ~new_P2_U3037;
  assign new_P2_U4754 = ~new_P2_U4753 | ~new_P2_U4752 | ~new_P2_U4751;
  assign new_P2_U4755 = ~new_P2_U3906 | ~new_P2_U5436;
  assign new_P2_U4756 = ~new_P2_U3366;
  assign new_P2_U4757 = ~new_P2_U3829 | ~new_P2_U3892;
  assign new_P2_U4758 = ~new_P2_R1054_U67 | ~new_P2_U3051;
  assign new_P2_U4759 = ~new_P2_U5764 | ~new_P2_U3379;
  assign new_P2_U4760 = ~new_P2_U3042 | ~new_P2_U4754;
  assign new_P2_U4761 = ~new_P2_U3041 | ~new_P2_R1212_U6;
  assign new_P2_U4762 = ~P2_REG3_REG_19_ | ~n2555;
  assign new_P2_U4763 = ~new_P2_U3038 | ~new_P2_R1209_U6;
  assign new_P2_U4764 = ~P2_ADDR_REG_19_ | ~new_P2_U4756;
  assign new_P2_U4765 = ~new_P2_R1212_U58 | ~new_P2_U3040;
  assign new_P2_U4766 = ~new_P2_U3039 | ~new_P2_U3442;
  assign new_P2_U4767 = ~new_P2_R1209_U58 | ~new_P2_U3037;
  assign new_P2_U4768 = ~new_P2_U4767 | ~new_P2_U4766 | ~new_P2_U4765;
  assign new_P2_U4769 = ~new_P2_R1054_U68 | ~new_P2_U3051;
  assign new_P2_U4770 = ~new_P2_U5764 | ~new_P2_U3442;
  assign new_P2_U4771 = ~new_P2_U3042 | ~new_P2_U4768;
  assign new_P2_U4772 = ~new_P2_R1212_U58 | ~new_P2_U3041;
  assign new_P2_U4773 = ~P2_REG3_REG_18_ | ~n2555;
  assign new_P2_U4774 = ~new_P2_R1209_U58 | ~new_P2_U3038;
  assign new_P2_U4775 = ~P2_ADDR_REG_18_ | ~new_P2_U4756;
  assign new_P2_U4776 = ~new_P2_R1212_U59 | ~new_P2_U3040;
  assign new_P2_U4777 = ~new_P2_U3039 | ~new_P2_U3439;
  assign new_P2_U4778 = ~new_P2_R1209_U59 | ~new_P2_U3037;
  assign new_P2_U4779 = ~new_P2_U4778 | ~new_P2_U4777 | ~new_P2_U4776;
  assign new_P2_U4780 = ~new_P2_R1054_U69 | ~new_P2_U3051;
  assign new_P2_U4781 = ~new_P2_U5764 | ~new_P2_U3439;
  assign new_P2_U4782 = ~new_P2_U3042 | ~new_P2_U4779;
  assign new_P2_U4783 = ~new_P2_R1212_U59 | ~new_P2_U3041;
  assign new_P2_U4784 = ~P2_REG3_REG_17_ | ~n2555;
  assign new_P2_U4785 = ~new_P2_R1209_U59 | ~new_P2_U3038;
  assign new_P2_U4786 = ~P2_ADDR_REG_17_ | ~new_P2_U4756;
  assign new_P2_U4787 = ~new_P2_R1212_U60 | ~new_P2_U3040;
  assign new_P2_U4788 = ~new_P2_U3039 | ~new_P2_U3436;
  assign new_P2_U4789 = ~new_P2_R1209_U60 | ~new_P2_U3037;
  assign new_P2_U4790 = ~new_P2_U4789 | ~new_P2_U4788 | ~new_P2_U4787;
  assign new_P2_U4791 = ~new_P2_R1054_U13 | ~new_P2_U3051;
  assign new_P2_U4792 = ~new_P2_U5764 | ~new_P2_U3436;
  assign new_P2_U4793 = ~new_P2_U3042 | ~new_P2_U4790;
  assign new_P2_U4794 = ~new_P2_R1212_U60 | ~new_P2_U3041;
  assign new_P2_U4795 = ~P2_REG3_REG_16_ | ~n2555;
  assign new_P2_U4796 = ~new_P2_R1209_U60 | ~new_P2_U3038;
  assign new_P2_U4797 = ~P2_ADDR_REG_16_ | ~new_P2_U4756;
  assign new_P2_U4798 = ~new_P2_R1212_U61 | ~new_P2_U3040;
  assign new_P2_U4799 = ~new_P2_U3039 | ~new_P2_U3433;
  assign new_P2_U4800 = ~new_P2_R1209_U61 | ~new_P2_U3037;
  assign new_P2_U4801 = ~new_P2_U4800 | ~new_P2_U4799 | ~new_P2_U4798;
  assign new_P2_U4802 = ~new_P2_R1054_U77 | ~new_P2_U3051;
  assign new_P2_U4803 = ~new_P2_U5764 | ~new_P2_U3433;
  assign new_P2_U4804 = ~new_P2_U3042 | ~new_P2_U4801;
  assign new_P2_U4805 = ~new_P2_R1212_U61 | ~new_P2_U3041;
  assign new_P2_U4806 = ~P2_REG3_REG_15_ | ~n2555;
  assign new_P2_U4807 = ~new_P2_R1209_U61 | ~new_P2_U3038;
  assign new_P2_U4808 = ~P2_ADDR_REG_15_ | ~new_P2_U4756;
  assign new_P2_U4809 = ~new_P2_R1212_U62 | ~new_P2_U3040;
  assign new_P2_U4810 = ~new_P2_U3039 | ~new_P2_U3430;
  assign new_P2_U4811 = ~new_P2_R1209_U62 | ~new_P2_U3037;
  assign new_P2_U4812 = ~new_P2_U4811 | ~new_P2_U4810 | ~new_P2_U4809;
  assign new_P2_U4813 = ~new_P2_R1054_U78 | ~new_P2_U3051;
  assign new_P2_U4814 = ~new_P2_U5764 | ~new_P2_U3430;
  assign new_P2_U4815 = ~new_P2_U3042 | ~new_P2_U4812;
  assign new_P2_U4816 = ~new_P2_R1212_U62 | ~new_P2_U3041;
  assign new_P2_U4817 = ~P2_REG3_REG_14_ | ~n2555;
  assign new_P2_U4818 = ~new_P2_R1209_U62 | ~new_P2_U3038;
  assign new_P2_U4819 = ~P2_ADDR_REG_14_ | ~new_P2_U4756;
  assign new_P2_U4820 = ~new_P2_R1212_U63 | ~new_P2_U3040;
  assign new_P2_U4821 = ~new_P2_U3039 | ~new_P2_U3427;
  assign new_P2_U4822 = ~new_P2_R1209_U63 | ~new_P2_U3037;
  assign new_P2_U4823 = ~new_P2_U4822 | ~new_P2_U4821 | ~new_P2_U4820;
  assign new_P2_U4824 = ~new_P2_R1054_U70 | ~new_P2_U3051;
  assign new_P2_U4825 = ~new_P2_U5764 | ~new_P2_U3427;
  assign new_P2_U4826 = ~new_P2_U3042 | ~new_P2_U4823;
  assign new_P2_U4827 = ~new_P2_R1212_U63 | ~new_P2_U3041;
  assign new_P2_U4828 = ~P2_REG3_REG_13_ | ~n2555;
  assign new_P2_U4829 = ~new_P2_R1209_U63 | ~new_P2_U3038;
  assign new_P2_U4830 = ~P2_ADDR_REG_13_ | ~new_P2_U4756;
  assign new_P2_U4831 = ~new_P2_R1212_U64 | ~new_P2_U3040;
  assign new_P2_U4832 = ~new_P2_U3039 | ~new_P2_U3424;
  assign new_P2_U4833 = ~new_P2_R1209_U64 | ~new_P2_U3037;
  assign new_P2_U4834 = ~new_P2_U4833 | ~new_P2_U4832 | ~new_P2_U4831;
  assign new_P2_U4835 = ~new_P2_R1054_U71 | ~new_P2_U3051;
  assign new_P2_U4836 = ~new_P2_U5764 | ~new_P2_U3424;
  assign new_P2_U4837 = ~new_P2_U3042 | ~new_P2_U4834;
  assign new_P2_U4838 = ~new_P2_R1212_U64 | ~new_P2_U3041;
  assign new_P2_U4839 = ~P2_REG3_REG_12_ | ~n2555;
  assign new_P2_U4840 = ~new_P2_R1209_U64 | ~new_P2_U3038;
  assign new_P2_U4841 = ~P2_ADDR_REG_12_ | ~new_P2_U4756;
  assign new_P2_U4842 = ~new_P2_R1212_U65 | ~new_P2_U3040;
  assign new_P2_U4843 = ~new_P2_U3039 | ~new_P2_U3421;
  assign new_P2_U4844 = ~new_P2_R1209_U65 | ~new_P2_U3037;
  assign new_P2_U4845 = ~new_P2_U4844 | ~new_P2_U4843 | ~new_P2_U4842;
  assign new_P2_U4846 = ~new_P2_R1054_U12 | ~new_P2_U3051;
  assign new_P2_U4847 = ~new_P2_U5764 | ~new_P2_U3421;
  assign new_P2_U4848 = ~new_P2_U3042 | ~new_P2_U4845;
  assign new_P2_U4849 = ~new_P2_R1212_U65 | ~new_P2_U3041;
  assign new_P2_U4850 = ~P2_REG3_REG_11_ | ~n2555;
  assign new_P2_U4851 = ~new_P2_R1209_U65 | ~new_P2_U3038;
  assign new_P2_U4852 = ~P2_ADDR_REG_11_ | ~new_P2_U4756;
  assign new_P2_U4853 = ~new_P2_R1212_U66 | ~new_P2_U3040;
  assign new_P2_U4854 = ~new_P2_U3039 | ~new_P2_U3418;
  assign new_P2_U4855 = ~new_P2_R1209_U66 | ~new_P2_U3037;
  assign new_P2_U4856 = ~new_P2_U4855 | ~new_P2_U4854 | ~new_P2_U4853;
  assign new_P2_U4857 = ~new_P2_R1054_U79 | ~new_P2_U3051;
  assign new_P2_U4858 = ~new_P2_U5764 | ~new_P2_U3418;
  assign new_P2_U4859 = ~new_P2_U3042 | ~new_P2_U4856;
  assign new_P2_U4860 = ~new_P2_R1212_U66 | ~new_P2_U3041;
  assign new_P2_U4861 = ~P2_REG3_REG_10_ | ~n2555;
  assign new_P2_U4862 = ~new_P2_R1209_U66 | ~new_P2_U3038;
  assign new_P2_U4863 = ~P2_ADDR_REG_10_ | ~new_P2_U4756;
  assign new_P2_U4864 = ~new_P2_R1212_U49 | ~new_P2_U3040;
  assign new_P2_U4865 = ~new_P2_U3039 | ~new_P2_U3415;
  assign new_P2_U4866 = ~new_P2_R1209_U49 | ~new_P2_U3037;
  assign new_P2_U4867 = ~new_P2_U4866 | ~new_P2_U4865 | ~new_P2_U4864;
  assign new_P2_U4868 = ~new_P2_R1054_U72 | ~new_P2_U3051;
  assign new_P2_U4869 = ~new_P2_U5764 | ~new_P2_U3415;
  assign new_P2_U4870 = ~new_P2_U3042 | ~new_P2_U4867;
  assign new_P2_U4871 = ~new_P2_R1212_U49 | ~new_P2_U3041;
  assign new_P2_U4872 = ~P2_REG3_REG_9_ | ~n2555;
  assign new_P2_U4873 = ~new_P2_R1209_U49 | ~new_P2_U3038;
  assign new_P2_U4874 = ~P2_ADDR_REG_9_ | ~new_P2_U4756;
  assign new_P2_U4875 = ~new_P2_R1212_U50 | ~new_P2_U3040;
  assign new_P2_U4876 = ~new_P2_U3039 | ~new_P2_U3412;
  assign new_P2_U4877 = ~new_P2_R1209_U50 | ~new_P2_U3037;
  assign new_P2_U4878 = ~new_P2_U4877 | ~new_P2_U4876 | ~new_P2_U4875;
  assign new_P2_U4879 = ~new_P2_R1054_U16 | ~new_P2_U3051;
  assign new_P2_U4880 = ~new_P2_U5764 | ~new_P2_U3412;
  assign new_P2_U4881 = ~new_P2_U3042 | ~new_P2_U4878;
  assign new_P2_U4882 = ~new_P2_R1212_U50 | ~new_P2_U3041;
  assign new_P2_U4883 = ~P2_REG3_REG_8_ | ~n2555;
  assign new_P2_U4884 = ~new_P2_R1209_U50 | ~new_P2_U3038;
  assign new_P2_U4885 = ~P2_ADDR_REG_8_ | ~new_P2_U4756;
  assign new_P2_U4886 = ~new_P2_R1212_U51 | ~new_P2_U3040;
  assign new_P2_U4887 = ~new_P2_U3039 | ~new_P2_U3409;
  assign new_P2_U4888 = ~new_P2_R1209_U51 | ~new_P2_U3037;
  assign new_P2_U4889 = ~new_P2_U4888 | ~new_P2_U4887 | ~new_P2_U4886;
  assign new_P2_U4890 = ~new_P2_R1054_U73 | ~new_P2_U3051;
  assign new_P2_U4891 = ~new_P2_U5764 | ~new_P2_U3409;
  assign new_P2_U4892 = ~new_P2_U3042 | ~new_P2_U4889;
  assign new_P2_U4893 = ~new_P2_R1212_U51 | ~new_P2_U3041;
  assign new_P2_U4894 = ~P2_REG3_REG_7_ | ~n2555;
  assign new_P2_U4895 = ~new_P2_R1209_U51 | ~new_P2_U3038;
  assign new_P2_U4896 = ~P2_ADDR_REG_7_ | ~new_P2_U4756;
  assign new_P2_U4897 = ~new_P2_R1212_U52 | ~new_P2_U3040;
  assign new_P2_U4898 = ~new_P2_U3039 | ~new_P2_U3406;
  assign new_P2_U4899 = ~new_P2_R1209_U52 | ~new_P2_U3037;
  assign new_P2_U4900 = ~new_P2_U4899 | ~new_P2_U4898 | ~new_P2_U4897;
  assign new_P2_U4901 = ~new_P2_R1054_U15 | ~new_P2_U3051;
  assign new_P2_U4902 = ~new_P2_U5764 | ~new_P2_U3406;
  assign new_P2_U4903 = ~new_P2_U3042 | ~new_P2_U4900;
  assign new_P2_U4904 = ~new_P2_R1212_U52 | ~new_P2_U3041;
  assign new_P2_U4905 = ~P2_REG3_REG_6_ | ~n2555;
  assign new_P2_U4906 = ~new_P2_R1209_U52 | ~new_P2_U3038;
  assign new_P2_U4907 = ~P2_ADDR_REG_6_ | ~new_P2_U4756;
  assign new_P2_U4908 = ~new_P2_R1212_U53 | ~new_P2_U3040;
  assign new_P2_U4909 = ~new_P2_U3039 | ~new_P2_U3403;
  assign new_P2_U4910 = ~new_P2_R1209_U53 | ~new_P2_U3037;
  assign new_P2_U4911 = ~new_P2_U4910 | ~new_P2_U4909 | ~new_P2_U4908;
  assign new_P2_U4912 = ~new_P2_R1054_U74 | ~new_P2_U3051;
  assign new_P2_U4913 = ~new_P2_U5764 | ~new_P2_U3403;
  assign new_P2_U4914 = ~new_P2_U3042 | ~new_P2_U4911;
  assign new_P2_U4915 = ~new_P2_R1212_U53 | ~new_P2_U3041;
  assign new_P2_U4916 = ~P2_REG3_REG_5_ | ~n2555;
  assign new_P2_U4917 = ~new_P2_R1209_U53 | ~new_P2_U3038;
  assign new_P2_U4918 = ~P2_ADDR_REG_5_ | ~new_P2_U4756;
  assign new_P2_U4919 = ~new_P2_R1212_U54 | ~new_P2_U3040;
  assign new_P2_U4920 = ~new_P2_U3039 | ~new_P2_U3400;
  assign new_P2_U4921 = ~new_P2_R1209_U54 | ~new_P2_U3037;
  assign new_P2_U4922 = ~new_P2_U4921 | ~new_P2_U4920 | ~new_P2_U4919;
  assign new_P2_U4923 = ~new_P2_R1054_U75 | ~new_P2_U3051;
  assign new_P2_U4924 = ~new_P2_U5764 | ~new_P2_U3400;
  assign new_P2_U4925 = ~new_P2_U3042 | ~new_P2_U4922;
  assign new_P2_U4926 = ~new_P2_R1212_U54 | ~new_P2_U3041;
  assign new_P2_U4927 = ~P2_REG3_REG_4_ | ~n2555;
  assign new_P2_U4928 = ~new_P2_R1209_U54 | ~new_P2_U3038;
  assign new_P2_U4929 = ~P2_ADDR_REG_4_ | ~new_P2_U4756;
  assign new_P2_U4930 = ~new_P2_R1212_U55 | ~new_P2_U3040;
  assign new_P2_U4931 = ~new_P2_U3039 | ~new_P2_U3397;
  assign new_P2_U4932 = ~new_P2_R1209_U55 | ~new_P2_U3037;
  assign new_P2_U4933 = ~new_P2_U4932 | ~new_P2_U4931 | ~new_P2_U4930;
  assign new_P2_U4934 = ~new_P2_R1054_U14 | ~new_P2_U3051;
  assign new_P2_U4935 = ~new_P2_U5764 | ~new_P2_U3397;
  assign new_P2_U4936 = ~new_P2_U3042 | ~new_P2_U4933;
  assign new_P2_U4937 = ~new_P2_R1212_U55 | ~new_P2_U3041;
  assign new_P2_U4938 = ~P2_REG3_REG_3_ | ~n2555;
  assign new_P2_U4939 = ~new_P2_R1209_U55 | ~new_P2_U3038;
  assign new_P2_U4940 = ~P2_ADDR_REG_3_ | ~new_P2_U4756;
  assign new_P2_U4941 = ~new_P2_R1212_U56 | ~new_P2_U3040;
  assign new_P2_U4942 = ~new_P2_U3039 | ~new_P2_U3394;
  assign new_P2_U4943 = ~new_P2_R1209_U56 | ~new_P2_U3037;
  assign new_P2_U4944 = ~new_P2_U4943 | ~new_P2_U4942 | ~new_P2_U4941;
  assign new_P2_U4945 = ~new_P2_R1054_U76 | ~new_P2_U3051;
  assign new_P2_U4946 = ~new_P2_U5764 | ~new_P2_U3394;
  assign new_P2_U4947 = ~new_P2_U3042 | ~new_P2_U4944;
  assign new_P2_U4948 = ~new_P2_R1212_U56 | ~new_P2_U3041;
  assign new_P2_U4949 = ~P2_REG3_REG_2_ | ~n2555;
  assign new_P2_U4950 = ~new_P2_R1209_U56 | ~new_P2_U3038;
  assign new_P2_U4951 = ~P2_ADDR_REG_2_ | ~new_P2_U4756;
  assign new_P2_U4952 = ~new_P2_R1212_U57 | ~new_P2_U3040;
  assign new_P2_U4953 = ~new_P2_U3039 | ~new_P2_U3391;
  assign new_P2_U4954 = ~new_P2_R1209_U57 | ~new_P2_U3037;
  assign new_P2_U4955 = ~new_P2_U4954 | ~new_P2_U4953 | ~new_P2_U4952;
  assign new_P2_U4956 = ~new_P2_R1054_U66 | ~new_P2_U3051;
  assign new_P2_U4957 = ~new_P2_U5764 | ~new_P2_U3391;
  assign new_P2_U4958 = ~new_P2_U3042 | ~new_P2_U4955;
  assign new_P2_U4959 = ~new_P2_R1212_U57 | ~new_P2_U3041;
  assign new_P2_U4960 = ~P2_REG3_REG_1_ | ~n2555;
  assign new_P2_U4961 = ~new_P2_R1209_U57 | ~new_P2_U3038;
  assign new_P2_U4962 = ~P2_ADDR_REG_1_ | ~new_P2_U4756;
  assign new_P2_U4963 = ~new_P2_R1212_U7 | ~new_P2_U3040;
  assign new_P2_U4964 = ~new_P2_U3039 | ~new_P2_U3386;
  assign new_P2_U4965 = ~new_P2_R1209_U7 | ~new_P2_U3037;
  assign new_P2_U4966 = ~new_P2_U4965 | ~new_P2_U4964 | ~new_P2_U4963;
  assign new_P2_U4967 = ~new_P2_R1054_U17 | ~new_P2_U3051;
  assign new_P2_U4968 = ~new_P2_U5764 | ~new_P2_U3386;
  assign new_P2_U4969 = ~new_P2_U3042 | ~new_P2_U4966;
  assign new_P2_U4970 = ~new_P2_R1212_U7 | ~new_P2_U3041;
  assign new_P2_U4971 = ~P2_REG3_REG_0_ | ~n2555;
  assign new_P2_U4972 = ~new_P2_R1209_U7 | ~new_P2_U3038;
  assign new_P2_U4973 = ~P2_ADDR_REG_0_ | ~new_P2_U4756;
  assign new_P2_U4974 = ~new_P2_U3864;
  assign new_P2_U4975 = ~new_P2_U3050 | ~new_P2_U5938 | ~new_P2_U5937;
  assign new_P2_U4976 = ~new_P2_U3863 | ~new_P2_U3023 | ~new_P2_U3905;
  assign new_P2_U4977 = ~P2_B_REG | ~new_P2_U4975;
  assign new_P2_U4978 = ~new_P2_U3036 | ~new_P2_U3078;
  assign new_P2_U4979 = ~new_P2_U3032 | ~new_P2_U3072;
  assign new_P2_U4980 = ~new_P2_SUB_605_U21 | ~new_P2_U3304;
  assign new_P2_U4981 = ~new_P2_U4980 | ~new_P2_U4979 | ~new_P2_U4978;
  assign new_P2_U4982 = ~new_P2_U3312 | ~new_P2_U5421 | ~new_P2_U3884 | ~new_P2_U3311 | ~new_P2_U3871;
  assign new_P2_U4983 = ~new_P2_U3890 | ~new_P2_U4982;
  assign new_P2_U4984 = ~new_P2_U3885 | ~new_P2_U3891;
  assign new_P2_U4985 = ~new_P2_U4984 | ~new_P2_U4983;
  assign new_P2_U4986 = ~new_P2_U3907 | ~new_P2_U3378;
  assign new_P2_U4987 = ~new_P2_U3885 | ~new_P2_U3304;
  assign new_P2_U4988 = ~new_P2_U4982 | ~new_P2_U3303;
  assign new_P2_U4989 = ~new_P2_U3370;
  assign new_P2_U4990 = ~new_P2_U3434 | ~new_P2_U5416;
  assign new_P2_U4991 = ~new_P2_SUB_605_U21 | ~new_P2_U3371;
  assign new_P2_U4992 = ~new_P2_R1158_U114 | ~new_P2_U3035;
  assign new_P2_U4993 = ~new_P2_U3031 | ~new_P2_U4981;
  assign new_P2_U4994 = ~P2_REG3_REG_15_ | ~n2555;
  assign new_P2_U4995 = ~new_P2_U3036 | ~new_P2_U3057;
  assign new_P2_U4996 = ~new_P2_U3032 | ~new_P2_U3052;
  assign new_P2_U4997 = ~new_P2_SUB_605_U27 | ~new_P2_U3304;
  assign new_P2_U4998 = ~new_P2_U4997 | ~new_P2_U4996 | ~new_P2_U4995;
  assign new_P2_U4999 = ~new_P2_U3365 | ~new_P2_U3303;
  assign new_P2_U5000 = ~new_P2_U4989 | ~new_P2_U4999;
  assign new_P2_U5001 = ~new_P2_U3890 | ~new_P2_U3365;
  assign new_P2_U5002 = ~new_P2_U3360 | ~new_P2_U5001;
  assign new_P2_U5003 = ~new_P2_U3045 | ~new_P2_U3897;
  assign new_P2_U5004 = ~new_P2_U3044 | ~new_P2_SUB_605_U27;
  assign new_P2_U5005 = ~new_P2_R1158_U17 | ~new_P2_U3035;
  assign new_P2_U5006 = ~new_P2_U3031 | ~new_P2_U4998;
  assign new_P2_U5007 = ~P2_REG3_REG_26_ | ~n2555;
  assign new_P2_U5008 = ~new_P2_U3036 | ~new_P2_U3066;
  assign new_P2_U5009 = ~new_P2_U3032 | ~new_P2_U3069;
  assign new_P2_U5010 = ~new_P2_SUB_605_U8 | ~new_P2_U3304;
  assign new_P2_U5011 = ~new_P2_U5010 | ~new_P2_U5009 | ~new_P2_U5008;
  assign new_P2_U5012 = ~new_P2_U3407 | ~new_P2_U5416;
  assign new_P2_U5013 = ~new_P2_SUB_605_U8 | ~new_P2_U3371;
  assign new_P2_U5014 = ~new_P2_R1158_U99 | ~new_P2_U3035;
  assign new_P2_U5015 = ~new_P2_U3031 | ~new_P2_U5011;
  assign new_P2_U5016 = ~P2_REG3_REG_6_ | ~n2555;
  assign new_P2_U5017 = ~new_P2_U3036 | ~new_P2_U3068;
  assign new_P2_U5018 = ~new_P2_U3032 | ~new_P2_U3080;
  assign new_P2_U5019 = ~new_P2_SUB_605_U11 | ~new_P2_U3304;
  assign new_P2_U5020 = ~new_P2_U5019 | ~new_P2_U5018 | ~new_P2_U5017;
  assign new_P2_U5021 = ~new_P2_U3443 | ~new_P2_U5416;
  assign new_P2_U5022 = ~new_P2_SUB_605_U11 | ~new_P2_U3371;
  assign new_P2_U5023 = ~new_P2_R1158_U112 | ~new_P2_U3035;
  assign new_P2_U5024 = ~new_P2_U3031 | ~new_P2_U5020;
  assign new_P2_U5025 = ~P2_REG3_REG_18_ | ~n2555;
  assign new_P2_U5026 = ~new_P2_U3036 | ~new_P2_U3077;
  assign new_P2_U5027 = ~new_P2_U3032 | ~new_P2_U3063;
  assign new_P2_U5028 = ~P2_REG3_REG_2_ | ~new_P2_U3304;
  assign new_P2_U5029 = ~new_P2_U5028 | ~new_P2_U5027 | ~new_P2_U5026;
  assign new_P2_U5030 = ~new_P2_U3395 | ~new_P2_U5416;
  assign new_P2_U5031 = ~P2_REG3_REG_2_ | ~new_P2_U3371;
  assign new_P2_U5032 = ~new_P2_R1158_U102 | ~new_P2_U3035;
  assign new_P2_U5033 = ~new_P2_U3031 | ~new_P2_U5029;
  assign new_P2_U5034 = ~P2_REG3_REG_2_ | ~n2555;
  assign new_P2_U5035 = ~new_P2_U3036 | ~new_P2_U3061;
  assign new_P2_U5036 = ~new_P2_U3032 | ~new_P2_U3071;
  assign new_P2_U5037 = ~new_P2_SUB_605_U9 | ~new_P2_U3304;
  assign new_P2_U5038 = ~new_P2_U5037 | ~new_P2_U5036 | ~new_P2_U5035;
  assign new_P2_U5039 = ~new_P2_U3422 | ~new_P2_U5416;
  assign new_P2_U5040 = ~new_P2_SUB_605_U9 | ~new_P2_U3371;
  assign new_P2_U5041 = ~new_P2_R1158_U117 | ~new_P2_U3035;
  assign new_P2_U5042 = ~new_P2_U3031 | ~new_P2_U5038;
  assign new_P2_U5043 = ~P2_REG3_REG_11_ | ~n2555;
  assign new_P2_U5044 = ~new_P2_U3036 | ~new_P2_U3074;
  assign new_P2_U5045 = ~new_P2_U3032 | ~new_P2_U3065;
  assign new_P2_U5046 = ~new_P2_SUB_605_U17 | ~new_P2_U3304;
  assign new_P2_U5047 = ~new_P2_U5046 | ~new_P2_U5045 | ~new_P2_U5044;
  assign new_P2_U5048 = ~new_P2_U3045 | ~new_P2_U3901;
  assign new_P2_U5049 = ~new_P2_U3044 | ~new_P2_SUB_605_U17;
  assign new_P2_U5050 = ~new_P2_R1158_U108 | ~new_P2_U3035;
  assign new_P2_U5051 = ~new_P2_U3031 | ~new_P2_U5047;
  assign new_P2_U5052 = ~P2_REG3_REG_22_ | ~n2555;
  assign new_P2_U5053 = ~new_P2_U3036 | ~new_P2_U3071;
  assign new_P2_U5054 = ~new_P2_U3032 | ~new_P2_U3078;
  assign new_P2_U5055 = ~new_P2_SUB_605_U25 | ~new_P2_U3304;
  assign new_P2_U5056 = ~new_P2_U5055 | ~new_P2_U5054 | ~new_P2_U5053;
  assign new_P2_U5057 = ~new_P2_U3428 | ~new_P2_U5416;
  assign new_P2_U5058 = ~new_P2_SUB_605_U25 | ~new_P2_U3371;
  assign new_P2_U5059 = ~new_P2_R1158_U14 | ~new_P2_U3035;
  assign new_P2_U5060 = ~new_P2_U3031 | ~new_P2_U5056;
  assign new_P2_U5061 = ~P2_REG3_REG_13_ | ~n2555;
  assign new_P2_U5062 = ~new_P2_U3036 | ~new_P2_U3080;
  assign new_P2_U5063 = ~new_P2_U3032 | ~new_P2_U3074;
  assign new_P2_U5064 = ~new_P2_SUB_605_U20 | ~new_P2_U3304;
  assign new_P2_U5065 = ~new_P2_U5064 | ~new_P2_U5063 | ~new_P2_U5062;
  assign new_P2_U5066 = ~new_P2_U3045 | ~new_P2_U3903;
  assign new_P2_U5067 = ~new_P2_U3044 | ~new_P2_SUB_605_U20;
  assign new_P2_U5068 = ~new_P2_R1158_U109 | ~new_P2_U3035;
  assign new_P2_U5069 = ~new_P2_U3031 | ~new_P2_U5065;
  assign new_P2_U5070 = ~P2_REG3_REG_20_ | ~n2555;
  assign new_P2_U5071 = ~new_P2_U3031 | ~new_P2_U3304;
  assign new_P2_U5072 = ~new_P2_U5415 | ~new_P2_U5071;
  assign new_P2_U5073 = ~new_P2_U3792 | ~new_P2_U3032;
  assign new_P2_U5074 = ~new_P2_U3387 | ~new_P2_U5416;
  assign new_P2_U5075 = ~P2_REG3_REG_0_ | ~new_P2_U5072;
  assign new_P2_U5076 = ~new_P2_R1158_U96 | ~new_P2_U3035;
  assign new_P2_U5077 = ~P2_REG3_REG_0_ | ~n2555;
  assign new_P2_U5078 = ~new_P2_U3036 | ~new_P2_U3083;
  assign new_P2_U5079 = ~new_P2_U3032 | ~new_P2_U3061;
  assign new_P2_U5080 = ~new_P2_SUB_605_U14 | ~new_P2_U3304;
  assign new_P2_U5081 = ~new_P2_U5080 | ~new_P2_U5079 | ~new_P2_U5078;
  assign new_P2_U5082 = ~new_P2_U3416 | ~new_P2_U5416;
  assign new_P2_U5083 = ~new_P2_SUB_605_U14 | ~new_P2_U3371;
  assign new_P2_U5084 = ~new_P2_R1158_U97 | ~new_P2_U3035;
  assign new_P2_U5085 = ~new_P2_U3031 | ~new_P2_U5081;
  assign new_P2_U5086 = ~P2_REG3_REG_9_ | ~n2555;
  assign new_P2_U5087 = ~new_P2_U3036 | ~new_P2_U3063;
  assign new_P2_U5088 = ~new_P2_U3032 | ~new_P2_U3066;
  assign new_P2_U5089 = ~new_P2_SUB_605_U30 | ~new_P2_U3304;
  assign new_P2_U5090 = ~new_P2_U5089 | ~new_P2_U5088 | ~new_P2_U5087;
  assign new_P2_U5091 = ~new_P2_U3401 | ~new_P2_U5416;
  assign new_P2_U5092 = ~new_P2_SUB_605_U30 | ~new_P2_U3371;
  assign new_P2_U5093 = ~new_P2_R1158_U101 | ~new_P2_U3035;
  assign new_P2_U5094 = ~new_P2_U3031 | ~new_P2_U5090;
  assign new_P2_U5095 = ~P2_REG3_REG_4_ | ~n2555;
  assign new_P2_U5096 = ~new_P2_U3036 | ~new_P2_U3065;
  assign new_P2_U5097 = ~new_P2_U3032 | ~new_P2_U3057;
  assign new_P2_U5098 = ~new_P2_SUB_605_U10 | ~new_P2_U3304;
  assign new_P2_U5099 = ~new_P2_U5098 | ~new_P2_U5097 | ~new_P2_U5096;
  assign new_P2_U5100 = ~new_P2_U3045 | ~new_P2_U3899;
  assign new_P2_U5101 = ~new_P2_U3044 | ~new_P2_SUB_605_U10;
  assign new_P2_U5102 = ~new_P2_R1158_U106 | ~new_P2_U3035;
  assign new_P2_U5103 = ~new_P2_U3031 | ~new_P2_U5099;
  assign new_P2_U5104 = ~P2_REG3_REG_24_ | ~n2555;
  assign new_P2_U5105 = ~new_P2_U3036 | ~new_P2_U3072;
  assign new_P2_U5106 = ~new_P2_U3032 | ~new_P2_U3081;
  assign new_P2_U5107 = ~new_P2_SUB_605_U19 | ~new_P2_U3304;
  assign new_P2_U5108 = ~new_P2_U5107 | ~new_P2_U5106 | ~new_P2_U5105;
  assign new_P2_U5109 = ~new_P2_U3440 | ~new_P2_U5416;
  assign new_P2_U5110 = ~new_P2_SUB_605_U19 | ~new_P2_U3371;
  assign new_P2_U5111 = ~new_P2_R1158_U15 | ~new_P2_U3035;
  assign new_P2_U5112 = ~new_P2_U3031 | ~new_P2_U5108;
  assign new_P2_U5113 = ~P2_REG3_REG_17_ | ~n2555;
  assign new_P2_U5114 = ~new_P2_U3036 | ~new_P2_U3059;
  assign new_P2_U5115 = ~new_P2_U3032 | ~new_P2_U3070;
  assign new_P2_U5116 = ~new_P2_SUB_605_U22 | ~new_P2_U3304;
  assign new_P2_U5117 = ~new_P2_U5116 | ~new_P2_U5115 | ~new_P2_U5114;
  assign new_P2_U5118 = ~new_P2_U3404 | ~new_P2_U5416;
  assign new_P2_U5119 = ~new_P2_SUB_605_U22 | ~new_P2_U3371;
  assign new_P2_U5120 = ~new_P2_R1158_U100 | ~new_P2_U3035;
  assign new_P2_U5121 = ~new_P2_U3031 | ~new_P2_U5117;
  assign new_P2_U5122 = ~P2_REG3_REG_5_ | ~n2555;
  assign new_P2_U5123 = ~new_P2_U3036 | ~new_P2_U3073;
  assign new_P2_U5124 = ~new_P2_U3032 | ~new_P2_U3068;
  assign new_P2_U5125 = ~new_P2_SUB_605_U7 | ~new_P2_U3304;
  assign new_P2_U5126 = ~new_P2_U5125 | ~new_P2_U5124 | ~new_P2_U5123;
  assign new_P2_U5127 = ~new_P2_U3437 | ~new_P2_U5416;
  assign new_P2_U5128 = ~new_P2_SUB_605_U7 | ~new_P2_U3371;
  assign new_P2_U5129 = ~new_P2_R1158_U113 | ~new_P2_U3035;
  assign new_P2_U5130 = ~new_P2_U3031 | ~new_P2_U5126;
  assign new_P2_U5131 = ~P2_REG3_REG_16_ | ~n2555;
  assign new_P2_U5132 = ~new_P2_U3036 | ~new_P2_U3064;
  assign new_P2_U5133 = ~new_P2_U3032 | ~new_P2_U3056;
  assign new_P2_U5134 = ~new_P2_SUB_605_U16 | ~new_P2_U3304;
  assign new_P2_U5135 = ~new_P2_U5134 | ~new_P2_U5133 | ~new_P2_U5132;
  assign new_P2_U5136 = ~new_P2_U3045 | ~new_P2_U3898;
  assign new_P2_U5137 = ~new_P2_U3044 | ~new_P2_SUB_605_U16;
  assign new_P2_U5138 = ~new_P2_R1158_U105 | ~new_P2_U3035;
  assign new_P2_U5139 = ~new_P2_U3031 | ~new_P2_U5135;
  assign new_P2_U5140 = ~P2_REG3_REG_25_ | ~n2555;
  assign new_P2_U5141 = ~new_P2_U3036 | ~new_P2_U3062;
  assign new_P2_U5142 = ~new_P2_U3032 | ~new_P2_U3079;
  assign new_P2_U5143 = ~new_P2_SUB_605_U24 | ~new_P2_U3304;
  assign new_P2_U5144 = ~new_P2_U5143 | ~new_P2_U5142 | ~new_P2_U5141;
  assign new_P2_U5145 = ~new_P2_U3425 | ~new_P2_U5416;
  assign new_P2_U5146 = ~new_P2_SUB_605_U24 | ~new_P2_U3371;
  assign new_P2_U5147 = ~new_P2_R1158_U116 | ~new_P2_U3035;
  assign new_P2_U5148 = ~new_P2_U3031 | ~new_P2_U5144;
  assign new_P2_U5149 = ~P2_REG3_REG_12_ | ~n2555;
  assign new_P2_U5150 = ~new_P2_U3036 | ~new_P2_U3075;
  assign new_P2_U5151 = ~new_P2_U3032 | ~new_P2_U3060;
  assign new_P2_U5152 = ~new_P2_SUB_605_U28 | ~new_P2_U3304;
  assign new_P2_U5153 = ~new_P2_U5152 | ~new_P2_U5151 | ~new_P2_U5150;
  assign new_P2_U5154 = ~new_P2_U3045 | ~new_P2_U3902;
  assign new_P2_U5155 = ~new_P2_U3044 | ~new_P2_SUB_605_U28;
  assign new_P2_U5156 = ~new_P2_R1158_U16 | ~new_P2_U3035;
  assign new_P2_U5157 = ~new_P2_U3031 | ~new_P2_U5153;
  assign new_P2_U5158 = ~P2_REG3_REG_21_ | ~n2555;
  assign new_P2_U5159 = ~new_P2_U3036 | ~new_P2_U3076;
  assign new_P2_U5160 = ~new_P2_U3032 | ~new_P2_U3067;
  assign new_P2_U5161 = ~P2_REG3_REG_1_ | ~new_P2_U3304;
  assign new_P2_U5162 = ~new_P2_U5161 | ~new_P2_U5160 | ~new_P2_U5159;
  assign new_P2_U5163 = ~new_P2_U3392 | ~new_P2_U5416;
  assign new_P2_U5164 = ~P2_REG3_REG_1_ | ~new_P2_U3371;
  assign new_P2_U5165 = ~new_P2_R1158_U110 | ~new_P2_U3035;
  assign new_P2_U5166 = ~new_P2_U3031 | ~new_P2_U5162;
  assign new_P2_U5167 = ~P2_REG3_REG_1_ | ~n2555;
  assign new_P2_U5168 = ~new_P2_U3036 | ~new_P2_U3069;
  assign new_P2_U5169 = ~new_P2_U3032 | ~new_P2_U3082;
  assign new_P2_U5170 = ~new_P2_SUB_605_U12 | ~new_P2_U3304;
  assign new_P2_U5171 = ~new_P2_U5170 | ~new_P2_U5169 | ~new_P2_U5168;
  assign new_P2_U5172 = ~new_P2_U3413 | ~new_P2_U5416;
  assign new_P2_U5173 = ~new_P2_SUB_605_U12 | ~new_P2_U3371;
  assign new_P2_U5174 = ~new_P2_R1158_U98 | ~new_P2_U3035;
  assign new_P2_U5175 = ~new_P2_U3031 | ~new_P2_U5171;
  assign new_P2_U5176 = ~P2_REG3_REG_8_ | ~n2555;
  assign new_P2_U5177 = ~new_P2_U3036 | ~new_P2_U3052;
  assign new_P2_U5178 = ~new_P2_U3032 | ~new_P2_U3054;
  assign new_P2_U5179 = ~new_P2_SUB_605_U29 | ~new_P2_U3304;
  assign new_P2_U5180 = ~new_P2_U5179 | ~new_P2_U5178 | ~new_P2_U5177;
  assign new_P2_U5181 = ~new_P2_U3045 | ~new_P2_U3895;
  assign new_P2_U5182 = ~new_P2_U3044 | ~new_P2_SUB_605_U29;
  assign new_P2_U5183 = ~new_P2_R1158_U103 | ~new_P2_U3035;
  assign new_P2_U5184 = ~new_P2_U3031 | ~new_P2_U5180;
  assign new_P2_U5185 = ~P2_REG3_REG_28_ | ~n2555;
  assign new_P2_U5186 = ~new_P2_U3036 | ~new_P2_U3081;
  assign new_P2_U5187 = ~new_P2_U3032 | ~new_P2_U3075;
  assign new_P2_U5188 = ~new_P2_SUB_605_U15 | ~new_P2_U3304;
  assign new_P2_U5189 = ~new_P2_U5188 | ~new_P2_U5187 | ~new_P2_U5186;
  assign new_P2_U5190 = ~new_P2_U3445 | ~new_P2_U5416;
  assign new_P2_U5191 = ~new_P2_SUB_605_U15 | ~new_P2_U3371;
  assign new_P2_U5192 = ~new_P2_R1158_U111 | ~new_P2_U3035;
  assign new_P2_U5193 = ~new_P2_U3031 | ~new_P2_U5189;
  assign new_P2_U5194 = ~P2_REG3_REG_19_ | ~n2555;
  assign new_P2_U5195 = ~new_P2_U3036 | ~new_P2_U3067;
  assign new_P2_U5196 = ~new_P2_U3032 | ~new_P2_U3059;
  assign new_P2_U5197 = ~new_P2_SUB_605_U26 | ~new_P2_U3304;
  assign new_P2_U5198 = ~new_P2_U5197 | ~new_P2_U5196 | ~new_P2_U5195;
  assign new_P2_U5199 = ~new_P2_U3398 | ~new_P2_U5416;
  assign new_P2_U5200 = ~new_P2_SUB_605_U26 | ~new_P2_U3371;
  assign new_P2_U5201 = ~new_P2_R1158_U18 | ~new_P2_U3035;
  assign new_P2_U5202 = ~new_P2_U3031 | ~new_P2_U5198;
  assign new_P2_U5203 = ~P2_REG3_REG_3_ | ~n2555;
  assign new_P2_U5204 = ~new_P2_U3036 | ~new_P2_U3082;
  assign new_P2_U5205 = ~new_P2_U3032 | ~new_P2_U3062;
  assign new_P2_U5206 = ~new_P2_SUB_605_U13 | ~new_P2_U3304;
  assign new_P2_U5207 = ~new_P2_U5206 | ~new_P2_U5205 | ~new_P2_U5204;
  assign new_P2_U5208 = ~new_P2_U3419 | ~new_P2_U5416;
  assign new_P2_U5209 = ~new_P2_SUB_605_U13 | ~new_P2_U3371;
  assign new_P2_U5210 = ~new_P2_R1158_U118 | ~new_P2_U3035;
  assign new_P2_U5211 = ~new_P2_U3031 | ~new_P2_U5207;
  assign new_P2_U5212 = ~P2_REG3_REG_10_ | ~n2555;
  assign new_P2_U5213 = ~new_P2_U3036 | ~new_P2_U3060;
  assign new_P2_U5214 = ~new_P2_U3032 | ~new_P2_U3064;
  assign new_P2_U5215 = ~new_P2_SUB_605_U6 | ~new_P2_U3304;
  assign new_P2_U5216 = ~new_P2_U5215 | ~new_P2_U5214 | ~new_P2_U5213;
  assign new_P2_U5217 = ~new_P2_U3045 | ~new_P2_U3900;
  assign new_P2_U5218 = ~new_P2_U3044 | ~new_P2_SUB_605_U6;
  assign new_P2_U5219 = ~new_P2_R1158_U107 | ~new_P2_U3035;
  assign new_P2_U5220 = ~new_P2_U3031 | ~new_P2_U5216;
  assign new_P2_U5221 = ~P2_REG3_REG_23_ | ~n2555;
  assign new_P2_U5222 = ~new_P2_U3036 | ~new_P2_U3079;
  assign new_P2_U5223 = ~new_P2_U3032 | ~new_P2_U3073;
  assign new_P2_U5224 = ~new_P2_SUB_605_U31 | ~new_P2_U3304;
  assign new_P2_U5225 = ~new_P2_U5224 | ~new_P2_U5223 | ~new_P2_U5222;
  assign new_P2_U5226 = ~new_P2_U3431 | ~new_P2_U5416;
  assign new_P2_U5227 = ~new_P2_SUB_605_U31 | ~new_P2_U3371;
  assign new_P2_U5228 = ~new_P2_R1158_U115 | ~new_P2_U3035;
  assign new_P2_U5229 = ~new_P2_U3031 | ~new_P2_U5225;
  assign new_P2_U5230 = ~P2_REG3_REG_14_ | ~n2555;
  assign new_P2_U5231 = ~new_P2_U3036 | ~new_P2_U3056;
  assign new_P2_U5232 = ~new_P2_U3032 | ~new_P2_U3053;
  assign new_P2_U5233 = ~new_P2_SUB_605_U23 | ~new_P2_U3304;
  assign new_P2_U5234 = ~new_P2_U5233 | ~new_P2_U5232 | ~new_P2_U5231;
  assign new_P2_U5235 = ~new_P2_U3045 | ~new_P2_U3896;
  assign new_P2_U5236 = ~new_P2_U3044 | ~new_P2_SUB_605_U23;
  assign new_P2_U5237 = ~new_P2_R1158_U104 | ~new_P2_U3035;
  assign new_P2_U5238 = ~new_P2_U3031 | ~new_P2_U5234;
  assign new_P2_U5239 = ~P2_REG3_REG_27_ | ~n2555;
  assign new_P2_U5240 = ~new_P2_U3036 | ~new_P2_U3070;
  assign new_P2_U5241 = ~new_P2_U3032 | ~new_P2_U3083;
  assign new_P2_U5242 = ~new_P2_SUB_605_U18 | ~new_P2_U3304;
  assign new_P2_U5243 = ~new_P2_U5242 | ~new_P2_U5241 | ~new_P2_U5240;
  assign new_P2_U5244 = ~new_P2_U3410 | ~new_P2_U5416;
  assign new_P2_U5245 = ~new_P2_SUB_605_U18 | ~new_P2_U3371;
  assign new_P2_U5246 = ~new_P2_R1158_U19 | ~new_P2_U3035;
  assign new_P2_U5247 = ~new_P2_U3031 | ~new_P2_U5243;
  assign new_P2_U5248 = ~P2_REG3_REG_7_ | ~n2555;
  assign new_P2_U5249 = ~new_P2_U3894 | ~new_P2_U3046;
  assign new_P2_U5250 = ~new_P2_U3375 | ~new_P2_U3829;
  assign new_P2_U5251 = ~new_P2_U3821 | ~new_P2_U3820;
  assign new_P2_U5252 = ~new_P2_U3819 | ~new_P2_U3013;
  assign new_P2_U5253 = ~new_P2_U3876 | ~new_P2_U5252;
  assign new_P2_U5254 = ~new_P2_U3416 | ~new_P2_U5253;
  assign new_P2_U5255 = ~new_P2_U5251 | ~new_P2_U3082;
  assign new_P2_U5256 = ~new_P2_U3413 | ~new_P2_U5253;
  assign new_P2_U5257 = ~new_P2_U5251 | ~new_P2_U3083;
  assign new_P2_U5258 = ~new_P2_U3410 | ~new_P2_U5253;
  assign new_P2_U5259 = ~new_P2_U5251 | ~new_P2_U3069;
  assign new_P2_U5260 = ~new_P2_U3407 | ~new_P2_U5253;
  assign new_P2_U5261 = ~new_P2_U5251 | ~new_P2_U3070;
  assign new_P2_U5262 = ~new_P2_U3404 | ~new_P2_U5253;
  assign new_P2_U5263 = ~new_P2_U5251 | ~new_P2_U3066;
  assign new_P2_U5264 = ~new_P2_U3401 | ~new_P2_U5253;
  assign new_P2_U5265 = ~new_P2_U5251 | ~new_P2_U3059;
  assign new_P2_U5266 = ~new_P2_U3868 | ~new_P2_U5253;
  assign new_P2_U5267 = ~new_P2_U5251 | ~new_P2_U3055;
  assign new_P2_U5268 = ~new_P2_U3869 | ~new_P2_U5253;
  assign new_P2_U5269 = ~new_P2_U5251 | ~new_P2_U3058;
  assign new_P2_U5270 = ~new_P2_U3398 | ~new_P2_U5253;
  assign new_P2_U5271 = ~new_P2_U5251 | ~new_P2_U3063;
  assign new_P2_U5272 = ~new_P2_U3904 | ~new_P2_U5253;
  assign new_P2_U5273 = ~new_P2_U5251 | ~new_P2_U3054;
  assign new_P2_U5274 = ~new_P2_U3895 | ~new_P2_U5253;
  assign new_P2_U5275 = ~new_P2_U5251 | ~new_P2_U3053;
  assign new_P2_U5276 = ~new_P2_U3896 | ~new_P2_U5253;
  assign new_P2_U5277 = ~new_P2_U5251 | ~new_P2_U3052;
  assign new_P2_U5278 = ~new_P2_U3897 | ~new_P2_U5253;
  assign new_P2_U5279 = ~new_P2_U5251 | ~new_P2_U3056;
  assign new_P2_U5280 = ~new_P2_U3898 | ~new_P2_U5253;
  assign new_P2_U5281 = ~new_P2_U5251 | ~new_P2_U3057;
  assign new_P2_U5282 = ~new_P2_U3899 | ~new_P2_U5253;
  assign new_P2_U5283 = ~new_P2_U5251 | ~new_P2_U3064;
  assign new_P2_U5284 = ~new_P2_U3900 | ~new_P2_U5253;
  assign new_P2_U5285 = ~new_P2_U5251 | ~new_P2_U3065;
  assign new_P2_U5286 = ~new_P2_U3901 | ~new_P2_U5253;
  assign new_P2_U5287 = ~new_P2_U5251 | ~new_P2_U3060;
  assign new_P2_U5288 = ~new_P2_U3902 | ~new_P2_U5253;
  assign new_P2_U5289 = ~new_P2_U5251 | ~new_P2_U3074;
  assign new_P2_U5290 = ~new_P2_U3903 | ~new_P2_U5253;
  assign new_P2_U5291 = ~new_P2_U5251 | ~new_P2_U3075;
  assign new_P2_U5292 = ~new_P2_U3395 | ~new_P2_U5253;
  assign new_P2_U5293 = ~new_P2_U5251 | ~new_P2_U3067;
  assign new_P2_U5294 = ~new_P2_U3445 | ~new_P2_U5253;
  assign new_P2_U5295 = ~new_P2_U5251 | ~new_P2_U3080;
  assign new_P2_U5296 = ~new_P2_U3443 | ~new_P2_U5253;
  assign new_P2_U5297 = ~new_P2_U5251 | ~new_P2_U3081;
  assign new_P2_U5298 = ~new_P2_U3440 | ~new_P2_U5253;
  assign new_P2_U5299 = ~new_P2_U5251 | ~new_P2_U3068;
  assign new_P2_U5300 = ~new_P2_U3437 | ~new_P2_U5253;
  assign new_P2_U5301 = ~new_P2_U5251 | ~new_P2_U3072;
  assign new_P2_U5302 = ~new_P2_U3434 | ~new_P2_U5253;
  assign new_P2_U5303 = ~new_P2_U5251 | ~new_P2_U3073;
  assign new_P2_U5304 = ~new_P2_U3431 | ~new_P2_U5253;
  assign new_P2_U5305 = ~new_P2_U5251 | ~new_P2_U3078;
  assign new_P2_U5306 = ~new_P2_U3428 | ~new_P2_U5253;
  assign new_P2_U5307 = ~new_P2_U5251 | ~new_P2_U3079;
  assign new_P2_U5308 = ~new_P2_U3425 | ~new_P2_U5253;
  assign new_P2_U5309 = ~new_P2_U5251 | ~new_P2_U3071;
  assign new_P2_U5310 = ~new_P2_U3422 | ~new_P2_U5253;
  assign new_P2_U5311 = ~new_P2_U5251 | ~new_P2_U3062;
  assign new_P2_U5312 = ~new_P2_U3419 | ~new_P2_U5253;
  assign new_P2_U5313 = ~new_P2_U5251 | ~new_P2_U3061;
  assign new_P2_U5314 = ~new_P2_U3392 | ~new_P2_U5253;
  assign new_P2_U5315 = ~new_P2_U5251 | ~new_P2_U3077;
  assign new_P2_U5316 = ~new_P2_U3387 | ~new_P2_U5253;
  assign new_P2_U5317 = ~new_P2_U5251 | ~new_P2_U3076;
  assign new_P2_U5318 = ~new_P2_U3416 | ~new_P2_U5251;
  assign new_P2_U5319 = ~new_P2_U5253 | ~new_P2_U3082;
  assign new_P2_U5320 = ~new_P2_U5436 | ~new_P2_U3083;
  assign new_P2_U5321 = ~new_P2_U3413 | ~new_P2_U5251;
  assign new_P2_U5322 = ~new_P2_U5253 | ~new_P2_U3083;
  assign new_P2_U5323 = ~new_P2_U5436 | ~new_P2_U3069;
  assign new_P2_U5324 = ~new_P2_U3410 | ~new_P2_U5251;
  assign new_P2_U5325 = ~new_P2_U5253 | ~new_P2_U3069;
  assign new_P2_U5326 = ~new_P2_U5436 | ~new_P2_U3070;
  assign new_P2_U5327 = ~new_P2_U3407 | ~new_P2_U5251;
  assign new_P2_U5328 = ~new_P2_U5253 | ~new_P2_U3070;
  assign new_P2_U5329 = ~new_P2_U5436 | ~new_P2_U3066;
  assign new_P2_U5330 = ~new_P2_U3404 | ~new_P2_U5251;
  assign new_P2_U5331 = ~new_P2_U5253 | ~new_P2_U3066;
  assign new_P2_U5332 = ~new_P2_U5436 | ~new_P2_U3059;
  assign new_P2_U5333 = ~new_P2_U3401 | ~new_P2_U5251;
  assign new_P2_U5334 = ~new_P2_U5253 | ~new_P2_U3059;
  assign new_P2_U5335 = ~new_P2_U5436 | ~new_P2_U3063;
  assign new_P2_U5336 = ~new_P2_U5253 | ~new_P2_U3055;
  assign new_P2_U5337 = ~new_P2_U3868 | ~new_P2_U5251;
  assign new_P2_U5338 = ~new_P2_U5253 | ~new_P2_U3058;
  assign new_P2_U5339 = ~new_P2_U3869 | ~new_P2_U5251;
  assign new_P2_U5340 = ~new_P2_U3398 | ~new_P2_U5251;
  assign new_P2_U5341 = ~new_P2_U5253 | ~new_P2_U3063;
  assign new_P2_U5342 = ~new_P2_U5436 | ~new_P2_U3067;
  assign new_P2_U5343 = ~new_P2_U5253 | ~new_P2_U3054;
  assign new_P2_U5344 = ~new_P2_U3904 | ~new_P2_U5251;
  assign new_P2_U5345 = ~new_P2_U5436 | ~new_P2_U3053;
  assign new_P2_U5346 = ~new_P2_U5253 | ~new_P2_U3053;
  assign new_P2_U5347 = ~new_P2_U3895 | ~new_P2_U5251;
  assign new_P2_U5348 = ~new_P2_U5436 | ~new_P2_U3052;
  assign new_P2_U5349 = ~new_P2_U5253 | ~new_P2_U3052;
  assign new_P2_U5350 = ~new_P2_U3896 | ~new_P2_U5251;
  assign new_P2_U5351 = ~new_P2_U5436 | ~new_P2_U3056;
  assign new_P2_U5352 = ~new_P2_U5253 | ~new_P2_U3056;
  assign new_P2_U5353 = ~new_P2_U3897 | ~new_P2_U5251;
  assign new_P2_U5354 = ~new_P2_U5436 | ~new_P2_U3057;
  assign new_P2_U5355 = ~new_P2_U5253 | ~new_P2_U3057;
  assign new_P2_U5356 = ~new_P2_U3898 | ~new_P2_U5251;
  assign new_P2_U5357 = ~new_P2_U5436 | ~new_P2_U3064;
  assign new_P2_U5358 = ~new_P2_U5253 | ~new_P2_U3064;
  assign new_P2_U5359 = ~new_P2_U3899 | ~new_P2_U5251;
  assign new_P2_U5360 = ~new_P2_U5436 | ~new_P2_U3065;
  assign new_P2_U5361 = ~new_P2_U5253 | ~new_P2_U3065;
  assign new_P2_U5362 = ~new_P2_U3900 | ~new_P2_U5251;
  assign new_P2_U5363 = ~new_P2_U5436 | ~new_P2_U3060;
  assign new_P2_U5364 = ~new_P2_U5253 | ~new_P2_U3060;
  assign new_P2_U5365 = ~new_P2_U3901 | ~new_P2_U5251;
  assign new_P2_U5366 = ~new_P2_U5436 | ~new_P2_U3074;
  assign new_P2_U5367 = ~new_P2_U5253 | ~new_P2_U3074;
  assign new_P2_U5368 = ~new_P2_U3902 | ~new_P2_U5251;
  assign new_P2_U5369 = ~new_P2_U5436 | ~new_P2_U3075;
  assign new_P2_U5370 = ~new_P2_U5253 | ~new_P2_U3075;
  assign new_P2_U5371 = ~new_P2_U3903 | ~new_P2_U5251;
  assign new_P2_U5372 = ~new_P2_U5436 | ~new_P2_U3080;
  assign new_P2_U5373 = ~new_P2_U3395 | ~new_P2_U5251;
  assign new_P2_U5374 = ~new_P2_U5253 | ~new_P2_U3067;
  assign new_P2_U5375 = ~new_P2_U5436 | ~new_P2_U3077;
  assign new_P2_U5376 = ~new_P2_U3445 | ~new_P2_U5251;
  assign new_P2_U5377 = ~new_P2_U5253 | ~new_P2_U3080;
  assign new_P2_U5378 = ~new_P2_U5436 | ~new_P2_U3081;
  assign new_P2_U5379 = ~new_P2_U3443 | ~new_P2_U5251;
  assign new_P2_U5380 = ~new_P2_U5253 | ~new_P2_U3081;
  assign new_P2_U5381 = ~new_P2_U5436 | ~new_P2_U3068;
  assign new_P2_U5382 = ~new_P2_U3440 | ~new_P2_U5251;
  assign new_P2_U5383 = ~new_P2_U5253 | ~new_P2_U3068;
  assign new_P2_U5384 = ~new_P2_U5436 | ~new_P2_U3072;
  assign new_P2_U5385 = ~new_P2_U3437 | ~new_P2_U5251;
  assign new_P2_U5386 = ~new_P2_U5253 | ~new_P2_U3072;
  assign new_P2_U5387 = ~new_P2_U5436 | ~new_P2_U3073;
  assign new_P2_U5388 = ~new_P2_U3434 | ~new_P2_U5251;
  assign new_P2_U5389 = ~new_P2_U5253 | ~new_P2_U3073;
  assign new_P2_U5390 = ~new_P2_U5436 | ~new_P2_U3078;
  assign new_P2_U5391 = ~new_P2_U3431 | ~new_P2_U5251;
  assign new_P2_U5392 = ~new_P2_U5253 | ~new_P2_U3078;
  assign new_P2_U5393 = ~new_P2_U5436 | ~new_P2_U3079;
  assign new_P2_U5394 = ~new_P2_U3428 | ~new_P2_U5251;
  assign new_P2_U5395 = ~new_P2_U5253 | ~new_P2_U3079;
  assign new_P2_U5396 = ~new_P2_U5436 | ~new_P2_U3071;
  assign new_P2_U5397 = ~new_P2_U3425 | ~new_P2_U5251;
  assign new_P2_U5398 = ~new_P2_U5253 | ~new_P2_U3071;
  assign new_P2_U5399 = ~new_P2_U5436 | ~new_P2_U3062;
  assign new_P2_U5400 = ~new_P2_U3422 | ~new_P2_U5251;
  assign new_P2_U5401 = ~new_P2_U5253 | ~new_P2_U3062;
  assign new_P2_U5402 = ~new_P2_U5436 | ~new_P2_U3061;
  assign new_P2_U5403 = ~new_P2_U3419 | ~new_P2_U5251;
  assign new_P2_U5404 = ~new_P2_U5253 | ~new_P2_U3061;
  assign new_P2_U5405 = ~new_P2_U5436 | ~new_P2_U3082;
  assign new_P2_U5406 = ~new_P2_U3392 | ~new_P2_U5251;
  assign new_P2_U5407 = ~new_P2_U5253 | ~new_P2_U3077;
  assign new_P2_U5408 = ~new_P2_U5436 | ~new_P2_U3076;
  assign new_P2_U5409 = ~new_P2_U3387 | ~new_P2_U5251;
  assign new_P2_U5410 = ~new_P2_U5253 | ~new_P2_U3076;
  assign new_P2_U5411 = ~new_P2_U4977 | ~n2555;
  assign new_P2_U5412 = ~new_P2_U4976 | ~new_P2_U4977 | ~new_P2_U5436;
  assign new_P2_U5413 = ~new_P2_U3043 | ~new_P2_U3303;
  assign new_P2_U5414 = ~new_P2_U3043 | ~new_P2_U3890;
  assign new_P2_U5415 = ~new_P2_U3371;
  assign new_P2_U5416 = ~new_P2_U5414 | ~new_P2_U3914;
  assign new_P2_U5417 = ~new_P2_U3779 | ~new_P2_U5934 | ~new_P2_U5933;
  assign new_P2_U5418 = ~new_P2_U5430 | ~new_P2_U5424;
  assign new_P2_U5419 = ~new_P2_U3875 | ~new_P2_U3378;
  assign new_P2_U5420 = ~new_P2_U3375 | ~new_P2_U3829;
  assign new_P2_U5421 = ~new_P2_U3872 | ~new_P2_U5443;
  assign new_P2_U5422 = ~P2_IR_REG_24_ | ~new_P2_U3827;
  assign new_P2_U5423 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U19;
  assign new_P2_U5424 = ~new_P2_U3372;
  assign new_P2_U5425 = ~P2_IR_REG_25_ | ~new_P2_U3827;
  assign new_P2_U5426 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U79;
  assign new_P2_U5427 = ~new_P2_U3373;
  assign new_P2_U5428 = ~P2_IR_REG_26_ | ~new_P2_U3827;
  assign new_P2_U5429 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U20;
  assign new_P2_U5430 = ~new_P2_U3374;
  assign new_P2_U5431 = ~new_P2_U5424 | ~P2_B_REG;
  assign new_P2_U5432 = ~new_P2_U3372 | ~new_P2_U3298;
  assign new_P2_U5433 = ~new_P2_U5432 | ~new_P2_U5431;
  assign new_P2_U5434 = ~P2_IR_REG_23_ | ~new_P2_U3827;
  assign new_P2_U5435 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U18;
  assign new_P2_U5436 = ~new_P2_U3375;
  assign new_P2_U5437 = ~P2_D_REG_0_ | ~new_P2_U3828;
  assign new_P2_U5438 = ~new_P2_U3911 | ~new_P2_U4016;
  assign new_P2_U5439 = ~P2_D_REG_1_ | ~new_P2_U3828;
  assign new_P2_U5440 = ~new_P2_U3911 | ~new_P2_U4017;
  assign new_P2_U5441 = ~P2_IR_REG_20_ | ~new_P2_U3827;
  assign new_P2_U5442 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U16;
  assign new_P2_U5443 = ~new_P2_U3378;
  assign new_P2_U5444 = ~P2_IR_REG_19_ | ~new_P2_U3827;
  assign new_P2_U5445 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U15;
  assign new_P2_U5446 = ~new_P2_U3379;
  assign new_P2_U5447 = ~P2_IR_REG_22_ | ~new_P2_U3827;
  assign new_P2_U5448 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U17;
  assign new_P2_U5449 = ~new_P2_U3380;
  assign new_P2_U5450 = ~P2_IR_REG_21_ | ~new_P2_U3827;
  assign new_P2_U5451 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U81;
  assign new_P2_U5452 = ~new_P2_U3385;
  assign new_P2_U5453 = ~P2_IR_REG_30_ | ~new_P2_U3827;
  assign new_P2_U5454 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U75;
  assign new_P2_U5455 = ~new_P2_U3381;
  assign new_P2_U5456 = ~P2_IR_REG_29_ | ~new_P2_U3827;
  assign new_P2_U5457 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U22;
  assign new_P2_U5458 = ~new_P2_U3382;
  assign new_P2_U5459 = ~P2_IR_REG_28_ | ~new_P2_U3827;
  assign new_P2_U5460 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U21;
  assign new_P2_U5461 = ~new_P2_U3383;
  assign new_P2_U5462 = ~P2_IR_REG_27_ | ~new_P2_U3827;
  assign new_P2_U5463 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U77;
  assign new_P2_U5464 = ~new_P2_U3384;
  assign new_P2_U5465 = ~P2_IR_REG_0_ | ~new_P2_U3827;
  assign new_P2_U5466 = ~P2_IR_REG_31_ | ~P2_IR_REG_0_;
  assign new_P2_U5467 = ~new_U56 | ~new_P2_U3829;
  assign new_P2_U5468 = ~new_P2_U3889 | ~new_P2_U3386;
  assign new_P2_U5469 = ~new_P2_U3387;
  assign new_P2_U5470 = ~new_P2_U5418 | ~new_P2_U3300;
  assign new_P2_U5471 = ~P2_D_REG_0_ | ~new_P2_U4015;
  assign new_P2_U5472 = ~new_P2_U3388;
  assign new_P2_U5473 = ~P2_D_REG_1_ | ~new_P2_U4015;
  assign new_P2_U5474 = ~new_P2_U4017 | ~new_P2_U3300;
  assign new_P2_U5475 = ~new_P2_U3389;
  assign new_P2_U5476 = ~new_P2_U4048 | ~new_P2_U5449;
  assign new_P2_U5477 = ~new_P2_U3380 | ~new_P2_U3830;
  assign new_P2_U5478 = ~new_P2_U5477 | ~new_P2_U5476;
  assign new_P2_U5479 = ~P2_REG0_REG_0_ | ~new_P2_U3831;
  assign new_P2_U5480 = ~new_P2_U3910 | ~new_P2_U4073;
  assign new_P2_U5481 = ~P2_IR_REG_1_ | ~new_P2_U3827;
  assign new_P2_U5482 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U53;
  assign new_P2_U5483 = ~new_U45 | ~new_P2_U3829;
  assign new_P2_U5484 = ~new_P2_U3391 | ~new_P2_U3889;
  assign new_P2_U5485 = ~new_P2_U3392;
  assign new_P2_U5486 = ~P2_REG0_REG_1_ | ~new_P2_U3831;
  assign new_P2_U5487 = ~new_P2_U3910 | ~new_P2_U4098;
  assign new_P2_U5488 = ~P2_IR_REG_2_ | ~new_P2_U3827;
  assign new_P2_U5489 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U23;
  assign new_P2_U5490 = ~new_U34 | ~new_P2_U3829;
  assign new_P2_U5491 = ~new_P2_U3394 | ~new_P2_U3889;
  assign new_P2_U5492 = ~new_P2_U3395;
  assign new_P2_U5493 = ~P2_REG0_REG_2_ | ~new_P2_U3831;
  assign new_P2_U5494 = ~new_P2_U3910 | ~new_P2_U4116;
  assign new_P2_U5495 = ~P2_IR_REG_3_ | ~new_P2_U3827;
  assign new_P2_U5496 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U24;
  assign new_P2_U5497 = ~new_U31 | ~new_P2_U3829;
  assign new_P2_U5498 = ~new_P2_U3397 | ~new_P2_U3889;
  assign new_P2_U5499 = ~new_P2_U3398;
  assign new_P2_U5500 = ~P2_REG0_REG_3_ | ~new_P2_U3831;
  assign new_P2_U5501 = ~new_P2_U3910 | ~new_P2_U4134;
  assign new_P2_U5502 = ~P2_IR_REG_4_ | ~new_P2_U3827;
  assign new_P2_U5503 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U25;
  assign new_P2_U5504 = ~new_U30 | ~new_P2_U3829;
  assign new_P2_U5505 = ~new_P2_U3400 | ~new_P2_U3889;
  assign new_P2_U5506 = ~new_P2_U3401;
  assign new_P2_U5507 = ~P2_REG0_REG_4_ | ~new_P2_U3831;
  assign new_P2_U5508 = ~new_P2_U3910 | ~new_P2_U4152;
  assign new_P2_U5509 = ~P2_IR_REG_5_ | ~new_P2_U3827;
  assign new_P2_U5510 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U72;
  assign new_P2_U5511 = ~new_U29 | ~new_P2_U3829;
  assign new_P2_U5512 = ~new_P2_U3403 | ~new_P2_U3889;
  assign new_P2_U5513 = ~new_P2_U3404;
  assign new_P2_U5514 = ~P2_REG0_REG_5_ | ~new_P2_U3831;
  assign new_P2_U5515 = ~new_P2_U3910 | ~new_P2_U4170;
  assign new_P2_U5516 = ~P2_IR_REG_6_ | ~new_P2_U3827;
  assign new_P2_U5517 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U26;
  assign new_P2_U5518 = ~new_U28 | ~new_P2_U3829;
  assign new_P2_U5519 = ~new_P2_U3406 | ~new_P2_U3889;
  assign new_P2_U5520 = ~new_P2_U3407;
  assign new_P2_U5521 = ~P2_REG0_REG_6_ | ~new_P2_U3831;
  assign new_P2_U5522 = ~new_P2_U3910 | ~new_P2_U4188;
  assign new_P2_U5523 = ~P2_IR_REG_7_ | ~new_P2_U3827;
  assign new_P2_U5524 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U27;
  assign new_P2_U5525 = ~new_U27 | ~new_P2_U3829;
  assign new_P2_U5526 = ~new_P2_U3409 | ~new_P2_U3889;
  assign new_P2_U5527 = ~new_P2_U3410;
  assign new_P2_U5528 = ~P2_REG0_REG_7_ | ~new_P2_U3831;
  assign new_P2_U5529 = ~new_P2_U3910 | ~new_P2_U4206;
  assign new_P2_U5530 = ~P2_IR_REG_8_ | ~new_P2_U3827;
  assign new_P2_U5531 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U28;
  assign new_P2_U5532 = ~new_U26 | ~new_P2_U3829;
  assign new_P2_U5533 = ~new_P2_U3412 | ~new_P2_U3889;
  assign new_P2_U5534 = ~new_P2_U3413;
  assign new_P2_U5535 = ~P2_REG0_REG_8_ | ~new_P2_U3831;
  assign new_P2_U5536 = ~new_P2_U3910 | ~new_P2_U4224;
  assign new_P2_U5537 = ~P2_IR_REG_9_ | ~new_P2_U3827;
  assign new_P2_U5538 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U70;
  assign new_P2_U5539 = ~new_U25 | ~new_P2_U3829;
  assign new_P2_U5540 = ~new_P2_U3415 | ~new_P2_U3889;
  assign new_P2_U5541 = ~new_P2_U3416;
  assign new_P2_U5542 = ~P2_REG0_REG_9_ | ~new_P2_U3831;
  assign new_P2_U5543 = ~new_P2_U3910 | ~new_P2_U4242;
  assign new_P2_U5544 = ~P2_IR_REG_10_ | ~new_P2_U3827;
  assign new_P2_U5545 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U8;
  assign new_P2_U5546 = ~new_U55 | ~new_P2_U3829;
  assign new_P2_U5547 = ~new_P2_U3418 | ~new_P2_U3889;
  assign new_P2_U5548 = ~new_P2_U3419;
  assign new_P2_U5549 = ~P2_REG0_REG_10_ | ~new_P2_U3831;
  assign new_P2_U5550 = ~new_P2_U3910 | ~new_P2_U4260;
  assign new_P2_U5551 = ~P2_IR_REG_11_ | ~new_P2_U3827;
  assign new_P2_U5552 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U9;
  assign new_P2_U5553 = ~new_U54 | ~new_P2_U3829;
  assign new_P2_U5554 = ~new_P2_U3421 | ~new_P2_U3889;
  assign new_P2_U5555 = ~new_P2_U3422;
  assign new_P2_U5556 = ~P2_REG0_REG_11_ | ~new_P2_U3831;
  assign new_P2_U5557 = ~new_P2_U3910 | ~new_P2_U4278;
  assign new_P2_U5558 = ~P2_IR_REG_12_ | ~new_P2_U3827;
  assign new_P2_U5559 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U10;
  assign new_P2_U5560 = ~new_U53 | ~new_P2_U3829;
  assign new_P2_U5561 = ~new_P2_U3424 | ~new_P2_U3889;
  assign new_P2_U5562 = ~new_P2_U3425;
  assign new_P2_U5563 = ~P2_REG0_REG_12_ | ~new_P2_U3831;
  assign new_P2_U5564 = ~new_P2_U3910 | ~new_P2_U4296;
  assign new_P2_U5565 = ~P2_IR_REG_13_ | ~new_P2_U3827;
  assign new_P2_U5566 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U87;
  assign new_P2_U5567 = ~new_U52 | ~new_P2_U3829;
  assign new_P2_U5568 = ~new_P2_U3427 | ~new_P2_U3889;
  assign new_P2_U5569 = ~new_P2_U3428;
  assign new_P2_U5570 = ~P2_REG0_REG_13_ | ~new_P2_U3831;
  assign new_P2_U5571 = ~new_P2_U3910 | ~new_P2_U4314;
  assign new_P2_U5572 = ~P2_IR_REG_14_ | ~new_P2_U3827;
  assign new_P2_U5573 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U11;
  assign new_P2_U5574 = ~new_U51 | ~new_P2_U3829;
  assign new_P2_U5575 = ~new_P2_U3430 | ~new_P2_U3889;
  assign new_P2_U5576 = ~new_P2_U3431;
  assign new_P2_U5577 = ~P2_REG0_REG_14_ | ~new_P2_U3831;
  assign new_P2_U5578 = ~new_P2_U3910 | ~new_P2_U4332;
  assign new_P2_U5579 = ~P2_IR_REG_15_ | ~new_P2_U3827;
  assign new_P2_U5580 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U12;
  assign new_P2_U5581 = ~new_U50 | ~new_P2_U3829;
  assign new_P2_U5582 = ~new_P2_U3433 | ~new_P2_U3889;
  assign new_P2_U5583 = ~new_P2_U3434;
  assign new_P2_U5584 = ~P2_REG0_REG_15_ | ~new_P2_U3831;
  assign new_P2_U5585 = ~new_P2_U3910 | ~new_P2_U4350;
  assign new_P2_U5586 = ~P2_IR_REG_16_ | ~new_P2_U3827;
  assign new_P2_U5587 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U13;
  assign new_P2_U5588 = ~new_U49 | ~new_P2_U3829;
  assign new_P2_U5589 = ~new_P2_U3436 | ~new_P2_U3889;
  assign new_P2_U5590 = ~new_P2_U3437;
  assign new_P2_U5591 = ~P2_REG0_REG_16_ | ~new_P2_U3831;
  assign new_P2_U5592 = ~new_P2_U3910 | ~new_P2_U4368;
  assign new_P2_U5593 = ~P2_IR_REG_17_ | ~new_P2_U3827;
  assign new_P2_U5594 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U85;
  assign new_P2_U5595 = ~new_U48 | ~new_P2_U3829;
  assign new_P2_U5596 = ~new_P2_U3439 | ~new_P2_U3889;
  assign new_P2_U5597 = ~new_P2_U3440;
  assign new_P2_U5598 = ~P2_REG0_REG_17_ | ~new_P2_U3831;
  assign new_P2_U5599 = ~new_P2_U3910 | ~new_P2_U4386;
  assign new_P2_U5600 = ~P2_IR_REG_18_ | ~new_P2_U3827;
  assign new_P2_U5601 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U14;
  assign new_P2_U5602 = ~new_U47 | ~new_P2_U3829;
  assign new_P2_U5603 = ~new_P2_U3442 | ~new_P2_U3889;
  assign new_P2_U5604 = ~new_P2_U3443;
  assign new_P2_U5605 = ~P2_REG0_REG_18_ | ~new_P2_U3831;
  assign new_P2_U5606 = ~new_P2_U3910 | ~new_P2_U4404;
  assign new_P2_U5607 = ~new_U46 | ~new_P2_U3829;
  assign new_P2_U5608 = ~new_P2_U3889 | ~new_P2_U3379;
  assign new_P2_U5609 = ~new_P2_U3445;
  assign new_P2_U5610 = ~P2_REG0_REG_19_ | ~new_P2_U3831;
  assign new_P2_U5611 = ~new_P2_U3910 | ~new_P2_U4422;
  assign new_P2_U5612 = ~P2_REG0_REG_20_ | ~new_P2_U3831;
  assign new_P2_U5613 = ~new_P2_U3910 | ~new_P2_U4440;
  assign new_P2_U5614 = ~P2_REG0_REG_21_ | ~new_P2_U3831;
  assign new_P2_U5615 = ~new_P2_U3910 | ~new_P2_U4458;
  assign new_P2_U5616 = ~P2_REG0_REG_22_ | ~new_P2_U3831;
  assign new_P2_U5617 = ~new_P2_U3910 | ~new_P2_U4476;
  assign new_P2_U5618 = ~P2_REG0_REG_23_ | ~new_P2_U3831;
  assign new_P2_U5619 = ~new_P2_U3910 | ~new_P2_U4494;
  assign new_P2_U5620 = ~P2_REG0_REG_24_ | ~new_P2_U3831;
  assign new_P2_U5621 = ~new_P2_U3910 | ~new_P2_U4512;
  assign new_P2_U5622 = ~P2_REG0_REG_25_ | ~new_P2_U3831;
  assign new_P2_U5623 = ~new_P2_U3910 | ~new_P2_U4530;
  assign new_P2_U5624 = ~P2_REG0_REG_26_ | ~new_P2_U3831;
  assign new_P2_U5625 = ~new_P2_U3910 | ~new_P2_U4548;
  assign new_P2_U5626 = ~P2_REG0_REG_27_ | ~new_P2_U3831;
  assign new_P2_U5627 = ~new_P2_U3910 | ~new_P2_U4566;
  assign new_P2_U5628 = ~P2_REG0_REG_28_ | ~new_P2_U3831;
  assign new_P2_U5629 = ~new_P2_U3910 | ~new_P2_U4584;
  assign new_P2_U5630 = ~P2_REG0_REG_29_ | ~new_P2_U3831;
  assign new_P2_U5631 = ~new_P2_U3910 | ~new_P2_U4604;
  assign new_P2_U5632 = ~P2_REG0_REG_30_ | ~new_P2_U3831;
  assign new_P2_U5633 = ~new_P2_U3910 | ~new_P2_U4611;
  assign new_P2_U5634 = ~P2_REG0_REG_31_ | ~new_P2_U3831;
  assign new_P2_U5635 = ~new_P2_U3910 | ~new_P2_U4613;
  assign new_P2_U5636 = ~new_P2_U5449 | ~new_P2_U3830;
  assign new_P2_U5637 = ~new_P2_U4048 | ~new_P2_U5446;
  assign new_P2_U5638 = ~P2_REG1_REG_0_ | ~new_P2_U3832;
  assign new_P2_U5639 = ~new_P2_U3909 | ~new_P2_U4073;
  assign new_P2_U5640 = ~P2_REG1_REG_1_ | ~new_P2_U3832;
  assign new_P2_U5641 = ~new_P2_U3909 | ~new_P2_U4098;
  assign new_P2_U5642 = ~P2_REG1_REG_2_ | ~new_P2_U3832;
  assign new_P2_U5643 = ~new_P2_U3909 | ~new_P2_U4116;
  assign new_P2_U5644 = ~P2_REG1_REG_3_ | ~new_P2_U3832;
  assign new_P2_U5645 = ~new_P2_U3909 | ~new_P2_U4134;
  assign new_P2_U5646 = ~P2_REG1_REG_4_ | ~new_P2_U3832;
  assign new_P2_U5647 = ~new_P2_U3909 | ~new_P2_U4152;
  assign new_P2_U5648 = ~P2_REG1_REG_5_ | ~new_P2_U3832;
  assign new_P2_U5649 = ~new_P2_U3909 | ~new_P2_U4170;
  assign new_P2_U5650 = ~P2_REG1_REG_6_ | ~new_P2_U3832;
  assign new_P2_U5651 = ~new_P2_U3909 | ~new_P2_U4188;
  assign new_P2_U5652 = ~P2_REG1_REG_7_ | ~new_P2_U3832;
  assign new_P2_U5653 = ~new_P2_U3909 | ~new_P2_U4206;
  assign new_P2_U5654 = ~P2_REG1_REG_8_ | ~new_P2_U3832;
  assign new_P2_U5655 = ~new_P2_U3909 | ~new_P2_U4224;
  assign new_P2_U5656 = ~P2_REG1_REG_9_ | ~new_P2_U3832;
  assign new_P2_U5657 = ~new_P2_U3909 | ~new_P2_U4242;
  assign new_P2_U5658 = ~P2_REG1_REG_10_ | ~new_P2_U3832;
  assign new_P2_U5659 = ~new_P2_U3909 | ~new_P2_U4260;
  assign new_P2_U5660 = ~P2_REG1_REG_11_ | ~new_P2_U3832;
  assign new_P2_U5661 = ~new_P2_U3909 | ~new_P2_U4278;
  assign new_P2_U5662 = ~P2_REG1_REG_12_ | ~new_P2_U3832;
  assign new_P2_U5663 = ~new_P2_U3909 | ~new_P2_U4296;
  assign new_P2_U5664 = ~P2_REG1_REG_13_ | ~new_P2_U3832;
  assign new_P2_U5665 = ~new_P2_U3909 | ~new_P2_U4314;
  assign new_P2_U5666 = ~P2_REG1_REG_14_ | ~new_P2_U3832;
  assign new_P2_U5667 = ~new_P2_U3909 | ~new_P2_U4332;
  assign new_P2_U5668 = ~P2_REG1_REG_15_ | ~new_P2_U3832;
  assign new_P2_U5669 = ~new_P2_U3909 | ~new_P2_U4350;
  assign new_P2_U5670 = ~P2_REG1_REG_16_ | ~new_P2_U3832;
  assign new_P2_U5671 = ~new_P2_U3909 | ~new_P2_U4368;
  assign new_P2_U5672 = ~P2_REG1_REG_17_ | ~new_P2_U3832;
  assign new_P2_U5673 = ~new_P2_U3909 | ~new_P2_U4386;
  assign new_P2_U5674 = ~P2_REG1_REG_18_ | ~new_P2_U3832;
  assign new_P2_U5675 = ~new_P2_U3909 | ~new_P2_U4404;
  assign new_P2_U5676 = ~P2_REG1_REG_19_ | ~new_P2_U3832;
  assign new_P2_U5677 = ~new_P2_U3909 | ~new_P2_U4422;
  assign new_P2_U5678 = ~P2_REG1_REG_20_ | ~new_P2_U3832;
  assign new_P2_U5679 = ~new_P2_U3909 | ~new_P2_U4440;
  assign new_P2_U5680 = ~P2_REG1_REG_21_ | ~new_P2_U3832;
  assign new_P2_U5681 = ~new_P2_U3909 | ~new_P2_U4458;
  assign new_P2_U5682 = ~P2_REG1_REG_22_ | ~new_P2_U3832;
  assign new_P2_U5683 = ~new_P2_U3909 | ~new_P2_U4476;
  assign new_P2_U5684 = ~P2_REG1_REG_23_ | ~new_P2_U3832;
  assign new_P2_U5685 = ~new_P2_U3909 | ~new_P2_U4494;
  assign new_P2_U5686 = ~P2_REG1_REG_24_ | ~new_P2_U3832;
  assign new_P2_U5687 = ~new_P2_U3909 | ~new_P2_U4512;
  assign new_P2_U5688 = ~P2_REG1_REG_25_ | ~new_P2_U3832;
  assign new_P2_U5689 = ~new_P2_U3909 | ~new_P2_U4530;
  assign new_P2_U5690 = ~P2_REG1_REG_26_ | ~new_P2_U3832;
  assign new_P2_U5691 = ~new_P2_U3909 | ~new_P2_U4548;
  assign new_P2_U5692 = ~P2_REG1_REG_27_ | ~new_P2_U3832;
  assign new_P2_U5693 = ~new_P2_U3909 | ~new_P2_U4566;
  assign new_P2_U5694 = ~P2_REG1_REG_28_ | ~new_P2_U3832;
  assign new_P2_U5695 = ~new_P2_U3909 | ~new_P2_U4584;
  assign new_P2_U5696 = ~P2_REG1_REG_29_ | ~new_P2_U3832;
  assign new_P2_U5697 = ~new_P2_U3909 | ~new_P2_U4604;
  assign new_P2_U5698 = ~P2_REG1_REG_30_ | ~new_P2_U3832;
  assign new_P2_U5699 = ~new_P2_U3909 | ~new_P2_U4611;
  assign new_P2_U5700 = ~P2_REG1_REG_31_ | ~new_P2_U3832;
  assign new_P2_U5701 = ~new_P2_U3909 | ~new_P2_U4613;
  assign new_P2_U5702 = ~P2_REG2_REG_0_ | ~new_P2_U3358;
  assign new_P2_U5703 = ~new_P2_U3908 | ~new_P2_U3314;
  assign new_P2_U5704 = ~P2_REG2_REG_1_ | ~new_P2_U3358;
  assign new_P2_U5705 = ~new_P2_U3908 | ~new_P2_U3315;
  assign new_P2_U5706 = ~P2_REG2_REG_2_ | ~new_P2_U3358;
  assign new_P2_U5707 = ~new_P2_U3908 | ~new_P2_U3316;
  assign new_P2_U5708 = ~P2_REG2_REG_3_ | ~new_P2_U3358;
  assign new_P2_U5709 = ~new_P2_U3908 | ~new_P2_U3317;
  assign new_P2_U5710 = ~P2_REG2_REG_4_ | ~new_P2_U3358;
  assign new_P2_U5711 = ~new_P2_U3908 | ~new_P2_U3318;
  assign new_P2_U5712 = ~P2_REG2_REG_5_ | ~new_P2_U3358;
  assign new_P2_U5713 = ~new_P2_U3908 | ~new_P2_U3319;
  assign new_P2_U5714 = ~P2_REG2_REG_6_ | ~new_P2_U3358;
  assign new_P2_U5715 = ~new_P2_U3908 | ~new_P2_U3320;
  assign new_P2_U5716 = ~P2_REG2_REG_7_ | ~new_P2_U3358;
  assign new_P2_U5717 = ~new_P2_U3908 | ~new_P2_U3321;
  assign new_P2_U5718 = ~P2_REG2_REG_8_ | ~new_P2_U3358;
  assign new_P2_U5719 = ~new_P2_U3908 | ~new_P2_U3322;
  assign new_P2_U5720 = ~P2_REG2_REG_9_ | ~new_P2_U3358;
  assign new_P2_U5721 = ~new_P2_U3908 | ~new_P2_U3323;
  assign new_P2_U5722 = ~P2_REG2_REG_10_ | ~new_P2_U3358;
  assign new_P2_U5723 = ~new_P2_U3908 | ~new_P2_U3324;
  assign new_P2_U5724 = ~P2_REG2_REG_11_ | ~new_P2_U3358;
  assign new_P2_U5725 = ~new_P2_U3908 | ~new_P2_U3325;
  assign new_P2_U5726 = ~P2_REG2_REG_12_ | ~new_P2_U3358;
  assign new_P2_U5727 = ~new_P2_U3908 | ~new_P2_U3326;
  assign new_P2_U5728 = ~P2_REG2_REG_13_ | ~new_P2_U3358;
  assign new_P2_U5729 = ~new_P2_U3908 | ~new_P2_U3327;
  assign new_P2_U5730 = ~P2_REG2_REG_14_ | ~new_P2_U3358;
  assign new_P2_U5731 = ~new_P2_U3908 | ~new_P2_U3328;
  assign new_P2_U5732 = ~P2_REG2_REG_15_ | ~new_P2_U3358;
  assign new_P2_U5733 = ~new_P2_U3908 | ~new_P2_U3329;
  assign new_P2_U5734 = ~P2_REG2_REG_16_ | ~new_P2_U3358;
  assign new_P2_U5735 = ~new_P2_U3908 | ~new_P2_U3330;
  assign new_P2_U5736 = ~P2_REG2_REG_17_ | ~new_P2_U3358;
  assign new_P2_U5737 = ~new_P2_U3908 | ~new_P2_U3331;
  assign new_P2_U5738 = ~P2_REG2_REG_18_ | ~new_P2_U3358;
  assign new_P2_U5739 = ~new_P2_U3908 | ~new_P2_U3332;
  assign new_P2_U5740 = ~P2_REG2_REG_19_ | ~new_P2_U3358;
  assign new_P2_U5741 = ~new_P2_U3908 | ~new_P2_U3333;
  assign new_P2_U5742 = ~P2_REG2_REG_20_ | ~new_P2_U3358;
  assign new_P2_U5743 = ~new_P2_U3908 | ~new_P2_U3335;
  assign new_P2_U5744 = ~P2_REG2_REG_21_ | ~new_P2_U3358;
  assign new_P2_U5745 = ~new_P2_U3908 | ~new_P2_U3337;
  assign new_P2_U5746 = ~P2_REG2_REG_22_ | ~new_P2_U3358;
  assign new_P2_U5747 = ~new_P2_U3908 | ~new_P2_U3339;
  assign new_P2_U5748 = ~P2_REG2_REG_23_ | ~new_P2_U3358;
  assign new_P2_U5749 = ~new_P2_U3908 | ~new_P2_U3341;
  assign new_P2_U5750 = ~P2_REG2_REG_24_ | ~new_P2_U3358;
  assign new_P2_U5751 = ~new_P2_U3908 | ~new_P2_U3343;
  assign new_P2_U5752 = ~P2_REG2_REG_25_ | ~new_P2_U3358;
  assign new_P2_U5753 = ~new_P2_U3908 | ~new_P2_U3345;
  assign new_P2_U5754 = ~P2_REG2_REG_26_ | ~new_P2_U3358;
  assign new_P2_U5755 = ~new_P2_U3908 | ~new_P2_U3347;
  assign new_P2_U5756 = ~P2_REG2_REG_27_ | ~new_P2_U3358;
  assign new_P2_U5757 = ~new_P2_U3908 | ~new_P2_U3349;
  assign new_P2_U5758 = ~P2_REG2_REG_28_ | ~new_P2_U3358;
  assign new_P2_U5759 = ~new_P2_U3908 | ~new_P2_U3351;
  assign new_P2_U5760 = ~P2_REG2_REG_29_ | ~new_P2_U3358;
  assign new_P2_U5761 = ~new_P2_U3908 | ~new_P2_U3354;
  assign new_P2_U5762 = ~new_P2_U5461 | ~new_P2_U3024;
  assign new_P2_U5763 = ~new_P2_U3383 | ~n2565;
  assign new_P2_U5764 = ~new_P2_U5763 | ~new_P2_U5762;
  assign new_P2_U5765 = ~P2_DATAO_REG_0_ | ~new_P2_U3363;
  assign new_P2_U5766 = ~n2565 | ~new_P2_U3076;
  assign new_P2_U5767 = ~P2_DATAO_REG_1_ | ~new_P2_U3363;
  assign new_P2_U5768 = ~n2565 | ~new_P2_U3077;
  assign new_P2_U5769 = ~P2_DATAO_REG_2_ | ~new_P2_U3363;
  assign new_P2_U5770 = ~n2565 | ~new_P2_U3067;
  assign new_P2_U5771 = ~P2_DATAO_REG_3_ | ~new_P2_U3363;
  assign new_P2_U5772 = ~n2565 | ~new_P2_U3063;
  assign new_P2_U5773 = ~P2_DATAO_REG_4_ | ~new_P2_U3363;
  assign new_P2_U5774 = ~n2565 | ~new_P2_U3059;
  assign new_P2_U5775 = ~P2_DATAO_REG_5_ | ~new_P2_U3363;
  assign new_P2_U5776 = ~n2565 | ~new_P2_U3066;
  assign new_P2_U5777 = ~P2_DATAO_REG_6_ | ~new_P2_U3363;
  assign new_P2_U5778 = ~n2565 | ~new_P2_U3070;
  assign new_P2_U5779 = ~P2_DATAO_REG_7_ | ~new_P2_U3363;
  assign new_P2_U5780 = ~n2565 | ~new_P2_U3069;
  assign new_P2_U5781 = ~P2_DATAO_REG_8_ | ~new_P2_U3363;
  assign new_P2_U5782 = ~n2565 | ~new_P2_U3083;
  assign new_P2_U5783 = ~P2_DATAO_REG_9_ | ~new_P2_U3363;
  assign new_P2_U5784 = ~n2565 | ~new_P2_U3082;
  assign new_P2_U5785 = ~P2_DATAO_REG_10_ | ~new_P2_U3363;
  assign new_P2_U5786 = ~n2565 | ~new_P2_U3061;
  assign new_P2_U5787 = ~P2_DATAO_REG_11_ | ~new_P2_U3363;
  assign new_P2_U5788 = ~n2565 | ~new_P2_U3062;
  assign new_P2_U5789 = ~P2_DATAO_REG_12_ | ~new_P2_U3363;
  assign new_P2_U5790 = ~n2565 | ~new_P2_U3071;
  assign new_P2_U5791 = ~P2_DATAO_REG_13_ | ~new_P2_U3363;
  assign new_P2_U5792 = ~n2565 | ~new_P2_U3079;
  assign new_P2_U5793 = ~P2_DATAO_REG_14_ | ~new_P2_U3363;
  assign new_P2_U5794 = ~n2565 | ~new_P2_U3078;
  assign new_P2_U5795 = ~P2_DATAO_REG_15_ | ~new_P2_U3363;
  assign new_P2_U5796 = ~n2565 | ~new_P2_U3073;
  assign new_P2_U5797 = ~P2_DATAO_REG_16_ | ~new_P2_U3363;
  assign new_P2_U5798 = ~n2565 | ~new_P2_U3072;
  assign new_P2_U5799 = ~P2_DATAO_REG_17_ | ~new_P2_U3363;
  assign new_P2_U5800 = ~n2565 | ~new_P2_U3068;
  assign new_P2_U5801 = ~P2_DATAO_REG_18_ | ~new_P2_U3363;
  assign new_P2_U5802 = ~n2565 | ~new_P2_U3081;
  assign new_P2_U5803 = ~P2_DATAO_REG_19_ | ~new_P2_U3363;
  assign new_P2_U5804 = ~n2565 | ~new_P2_U3080;
  assign new_P2_U5805 = ~P2_DATAO_REG_20_ | ~new_P2_U3363;
  assign new_P2_U5806 = ~n2565 | ~new_P2_U3075;
  assign new_P2_U5807 = ~P2_DATAO_REG_21_ | ~new_P2_U3363;
  assign new_P2_U5808 = ~n2565 | ~new_P2_U3074;
  assign new_P2_U5809 = ~P2_DATAO_REG_22_ | ~new_P2_U3363;
  assign new_P2_U5810 = ~n2565 | ~new_P2_U3060;
  assign new_P2_U5811 = ~P2_DATAO_REG_23_ | ~new_P2_U3363;
  assign new_P2_U5812 = ~n2565 | ~new_P2_U3065;
  assign new_P2_U5813 = ~P2_DATAO_REG_24_ | ~new_P2_U3363;
  assign new_P2_U5814 = ~n2565 | ~new_P2_U3064;
  assign new_P2_U5815 = ~P2_DATAO_REG_25_ | ~new_P2_U3363;
  assign new_P2_U5816 = ~n2565 | ~new_P2_U3057;
  assign new_P2_U5817 = ~P2_DATAO_REG_26_ | ~new_P2_U3363;
  assign new_P2_U5818 = ~n2565 | ~new_P2_U3056;
  assign new_P2_U5819 = ~P2_DATAO_REG_27_ | ~new_P2_U3363;
  assign new_P2_U5820 = ~n2565 | ~new_P2_U3052;
  assign new_P2_U5821 = ~P2_DATAO_REG_28_ | ~new_P2_U3363;
  assign new_P2_U5822 = ~n2565 | ~new_P2_U3053;
  assign new_P2_U5823 = ~P2_DATAO_REG_29_ | ~new_P2_U3363;
  assign new_P2_U5824 = ~n2565 | ~new_P2_U3054;
  assign new_P2_U5825 = ~P2_DATAO_REG_30_ | ~new_P2_U3363;
  assign new_P2_U5826 = ~n2565 | ~new_P2_U3058;
  assign new_P2_U5827 = ~P2_DATAO_REG_31_ | ~new_P2_U3363;
  assign new_P2_U5828 = ~n2565 | ~new_P2_U3055;
  assign new_P2_U5829 = ~new_P2_U3379 | ~new_P2_U3313;
  assign new_P2_U5830 = ~new_P2_U5446 | ~new_P2_U3907;
  assign new_P2_U5831 = ~new_P2_U3765;
  assign new_P2_U5832 = ~new_P2_R1269_U22 | ~new_P2_U5831;
  assign new_P2_U5833 = ~new_P2_U3765 | ~new_P2_U3863;
  assign new_P2_U5834 = ~new_P2_U3896 | ~new_P2_U3052;
  assign new_P2_U5835 = ~new_P2_U3348 | ~new_P2_U4535;
  assign new_P2_U5836 = ~new_P2_U5835 | ~new_P2_U5834;
  assign new_P2_U5837 = ~new_P2_U3895 | ~new_P2_U3053;
  assign new_P2_U5838 = ~new_P2_U3350 | ~new_P2_U4553;
  assign new_P2_U5839 = ~new_P2_U5838 | ~new_P2_U5837;
  assign new_P2_U5840 = ~new_P2_U3868 | ~new_P2_U3055;
  assign new_P2_U5841 = ~new_P2_U3356 | ~new_P2_U4609;
  assign new_P2_U5842 = ~new_P2_U5841 | ~new_P2_U5840;
  assign new_P2_U5843 = ~new_P2_U3904 | ~new_P2_U3054;
  assign new_P2_U5844 = ~new_P2_U3353 | ~new_P2_U4571;
  assign new_P2_U5845 = ~new_P2_U5844 | ~new_P2_U5843;
  assign new_P2_U5846 = ~new_P2_U3902 | ~new_P2_U3074;
  assign new_P2_U5847 = ~new_P2_U3336 | ~new_P2_U4427;
  assign new_P2_U5848 = ~new_P2_U5847 | ~new_P2_U5846;
  assign new_P2_U5849 = ~new_P2_U3903 | ~new_P2_U3075;
  assign new_P2_U5850 = ~new_P2_U3334 | ~new_P2_U4409;
  assign new_P2_U5851 = ~new_P2_U5850 | ~new_P2_U5849;
  assign new_P2_U5852 = ~new_P2_U5499 | ~new_P2_U4103;
  assign new_P2_U5853 = ~new_P2_U3398 | ~new_P2_U3063;
  assign new_P2_U5854 = ~new_P2_U5853 | ~new_P2_U5852;
  assign new_P2_U5855 = ~new_P2_U5555 | ~new_P2_U4247;
  assign new_P2_U5856 = ~new_P2_U3422 | ~new_P2_U3062;
  assign new_P2_U5857 = ~new_P2_U5856 | ~new_P2_U5855;
  assign new_P2_U5858 = ~new_P2_U5548 | ~new_P2_U4229;
  assign new_P2_U5859 = ~new_P2_U3419 | ~new_P2_U3061;
  assign new_P2_U5860 = ~new_P2_U5859 | ~new_P2_U5858;
  assign new_P2_U5861 = ~new_P2_U5506 | ~new_P2_U4121;
  assign new_P2_U5862 = ~new_P2_U3401 | ~new_P2_U3059;
  assign new_P2_U5863 = ~new_P2_U5862 | ~new_P2_U5861;
  assign new_P2_U5864 = ~new_P2_U3901 | ~new_P2_U3060;
  assign new_P2_U5865 = ~new_P2_U3338 | ~new_P2_U4445;
  assign new_P2_U5866 = ~new_P2_U5865 | ~new_P2_U5864;
  assign new_P2_U5867 = ~new_P2_U5597 | ~new_P2_U4355;
  assign new_P2_U5868 = ~new_P2_U3440 | ~new_P2_U3068;
  assign new_P2_U5869 = ~new_P2_U5868 | ~new_P2_U5867;
  assign new_P2_U5870 = ~new_P2_U5583 | ~new_P2_U4319;
  assign new_P2_U5871 = ~new_P2_U3434 | ~new_P2_U3073;
  assign new_P2_U5872 = ~new_P2_U5871 | ~new_P2_U5870;
  assign new_P2_U5873 = ~new_P2_U5562 | ~new_P2_U4265;
  assign new_P2_U5874 = ~new_P2_U3425 | ~new_P2_U3071;
  assign new_P2_U5875 = ~new_P2_U5874 | ~new_P2_U5873;
  assign new_P2_U5876 = ~new_P2_U5520 | ~new_P2_U4157;
  assign new_P2_U5877 = ~new_P2_U3407 | ~new_P2_U3070;
  assign new_P2_U5878 = ~new_P2_U5877 | ~new_P2_U5876;
  assign new_P2_U5879 = ~new_P2_U5527 | ~new_P2_U4175;
  assign new_P2_U5880 = ~new_P2_U3410 | ~new_P2_U3069;
  assign new_P2_U5881 = ~new_P2_U5880 | ~new_P2_U5879;
  assign new_P2_U5882 = ~new_P2_U5492 | ~new_P2_U4078;
  assign new_P2_U5883 = ~new_P2_U3395 | ~new_P2_U3067;
  assign new_P2_U5884 = ~new_P2_U5883 | ~new_P2_U5882;
  assign new_P2_U5885 = ~new_P2_U5513 | ~new_P2_U4139;
  assign new_P2_U5886 = ~new_P2_U3404 | ~new_P2_U3066;
  assign new_P2_U5887 = ~new_P2_U5886 | ~new_P2_U5885;
  assign new_P2_U5888 = ~new_P2_U5590 | ~new_P2_U4337;
  assign new_P2_U5889 = ~new_P2_U3437 | ~new_P2_U3072;
  assign new_P2_U5890 = ~new_P2_U5889 | ~new_P2_U5888;
  assign new_P2_U5891 = ~new_P2_U5604 | ~new_P2_U4373;
  assign new_P2_U5892 = ~new_P2_U3443 | ~new_P2_U3081;
  assign new_P2_U5893 = ~new_P2_U5892 | ~new_P2_U5891;
  assign new_P2_U5894 = ~new_P2_U5569 | ~new_P2_U4283;
  assign new_P2_U5895 = ~new_P2_U3428 | ~new_P2_U3079;
  assign new_P2_U5896 = ~new_P2_U5895 | ~new_P2_U5894;
  assign new_P2_U5897 = ~new_P2_U5576 | ~new_P2_U4301;
  assign new_P2_U5898 = ~new_P2_U3431 | ~new_P2_U3078;
  assign new_P2_U5899 = ~new_P2_U5898 | ~new_P2_U5897;
  assign new_P2_U5900 = ~new_P2_U5485 | ~new_P2_U4059;
  assign new_P2_U5901 = ~new_P2_U3392 | ~new_P2_U3077;
  assign new_P2_U5902 = ~new_P2_U5901 | ~new_P2_U5900;
  assign new_P2_U5903 = ~new_P2_U5469 | ~new_P2_U4083;
  assign new_P2_U5904 = ~new_P2_U3387 | ~new_P2_U3076;
  assign new_P2_U5905 = ~new_P2_U5904 | ~new_P2_U5903;
  assign new_P2_U5906 = ~new_P2_U5534 | ~new_P2_U4193;
  assign new_P2_U5907 = ~new_P2_U3413 | ~new_P2_U3083;
  assign new_P2_U5908 = ~new_P2_U5907 | ~new_P2_U5906;
  assign new_P2_U5909 = ~new_P2_U5541 | ~new_P2_U4211;
  assign new_P2_U5910 = ~new_P2_U3416 | ~new_P2_U3082;
  assign new_P2_U5911 = ~new_P2_U5910 | ~new_P2_U5909;
  assign new_P2_U5912 = ~new_P2_U5609 | ~new_P2_U4391;
  assign new_P2_U5913 = ~new_P2_U3445 | ~new_P2_U3080;
  assign new_P2_U5914 = ~new_P2_U5913 | ~new_P2_U5912;
  assign new_P2_U5915 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_U5916 = ~new_P2_U3346 | ~new_P2_U4517;
  assign new_P2_U5917 = ~new_P2_U5916 | ~new_P2_U5915;
  assign new_P2_U5918 = ~new_P2_U3898 | ~new_P2_U3057;
  assign new_P2_U5919 = ~new_P2_U3344 | ~new_P2_U4499;
  assign new_P2_U5920 = ~new_P2_U5919 | ~new_P2_U5918;
  assign new_P2_U5921 = ~new_P2_U3900 | ~new_P2_U3065;
  assign new_P2_U5922 = ~new_P2_U3340 | ~new_P2_U4463;
  assign new_P2_U5923 = ~new_P2_U5922 | ~new_P2_U5921;
  assign new_P2_U5924 = ~new_P2_U3899 | ~new_P2_U3064;
  assign new_P2_U5925 = ~new_P2_U3342 | ~new_P2_U4481;
  assign new_P2_U5926 = ~new_P2_U5925 | ~new_P2_U5924;
  assign new_P2_U5927 = ~new_P2_U3869 | ~new_P2_U3058;
  assign new_P2_U5928 = ~new_P2_U3355 | ~new_P2_U4589;
  assign new_P2_U5929 = ~new_P2_U5928 | ~new_P2_U5927;
  assign new_P2_U5930 = ~new_P2_U4974 | ~new_P2_U5446;
  assign new_P2_U5931 = ~new_P2_U3379 | ~new_P2_U3864;
  assign new_P2_U5932 = ~new_P2_U5931 | ~new_P2_U5930;
  assign new_P2_U5933 = ~new_P2_U5443 | ~new_P2_U5833 | ~new_P2_U5832;
  assign new_P2_U5934 = ~new_P2_U3378 | ~new_P2_U5452 | ~new_P2_U5932;
  assign new_P2_U5935 = ~new_P2_U3877 | ~new_P2_U3865;
  assign new_P2_U5936 = ~new_P2_R693_U14 | ~new_P2_U3887;
  assign new_P2_U5937 = ~new_P2_U5436 | ~new_P2_U3368;
  assign new_P2_U5938 = ~new_P2_U3380 | ~new_P2_U3375;
  assign new_P2_U5939 = ~new_P2_U5446 | ~new_P2_U5443;
  assign new_P2_U5940 = ~new_P2_U3378 | ~new_P2_U3388 | ~new_P2_U5452;
  assign new_P2_U5941 = ~new_P2_U3082 | ~new_P2_R1297_U6;
  assign new_P2_U5942 = ~new_P2_U3082 | ~new_P2_U3867;
  assign new_P2_U5943 = ~new_P2_U3083 | ~new_P2_R1297_U6;
  assign new_P2_U5944 = ~new_P2_U3083 | ~new_P2_U3867;
  assign new_P2_U5945 = ~new_P2_U3069 | ~new_P2_R1297_U6;
  assign new_P2_U5946 = ~new_P2_U3069 | ~new_P2_U3867;
  assign new_P2_U5947 = ~new_P2_U3070 | ~new_P2_R1297_U6;
  assign new_P2_U5948 = ~new_P2_U3070 | ~new_P2_U3867;
  assign new_P2_U5949 = ~new_P2_U3066 | ~new_P2_R1297_U6;
  assign new_P2_U5950 = ~new_P2_U3066 | ~new_P2_U3867;
  assign new_P2_U5951 = ~new_P2_U3059 | ~new_P2_R1297_U6;
  assign new_P2_U5952 = ~new_P2_U3059 | ~new_P2_U3867;
  assign new_P2_U5953 = ~new_P2_R1300_U8 | ~new_P2_R1297_U6;
  assign new_P2_U5954 = ~new_P2_U3055 | ~new_P2_U3867;
  assign new_P2_U5955 = ~new_P2_R1300_U6 | ~new_P2_R1297_U6;
  assign new_P2_U5956 = ~new_P2_U3058 | ~new_P2_U3867;
  assign new_P2_U5957 = ~new_P2_U3063 | ~new_P2_R1297_U6;
  assign new_P2_U5958 = ~new_P2_U3063 | ~new_P2_U3867;
  assign new_P2_U5959 = ~new_P2_U3054 | ~new_P2_R1297_U6;
  assign new_P2_U5960 = ~new_P2_U3054 | ~new_P2_U3867;
  assign new_P2_U5961 = ~new_P2_U3053 | ~new_P2_R1297_U6;
  assign new_P2_U5962 = ~new_P2_U3053 | ~new_P2_U3867;
  assign new_P2_U5963 = ~new_P2_U3052 | ~new_P2_R1297_U6;
  assign new_P2_U5964 = ~new_P2_U3052 | ~new_P2_U3867;
  assign new_P2_U5965 = ~new_P2_U3056 | ~new_P2_R1297_U6;
  assign new_P2_U5966 = ~new_P2_U3056 | ~new_P2_U3867;
  assign new_P2_U5967 = ~new_P2_U3057 | ~new_P2_R1297_U6;
  assign new_P2_U5968 = ~new_P2_U3057 | ~new_P2_U3867;
  assign new_P2_U5969 = ~new_P2_U3064 | ~new_P2_R1297_U6;
  assign new_P2_U5970 = ~new_P2_U3064 | ~new_P2_U3867;
  assign new_P2_U5971 = ~new_P2_U3065 | ~new_P2_R1297_U6;
  assign new_P2_U5972 = ~new_P2_U3065 | ~new_P2_U3867;
  assign new_P2_U5973 = ~new_P2_U3060 | ~new_P2_R1297_U6;
  assign new_P2_U5974 = ~new_P2_U3060 | ~new_P2_U3867;
  assign new_P2_U5975 = ~new_P2_U3074 | ~new_P2_R1297_U6;
  assign new_P2_U5976 = ~new_P2_U3074 | ~new_P2_U3867;
  assign new_P2_U5977 = ~new_P2_U3075 | ~new_P2_R1297_U6;
  assign new_P2_U5978 = ~new_P2_U3075 | ~new_P2_U3867;
  assign new_P2_U5979 = ~new_P2_U3067 | ~new_P2_R1297_U6;
  assign new_P2_U5980 = ~new_P2_U3067 | ~new_P2_U3867;
  assign new_P2_U5981 = ~new_P2_U3080 | ~new_P2_R1297_U6;
  assign new_P2_U5982 = ~new_P2_U3080 | ~new_P2_U3867;
  assign new_P2_U5983 = ~new_P2_U3081 | ~new_P2_R1297_U6;
  assign new_P2_U5984 = ~new_P2_U3081 | ~new_P2_U3867;
  assign new_P2_U5985 = ~new_P2_U3068 | ~new_P2_R1297_U6;
  assign new_P2_U5986 = ~new_P2_U3068 | ~new_P2_U3867;
  assign new_P2_U5987 = ~new_P2_U3072 | ~new_P2_R1297_U6;
  assign new_P2_U5988 = ~new_P2_U3072 | ~new_P2_U3867;
  assign new_P2_U5989 = ~new_P2_U3073 | ~new_P2_R1297_U6;
  assign new_P2_U5990 = ~new_P2_U3073 | ~new_P2_U3867;
  assign new_P2_U5991 = ~new_P2_U3078 | ~new_P2_R1297_U6;
  assign new_P2_U5992 = ~new_P2_U3078 | ~new_P2_U3867;
  assign new_P2_U5993 = ~new_P2_U3079 | ~new_P2_R1297_U6;
  assign new_P2_U5994 = ~new_P2_U3079 | ~new_P2_U3867;
  assign new_P2_U5995 = ~new_P2_U3071 | ~new_P2_R1297_U6;
  assign new_P2_U5996 = ~new_P2_U3071 | ~new_P2_U3867;
  assign new_P2_U5997 = ~new_P2_U3062 | ~new_P2_R1297_U6;
  assign new_P2_U5998 = ~new_P2_U3062 | ~new_P2_U3867;
  assign new_P2_U5999 = ~new_P2_U3061 | ~new_P2_R1297_U6;
  assign new_P2_U6000 = ~new_P2_U3061 | ~new_P2_U3867;
  assign new_P2_U6001 = ~new_P2_U3077 | ~new_P2_R1297_U6;
  assign new_P2_U6002 = ~new_P2_U3077 | ~new_P2_U3867;
  assign new_P2_U6003 = ~new_P2_U3076 | ~new_P2_R1297_U6;
  assign new_P2_U6004 = ~new_P2_U3076 | ~new_P2_U3867;
  assign new_P2_U6005 = ~new_P2_U5464 | ~P2_REG1_REG_9_;
  assign new_P2_U6006 = ~new_P2_U3384 | ~P2_REG2_REG_9_;
  assign new_P2_U6007 = ~new_P2_U5464 | ~P2_REG1_REG_8_;
  assign new_P2_U6008 = ~new_P2_U3384 | ~P2_REG2_REG_8_;
  assign new_P2_U6009 = ~new_P2_U5464 | ~P2_REG1_REG_7_;
  assign new_P2_U6010 = ~new_P2_U3384 | ~P2_REG2_REG_7_;
  assign new_P2_U6011 = ~new_P2_U5464 | ~P2_REG1_REG_6_;
  assign new_P2_U6012 = ~new_P2_U3384 | ~P2_REG2_REG_6_;
  assign new_P2_U6013 = ~new_P2_U5464 | ~P2_REG1_REG_5_;
  assign new_P2_U6014 = ~new_P2_U3384 | ~P2_REG2_REG_5_;
  assign new_P2_U6015 = ~new_P2_U5464 | ~P2_REG1_REG_4_;
  assign new_P2_U6016 = ~new_P2_U3384 | ~P2_REG2_REG_4_;
  assign new_P2_U6017 = ~new_P2_U5464 | ~P2_REG1_REG_3_;
  assign new_P2_U6018 = ~new_P2_U3384 | ~P2_REG2_REG_3_;
  assign new_P2_U6019 = ~new_P2_U5464 | ~P2_REG1_REG_2_;
  assign new_P2_U6020 = ~new_P2_U3384 | ~P2_REG2_REG_2_;
  assign new_P2_U6021 = ~new_P2_U5464 | ~P2_REG1_REG_19_;
  assign new_P2_U6022 = ~new_P2_U3384 | ~P2_REG2_REG_19_;
  assign new_P2_U6023 = ~new_P2_U5464 | ~P2_REG1_REG_18_;
  assign new_P2_U6024 = ~new_P2_U3384 | ~P2_REG2_REG_18_;
  assign new_P2_U6025 = ~new_P2_U5464 | ~P2_REG1_REG_17_;
  assign new_P2_U6026 = ~new_P2_U3384 | ~P2_REG2_REG_17_;
  assign new_P2_U6027 = ~new_P2_U5464 | ~P2_REG1_REG_16_;
  assign new_P2_U6028 = ~new_P2_U3384 | ~P2_REG2_REG_16_;
  assign new_P2_U6029 = ~new_P2_U5464 | ~P2_REG1_REG_15_;
  assign new_P2_U6030 = ~new_P2_U3384 | ~P2_REG2_REG_15_;
  assign new_P2_U6031 = ~new_P2_U5464 | ~P2_REG1_REG_14_;
  assign new_P2_U6032 = ~new_P2_U3384 | ~P2_REG2_REG_14_;
  assign new_P2_U6033 = ~new_P2_U5464 | ~P2_REG1_REG_13_;
  assign new_P2_U6034 = ~new_P2_U3384 | ~P2_REG2_REG_13_;
  assign new_P2_U6035 = ~new_P2_U5464 | ~P2_REG1_REG_12_;
  assign new_P2_U6036 = ~new_P2_U3384 | ~P2_REG2_REG_12_;
  assign new_P2_U6037 = ~new_P2_U5464 | ~P2_REG1_REG_11_;
  assign new_P2_U6038 = ~new_P2_U3384 | ~P2_REG2_REG_11_;
  assign new_P2_U6039 = ~new_P2_U5464 | ~P2_REG1_REG_10_;
  assign new_P2_U6040 = ~new_P2_U3384 | ~P2_REG2_REG_10_;
  assign new_P2_U6041 = ~new_P2_U5464 | ~P2_REG1_REG_1_;
  assign new_P2_U6042 = ~new_P2_U3384 | ~P2_REG2_REG_1_;
  assign new_P2_U6043 = ~new_P2_U5464 | ~P2_REG1_REG_0_;
  assign new_P2_U6044 = ~new_P2_U3384 | ~P2_REG2_REG_0_;
  assign new_P2_R1161_U465 = ~new_P2_R1161_U464 | ~new_P2_R1161_U463;
  assign new_P2_R1161_U464 = ~new_P2_U3443 | ~new_P2_R1161_U76;
  assign new_P2_R1161_U463 = ~new_P2_U3081 | ~new_P2_R1161_U75;
  assign new_P2_R1161_U462 = ~new_P2_R1161_U460 | ~new_P2_R1161_U316;
  assign new_P2_R1161_U461 = ~new_P2_R1161_U359 | ~new_P2_R1161_U91;
  assign new_P2_R1161_U460 = ~new_P2_R1161_U459 | ~new_P2_R1161_U458;
  assign new_P2_R1161_U459 = ~new_P2_U3445 | ~new_P2_R1161_U79;
  assign new_P2_R1161_U458 = ~new_P2_U3080 | ~new_P2_R1161_U78;
  assign new_P2_R1161_U457 = ~new_P2_R1161_U328 | ~new_P2_R1161_U31;
  assign new_P2_R1161_U456 = ~new_P2_R1161_U182 | ~new_P2_R1161_U161;
  assign new_P2_R1161_U455 = ~new_P2_U3903 | ~new_P2_R1161_U90;
  assign new_P2_R1161_U454 = ~new_P2_U3075 | ~new_P2_R1161_U81;
  assign new_P2_R1161_U453 = ~new_P2_R1161_U452 | ~new_P2_R1161_U451;
  assign new_P2_R1161_U452 = ~new_P2_U3902 | ~new_P2_R1161_U55;
  assign new_P2_R1161_U451 = ~new_P2_U3074 | ~new_P2_R1161_U54;
  assign new_P2_R1161_U450 = ~new_P2_U3902 | ~new_P2_R1161_U55;
  assign new_P2_R1161_U449 = ~new_P2_U3074 | ~new_P2_R1161_U54;
  assign new_P2_R1161_U448 = ~new_P2_R1161_U286 | ~new_P2_R1161_U446;
  assign new_P2_R1161_U447 = ~new_P2_R1161_U158 | ~new_P2_R1161_U159;
  assign new_LT_1075_U6 = ~P1_ADDR_REG_19_;
  assign ADD_1068_U4 = new_ADD_1068_U159 & new_ADD_1068_U155;
  assign ADD_1068_U5 = ~new_ADD_1068_U160 | ~new_ADD_1068_U221 | ~new_ADD_1068_U220;
  assign new_ADD_1068_U6 = ~P1_ADDR_REG_0_;
  assign new_ADD_1068_U7 = ~P2_ADDR_REG_0_;
  assign new_ADD_1068_U8 = ~P2_ADDR_REG_1_;
  assign new_ADD_1068_U9 = ~P2_ADDR_REG_0_ | ~P1_ADDR_REG_0_;
  assign new_ADD_1068_U10 = ~P1_ADDR_REG_1_;
  assign new_ADD_1068_U11 = ~P1_ADDR_REG_2_;
  assign new_ADD_1068_U12 = ~P2_ADDR_REG_2_;
  assign new_ADD_1068_U13 = ~P1_ADDR_REG_3_;
  assign new_ADD_1068_U14 = ~P2_ADDR_REG_3_;
  assign new_ADD_1068_U15 = ~P1_ADDR_REG_4_;
  assign new_ADD_1068_U16 = ~P2_ADDR_REG_4_;
  assign new_ADD_1068_U17 = ~P1_ADDR_REG_5_;
  assign new_ADD_1068_U18 = ~P2_ADDR_REG_5_;
  assign new_ADD_1068_U19 = ~P1_ADDR_REG_6_;
  assign new_ADD_1068_U20 = ~P2_ADDR_REG_6_;
  assign new_ADD_1068_U21 = ~P1_ADDR_REG_7_;
  assign new_ADD_1068_U22 = ~P2_ADDR_REG_7_;
  assign new_ADD_1068_U23 = ~P1_ADDR_REG_8_;
  assign new_ADD_1068_U24 = ~P2_ADDR_REG_8_;
  assign new_ADD_1068_U25 = ~P2_ADDR_REG_9_;
  assign new_ADD_1068_U26 = ~P1_ADDR_REG_9_;
  assign new_ADD_1068_U27 = ~P1_ADDR_REG_10_;
  assign new_ADD_1068_U28 = ~P2_ADDR_REG_10_;
  assign new_ADD_1068_U29 = ~P1_ADDR_REG_11_;
  assign new_ADD_1068_U30 = ~P2_ADDR_REG_11_;
  assign new_ADD_1068_U31 = ~P1_ADDR_REG_12_;
  assign new_ADD_1068_U32 = ~P2_ADDR_REG_12_;
  assign new_ADD_1068_U33 = ~P1_ADDR_REG_13_;
  assign new_ADD_1068_U34 = ~P2_ADDR_REG_13_;
  assign new_ADD_1068_U35 = ~P1_ADDR_REG_14_;
  assign new_ADD_1068_U36 = ~P2_ADDR_REG_14_;
  assign new_ADD_1068_U37 = ~P1_ADDR_REG_15_;
  assign new_ADD_1068_U38 = ~P2_ADDR_REG_15_;
  assign new_ADD_1068_U39 = ~P1_ADDR_REG_16_;
  assign new_ADD_1068_U40 = ~P2_ADDR_REG_16_;
  assign new_ADD_1068_U41 = ~P1_ADDR_REG_17_;
  assign new_ADD_1068_U42 = ~P2_ADDR_REG_17_;
  assign new_ADD_1068_U43 = ~P1_ADDR_REG_18_;
  assign new_ADD_1068_U44 = ~P2_ADDR_REG_18_;
  assign new_ADD_1068_U45 = ~new_ADD_1068_U150 | ~new_ADD_1068_U149;
  assign ADD_1068_U46 = ~new_ADD_1068_U291 | ~new_ADD_1068_U290;
  assign ADD_1068_U47 = ~new_ADD_1068_U167 | ~new_ADD_1068_U166;
  assign ADD_1068_U48 = ~new_ADD_1068_U174 | ~new_ADD_1068_U173;
  assign ADD_1068_U49 = ~new_ADD_1068_U181 | ~new_ADD_1068_U180;
  assign ADD_1068_U50 = ~new_ADD_1068_U188 | ~new_ADD_1068_U187;
  assign ADD_1068_U51 = ~new_ADD_1068_U195 | ~new_ADD_1068_U194;
  assign ADD_1068_U52 = ~new_ADD_1068_U202 | ~new_ADD_1068_U201;
  assign ADD_1068_U53 = ~new_ADD_1068_U209 | ~new_ADD_1068_U208;
  assign ADD_1068_U54 = ~new_ADD_1068_U216 | ~new_ADD_1068_U215;
  assign ADD_1068_U55 = ~new_ADD_1068_U233 | ~new_ADD_1068_U232;
  assign ADD_1068_U56 = ~new_ADD_1068_U240 | ~new_ADD_1068_U239;
  assign ADD_1068_U57 = ~new_ADD_1068_U247 | ~new_ADD_1068_U246;
  assign ADD_1068_U58 = ~new_ADD_1068_U254 | ~new_ADD_1068_U253;
  assign ADD_1068_U59 = ~new_ADD_1068_U261 | ~new_ADD_1068_U260;
  assign ADD_1068_U60 = ~new_ADD_1068_U268 | ~new_ADD_1068_U267;
  assign ADD_1068_U61 = ~new_ADD_1068_U275 | ~new_ADD_1068_U274;
  assign ADD_1068_U62 = ~new_ADD_1068_U282 | ~new_ADD_1068_U281;
  assign ADD_1068_U63 = ~new_ADD_1068_U289 | ~new_ADD_1068_U288;
  assign new_ADD_1068_U64 = ~new_ADD_1068_U114 | ~new_ADD_1068_U113;
  assign new_ADD_1068_U65 = ~new_ADD_1068_U110 | ~new_ADD_1068_U109;
  assign new_ADD_1068_U66 = ~new_ADD_1068_U106 | ~new_ADD_1068_U105;
  assign new_ADD_1068_U67 = ~new_ADD_1068_U102 | ~new_ADD_1068_U101;
  assign new_ADD_1068_U68 = ~new_ADD_1068_U98 | ~new_ADD_1068_U97;
  assign new_ADD_1068_U69 = ~new_ADD_1068_U94 | ~new_ADD_1068_U93;
  assign new_ADD_1068_U70 = ~new_ADD_1068_U90 | ~new_ADD_1068_U89;
  assign new_ADD_1068_U71 = ~new_ADD_1068_U72 | ~new_ADD_1068_U86;
  assign new_ADD_1068_U72 = ~P1_ADDR_REG_1_ | ~new_ADD_1068_U84;
  assign new_ADD_1068_U73 = ~P2_ADDR_REG_19_;
  assign new_ADD_1068_U74 = ~P1_ADDR_REG_19_;
  assign new_ADD_1068_U75 = ~new_ADD_1068_U146 | ~new_ADD_1068_U145;
  assign new_ADD_1068_U76 = ~new_ADD_1068_U142 | ~new_ADD_1068_U141;
  assign new_ADD_1068_U77 = ~new_ADD_1068_U138 | ~new_ADD_1068_U137;
  assign new_ADD_1068_U78 = ~new_ADD_1068_U134 | ~new_ADD_1068_U133;
  assign new_ADD_1068_U79 = ~new_ADD_1068_U130 | ~new_ADD_1068_U129;
  assign new_ADD_1068_U80 = ~new_ADD_1068_U126 | ~new_ADD_1068_U125;
  assign new_ADD_1068_U81 = ~new_ADD_1068_U122 | ~new_ADD_1068_U121;
  assign new_ADD_1068_U82 = ~new_ADD_1068_U118 | ~new_ADD_1068_U117;
  assign new_ADD_1068_U83 = ~new_ADD_1068_U72;
  assign new_ADD_1068_U84 = ~new_ADD_1068_U9;
  assign new_ADD_1068_U85 = ~new_ADD_1068_U10 | ~new_ADD_1068_U9;
  assign new_ADD_1068_U86 = ~P2_ADDR_REG_1_ | ~new_ADD_1068_U85;
  assign new_ADD_1068_U87 = ~new_ADD_1068_U71;
  assign new_ADD_1068_U88 = P1_ADDR_REG_2_ | P2_ADDR_REG_2_;
  assign new_ADD_1068_U89 = ~new_ADD_1068_U88 | ~new_ADD_1068_U71;
  assign new_ADD_1068_U90 = ~P2_ADDR_REG_2_ | ~P1_ADDR_REG_2_;
  assign new_ADD_1068_U91 = ~new_ADD_1068_U70;
  assign new_ADD_1068_U92 = P1_ADDR_REG_3_ | P2_ADDR_REG_3_;
  assign new_ADD_1068_U93 = ~new_ADD_1068_U92 | ~new_ADD_1068_U70;
  assign new_ADD_1068_U94 = ~P2_ADDR_REG_3_ | ~P1_ADDR_REG_3_;
  assign new_ADD_1068_U95 = ~new_ADD_1068_U69;
  assign new_ADD_1068_U96 = P1_ADDR_REG_4_ | P2_ADDR_REG_4_;
  assign new_ADD_1068_U97 = ~new_ADD_1068_U96 | ~new_ADD_1068_U69;
  assign new_ADD_1068_U98 = ~P2_ADDR_REG_4_ | ~P1_ADDR_REG_4_;
  assign new_ADD_1068_U99 = ~new_ADD_1068_U68;
  assign new_ADD_1068_U100 = P1_ADDR_REG_5_ | P2_ADDR_REG_5_;
  assign new_ADD_1068_U101 = ~new_ADD_1068_U100 | ~new_ADD_1068_U68;
  assign new_ADD_1068_U102 = ~P2_ADDR_REG_5_ | ~P1_ADDR_REG_5_;
  assign new_ADD_1068_U103 = ~new_ADD_1068_U67;
  assign new_ADD_1068_U104 = P1_ADDR_REG_6_ | P2_ADDR_REG_6_;
  assign new_ADD_1068_U105 = ~new_ADD_1068_U104 | ~new_ADD_1068_U67;
  assign new_ADD_1068_U106 = ~P2_ADDR_REG_6_ | ~P1_ADDR_REG_6_;
  assign new_ADD_1068_U107 = ~new_ADD_1068_U66;
  assign new_ADD_1068_U108 = P1_ADDR_REG_7_ | P2_ADDR_REG_7_;
  assign new_ADD_1068_U109 = ~new_ADD_1068_U108 | ~new_ADD_1068_U66;
  assign new_ADD_1068_U110 = ~P2_ADDR_REG_7_ | ~P1_ADDR_REG_7_;
  assign new_ADD_1068_U111 = ~new_ADD_1068_U65;
  assign new_ADD_1068_U112 = P1_ADDR_REG_8_ | P2_ADDR_REG_8_;
  assign new_ADD_1068_U113 = ~new_ADD_1068_U112 | ~new_ADD_1068_U65;
  assign new_ADD_1068_U114 = ~P2_ADDR_REG_8_ | ~P1_ADDR_REG_8_;
  assign new_ADD_1068_U115 = ~new_ADD_1068_U64;
  assign new_ADD_1068_U116 = P1_ADDR_REG_9_ | P2_ADDR_REG_9_;
  assign new_ADD_1068_U117 = ~new_ADD_1068_U116 | ~new_ADD_1068_U64;
  assign new_ADD_1068_U118 = ~P1_ADDR_REG_9_ | ~P2_ADDR_REG_9_;
  assign new_ADD_1068_U119 = ~new_ADD_1068_U82;
  assign new_ADD_1068_U120 = P1_ADDR_REG_10_ | P2_ADDR_REG_10_;
  assign new_ADD_1068_U121 = ~new_ADD_1068_U120 | ~new_ADD_1068_U82;
  assign new_ADD_1068_U122 = ~P2_ADDR_REG_10_ | ~P1_ADDR_REG_10_;
  assign new_ADD_1068_U123 = ~new_ADD_1068_U81;
  assign new_ADD_1068_U124 = P1_ADDR_REG_11_ | P2_ADDR_REG_11_;
  assign new_ADD_1068_U125 = ~new_ADD_1068_U124 | ~new_ADD_1068_U81;
  assign new_ADD_1068_U126 = ~P2_ADDR_REG_11_ | ~P1_ADDR_REG_11_;
  assign new_ADD_1068_U127 = ~new_ADD_1068_U80;
  assign new_ADD_1068_U128 = P1_ADDR_REG_12_ | P2_ADDR_REG_12_;
  assign new_ADD_1068_U129 = ~new_ADD_1068_U128 | ~new_ADD_1068_U80;
  assign new_ADD_1068_U130 = ~P2_ADDR_REG_12_ | ~P1_ADDR_REG_12_;
  assign new_ADD_1068_U131 = ~new_ADD_1068_U79;
  assign new_ADD_1068_U132 = P1_ADDR_REG_13_ | P2_ADDR_REG_13_;
  assign new_ADD_1068_U133 = ~new_ADD_1068_U132 | ~new_ADD_1068_U79;
  assign new_ADD_1068_U134 = ~P2_ADDR_REG_13_ | ~P1_ADDR_REG_13_;
  assign new_ADD_1068_U135 = ~new_ADD_1068_U78;
  assign new_ADD_1068_U136 = P1_ADDR_REG_14_ | P2_ADDR_REG_14_;
  assign new_ADD_1068_U137 = ~new_ADD_1068_U136 | ~new_ADD_1068_U78;
  assign new_ADD_1068_U138 = ~P2_ADDR_REG_14_ | ~P1_ADDR_REG_14_;
  assign new_ADD_1068_U139 = ~new_ADD_1068_U77;
  assign new_ADD_1068_U140 = P1_ADDR_REG_15_ | P2_ADDR_REG_15_;
  assign new_ADD_1068_U141 = ~new_ADD_1068_U140 | ~new_ADD_1068_U77;
  assign new_ADD_1068_U142 = ~P2_ADDR_REG_15_ | ~P1_ADDR_REG_15_;
  assign new_ADD_1068_U143 = ~new_ADD_1068_U76;
  assign new_ADD_1068_U144 = P1_ADDR_REG_16_ | P2_ADDR_REG_16_;
  assign new_ADD_1068_U145 = ~new_ADD_1068_U144 | ~new_ADD_1068_U76;
  assign new_ADD_1068_U146 = ~P2_ADDR_REG_16_ | ~P1_ADDR_REG_16_;
  assign new_ADD_1068_U147 = ~new_ADD_1068_U75;
  assign new_ADD_1068_U148 = P1_ADDR_REG_17_ | P2_ADDR_REG_17_;
  assign new_ADD_1068_U149 = ~new_ADD_1068_U148 | ~new_ADD_1068_U75;
  assign new_ADD_1068_U150 = ~P2_ADDR_REG_17_ | ~P1_ADDR_REG_17_;
  assign new_ADD_1068_U151 = ~new_ADD_1068_U45;
  assign new_ADD_1068_U152 = P1_ADDR_REG_18_ | P2_ADDR_REG_18_;
  assign new_ADD_1068_U153 = ~new_ADD_1068_U152 | ~new_ADD_1068_U45;
  assign new_ADD_1068_U154 = ~P2_ADDR_REG_18_ | ~P1_ADDR_REG_18_;
  assign new_ADD_1068_U155 = ~new_ADD_1068_U153 | ~new_ADD_1068_U154 | ~new_ADD_1068_U223 | ~new_ADD_1068_U222;
  assign new_ADD_1068_U156 = ~P2_ADDR_REG_18_ | ~P1_ADDR_REG_18_;
  assign new_ADD_1068_U157 = ~new_ADD_1068_U151 | ~new_ADD_1068_U156;
  assign new_ADD_1068_U158 = P2_ADDR_REG_18_ | P1_ADDR_REG_18_;
  assign new_ADD_1068_U159 = ~new_ADD_1068_U157 | ~new_ADD_1068_U158 | ~new_ADD_1068_U226;
  assign new_ADD_1068_U160 = ~new_ADD_1068_U219 | ~new_ADD_1068_U10;
  assign new_ADD_1068_U161 = ~P2_ADDR_REG_9_ | ~new_ADD_1068_U26;
  assign new_ADD_1068_U162 = ~P1_ADDR_REG_9_ | ~new_ADD_1068_U25;
  assign new_ADD_1068_U163 = ~P2_ADDR_REG_9_ | ~new_ADD_1068_U26;
  assign new_ADD_1068_U164 = ~P1_ADDR_REG_9_ | ~new_ADD_1068_U25;
  assign new_ADD_1068_U165 = ~new_ADD_1068_U164 | ~new_ADD_1068_U163;
  assign new_ADD_1068_U166 = ~new_ADD_1068_U64 | ~new_ADD_1068_U162 | ~new_ADD_1068_U161;
  assign new_ADD_1068_U167 = ~new_ADD_1068_U115 | ~new_ADD_1068_U165;
  assign new_ADD_1068_U168 = ~P2_ADDR_REG_8_ | ~new_ADD_1068_U23;
  assign new_ADD_1068_U169 = ~P1_ADDR_REG_8_ | ~new_ADD_1068_U24;
  assign new_ADD_1068_U170 = ~P2_ADDR_REG_8_ | ~new_ADD_1068_U23;
  assign new_ADD_1068_U171 = ~P1_ADDR_REG_8_ | ~new_ADD_1068_U24;
  assign new_ADD_1068_U172 = ~new_ADD_1068_U171 | ~new_ADD_1068_U170;
  assign new_ADD_1068_U173 = ~new_ADD_1068_U65 | ~new_ADD_1068_U169 | ~new_ADD_1068_U168;
  assign new_ADD_1068_U174 = ~new_ADD_1068_U111 | ~new_ADD_1068_U172;
  assign new_ADD_1068_U175 = ~P2_ADDR_REG_7_ | ~new_ADD_1068_U21;
  assign new_ADD_1068_U176 = ~P1_ADDR_REG_7_ | ~new_ADD_1068_U22;
  assign new_ADD_1068_U177 = ~P2_ADDR_REG_7_ | ~new_ADD_1068_U21;
  assign new_ADD_1068_U178 = ~P1_ADDR_REG_7_ | ~new_ADD_1068_U22;
  assign new_ADD_1068_U179 = ~new_ADD_1068_U178 | ~new_ADD_1068_U177;
  assign new_ADD_1068_U180 = ~new_ADD_1068_U66 | ~new_ADD_1068_U176 | ~new_ADD_1068_U175;
  assign new_ADD_1068_U181 = ~new_ADD_1068_U107 | ~new_ADD_1068_U179;
  assign new_ADD_1068_U182 = ~P2_ADDR_REG_6_ | ~new_ADD_1068_U19;
  assign new_ADD_1068_U183 = ~P1_ADDR_REG_6_ | ~new_ADD_1068_U20;
  assign new_ADD_1068_U184 = ~P2_ADDR_REG_6_ | ~new_ADD_1068_U19;
  assign new_ADD_1068_U185 = ~P1_ADDR_REG_6_ | ~new_ADD_1068_U20;
  assign new_ADD_1068_U186 = ~new_ADD_1068_U185 | ~new_ADD_1068_U184;
  assign new_ADD_1068_U187 = ~new_ADD_1068_U67 | ~new_ADD_1068_U183 | ~new_ADD_1068_U182;
  assign new_ADD_1068_U188 = ~new_ADD_1068_U103 | ~new_ADD_1068_U186;
  assign new_ADD_1068_U189 = ~P2_ADDR_REG_5_ | ~new_ADD_1068_U17;
  assign new_ADD_1068_U190 = ~P1_ADDR_REG_5_ | ~new_ADD_1068_U18;
  assign new_ADD_1068_U191 = ~P2_ADDR_REG_5_ | ~new_ADD_1068_U17;
  assign new_ADD_1068_U192 = ~P1_ADDR_REG_5_ | ~new_ADD_1068_U18;
  assign new_ADD_1068_U193 = ~new_ADD_1068_U192 | ~new_ADD_1068_U191;
  assign new_ADD_1068_U194 = ~new_ADD_1068_U68 | ~new_ADD_1068_U190 | ~new_ADD_1068_U189;
  assign new_ADD_1068_U195 = ~new_ADD_1068_U99 | ~new_ADD_1068_U193;
  assign new_ADD_1068_U196 = ~P2_ADDR_REG_4_ | ~new_ADD_1068_U15;
  assign new_ADD_1068_U197 = ~P1_ADDR_REG_4_ | ~new_ADD_1068_U16;
  assign new_ADD_1068_U198 = ~P2_ADDR_REG_4_ | ~new_ADD_1068_U15;
  assign new_ADD_1068_U199 = ~P1_ADDR_REG_4_ | ~new_ADD_1068_U16;
  assign new_ADD_1068_U200 = ~new_ADD_1068_U199 | ~new_ADD_1068_U198;
  assign new_ADD_1068_U201 = ~new_ADD_1068_U69 | ~new_ADD_1068_U197 | ~new_ADD_1068_U196;
  assign new_ADD_1068_U202 = ~new_ADD_1068_U95 | ~new_ADD_1068_U200;
  assign new_ADD_1068_U203 = ~P2_ADDR_REG_3_ | ~new_ADD_1068_U13;
  assign new_ADD_1068_U204 = ~P1_ADDR_REG_3_ | ~new_ADD_1068_U14;
  assign new_ADD_1068_U205 = ~P2_ADDR_REG_3_ | ~new_ADD_1068_U13;
  assign new_ADD_1068_U206 = ~P1_ADDR_REG_3_ | ~new_ADD_1068_U14;
  assign new_ADD_1068_U207 = ~new_ADD_1068_U206 | ~new_ADD_1068_U205;
  assign new_ADD_1068_U208 = ~new_ADD_1068_U70 | ~new_ADD_1068_U204 | ~new_ADD_1068_U203;
  assign new_ADD_1068_U209 = ~new_ADD_1068_U91 | ~new_ADD_1068_U207;
  assign new_ADD_1068_U210 = ~P2_ADDR_REG_2_ | ~new_ADD_1068_U11;
  assign new_ADD_1068_U211 = ~P1_ADDR_REG_2_ | ~new_ADD_1068_U12;
  assign new_ADD_1068_U212 = ~P2_ADDR_REG_2_ | ~new_ADD_1068_U11;
  assign new_ADD_1068_U213 = ~P1_ADDR_REG_2_ | ~new_ADD_1068_U12;
  assign new_ADD_1068_U214 = ~new_ADD_1068_U213 | ~new_ADD_1068_U212;
  assign new_ADD_1068_U215 = ~new_ADD_1068_U71 | ~new_ADD_1068_U211 | ~new_ADD_1068_U210;
  assign new_ADD_1068_U216 = ~new_ADD_1068_U87 | ~new_ADD_1068_U214;
  assign new_ADD_1068_U217 = ~P2_ADDR_REG_1_ | ~new_ADD_1068_U9;
  assign new_ADD_1068_U218 = ~new_ADD_1068_U84 | ~new_ADD_1068_U8;
  assign new_ADD_1068_U219 = ~new_ADD_1068_U218 | ~new_ADD_1068_U217;
  assign new_ADD_1068_U220 = ~new_ADD_1068_U8 | ~P1_ADDR_REG_1_ | ~new_ADD_1068_U9;
  assign new_ADD_1068_U221 = ~new_ADD_1068_U83 | ~P2_ADDR_REG_1_;
  assign new_ADD_1068_U222 = ~P2_ADDR_REG_19_ | ~new_ADD_1068_U74;
  assign new_ADD_1068_U223 = ~P1_ADDR_REG_19_ | ~new_ADD_1068_U73;
  assign new_ADD_1068_U224 = ~P2_ADDR_REG_19_ | ~new_ADD_1068_U74;
  assign new_ADD_1068_U225 = ~P1_ADDR_REG_19_ | ~new_ADD_1068_U73;
  assign new_ADD_1068_U226 = ~new_ADD_1068_U225 | ~new_ADD_1068_U224;
  assign new_ADD_1068_U227 = ~P2_ADDR_REG_18_ | ~new_ADD_1068_U43;
  assign new_ADD_1068_U228 = ~P1_ADDR_REG_18_ | ~new_ADD_1068_U44;
  assign new_ADD_1068_U229 = ~P2_ADDR_REG_18_ | ~new_ADD_1068_U43;
  assign new_ADD_1068_U230 = ~P1_ADDR_REG_18_ | ~new_ADD_1068_U44;
  assign new_ADD_1068_U231 = ~new_ADD_1068_U230 | ~new_ADD_1068_U229;
  assign new_ADD_1068_U232 = ~new_ADD_1068_U45 | ~new_ADD_1068_U228 | ~new_ADD_1068_U227;
  assign new_ADD_1068_U233 = ~new_ADD_1068_U231 | ~new_ADD_1068_U151;
  assign new_ADD_1068_U234 = ~P2_ADDR_REG_17_ | ~new_ADD_1068_U41;
  assign new_ADD_1068_U235 = ~P1_ADDR_REG_17_ | ~new_ADD_1068_U42;
  assign new_ADD_1068_U236 = ~P2_ADDR_REG_17_ | ~new_ADD_1068_U41;
  assign new_ADD_1068_U237 = ~P1_ADDR_REG_17_ | ~new_ADD_1068_U42;
  assign new_ADD_1068_U238 = ~new_ADD_1068_U237 | ~new_ADD_1068_U236;
  assign new_ADD_1068_U239 = ~new_ADD_1068_U75 | ~new_ADD_1068_U235 | ~new_ADD_1068_U234;
  assign new_ADD_1068_U240 = ~new_ADD_1068_U147 | ~new_ADD_1068_U238;
  assign new_ADD_1068_U241 = ~P2_ADDR_REG_16_ | ~new_ADD_1068_U39;
  assign new_ADD_1068_U242 = ~P1_ADDR_REG_16_ | ~new_ADD_1068_U40;
  assign new_ADD_1068_U243 = ~P2_ADDR_REG_16_ | ~new_ADD_1068_U39;
  assign new_ADD_1068_U244 = ~P1_ADDR_REG_16_ | ~new_ADD_1068_U40;
  assign new_ADD_1068_U245 = ~new_ADD_1068_U244 | ~new_ADD_1068_U243;
  assign new_ADD_1068_U246 = ~new_ADD_1068_U76 | ~new_ADD_1068_U242 | ~new_ADD_1068_U241;
  assign new_ADD_1068_U247 = ~new_ADD_1068_U143 | ~new_ADD_1068_U245;
  assign new_ADD_1068_U248 = ~P2_ADDR_REG_15_ | ~new_ADD_1068_U37;
  assign new_ADD_1068_U249 = ~P1_ADDR_REG_15_ | ~new_ADD_1068_U38;
  assign new_ADD_1068_U250 = ~P2_ADDR_REG_15_ | ~new_ADD_1068_U37;
  assign new_ADD_1068_U251 = ~P1_ADDR_REG_15_ | ~new_ADD_1068_U38;
  assign new_ADD_1068_U252 = ~new_ADD_1068_U251 | ~new_ADD_1068_U250;
  assign new_ADD_1068_U253 = ~new_ADD_1068_U77 | ~new_ADD_1068_U249 | ~new_ADD_1068_U248;
  assign new_ADD_1068_U254 = ~new_ADD_1068_U139 | ~new_ADD_1068_U252;
  assign new_ADD_1068_U255 = ~P2_ADDR_REG_14_ | ~new_ADD_1068_U35;
  assign new_ADD_1068_U256 = ~P1_ADDR_REG_14_ | ~new_ADD_1068_U36;
  assign new_ADD_1068_U257 = ~P2_ADDR_REG_14_ | ~new_ADD_1068_U35;
  assign new_ADD_1068_U258 = ~P1_ADDR_REG_14_ | ~new_ADD_1068_U36;
  assign new_ADD_1068_U259 = ~new_ADD_1068_U258 | ~new_ADD_1068_U257;
  assign new_ADD_1068_U260 = ~new_ADD_1068_U78 | ~new_ADD_1068_U256 | ~new_ADD_1068_U255;
  assign new_ADD_1068_U261 = ~new_ADD_1068_U135 | ~new_ADD_1068_U259;
  assign new_ADD_1068_U262 = ~P2_ADDR_REG_13_ | ~new_ADD_1068_U33;
  assign new_ADD_1068_U263 = ~P1_ADDR_REG_13_ | ~new_ADD_1068_U34;
  assign new_ADD_1068_U264 = ~P2_ADDR_REG_13_ | ~new_ADD_1068_U33;
  assign new_ADD_1068_U265 = ~P1_ADDR_REG_13_ | ~new_ADD_1068_U34;
  assign new_ADD_1068_U266 = ~new_ADD_1068_U265 | ~new_ADD_1068_U264;
  assign new_ADD_1068_U267 = ~new_ADD_1068_U79 | ~new_ADD_1068_U263 | ~new_ADD_1068_U262;
  assign new_ADD_1068_U268 = ~new_ADD_1068_U131 | ~new_ADD_1068_U266;
  assign new_ADD_1068_U269 = ~P2_ADDR_REG_12_ | ~new_ADD_1068_U31;
  assign new_ADD_1068_U270 = ~P1_ADDR_REG_12_ | ~new_ADD_1068_U32;
  assign new_ADD_1068_U271 = ~P2_ADDR_REG_12_ | ~new_ADD_1068_U31;
  assign new_ADD_1068_U272 = ~P1_ADDR_REG_12_ | ~new_ADD_1068_U32;
  assign new_ADD_1068_U273 = ~new_ADD_1068_U272 | ~new_ADD_1068_U271;
  assign new_ADD_1068_U274 = ~new_ADD_1068_U80 | ~new_ADD_1068_U270 | ~new_ADD_1068_U269;
  assign new_ADD_1068_U275 = ~new_ADD_1068_U127 | ~new_ADD_1068_U273;
  assign new_ADD_1068_U276 = ~P2_ADDR_REG_11_ | ~new_ADD_1068_U29;
  assign new_ADD_1068_U277 = ~P1_ADDR_REG_11_ | ~new_ADD_1068_U30;
  assign new_ADD_1068_U278 = ~P2_ADDR_REG_11_ | ~new_ADD_1068_U29;
  assign new_ADD_1068_U279 = ~P1_ADDR_REG_11_ | ~new_ADD_1068_U30;
  assign new_ADD_1068_U280 = ~new_ADD_1068_U279 | ~new_ADD_1068_U278;
  assign new_ADD_1068_U281 = ~new_ADD_1068_U81 | ~new_ADD_1068_U277 | ~new_ADD_1068_U276;
  assign new_ADD_1068_U282 = ~new_ADD_1068_U123 | ~new_ADD_1068_U280;
  assign new_ADD_1068_U283 = ~P2_ADDR_REG_10_ | ~new_ADD_1068_U27;
  assign new_ADD_1068_U284 = ~P1_ADDR_REG_10_ | ~new_ADD_1068_U28;
  assign new_ADD_1068_U285 = ~P2_ADDR_REG_10_ | ~new_ADD_1068_U27;
  assign new_ADD_1068_U286 = ~P1_ADDR_REG_10_ | ~new_ADD_1068_U28;
  assign new_ADD_1068_U287 = ~new_ADD_1068_U286 | ~new_ADD_1068_U285;
  assign new_ADD_1068_U288 = ~new_ADD_1068_U82 | ~new_ADD_1068_U284 | ~new_ADD_1068_U283;
  assign new_ADD_1068_U289 = ~new_ADD_1068_U119 | ~new_ADD_1068_U287;
  assign new_ADD_1068_U290 = ~P2_ADDR_REG_0_ | ~new_ADD_1068_U6;
  assign new_ADD_1068_U291 = ~P1_ADDR_REG_0_ | ~new_ADD_1068_U7;
  assign new_R140_U4 = new_R140_U197 & new_R140_U195;
  assign new_R140_U5 = new_R140_U203 & new_R140_U201;
  assign new_R140_U6 = new_R140_U5 & new_R140_U205;
  assign new_R140_U7 = new_R140_U213 & new_R140_U209;
  assign new_R140_U8 = new_R140_U7 & new_R140_U216;
  assign new_R140_U9 = new_R140_U378 & new_R140_U377;
  assign new_R140_U10 = ~new_R140_U324 | ~new_R140_U469 | ~new_R140_U468;
  assign new_R140_U11 = new_R140_U124 & new_R140_U323;
  assign new_R140_U12 = ~SI_8_;
  assign new_R140_U13 = ~new_U90;
  assign new_R140_U14 = ~SI_7_;
  assign new_R140_U15 = ~new_U91;
  assign new_R140_U16 = ~new_U91 | ~SI_7_;
  assign new_R140_U17 = ~SI_6_;
  assign new_R140_U18 = ~new_U92;
  assign new_R140_U19 = ~SI_5_;
  assign new_R140_U20 = ~new_U93;
  assign new_R140_U21 = ~SI_4_;
  assign new_R140_U22 = ~new_U94;
  assign new_R140_U23 = ~new_U94 | ~SI_4_;
  assign new_R140_U24 = ~SI_3_;
  assign new_R140_U25 = ~new_U97;
  assign new_R140_U26 = ~SI_2_;
  assign new_R140_U27 = ~new_U108;
  assign new_R140_U28 = ~new_U108 | ~SI_2_;
  assign new_R140_U29 = ~SI_1_;
  assign new_R140_U30 = ~SI_0_;
  assign new_R140_U31 = ~new_U120;
  assign new_R140_U32 = ~new_U119;
  assign new_R140_U33 = ~new_U89;
  assign new_R140_U34 = ~SI_9_;
  assign new_R140_U35 = ~new_R140_U288 | ~new_R140_U198;
  assign new_R140_U36 = ~SI_14_;
  assign new_R140_U37 = ~new_U114;
  assign new_R140_U38 = ~SI_10_;
  assign new_R140_U39 = ~new_U118;
  assign new_R140_U40 = ~SI_13_;
  assign new_R140_U41 = ~new_U115;
  assign new_R140_U42 = ~SI_12_;
  assign new_R140_U43 = ~new_U116;
  assign new_R140_U44 = ~SI_11_;
  assign new_R140_U45 = ~new_U117;
  assign new_R140_U46 = ~new_U117 | ~SI_11_;
  assign new_R140_U47 = ~SI_15_;
  assign new_R140_U48 = ~new_U113;
  assign new_R140_U49 = ~SI_16_;
  assign new_R140_U50 = ~new_U112;
  assign new_R140_U51 = ~SI_17_;
  assign new_R140_U52 = ~new_U111;
  assign new_R140_U53 = ~SI_18_;
  assign new_R140_U54 = ~new_U110;
  assign new_R140_U55 = ~SI_19_;
  assign new_R140_U56 = ~new_U109;
  assign new_R140_U57 = ~SI_20_;
  assign new_R140_U58 = ~new_U107;
  assign new_R140_U59 = ~SI_21_;
  assign new_R140_U60 = ~new_U106;
  assign new_R140_U61 = ~SI_22_;
  assign new_R140_U62 = ~new_U105;
  assign new_R140_U63 = ~SI_23_;
  assign new_R140_U64 = ~new_U104;
  assign new_R140_U65 = ~SI_24_;
  assign new_R140_U66 = ~new_U103;
  assign new_R140_U67 = ~SI_25_;
  assign new_R140_U68 = ~new_U102;
  assign new_R140_U69 = ~SI_26_;
  assign new_R140_U70 = ~new_U101;
  assign new_R140_U71 = ~SI_27_;
  assign new_R140_U72 = ~new_U100;
  assign new_R140_U73 = ~SI_28_;
  assign new_R140_U74 = ~new_U99;
  assign new_R140_U75 = ~SI_29_;
  assign new_R140_U76 = ~new_U98;
  assign new_R140_U77 = ~SI_30_;
  assign new_R140_U78 = ~new_U96;
  assign new_R140_U79 = ~new_U120 | ~SI_0_ | ~SI_1_;
  assign new_R140_U80 = ~new_R140_U300 | ~new_R140_U217;
  assign new_R140_U81 = ~new_R140_U297 | ~new_R140_U214;
  assign new_R140_U82 = ~new_R140_U293 | ~new_R140_U206;
  assign new_R140_U83 = ~new_R140_U541 | ~new_R140_U540;
  assign new_R140_U84 = ~new_R140_U331 | ~new_R140_U330;
  assign new_R140_U85 = ~new_R140_U338 | ~new_R140_U337;
  assign new_R140_U86 = ~new_R140_U345 | ~new_R140_U344;
  assign new_R140_U87 = ~new_R140_U352 | ~new_R140_U351;
  assign new_R140_U88 = ~new_R140_U359 | ~new_R140_U358;
  assign new_R140_U89 = ~new_R140_U366 | ~new_R140_U365;
  assign new_R140_U90 = ~new_R140_U373 | ~new_R140_U372;
  assign new_R140_U91 = ~new_R140_U387 | ~new_R140_U386;
  assign new_R140_U92 = ~new_R140_U394 | ~new_R140_U393;
  assign new_R140_U93 = ~new_R140_U401 | ~new_R140_U400;
  assign new_R140_U94 = ~new_R140_U408 | ~new_R140_U407;
  assign new_R140_U95 = ~new_R140_U415 | ~new_R140_U414;
  assign new_R140_U96 = ~new_R140_U422 | ~new_R140_U421;
  assign new_R140_U97 = ~new_R140_U429 | ~new_R140_U428;
  assign new_R140_U98 = ~new_R140_U436 | ~new_R140_U435;
  assign new_R140_U99 = ~new_R140_U443 | ~new_R140_U442;
  assign new_R140_U100 = ~new_R140_U450 | ~new_R140_U449;
  assign new_R140_U101 = ~new_R140_U457 | ~new_R140_U456;
  assign new_R140_U102 = ~new_R140_U464 | ~new_R140_U463;
  assign new_R140_U103 = ~new_R140_U476 | ~new_R140_U475;
  assign new_R140_U104 = ~new_R140_U483 | ~new_R140_U482;
  assign new_R140_U105 = ~new_R140_U490 | ~new_R140_U489;
  assign new_R140_U106 = ~new_R140_U497 | ~new_R140_U496;
  assign new_R140_U107 = ~new_R140_U504 | ~new_R140_U503;
  assign new_R140_U108 = ~new_R140_U511 | ~new_R140_U510;
  assign new_R140_U109 = ~new_R140_U518 | ~new_R140_U517;
  assign new_R140_U110 = ~new_R140_U525 | ~new_R140_U524;
  assign new_R140_U111 = ~new_R140_U532 | ~new_R140_U531;
  assign new_R140_U112 = ~new_R140_U539 | ~new_R140_U538;
  assign new_R140_U113 = new_R140_U189 & new_R140_U193;
  assign new_R140_U114 = new_R140_U287 & new_R140_U194;
  assign new_R140_U115 = new_R140_U4 & new_R140_U199;
  assign new_R140_U116 = new_R140_U290 & new_R140_U200;
  assign new_R140_U117 = new_R140_U291 & new_R140_U204;
  assign new_R140_U118 = new_R140_U6 & new_R140_U207;
  assign new_R140_U119 = new_R140_U295 & new_R140_U208;
  assign new_R140_U120 = new_R140_U8 & new_R140_U219;
  assign new_R140_U121 = new_R140_U303 & new_R140_U220;
  assign new_R140_U122 = new_R140_U280 & new_R140_U9 & new_R140_U282;
  assign new_R140_U123 = new_R140_U283 & new_R140_U376;
  assign new_R140_U124 = new_R140_U141 & new_R140_U284;
  assign new_R140_U125 = new_R140_U326 & new_R140_U325;
  assign new_R140_U126 = ~new_R140_U117 | ~new_R140_U309;
  assign new_R140_U127 = new_R140_U333 & new_R140_U332;
  assign new_R140_U128 = ~new_R140_U307 | ~new_R140_U16;
  assign new_R140_U129 = new_R140_U340 & new_R140_U339;
  assign new_R140_U130 = ~new_R140_U116 | ~new_R140_U319;
  assign new_R140_U131 = new_R140_U347 & new_R140_U346;
  assign new_R140_U132 = ~new_R140_U289 | ~new_R140_U317;
  assign new_R140_U133 = new_R140_U354 & new_R140_U353;
  assign new_R140_U134 = ~new_R140_U315 | ~new_R140_U23;
  assign new_R140_U135 = new_R140_U361 & new_R140_U360;
  assign new_R140_U136 = ~new_R140_U114 | ~new_R140_U321;
  assign new_R140_U137 = new_R140_U368 & new_R140_U367;
  assign new_R140_U138 = ~new_R140_U28 | ~new_R140_U190;
  assign new_R140_U139 = ~new_U95;
  assign new_R140_U140 = ~SI_31_;
  assign new_R140_U141 = new_R140_U380 & new_R140_U379;
  assign new_R140_U142 = new_R140_U382 & new_R140_U381;
  assign new_R140_U143 = ~new_R140_U280 | ~new_R140_U279;
  assign new_R140_U144 = ~new_R140_U285 | ~new_R140_U286 | ~new_R140_U79;
  assign new_R140_U145 = new_R140_U396 & new_R140_U395;
  assign new_R140_U146 = ~new_R140_U276 | ~new_R140_U275;
  assign new_R140_U147 = new_R140_U403 & new_R140_U402;
  assign new_R140_U148 = ~new_R140_U272 | ~new_R140_U271;
  assign new_R140_U149 = new_R140_U410 & new_R140_U409;
  assign new_R140_U150 = ~new_R140_U268 | ~new_R140_U267;
  assign new_R140_U151 = new_R140_U417 & new_R140_U416;
  assign new_R140_U152 = ~new_R140_U264 | ~new_R140_U263;
  assign new_R140_U153 = new_R140_U424 & new_R140_U423;
  assign new_R140_U154 = ~new_R140_U260 | ~new_R140_U259;
  assign new_R140_U155 = new_R140_U431 & new_R140_U430;
  assign new_R140_U156 = ~new_R140_U256 | ~new_R140_U255;
  assign new_R140_U157 = new_R140_U438 & new_R140_U437;
  assign new_R140_U158 = ~new_R140_U252 | ~new_R140_U251;
  assign new_R140_U159 = new_R140_U445 & new_R140_U444;
  assign new_R140_U160 = ~new_R140_U248 | ~new_R140_U247;
  assign new_R140_U161 = new_R140_U452 & new_R140_U451;
  assign new_R140_U162 = ~new_R140_U244 | ~new_R140_U243;
  assign new_R140_U163 = new_R140_U459 & new_R140_U458;
  assign new_R140_U164 = ~new_R140_U240 | ~new_R140_U239;
  assign new_R140_U165 = ~new_U120 | ~SI_0_;
  assign new_R140_U166 = new_R140_U471 & new_R140_U470;
  assign new_R140_U167 = ~new_R140_U236 | ~new_R140_U235;
  assign new_R140_U168 = new_R140_U478 & new_R140_U477;
  assign new_R140_U169 = ~new_R140_U232 | ~new_R140_U231;
  assign new_R140_U170 = new_R140_U485 & new_R140_U484;
  assign new_R140_U171 = ~new_R140_U228 | ~new_R140_U227;
  assign new_R140_U172 = new_R140_U492 & new_R140_U491;
  assign new_R140_U173 = ~new_R140_U224 | ~new_R140_U223;
  assign new_R140_U174 = new_R140_U499 & new_R140_U498;
  assign new_R140_U175 = ~new_R140_U121 | ~new_R140_U302;
  assign new_R140_U176 = new_R140_U506 & new_R140_U505;
  assign new_R140_U177 = ~new_R140_U301 | ~new_R140_U299;
  assign new_R140_U178 = new_R140_U513 & new_R140_U512;
  assign new_R140_U179 = ~new_R140_U298 | ~new_R140_U296;
  assign new_R140_U180 = new_R140_U520 & new_R140_U519;
  assign new_R140_U181 = ~new_R140_U46 | ~new_R140_U210;
  assign new_R140_U182 = new_R140_U527 & new_R140_U526;
  assign new_R140_U183 = ~new_R140_U119 | ~new_R140_U313;
  assign new_R140_U184 = new_R140_U534 & new_R140_U533;
  assign new_R140_U185 = ~new_R140_U294 | ~new_R140_U311;
  assign new_R140_U186 = ~new_R140_U79;
  assign new_R140_U187 = ~new_R140_U165;
  assign new_R140_U188 = ~new_R140_U144;
  assign new_R140_U189 = SI_2_ | new_U108;
  assign new_R140_U190 = ~new_R140_U304 | ~new_R140_U189;
  assign new_R140_U191 = ~new_R140_U28;
  assign new_R140_U192 = ~new_R140_U138;
  assign new_R140_U193 = SI_3_ | new_U97;
  assign new_R140_U194 = ~new_U97 | ~SI_3_;
  assign new_R140_U195 = SI_4_ | new_U94;
  assign new_R140_U196 = ~new_R140_U23;
  assign new_R140_U197 = SI_5_ | new_U93;
  assign new_R140_U198 = ~new_U93 | ~SI_5_;
  assign new_R140_U199 = SI_6_ | new_U92;
  assign new_R140_U200 = ~new_U92 | ~SI_6_;
  assign new_R140_U201 = SI_7_ | new_U91;
  assign new_R140_U202 = ~new_R140_U16;
  assign new_R140_U203 = SI_8_ | new_U90;
  assign new_R140_U204 = ~new_U90 | ~SI_8_;
  assign new_R140_U205 = SI_9_ | new_U89;
  assign new_R140_U206 = ~SI_9_ | ~new_U89;
  assign new_R140_U207 = SI_10_ | new_U118;
  assign new_R140_U208 = ~new_U118 | ~SI_10_;
  assign new_R140_U209 = SI_11_ | new_U117;
  assign new_R140_U210 = ~new_R140_U209 | ~new_R140_U183;
  assign new_R140_U211 = ~new_R140_U46;
  assign new_R140_U212 = ~new_R140_U181;
  assign new_R140_U213 = SI_12_ | new_U116;
  assign new_R140_U214 = ~new_U116 | ~SI_12_;
  assign new_R140_U215 = ~new_R140_U179;
  assign new_R140_U216 = SI_13_ | new_U115;
  assign new_R140_U217 = ~new_U115 | ~SI_13_;
  assign new_R140_U218 = ~new_R140_U177;
  assign new_R140_U219 = SI_14_ | new_U114;
  assign new_R140_U220 = ~new_U114 | ~SI_14_;
  assign new_R140_U221 = ~new_R140_U175;
  assign new_R140_U222 = SI_15_ | new_U113;
  assign new_R140_U223 = ~new_R140_U222 | ~new_R140_U175;
  assign new_R140_U224 = ~new_U113 | ~SI_15_;
  assign new_R140_U225 = ~new_R140_U173;
  assign new_R140_U226 = SI_16_ | new_U112;
  assign new_R140_U227 = ~new_R140_U226 | ~new_R140_U173;
  assign new_R140_U228 = ~new_U112 | ~SI_16_;
  assign new_R140_U229 = ~new_R140_U171;
  assign new_R140_U230 = SI_17_ | new_U111;
  assign new_R140_U231 = ~new_R140_U230 | ~new_R140_U171;
  assign new_R140_U232 = ~new_U111 | ~SI_17_;
  assign new_R140_U233 = ~new_R140_U169;
  assign new_R140_U234 = SI_18_ | new_U110;
  assign new_R140_U235 = ~new_R140_U234 | ~new_R140_U169;
  assign new_R140_U236 = ~new_U110 | ~SI_18_;
  assign new_R140_U237 = ~new_R140_U167;
  assign new_R140_U238 = SI_19_ | new_U109;
  assign new_R140_U239 = ~new_R140_U238 | ~new_R140_U167;
  assign new_R140_U240 = ~new_U109 | ~SI_19_;
  assign new_R140_U241 = ~new_R140_U164;
  assign new_R140_U242 = SI_20_ | new_U107;
  assign new_R140_U243 = ~new_R140_U242 | ~new_R140_U164;
  assign new_R140_U244 = ~new_U107 | ~SI_20_;
  assign new_R140_U245 = ~new_R140_U162;
  assign new_R140_U246 = SI_21_ | new_U106;
  assign new_R140_U247 = ~new_R140_U246 | ~new_R140_U162;
  assign new_R140_U248 = ~new_U106 | ~SI_21_;
  assign new_R140_U249 = ~new_R140_U160;
  assign new_R140_U250 = SI_22_ | new_U105;
  assign new_R140_U251 = ~new_R140_U250 | ~new_R140_U160;
  assign new_R140_U252 = ~new_U105 | ~SI_22_;
  assign new_R140_U253 = ~new_R140_U158;
  assign new_R140_U254 = SI_23_ | new_U104;
  assign new_R140_U255 = ~new_R140_U254 | ~new_R140_U158;
  assign new_R140_U256 = ~new_U104 | ~SI_23_;
  assign new_R140_U257 = ~new_R140_U156;
  assign new_R140_U258 = SI_24_ | new_U103;
  assign new_R140_U259 = ~new_R140_U258 | ~new_R140_U156;
  assign new_R140_U260 = ~new_U103 | ~SI_24_;
  assign new_R140_U261 = ~new_R140_U154;
  assign new_R140_U262 = SI_25_ | new_U102;
  assign new_R140_U263 = ~new_R140_U262 | ~new_R140_U154;
  assign new_R140_U264 = ~new_U102 | ~SI_25_;
  assign new_R140_U265 = ~new_R140_U152;
  assign new_R140_U266 = SI_26_ | new_U101;
  assign new_R140_U267 = ~new_R140_U266 | ~new_R140_U152;
  assign new_R140_U268 = ~new_U101 | ~SI_26_;
  assign new_R140_U269 = ~new_R140_U150;
  assign new_R140_U270 = SI_27_ | new_U100;
  assign new_R140_U271 = ~new_R140_U270 | ~new_R140_U150;
  assign new_R140_U272 = ~new_U100 | ~SI_27_;
  assign new_R140_U273 = ~new_R140_U148;
  assign new_R140_U274 = SI_28_ | new_U99;
  assign new_R140_U275 = ~new_R140_U274 | ~new_R140_U148;
  assign new_R140_U276 = ~new_U99 | ~SI_28_;
  assign new_R140_U277 = ~new_R140_U146;
  assign new_R140_U278 = SI_29_ | new_U98;
  assign new_R140_U279 = ~new_R140_U278 | ~new_R140_U146;
  assign new_R140_U280 = ~new_U98 | ~SI_29_;
  assign new_R140_U281 = ~new_R140_U143;
  assign new_R140_U282 = ~new_U96 | ~SI_30_;
  assign new_R140_U283 = new_U96 | SI_30_;
  assign new_R140_U284 = ~new_R140_U279 | ~new_R140_U122;
  assign new_R140_U285 = ~new_U119 | ~new_U120 | ~SI_0_;
  assign new_R140_U286 = ~new_U119 | ~SI_1_;
  assign new_R140_U287 = ~new_R140_U191 | ~new_R140_U193;
  assign new_R140_U288 = ~new_R140_U196 | ~new_R140_U197;
  assign new_R140_U289 = ~new_R140_U35;
  assign new_R140_U290 = ~new_R140_U35 | ~new_R140_U199;
  assign new_R140_U291 = ~new_R140_U202 | ~new_R140_U203;
  assign new_R140_U292 = ~new_R140_U291 | ~new_R140_U204;
  assign new_R140_U293 = ~new_R140_U292 | ~new_R140_U205;
  assign new_R140_U294 = ~new_R140_U82;
  assign new_R140_U295 = ~new_R140_U82 | ~new_R140_U207;
  assign new_R140_U296 = ~new_R140_U7 | ~new_R140_U183;
  assign new_R140_U297 = ~new_R140_U211 | ~new_R140_U213;
  assign new_R140_U298 = ~new_R140_U81;
  assign new_R140_U299 = ~new_R140_U8 | ~new_R140_U183;
  assign new_R140_U300 = ~new_R140_U81 | ~new_R140_U216;
  assign new_R140_U301 = ~new_R140_U80;
  assign new_R140_U302 = ~new_R140_U120 | ~new_R140_U183;
  assign new_R140_U303 = ~new_R140_U80 | ~new_R140_U219;
  assign new_R140_U304 = ~new_R140_U305 | ~new_R140_U306 | ~new_R140_U286;
  assign new_R140_U305 = ~new_U119 | ~new_U120 | ~SI_0_;
  assign new_R140_U306 = ~new_U120 | ~SI_0_ | ~SI_1_;
  assign new_R140_U307 = ~new_R140_U201 | ~new_R140_U130;
  assign new_R140_U308 = ~new_R140_U128;
  assign new_R140_U309 = ~new_R140_U5 | ~new_R140_U130;
  assign new_R140_U310 = ~new_R140_U126;
  assign new_R140_U311 = ~new_R140_U6 | ~new_R140_U130;
  assign new_R140_U312 = ~new_R140_U185;
  assign new_R140_U313 = ~new_R140_U118 | ~new_R140_U130;
  assign new_R140_U314 = ~new_R140_U183;
  assign new_R140_U315 = ~new_R140_U195 | ~new_R140_U136;
  assign new_R140_U316 = ~new_R140_U134;
  assign new_R140_U317 = ~new_R140_U4 | ~new_R140_U136;
  assign new_R140_U318 = ~new_R140_U132;
  assign new_R140_U319 = ~new_R140_U115 | ~new_R140_U136;
  assign new_R140_U320 = ~new_R140_U130;
  assign new_R140_U321 = ~new_R140_U113 | ~new_R140_U144;
  assign new_R140_U322 = ~new_R140_U136;
  assign new_R140_U323 = ~new_R140_U123 | ~new_R140_U143;
  assign new_R140_U324 = ~new_R140_U186 | ~new_U119;
  assign new_R140_U325 = ~new_U89 | ~new_R140_U34;
  assign new_R140_U326 = ~SI_9_ | ~new_R140_U33;
  assign new_R140_U327 = ~new_U89 | ~new_R140_U34;
  assign new_R140_U328 = ~SI_9_ | ~new_R140_U33;
  assign new_R140_U329 = ~new_R140_U328 | ~new_R140_U327;
  assign new_R140_U330 = ~new_R140_U125 | ~new_R140_U126;
  assign new_R140_U331 = ~new_R140_U310 | ~new_R140_U329;
  assign new_R140_U332 = ~new_U90 | ~new_R140_U12;
  assign new_R140_U333 = ~SI_8_ | ~new_R140_U13;
  assign new_R140_U334 = ~new_U90 | ~new_R140_U12;
  assign new_R140_U335 = ~SI_8_ | ~new_R140_U13;
  assign new_R140_U336 = ~new_R140_U335 | ~new_R140_U334;
  assign new_R140_U337 = ~new_R140_U127 | ~new_R140_U128;
  assign new_R140_U338 = ~new_R140_U308 | ~new_R140_U336;
  assign new_R140_U339 = ~new_U91 | ~new_R140_U14;
  assign new_R140_U340 = ~SI_7_ | ~new_R140_U15;
  assign new_R140_U341 = ~new_U91 | ~new_R140_U14;
  assign new_R140_U342 = ~SI_7_ | ~new_R140_U15;
  assign new_R140_U343 = ~new_R140_U342 | ~new_R140_U341;
  assign new_R140_U344 = ~new_R140_U129 | ~new_R140_U130;
  assign new_R140_U345 = ~new_R140_U320 | ~new_R140_U343;
  assign new_R140_U346 = ~new_U92 | ~new_R140_U17;
  assign new_R140_U347 = ~SI_6_ | ~new_R140_U18;
  assign new_R140_U348 = ~new_U92 | ~new_R140_U17;
  assign new_R140_U349 = ~SI_6_ | ~new_R140_U18;
  assign new_R140_U350 = ~new_R140_U349 | ~new_R140_U348;
  assign new_R140_U351 = ~new_R140_U131 | ~new_R140_U132;
  assign new_R140_U352 = ~new_R140_U318 | ~new_R140_U350;
  assign new_R140_U353 = ~new_U93 | ~new_R140_U19;
  assign new_R140_U354 = ~SI_5_ | ~new_R140_U20;
  assign new_R140_U355 = ~new_U93 | ~new_R140_U19;
  assign new_R140_U356 = ~SI_5_ | ~new_R140_U20;
  assign new_R140_U357 = ~new_R140_U356 | ~new_R140_U355;
  assign new_R140_U358 = ~new_R140_U133 | ~new_R140_U134;
  assign new_R140_U359 = ~new_R140_U316 | ~new_R140_U357;
  assign new_R140_U360 = ~new_U94 | ~new_R140_U21;
  assign new_R140_U361 = ~SI_4_ | ~new_R140_U22;
  assign new_R140_U362 = ~new_U94 | ~new_R140_U21;
  assign new_R140_U363 = ~SI_4_ | ~new_R140_U22;
  assign new_R140_U364 = ~new_R140_U363 | ~new_R140_U362;
  assign new_R140_U365 = ~new_R140_U135 | ~new_R140_U136;
  assign new_R140_U366 = ~new_R140_U322 | ~new_R140_U364;
  assign new_R140_U367 = ~new_U97 | ~new_R140_U24;
  assign new_R140_U368 = ~SI_3_ | ~new_R140_U25;
  assign new_R140_U369 = ~new_U97 | ~new_R140_U24;
  assign new_R140_U370 = ~SI_3_ | ~new_R140_U25;
  assign new_R140_U371 = ~new_R140_U370 | ~new_R140_U369;
  assign new_R140_U372 = ~new_R140_U137 | ~new_R140_U138;
  assign new_R140_U373 = ~new_R140_U192 | ~new_R140_U371;
  assign new_R140_U374 = ~new_U95 | ~new_R140_U140;
  assign new_R140_U375 = ~SI_31_ | ~new_R140_U139;
  assign new_R140_U376 = ~new_R140_U375 | ~new_R140_U374;
  assign new_R140_U377 = ~new_U95 | ~new_R140_U140;
  assign new_R140_U378 = ~SI_31_ | ~new_R140_U139;
  assign new_R140_U379 = ~new_R140_U78 | ~new_R140_U9 | ~new_R140_U77;
  assign new_R140_U380 = ~new_U96 | ~SI_30_ | ~new_R140_U376;
  assign new_R140_U381 = ~new_U96 | ~new_R140_U77;
  assign new_R140_U382 = ~SI_30_ | ~new_R140_U78;
  assign new_R140_U383 = ~new_U96 | ~new_R140_U77;
  assign new_R140_U384 = ~SI_30_ | ~new_R140_U78;
  assign new_R140_U385 = ~new_R140_U384 | ~new_R140_U383;
  assign new_R140_U386 = ~new_R140_U142 | ~new_R140_U143;
  assign new_R140_U387 = ~new_R140_U281 | ~new_R140_U385;
  assign new_R140_U388 = ~new_U108 | ~new_R140_U26;
  assign new_R140_U389 = ~SI_2_ | ~new_R140_U27;
  assign new_R140_U390 = ~new_U108 | ~new_R140_U26;
  assign new_R140_U391 = ~SI_2_ | ~new_R140_U27;
  assign new_R140_U392 = ~new_R140_U391 | ~new_R140_U390;
  assign new_R140_U393 = ~new_R140_U144 | ~new_R140_U389 | ~new_R140_U388;
  assign new_R140_U394 = ~new_R140_U188 | ~new_R140_U392;
  assign new_R140_U395 = ~new_U98 | ~new_R140_U75;
  assign new_R140_U396 = ~SI_29_ | ~new_R140_U76;
  assign new_R140_U397 = ~new_U98 | ~new_R140_U75;
  assign new_R140_U398 = ~SI_29_ | ~new_R140_U76;
  assign new_R140_U399 = ~new_R140_U398 | ~new_R140_U397;
  assign new_R140_U400 = ~new_R140_U145 | ~new_R140_U146;
  assign new_R140_U401 = ~new_R140_U277 | ~new_R140_U399;
  assign new_R140_U402 = ~new_U99 | ~new_R140_U73;
  assign new_R140_U403 = ~SI_28_ | ~new_R140_U74;
  assign new_R140_U404 = ~new_U99 | ~new_R140_U73;
  assign new_R140_U405 = ~SI_28_ | ~new_R140_U74;
  assign new_R140_U406 = ~new_R140_U405 | ~new_R140_U404;
  assign new_R140_U407 = ~new_R140_U147 | ~new_R140_U148;
  assign new_R140_U408 = ~new_R140_U273 | ~new_R140_U406;
  assign new_R140_U409 = ~new_U100 | ~new_R140_U71;
  assign new_R140_U410 = ~SI_27_ | ~new_R140_U72;
  assign new_R140_U411 = ~new_U100 | ~new_R140_U71;
  assign new_R140_U412 = ~SI_27_ | ~new_R140_U72;
  assign new_R140_U413 = ~new_R140_U412 | ~new_R140_U411;
  assign new_R140_U414 = ~new_R140_U149 | ~new_R140_U150;
  assign new_R140_U415 = ~new_R140_U269 | ~new_R140_U413;
  assign new_R140_U416 = ~new_U101 | ~new_R140_U69;
  assign new_R140_U417 = ~SI_26_ | ~new_R140_U70;
  assign new_R140_U418 = ~new_U101 | ~new_R140_U69;
  assign new_R140_U419 = ~SI_26_ | ~new_R140_U70;
  assign new_R140_U420 = ~new_R140_U419 | ~new_R140_U418;
  assign new_R140_U421 = ~new_R140_U151 | ~new_R140_U152;
  assign new_R140_U422 = ~new_R140_U265 | ~new_R140_U420;
  assign new_R140_U423 = ~new_U102 | ~new_R140_U67;
  assign new_R140_U424 = ~SI_25_ | ~new_R140_U68;
  assign new_R140_U425 = ~new_U102 | ~new_R140_U67;
  assign new_R140_U426 = ~SI_25_ | ~new_R140_U68;
  assign new_R140_U427 = ~new_R140_U426 | ~new_R140_U425;
  assign new_R140_U428 = ~new_R140_U153 | ~new_R140_U154;
  assign new_R140_U429 = ~new_R140_U261 | ~new_R140_U427;
  assign new_R140_U430 = ~new_U103 | ~new_R140_U65;
  assign new_R140_U431 = ~SI_24_ | ~new_R140_U66;
  assign new_R140_U432 = ~new_U103 | ~new_R140_U65;
  assign new_R140_U433 = ~SI_24_ | ~new_R140_U66;
  assign new_R140_U434 = ~new_R140_U433 | ~new_R140_U432;
  assign new_R140_U435 = ~new_R140_U155 | ~new_R140_U156;
  assign new_R140_U436 = ~new_R140_U257 | ~new_R140_U434;
  assign new_R140_U437 = ~new_U104 | ~new_R140_U63;
  assign new_R140_U438 = ~SI_23_ | ~new_R140_U64;
  assign new_R140_U439 = ~new_U104 | ~new_R140_U63;
  assign new_R140_U440 = ~SI_23_ | ~new_R140_U64;
  assign new_R140_U441 = ~new_R140_U440 | ~new_R140_U439;
  assign new_R140_U442 = ~new_R140_U157 | ~new_R140_U158;
  assign new_R140_U443 = ~new_R140_U253 | ~new_R140_U441;
  assign new_R140_U444 = ~new_U105 | ~new_R140_U61;
  assign new_R140_U445 = ~SI_22_ | ~new_R140_U62;
  assign new_R140_U446 = ~new_U105 | ~new_R140_U61;
  assign new_R140_U447 = ~SI_22_ | ~new_R140_U62;
  assign new_R140_U448 = ~new_R140_U447 | ~new_R140_U446;
  assign new_R140_U449 = ~new_R140_U159 | ~new_R140_U160;
  assign new_R140_U450 = ~new_R140_U249 | ~new_R140_U448;
  assign new_R140_U451 = ~new_U106 | ~new_R140_U59;
  assign new_R140_U452 = ~SI_21_ | ~new_R140_U60;
  assign new_R140_U453 = ~new_U106 | ~new_R140_U59;
  assign new_R140_U454 = ~SI_21_ | ~new_R140_U60;
  assign new_R140_U455 = ~new_R140_U454 | ~new_R140_U453;
  assign new_R140_U456 = ~new_R140_U161 | ~new_R140_U162;
  assign new_R140_U457 = ~new_R140_U245 | ~new_R140_U455;
  assign new_R140_U458 = ~new_U107 | ~new_R140_U57;
  assign new_R140_U459 = ~SI_20_ | ~new_R140_U58;
  assign new_R140_U460 = ~new_U107 | ~new_R140_U57;
  assign new_R140_U461 = ~SI_20_ | ~new_R140_U58;
  assign new_R140_U462 = ~new_R140_U461 | ~new_R140_U460;
  assign new_R140_U463 = ~new_R140_U163 | ~new_R140_U164;
  assign new_R140_U464 = ~new_R140_U241 | ~new_R140_U462;
  assign new_R140_U465 = ~new_U119 | ~new_R140_U165;
  assign new_R140_U466 = ~new_R140_U187 | ~new_R140_U32;
  assign new_R140_U467 = ~new_R140_U466 | ~new_R140_U465;
  assign new_R140_U468 = ~SI_1_ | ~new_R140_U165 | ~new_R140_U32;
  assign new_R140_U469 = ~new_R140_U467 | ~new_R140_U29;
  assign new_R140_U470 = ~new_U109 | ~new_R140_U55;
  assign new_R140_U471 = ~SI_19_ | ~new_R140_U56;
  assign new_R140_U472 = ~new_U109 | ~new_R140_U55;
  assign new_R140_U473 = ~SI_19_ | ~new_R140_U56;
  assign new_R140_U474 = ~new_R140_U473 | ~new_R140_U472;
  assign new_R140_U475 = ~new_R140_U166 | ~new_R140_U167;
  assign new_R140_U476 = ~new_R140_U237 | ~new_R140_U474;
  assign new_R140_U477 = ~new_U110 | ~new_R140_U53;
  assign new_R140_U478 = ~SI_18_ | ~new_R140_U54;
  assign new_R140_U479 = ~new_U110 | ~new_R140_U53;
  assign new_R140_U480 = ~SI_18_ | ~new_R140_U54;
  assign new_R140_U481 = ~new_R140_U480 | ~new_R140_U479;
  assign new_R140_U482 = ~new_R140_U168 | ~new_R140_U169;
  assign new_R140_U483 = ~new_R140_U233 | ~new_R140_U481;
  assign new_R140_U484 = ~new_U111 | ~new_R140_U51;
  assign new_R140_U485 = ~SI_17_ | ~new_R140_U52;
  assign new_R140_U486 = ~new_U111 | ~new_R140_U51;
  assign new_R140_U487 = ~SI_17_ | ~new_R140_U52;
  assign new_R140_U488 = ~new_R140_U487 | ~new_R140_U486;
  assign new_R140_U489 = ~new_R140_U170 | ~new_R140_U171;
  assign new_R140_U490 = ~new_R140_U229 | ~new_R140_U488;
  assign new_R140_U491 = ~new_U112 | ~new_R140_U49;
  assign new_R140_U492 = ~SI_16_ | ~new_R140_U50;
  assign new_R140_U493 = ~new_U112 | ~new_R140_U49;
  assign new_R140_U494 = ~SI_16_ | ~new_R140_U50;
  assign new_R140_U495 = ~new_R140_U494 | ~new_R140_U493;
  assign new_R140_U496 = ~new_R140_U172 | ~new_R140_U173;
  assign new_R140_U497 = ~new_R140_U225 | ~new_R140_U495;
  assign new_R140_U498 = ~new_U113 | ~new_R140_U47;
  assign new_R140_U499 = ~SI_15_ | ~new_R140_U48;
  assign new_R140_U500 = ~new_U113 | ~new_R140_U47;
  assign new_R140_U501 = ~SI_15_ | ~new_R140_U48;
  assign new_R140_U502 = ~new_R140_U501 | ~new_R140_U500;
  assign new_R140_U503 = ~new_R140_U174 | ~new_R140_U175;
  assign new_R140_U504 = ~new_R140_U221 | ~new_R140_U502;
  assign new_R140_U505 = ~new_U114 | ~new_R140_U36;
  assign new_R140_U506 = ~SI_14_ | ~new_R140_U37;
  assign new_R140_U507 = ~new_U114 | ~new_R140_U36;
  assign new_R140_U508 = ~SI_14_ | ~new_R140_U37;
  assign new_R140_U509 = ~new_R140_U508 | ~new_R140_U507;
  assign new_R140_U510 = ~new_R140_U176 | ~new_R140_U177;
  assign new_R140_U511 = ~new_R140_U218 | ~new_R140_U509;
  assign new_R140_U512 = ~new_U115 | ~new_R140_U40;
  assign new_R140_U513 = ~SI_13_ | ~new_R140_U41;
  assign new_R140_U514 = ~new_U115 | ~new_R140_U40;
  assign new_R140_U515 = ~SI_13_ | ~new_R140_U41;
  assign new_R140_U516 = ~new_R140_U515 | ~new_R140_U514;
  assign new_R140_U517 = ~new_R140_U178 | ~new_R140_U179;
  assign new_R140_U518 = ~new_R140_U215 | ~new_R140_U516;
  assign new_R140_U519 = ~new_U116 | ~new_R140_U42;
  assign new_R140_U520 = ~SI_12_ | ~new_R140_U43;
  assign new_R140_U521 = ~new_U116 | ~new_R140_U42;
  assign new_R140_U522 = ~SI_12_ | ~new_R140_U43;
  assign new_R140_U523 = ~new_R140_U522 | ~new_R140_U521;
  assign new_R140_U524 = ~new_R140_U180 | ~new_R140_U181;
  assign new_R140_U525 = ~new_R140_U212 | ~new_R140_U523;
  assign new_R140_U526 = ~new_U117 | ~new_R140_U44;
  assign new_R140_U527 = ~SI_11_ | ~new_R140_U45;
  assign new_R140_U528 = ~new_U117 | ~new_R140_U44;
  assign new_R140_U529 = ~SI_11_ | ~new_R140_U45;
  assign new_R140_U530 = ~new_R140_U529 | ~new_R140_U528;
  assign new_R140_U531 = ~new_R140_U182 | ~new_R140_U183;
  assign new_R140_U532 = ~new_R140_U314 | ~new_R140_U530;
  assign new_R140_U533 = ~new_U118 | ~new_R140_U38;
  assign new_R140_U534 = ~SI_10_ | ~new_R140_U39;
  assign new_R140_U535 = ~new_U118 | ~new_R140_U38;
  assign new_R140_U536 = ~SI_10_ | ~new_R140_U39;
  assign new_R140_U537 = ~new_R140_U536 | ~new_R140_U535;
  assign new_R140_U538 = ~new_R140_U184 | ~new_R140_U185;
  assign new_R140_U539 = ~new_R140_U312 | ~new_R140_U537;
  assign new_R140_U540 = ~new_U120 | ~new_R140_U30;
  assign new_R140_U541 = ~SI_0_ | ~new_R140_U31;
  assign new_LT_1075_19_U6 = ~P2_ADDR_REG_19_;
  assign new_P1_ADD_95_U4 = ~P1_REG3_REG_3_;
  assign new_P1_ADD_95_U5 = new_P1_ADD_95_U102 & P1_REG3_REG_28_ & P1_REG3_REG_27_;
  assign new_P1_ADD_95_U6 = ~P1_REG3_REG_4_;
  assign new_P1_ADD_95_U7 = ~P1_REG3_REG_4_ | ~P1_REG3_REG_3_;
  assign new_P1_ADD_95_U8 = ~P1_REG3_REG_5_;
  assign new_P1_ADD_95_U9 = ~P1_REG3_REG_5_ | ~new_P1_ADD_95_U80;
  assign new_P1_ADD_95_U10 = ~P1_REG3_REG_6_;
  assign new_P1_ADD_95_U11 = ~P1_REG3_REG_6_ | ~new_P1_ADD_95_U81;
  assign new_P1_ADD_95_U12 = ~P1_REG3_REG_7_;
  assign new_P1_ADD_95_U13 = ~P1_REG3_REG_7_ | ~new_P1_ADD_95_U82;
  assign new_P1_ADD_95_U14 = ~P1_REG3_REG_8_;
  assign new_P1_ADD_95_U15 = ~P1_REG3_REG_9_;
  assign new_P1_ADD_95_U16 = ~P1_REG3_REG_8_ | ~new_P1_ADD_95_U83;
  assign new_P1_ADD_95_U17 = ~new_P1_ADD_95_U84 | ~P1_REG3_REG_9_;
  assign new_P1_ADD_95_U18 = ~P1_REG3_REG_10_;
  assign new_P1_ADD_95_U19 = ~P1_REG3_REG_10_ | ~new_P1_ADD_95_U85;
  assign new_P1_ADD_95_U20 = ~P1_REG3_REG_11_;
  assign new_P1_ADD_95_U21 = ~P1_REG3_REG_11_ | ~new_P1_ADD_95_U86;
  assign new_P1_ADD_95_U22 = ~P1_REG3_REG_12_;
  assign new_P1_ADD_95_U23 = ~P1_REG3_REG_12_ | ~new_P1_ADD_95_U87;
  assign new_P1_ADD_95_U24 = ~P1_REG3_REG_13_;
  assign new_P1_ADD_95_U25 = ~P1_REG3_REG_13_ | ~new_P1_ADD_95_U88;
  assign new_P1_ADD_95_U26 = ~P1_REG3_REG_14_;
  assign new_P1_ADD_95_U27 = ~P1_REG3_REG_14_ | ~new_P1_ADD_95_U89;
  assign new_P1_ADD_95_U28 = ~P1_REG3_REG_15_;
  assign new_P1_ADD_95_U29 = ~P1_REG3_REG_15_ | ~new_P1_ADD_95_U90;
  assign new_P1_ADD_95_U30 = ~P1_REG3_REG_16_;
  assign new_P1_ADD_95_U31 = ~P1_REG3_REG_16_ | ~new_P1_ADD_95_U91;
  assign new_P1_ADD_95_U32 = ~P1_REG3_REG_17_;
  assign new_P1_ADD_95_U33 = ~P1_REG3_REG_17_ | ~new_P1_ADD_95_U92;
  assign new_P1_ADD_95_U34 = ~P1_REG3_REG_18_;
  assign new_P1_ADD_95_U35 = ~P1_REG3_REG_18_ | ~new_P1_ADD_95_U93;
  assign new_P1_ADD_95_U36 = ~P1_REG3_REG_19_;
  assign new_P1_ADD_95_U37 = ~P1_REG3_REG_19_ | ~new_P1_ADD_95_U94;
  assign new_P1_ADD_95_U38 = ~P1_REG3_REG_20_;
  assign new_P1_ADD_95_U39 = ~P1_REG3_REG_20_ | ~new_P1_ADD_95_U95;
  assign new_P1_ADD_95_U40 = ~P1_REG3_REG_21_;
  assign new_P1_ADD_95_U41 = ~P1_REG3_REG_21_ | ~new_P1_ADD_95_U96;
  assign new_P1_ADD_95_U42 = ~P1_REG3_REG_22_;
  assign new_P1_ADD_95_U43 = ~P1_REG3_REG_22_ | ~new_P1_ADD_95_U97;
  assign new_P1_ADD_95_U44 = ~P1_REG3_REG_23_;
  assign new_P1_ADD_95_U45 = ~P1_REG3_REG_23_ | ~new_P1_ADD_95_U98;
  assign new_P1_ADD_95_U46 = ~P1_REG3_REG_24_;
  assign new_P1_ADD_95_U47 = ~P1_REG3_REG_24_ | ~new_P1_ADD_95_U99;
  assign new_P1_ADD_95_U48 = ~P1_REG3_REG_25_;
  assign new_P1_ADD_95_U49 = ~P1_REG3_REG_25_ | ~new_P1_ADD_95_U100;
  assign new_P1_ADD_95_U50 = ~P1_REG3_REG_26_;
  assign new_P1_ADD_95_U51 = ~P1_REG3_REG_26_ | ~new_P1_ADD_95_U101;
  assign new_P1_ADD_95_U52 = ~P1_REG3_REG_28_;
  assign new_P1_ADD_95_U53 = ~P1_REG3_REG_27_;
  assign new_P1_ADD_95_U54 = ~new_P1_ADD_95_U105 | ~new_P1_ADD_95_U104;
  assign new_P1_ADD_95_U55 = ~new_P1_ADD_95_U107 | ~new_P1_ADD_95_U106;
  assign new_P1_ADD_95_U56 = ~new_P1_ADD_95_U109 | ~new_P1_ADD_95_U108;
  assign new_P1_ADD_95_U57 = ~new_P1_ADD_95_U111 | ~new_P1_ADD_95_U110;
  assign new_P1_ADD_95_U58 = ~new_P1_ADD_95_U113 | ~new_P1_ADD_95_U112;
  assign new_P1_ADD_95_U59 = ~new_P1_ADD_95_U115 | ~new_P1_ADD_95_U114;
  assign new_P1_ADD_95_U60 = ~new_P1_ADD_95_U117 | ~new_P1_ADD_95_U116;
  assign new_P1_ADD_95_U61 = ~new_P1_ADD_95_U119 | ~new_P1_ADD_95_U118;
  assign new_P1_ADD_95_U62 = ~new_P1_ADD_95_U121 | ~new_P1_ADD_95_U120;
  assign new_P1_ADD_95_U63 = ~new_P1_ADD_95_U123 | ~new_P1_ADD_95_U122;
  assign new_P1_ADD_95_U64 = ~new_P1_ADD_95_U125 | ~new_P1_ADD_95_U124;
  assign new_P1_ADD_95_U65 = ~new_P1_ADD_95_U127 | ~new_P1_ADD_95_U126;
  assign new_P1_ADD_95_U66 = ~new_P1_ADD_95_U129 | ~new_P1_ADD_95_U128;
  assign new_P1_ADD_95_U67 = ~new_P1_ADD_95_U131 | ~new_P1_ADD_95_U130;
  assign new_P1_ADD_95_U68 = ~new_P1_ADD_95_U133 | ~new_P1_ADD_95_U132;
  assign new_P1_ADD_95_U69 = ~new_P1_ADD_95_U135 | ~new_P1_ADD_95_U134;
  assign new_P1_ADD_95_U70 = ~new_P1_ADD_95_U137 | ~new_P1_ADD_95_U136;
  assign new_P1_ADD_95_U71 = ~new_P1_ADD_95_U139 | ~new_P1_ADD_95_U138;
  assign new_P1_ADD_95_U72 = ~new_P1_ADD_95_U141 | ~new_P1_ADD_95_U140;
  assign new_P1_ADD_95_U73 = ~new_P1_ADD_95_U143 | ~new_P1_ADD_95_U142;
  assign new_P1_ADD_95_U74 = ~new_P1_ADD_95_U145 | ~new_P1_ADD_95_U144;
  assign new_P1_ADD_95_U75 = ~new_P1_ADD_95_U147 | ~new_P1_ADD_95_U146;
  assign new_P1_ADD_95_U76 = ~new_P1_ADD_95_U149 | ~new_P1_ADD_95_U148;
  assign new_P1_ADD_95_U77 = ~new_P1_ADD_95_U151 | ~new_P1_ADD_95_U150;
  assign new_P1_ADD_95_U78 = ~new_P1_ADD_95_U153 | ~new_P1_ADD_95_U152;
  assign new_P1_ADD_95_U79 = ~P1_REG3_REG_27_ | ~new_P1_ADD_95_U102;
  assign new_P1_ADD_95_U80 = ~new_P1_ADD_95_U7;
  assign new_P1_ADD_95_U81 = ~new_P1_ADD_95_U9;
  assign new_P1_ADD_95_U82 = ~new_P1_ADD_95_U11;
  assign new_P1_ADD_95_U83 = ~new_P1_ADD_95_U13;
  assign new_P1_ADD_95_U84 = ~new_P1_ADD_95_U16;
  assign new_P1_ADD_95_U85 = ~new_P1_ADD_95_U17;
  assign new_P1_ADD_95_U86 = ~new_P1_ADD_95_U19;
  assign new_P1_ADD_95_U87 = ~new_P1_ADD_95_U21;
  assign new_P1_ADD_95_U88 = ~new_P1_ADD_95_U23;
  assign new_P1_ADD_95_U89 = ~new_P1_ADD_95_U25;
  assign new_P1_ADD_95_U90 = ~new_P1_ADD_95_U27;
  assign new_P1_ADD_95_U91 = ~new_P1_ADD_95_U29;
  assign new_P1_ADD_95_U92 = ~new_P1_ADD_95_U31;
  assign new_P1_ADD_95_U93 = ~new_P1_ADD_95_U33;
  assign new_P1_ADD_95_U94 = ~new_P1_ADD_95_U35;
  assign new_P1_ADD_95_U95 = ~new_P1_ADD_95_U37;
  assign new_P1_ADD_95_U96 = ~new_P1_ADD_95_U39;
  assign new_P1_ADD_95_U97 = ~new_P1_ADD_95_U41;
  assign new_P1_ADD_95_U98 = ~new_P1_ADD_95_U43;
  assign new_P1_ADD_95_U99 = ~new_P1_ADD_95_U45;
  assign new_P1_ADD_95_U100 = ~new_P1_ADD_95_U47;
  assign new_P1_ADD_95_U101 = ~new_P1_ADD_95_U49;
  assign new_P1_ADD_95_U102 = ~new_P1_ADD_95_U51;
  assign new_P1_ADD_95_U103 = ~new_P1_ADD_95_U79;
  assign new_P1_ADD_95_U104 = ~P1_REG3_REG_9_ | ~new_P1_ADD_95_U16;
  assign new_P1_ADD_95_U105 = ~new_P1_ADD_95_U84 | ~new_P1_ADD_95_U15;
  assign new_P1_ADD_95_U106 = ~P1_REG3_REG_8_ | ~new_P1_ADD_95_U13;
  assign new_P1_ADD_95_U107 = ~new_P1_ADD_95_U83 | ~new_P1_ADD_95_U14;
  assign new_P1_ADD_95_U108 = ~P1_REG3_REG_7_ | ~new_P1_ADD_95_U11;
  assign new_P1_ADD_95_U109 = ~new_P1_ADD_95_U82 | ~new_P1_ADD_95_U12;
  assign new_P1_ADD_95_U110 = ~P1_REG3_REG_6_ | ~new_P1_ADD_95_U9;
  assign new_P1_ADD_95_U111 = ~new_P1_ADD_95_U81 | ~new_P1_ADD_95_U10;
  assign new_P1_ADD_95_U112 = ~P1_REG3_REG_5_ | ~new_P1_ADD_95_U7;
  assign new_P1_ADD_95_U113 = ~new_P1_ADD_95_U80 | ~new_P1_ADD_95_U8;
  assign new_P1_ADD_95_U114 = ~P1_REG3_REG_4_ | ~new_P1_ADD_95_U4;
  assign new_P1_ADD_95_U115 = ~P1_REG3_REG_3_ | ~new_P1_ADD_95_U6;
  assign new_P1_ADD_95_U116 = ~P1_REG3_REG_28_ | ~new_P1_ADD_95_U79;
  assign new_P1_ADD_95_U117 = ~new_P1_ADD_95_U103 | ~new_P1_ADD_95_U52;
  assign new_P1_ADD_95_U118 = ~P1_REG3_REG_27_ | ~new_P1_ADD_95_U51;
  assign new_P1_ADD_95_U119 = ~new_P1_ADD_95_U102 | ~new_P1_ADD_95_U53;
  assign new_P1_ADD_95_U120 = ~P1_REG3_REG_26_ | ~new_P1_ADD_95_U49;
  assign new_P1_ADD_95_U121 = ~new_P1_ADD_95_U101 | ~new_P1_ADD_95_U50;
  assign new_P1_ADD_95_U122 = ~P1_REG3_REG_25_ | ~new_P1_ADD_95_U47;
  assign new_P1_ADD_95_U123 = ~new_P1_ADD_95_U100 | ~new_P1_ADD_95_U48;
  assign new_P1_ADD_95_U124 = ~P1_REG3_REG_24_ | ~new_P1_ADD_95_U45;
  assign new_P1_ADD_95_U125 = ~new_P1_ADD_95_U99 | ~new_P1_ADD_95_U46;
  assign new_P1_ADD_95_U126 = ~P1_REG3_REG_23_ | ~new_P1_ADD_95_U43;
  assign new_P1_ADD_95_U127 = ~new_P1_ADD_95_U98 | ~new_P1_ADD_95_U44;
  assign new_P1_ADD_95_U128 = ~P1_REG3_REG_22_ | ~new_P1_ADD_95_U41;
  assign new_P1_ADD_95_U129 = ~new_P1_ADD_95_U97 | ~new_P1_ADD_95_U42;
  assign new_P1_ADD_95_U130 = ~P1_REG3_REG_21_ | ~new_P1_ADD_95_U39;
  assign new_P1_ADD_95_U131 = ~new_P1_ADD_95_U96 | ~new_P1_ADD_95_U40;
  assign new_P1_ADD_95_U132 = ~P1_REG3_REG_20_ | ~new_P1_ADD_95_U37;
  assign new_P1_ADD_95_U133 = ~new_P1_ADD_95_U95 | ~new_P1_ADD_95_U38;
  assign new_P1_ADD_95_U134 = ~P1_REG3_REG_19_ | ~new_P1_ADD_95_U35;
  assign new_P1_ADD_95_U135 = ~new_P1_ADD_95_U94 | ~new_P1_ADD_95_U36;
  assign new_P1_ADD_95_U136 = ~P1_REG3_REG_18_ | ~new_P1_ADD_95_U33;
  assign new_P1_ADD_95_U137 = ~new_P1_ADD_95_U93 | ~new_P1_ADD_95_U34;
  assign new_P1_ADD_95_U138 = ~P1_REG3_REG_17_ | ~new_P1_ADD_95_U31;
  assign new_P1_ADD_95_U139 = ~new_P1_ADD_95_U92 | ~new_P1_ADD_95_U32;
  assign new_P1_ADD_95_U140 = ~P1_REG3_REG_16_ | ~new_P1_ADD_95_U29;
  assign new_P1_ADD_95_U141 = ~new_P1_ADD_95_U91 | ~new_P1_ADD_95_U30;
  assign new_P1_ADD_95_U142 = ~P1_REG3_REG_15_ | ~new_P1_ADD_95_U27;
  assign new_P1_ADD_95_U143 = ~new_P1_ADD_95_U90 | ~new_P1_ADD_95_U28;
  assign new_P1_ADD_95_U144 = ~P1_REG3_REG_14_ | ~new_P1_ADD_95_U25;
  assign new_P1_ADD_95_U145 = ~new_P1_ADD_95_U89 | ~new_P1_ADD_95_U26;
  assign new_P1_ADD_95_U146 = ~P1_REG3_REG_13_ | ~new_P1_ADD_95_U23;
  assign new_P1_ADD_95_U147 = ~new_P1_ADD_95_U88 | ~new_P1_ADD_95_U24;
  assign new_P1_ADD_95_U148 = ~P1_REG3_REG_12_ | ~new_P1_ADD_95_U21;
  assign new_P1_ADD_95_U149 = ~new_P1_ADD_95_U87 | ~new_P1_ADD_95_U22;
  assign new_P1_ADD_95_U150 = ~P1_REG3_REG_11_ | ~new_P1_ADD_95_U19;
  assign new_P1_ADD_95_U151 = ~new_P1_ADD_95_U86 | ~new_P1_ADD_95_U20;
  assign new_P1_ADD_95_U152 = ~P1_REG3_REG_10_ | ~new_P1_ADD_95_U17;
  assign new_P1_ADD_95_U153 = ~new_P1_ADD_95_U85 | ~new_P1_ADD_95_U18;
  assign new_P1_R1105_U4 = new_P1_R1105_U95 & new_P1_R1105_U94;
  assign new_P1_R1105_U5 = new_P1_R1105_U96 & new_P1_R1105_U97;
  assign new_P1_R1105_U6 = new_P1_R1105_U113 & new_P1_R1105_U112;
  assign new_P1_R1105_U7 = new_P1_R1105_U155 & new_P1_R1105_U154;
  assign new_P1_R1105_U8 = new_P1_R1105_U164 & new_P1_R1105_U163;
  assign new_P1_R1105_U9 = new_P1_R1105_U182 & new_P1_R1105_U181;
  assign new_P1_R1105_U10 = new_P1_R1105_U218 & new_P1_R1105_U215;
  assign new_P1_R1105_U11 = new_P1_R1105_U211 & new_P1_R1105_U208;
  assign new_P1_R1105_U12 = new_P1_R1105_U202 & new_P1_R1105_U199;
  assign new_P1_R1105_U13 = new_P1_R1105_U196 & new_P1_R1105_U192;
  assign new_P1_R1105_U14 = new_P1_R1105_U151 & new_P1_R1105_U148;
  assign new_P1_R1105_U15 = new_P1_R1105_U143 & new_P1_R1105_U140;
  assign new_P1_R1105_U16 = new_P1_R1105_U129 & new_P1_R1105_U126;
  assign new_P1_R1105_U17 = ~P1_REG2_REG_6_;
  assign new_P1_R1105_U18 = ~new_P1_U3469;
  assign new_P1_R1105_U19 = ~new_P1_U3472;
  assign new_P1_R1105_U20 = ~new_P1_U3469 | ~P1_REG2_REG_6_;
  assign new_P1_R1105_U21 = ~P1_REG2_REG_7_;
  assign new_P1_R1105_U22 = ~P1_REG2_REG_4_;
  assign new_P1_R1105_U23 = ~new_P1_U3463;
  assign new_P1_R1105_U24 = ~new_P1_U3466;
  assign new_P1_R1105_U25 = ~P1_REG2_REG_2_;
  assign new_P1_R1105_U26 = ~new_P1_U3457;
  assign new_P1_R1105_U27 = ~P1_REG2_REG_0_;
  assign new_P1_R1105_U28 = ~new_P1_U3448;
  assign new_P1_R1105_U29 = ~new_P1_U3448 | ~P1_REG2_REG_0_;
  assign new_P1_R1105_U30 = ~P1_REG2_REG_3_;
  assign new_P1_R1105_U31 = ~new_P1_U3460;
  assign new_P1_R1105_U32 = ~new_P1_U3463 | ~P1_REG2_REG_4_;
  assign new_P1_R1105_U33 = ~P1_REG2_REG_5_;
  assign new_P1_R1105_U34 = ~P1_REG2_REG_8_;
  assign new_P1_R1105_U35 = ~new_P1_U3475;
  assign new_P1_R1105_U36 = ~new_P1_U3478;
  assign new_P1_R1105_U37 = ~P1_REG2_REG_9_;
  assign new_P1_R1105_U38 = ~new_P1_R1105_U49 | ~new_P1_R1105_U121;
  assign new_P1_R1105_U39 = ~new_P1_R1105_U109 | ~new_P1_R1105_U110 | ~new_P1_R1105_U108;
  assign new_P1_R1105_U40 = ~new_P1_R1105_U98 | ~new_P1_R1105_U99;
  assign new_P1_R1105_U41 = ~P1_REG2_REG_1_ | ~new_P1_U3454;
  assign new_P1_R1105_U42 = ~new_P1_R1105_U135 | ~new_P1_R1105_U136 | ~new_P1_R1105_U134;
  assign new_P1_R1105_U43 = ~new_P1_R1105_U132 | ~new_P1_R1105_U131;
  assign new_P1_R1105_U44 = ~P1_REG2_REG_16_;
  assign new_P1_R1105_U45 = ~new_P1_U3499;
  assign new_P1_R1105_U46 = ~new_P1_U3502;
  assign new_P1_R1105_U47 = ~new_P1_U3499 | ~P1_REG2_REG_16_;
  assign new_P1_R1105_U48 = ~P1_REG2_REG_17_;
  assign new_P1_R1105_U49 = ~new_P1_U3475 | ~P1_REG2_REG_8_;
  assign new_P1_R1105_U50 = ~P1_REG2_REG_10_;
  assign new_P1_R1105_U51 = ~new_P1_U3481;
  assign new_P1_R1105_U52 = ~P1_REG2_REG_12_;
  assign new_P1_R1105_U53 = ~new_P1_U3487;
  assign new_P1_R1105_U54 = ~P1_REG2_REG_11_;
  assign new_P1_R1105_U55 = ~new_P1_U3484;
  assign new_P1_R1105_U56 = ~new_P1_U3484 | ~P1_REG2_REG_11_;
  assign new_P1_R1105_U57 = ~P1_REG2_REG_13_;
  assign new_P1_R1105_U58 = ~new_P1_U3490;
  assign new_P1_R1105_U59 = ~P1_REG2_REG_14_;
  assign new_P1_R1105_U60 = ~new_P1_U3493;
  assign new_P1_R1105_U61 = ~P1_REG2_REG_15_;
  assign new_P1_R1105_U62 = ~new_P1_U3496;
  assign new_P1_R1105_U63 = ~P1_REG2_REG_18_;
  assign new_P1_R1105_U64 = ~new_P1_U3505;
  assign new_P1_R1105_U65 = ~new_P1_R1105_U187 | ~new_P1_R1105_U186 | ~new_P1_R1105_U185;
  assign new_P1_R1105_U66 = ~new_P1_R1105_U179 | ~new_P1_R1105_U178;
  assign new_P1_R1105_U67 = ~new_P1_R1105_U56 | ~new_P1_R1105_U204;
  assign new_P1_R1105_U68 = ~new_P1_R1105_U259 | ~new_P1_R1105_U258;
  assign new_P1_R1105_U69 = ~new_P1_R1105_U308 | ~new_P1_R1105_U307;
  assign new_P1_R1105_U70 = ~new_P1_R1105_U231 | ~new_P1_R1105_U230;
  assign new_P1_R1105_U71 = ~new_P1_R1105_U236 | ~new_P1_R1105_U235;
  assign new_P1_R1105_U72 = ~new_P1_R1105_U243 | ~new_P1_R1105_U242;
  assign new_P1_R1105_U73 = ~new_P1_R1105_U250 | ~new_P1_R1105_U249;
  assign new_P1_R1105_U74 = ~new_P1_R1105_U255 | ~new_P1_R1105_U254;
  assign new_P1_R1105_U75 = ~new_P1_R1105_U271 | ~new_P1_R1105_U270;
  assign new_P1_R1105_U76 = ~new_P1_R1105_U278 | ~new_P1_R1105_U277;
  assign new_P1_R1105_U77 = ~new_P1_R1105_U285 | ~new_P1_R1105_U284;
  assign new_P1_R1105_U78 = ~new_P1_R1105_U292 | ~new_P1_R1105_U291;
  assign new_P1_R1105_U79 = ~new_P1_R1105_U299 | ~new_P1_R1105_U298;
  assign new_P1_R1105_U80 = ~new_P1_R1105_U304 | ~new_P1_R1105_U303;
  assign new_P1_R1105_U81 = ~new_P1_R1105_U118 | ~new_P1_R1105_U117 | ~new_P1_R1105_U116;
  assign new_P1_R1105_U82 = ~new_P1_R1105_U133 | ~new_P1_R1105_U145;
  assign new_P1_R1105_U83 = ~new_P1_R1105_U41 | ~new_P1_R1105_U152;
  assign new_P1_R1105_U84 = ~new_P1_U3442;
  assign new_P1_R1105_U85 = ~P1_REG2_REG_19_;
  assign new_P1_R1105_U86 = ~new_P1_R1105_U175 | ~new_P1_R1105_U174;
  assign new_P1_R1105_U87 = ~new_P1_R1105_U171 | ~new_P1_R1105_U170;
  assign new_P1_R1105_U88 = ~new_P1_R1105_U161 | ~new_P1_R1105_U160;
  assign new_P1_R1105_U89 = ~new_P1_R1105_U32;
  assign new_P1_R1105_U90 = ~P1_REG2_REG_9_ | ~new_P1_U3478;
  assign new_P1_R1105_U91 = ~new_P1_U3487 | ~P1_REG2_REG_12_;
  assign new_P1_R1105_U92 = ~new_P1_R1105_U56;
  assign new_P1_R1105_U93 = ~new_P1_R1105_U49;
  assign new_P1_R1105_U94 = new_P1_U3466 | P1_REG2_REG_5_;
  assign new_P1_R1105_U95 = new_P1_U3463 | P1_REG2_REG_4_;
  assign new_P1_R1105_U96 = P1_REG2_REG_3_ | new_P1_U3460;
  assign new_P1_R1105_U97 = P1_REG2_REG_2_ | new_P1_U3457;
  assign new_P1_R1105_U98 = ~new_P1_R1105_U29;
  assign new_P1_R1105_U99 = P1_REG2_REG_1_ | new_P1_U3454;
  assign new_P1_R1105_U100 = ~new_P1_R1105_U40;
  assign new_P1_R1105_U101 = ~new_P1_R1105_U41;
  assign new_P1_R1105_U102 = ~new_P1_R1105_U40 | ~new_P1_R1105_U41;
  assign new_P1_R1105_U103 = ~new_P1_R1105_U96 | ~P1_REG2_REG_2_ | ~new_P1_U3457;
  assign new_P1_R1105_U104 = ~new_P1_R1105_U5 | ~new_P1_R1105_U102;
  assign new_P1_R1105_U105 = ~new_P1_U3460 | ~P1_REG2_REG_3_;
  assign new_P1_R1105_U106 = ~new_P1_R1105_U104 | ~new_P1_R1105_U105 | ~new_P1_R1105_U103;
  assign new_P1_R1105_U107 = ~new_P1_R1105_U33 | ~new_P1_R1105_U32;
  assign new_P1_R1105_U108 = ~new_P1_U3466 | ~new_P1_R1105_U107;
  assign new_P1_R1105_U109 = ~new_P1_R1105_U4 | ~new_P1_R1105_U106;
  assign new_P1_R1105_U110 = ~P1_REG2_REG_5_ | ~new_P1_R1105_U89;
  assign new_P1_R1105_U111 = ~new_P1_R1105_U39;
  assign new_P1_R1105_U112 = new_P1_U3472 | P1_REG2_REG_7_;
  assign new_P1_R1105_U113 = new_P1_U3469 | P1_REG2_REG_6_;
  assign new_P1_R1105_U114 = ~new_P1_R1105_U20;
  assign new_P1_R1105_U115 = ~new_P1_R1105_U21 | ~new_P1_R1105_U20;
  assign new_P1_R1105_U116 = ~new_P1_U3472 | ~new_P1_R1105_U115;
  assign new_P1_R1105_U117 = ~P1_REG2_REG_7_ | ~new_P1_R1105_U114;
  assign new_P1_R1105_U118 = ~new_P1_R1105_U6 | ~new_P1_R1105_U39;
  assign new_P1_R1105_U119 = ~new_P1_R1105_U81;
  assign new_P1_R1105_U120 = P1_REG2_REG_8_ | new_P1_U3475;
  assign new_P1_R1105_U121 = ~new_P1_R1105_U120 | ~new_P1_R1105_U81;
  assign new_P1_R1105_U122 = ~new_P1_R1105_U38;
  assign new_P1_R1105_U123 = new_P1_U3478 | P1_REG2_REG_9_;
  assign new_P1_R1105_U124 = P1_REG2_REG_6_ | new_P1_U3469;
  assign new_P1_R1105_U125 = ~new_P1_R1105_U124 | ~new_P1_R1105_U39;
  assign new_P1_R1105_U126 = ~new_P1_R1105_U125 | ~new_P1_R1105_U20 | ~new_P1_R1105_U238 | ~new_P1_R1105_U237;
  assign new_P1_R1105_U127 = ~new_P1_R1105_U111 | ~new_P1_R1105_U20;
  assign new_P1_R1105_U128 = ~P1_REG2_REG_7_ | ~new_P1_U3472;
  assign new_P1_R1105_U129 = ~new_P1_R1105_U127 | ~new_P1_R1105_U128 | ~new_P1_R1105_U6;
  assign new_P1_R1105_U130 = new_P1_U3469 | P1_REG2_REG_6_;
  assign new_P1_R1105_U131 = ~new_P1_R1105_U101 | ~new_P1_R1105_U97;
  assign new_P1_R1105_U132 = ~new_P1_U3457 | ~P1_REG2_REG_2_;
  assign new_P1_R1105_U133 = ~new_P1_R1105_U43;
  assign new_P1_R1105_U134 = ~new_P1_R1105_U100 | ~new_P1_R1105_U5;
  assign new_P1_R1105_U135 = ~new_P1_R1105_U43 | ~new_P1_R1105_U96;
  assign new_P1_R1105_U136 = ~new_P1_U3460 | ~P1_REG2_REG_3_;
  assign new_P1_R1105_U137 = ~new_P1_R1105_U42;
  assign new_P1_R1105_U138 = P1_REG2_REG_4_ | new_P1_U3463;
  assign new_P1_R1105_U139 = ~new_P1_R1105_U138 | ~new_P1_R1105_U42;
  assign new_P1_R1105_U140 = ~new_P1_R1105_U139 | ~new_P1_R1105_U32 | ~new_P1_R1105_U245 | ~new_P1_R1105_U244;
  assign new_P1_R1105_U141 = ~new_P1_R1105_U137 | ~new_P1_R1105_U32;
  assign new_P1_R1105_U142 = ~P1_REG2_REG_5_ | ~new_P1_U3466;
  assign new_P1_R1105_U143 = ~new_P1_R1105_U141 | ~new_P1_R1105_U142 | ~new_P1_R1105_U4;
  assign new_P1_R1105_U144 = new_P1_U3463 | P1_REG2_REG_4_;
  assign new_P1_R1105_U145 = ~new_P1_R1105_U100 | ~new_P1_R1105_U97;
  assign new_P1_R1105_U146 = ~new_P1_R1105_U82;
  assign new_P1_R1105_U147 = ~new_P1_U3460 | ~P1_REG2_REG_3_;
  assign new_P1_R1105_U148 = ~new_P1_R1105_U256 | ~new_P1_R1105_U257 | ~new_P1_R1105_U41 | ~new_P1_R1105_U40;
  assign new_P1_R1105_U149 = ~new_P1_R1105_U41 | ~new_P1_R1105_U40;
  assign new_P1_R1105_U150 = ~new_P1_U3457 | ~P1_REG2_REG_2_;
  assign new_P1_R1105_U151 = ~new_P1_R1105_U149 | ~new_P1_R1105_U150 | ~new_P1_R1105_U97;
  assign new_P1_R1105_U152 = P1_REG2_REG_1_ | new_P1_U3454;
  assign new_P1_R1105_U153 = ~new_P1_R1105_U83;
  assign new_P1_R1105_U154 = new_P1_U3478 | P1_REG2_REG_9_;
  assign new_P1_R1105_U155 = new_P1_U3481 | P1_REG2_REG_10_;
  assign new_P1_R1105_U156 = ~new_P1_R1105_U93 | ~new_P1_R1105_U7;
  assign new_P1_R1105_U157 = ~new_P1_U3481 | ~P1_REG2_REG_10_;
  assign new_P1_R1105_U158 = ~new_P1_R1105_U156 | ~new_P1_R1105_U157 | ~new_P1_R1105_U90;
  assign new_P1_R1105_U159 = P1_REG2_REG_10_ | new_P1_U3481;
  assign new_P1_R1105_U160 = ~new_P1_R1105_U81 | ~new_P1_R1105_U120 | ~new_P1_R1105_U7;
  assign new_P1_R1105_U161 = ~new_P1_R1105_U159 | ~new_P1_R1105_U158;
  assign new_P1_R1105_U162 = ~new_P1_R1105_U88;
  assign new_P1_R1105_U163 = new_P1_U3490 | P1_REG2_REG_13_;
  assign new_P1_R1105_U164 = new_P1_U3487 | P1_REG2_REG_12_;
  assign new_P1_R1105_U165 = ~new_P1_R1105_U92 | ~new_P1_R1105_U8;
  assign new_P1_R1105_U166 = ~new_P1_U3490 | ~P1_REG2_REG_13_;
  assign new_P1_R1105_U167 = ~new_P1_R1105_U165 | ~new_P1_R1105_U166 | ~new_P1_R1105_U91;
  assign new_P1_R1105_U168 = P1_REG2_REG_11_ | new_P1_U3484;
  assign new_P1_R1105_U169 = P1_REG2_REG_13_ | new_P1_U3490;
  assign new_P1_R1105_U170 = ~new_P1_R1105_U88 | ~new_P1_R1105_U168 | ~new_P1_R1105_U8;
  assign new_P1_R1105_U171 = ~new_P1_R1105_U169 | ~new_P1_R1105_U167;
  assign new_P1_R1105_U172 = ~new_P1_R1105_U87;
  assign new_P1_R1105_U173 = P1_REG2_REG_14_ | new_P1_U3493;
  assign new_P1_R1105_U174 = ~new_P1_R1105_U173 | ~new_P1_R1105_U87;
  assign new_P1_R1105_U175 = ~new_P1_U3493 | ~P1_REG2_REG_14_;
  assign new_P1_R1105_U176 = ~new_P1_R1105_U86;
  assign new_P1_R1105_U177 = P1_REG2_REG_15_ | new_P1_U3496;
  assign new_P1_R1105_U178 = ~new_P1_R1105_U177 | ~new_P1_R1105_U86;
  assign new_P1_R1105_U179 = ~new_P1_U3496 | ~P1_REG2_REG_15_;
  assign new_P1_R1105_U180 = ~new_P1_R1105_U66;
  assign new_P1_R1105_U181 = new_P1_U3502 | P1_REG2_REG_17_;
  assign new_P1_R1105_U182 = new_P1_U3499 | P1_REG2_REG_16_;
  assign new_P1_R1105_U183 = ~new_P1_R1105_U47;
  assign new_P1_R1105_U184 = ~new_P1_R1105_U48 | ~new_P1_R1105_U47;
  assign new_P1_R1105_U185 = ~new_P1_U3502 | ~new_P1_R1105_U184;
  assign new_P1_R1105_U186 = ~P1_REG2_REG_17_ | ~new_P1_R1105_U183;
  assign new_P1_R1105_U187 = ~new_P1_R1105_U9 | ~new_P1_R1105_U66;
  assign new_P1_R1105_U188 = ~new_P1_R1105_U65;
  assign new_P1_R1105_U189 = P1_REG2_REG_18_ | new_P1_U3505;
  assign new_P1_R1105_U190 = ~new_P1_R1105_U189 | ~new_P1_R1105_U65;
  assign new_P1_R1105_U191 = ~new_P1_U3505 | ~P1_REG2_REG_18_;
  assign new_P1_R1105_U192 = ~new_P1_R1105_U190 | ~new_P1_R1105_U191 | ~new_P1_R1105_U261 | ~new_P1_R1105_U260;
  assign new_P1_R1105_U193 = ~new_P1_U3505 | ~P1_REG2_REG_18_;
  assign new_P1_R1105_U194 = ~new_P1_R1105_U188 | ~new_P1_R1105_U193;
  assign new_P1_R1105_U195 = new_P1_U3505 | P1_REG2_REG_18_;
  assign new_P1_R1105_U196 = ~new_P1_R1105_U194 | ~new_P1_R1105_U195 | ~new_P1_R1105_U264;
  assign new_P1_R1105_U197 = P1_REG2_REG_16_ | new_P1_U3499;
  assign new_P1_R1105_U198 = ~new_P1_R1105_U197 | ~new_P1_R1105_U66;
  assign new_P1_R1105_U199 = ~new_P1_R1105_U198 | ~new_P1_R1105_U47 | ~new_P1_R1105_U273 | ~new_P1_R1105_U272;
  assign new_P1_R1105_U200 = ~new_P1_R1105_U180 | ~new_P1_R1105_U47;
  assign new_P1_R1105_U201 = ~P1_REG2_REG_17_ | ~new_P1_U3502;
  assign new_P1_R1105_U202 = ~new_P1_R1105_U200 | ~new_P1_R1105_U201 | ~new_P1_R1105_U9;
  assign new_P1_R1105_U203 = new_P1_U3499 | P1_REG2_REG_16_;
  assign new_P1_R1105_U204 = ~new_P1_R1105_U168 | ~new_P1_R1105_U88;
  assign new_P1_R1105_U205 = ~new_P1_R1105_U67;
  assign new_P1_R1105_U206 = P1_REG2_REG_12_ | new_P1_U3487;
  assign new_P1_R1105_U207 = ~new_P1_R1105_U206 | ~new_P1_R1105_U67;
  assign new_P1_R1105_U208 = ~new_P1_R1105_U207 | ~new_P1_R1105_U91 | ~new_P1_R1105_U294 | ~new_P1_R1105_U293;
  assign new_P1_R1105_U209 = ~new_P1_R1105_U205 | ~new_P1_R1105_U91;
  assign new_P1_R1105_U210 = ~new_P1_U3490 | ~P1_REG2_REG_13_;
  assign new_P1_R1105_U211 = ~new_P1_R1105_U209 | ~new_P1_R1105_U210 | ~new_P1_R1105_U8;
  assign new_P1_R1105_U212 = new_P1_U3487 | P1_REG2_REG_12_;
  assign new_P1_R1105_U213 = P1_REG2_REG_9_ | new_P1_U3478;
  assign new_P1_R1105_U214 = ~new_P1_R1105_U213 | ~new_P1_R1105_U38;
  assign new_P1_R1105_U215 = ~new_P1_R1105_U214 | ~new_P1_R1105_U90 | ~new_P1_R1105_U306 | ~new_P1_R1105_U305;
  assign new_P1_R1105_U216 = ~new_P1_R1105_U122 | ~new_P1_R1105_U90;
  assign new_P1_R1105_U217 = ~new_P1_U3481 | ~P1_REG2_REG_10_;
  assign new_P1_R1105_U218 = ~new_P1_R1105_U216 | ~new_P1_R1105_U217 | ~new_P1_R1105_U7;
  assign new_P1_R1105_U219 = ~new_P1_R1105_U123 | ~new_P1_R1105_U90;
  assign new_P1_R1105_U220 = ~new_P1_R1105_U120 | ~new_P1_R1105_U49;
  assign new_P1_R1105_U221 = ~new_P1_R1105_U130 | ~new_P1_R1105_U20;
  assign new_P1_R1105_U222 = ~new_P1_R1105_U144 | ~new_P1_R1105_U32;
  assign new_P1_R1105_U223 = ~new_P1_R1105_U147 | ~new_P1_R1105_U96;
  assign new_P1_R1105_U224 = ~new_P1_R1105_U203 | ~new_P1_R1105_U47;
  assign new_P1_R1105_U225 = ~new_P1_R1105_U212 | ~new_P1_R1105_U91;
  assign new_P1_R1105_U226 = ~new_P1_R1105_U168 | ~new_P1_R1105_U56;
  assign new_P1_R1105_U227 = ~new_P1_U3478 | ~new_P1_R1105_U37;
  assign new_P1_R1105_U228 = ~P1_REG2_REG_9_ | ~new_P1_R1105_U36;
  assign new_P1_R1105_U229 = ~new_P1_R1105_U228 | ~new_P1_R1105_U227;
  assign new_P1_R1105_U230 = ~new_P1_R1105_U219 | ~new_P1_R1105_U38;
  assign new_P1_R1105_U231 = ~new_P1_R1105_U229 | ~new_P1_R1105_U122;
  assign new_P1_R1105_U232 = ~new_P1_U3475 | ~new_P1_R1105_U34;
  assign new_P1_R1105_U233 = ~P1_REG2_REG_8_ | ~new_P1_R1105_U35;
  assign new_P1_R1105_U234 = ~new_P1_R1105_U233 | ~new_P1_R1105_U232;
  assign new_P1_R1105_U235 = ~new_P1_R1105_U220 | ~new_P1_R1105_U81;
  assign new_P1_R1105_U236 = ~new_P1_R1105_U119 | ~new_P1_R1105_U234;
  assign new_P1_R1105_U237 = ~new_P1_U3472 | ~new_P1_R1105_U21;
  assign new_P1_R1105_U238 = ~P1_REG2_REG_7_ | ~new_P1_R1105_U19;
  assign new_P1_R1105_U239 = ~new_P1_U3469 | ~new_P1_R1105_U17;
  assign new_P1_R1105_U240 = ~P1_REG2_REG_6_ | ~new_P1_R1105_U18;
  assign new_P1_R1105_U241 = ~new_P1_R1105_U240 | ~new_P1_R1105_U239;
  assign new_P1_R1105_U242 = ~new_P1_R1105_U221 | ~new_P1_R1105_U39;
  assign new_P1_R1105_U243 = ~new_P1_R1105_U241 | ~new_P1_R1105_U111;
  assign new_P1_R1105_U244 = ~new_P1_U3466 | ~new_P1_R1105_U33;
  assign new_P1_R1105_U245 = ~P1_REG2_REG_5_ | ~new_P1_R1105_U24;
  assign new_P1_R1105_U246 = ~new_P1_U3463 | ~new_P1_R1105_U22;
  assign new_P1_R1105_U247 = ~P1_REG2_REG_4_ | ~new_P1_R1105_U23;
  assign new_P1_R1105_U248 = ~new_P1_R1105_U247 | ~new_P1_R1105_U246;
  assign new_P1_R1105_U249 = ~new_P1_R1105_U222 | ~new_P1_R1105_U42;
  assign new_P1_R1105_U250 = ~new_P1_R1105_U248 | ~new_P1_R1105_U137;
  assign new_P1_R1105_U251 = ~new_P1_U3460 | ~new_P1_R1105_U30;
  assign new_P1_R1105_U252 = ~P1_REG2_REG_3_ | ~new_P1_R1105_U31;
  assign new_P1_R1105_U253 = ~new_P1_R1105_U252 | ~new_P1_R1105_U251;
  assign new_P1_R1105_U254 = ~new_P1_R1105_U223 | ~new_P1_R1105_U82;
  assign new_P1_R1105_U255 = ~new_P1_R1105_U146 | ~new_P1_R1105_U253;
  assign new_P1_R1105_U256 = ~new_P1_U3457 | ~new_P1_R1105_U25;
  assign new_P1_R1105_U257 = ~P1_REG2_REG_2_ | ~new_P1_R1105_U26;
  assign new_P1_R1105_U258 = ~new_P1_R1105_U98 | ~new_P1_R1105_U83;
  assign new_P1_R1105_U259 = ~new_P1_R1105_U153 | ~new_P1_R1105_U29;
  assign new_P1_R1105_U260 = ~new_P1_U3442 | ~new_P1_R1105_U85;
  assign new_P1_R1105_U261 = ~P1_REG2_REG_19_ | ~new_P1_R1105_U84;
  assign new_P1_R1105_U262 = ~new_P1_U3442 | ~new_P1_R1105_U85;
  assign new_P1_R1105_U263 = ~P1_REG2_REG_19_ | ~new_P1_R1105_U84;
  assign new_P1_R1105_U264 = ~new_P1_R1105_U263 | ~new_P1_R1105_U262;
  assign new_P1_R1105_U265 = ~new_P1_U3505 | ~new_P1_R1105_U63;
  assign new_P1_R1105_U266 = ~P1_REG2_REG_18_ | ~new_P1_R1105_U64;
  assign new_P1_R1105_U267 = ~new_P1_U3505 | ~new_P1_R1105_U63;
  assign new_P1_R1105_U268 = ~P1_REG2_REG_18_ | ~new_P1_R1105_U64;
  assign new_P1_R1105_U269 = ~new_P1_R1105_U268 | ~new_P1_R1105_U267;
  assign new_P1_R1105_U270 = ~new_P1_R1105_U65 | ~new_P1_R1105_U266 | ~new_P1_R1105_U265;
  assign new_P1_R1105_U271 = ~new_P1_R1105_U269 | ~new_P1_R1105_U188;
  assign new_P1_R1105_U272 = ~new_P1_U3502 | ~new_P1_R1105_U48;
  assign new_P1_R1105_U273 = ~P1_REG2_REG_17_ | ~new_P1_R1105_U46;
  assign new_P1_R1105_U274 = ~new_P1_U3499 | ~new_P1_R1105_U44;
  assign new_P1_R1105_U275 = ~P1_REG2_REG_16_ | ~new_P1_R1105_U45;
  assign new_P1_R1105_U276 = ~new_P1_R1105_U275 | ~new_P1_R1105_U274;
  assign new_P1_R1105_U277 = ~new_P1_R1105_U224 | ~new_P1_R1105_U66;
  assign new_P1_R1105_U278 = ~new_P1_R1105_U276 | ~new_P1_R1105_U180;
  assign new_P1_R1105_U279 = ~new_P1_U3496 | ~new_P1_R1105_U61;
  assign new_P1_R1105_U280 = ~P1_REG2_REG_15_ | ~new_P1_R1105_U62;
  assign new_P1_R1105_U281 = ~new_P1_U3496 | ~new_P1_R1105_U61;
  assign new_P1_R1105_U282 = ~P1_REG2_REG_15_ | ~new_P1_R1105_U62;
  assign new_P1_R1105_U283 = ~new_P1_R1105_U282 | ~new_P1_R1105_U281;
  assign new_P1_R1105_U284 = ~new_P1_R1105_U86 | ~new_P1_R1105_U280 | ~new_P1_R1105_U279;
  assign new_P1_R1105_U285 = ~new_P1_R1105_U176 | ~new_P1_R1105_U283;
  assign new_P1_R1105_U286 = ~new_P1_U3493 | ~new_P1_R1105_U59;
  assign new_P1_R1105_U287 = ~P1_REG2_REG_14_ | ~new_P1_R1105_U60;
  assign new_P1_R1105_U288 = ~new_P1_U3493 | ~new_P1_R1105_U59;
  assign new_P1_R1105_U289 = ~P1_REG2_REG_14_ | ~new_P1_R1105_U60;
  assign new_P1_R1105_U290 = ~new_P1_R1105_U289 | ~new_P1_R1105_U288;
  assign new_P1_R1105_U291 = ~new_P1_R1105_U87 | ~new_P1_R1105_U287 | ~new_P1_R1105_U286;
  assign new_P1_R1105_U292 = ~new_P1_R1105_U172 | ~new_P1_R1105_U290;
  assign new_P1_R1105_U293 = ~new_P1_U3490 | ~new_P1_R1105_U57;
  assign new_P1_R1105_U294 = ~P1_REG2_REG_13_ | ~new_P1_R1105_U58;
  assign new_P1_R1105_U295 = ~new_P1_U3487 | ~new_P1_R1105_U52;
  assign new_P1_R1105_U296 = ~P1_REG2_REG_12_ | ~new_P1_R1105_U53;
  assign new_P1_R1105_U297 = ~new_P1_R1105_U296 | ~new_P1_R1105_U295;
  assign new_P1_R1105_U298 = ~new_P1_R1105_U225 | ~new_P1_R1105_U67;
  assign new_P1_R1105_U299 = ~new_P1_R1105_U297 | ~new_P1_R1105_U205;
  assign new_P1_R1105_U300 = ~new_P1_U3484 | ~new_P1_R1105_U54;
  assign new_P1_R1105_U301 = ~P1_REG2_REG_11_ | ~new_P1_R1105_U55;
  assign new_P1_R1105_U302 = ~new_P1_R1105_U301 | ~new_P1_R1105_U300;
  assign new_P1_R1105_U303 = ~new_P1_R1105_U226 | ~new_P1_R1105_U88;
  assign new_P1_R1105_U304 = ~new_P1_R1105_U162 | ~new_P1_R1105_U302;
  assign new_P1_R1105_U305 = ~new_P1_U3481 | ~new_P1_R1105_U50;
  assign new_P1_R1105_U306 = ~P1_REG2_REG_10_ | ~new_P1_R1105_U51;
  assign new_P1_R1105_U307 = ~new_P1_U3448 | ~new_P1_R1105_U27;
  assign new_P1_R1105_U308 = ~P1_REG2_REG_0_ | ~new_P1_R1105_U28;
  assign new_P1_SUB_84_U6 = new_P1_SUB_84_U227 & new_P1_SUB_84_U38;
  assign new_P1_SUB_84_U7 = new_P1_SUB_84_U225 & new_P1_SUB_84_U192;
  assign new_P1_SUB_84_U8 = new_P1_SUB_84_U224 & new_P1_SUB_84_U35;
  assign new_P1_SUB_84_U9 = new_P1_SUB_84_U223 & new_P1_SUB_84_U36;
  assign new_P1_SUB_84_U10 = new_P1_SUB_84_U221 & new_P1_SUB_84_U195;
  assign new_P1_SUB_84_U11 = new_P1_SUB_84_U220 & new_P1_SUB_84_U34;
  assign new_P1_SUB_84_U12 = new_P1_SUB_84_U219 & new_P1_SUB_84_U197;
  assign new_P1_SUB_84_U13 = new_P1_SUB_84_U217 & new_P1_SUB_84_U198;
  assign new_P1_SUB_84_U14 = new_P1_SUB_84_U216 & new_P1_SUB_84_U172;
  assign new_P1_SUB_84_U15 = new_P1_SUB_84_U215 & new_P1_SUB_84_U200;
  assign new_P1_SUB_84_U16 = new_P1_SUB_84_U213 & new_P1_SUB_84_U201;
  assign new_P1_SUB_84_U17 = new_P1_SUB_84_U212 & new_P1_SUB_84_U169;
  assign new_P1_SUB_84_U18 = new_P1_SUB_84_U211 & new_P1_SUB_84_U167;
  assign new_P1_SUB_84_U19 = new_P1_SUB_84_U209 & new_P1_SUB_84_U204;
  assign new_P1_SUB_84_U20 = new_P1_SUB_84_U208 & new_P1_SUB_84_U33;
  assign new_P1_SUB_84_U21 = new_P1_SUB_84_U207 & new_P1_SUB_84_U27;
  assign new_P1_SUB_84_U22 = new_P1_SUB_84_U190 & new_P1_SUB_84_U180;
  assign new_P1_SUB_84_U23 = new_P1_SUB_84_U189 & new_P1_SUB_84_U29;
  assign new_P1_SUB_84_U24 = new_P1_SUB_84_U188 & new_P1_SUB_84_U30;
  assign new_P1_SUB_84_U25 = new_P1_SUB_84_U186 & new_P1_SUB_84_U183;
  assign new_P1_SUB_84_U26 = new_P1_SUB_84_U185 & new_P1_SUB_84_U28;
  assign new_P1_SUB_84_U27 = P1_IR_REG_2_ | P1_IR_REG_1_ | P1_IR_REG_0_;
  assign new_P1_SUB_84_U28 = ~new_P1_SUB_84_U43 | ~new_P1_SUB_84_U44 | ~new_P1_SUB_84_U230;
  assign new_P1_SUB_84_U29 = ~new_P1_SUB_84_U45 | ~new_P1_SUB_84_U230;
  assign new_P1_SUB_84_U30 = ~new_P1_SUB_84_U46 | ~new_P1_SUB_84_U181;
  assign new_P1_SUB_84_U31 = ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U32 = ~P1_IR_REG_3_;
  assign new_P1_SUB_84_U33 = ~new_P1_SUB_84_U56 | ~new_P1_SUB_84_U51;
  assign new_P1_SUB_84_U34 = ~new_P1_SUB_84_U127 | ~new_P1_SUB_84_U128 | ~new_P1_SUB_84_U130 | ~new_P1_SUB_84_U129;
  assign new_P1_SUB_84_U35 = ~new_P1_SUB_84_U156 | ~new_P1_SUB_84_U184;
  assign new_P1_SUB_84_U36 = ~new_P1_SUB_84_U157 | ~new_P1_SUB_84_U193;
  assign new_P1_SUB_84_U37 = ~P1_IR_REG_15_;
  assign new_P1_SUB_84_U38 = ~new_P1_SUB_84_U158 | ~new_P1_SUB_84_U184;
  assign new_P1_SUB_84_U39 = ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U40 = ~new_P1_SUB_84_U247 | ~new_P1_SUB_84_U246;
  assign new_P1_SUB_84_U41 = ~new_P1_SUB_84_U237 | ~new_P1_SUB_84_U236;
  assign new_P1_SUB_84_U42 = ~new_P1_SUB_84_U241 | ~new_P1_SUB_84_U240;
  assign new_P1_SUB_84_U43 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U44 = ~P1_IR_REG_7_ & ~P1_IR_REG_8_;
  assign new_P1_SUB_84_U45 = ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U46 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_;
  assign new_P1_SUB_84_U47 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U48 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_ & ~P1_IR_REG_15_;
  assign new_P1_SUB_84_U49 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_84_U50 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_84_U51 = new_P1_SUB_84_U47 & new_P1_SUB_84_U48 & new_P1_SUB_84_U50 & new_P1_SUB_84_U49;
  assign new_P1_SUB_84_U52 = ~P1_IR_REG_26_ & ~P1_IR_REG_25_ & ~P1_IR_REG_23_ & ~P1_IR_REG_24_;
  assign new_P1_SUB_84_U53 = ~P1_IR_REG_2_ & ~P1_IR_REG_29_ & ~P1_IR_REG_27_ & ~P1_IR_REG_28_;
  assign new_P1_SUB_84_U54 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U55 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U56 = new_P1_SUB_84_U52 & new_P1_SUB_84_U53 & new_P1_SUB_84_U55 & new_P1_SUB_84_U54;
  assign new_P1_SUB_84_U57 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U58 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_ & ~P1_IR_REG_15_;
  assign new_P1_SUB_84_U59 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_84_U60 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_84_U61 = new_P1_SUB_84_U57 & new_P1_SUB_84_U58 & new_P1_SUB_84_U60 & new_P1_SUB_84_U59;
  assign new_P1_SUB_84_U62 = ~P1_IR_REG_26_ & ~P1_IR_REG_25_ & ~P1_IR_REG_23_ & ~P1_IR_REG_24_;
  assign new_P1_SUB_84_U63 = ~P1_IR_REG_28_ & ~P1_IR_REG_2_ & ~P1_IR_REG_27_;
  assign new_P1_SUB_84_U64 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U65 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U66 = new_P1_SUB_84_U62 & new_P1_SUB_84_U63 & new_P1_SUB_84_U65 & new_P1_SUB_84_U64;
  assign new_P1_SUB_84_U67 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U68 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U69 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_84_U70 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_84_U71 = new_P1_SUB_84_U67 & new_P1_SUB_84_U68 & new_P1_SUB_84_U70 & new_P1_SUB_84_U69;
  assign new_P1_SUB_84_U72 = ~P1_IR_REG_25_ & ~P1_IR_REG_24_ & ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_84_U73 = ~P1_IR_REG_27_ & ~P1_IR_REG_2_ & ~P1_IR_REG_26_;
  assign new_P1_SUB_84_U74 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U75 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U76 = new_P1_SUB_84_U72 & new_P1_SUB_84_U73 & new_P1_SUB_84_U75 & new_P1_SUB_84_U74;
  assign new_P1_SUB_84_U77 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U78 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U79 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_84_U80 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_84_U81 = new_P1_SUB_84_U77 & new_P1_SUB_84_U78 & new_P1_SUB_84_U80 & new_P1_SUB_84_U79;
  assign new_P1_SUB_84_U82 = ~P1_IR_REG_25_ & ~P1_IR_REG_24_ & ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_84_U83 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_26_;
  assign new_P1_SUB_84_U84 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U85 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U86 = new_P1_SUB_84_U82 & new_P1_SUB_84_U83 & new_P1_SUB_84_U85 & new_P1_SUB_84_U84;
  assign new_P1_SUB_84_U87 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U88 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U89 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_84_U90 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_84_U91 = new_P1_SUB_84_U87 & new_P1_SUB_84_U88 & new_P1_SUB_84_U90 & new_P1_SUB_84_U89;
  assign new_P1_SUB_84_U92 = ~P1_IR_REG_25_ & ~P1_IR_REG_24_ & ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_84_U93 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_26_;
  assign new_P1_SUB_84_U94 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U95 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U96 = new_P1_SUB_84_U92 & new_P1_SUB_84_U93 & new_P1_SUB_84_U95 & new_P1_SUB_84_U94;
  assign new_P1_SUB_84_U97 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U98 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U99 = ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_;
  assign new_P1_SUB_84_U100 = ~P1_IR_REG_0_ & ~P1_IR_REG_20_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_84_U101 = new_P1_SUB_84_U97 & new_P1_SUB_84_U98 & new_P1_SUB_84_U100 & new_P1_SUB_84_U99;
  assign new_P1_SUB_84_U102 = ~P1_IR_REG_24_ & ~P1_IR_REG_23_ & ~P1_IR_REG_21_ & ~P1_IR_REG_22_;
  assign new_P1_SUB_84_U103 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_25_;
  assign new_P1_SUB_84_U104 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U105 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U106 = new_P1_SUB_84_U102 & new_P1_SUB_84_U103 & new_P1_SUB_84_U105 & new_P1_SUB_84_U104;
  assign new_P1_SUB_84_U107 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U108 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U109 = ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_;
  assign new_P1_SUB_84_U110 = ~P1_IR_REG_0_ & ~P1_IR_REG_20_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_84_U111 = new_P1_SUB_84_U107 & new_P1_SUB_84_U108 & new_P1_SUB_84_U110 & new_P1_SUB_84_U109;
  assign new_P1_SUB_84_U112 = ~P1_IR_REG_22_ & ~P1_IR_REG_23_ & ~P1_IR_REG_21_;
  assign new_P1_SUB_84_U113 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_24_;
  assign new_P1_SUB_84_U114 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U115 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U116 = new_P1_SUB_84_U112 & new_P1_SUB_84_U113 & new_P1_SUB_84_U115 & new_P1_SUB_84_U114;
  assign new_P1_SUB_84_U117 = ~P1_IR_REG_11_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_;
  assign new_P1_SUB_84_U118 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_ & ~P1_IR_REG_13_;
  assign new_P1_SUB_84_U119 = ~P1_IR_REG_17_ & ~P1_IR_REG_18_ & ~P1_IR_REG_16_;
  assign new_P1_SUB_84_U120 = ~P1_IR_REG_1_ & ~P1_IR_REG_0_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_84_U121 = new_P1_SUB_84_U117 & new_P1_SUB_84_U118 & new_P1_SUB_84_U120 & new_P1_SUB_84_U119;
  assign new_P1_SUB_84_U122 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_84_U123 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_84_U124 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U125 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U126 = new_P1_SUB_84_U122 & new_P1_SUB_84_U123 & new_P1_SUB_84_U125 & new_P1_SUB_84_U124;
  assign new_P1_SUB_84_U127 = ~P1_IR_REG_11_ & ~P1_IR_REG_10_ & ~P1_IR_REG_12_ & ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U128 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_15_ & ~P1_IR_REG_16_;
  assign new_P1_SUB_84_U129 = ~P1_IR_REG_5_ & ~P1_IR_REG_4_ & ~P1_IR_REG_2_ & ~P1_IR_REG_3_;
  assign new_P1_SUB_84_U130 = ~P1_IR_REG_9_ & ~P1_IR_REG_8_ & ~P1_IR_REG_6_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U131 = ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_84_U132 = ~P1_IR_REG_19_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_84_U133 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_;
  assign new_P1_SUB_84_U134 = new_P1_SUB_84_U133 & new_P1_SUB_84_U132 & new_P1_SUB_84_U131;
  assign new_P1_SUB_84_U135 = ~P1_IR_REG_11_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_;
  assign new_P1_SUB_84_U136 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_ & ~P1_IR_REG_13_;
  assign new_P1_SUB_84_U137 = new_P1_SUB_84_U136 & new_P1_SUB_84_U135;
  assign new_P1_SUB_84_U138 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_84_U139 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_84_U140 = ~P1_IR_REG_3_ & ~P1_IR_REG_4_ & ~P1_IR_REG_2_;
  assign new_P1_SUB_84_U141 = new_P1_SUB_84_U140 & new_P1_SUB_84_U139;
  assign new_P1_SUB_84_U142 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_7_ & ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_84_U143 = ~P1_IR_REG_11_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_;
  assign new_P1_SUB_84_U144 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_ & ~P1_IR_REG_13_;
  assign new_P1_SUB_84_U145 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_84_U146 = ~P1_IR_REG_20_ & ~P1_IR_REG_0_ & ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U147 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_7_ & ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_84_U148 = ~P1_IR_REG_11_ & ~P1_IR_REG_10_ & ~P1_IR_REG_12_ & ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U149 = ~P1_IR_REG_16_ & ~P1_IR_REG_15_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_84_U150 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_84_U151 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_7_ & ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_84_U152 = ~P1_IR_REG_11_ & ~P1_IR_REG_10_ & ~P1_IR_REG_12_ & ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U153 = ~P1_IR_REG_16_ & ~P1_IR_REG_15_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_84_U154 = ~P1_IR_REG_2_ & ~P1_IR_REG_0_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_ & ~P1_IR_REG_5_;
  assign new_P1_SUB_84_U155 = ~P1_IR_REG_9_ & ~P1_IR_REG_8_ & ~P1_IR_REG_6_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_84_U156 = ~P1_IR_REG_9_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_84_U157 = ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_84_U158 = ~P1_IR_REG_10_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_84_U159 = ~P1_IR_REG_9_;
  assign new_P1_SUB_84_U160 = new_P1_SUB_84_U233 & new_P1_SUB_84_U232;
  assign new_P1_SUB_84_U161 = ~P1_IR_REG_5_;
  assign new_P1_SUB_84_U162 = new_P1_SUB_84_U235 & new_P1_SUB_84_U234;
  assign new_P1_SUB_84_U163 = ~P1_IR_REG_31_;
  assign new_P1_SUB_84_U164 = ~P1_IR_REG_30_;
  assign new_P1_SUB_84_U165 = new_P1_SUB_84_U239 & new_P1_SUB_84_U238;
  assign new_P1_SUB_84_U166 = ~P1_IR_REG_27_;
  assign new_P1_SUB_84_U167 = ~new_P1_SUB_84_U96 | ~new_P1_SUB_84_U91;
  assign new_P1_SUB_84_U168 = ~P1_IR_REG_25_;
  assign new_P1_SUB_84_U169 = ~new_P1_SUB_84_U116 | ~new_P1_SUB_84_U111;
  assign new_P1_SUB_84_U170 = new_P1_SUB_84_U243 & new_P1_SUB_84_U242;
  assign new_P1_SUB_84_U171 = ~P1_IR_REG_21_;
  assign new_P1_SUB_84_U172 = ~new_P1_SUB_84_U146 | ~new_P1_SUB_84_U147 | ~new_P1_SUB_84_U145 | ~new_P1_SUB_84_U144 | ~new_P1_SUB_84_U143;
  assign new_P1_SUB_84_U173 = new_P1_SUB_84_U245 & new_P1_SUB_84_U244;
  assign new_P1_SUB_84_U174 = ~P1_IR_REG_1_;
  assign new_P1_SUB_84_U175 = ~P1_IR_REG_0_;
  assign new_P1_SUB_84_U176 = ~P1_IR_REG_17_;
  assign new_P1_SUB_84_U177 = new_P1_SUB_84_U249 & new_P1_SUB_84_U248;
  assign new_P1_SUB_84_U178 = ~P1_IR_REG_13_;
  assign new_P1_SUB_84_U179 = new_P1_SUB_84_U251 & new_P1_SUB_84_U250;
  assign new_P1_SUB_84_U180 = ~new_P1_SUB_84_U230 | ~new_P1_SUB_84_U32;
  assign new_P1_SUB_84_U181 = ~new_P1_SUB_84_U29;
  assign new_P1_SUB_84_U182 = ~new_P1_SUB_84_U30;
  assign new_P1_SUB_84_U183 = ~new_P1_SUB_84_U182 | ~new_P1_SUB_84_U31;
  assign new_P1_SUB_84_U184 = ~new_P1_SUB_84_U28;
  assign new_P1_SUB_84_U185 = ~P1_IR_REG_8_ | ~new_P1_SUB_84_U183;
  assign new_P1_SUB_84_U186 = ~P1_IR_REG_7_ | ~new_P1_SUB_84_U30;
  assign new_P1_SUB_84_U187 = ~new_P1_SUB_84_U181 | ~new_P1_SUB_84_U161;
  assign new_P1_SUB_84_U188 = ~P1_IR_REG_6_ | ~new_P1_SUB_84_U187;
  assign new_P1_SUB_84_U189 = ~P1_IR_REG_4_ | ~new_P1_SUB_84_U180;
  assign new_P1_SUB_84_U190 = ~P1_IR_REG_3_ | ~new_P1_SUB_84_U27;
  assign new_P1_SUB_84_U191 = ~new_P1_SUB_84_U38;
  assign new_P1_SUB_84_U192 = ~new_P1_SUB_84_U191 | ~new_P1_SUB_84_U39;
  assign new_P1_SUB_84_U193 = ~new_P1_SUB_84_U35;
  assign new_P1_SUB_84_U194 = ~new_P1_SUB_84_U36;
  assign new_P1_SUB_84_U195 = ~new_P1_SUB_84_U194 | ~new_P1_SUB_84_U37;
  assign new_P1_SUB_84_U196 = ~new_P1_SUB_84_U34;
  assign new_P1_SUB_84_U197 = ~new_P1_SUB_84_U152 | ~new_P1_SUB_84_U153 | ~new_P1_SUB_84_U155 | ~new_P1_SUB_84_U154;
  assign new_P1_SUB_84_U198 = ~new_P1_SUB_84_U148 | ~new_P1_SUB_84_U149 | ~new_P1_SUB_84_U151 | ~new_P1_SUB_84_U150;
  assign new_P1_SUB_84_U199 = ~new_P1_SUB_84_U172;
  assign new_P1_SUB_84_U200 = ~new_P1_SUB_84_U134 | ~new_P1_SUB_84_U196;
  assign new_P1_SUB_84_U201 = ~new_P1_SUB_84_U126 | ~new_P1_SUB_84_U121;
  assign new_P1_SUB_84_U202 = ~new_P1_SUB_84_U169;
  assign new_P1_SUB_84_U203 = ~new_P1_SUB_84_U167;
  assign new_P1_SUB_84_U204 = ~new_P1_SUB_84_U66 | ~new_P1_SUB_84_U61;
  assign new_P1_SUB_84_U205 = ~new_P1_SUB_84_U33;
  assign new_P1_SUB_84_U206 = P1_IR_REG_1_ | P1_IR_REG_0_;
  assign new_P1_SUB_84_U207 = ~P1_IR_REG_2_ | ~new_P1_SUB_84_U206;
  assign new_P1_SUB_84_U208 = ~P1_IR_REG_29_ | ~new_P1_SUB_84_U204;
  assign new_P1_SUB_84_U209 = ~P1_IR_REG_28_ | ~new_P1_SUB_84_U229;
  assign new_P1_SUB_84_U210 = ~new_P1_SUB_84_U106 | ~new_P1_SUB_84_U101;
  assign new_P1_SUB_84_U211 = ~P1_IR_REG_26_ | ~new_P1_SUB_84_U210;
  assign new_P1_SUB_84_U212 = ~P1_IR_REG_24_ | ~new_P1_SUB_84_U201;
  assign new_P1_SUB_84_U213 = ~P1_IR_REG_23_ | ~new_P1_SUB_84_U200;
  assign new_P1_SUB_84_U214 = ~new_P1_SUB_84_U137 | ~new_P1_SUB_84_U138 | ~new_P1_SUB_84_U142 | ~new_P1_SUB_84_U141;
  assign new_P1_SUB_84_U215 = ~P1_IR_REG_22_ | ~new_P1_SUB_84_U214;
  assign new_P1_SUB_84_U216 = ~P1_IR_REG_20_ | ~new_P1_SUB_84_U198;
  assign new_P1_SUB_84_U217 = ~P1_IR_REG_19_ | ~new_P1_SUB_84_U197;
  assign new_P1_SUB_84_U218 = ~new_P1_SUB_84_U196 | ~new_P1_SUB_84_U176;
  assign new_P1_SUB_84_U219 = ~P1_IR_REG_18_ | ~new_P1_SUB_84_U218;
  assign new_P1_SUB_84_U220 = ~P1_IR_REG_16_ | ~new_P1_SUB_84_U195;
  assign new_P1_SUB_84_U221 = ~P1_IR_REG_15_ | ~new_P1_SUB_84_U36;
  assign new_P1_SUB_84_U222 = ~new_P1_SUB_84_U193 | ~new_P1_SUB_84_U178;
  assign new_P1_SUB_84_U223 = ~P1_IR_REG_14_ | ~new_P1_SUB_84_U222;
  assign new_P1_SUB_84_U224 = ~P1_IR_REG_12_ | ~new_P1_SUB_84_U192;
  assign new_P1_SUB_84_U225 = ~P1_IR_REG_11_ | ~new_P1_SUB_84_U38;
  assign new_P1_SUB_84_U226 = ~new_P1_SUB_84_U184 | ~new_P1_SUB_84_U159;
  assign new_P1_SUB_84_U227 = ~P1_IR_REG_10_ | ~new_P1_SUB_84_U226;
  assign new_P1_SUB_84_U228 = ~new_P1_SUB_84_U205 | ~new_P1_SUB_84_U164;
  assign new_P1_SUB_84_U229 = ~new_P1_SUB_84_U76 | ~new_P1_SUB_84_U71;
  assign new_P1_SUB_84_U230 = ~new_P1_SUB_84_U27;
  assign new_P1_SUB_84_U231 = ~new_P1_SUB_84_U86 | ~new_P1_SUB_84_U81;
  assign new_P1_SUB_84_U232 = ~P1_IR_REG_9_ | ~new_P1_SUB_84_U28;
  assign new_P1_SUB_84_U233 = ~new_P1_SUB_84_U184 | ~new_P1_SUB_84_U159;
  assign new_P1_SUB_84_U234 = ~P1_IR_REG_5_ | ~new_P1_SUB_84_U29;
  assign new_P1_SUB_84_U235 = ~new_P1_SUB_84_U181 | ~new_P1_SUB_84_U161;
  assign new_P1_SUB_84_U236 = ~new_P1_SUB_84_U228 | ~new_P1_SUB_84_U163;
  assign new_P1_SUB_84_U237 = ~P1_IR_REG_31_ | ~new_P1_SUB_84_U205 | ~new_P1_SUB_84_U164;
  assign new_P1_SUB_84_U238 = ~P1_IR_REG_30_ | ~new_P1_SUB_84_U33;
  assign new_P1_SUB_84_U239 = ~new_P1_SUB_84_U205 | ~new_P1_SUB_84_U164;
  assign new_P1_SUB_84_U240 = ~new_P1_SUB_84_U203 | ~P1_IR_REG_27_;
  assign new_P1_SUB_84_U241 = ~new_P1_SUB_84_U231 | ~new_P1_SUB_84_U166;
  assign new_P1_SUB_84_U242 = ~P1_IR_REG_25_ | ~new_P1_SUB_84_U169;
  assign new_P1_SUB_84_U243 = ~new_P1_SUB_84_U202 | ~new_P1_SUB_84_U168;
  assign new_P1_SUB_84_U244 = ~P1_IR_REG_21_ | ~new_P1_SUB_84_U172;
  assign new_P1_SUB_84_U245 = ~new_P1_SUB_84_U199 | ~new_P1_SUB_84_U171;
  assign new_P1_SUB_84_U246 = ~P1_IR_REG_1_ | ~new_P1_SUB_84_U175;
  assign new_P1_SUB_84_U247 = ~P1_IR_REG_0_ | ~new_P1_SUB_84_U174;
  assign new_P1_SUB_84_U248 = ~P1_IR_REG_17_ | ~new_P1_SUB_84_U34;
  assign new_P1_SUB_84_U249 = ~new_P1_SUB_84_U196 | ~new_P1_SUB_84_U176;
  assign new_P1_SUB_84_U250 = ~P1_IR_REG_13_ | ~new_P1_SUB_84_U35;
  assign new_P1_SUB_84_U251 = ~new_P1_SUB_84_U193 | ~new_P1_SUB_84_U178;
  assign new_P1_R1309_U6 = ~new_P1_U3059;
  assign new_P1_R1309_U7 = ~new_P1_U3056;
  assign new_P1_R1309_U8 = new_P1_R1309_U10 & new_P1_R1309_U9;
  assign new_P1_R1309_U9 = ~new_P1_U3056 | ~new_P1_R1309_U6;
  assign new_P1_R1309_U10 = ~new_P1_U3059 | ~new_P1_R1309_U7;
  assign new_P1_R1282_U6 = new_P1_R1282_U135 & new_P1_R1282_U35;
  assign new_P1_R1282_U7 = new_P1_R1282_U133 & new_P1_R1282_U36;
  assign new_P1_R1282_U8 = new_P1_R1282_U132 & new_P1_R1282_U37;
  assign new_P1_R1282_U9 = new_P1_R1282_U131 & new_P1_R1282_U38;
  assign new_P1_R1282_U10 = new_P1_R1282_U129 & new_P1_R1282_U39;
  assign new_P1_R1282_U11 = new_P1_R1282_U128 & new_P1_R1282_U40;
  assign new_P1_R1282_U12 = new_P1_R1282_U127 & new_P1_R1282_U41;
  assign new_P1_R1282_U13 = new_P1_R1282_U125 & new_P1_R1282_U42;
  assign new_P1_R1282_U14 = new_P1_R1282_U123 & new_P1_R1282_U43;
  assign new_P1_R1282_U15 = new_P1_R1282_U121 & new_P1_R1282_U44;
  assign new_P1_R1282_U16 = new_P1_R1282_U119 & new_P1_R1282_U45;
  assign new_P1_R1282_U17 = new_P1_R1282_U117 & new_P1_R1282_U46;
  assign new_P1_R1282_U18 = new_P1_R1282_U115 & new_P1_R1282_U25;
  assign new_P1_R1282_U19 = new_P1_R1282_U113 & new_P1_R1282_U67;
  assign new_P1_R1282_U20 = new_P1_R1282_U98 & new_P1_R1282_U26;
  assign new_P1_R1282_U21 = new_P1_R1282_U97 & new_P1_R1282_U27;
  assign new_P1_R1282_U22 = new_P1_R1282_U96 & new_P1_R1282_U28;
  assign new_P1_R1282_U23 = new_P1_R1282_U94 & new_P1_R1282_U29;
  assign new_P1_R1282_U24 = new_P1_R1282_U93 & new_P1_R1282_U30;
  assign new_P1_R1282_U25 = new_P1_U3455 | new_P1_U3458 | new_P1_U3450;
  assign new_P1_R1282_U26 = ~new_P1_R1282_U87 | ~new_P1_R1282_U34;
  assign new_P1_R1282_U27 = ~new_P1_R1282_U88 | ~new_P1_R1282_U33;
  assign new_P1_R1282_U28 = ~new_P1_R1282_U58 | ~new_P1_R1282_U89;
  assign new_P1_R1282_U29 = ~new_P1_R1282_U90 | ~new_P1_R1282_U32;
  assign new_P1_R1282_U30 = ~new_P1_R1282_U91 | ~new_P1_R1282_U31;
  assign new_P1_R1282_U31 = ~new_P1_U3476;
  assign new_P1_R1282_U32 = ~new_P1_U3473;
  assign new_P1_R1282_U33 = ~new_P1_U3464;
  assign new_P1_R1282_U34 = ~new_P1_U3461;
  assign new_P1_R1282_U35 = ~new_P1_R1282_U59 | ~new_P1_R1282_U92;
  assign new_P1_R1282_U36 = ~new_P1_R1282_U99 | ~new_P1_R1282_U56;
  assign new_P1_R1282_U37 = ~new_P1_R1282_U100 | ~new_P1_R1282_U55;
  assign new_P1_R1282_U38 = ~new_P1_R1282_U60 | ~new_P1_R1282_U101;
  assign new_P1_R1282_U39 = ~new_P1_R1282_U102 | ~new_P1_R1282_U54;
  assign new_P1_R1282_U40 = ~new_P1_R1282_U103 | ~new_P1_R1282_U53;
  assign new_P1_R1282_U41 = ~new_P1_R1282_U61 | ~new_P1_R1282_U104;
  assign new_P1_R1282_U42 = ~new_P1_R1282_U52 | ~new_P1_R1282_U105 | ~new_P1_R1282_U81;
  assign new_P1_R1282_U43 = ~new_P1_R1282_U51 | ~new_P1_R1282_U106 | ~new_P1_R1282_U77;
  assign new_P1_R1282_U44 = ~new_P1_R1282_U50 | ~new_P1_R1282_U107 | ~new_P1_R1282_U75;
  assign new_P1_R1282_U45 = ~new_P1_R1282_U49 | ~new_P1_R1282_U108 | ~new_P1_R1282_U73;
  assign new_P1_R1282_U46 = ~new_P1_R1282_U48 | ~new_P1_R1282_U109 | ~new_P1_R1282_U71;
  assign new_P1_R1282_U47 = ~new_P1_U3984;
  assign new_P1_R1282_U48 = ~new_P1_U3974;
  assign new_P1_R1282_U49 = ~new_P1_U3976;
  assign new_P1_R1282_U50 = ~new_P1_U3978;
  assign new_P1_R1282_U51 = ~new_P1_U3980;
  assign new_P1_R1282_U52 = ~new_P1_U3982;
  assign new_P1_R1282_U53 = ~new_P1_U3500;
  assign new_P1_R1282_U54 = ~new_P1_U3497;
  assign new_P1_R1282_U55 = ~new_P1_U3488;
  assign new_P1_R1282_U56 = ~new_P1_U3485;
  assign new_P1_R1282_U57 = ~new_P1_R1282_U153 | ~new_P1_R1282_U152;
  assign new_P1_R1282_U58 = ~new_P1_U3467 & ~new_P1_U3470;
  assign new_P1_R1282_U59 = ~new_P1_U3482 & ~new_P1_U3479;
  assign new_P1_R1282_U60 = ~new_P1_U3491 & ~new_P1_U3494;
  assign new_P1_R1282_U61 = ~new_P1_U3503 & ~new_P1_U3506;
  assign new_P1_R1282_U62 = ~new_P1_U3479;
  assign new_P1_R1282_U63 = new_P1_R1282_U137 & new_P1_R1282_U136;
  assign new_P1_R1282_U64 = ~new_P1_U3467;
  assign new_P1_R1282_U65 = new_P1_R1282_U139 & new_P1_R1282_U138;
  assign new_P1_R1282_U66 = ~new_P1_U3983;
  assign new_P1_R1282_U67 = ~new_P1_R1282_U47 | ~new_P1_R1282_U110 | ~new_P1_R1282_U69;
  assign new_P1_R1282_U68 = new_P1_R1282_U141 & new_P1_R1282_U140;
  assign new_P1_R1282_U69 = ~new_P1_U3985;
  assign new_P1_R1282_U70 = new_P1_R1282_U143 & new_P1_R1282_U142;
  assign new_P1_R1282_U71 = ~new_P1_U3975;
  assign new_P1_R1282_U72 = new_P1_R1282_U145 & new_P1_R1282_U144;
  assign new_P1_R1282_U73 = ~new_P1_U3977;
  assign new_P1_R1282_U74 = new_P1_R1282_U147 & new_P1_R1282_U146;
  assign new_P1_R1282_U75 = ~new_P1_U3979;
  assign new_P1_R1282_U76 = new_P1_R1282_U149 & new_P1_R1282_U148;
  assign new_P1_R1282_U77 = ~new_P1_U3981;
  assign new_P1_R1282_U78 = new_P1_R1282_U151 & new_P1_R1282_U150;
  assign new_P1_R1282_U79 = ~new_P1_U3455;
  assign new_P1_R1282_U80 = ~new_P1_U3450;
  assign new_P1_R1282_U81 = ~new_P1_U3508;
  assign new_P1_R1282_U82 = new_P1_R1282_U155 & new_P1_R1282_U154;
  assign new_P1_R1282_U83 = ~new_P1_U3503;
  assign new_P1_R1282_U84 = new_P1_R1282_U157 & new_P1_R1282_U156;
  assign new_P1_R1282_U85 = ~new_P1_U3491;
  assign new_P1_R1282_U86 = new_P1_R1282_U159 & new_P1_R1282_U158;
  assign new_P1_R1282_U87 = ~new_P1_R1282_U25;
  assign new_P1_R1282_U88 = ~new_P1_R1282_U26;
  assign new_P1_R1282_U89 = ~new_P1_R1282_U27;
  assign new_P1_R1282_U90 = ~new_P1_R1282_U28;
  assign new_P1_R1282_U91 = ~new_P1_R1282_U29;
  assign new_P1_R1282_U92 = ~new_P1_R1282_U30;
  assign new_P1_R1282_U93 = ~new_P1_U3476 | ~new_P1_R1282_U29;
  assign new_P1_R1282_U94 = ~new_P1_U3473 | ~new_P1_R1282_U28;
  assign new_P1_R1282_U95 = ~new_P1_R1282_U89 | ~new_P1_R1282_U64;
  assign new_P1_R1282_U96 = ~new_P1_U3470 | ~new_P1_R1282_U95;
  assign new_P1_R1282_U97 = ~new_P1_U3464 | ~new_P1_R1282_U26;
  assign new_P1_R1282_U98 = ~new_P1_U3461 | ~new_P1_R1282_U25;
  assign new_P1_R1282_U99 = ~new_P1_R1282_U35;
  assign new_P1_R1282_U100 = ~new_P1_R1282_U36;
  assign new_P1_R1282_U101 = ~new_P1_R1282_U37;
  assign new_P1_R1282_U102 = ~new_P1_R1282_U38;
  assign new_P1_R1282_U103 = ~new_P1_R1282_U39;
  assign new_P1_R1282_U104 = ~new_P1_R1282_U40;
  assign new_P1_R1282_U105 = ~new_P1_R1282_U41;
  assign new_P1_R1282_U106 = ~new_P1_R1282_U42;
  assign new_P1_R1282_U107 = ~new_P1_R1282_U43;
  assign new_P1_R1282_U108 = ~new_P1_R1282_U44;
  assign new_P1_R1282_U109 = ~new_P1_R1282_U45;
  assign new_P1_R1282_U110 = ~new_P1_R1282_U46;
  assign new_P1_R1282_U111 = ~new_P1_R1282_U67;
  assign new_P1_R1282_U112 = ~new_P1_R1282_U110 | ~new_P1_R1282_U69;
  assign new_P1_R1282_U113 = ~new_P1_U3984 | ~new_P1_R1282_U112;
  assign new_P1_R1282_U114 = new_P1_U3455 | new_P1_U3450;
  assign new_P1_R1282_U115 = ~new_P1_U3458 | ~new_P1_R1282_U114;
  assign new_P1_R1282_U116 = ~new_P1_R1282_U109 | ~new_P1_R1282_U71;
  assign new_P1_R1282_U117 = ~new_P1_U3974 | ~new_P1_R1282_U116;
  assign new_P1_R1282_U118 = ~new_P1_R1282_U108 | ~new_P1_R1282_U73;
  assign new_P1_R1282_U119 = ~new_P1_U3976 | ~new_P1_R1282_U118;
  assign new_P1_R1282_U120 = ~new_P1_R1282_U107 | ~new_P1_R1282_U75;
  assign new_P1_R1282_U121 = ~new_P1_U3978 | ~new_P1_R1282_U120;
  assign new_P1_R1282_U122 = ~new_P1_R1282_U106 | ~new_P1_R1282_U77;
  assign new_P1_R1282_U123 = ~new_P1_U3980 | ~new_P1_R1282_U122;
  assign new_P1_R1282_U124 = ~new_P1_R1282_U105 | ~new_P1_R1282_U81;
  assign new_P1_R1282_U125 = ~new_P1_U3982 | ~new_P1_R1282_U124;
  assign new_P1_R1282_U126 = ~new_P1_R1282_U104 | ~new_P1_R1282_U83;
  assign new_P1_R1282_U127 = ~new_P1_U3506 | ~new_P1_R1282_U126;
  assign new_P1_R1282_U128 = ~new_P1_U3500 | ~new_P1_R1282_U39;
  assign new_P1_R1282_U129 = ~new_P1_U3497 | ~new_P1_R1282_U38;
  assign new_P1_R1282_U130 = ~new_P1_R1282_U101 | ~new_P1_R1282_U85;
  assign new_P1_R1282_U131 = ~new_P1_U3494 | ~new_P1_R1282_U130;
  assign new_P1_R1282_U132 = ~new_P1_U3488 | ~new_P1_R1282_U36;
  assign new_P1_R1282_U133 = ~new_P1_U3485 | ~new_P1_R1282_U35;
  assign new_P1_R1282_U134 = ~new_P1_R1282_U92 | ~new_P1_R1282_U62;
  assign new_P1_R1282_U135 = ~new_P1_U3482 | ~new_P1_R1282_U134;
  assign new_P1_R1282_U136 = ~new_P1_U3479 | ~new_P1_R1282_U30;
  assign new_P1_R1282_U137 = ~new_P1_R1282_U92 | ~new_P1_R1282_U62;
  assign new_P1_R1282_U138 = ~new_P1_U3467 | ~new_P1_R1282_U27;
  assign new_P1_R1282_U139 = ~new_P1_R1282_U89 | ~new_P1_R1282_U64;
  assign new_P1_R1282_U140 = ~new_P1_U3983 | ~new_P1_R1282_U67;
  assign new_P1_R1282_U141 = ~new_P1_R1282_U111 | ~new_P1_R1282_U66;
  assign new_P1_R1282_U142 = ~new_P1_U3985 | ~new_P1_R1282_U46;
  assign new_P1_R1282_U143 = ~new_P1_R1282_U110 | ~new_P1_R1282_U69;
  assign new_P1_R1282_U144 = ~new_P1_U3975 | ~new_P1_R1282_U45;
  assign new_P1_R1282_U145 = ~new_P1_R1282_U109 | ~new_P1_R1282_U71;
  assign new_P1_R1282_U146 = ~new_P1_U3977 | ~new_P1_R1282_U44;
  assign new_P1_R1282_U147 = ~new_P1_R1282_U108 | ~new_P1_R1282_U73;
  assign new_P1_R1282_U148 = ~new_P1_U3979 | ~new_P1_R1282_U43;
  assign new_P1_R1282_U149 = ~new_P1_R1282_U107 | ~new_P1_R1282_U75;
  assign new_P1_R1282_U150 = ~new_P1_U3981 | ~new_P1_R1282_U42;
  assign new_P1_R1282_U151 = ~new_P1_R1282_U106 | ~new_P1_R1282_U77;
  assign new_P1_R1282_U152 = ~new_P1_U3455 | ~new_P1_R1282_U80;
  assign new_P1_R1282_U153 = ~new_P1_U3450 | ~new_P1_R1282_U79;
  assign new_P1_R1282_U154 = ~new_P1_U3508 | ~new_P1_R1282_U41;
  assign new_P1_R1282_U155 = ~new_P1_R1282_U105 | ~new_P1_R1282_U81;
  assign new_P1_R1282_U156 = ~new_P1_U3503 | ~new_P1_R1282_U40;
  assign new_P1_R1282_U157 = ~new_P1_R1282_U104 | ~new_P1_R1282_U83;
  assign new_P1_R1282_U158 = ~new_P1_U3491 | ~new_P1_R1282_U37;
  assign new_P1_R1282_U159 = ~new_P1_R1282_U101 | ~new_P1_R1282_U85;
  assign new_P1_R1240_U4 = new_P1_R1240_U178 & new_P1_R1240_U177;
  assign new_P1_R1240_U5 = new_P1_R1240_U179 & new_P1_R1240_U180;
  assign new_P1_R1240_U6 = new_P1_R1240_U196 & new_P1_R1240_U195;
  assign new_P1_R1240_U7 = new_P1_R1240_U236 & new_P1_R1240_U235;
  assign new_P1_R1240_U8 = new_P1_R1240_U245 & new_P1_R1240_U244;
  assign new_P1_R1240_U9 = new_P1_R1240_U263 & new_P1_R1240_U262;
  assign new_P1_R1240_U10 = new_P1_R1240_U271 & new_P1_R1240_U270;
  assign new_P1_R1240_U11 = new_P1_R1240_U350 & new_P1_R1240_U347;
  assign new_P1_R1240_U12 = new_P1_R1240_U343 & new_P1_R1240_U340;
  assign new_P1_R1240_U13 = new_P1_R1240_U334 & new_P1_R1240_U331;
  assign new_P1_R1240_U14 = new_P1_R1240_U325 & new_P1_R1240_U322;
  assign new_P1_R1240_U15 = new_P1_R1240_U319 & new_P1_R1240_U317;
  assign new_P1_R1240_U16 = new_P1_R1240_U312 & new_P1_R1240_U309;
  assign new_P1_R1240_U17 = new_P1_R1240_U234 & new_P1_R1240_U231;
  assign new_P1_R1240_U18 = new_P1_R1240_U226 & new_P1_R1240_U223;
  assign new_P1_R1240_U19 = new_P1_R1240_U212 & new_P1_R1240_U209;
  assign new_P1_R1240_U20 = ~new_P1_U3470;
  assign new_P1_R1240_U21 = ~new_P1_U3071;
  assign new_P1_R1240_U22 = ~new_P1_U3070;
  assign new_P1_R1240_U23 = ~new_P1_U3071 | ~new_P1_U3470;
  assign new_P1_R1240_U24 = ~new_P1_U3473;
  assign new_P1_R1240_U25 = ~new_P1_U3464;
  assign new_P1_R1240_U26 = ~new_P1_U3060;
  assign new_P1_R1240_U27 = ~new_P1_U3067;
  assign new_P1_R1240_U28 = ~new_P1_U3458;
  assign new_P1_R1240_U29 = ~new_P1_U3068;
  assign new_P1_R1240_U30 = ~new_P1_U3450;
  assign new_P1_R1240_U31 = ~new_P1_U3077;
  assign new_P1_R1240_U32 = ~new_P1_U3077 | ~new_P1_U3450;
  assign new_P1_R1240_U33 = ~new_P1_U3461;
  assign new_P1_R1240_U34 = ~new_P1_U3064;
  assign new_P1_R1240_U35 = ~new_P1_U3060 | ~new_P1_U3464;
  assign new_P1_R1240_U36 = ~new_P1_U3467;
  assign new_P1_R1240_U37 = ~new_P1_U3476;
  assign new_P1_R1240_U38 = ~new_P1_U3084;
  assign new_P1_R1240_U39 = ~new_P1_U3083;
  assign new_P1_R1240_U40 = ~new_P1_U3479;
  assign new_P1_R1240_U41 = ~new_P1_R1240_U62 | ~new_P1_R1240_U204;
  assign new_P1_R1240_U42 = ~new_P1_R1240_U118 | ~new_P1_R1240_U192;
  assign new_P1_R1240_U43 = ~new_P1_R1240_U181 | ~new_P1_R1240_U182;
  assign new_P1_R1240_U44 = ~new_P1_U3455 | ~new_P1_U3078;
  assign new_P1_R1240_U45 = ~new_P1_R1240_U122 | ~new_P1_R1240_U218;
  assign new_P1_R1240_U46 = ~new_P1_R1240_U215 | ~new_P1_R1240_U214;
  assign new_P1_R1240_U47 = ~new_P1_U3975;
  assign new_P1_R1240_U48 = ~new_P1_U3053;
  assign new_P1_R1240_U49 = ~new_P1_U3057;
  assign new_P1_R1240_U50 = ~new_P1_U3976;
  assign new_P1_R1240_U51 = ~new_P1_U3977;
  assign new_P1_R1240_U52 = ~new_P1_U3058;
  assign new_P1_R1240_U53 = ~new_P1_U3978;
  assign new_P1_R1240_U54 = ~new_P1_U3065;
  assign new_P1_R1240_U55 = ~new_P1_U3981;
  assign new_P1_R1240_U56 = ~new_P1_U3075;
  assign new_P1_R1240_U57 = ~new_P1_U3500;
  assign new_P1_R1240_U58 = ~new_P1_U3073;
  assign new_P1_R1240_U59 = ~new_P1_U3069;
  assign new_P1_R1240_U60 = ~new_P1_U3073 | ~new_P1_U3500;
  assign new_P1_R1240_U61 = ~new_P1_U3503;
  assign new_P1_R1240_U62 = ~new_P1_U3084 | ~new_P1_U3476;
  assign new_P1_R1240_U63 = ~new_P1_U3482;
  assign new_P1_R1240_U64 = ~new_P1_U3062;
  assign new_P1_R1240_U65 = ~new_P1_U3488;
  assign new_P1_R1240_U66 = ~new_P1_U3072;
  assign new_P1_R1240_U67 = ~new_P1_U3485;
  assign new_P1_R1240_U68 = ~new_P1_U3063;
  assign new_P1_R1240_U69 = ~new_P1_U3063 | ~new_P1_U3485;
  assign new_P1_R1240_U70 = ~new_P1_U3491;
  assign new_P1_R1240_U71 = ~new_P1_U3080;
  assign new_P1_R1240_U72 = ~new_P1_U3494;
  assign new_P1_R1240_U73 = ~new_P1_U3079;
  assign new_P1_R1240_U74 = ~new_P1_U3497;
  assign new_P1_R1240_U75 = ~new_P1_U3074;
  assign new_P1_R1240_U76 = ~new_P1_U3506;
  assign new_P1_R1240_U77 = ~new_P1_U3082;
  assign new_P1_R1240_U78 = ~new_P1_U3082 | ~new_P1_U3506;
  assign new_P1_R1240_U79 = ~new_P1_U3508;
  assign new_P1_R1240_U80 = ~new_P1_U3081;
  assign new_P1_R1240_U81 = ~new_P1_U3081 | ~new_P1_U3508;
  assign new_P1_R1240_U82 = ~new_P1_U3982;
  assign new_P1_R1240_U83 = ~new_P1_U3980;
  assign new_P1_R1240_U84 = ~new_P1_U3061;
  assign new_P1_R1240_U85 = ~new_P1_U3979;
  assign new_P1_R1240_U86 = ~new_P1_U3066;
  assign new_P1_R1240_U87 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1240_U88 = ~new_P1_U3054;
  assign new_P1_R1240_U89 = ~new_P1_U3974;
  assign new_P1_R1240_U90 = ~new_P1_R1240_U305 | ~new_P1_R1240_U175;
  assign new_P1_R1240_U91 = ~new_P1_U3076;
  assign new_P1_R1240_U92 = ~new_P1_R1240_U78 | ~new_P1_R1240_U314;
  assign new_P1_R1240_U93 = ~new_P1_R1240_U260 | ~new_P1_R1240_U259;
  assign new_P1_R1240_U94 = ~new_P1_R1240_U69 | ~new_P1_R1240_U336;
  assign new_P1_R1240_U95 = ~new_P1_R1240_U456 | ~new_P1_R1240_U455;
  assign new_P1_R1240_U96 = ~new_P1_R1240_U503 | ~new_P1_R1240_U502;
  assign new_P1_R1240_U97 = ~new_P1_R1240_U374 | ~new_P1_R1240_U373;
  assign new_P1_R1240_U98 = ~new_P1_R1240_U379 | ~new_P1_R1240_U378;
  assign new_P1_R1240_U99 = ~new_P1_R1240_U386 | ~new_P1_R1240_U385;
  assign new_P1_R1240_U100 = ~new_P1_R1240_U393 | ~new_P1_R1240_U392;
  assign new_P1_R1240_U101 = ~new_P1_R1240_U398 | ~new_P1_R1240_U397;
  assign new_P1_R1240_U102 = ~new_P1_R1240_U407 | ~new_P1_R1240_U406;
  assign new_P1_R1240_U103 = ~new_P1_R1240_U414 | ~new_P1_R1240_U413;
  assign new_P1_R1240_U104 = ~new_P1_R1240_U421 | ~new_P1_R1240_U420;
  assign new_P1_R1240_U105 = ~new_P1_R1240_U428 | ~new_P1_R1240_U427;
  assign new_P1_R1240_U106 = ~new_P1_R1240_U433 | ~new_P1_R1240_U432;
  assign new_P1_R1240_U107 = ~new_P1_R1240_U440 | ~new_P1_R1240_U439;
  assign new_P1_R1240_U108 = ~new_P1_R1240_U447 | ~new_P1_R1240_U446;
  assign new_P1_R1240_U109 = ~new_P1_R1240_U461 | ~new_P1_R1240_U460;
  assign new_P1_R1240_U110 = ~new_P1_R1240_U466 | ~new_P1_R1240_U465;
  assign new_P1_R1240_U111 = ~new_P1_R1240_U473 | ~new_P1_R1240_U472;
  assign new_P1_R1240_U112 = ~new_P1_R1240_U480 | ~new_P1_R1240_U479;
  assign new_P1_R1240_U113 = ~new_P1_R1240_U487 | ~new_P1_R1240_U486;
  assign new_P1_R1240_U114 = ~new_P1_R1240_U494 | ~new_P1_R1240_U493;
  assign new_P1_R1240_U115 = ~new_P1_R1240_U499 | ~new_P1_R1240_U498;
  assign new_P1_R1240_U116 = new_P1_U3458 & new_P1_U3068;
  assign new_P1_R1240_U117 = new_P1_R1240_U188 & new_P1_R1240_U186;
  assign new_P1_R1240_U118 = new_P1_R1240_U193 & new_P1_R1240_U191;
  assign new_P1_R1240_U119 = new_P1_R1240_U200 & new_P1_R1240_U199;
  assign new_P1_R1240_U120 = new_P1_R1240_U23 & new_P1_R1240_U381 & new_P1_R1240_U380;
  assign new_P1_R1240_U121 = new_P1_R1240_U211 & new_P1_R1240_U6;
  assign new_P1_R1240_U122 = new_P1_R1240_U219 & new_P1_R1240_U217;
  assign new_P1_R1240_U123 = new_P1_R1240_U35 & new_P1_R1240_U388 & new_P1_R1240_U387;
  assign new_P1_R1240_U124 = new_P1_R1240_U225 & new_P1_R1240_U4;
  assign new_P1_R1240_U125 = new_P1_R1240_U233 & new_P1_R1240_U180;
  assign new_P1_R1240_U126 = new_P1_R1240_U203 & new_P1_R1240_U7;
  assign new_P1_R1240_U127 = new_P1_R1240_U238 & new_P1_R1240_U170;
  assign new_P1_R1240_U128 = new_P1_R1240_U249 & new_P1_R1240_U8;
  assign new_P1_R1240_U129 = new_P1_R1240_U247 & new_P1_R1240_U171;
  assign new_P1_R1240_U130 = new_P1_R1240_U267 & new_P1_R1240_U266;
  assign new_P1_R1240_U131 = new_P1_R1240_U10 & new_P1_R1240_U281;
  assign new_P1_R1240_U132 = new_P1_R1240_U284 & new_P1_R1240_U279;
  assign new_P1_R1240_U133 = new_P1_R1240_U300 & new_P1_R1240_U297;
  assign new_P1_R1240_U134 = new_P1_R1240_U367 & new_P1_R1240_U301;
  assign new_P1_R1240_U135 = new_P1_R1240_U159 & new_P1_R1240_U277;
  assign new_P1_R1240_U136 = new_P1_R1240_U81 & new_P1_R1240_U454 & new_P1_R1240_U453;
  assign new_P1_R1240_U137 = new_P1_R1240_U60 & new_P1_R1240_U468 & new_P1_R1240_U467;
  assign new_P1_R1240_U138 = new_P1_R1240_U333 & new_P1_R1240_U9;
  assign new_P1_R1240_U139 = new_P1_R1240_U171 & new_P1_R1240_U489 & new_P1_R1240_U488;
  assign new_P1_R1240_U140 = new_P1_R1240_U342 & new_P1_R1240_U8;
  assign new_P1_R1240_U141 = new_P1_R1240_U170 & new_P1_R1240_U501 & new_P1_R1240_U500;
  assign new_P1_R1240_U142 = new_P1_R1240_U349 & new_P1_R1240_U7;
  assign new_P1_R1240_U143 = ~new_P1_R1240_U119 | ~new_P1_R1240_U201;
  assign new_P1_R1240_U144 = ~new_P1_R1240_U216 | ~new_P1_R1240_U228;
  assign new_P1_R1240_U145 = ~new_P1_U3055;
  assign new_P1_R1240_U146 = ~new_P1_U3985;
  assign new_P1_R1240_U147 = new_P1_R1240_U402 & new_P1_R1240_U401;
  assign new_P1_R1240_U148 = ~new_P1_R1240_U363 | ~new_P1_R1240_U303 | ~new_P1_R1240_U168;
  assign new_P1_R1240_U149 = new_P1_R1240_U409 & new_P1_R1240_U408;
  assign new_P1_R1240_U150 = ~new_P1_R1240_U134 | ~new_P1_R1240_U369 | ~new_P1_R1240_U368;
  assign new_P1_R1240_U151 = new_P1_R1240_U416 & new_P1_R1240_U415;
  assign new_P1_R1240_U152 = ~new_P1_R1240_U87 | ~new_P1_R1240_U364 | ~new_P1_R1240_U298;
  assign new_P1_R1240_U153 = new_P1_R1240_U423 & new_P1_R1240_U422;
  assign new_P1_R1240_U154 = ~new_P1_R1240_U292 | ~new_P1_R1240_U291;
  assign new_P1_R1240_U155 = new_P1_R1240_U435 & new_P1_R1240_U434;
  assign new_P1_R1240_U156 = ~new_P1_R1240_U288 | ~new_P1_R1240_U287;
  assign new_P1_R1240_U157 = new_P1_R1240_U442 & new_P1_R1240_U441;
  assign new_P1_R1240_U158 = ~new_P1_R1240_U132 | ~new_P1_R1240_U283;
  assign new_P1_R1240_U159 = new_P1_R1240_U449 & new_P1_R1240_U448;
  assign new_P1_R1240_U160 = ~new_P1_R1240_U44 | ~new_P1_R1240_U326;
  assign new_P1_R1240_U161 = ~new_P1_R1240_U130 | ~new_P1_R1240_U268;
  assign new_P1_R1240_U162 = new_P1_R1240_U475 & new_P1_R1240_U474;
  assign new_P1_R1240_U163 = ~new_P1_R1240_U256 | ~new_P1_R1240_U255;
  assign new_P1_R1240_U164 = new_P1_R1240_U482 & new_P1_R1240_U481;
  assign new_P1_R1240_U165 = ~new_P1_R1240_U252 | ~new_P1_R1240_U251;
  assign new_P1_R1240_U166 = ~new_P1_R1240_U242 | ~new_P1_R1240_U241;
  assign new_P1_R1240_U167 = ~new_P1_R1240_U366 | ~new_P1_R1240_U365;
  assign new_P1_R1240_U168 = ~new_P1_U3054 | ~new_P1_R1240_U150;
  assign new_P1_R1240_U169 = ~new_P1_R1240_U35;
  assign new_P1_R1240_U170 = ~new_P1_U3479 | ~new_P1_U3083;
  assign new_P1_R1240_U171 = ~new_P1_U3072 | ~new_P1_U3488;
  assign new_P1_R1240_U172 = ~new_P1_U3058 | ~new_P1_U3977;
  assign new_P1_R1240_U173 = ~new_P1_R1240_U69;
  assign new_P1_R1240_U174 = ~new_P1_R1240_U78;
  assign new_P1_R1240_U175 = ~new_P1_U3065 | ~new_P1_U3978;
  assign new_P1_R1240_U176 = ~new_P1_R1240_U62;
  assign new_P1_R1240_U177 = new_P1_U3067 | new_P1_U3467;
  assign new_P1_R1240_U178 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1240_U179 = new_P1_U3461 | new_P1_U3064;
  assign new_P1_R1240_U180 = new_P1_U3458 | new_P1_U3068;
  assign new_P1_R1240_U181 = ~new_P1_R1240_U32;
  assign new_P1_R1240_U182 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1240_U183 = ~new_P1_R1240_U43;
  assign new_P1_R1240_U184 = ~new_P1_R1240_U44;
  assign new_P1_R1240_U185 = ~new_P1_R1240_U43 | ~new_P1_R1240_U44;
  assign new_P1_R1240_U186 = ~new_P1_R1240_U116 | ~new_P1_R1240_U179;
  assign new_P1_R1240_U187 = ~new_P1_R1240_U5 | ~new_P1_R1240_U185;
  assign new_P1_R1240_U188 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1240_U189 = ~new_P1_R1240_U117 | ~new_P1_R1240_U187;
  assign new_P1_R1240_U190 = ~new_P1_R1240_U36 | ~new_P1_R1240_U35;
  assign new_P1_R1240_U191 = ~new_P1_U3067 | ~new_P1_R1240_U190;
  assign new_P1_R1240_U192 = ~new_P1_R1240_U4 | ~new_P1_R1240_U189;
  assign new_P1_R1240_U193 = ~new_P1_U3467 | ~new_P1_R1240_U169;
  assign new_P1_R1240_U194 = ~new_P1_R1240_U42;
  assign new_P1_R1240_U195 = new_P1_U3070 | new_P1_U3473;
  assign new_P1_R1240_U196 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1240_U197 = ~new_P1_R1240_U23;
  assign new_P1_R1240_U198 = ~new_P1_R1240_U24 | ~new_P1_R1240_U23;
  assign new_P1_R1240_U199 = ~new_P1_U3070 | ~new_P1_R1240_U198;
  assign new_P1_R1240_U200 = ~new_P1_U3473 | ~new_P1_R1240_U197;
  assign new_P1_R1240_U201 = ~new_P1_R1240_U6 | ~new_P1_R1240_U42;
  assign new_P1_R1240_U202 = ~new_P1_R1240_U143;
  assign new_P1_R1240_U203 = new_P1_U3476 | new_P1_U3084;
  assign new_P1_R1240_U204 = ~new_P1_R1240_U203 | ~new_P1_R1240_U143;
  assign new_P1_R1240_U205 = ~new_P1_R1240_U41;
  assign new_P1_R1240_U206 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1240_U207 = new_P1_U3470 | new_P1_U3071;
  assign new_P1_R1240_U208 = ~new_P1_R1240_U207 | ~new_P1_R1240_U42;
  assign new_P1_R1240_U209 = ~new_P1_R1240_U120 | ~new_P1_R1240_U208;
  assign new_P1_R1240_U210 = ~new_P1_R1240_U194 | ~new_P1_R1240_U23;
  assign new_P1_R1240_U211 = ~new_P1_U3473 | ~new_P1_U3070;
  assign new_P1_R1240_U212 = ~new_P1_R1240_U121 | ~new_P1_R1240_U210;
  assign new_P1_R1240_U213 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1240_U214 = ~new_P1_R1240_U184 | ~new_P1_R1240_U180;
  assign new_P1_R1240_U215 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1240_U216 = ~new_P1_R1240_U46;
  assign new_P1_R1240_U217 = ~new_P1_R1240_U183 | ~new_P1_R1240_U5;
  assign new_P1_R1240_U218 = ~new_P1_R1240_U46 | ~new_P1_R1240_U179;
  assign new_P1_R1240_U219 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1240_U220 = ~new_P1_R1240_U45;
  assign new_P1_R1240_U221 = new_P1_U3464 | new_P1_U3060;
  assign new_P1_R1240_U222 = ~new_P1_R1240_U221 | ~new_P1_R1240_U45;
  assign new_P1_R1240_U223 = ~new_P1_R1240_U123 | ~new_P1_R1240_U222;
  assign new_P1_R1240_U224 = ~new_P1_R1240_U220 | ~new_P1_R1240_U35;
  assign new_P1_R1240_U225 = ~new_P1_U3467 | ~new_P1_U3067;
  assign new_P1_R1240_U226 = ~new_P1_R1240_U124 | ~new_P1_R1240_U224;
  assign new_P1_R1240_U227 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1240_U228 = ~new_P1_R1240_U183 | ~new_P1_R1240_U180;
  assign new_P1_R1240_U229 = ~new_P1_R1240_U144;
  assign new_P1_R1240_U230 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1240_U231 = ~new_P1_R1240_U43 | ~new_P1_R1240_U44 | ~new_P1_R1240_U400 | ~new_P1_R1240_U399;
  assign new_P1_R1240_U232 = ~new_P1_R1240_U44 | ~new_P1_R1240_U43;
  assign new_P1_R1240_U233 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1240_U234 = ~new_P1_R1240_U125 | ~new_P1_R1240_U232;
  assign new_P1_R1240_U235 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1240_U236 = new_P1_U3062 | new_P1_U3482;
  assign new_P1_R1240_U237 = ~new_P1_R1240_U176 | ~new_P1_R1240_U7;
  assign new_P1_R1240_U238 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1240_U239 = ~new_P1_R1240_U127 | ~new_P1_R1240_U237;
  assign new_P1_R1240_U240 = new_P1_U3482 | new_P1_U3062;
  assign new_P1_R1240_U241 = ~new_P1_R1240_U126 | ~new_P1_R1240_U143;
  assign new_P1_R1240_U242 = ~new_P1_R1240_U240 | ~new_P1_R1240_U239;
  assign new_P1_R1240_U243 = ~new_P1_R1240_U166;
  assign new_P1_R1240_U244 = new_P1_U3080 | new_P1_U3491;
  assign new_P1_R1240_U245 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1240_U246 = ~new_P1_R1240_U173 | ~new_P1_R1240_U8;
  assign new_P1_R1240_U247 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1240_U248 = ~new_P1_R1240_U129 | ~new_P1_R1240_U246;
  assign new_P1_R1240_U249 = new_P1_U3485 | new_P1_U3063;
  assign new_P1_R1240_U250 = new_P1_U3491 | new_P1_U3080;
  assign new_P1_R1240_U251 = ~new_P1_R1240_U128 | ~new_P1_R1240_U166;
  assign new_P1_R1240_U252 = ~new_P1_R1240_U250 | ~new_P1_R1240_U248;
  assign new_P1_R1240_U253 = ~new_P1_R1240_U165;
  assign new_P1_R1240_U254 = new_P1_U3494 | new_P1_U3079;
  assign new_P1_R1240_U255 = ~new_P1_R1240_U254 | ~new_P1_R1240_U165;
  assign new_P1_R1240_U256 = ~new_P1_U3079 | ~new_P1_U3494;
  assign new_P1_R1240_U257 = ~new_P1_R1240_U163;
  assign new_P1_R1240_U258 = new_P1_U3497 | new_P1_U3074;
  assign new_P1_R1240_U259 = ~new_P1_R1240_U258 | ~new_P1_R1240_U163;
  assign new_P1_R1240_U260 = ~new_P1_U3074 | ~new_P1_U3497;
  assign new_P1_R1240_U261 = ~new_P1_R1240_U93;
  assign new_P1_R1240_U262 = new_P1_U3069 | new_P1_U3503;
  assign new_P1_R1240_U263 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1240_U264 = ~new_P1_R1240_U60;
  assign new_P1_R1240_U265 = ~new_P1_R1240_U61 | ~new_P1_R1240_U60;
  assign new_P1_R1240_U266 = ~new_P1_U3069 | ~new_P1_R1240_U265;
  assign new_P1_R1240_U267 = ~new_P1_U3503 | ~new_P1_R1240_U264;
  assign new_P1_R1240_U268 = ~new_P1_R1240_U9 | ~new_P1_R1240_U93;
  assign new_P1_R1240_U269 = ~new_P1_R1240_U161;
  assign new_P1_R1240_U270 = new_P1_U3076 | new_P1_U3982;
  assign new_P1_R1240_U271 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1240_U272 = new_P1_U3075 | new_P1_U3981;
  assign new_P1_R1240_U273 = ~new_P1_R1240_U81;
  assign new_P1_R1240_U274 = ~new_P1_U3982 | ~new_P1_R1240_U273;
  assign new_P1_R1240_U275 = ~new_P1_R1240_U274 | ~new_P1_R1240_U91;
  assign new_P1_R1240_U276 = ~new_P1_R1240_U81 | ~new_P1_R1240_U82;
  assign new_P1_R1240_U277 = ~new_P1_R1240_U276 | ~new_P1_R1240_U275;
  assign new_P1_R1240_U278 = ~new_P1_R1240_U174 | ~new_P1_R1240_U10;
  assign new_P1_R1240_U279 = ~new_P1_U3075 | ~new_P1_U3981;
  assign new_P1_R1240_U280 = ~new_P1_R1240_U277 | ~new_P1_R1240_U278;
  assign new_P1_R1240_U281 = new_P1_U3506 | new_P1_U3082;
  assign new_P1_R1240_U282 = new_P1_U3981 | new_P1_U3075;
  assign new_P1_R1240_U283 = ~new_P1_R1240_U131 | ~new_P1_R1240_U272 | ~new_P1_R1240_U161;
  assign new_P1_R1240_U284 = ~new_P1_R1240_U282 | ~new_P1_R1240_U280;
  assign new_P1_R1240_U285 = ~new_P1_R1240_U158;
  assign new_P1_R1240_U286 = new_P1_U3980 | new_P1_U3061;
  assign new_P1_R1240_U287 = ~new_P1_R1240_U286 | ~new_P1_R1240_U158;
  assign new_P1_R1240_U288 = ~new_P1_U3061 | ~new_P1_U3980;
  assign new_P1_R1240_U289 = ~new_P1_R1240_U156;
  assign new_P1_R1240_U290 = new_P1_U3979 | new_P1_U3066;
  assign new_P1_R1240_U291 = ~new_P1_R1240_U290 | ~new_P1_R1240_U156;
  assign new_P1_R1240_U292 = ~new_P1_U3066 | ~new_P1_U3979;
  assign new_P1_R1240_U293 = ~new_P1_R1240_U154;
  assign new_P1_R1240_U294 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1240_U295 = ~new_P1_R1240_U175 | ~new_P1_R1240_U172;
  assign new_P1_R1240_U296 = ~new_P1_R1240_U87;
  assign new_P1_R1240_U297 = new_P1_U3978 | new_P1_U3065;
  assign new_P1_R1240_U298 = ~new_P1_R1240_U167 | ~new_P1_R1240_U154 | ~new_P1_R1240_U297;
  assign new_P1_R1240_U299 = ~new_P1_R1240_U152;
  assign new_P1_R1240_U300 = new_P1_U3975 | new_P1_U3053;
  assign new_P1_R1240_U301 = ~new_P1_U3053 | ~new_P1_U3975;
  assign new_P1_R1240_U302 = ~new_P1_R1240_U150;
  assign new_P1_R1240_U303 = ~new_P1_U3974 | ~new_P1_R1240_U150;
  assign new_P1_R1240_U304 = ~new_P1_R1240_U148;
  assign new_P1_R1240_U305 = ~new_P1_R1240_U297 | ~new_P1_R1240_U154;
  assign new_P1_R1240_U306 = ~new_P1_R1240_U90;
  assign new_P1_R1240_U307 = new_P1_U3977 | new_P1_U3058;
  assign new_P1_R1240_U308 = ~new_P1_R1240_U307 | ~new_P1_R1240_U90;
  assign new_P1_R1240_U309 = ~new_P1_R1240_U153 | ~new_P1_R1240_U308 | ~new_P1_R1240_U172;
  assign new_P1_R1240_U310 = ~new_P1_R1240_U306 | ~new_P1_R1240_U172;
  assign new_P1_R1240_U311 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1240_U312 = ~new_P1_R1240_U167 | ~new_P1_R1240_U310 | ~new_P1_R1240_U311;
  assign new_P1_R1240_U313 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1240_U314 = ~new_P1_R1240_U281 | ~new_P1_R1240_U161;
  assign new_P1_R1240_U315 = ~new_P1_R1240_U92;
  assign new_P1_R1240_U316 = ~new_P1_R1240_U10 | ~new_P1_R1240_U92;
  assign new_P1_R1240_U317 = ~new_P1_R1240_U135 | ~new_P1_R1240_U316;
  assign new_P1_R1240_U318 = ~new_P1_R1240_U316 | ~new_P1_R1240_U277;
  assign new_P1_R1240_U319 = ~new_P1_R1240_U452 | ~new_P1_R1240_U318;
  assign new_P1_R1240_U320 = new_P1_U3508 | new_P1_U3081;
  assign new_P1_R1240_U321 = ~new_P1_R1240_U320 | ~new_P1_R1240_U92;
  assign new_P1_R1240_U322 = ~new_P1_R1240_U136 | ~new_P1_R1240_U321;
  assign new_P1_R1240_U323 = ~new_P1_R1240_U315 | ~new_P1_R1240_U81;
  assign new_P1_R1240_U324 = ~new_P1_U3076 | ~new_P1_U3982;
  assign new_P1_R1240_U325 = ~new_P1_R1240_U10 | ~new_P1_R1240_U324 | ~new_P1_R1240_U323;
  assign new_P1_R1240_U326 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1240_U327 = ~new_P1_R1240_U160;
  assign new_P1_R1240_U328 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1240_U329 = new_P1_U3500 | new_P1_U3073;
  assign new_P1_R1240_U330 = ~new_P1_R1240_U329 | ~new_P1_R1240_U93;
  assign new_P1_R1240_U331 = ~new_P1_R1240_U137 | ~new_P1_R1240_U330;
  assign new_P1_R1240_U332 = ~new_P1_R1240_U261 | ~new_P1_R1240_U60;
  assign new_P1_R1240_U333 = ~new_P1_U3503 | ~new_P1_U3069;
  assign new_P1_R1240_U334 = ~new_P1_R1240_U138 | ~new_P1_R1240_U332;
  assign new_P1_R1240_U335 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1240_U336 = ~new_P1_R1240_U249 | ~new_P1_R1240_U166;
  assign new_P1_R1240_U337 = ~new_P1_R1240_U94;
  assign new_P1_R1240_U338 = new_P1_U3488 | new_P1_U3072;
  assign new_P1_R1240_U339 = ~new_P1_R1240_U338 | ~new_P1_R1240_U94;
  assign new_P1_R1240_U340 = ~new_P1_R1240_U139 | ~new_P1_R1240_U339;
  assign new_P1_R1240_U341 = ~new_P1_R1240_U337 | ~new_P1_R1240_U171;
  assign new_P1_R1240_U342 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1240_U343 = ~new_P1_R1240_U140 | ~new_P1_R1240_U341;
  assign new_P1_R1240_U344 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1240_U345 = new_P1_U3479 | new_P1_U3083;
  assign new_P1_R1240_U346 = ~new_P1_R1240_U345 | ~new_P1_R1240_U41;
  assign new_P1_R1240_U347 = ~new_P1_R1240_U141 | ~new_P1_R1240_U346;
  assign new_P1_R1240_U348 = ~new_P1_R1240_U205 | ~new_P1_R1240_U170;
  assign new_P1_R1240_U349 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1240_U350 = ~new_P1_R1240_U142 | ~new_P1_R1240_U348;
  assign new_P1_R1240_U351 = ~new_P1_R1240_U206 | ~new_P1_R1240_U170;
  assign new_P1_R1240_U352 = ~new_P1_R1240_U203 | ~new_P1_R1240_U62;
  assign new_P1_R1240_U353 = ~new_P1_R1240_U213 | ~new_P1_R1240_U23;
  assign new_P1_R1240_U354 = ~new_P1_R1240_U227 | ~new_P1_R1240_U35;
  assign new_P1_R1240_U355 = ~new_P1_R1240_U230 | ~new_P1_R1240_U179;
  assign new_P1_R1240_U356 = ~new_P1_R1240_U313 | ~new_P1_R1240_U172;
  assign new_P1_R1240_U357 = ~new_P1_R1240_U297 | ~new_P1_R1240_U175;
  assign new_P1_R1240_U358 = ~new_P1_R1240_U328 | ~new_P1_R1240_U81;
  assign new_P1_R1240_U359 = ~new_P1_R1240_U281 | ~new_P1_R1240_U78;
  assign new_P1_R1240_U360 = ~new_P1_R1240_U335 | ~new_P1_R1240_U60;
  assign new_P1_R1240_U361 = ~new_P1_R1240_U344 | ~new_P1_R1240_U171;
  assign new_P1_R1240_U362 = ~new_P1_R1240_U249 | ~new_P1_R1240_U69;
  assign new_P1_R1240_U363 = ~new_P1_U3974 | ~new_P1_U3054;
  assign new_P1_R1240_U364 = ~new_P1_R1240_U295 | ~new_P1_R1240_U167;
  assign new_P1_R1240_U365 = ~new_P1_U3057 | ~new_P1_R1240_U294;
  assign new_P1_R1240_U366 = ~new_P1_U3976 | ~new_P1_R1240_U294;
  assign new_P1_R1240_U367 = ~new_P1_R1240_U300 | ~new_P1_R1240_U295 | ~new_P1_R1240_U167;
  assign new_P1_R1240_U368 = ~new_P1_R1240_U133 | ~new_P1_R1240_U154 | ~new_P1_R1240_U167;
  assign new_P1_R1240_U369 = ~new_P1_R1240_U296 | ~new_P1_R1240_U300;
  assign new_P1_R1240_U370 = ~new_P1_U3083 | ~new_P1_R1240_U40;
  assign new_P1_R1240_U371 = ~new_P1_U3479 | ~new_P1_R1240_U39;
  assign new_P1_R1240_U372 = ~new_P1_R1240_U371 | ~new_P1_R1240_U370;
  assign new_P1_R1240_U373 = ~new_P1_R1240_U351 | ~new_P1_R1240_U41;
  assign new_P1_R1240_U374 = ~new_P1_R1240_U372 | ~new_P1_R1240_U205;
  assign new_P1_R1240_U375 = ~new_P1_U3084 | ~new_P1_R1240_U37;
  assign new_P1_R1240_U376 = ~new_P1_U3476 | ~new_P1_R1240_U38;
  assign new_P1_R1240_U377 = ~new_P1_R1240_U376 | ~new_P1_R1240_U375;
  assign new_P1_R1240_U378 = ~new_P1_R1240_U352 | ~new_P1_R1240_U143;
  assign new_P1_R1240_U379 = ~new_P1_R1240_U202 | ~new_P1_R1240_U377;
  assign new_P1_R1240_U380 = ~new_P1_U3070 | ~new_P1_R1240_U24;
  assign new_P1_R1240_U381 = ~new_P1_U3473 | ~new_P1_R1240_U22;
  assign new_P1_R1240_U382 = ~new_P1_U3071 | ~new_P1_R1240_U20;
  assign new_P1_R1240_U383 = ~new_P1_U3470 | ~new_P1_R1240_U21;
  assign new_P1_R1240_U384 = ~new_P1_R1240_U383 | ~new_P1_R1240_U382;
  assign new_P1_R1240_U385 = ~new_P1_R1240_U353 | ~new_P1_R1240_U42;
  assign new_P1_R1240_U386 = ~new_P1_R1240_U384 | ~new_P1_R1240_U194;
  assign new_P1_R1240_U387 = ~new_P1_U3067 | ~new_P1_R1240_U36;
  assign new_P1_R1240_U388 = ~new_P1_U3467 | ~new_P1_R1240_U27;
  assign new_P1_R1240_U389 = ~new_P1_U3060 | ~new_P1_R1240_U25;
  assign new_P1_R1240_U390 = ~new_P1_U3464 | ~new_P1_R1240_U26;
  assign new_P1_R1240_U391 = ~new_P1_R1240_U390 | ~new_P1_R1240_U389;
  assign new_P1_R1240_U392 = ~new_P1_R1240_U354 | ~new_P1_R1240_U45;
  assign new_P1_R1240_U393 = ~new_P1_R1240_U391 | ~new_P1_R1240_U220;
  assign new_P1_R1240_U394 = ~new_P1_U3064 | ~new_P1_R1240_U33;
  assign new_P1_R1240_U395 = ~new_P1_U3461 | ~new_P1_R1240_U34;
  assign new_P1_R1240_U396 = ~new_P1_R1240_U395 | ~new_P1_R1240_U394;
  assign new_P1_R1240_U397 = ~new_P1_R1240_U355 | ~new_P1_R1240_U144;
  assign new_P1_R1240_U398 = ~new_P1_R1240_U229 | ~new_P1_R1240_U396;
  assign new_P1_R1240_U399 = ~new_P1_U3068 | ~new_P1_R1240_U28;
  assign new_P1_R1240_U400 = ~new_P1_U3458 | ~new_P1_R1240_U29;
  assign new_P1_R1240_U401 = ~new_P1_U3055 | ~new_P1_R1240_U146;
  assign new_P1_R1240_U402 = ~new_P1_U3985 | ~new_P1_R1240_U145;
  assign new_P1_R1240_U403 = ~new_P1_U3055 | ~new_P1_R1240_U146;
  assign new_P1_R1240_U404 = ~new_P1_U3985 | ~new_P1_R1240_U145;
  assign new_P1_R1240_U405 = ~new_P1_R1240_U404 | ~new_P1_R1240_U403;
  assign new_P1_R1240_U406 = ~new_P1_R1240_U147 | ~new_P1_R1240_U148;
  assign new_P1_R1240_U407 = ~new_P1_R1240_U304 | ~new_P1_R1240_U405;
  assign new_P1_R1240_U408 = ~new_P1_U3054 | ~new_P1_R1240_U89;
  assign new_P1_R1240_U409 = ~new_P1_U3974 | ~new_P1_R1240_U88;
  assign new_P1_R1240_U410 = ~new_P1_U3054 | ~new_P1_R1240_U89;
  assign new_P1_R1240_U411 = ~new_P1_U3974 | ~new_P1_R1240_U88;
  assign new_P1_R1240_U412 = ~new_P1_R1240_U411 | ~new_P1_R1240_U410;
  assign new_P1_R1240_U413 = ~new_P1_R1240_U149 | ~new_P1_R1240_U150;
  assign new_P1_R1240_U414 = ~new_P1_R1240_U302 | ~new_P1_R1240_U412;
  assign new_P1_R1240_U415 = ~new_P1_U3053 | ~new_P1_R1240_U47;
  assign new_P1_R1240_U416 = ~new_P1_U3975 | ~new_P1_R1240_U48;
  assign new_P1_R1240_U417 = ~new_P1_U3053 | ~new_P1_R1240_U47;
  assign new_P1_R1240_U418 = ~new_P1_U3975 | ~new_P1_R1240_U48;
  assign new_P1_R1240_U419 = ~new_P1_R1240_U418 | ~new_P1_R1240_U417;
  assign new_P1_R1240_U420 = ~new_P1_R1240_U151 | ~new_P1_R1240_U152;
  assign new_P1_R1240_U421 = ~new_P1_R1240_U299 | ~new_P1_R1240_U419;
  assign new_P1_R1240_U422 = ~new_P1_U3057 | ~new_P1_R1240_U50;
  assign new_P1_R1240_U423 = ~new_P1_U3976 | ~new_P1_R1240_U49;
  assign new_P1_R1240_U424 = ~new_P1_U3058 | ~new_P1_R1240_U51;
  assign new_P1_R1240_U425 = ~new_P1_U3977 | ~new_P1_R1240_U52;
  assign new_P1_R1240_U426 = ~new_P1_R1240_U425 | ~new_P1_R1240_U424;
  assign new_P1_R1240_U427 = ~new_P1_R1240_U356 | ~new_P1_R1240_U90;
  assign new_P1_R1240_U428 = ~new_P1_R1240_U426 | ~new_P1_R1240_U306;
  assign new_P1_R1240_U429 = ~new_P1_U3065 | ~new_P1_R1240_U53;
  assign new_P1_R1240_U430 = ~new_P1_U3978 | ~new_P1_R1240_U54;
  assign new_P1_R1240_U431 = ~new_P1_R1240_U430 | ~new_P1_R1240_U429;
  assign new_P1_R1240_U432 = ~new_P1_R1240_U357 | ~new_P1_R1240_U154;
  assign new_P1_R1240_U433 = ~new_P1_R1240_U293 | ~new_P1_R1240_U431;
  assign new_P1_R1240_U434 = ~new_P1_U3066 | ~new_P1_R1240_U85;
  assign new_P1_R1240_U435 = ~new_P1_U3979 | ~new_P1_R1240_U86;
  assign new_P1_R1240_U436 = ~new_P1_U3066 | ~new_P1_R1240_U85;
  assign new_P1_R1240_U437 = ~new_P1_U3979 | ~new_P1_R1240_U86;
  assign new_P1_R1240_U438 = ~new_P1_R1240_U437 | ~new_P1_R1240_U436;
  assign new_P1_R1240_U439 = ~new_P1_R1240_U155 | ~new_P1_R1240_U156;
  assign new_P1_R1240_U440 = ~new_P1_R1240_U289 | ~new_P1_R1240_U438;
  assign new_P1_R1240_U441 = ~new_P1_U3061 | ~new_P1_R1240_U83;
  assign new_P1_R1240_U442 = ~new_P1_U3980 | ~new_P1_R1240_U84;
  assign new_P1_R1240_U443 = ~new_P1_U3061 | ~new_P1_R1240_U83;
  assign new_P1_R1240_U444 = ~new_P1_U3980 | ~new_P1_R1240_U84;
  assign new_P1_R1240_U445 = ~new_P1_R1240_U444 | ~new_P1_R1240_U443;
  assign new_P1_R1240_U446 = ~new_P1_R1240_U157 | ~new_P1_R1240_U158;
  assign new_P1_R1240_U447 = ~new_P1_R1240_U285 | ~new_P1_R1240_U445;
  assign new_P1_R1240_U448 = ~new_P1_U3075 | ~new_P1_R1240_U55;
  assign new_P1_R1240_U449 = ~new_P1_U3981 | ~new_P1_R1240_U56;
  assign new_P1_R1240_U450 = ~new_P1_U3075 | ~new_P1_R1240_U55;
  assign new_P1_R1240_U451 = ~new_P1_U3981 | ~new_P1_R1240_U56;
  assign new_P1_R1240_U452 = ~new_P1_R1240_U451 | ~new_P1_R1240_U450;
  assign new_P1_R1240_U453 = ~new_P1_U3076 | ~new_P1_R1240_U82;
  assign new_P1_R1240_U454 = ~new_P1_U3982 | ~new_P1_R1240_U91;
  assign new_P1_R1240_U455 = ~new_P1_R1240_U181 | ~new_P1_R1240_U160;
  assign new_P1_R1240_U456 = ~new_P1_R1240_U327 | ~new_P1_R1240_U32;
  assign new_P1_R1240_U457 = ~new_P1_U3081 | ~new_P1_R1240_U79;
  assign new_P1_R1240_U458 = ~new_P1_U3508 | ~new_P1_R1240_U80;
  assign new_P1_R1240_U459 = ~new_P1_R1240_U458 | ~new_P1_R1240_U457;
  assign new_P1_R1240_U460 = ~new_P1_R1240_U358 | ~new_P1_R1240_U92;
  assign new_P1_R1240_U461 = ~new_P1_R1240_U459 | ~new_P1_R1240_U315;
  assign new_P1_R1240_U462 = ~new_P1_U3082 | ~new_P1_R1240_U76;
  assign new_P1_R1240_U463 = ~new_P1_U3506 | ~new_P1_R1240_U77;
  assign new_P1_R1240_U464 = ~new_P1_R1240_U463 | ~new_P1_R1240_U462;
  assign new_P1_R1240_U465 = ~new_P1_R1240_U359 | ~new_P1_R1240_U161;
  assign new_P1_R1240_U466 = ~new_P1_R1240_U269 | ~new_P1_R1240_U464;
  assign new_P1_R1240_U467 = ~new_P1_U3069 | ~new_P1_R1240_U61;
  assign new_P1_R1240_U468 = ~new_P1_U3503 | ~new_P1_R1240_U59;
  assign new_P1_R1240_U469 = ~new_P1_U3073 | ~new_P1_R1240_U57;
  assign new_P1_R1240_U470 = ~new_P1_U3500 | ~new_P1_R1240_U58;
  assign new_P1_R1240_U471 = ~new_P1_R1240_U470 | ~new_P1_R1240_U469;
  assign new_P1_R1240_U472 = ~new_P1_R1240_U360 | ~new_P1_R1240_U93;
  assign new_P1_R1240_U473 = ~new_P1_R1240_U471 | ~new_P1_R1240_U261;
  assign new_P1_R1240_U474 = ~new_P1_U3074 | ~new_P1_R1240_U74;
  assign new_P1_R1240_U475 = ~new_P1_U3497 | ~new_P1_R1240_U75;
  assign new_P1_R1240_U476 = ~new_P1_U3074 | ~new_P1_R1240_U74;
  assign new_P1_R1240_U477 = ~new_P1_U3497 | ~new_P1_R1240_U75;
  assign new_P1_R1240_U478 = ~new_P1_R1240_U477 | ~new_P1_R1240_U476;
  assign new_P1_R1240_U479 = ~new_P1_R1240_U162 | ~new_P1_R1240_U163;
  assign new_P1_R1240_U480 = ~new_P1_R1240_U257 | ~new_P1_R1240_U478;
  assign new_P1_R1240_U481 = ~new_P1_U3079 | ~new_P1_R1240_U72;
  assign new_P1_R1240_U482 = ~new_P1_U3494 | ~new_P1_R1240_U73;
  assign new_P1_R1240_U483 = ~new_P1_U3079 | ~new_P1_R1240_U72;
  assign new_P1_R1240_U484 = ~new_P1_U3494 | ~new_P1_R1240_U73;
  assign new_P1_R1240_U485 = ~new_P1_R1240_U484 | ~new_P1_R1240_U483;
  assign new_P1_R1240_U486 = ~new_P1_R1240_U164 | ~new_P1_R1240_U165;
  assign new_P1_R1240_U487 = ~new_P1_R1240_U253 | ~new_P1_R1240_U485;
  assign new_P1_R1240_U488 = ~new_P1_U3080 | ~new_P1_R1240_U70;
  assign new_P1_R1240_U489 = ~new_P1_U3491 | ~new_P1_R1240_U71;
  assign new_P1_R1240_U490 = ~new_P1_U3072 | ~new_P1_R1240_U65;
  assign new_P1_R1240_U491 = ~new_P1_U3488 | ~new_P1_R1240_U66;
  assign new_P1_R1240_U492 = ~new_P1_R1240_U491 | ~new_P1_R1240_U490;
  assign new_P1_R1240_U493 = ~new_P1_R1240_U361 | ~new_P1_R1240_U94;
  assign new_P1_R1240_U494 = ~new_P1_R1240_U492 | ~new_P1_R1240_U337;
  assign new_P1_R1240_U495 = ~new_P1_U3063 | ~new_P1_R1240_U67;
  assign new_P1_R1240_U496 = ~new_P1_U3485 | ~new_P1_R1240_U68;
  assign new_P1_R1240_U497 = ~new_P1_R1240_U496 | ~new_P1_R1240_U495;
  assign new_P1_R1240_U498 = ~new_P1_R1240_U362 | ~new_P1_R1240_U166;
  assign new_P1_R1240_U499 = ~new_P1_R1240_U243 | ~new_P1_R1240_U497;
  assign new_P1_R1240_U500 = ~new_P1_U3062 | ~new_P1_R1240_U63;
  assign new_P1_R1240_U501 = ~new_P1_U3482 | ~new_P1_R1240_U64;
  assign new_P1_R1240_U502 = ~new_P1_U3077 | ~new_P1_R1240_U30;
  assign new_P1_R1240_U503 = ~new_P1_U3450 | ~new_P1_R1240_U31;
  assign new_P1_R1162_U4 = new_P1_R1162_U95 & new_P1_R1162_U94;
  assign new_P1_R1162_U5 = new_P1_R1162_U96 & new_P1_R1162_U97;
  assign new_P1_R1162_U6 = new_P1_R1162_U113 & new_P1_R1162_U112;
  assign new_P1_R1162_U7 = new_P1_R1162_U155 & new_P1_R1162_U154;
  assign new_P1_R1162_U8 = new_P1_R1162_U164 & new_P1_R1162_U163;
  assign new_P1_R1162_U9 = new_P1_R1162_U182 & new_P1_R1162_U181;
  assign new_P1_R1162_U10 = new_P1_R1162_U218 & new_P1_R1162_U215;
  assign new_P1_R1162_U11 = new_P1_R1162_U211 & new_P1_R1162_U208;
  assign new_P1_R1162_U12 = new_P1_R1162_U202 & new_P1_R1162_U199;
  assign new_P1_R1162_U13 = new_P1_R1162_U196 & new_P1_R1162_U192;
  assign new_P1_R1162_U14 = new_P1_R1162_U151 & new_P1_R1162_U148;
  assign new_P1_R1162_U15 = new_P1_R1162_U143 & new_P1_R1162_U140;
  assign new_P1_R1162_U16 = new_P1_R1162_U129 & new_P1_R1162_U126;
  assign new_P1_R1162_U17 = ~P1_REG1_REG_6_;
  assign new_P1_R1162_U18 = ~new_P1_U3469;
  assign new_P1_R1162_U19 = ~new_P1_U3472;
  assign new_P1_R1162_U20 = ~new_P1_U3469 | ~P1_REG1_REG_6_;
  assign new_P1_R1162_U21 = ~P1_REG1_REG_7_;
  assign new_P1_R1162_U22 = ~P1_REG1_REG_4_;
  assign new_P1_R1162_U23 = ~new_P1_U3463;
  assign new_P1_R1162_U24 = ~new_P1_U3466;
  assign new_P1_R1162_U25 = ~P1_REG1_REG_2_;
  assign new_P1_R1162_U26 = ~new_P1_U3457;
  assign new_P1_R1162_U27 = ~P1_REG1_REG_0_;
  assign new_P1_R1162_U28 = ~new_P1_U3448;
  assign new_P1_R1162_U29 = ~new_P1_U3448 | ~P1_REG1_REG_0_;
  assign new_P1_R1162_U30 = ~P1_REG1_REG_3_;
  assign new_P1_R1162_U31 = ~new_P1_U3460;
  assign new_P1_R1162_U32 = ~new_P1_U3463 | ~P1_REG1_REG_4_;
  assign new_P1_R1162_U33 = ~P1_REG1_REG_5_;
  assign new_P1_R1162_U34 = ~P1_REG1_REG_8_;
  assign new_P1_R1162_U35 = ~new_P1_U3475;
  assign new_P1_R1162_U36 = ~new_P1_U3478;
  assign new_P1_R1162_U37 = ~P1_REG1_REG_9_;
  assign new_P1_R1162_U38 = ~new_P1_R1162_U49 | ~new_P1_R1162_U121;
  assign new_P1_R1162_U39 = ~new_P1_R1162_U109 | ~new_P1_R1162_U110 | ~new_P1_R1162_U108;
  assign new_P1_R1162_U40 = ~new_P1_R1162_U98 | ~new_P1_R1162_U99;
  assign new_P1_R1162_U41 = ~P1_REG1_REG_1_ | ~new_P1_U3454;
  assign new_P1_R1162_U42 = ~new_P1_R1162_U135 | ~new_P1_R1162_U136 | ~new_P1_R1162_U134;
  assign new_P1_R1162_U43 = ~new_P1_R1162_U132 | ~new_P1_R1162_U131;
  assign new_P1_R1162_U44 = ~P1_REG1_REG_16_;
  assign new_P1_R1162_U45 = ~new_P1_U3499;
  assign new_P1_R1162_U46 = ~new_P1_U3502;
  assign new_P1_R1162_U47 = ~new_P1_U3499 | ~P1_REG1_REG_16_;
  assign new_P1_R1162_U48 = ~P1_REG1_REG_17_;
  assign new_P1_R1162_U49 = ~new_P1_U3475 | ~P1_REG1_REG_8_;
  assign new_P1_R1162_U50 = ~P1_REG1_REG_10_;
  assign new_P1_R1162_U51 = ~new_P1_U3481;
  assign new_P1_R1162_U52 = ~P1_REG1_REG_12_;
  assign new_P1_R1162_U53 = ~new_P1_U3487;
  assign new_P1_R1162_U54 = ~P1_REG1_REG_11_;
  assign new_P1_R1162_U55 = ~new_P1_U3484;
  assign new_P1_R1162_U56 = ~new_P1_U3484 | ~P1_REG1_REG_11_;
  assign new_P1_R1162_U57 = ~P1_REG1_REG_13_;
  assign new_P1_R1162_U58 = ~new_P1_U3490;
  assign new_P1_R1162_U59 = ~P1_REG1_REG_14_;
  assign new_P1_R1162_U60 = ~new_P1_U3493;
  assign new_P1_R1162_U61 = ~P1_REG1_REG_15_;
  assign new_P1_R1162_U62 = ~new_P1_U3496;
  assign new_P1_R1162_U63 = ~P1_REG1_REG_18_;
  assign new_P1_R1162_U64 = ~new_P1_U3505;
  assign new_P1_R1162_U65 = ~new_P1_R1162_U187 | ~new_P1_R1162_U186 | ~new_P1_R1162_U185;
  assign new_P1_R1162_U66 = ~new_P1_R1162_U179 | ~new_P1_R1162_U178;
  assign new_P1_R1162_U67 = ~new_P1_R1162_U56 | ~new_P1_R1162_U204;
  assign new_P1_R1162_U68 = ~new_P1_R1162_U259 | ~new_P1_R1162_U258;
  assign new_P1_R1162_U69 = ~new_P1_R1162_U308 | ~new_P1_R1162_U307;
  assign new_P1_R1162_U70 = ~new_P1_R1162_U231 | ~new_P1_R1162_U230;
  assign new_P1_R1162_U71 = ~new_P1_R1162_U236 | ~new_P1_R1162_U235;
  assign new_P1_R1162_U72 = ~new_P1_R1162_U243 | ~new_P1_R1162_U242;
  assign new_P1_R1162_U73 = ~new_P1_R1162_U250 | ~new_P1_R1162_U249;
  assign new_P1_R1162_U74 = ~new_P1_R1162_U255 | ~new_P1_R1162_U254;
  assign new_P1_R1162_U75 = ~new_P1_R1162_U271 | ~new_P1_R1162_U270;
  assign new_P1_R1162_U76 = ~new_P1_R1162_U278 | ~new_P1_R1162_U277;
  assign new_P1_R1162_U77 = ~new_P1_R1162_U285 | ~new_P1_R1162_U284;
  assign new_P1_R1162_U78 = ~new_P1_R1162_U292 | ~new_P1_R1162_U291;
  assign new_P1_R1162_U79 = ~new_P1_R1162_U299 | ~new_P1_R1162_U298;
  assign new_P1_R1162_U80 = ~new_P1_R1162_U304 | ~new_P1_R1162_U303;
  assign new_P1_R1162_U81 = ~new_P1_R1162_U118 | ~new_P1_R1162_U117 | ~new_P1_R1162_U116;
  assign new_P1_R1162_U82 = ~new_P1_R1162_U133 | ~new_P1_R1162_U145;
  assign new_P1_R1162_U83 = ~new_P1_R1162_U41 | ~new_P1_R1162_U152;
  assign new_P1_R1162_U84 = ~new_P1_U3442;
  assign new_P1_R1162_U85 = ~P1_REG1_REG_19_;
  assign new_P1_R1162_U86 = ~new_P1_R1162_U175 | ~new_P1_R1162_U174;
  assign new_P1_R1162_U87 = ~new_P1_R1162_U171 | ~new_P1_R1162_U170;
  assign new_P1_R1162_U88 = ~new_P1_R1162_U161 | ~new_P1_R1162_U160;
  assign new_P1_R1162_U89 = ~new_P1_R1162_U32;
  assign new_P1_R1162_U90 = ~P1_REG1_REG_9_ | ~new_P1_U3478;
  assign new_P1_R1162_U91 = ~new_P1_U3487 | ~P1_REG1_REG_12_;
  assign new_P1_R1162_U92 = ~new_P1_R1162_U56;
  assign new_P1_R1162_U93 = ~new_P1_R1162_U49;
  assign new_P1_R1162_U94 = new_P1_U3466 | P1_REG1_REG_5_;
  assign new_P1_R1162_U95 = new_P1_U3463 | P1_REG1_REG_4_;
  assign new_P1_R1162_U96 = P1_REG1_REG_3_ | new_P1_U3460;
  assign new_P1_R1162_U97 = P1_REG1_REG_2_ | new_P1_U3457;
  assign new_P1_R1162_U98 = ~new_P1_R1162_U29;
  assign new_P1_R1162_U99 = P1_REG1_REG_1_ | new_P1_U3454;
  assign new_P1_R1162_U100 = ~new_P1_R1162_U40;
  assign new_P1_R1162_U101 = ~new_P1_R1162_U41;
  assign new_P1_R1162_U102 = ~new_P1_R1162_U40 | ~new_P1_R1162_U41;
  assign new_P1_R1162_U103 = ~new_P1_R1162_U96 | ~P1_REG1_REG_2_ | ~new_P1_U3457;
  assign new_P1_R1162_U104 = ~new_P1_R1162_U5 | ~new_P1_R1162_U102;
  assign new_P1_R1162_U105 = ~new_P1_U3460 | ~P1_REG1_REG_3_;
  assign new_P1_R1162_U106 = ~new_P1_R1162_U104 | ~new_P1_R1162_U105 | ~new_P1_R1162_U103;
  assign new_P1_R1162_U107 = ~new_P1_R1162_U33 | ~new_P1_R1162_U32;
  assign new_P1_R1162_U108 = ~new_P1_U3466 | ~new_P1_R1162_U107;
  assign new_P1_R1162_U109 = ~new_P1_R1162_U4 | ~new_P1_R1162_U106;
  assign new_P1_R1162_U110 = ~P1_REG1_REG_5_ | ~new_P1_R1162_U89;
  assign new_P1_R1162_U111 = ~new_P1_R1162_U39;
  assign new_P1_R1162_U112 = new_P1_U3472 | P1_REG1_REG_7_;
  assign new_P1_R1162_U113 = new_P1_U3469 | P1_REG1_REG_6_;
  assign new_P1_R1162_U114 = ~new_P1_R1162_U20;
  assign new_P1_R1162_U115 = ~new_P1_R1162_U21 | ~new_P1_R1162_U20;
  assign new_P1_R1162_U116 = ~new_P1_U3472 | ~new_P1_R1162_U115;
  assign new_P1_R1162_U117 = ~P1_REG1_REG_7_ | ~new_P1_R1162_U114;
  assign new_P1_R1162_U118 = ~new_P1_R1162_U6 | ~new_P1_R1162_U39;
  assign new_P1_R1162_U119 = ~new_P1_R1162_U81;
  assign new_P1_R1162_U120 = P1_REG1_REG_8_ | new_P1_U3475;
  assign new_P1_R1162_U121 = ~new_P1_R1162_U120 | ~new_P1_R1162_U81;
  assign new_P1_R1162_U122 = ~new_P1_R1162_U38;
  assign new_P1_R1162_U123 = new_P1_U3478 | P1_REG1_REG_9_;
  assign new_P1_R1162_U124 = P1_REG1_REG_6_ | new_P1_U3469;
  assign new_P1_R1162_U125 = ~new_P1_R1162_U124 | ~new_P1_R1162_U39;
  assign new_P1_R1162_U126 = ~new_P1_R1162_U125 | ~new_P1_R1162_U20 | ~new_P1_R1162_U238 | ~new_P1_R1162_U237;
  assign new_P1_R1162_U127 = ~new_P1_R1162_U111 | ~new_P1_R1162_U20;
  assign new_P1_R1162_U128 = ~P1_REG1_REG_7_ | ~new_P1_U3472;
  assign new_P1_R1162_U129 = ~new_P1_R1162_U127 | ~new_P1_R1162_U128 | ~new_P1_R1162_U6;
  assign new_P1_R1162_U130 = new_P1_U3469 | P1_REG1_REG_6_;
  assign new_P1_R1162_U131 = ~new_P1_R1162_U101 | ~new_P1_R1162_U97;
  assign new_P1_R1162_U132 = ~new_P1_U3457 | ~P1_REG1_REG_2_;
  assign new_P1_R1162_U133 = ~new_P1_R1162_U43;
  assign new_P1_R1162_U134 = ~new_P1_R1162_U100 | ~new_P1_R1162_U5;
  assign new_P1_R1162_U135 = ~new_P1_R1162_U43 | ~new_P1_R1162_U96;
  assign new_P1_R1162_U136 = ~new_P1_U3460 | ~P1_REG1_REG_3_;
  assign new_P1_R1162_U137 = ~new_P1_R1162_U42;
  assign new_P1_R1162_U138 = P1_REG1_REG_4_ | new_P1_U3463;
  assign new_P1_R1162_U139 = ~new_P1_R1162_U138 | ~new_P1_R1162_U42;
  assign new_P1_R1162_U140 = ~new_P1_R1162_U139 | ~new_P1_R1162_U32 | ~new_P1_R1162_U245 | ~new_P1_R1162_U244;
  assign new_P1_R1162_U141 = ~new_P1_R1162_U137 | ~new_P1_R1162_U32;
  assign new_P1_R1162_U142 = ~P1_REG1_REG_5_ | ~new_P1_U3466;
  assign new_P1_R1162_U143 = ~new_P1_R1162_U141 | ~new_P1_R1162_U142 | ~new_P1_R1162_U4;
  assign new_P1_R1162_U144 = new_P1_U3463 | P1_REG1_REG_4_;
  assign new_P1_R1162_U145 = ~new_P1_R1162_U100 | ~new_P1_R1162_U97;
  assign new_P1_R1162_U146 = ~new_P1_R1162_U82;
  assign new_P1_R1162_U147 = ~new_P1_U3460 | ~P1_REG1_REG_3_;
  assign new_P1_R1162_U148 = ~new_P1_R1162_U40 | ~new_P1_R1162_U41 | ~new_P1_R1162_U257 | ~new_P1_R1162_U256;
  assign new_P1_R1162_U149 = ~new_P1_R1162_U41 | ~new_P1_R1162_U40;
  assign new_P1_R1162_U150 = ~new_P1_U3457 | ~P1_REG1_REG_2_;
  assign new_P1_R1162_U151 = ~new_P1_R1162_U149 | ~new_P1_R1162_U150 | ~new_P1_R1162_U97;
  assign new_P1_R1162_U152 = P1_REG1_REG_1_ | new_P1_U3454;
  assign new_P1_R1162_U153 = ~new_P1_R1162_U83;
  assign new_P1_R1162_U154 = new_P1_U3478 | P1_REG1_REG_9_;
  assign new_P1_R1162_U155 = new_P1_U3481 | P1_REG1_REG_10_;
  assign new_P1_R1162_U156 = ~new_P1_R1162_U93 | ~new_P1_R1162_U7;
  assign new_P1_R1162_U157 = ~new_P1_U3481 | ~P1_REG1_REG_10_;
  assign new_P1_R1162_U158 = ~new_P1_R1162_U156 | ~new_P1_R1162_U157 | ~new_P1_R1162_U90;
  assign new_P1_R1162_U159 = P1_REG1_REG_10_ | new_P1_U3481;
  assign new_P1_R1162_U160 = ~new_P1_R1162_U81 | ~new_P1_R1162_U120 | ~new_P1_R1162_U7;
  assign new_P1_R1162_U161 = ~new_P1_R1162_U159 | ~new_P1_R1162_U158;
  assign new_P1_R1162_U162 = ~new_P1_R1162_U88;
  assign new_P1_R1162_U163 = new_P1_U3490 | P1_REG1_REG_13_;
  assign new_P1_R1162_U164 = new_P1_U3487 | P1_REG1_REG_12_;
  assign new_P1_R1162_U165 = ~new_P1_R1162_U92 | ~new_P1_R1162_U8;
  assign new_P1_R1162_U166 = ~new_P1_U3490 | ~P1_REG1_REG_13_;
  assign new_P1_R1162_U167 = ~new_P1_R1162_U165 | ~new_P1_R1162_U166 | ~new_P1_R1162_U91;
  assign new_P1_R1162_U168 = P1_REG1_REG_11_ | new_P1_U3484;
  assign new_P1_R1162_U169 = P1_REG1_REG_13_ | new_P1_U3490;
  assign new_P1_R1162_U170 = ~new_P1_R1162_U88 | ~new_P1_R1162_U168 | ~new_P1_R1162_U8;
  assign new_P1_R1162_U171 = ~new_P1_R1162_U169 | ~new_P1_R1162_U167;
  assign new_P1_R1162_U172 = ~new_P1_R1162_U87;
  assign new_P1_R1162_U173 = P1_REG1_REG_14_ | new_P1_U3493;
  assign new_P1_R1162_U174 = ~new_P1_R1162_U173 | ~new_P1_R1162_U87;
  assign new_P1_R1162_U175 = ~new_P1_U3493 | ~P1_REG1_REG_14_;
  assign new_P1_R1162_U176 = ~new_P1_R1162_U86;
  assign new_P1_R1162_U177 = P1_REG1_REG_15_ | new_P1_U3496;
  assign new_P1_R1162_U178 = ~new_P1_R1162_U177 | ~new_P1_R1162_U86;
  assign new_P1_R1162_U179 = ~new_P1_U3496 | ~P1_REG1_REG_15_;
  assign new_P1_R1162_U180 = ~new_P1_R1162_U66;
  assign new_P1_R1162_U181 = new_P1_U3502 | P1_REG1_REG_17_;
  assign new_P1_R1162_U182 = new_P1_U3499 | P1_REG1_REG_16_;
  assign new_P1_R1162_U183 = ~new_P1_R1162_U47;
  assign new_P1_R1162_U184 = ~new_P1_R1162_U48 | ~new_P1_R1162_U47;
  assign new_P1_R1162_U185 = ~new_P1_U3502 | ~new_P1_R1162_U184;
  assign new_P1_R1162_U186 = ~P1_REG1_REG_17_ | ~new_P1_R1162_U183;
  assign new_P1_R1162_U187 = ~new_P1_R1162_U9 | ~new_P1_R1162_U66;
  assign new_P1_R1162_U188 = ~new_P1_R1162_U65;
  assign new_P1_R1162_U189 = P1_REG1_REG_18_ | new_P1_U3505;
  assign new_P1_R1162_U190 = ~new_P1_R1162_U189 | ~new_P1_R1162_U65;
  assign new_P1_R1162_U191 = ~new_P1_U3505 | ~P1_REG1_REG_18_;
  assign new_P1_R1162_U192 = ~new_P1_R1162_U190 | ~new_P1_R1162_U191 | ~new_P1_R1162_U261 | ~new_P1_R1162_U260;
  assign new_P1_R1162_U193 = ~new_P1_U3505 | ~P1_REG1_REG_18_;
  assign new_P1_R1162_U194 = ~new_P1_R1162_U188 | ~new_P1_R1162_U193;
  assign new_P1_R1162_U195 = new_P1_U3505 | P1_REG1_REG_18_;
  assign new_P1_R1162_U196 = ~new_P1_R1162_U194 | ~new_P1_R1162_U195 | ~new_P1_R1162_U264;
  assign new_P1_R1162_U197 = P1_REG1_REG_16_ | new_P1_U3499;
  assign new_P1_R1162_U198 = ~new_P1_R1162_U197 | ~new_P1_R1162_U66;
  assign new_P1_R1162_U199 = ~new_P1_R1162_U198 | ~new_P1_R1162_U47 | ~new_P1_R1162_U273 | ~new_P1_R1162_U272;
  assign new_P1_R1162_U200 = ~new_P1_R1162_U180 | ~new_P1_R1162_U47;
  assign new_P1_R1162_U201 = ~P1_REG1_REG_17_ | ~new_P1_U3502;
  assign new_P1_R1162_U202 = ~new_P1_R1162_U200 | ~new_P1_R1162_U201 | ~new_P1_R1162_U9;
  assign new_P1_R1162_U203 = new_P1_U3499 | P1_REG1_REG_16_;
  assign new_P1_R1162_U204 = ~new_P1_R1162_U168 | ~new_P1_R1162_U88;
  assign new_P1_R1162_U205 = ~new_P1_R1162_U67;
  assign new_P1_R1162_U206 = P1_REG1_REG_12_ | new_P1_U3487;
  assign new_P1_R1162_U207 = ~new_P1_R1162_U206 | ~new_P1_R1162_U67;
  assign new_P1_R1162_U208 = ~new_P1_R1162_U207 | ~new_P1_R1162_U91 | ~new_P1_R1162_U294 | ~new_P1_R1162_U293;
  assign new_P1_R1162_U209 = ~new_P1_R1162_U205 | ~new_P1_R1162_U91;
  assign new_P1_R1162_U210 = ~new_P1_U3490 | ~P1_REG1_REG_13_;
  assign new_P1_R1162_U211 = ~new_P1_R1162_U209 | ~new_P1_R1162_U210 | ~new_P1_R1162_U8;
  assign new_P1_R1162_U212 = new_P1_U3487 | P1_REG1_REG_12_;
  assign new_P1_R1162_U213 = P1_REG1_REG_9_ | new_P1_U3478;
  assign new_P1_R1162_U214 = ~new_P1_R1162_U213 | ~new_P1_R1162_U38;
  assign new_P1_R1162_U215 = ~new_P1_R1162_U214 | ~new_P1_R1162_U90 | ~new_P1_R1162_U306 | ~new_P1_R1162_U305;
  assign new_P1_R1162_U216 = ~new_P1_R1162_U122 | ~new_P1_R1162_U90;
  assign new_P1_R1162_U217 = ~new_P1_U3481 | ~P1_REG1_REG_10_;
  assign new_P1_R1162_U218 = ~new_P1_R1162_U216 | ~new_P1_R1162_U217 | ~new_P1_R1162_U7;
  assign new_P1_R1162_U219 = ~new_P1_R1162_U123 | ~new_P1_R1162_U90;
  assign new_P1_R1162_U220 = ~new_P1_R1162_U120 | ~new_P1_R1162_U49;
  assign new_P1_R1162_U221 = ~new_P1_R1162_U130 | ~new_P1_R1162_U20;
  assign new_P1_R1162_U222 = ~new_P1_R1162_U144 | ~new_P1_R1162_U32;
  assign new_P1_R1162_U223 = ~new_P1_R1162_U147 | ~new_P1_R1162_U96;
  assign new_P1_R1162_U224 = ~new_P1_R1162_U203 | ~new_P1_R1162_U47;
  assign new_P1_R1162_U225 = ~new_P1_R1162_U212 | ~new_P1_R1162_U91;
  assign new_P1_R1162_U226 = ~new_P1_R1162_U168 | ~new_P1_R1162_U56;
  assign new_P1_R1162_U227 = ~new_P1_U3478 | ~new_P1_R1162_U37;
  assign new_P1_R1162_U228 = ~P1_REG1_REG_9_ | ~new_P1_R1162_U36;
  assign new_P1_R1162_U229 = ~new_P1_R1162_U228 | ~new_P1_R1162_U227;
  assign new_P1_R1162_U230 = ~new_P1_R1162_U219 | ~new_P1_R1162_U38;
  assign new_P1_R1162_U231 = ~new_P1_R1162_U229 | ~new_P1_R1162_U122;
  assign new_P1_R1162_U232 = ~new_P1_U3475 | ~new_P1_R1162_U34;
  assign new_P1_R1162_U233 = ~P1_REG1_REG_8_ | ~new_P1_R1162_U35;
  assign new_P1_R1162_U234 = ~new_P1_R1162_U233 | ~new_P1_R1162_U232;
  assign new_P1_R1162_U235 = ~new_P1_R1162_U220 | ~new_P1_R1162_U81;
  assign new_P1_R1162_U236 = ~new_P1_R1162_U119 | ~new_P1_R1162_U234;
  assign new_P1_R1162_U237 = ~new_P1_U3472 | ~new_P1_R1162_U21;
  assign new_P1_R1162_U238 = ~P1_REG1_REG_7_ | ~new_P1_R1162_U19;
  assign new_P1_R1162_U239 = ~new_P1_U3469 | ~new_P1_R1162_U17;
  assign new_P1_R1162_U240 = ~P1_REG1_REG_6_ | ~new_P1_R1162_U18;
  assign new_P1_R1162_U241 = ~new_P1_R1162_U240 | ~new_P1_R1162_U239;
  assign new_P1_R1162_U242 = ~new_P1_R1162_U221 | ~new_P1_R1162_U39;
  assign new_P1_R1162_U243 = ~new_P1_R1162_U241 | ~new_P1_R1162_U111;
  assign new_P1_R1162_U244 = ~new_P1_U3466 | ~new_P1_R1162_U33;
  assign new_P1_R1162_U245 = ~P1_REG1_REG_5_ | ~new_P1_R1162_U24;
  assign new_P1_R1162_U246 = ~new_P1_U3463 | ~new_P1_R1162_U22;
  assign new_P1_R1162_U247 = ~P1_REG1_REG_4_ | ~new_P1_R1162_U23;
  assign new_P1_R1162_U248 = ~new_P1_R1162_U247 | ~new_P1_R1162_U246;
  assign new_P1_R1162_U249 = ~new_P1_R1162_U222 | ~new_P1_R1162_U42;
  assign new_P1_R1162_U250 = ~new_P1_R1162_U248 | ~new_P1_R1162_U137;
  assign new_P1_R1162_U251 = ~new_P1_U3460 | ~new_P1_R1162_U30;
  assign new_P1_R1162_U252 = ~P1_REG1_REG_3_ | ~new_P1_R1162_U31;
  assign new_P1_R1162_U253 = ~new_P1_R1162_U252 | ~new_P1_R1162_U251;
  assign new_P1_R1162_U254 = ~new_P1_R1162_U223 | ~new_P1_R1162_U82;
  assign new_P1_R1162_U255 = ~new_P1_R1162_U146 | ~new_P1_R1162_U253;
  assign new_P1_R1162_U256 = ~new_P1_U3457 | ~new_P1_R1162_U25;
  assign new_P1_R1162_U257 = ~P1_REG1_REG_2_ | ~new_P1_R1162_U26;
  assign new_P1_R1162_U258 = ~new_P1_R1162_U98 | ~new_P1_R1162_U83;
  assign new_P1_R1162_U259 = ~new_P1_R1162_U153 | ~new_P1_R1162_U29;
  assign new_P1_R1162_U260 = ~new_P1_U3442 | ~new_P1_R1162_U85;
  assign new_P1_R1162_U261 = ~P1_REG1_REG_19_ | ~new_P1_R1162_U84;
  assign new_P1_R1162_U262 = ~new_P1_U3442 | ~new_P1_R1162_U85;
  assign new_P1_R1162_U263 = ~P1_REG1_REG_19_ | ~new_P1_R1162_U84;
  assign new_P1_R1162_U264 = ~new_P1_R1162_U263 | ~new_P1_R1162_U262;
  assign new_P1_R1162_U265 = ~new_P1_U3505 | ~new_P1_R1162_U63;
  assign new_P1_R1162_U266 = ~P1_REG1_REG_18_ | ~new_P1_R1162_U64;
  assign new_P1_R1162_U267 = ~new_P1_U3505 | ~new_P1_R1162_U63;
  assign new_P1_R1162_U268 = ~P1_REG1_REG_18_ | ~new_P1_R1162_U64;
  assign new_P1_R1162_U269 = ~new_P1_R1162_U268 | ~new_P1_R1162_U267;
  assign new_P1_R1162_U270 = ~new_P1_R1162_U65 | ~new_P1_R1162_U266 | ~new_P1_R1162_U265;
  assign new_P1_R1162_U271 = ~new_P1_R1162_U269 | ~new_P1_R1162_U188;
  assign new_P1_R1162_U272 = ~new_P1_U3502 | ~new_P1_R1162_U48;
  assign new_P1_R1162_U273 = ~P1_REG1_REG_17_ | ~new_P1_R1162_U46;
  assign new_P1_R1162_U274 = ~new_P1_U3499 | ~new_P1_R1162_U44;
  assign new_P1_R1162_U275 = ~P1_REG1_REG_16_ | ~new_P1_R1162_U45;
  assign new_P1_R1162_U276 = ~new_P1_R1162_U275 | ~new_P1_R1162_U274;
  assign new_P1_R1162_U277 = ~new_P1_R1162_U224 | ~new_P1_R1162_U66;
  assign new_P1_R1162_U278 = ~new_P1_R1162_U276 | ~new_P1_R1162_U180;
  assign new_P1_R1162_U279 = ~new_P1_U3496 | ~new_P1_R1162_U61;
  assign new_P1_R1162_U280 = ~P1_REG1_REG_15_ | ~new_P1_R1162_U62;
  assign new_P1_R1162_U281 = ~new_P1_U3496 | ~new_P1_R1162_U61;
  assign new_P1_R1162_U282 = ~P1_REG1_REG_15_ | ~new_P1_R1162_U62;
  assign new_P1_R1162_U283 = ~new_P1_R1162_U282 | ~new_P1_R1162_U281;
  assign new_P1_R1162_U284 = ~new_P1_R1162_U86 | ~new_P1_R1162_U280 | ~new_P1_R1162_U279;
  assign new_P1_R1162_U285 = ~new_P1_R1162_U176 | ~new_P1_R1162_U283;
  assign new_P1_R1162_U286 = ~new_P1_U3493 | ~new_P1_R1162_U59;
  assign new_P1_R1162_U287 = ~P1_REG1_REG_14_ | ~new_P1_R1162_U60;
  assign new_P1_R1162_U288 = ~new_P1_U3493 | ~new_P1_R1162_U59;
  assign new_P1_R1162_U289 = ~P1_REG1_REG_14_ | ~new_P1_R1162_U60;
  assign new_P1_R1162_U290 = ~new_P1_R1162_U289 | ~new_P1_R1162_U288;
  assign new_P1_R1162_U291 = ~new_P1_R1162_U87 | ~new_P1_R1162_U287 | ~new_P1_R1162_U286;
  assign new_P1_R1162_U292 = ~new_P1_R1162_U172 | ~new_P1_R1162_U290;
  assign new_P1_R1162_U293 = ~new_P1_U3490 | ~new_P1_R1162_U57;
  assign new_P1_R1162_U294 = ~P1_REG1_REG_13_ | ~new_P1_R1162_U58;
  assign new_P1_R1162_U295 = ~new_P1_U3487 | ~new_P1_R1162_U52;
  assign new_P1_R1162_U296 = ~P1_REG1_REG_12_ | ~new_P1_R1162_U53;
  assign new_P1_R1162_U297 = ~new_P1_R1162_U296 | ~new_P1_R1162_U295;
  assign new_P1_R1162_U298 = ~new_P1_R1162_U225 | ~new_P1_R1162_U67;
  assign new_P1_R1162_U299 = ~new_P1_R1162_U297 | ~new_P1_R1162_U205;
  assign new_P1_R1162_U300 = ~new_P1_U3484 | ~new_P1_R1162_U54;
  assign new_P1_R1162_U301 = ~P1_REG1_REG_11_ | ~new_P1_R1162_U55;
  assign new_P1_R1162_U302 = ~new_P1_R1162_U301 | ~new_P1_R1162_U300;
  assign new_P1_R1162_U303 = ~new_P1_R1162_U226 | ~new_P1_R1162_U88;
  assign new_P1_R1162_U304 = ~new_P1_R1162_U162 | ~new_P1_R1162_U302;
  assign new_P1_R1162_U305 = ~new_P1_U3481 | ~new_P1_R1162_U50;
  assign new_P1_R1162_U306 = ~P1_REG1_REG_10_ | ~new_P1_R1162_U51;
  assign new_P1_R1162_U307 = ~new_P1_U3448 | ~new_P1_R1162_U27;
  assign new_P1_R1162_U308 = ~P1_REG1_REG_0_ | ~new_P1_R1162_U28;
  assign new_P1_R1117_U6 = new_P1_R1117_U198 & new_P1_R1117_U197;
  assign new_P1_R1117_U7 = new_P1_R1117_U237 & new_P1_R1117_U236;
  assign new_P1_R1117_U8 = new_P1_R1117_U254 & new_P1_R1117_U253;
  assign new_P1_R1117_U9 = new_P1_R1117_U280 & new_P1_R1117_U279;
  assign new_P1_R1117_U10 = ~new_P1_R1117_U340 | ~new_P1_R1117_U343;
  assign new_P1_R1117_U11 = ~new_P1_R1117_U329 | ~new_P1_R1117_U332;
  assign new_P1_R1117_U12 = ~new_P1_R1117_U318 | ~new_P1_R1117_U321;
  assign new_P1_R1117_U13 = ~new_P1_R1117_U310 | ~new_P1_R1117_U312;
  assign new_P1_R1117_U14 = ~new_P1_R1117_U347 | ~new_P1_R1117_U308;
  assign new_P1_R1117_U15 = ~new_P1_R1117_U231 | ~new_P1_R1117_U233;
  assign new_P1_R1117_U16 = ~new_P1_R1117_U223 | ~new_P1_R1117_U226;
  assign new_P1_R1117_U17 = ~new_P1_R1117_U215 | ~new_P1_R1117_U217;
  assign new_P1_R1117_U18 = ~new_P1_R1117_U23 | ~new_P1_R1117_U346;
  assign new_P1_R1117_U19 = ~new_P1_U3473;
  assign new_P1_R1117_U20 = ~new_P1_U3467;
  assign new_P1_R1117_U21 = ~new_P1_U3458;
  assign new_P1_R1117_U22 = ~new_P1_U3450;
  assign new_P1_R1117_U23 = ~new_P1_U3450 | ~new_P1_R1117_U91;
  assign new_P1_R1117_U24 = ~new_P1_U3078;
  assign new_P1_R1117_U25 = ~new_P1_U3461;
  assign new_P1_R1117_U26 = ~new_P1_U3068;
  assign new_P1_R1117_U27 = ~new_P1_U3068 | ~new_P1_R1117_U21;
  assign new_P1_R1117_U28 = ~new_P1_U3064;
  assign new_P1_R1117_U29 = ~new_P1_U3470;
  assign new_P1_R1117_U30 = ~new_P1_U3464;
  assign new_P1_R1117_U31 = ~new_P1_U3071;
  assign new_P1_R1117_U32 = ~new_P1_U3067;
  assign new_P1_R1117_U33 = ~new_P1_U3060;
  assign new_P1_R1117_U34 = ~new_P1_U3060 | ~new_P1_R1117_U30;
  assign new_P1_R1117_U35 = ~new_P1_U3476;
  assign new_P1_R1117_U36 = ~new_P1_U3070;
  assign new_P1_R1117_U37 = ~new_P1_U3070 | ~new_P1_R1117_U19;
  assign new_P1_R1117_U38 = ~new_P1_U3084;
  assign new_P1_R1117_U39 = ~new_P1_U3479;
  assign new_P1_R1117_U40 = ~new_P1_U3083;
  assign new_P1_R1117_U41 = ~new_P1_R1117_U204 | ~new_P1_R1117_U203;
  assign new_P1_R1117_U42 = ~new_P1_R1117_U34 | ~new_P1_R1117_U219;
  assign new_P1_R1117_U43 = ~new_P1_R1117_U188 | ~new_P1_R1117_U187;
  assign new_P1_R1117_U44 = ~new_P1_U3976;
  assign new_P1_R1117_U45 = ~new_P1_U3980;
  assign new_P1_R1117_U46 = ~new_P1_U3497;
  assign new_P1_R1117_U47 = ~new_P1_U3482;
  assign new_P1_R1117_U48 = ~new_P1_U3485;
  assign new_P1_R1117_U49 = ~new_P1_U3063;
  assign new_P1_R1117_U50 = ~new_P1_U3062;
  assign new_P1_R1117_U51 = ~new_P1_U3083 | ~new_P1_R1117_U39;
  assign new_P1_R1117_U52 = ~new_P1_U3488;
  assign new_P1_R1117_U53 = ~new_P1_U3072;
  assign new_P1_R1117_U54 = ~new_P1_U3491;
  assign new_P1_R1117_U55 = ~new_P1_U3080;
  assign new_P1_R1117_U56 = ~new_P1_U3500;
  assign new_P1_R1117_U57 = ~new_P1_U3494;
  assign new_P1_R1117_U58 = ~new_P1_U3073;
  assign new_P1_R1117_U59 = ~new_P1_U3074;
  assign new_P1_R1117_U60 = ~new_P1_U3079;
  assign new_P1_R1117_U61 = ~new_P1_U3079 | ~new_P1_R1117_U57;
  assign new_P1_R1117_U62 = ~new_P1_U3503;
  assign new_P1_R1117_U63 = ~new_P1_U3069;
  assign new_P1_R1117_U64 = ~new_P1_R1117_U264 | ~new_P1_R1117_U263;
  assign new_P1_R1117_U65 = ~new_P1_U3082;
  assign new_P1_R1117_U66 = ~new_P1_U3508;
  assign new_P1_R1117_U67 = ~new_P1_U3081;
  assign new_P1_R1117_U68 = ~new_P1_U3982;
  assign new_P1_R1117_U69 = ~new_P1_U3076;
  assign new_P1_R1117_U70 = ~new_P1_U3979;
  assign new_P1_R1117_U71 = ~new_P1_U3981;
  assign new_P1_R1117_U72 = ~new_P1_U3066;
  assign new_P1_R1117_U73 = ~new_P1_U3061;
  assign new_P1_R1117_U74 = ~new_P1_U3075;
  assign new_P1_R1117_U75 = ~new_P1_U3075 | ~new_P1_R1117_U71;
  assign new_P1_R1117_U76 = ~new_P1_U3978;
  assign new_P1_R1117_U77 = ~new_P1_U3065;
  assign new_P1_R1117_U78 = ~new_P1_U3977;
  assign new_P1_R1117_U79 = ~new_P1_U3058;
  assign new_P1_R1117_U80 = ~new_P1_U3975;
  assign new_P1_R1117_U81 = ~new_P1_U3057;
  assign new_P1_R1117_U82 = ~new_P1_U3057 | ~new_P1_R1117_U44;
  assign new_P1_R1117_U83 = ~new_P1_U3053;
  assign new_P1_R1117_U84 = ~new_P1_U3974;
  assign new_P1_R1117_U85 = ~new_P1_U3054;
  assign new_P1_R1117_U86 = ~new_P1_R1117_U126 | ~new_P1_R1117_U297;
  assign new_P1_R1117_U87 = ~new_P1_R1117_U294 | ~new_P1_R1117_U293;
  assign new_P1_R1117_U88 = ~new_P1_R1117_U75 | ~new_P1_R1117_U314;
  assign new_P1_R1117_U89 = ~new_P1_R1117_U61 | ~new_P1_R1117_U325;
  assign new_P1_R1117_U90 = ~new_P1_R1117_U51 | ~new_P1_R1117_U336;
  assign new_P1_R1117_U91 = ~new_P1_U3077;
  assign new_P1_R1117_U92 = ~new_P1_R1117_U390 | ~new_P1_R1117_U389;
  assign new_P1_R1117_U93 = ~new_P1_R1117_U404 | ~new_P1_R1117_U403;
  assign new_P1_R1117_U94 = ~new_P1_R1117_U409 | ~new_P1_R1117_U408;
  assign new_P1_R1117_U95 = ~new_P1_R1117_U425 | ~new_P1_R1117_U424;
  assign new_P1_R1117_U96 = ~new_P1_R1117_U430 | ~new_P1_R1117_U429;
  assign new_P1_R1117_U97 = ~new_P1_R1117_U435 | ~new_P1_R1117_U434;
  assign new_P1_R1117_U98 = ~new_P1_R1117_U440 | ~new_P1_R1117_U439;
  assign new_P1_R1117_U99 = ~new_P1_R1117_U445 | ~new_P1_R1117_U444;
  assign new_P1_R1117_U100 = ~new_P1_R1117_U461 | ~new_P1_R1117_U460;
  assign new_P1_R1117_U101 = ~new_P1_R1117_U466 | ~new_P1_R1117_U465;
  assign new_P1_R1117_U102 = ~new_P1_R1117_U351 | ~new_P1_R1117_U350;
  assign new_P1_R1117_U103 = ~new_P1_R1117_U360 | ~new_P1_R1117_U359;
  assign new_P1_R1117_U104 = ~new_P1_R1117_U367 | ~new_P1_R1117_U366;
  assign new_P1_R1117_U105 = ~new_P1_R1117_U371 | ~new_P1_R1117_U370;
  assign new_P1_R1117_U106 = ~new_P1_R1117_U380 | ~new_P1_R1117_U379;
  assign new_P1_R1117_U107 = ~new_P1_R1117_U399 | ~new_P1_R1117_U398;
  assign new_P1_R1117_U108 = ~new_P1_R1117_U416 | ~new_P1_R1117_U415;
  assign new_P1_R1117_U109 = ~new_P1_R1117_U420 | ~new_P1_R1117_U419;
  assign new_P1_R1117_U110 = ~new_P1_R1117_U452 | ~new_P1_R1117_U451;
  assign new_P1_R1117_U111 = ~new_P1_R1117_U456 | ~new_P1_R1117_U455;
  assign new_P1_R1117_U112 = ~new_P1_R1117_U473 | ~new_P1_R1117_U472;
  assign new_P1_R1117_U113 = new_P1_R1117_U193 & new_P1_R1117_U194;
  assign new_P1_R1117_U114 = new_P1_R1117_U201 & new_P1_R1117_U196;
  assign new_P1_R1117_U115 = new_P1_R1117_U206 & new_P1_R1117_U180;
  assign new_P1_R1117_U116 = new_P1_R1117_U209 & new_P1_R1117_U210;
  assign new_P1_R1117_U117 = new_P1_R1117_U37 & new_P1_R1117_U353 & new_P1_R1117_U352;
  assign new_P1_R1117_U118 = new_P1_R1117_U356 & new_P1_R1117_U180;
  assign new_P1_R1117_U119 = new_P1_R1117_U225 & new_P1_R1117_U6;
  assign new_P1_R1117_U120 = new_P1_R1117_U363 & new_P1_R1117_U179;
  assign new_P1_R1117_U121 = new_P1_R1117_U27 & new_P1_R1117_U373 & new_P1_R1117_U372;
  assign new_P1_R1117_U122 = new_P1_R1117_U376 & new_P1_R1117_U178;
  assign new_P1_R1117_U123 = new_P1_R1117_U174 & new_P1_R1117_U235 & new_P1_R1117_U212;
  assign new_P1_R1117_U124 = new_P1_R1117_U252 & new_P1_R1117_U257 & new_P1_R1117_U175;
  assign new_P1_R1117_U125 = new_P1_R1117_U283 & new_P1_R1117_U176;
  assign new_P1_R1117_U126 = new_P1_R1117_U299 & new_P1_R1117_U300;
  assign new_P1_R1117_U127 = ~new_P1_R1117_U387 | ~new_P1_R1117_U386;
  assign new_P1_R1117_U128 = new_P1_R1117_U82 & new_P1_R1117_U392 & new_P1_R1117_U391;
  assign new_P1_R1117_U129 = new_P1_R1117_U395 & new_P1_R1117_U177;
  assign new_P1_R1117_U130 = ~new_P1_R1117_U401 | ~new_P1_R1117_U400;
  assign new_P1_R1117_U131 = ~new_P1_R1117_U406 | ~new_P1_R1117_U405;
  assign new_P1_R1117_U132 = new_P1_R1117_U412 & new_P1_R1117_U176;
  assign new_P1_R1117_U133 = ~new_P1_R1117_U422 | ~new_P1_R1117_U421;
  assign new_P1_R1117_U134 = ~new_P1_R1117_U427 | ~new_P1_R1117_U426;
  assign new_P1_R1117_U135 = ~new_P1_R1117_U432 | ~new_P1_R1117_U431;
  assign new_P1_R1117_U136 = ~new_P1_R1117_U437 | ~new_P1_R1117_U436;
  assign new_P1_R1117_U137 = ~new_P1_R1117_U442 | ~new_P1_R1117_U441;
  assign new_P1_R1117_U138 = new_P1_R1117_U331 & new_P1_R1117_U8;
  assign new_P1_R1117_U139 = new_P1_R1117_U448 & new_P1_R1117_U175;
  assign new_P1_R1117_U140 = ~new_P1_R1117_U458 | ~new_P1_R1117_U457;
  assign new_P1_R1117_U141 = ~new_P1_R1117_U463 | ~new_P1_R1117_U462;
  assign new_P1_R1117_U142 = new_P1_R1117_U342 & new_P1_R1117_U7;
  assign new_P1_R1117_U143 = new_P1_R1117_U469 & new_P1_R1117_U174;
  assign new_P1_R1117_U144 = new_P1_R1117_U349 & new_P1_R1117_U348;
  assign new_P1_R1117_U145 = ~new_P1_R1117_U116 | ~new_P1_R1117_U207;
  assign new_P1_R1117_U146 = new_P1_R1117_U358 & new_P1_R1117_U357;
  assign new_P1_R1117_U147 = new_P1_R1117_U365 & new_P1_R1117_U364;
  assign new_P1_R1117_U148 = new_P1_R1117_U369 & new_P1_R1117_U368;
  assign new_P1_R1117_U149 = ~new_P1_R1117_U113 | ~new_P1_R1117_U191;
  assign new_P1_R1117_U150 = new_P1_R1117_U378 & new_P1_R1117_U377;
  assign new_P1_R1117_U151 = ~new_P1_U3985;
  assign new_P1_R1117_U152 = ~new_P1_U3055;
  assign new_P1_R1117_U153 = new_P1_R1117_U382 & new_P1_R1117_U381;
  assign new_P1_R1117_U154 = new_P1_R1117_U397 & new_P1_R1117_U396;
  assign new_P1_R1117_U155 = ~new_P1_R1117_U290 | ~new_P1_R1117_U289;
  assign new_P1_R1117_U156 = ~new_P1_R1117_U286 | ~new_P1_R1117_U285;
  assign new_P1_R1117_U157 = new_P1_R1117_U414 & new_P1_R1117_U413;
  assign new_P1_R1117_U158 = new_P1_R1117_U418 & new_P1_R1117_U417;
  assign new_P1_R1117_U159 = ~new_P1_R1117_U276 | ~new_P1_R1117_U275;
  assign new_P1_R1117_U160 = ~new_P1_R1117_U272 | ~new_P1_R1117_U271;
  assign new_P1_R1117_U161 = ~new_P1_U3455;
  assign new_P1_R1117_U162 = ~new_P1_R1117_U268 | ~new_P1_R1117_U267;
  assign new_P1_R1117_U163 = ~new_P1_U3506;
  assign new_P1_R1117_U164 = ~new_P1_R1117_U260 | ~new_P1_R1117_U259;
  assign new_P1_R1117_U165 = new_P1_R1117_U450 & new_P1_R1117_U449;
  assign new_P1_R1117_U166 = new_P1_R1117_U454 & new_P1_R1117_U453;
  assign new_P1_R1117_U167 = ~new_P1_R1117_U250 | ~new_P1_R1117_U249;
  assign new_P1_R1117_U168 = ~new_P1_R1117_U246 | ~new_P1_R1117_U245;
  assign new_P1_R1117_U169 = ~new_P1_R1117_U242 | ~new_P1_R1117_U241;
  assign new_P1_R1117_U170 = new_P1_R1117_U471 & new_P1_R1117_U470;
  assign new_P1_R1117_U171 = ~new_P1_R1117_U82;
  assign new_P1_R1117_U172 = ~new_P1_R1117_U27;
  assign new_P1_R1117_U173 = ~new_P1_R1117_U37;
  assign new_P1_R1117_U174 = ~new_P1_U3482 | ~new_P1_R1117_U50;
  assign new_P1_R1117_U175 = ~new_P1_U3497 | ~new_P1_R1117_U59;
  assign new_P1_R1117_U176 = ~new_P1_U3980 | ~new_P1_R1117_U73;
  assign new_P1_R1117_U177 = ~new_P1_U3976 | ~new_P1_R1117_U81;
  assign new_P1_R1117_U178 = ~new_P1_U3458 | ~new_P1_R1117_U26;
  assign new_P1_R1117_U179 = ~new_P1_U3467 | ~new_P1_R1117_U32;
  assign new_P1_R1117_U180 = ~new_P1_U3473 | ~new_P1_R1117_U36;
  assign new_P1_R1117_U181 = ~new_P1_R1117_U61;
  assign new_P1_R1117_U182 = ~new_P1_R1117_U75;
  assign new_P1_R1117_U183 = ~new_P1_R1117_U34;
  assign new_P1_R1117_U184 = ~new_P1_R1117_U51;
  assign new_P1_R1117_U185 = ~new_P1_R1117_U23;
  assign new_P1_R1117_U186 = ~new_P1_R1117_U185 | ~new_P1_R1117_U24;
  assign new_P1_R1117_U187 = ~new_P1_R1117_U186 | ~new_P1_R1117_U161;
  assign new_P1_R1117_U188 = ~new_P1_U3078 | ~new_P1_R1117_U23;
  assign new_P1_R1117_U189 = ~new_P1_R1117_U43;
  assign new_P1_R1117_U190 = ~new_P1_U3461 | ~new_P1_R1117_U28;
  assign new_P1_R1117_U191 = ~new_P1_R1117_U190 | ~new_P1_R1117_U43 | ~new_P1_R1117_U178;
  assign new_P1_R1117_U192 = ~new_P1_R1117_U28 | ~new_P1_R1117_U27;
  assign new_P1_R1117_U193 = ~new_P1_R1117_U192 | ~new_P1_R1117_U25;
  assign new_P1_R1117_U194 = ~new_P1_U3064 | ~new_P1_R1117_U172;
  assign new_P1_R1117_U195 = ~new_P1_R1117_U149;
  assign new_P1_R1117_U196 = ~new_P1_U3470 | ~new_P1_R1117_U31;
  assign new_P1_R1117_U197 = ~new_P1_U3071 | ~new_P1_R1117_U29;
  assign new_P1_R1117_U198 = ~new_P1_U3067 | ~new_P1_R1117_U20;
  assign new_P1_R1117_U199 = ~new_P1_R1117_U183 | ~new_P1_R1117_U179;
  assign new_P1_R1117_U200 = ~new_P1_R1117_U6 | ~new_P1_R1117_U199;
  assign new_P1_R1117_U201 = ~new_P1_U3464 | ~new_P1_R1117_U33;
  assign new_P1_R1117_U202 = ~new_P1_U3470 | ~new_P1_R1117_U31;
  assign new_P1_R1117_U203 = ~new_P1_R1117_U114 | ~new_P1_R1117_U149 | ~new_P1_R1117_U179;
  assign new_P1_R1117_U204 = ~new_P1_R1117_U202 | ~new_P1_R1117_U200;
  assign new_P1_R1117_U205 = ~new_P1_R1117_U41;
  assign new_P1_R1117_U206 = ~new_P1_U3476 | ~new_P1_R1117_U38;
  assign new_P1_R1117_U207 = ~new_P1_R1117_U115 | ~new_P1_R1117_U41;
  assign new_P1_R1117_U208 = ~new_P1_R1117_U38 | ~new_P1_R1117_U37;
  assign new_P1_R1117_U209 = ~new_P1_R1117_U208 | ~new_P1_R1117_U35;
  assign new_P1_R1117_U210 = ~new_P1_U3084 | ~new_P1_R1117_U173;
  assign new_P1_R1117_U211 = ~new_P1_R1117_U145;
  assign new_P1_R1117_U212 = ~new_P1_U3479 | ~new_P1_R1117_U40;
  assign new_P1_R1117_U213 = ~new_P1_R1117_U212 | ~new_P1_R1117_U51;
  assign new_P1_R1117_U214 = ~new_P1_R1117_U205 | ~new_P1_R1117_U37;
  assign new_P1_R1117_U215 = ~new_P1_R1117_U118 | ~new_P1_R1117_U214;
  assign new_P1_R1117_U216 = ~new_P1_R1117_U41 | ~new_P1_R1117_U180;
  assign new_P1_R1117_U217 = ~new_P1_R1117_U117 | ~new_P1_R1117_U216;
  assign new_P1_R1117_U218 = ~new_P1_R1117_U37 | ~new_P1_R1117_U180;
  assign new_P1_R1117_U219 = ~new_P1_R1117_U201 | ~new_P1_R1117_U149;
  assign new_P1_R1117_U220 = ~new_P1_R1117_U42;
  assign new_P1_R1117_U221 = ~new_P1_U3067 | ~new_P1_R1117_U20;
  assign new_P1_R1117_U222 = ~new_P1_R1117_U220 | ~new_P1_R1117_U221;
  assign new_P1_R1117_U223 = ~new_P1_R1117_U120 | ~new_P1_R1117_U222;
  assign new_P1_R1117_U224 = ~new_P1_R1117_U42 | ~new_P1_R1117_U179;
  assign new_P1_R1117_U225 = ~new_P1_U3470 | ~new_P1_R1117_U31;
  assign new_P1_R1117_U226 = ~new_P1_R1117_U119 | ~new_P1_R1117_U224;
  assign new_P1_R1117_U227 = ~new_P1_U3067 | ~new_P1_R1117_U20;
  assign new_P1_R1117_U228 = ~new_P1_R1117_U179 | ~new_P1_R1117_U227;
  assign new_P1_R1117_U229 = ~new_P1_R1117_U201 | ~new_P1_R1117_U34;
  assign new_P1_R1117_U230 = ~new_P1_R1117_U189 | ~new_P1_R1117_U27;
  assign new_P1_R1117_U231 = ~new_P1_R1117_U122 | ~new_P1_R1117_U230;
  assign new_P1_R1117_U232 = ~new_P1_R1117_U43 | ~new_P1_R1117_U178;
  assign new_P1_R1117_U233 = ~new_P1_R1117_U121 | ~new_P1_R1117_U232;
  assign new_P1_R1117_U234 = ~new_P1_R1117_U27 | ~new_P1_R1117_U178;
  assign new_P1_R1117_U235 = ~new_P1_U3485 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U236 = ~new_P1_U3063 | ~new_P1_R1117_U48;
  assign new_P1_R1117_U237 = ~new_P1_U3062 | ~new_P1_R1117_U47;
  assign new_P1_R1117_U238 = ~new_P1_R1117_U184 | ~new_P1_R1117_U174;
  assign new_P1_R1117_U239 = ~new_P1_R1117_U7 | ~new_P1_R1117_U238;
  assign new_P1_R1117_U240 = ~new_P1_U3485 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U241 = ~new_P1_R1117_U145 | ~new_P1_R1117_U123;
  assign new_P1_R1117_U242 = ~new_P1_R1117_U240 | ~new_P1_R1117_U239;
  assign new_P1_R1117_U243 = ~new_P1_R1117_U169;
  assign new_P1_R1117_U244 = ~new_P1_U3488 | ~new_P1_R1117_U53;
  assign new_P1_R1117_U245 = ~new_P1_R1117_U244 | ~new_P1_R1117_U169;
  assign new_P1_R1117_U246 = ~new_P1_U3072 | ~new_P1_R1117_U52;
  assign new_P1_R1117_U247 = ~new_P1_R1117_U168;
  assign new_P1_R1117_U248 = ~new_P1_U3491 | ~new_P1_R1117_U55;
  assign new_P1_R1117_U249 = ~new_P1_R1117_U248 | ~new_P1_R1117_U168;
  assign new_P1_R1117_U250 = ~new_P1_U3080 | ~new_P1_R1117_U54;
  assign new_P1_R1117_U251 = ~new_P1_R1117_U167;
  assign new_P1_R1117_U252 = ~new_P1_U3500 | ~new_P1_R1117_U58;
  assign new_P1_R1117_U253 = ~new_P1_U3073 | ~new_P1_R1117_U56;
  assign new_P1_R1117_U254 = ~new_P1_U3074 | ~new_P1_R1117_U46;
  assign new_P1_R1117_U255 = ~new_P1_R1117_U181 | ~new_P1_R1117_U175;
  assign new_P1_R1117_U256 = ~new_P1_R1117_U8 | ~new_P1_R1117_U255;
  assign new_P1_R1117_U257 = ~new_P1_U3494 | ~new_P1_R1117_U60;
  assign new_P1_R1117_U258 = ~new_P1_U3500 | ~new_P1_R1117_U58;
  assign new_P1_R1117_U259 = ~new_P1_R1117_U167 | ~new_P1_R1117_U124;
  assign new_P1_R1117_U260 = ~new_P1_R1117_U258 | ~new_P1_R1117_U256;
  assign new_P1_R1117_U261 = ~new_P1_R1117_U164;
  assign new_P1_R1117_U262 = ~new_P1_U3503 | ~new_P1_R1117_U63;
  assign new_P1_R1117_U263 = ~new_P1_R1117_U262 | ~new_P1_R1117_U164;
  assign new_P1_R1117_U264 = ~new_P1_U3069 | ~new_P1_R1117_U62;
  assign new_P1_R1117_U265 = ~new_P1_R1117_U64;
  assign new_P1_R1117_U266 = ~new_P1_R1117_U265 | ~new_P1_R1117_U65;
  assign new_P1_R1117_U267 = ~new_P1_R1117_U266 | ~new_P1_R1117_U163;
  assign new_P1_R1117_U268 = ~new_P1_U3082 | ~new_P1_R1117_U64;
  assign new_P1_R1117_U269 = ~new_P1_R1117_U162;
  assign new_P1_R1117_U270 = ~new_P1_U3508 | ~new_P1_R1117_U67;
  assign new_P1_R1117_U271 = ~new_P1_R1117_U270 | ~new_P1_R1117_U162;
  assign new_P1_R1117_U272 = ~new_P1_U3081 | ~new_P1_R1117_U66;
  assign new_P1_R1117_U273 = ~new_P1_R1117_U160;
  assign new_P1_R1117_U274 = ~new_P1_U3982 | ~new_P1_R1117_U69;
  assign new_P1_R1117_U275 = ~new_P1_R1117_U274 | ~new_P1_R1117_U160;
  assign new_P1_R1117_U276 = ~new_P1_U3076 | ~new_P1_R1117_U68;
  assign new_P1_R1117_U277 = ~new_P1_R1117_U159;
  assign new_P1_R1117_U278 = ~new_P1_U3979 | ~new_P1_R1117_U72;
  assign new_P1_R1117_U279 = ~new_P1_U3066 | ~new_P1_R1117_U70;
  assign new_P1_R1117_U280 = ~new_P1_U3061 | ~new_P1_R1117_U45;
  assign new_P1_R1117_U281 = ~new_P1_R1117_U182 | ~new_P1_R1117_U176;
  assign new_P1_R1117_U282 = ~new_P1_R1117_U9 | ~new_P1_R1117_U281;
  assign new_P1_R1117_U283 = ~new_P1_U3981 | ~new_P1_R1117_U74;
  assign new_P1_R1117_U284 = ~new_P1_U3979 | ~new_P1_R1117_U72;
  assign new_P1_R1117_U285 = ~new_P1_R1117_U278 | ~new_P1_R1117_U159 | ~new_P1_R1117_U125;
  assign new_P1_R1117_U286 = ~new_P1_R1117_U284 | ~new_P1_R1117_U282;
  assign new_P1_R1117_U287 = ~new_P1_R1117_U156;
  assign new_P1_R1117_U288 = ~new_P1_U3978 | ~new_P1_R1117_U77;
  assign new_P1_R1117_U289 = ~new_P1_R1117_U288 | ~new_P1_R1117_U156;
  assign new_P1_R1117_U290 = ~new_P1_U3065 | ~new_P1_R1117_U76;
  assign new_P1_R1117_U291 = ~new_P1_R1117_U155;
  assign new_P1_R1117_U292 = ~new_P1_U3977 | ~new_P1_R1117_U79;
  assign new_P1_R1117_U293 = ~new_P1_R1117_U292 | ~new_P1_R1117_U155;
  assign new_P1_R1117_U294 = ~new_P1_U3058 | ~new_P1_R1117_U78;
  assign new_P1_R1117_U295 = ~new_P1_R1117_U87;
  assign new_P1_R1117_U296 = ~new_P1_U3975 | ~new_P1_R1117_U83;
  assign new_P1_R1117_U297 = ~new_P1_R1117_U296 | ~new_P1_R1117_U87 | ~new_P1_R1117_U177;
  assign new_P1_R1117_U298 = ~new_P1_R1117_U83 | ~new_P1_R1117_U82;
  assign new_P1_R1117_U299 = ~new_P1_R1117_U298 | ~new_P1_R1117_U80;
  assign new_P1_R1117_U300 = ~new_P1_U3053 | ~new_P1_R1117_U171;
  assign new_P1_R1117_U301 = ~new_P1_R1117_U86;
  assign new_P1_R1117_U302 = ~new_P1_U3054 | ~new_P1_R1117_U84;
  assign new_P1_R1117_U303 = ~new_P1_R1117_U301 | ~new_P1_R1117_U302;
  assign new_P1_R1117_U304 = ~new_P1_U3974 | ~new_P1_R1117_U85;
  assign new_P1_R1117_U305 = ~new_P1_U3974 | ~new_P1_R1117_U85;
  assign new_P1_R1117_U306 = ~new_P1_R1117_U305 | ~new_P1_R1117_U86;
  assign new_P1_R1117_U307 = ~new_P1_U3054 | ~new_P1_R1117_U84;
  assign new_P1_R1117_U308 = ~new_P1_R1117_U153 | ~new_P1_R1117_U307 | ~new_P1_R1117_U306;
  assign new_P1_R1117_U309 = ~new_P1_R1117_U295 | ~new_P1_R1117_U82;
  assign new_P1_R1117_U310 = ~new_P1_R1117_U129 | ~new_P1_R1117_U309;
  assign new_P1_R1117_U311 = ~new_P1_R1117_U87 | ~new_P1_R1117_U177;
  assign new_P1_R1117_U312 = ~new_P1_R1117_U128 | ~new_P1_R1117_U311;
  assign new_P1_R1117_U313 = ~new_P1_R1117_U82 | ~new_P1_R1117_U177;
  assign new_P1_R1117_U314 = ~new_P1_R1117_U283 | ~new_P1_R1117_U159;
  assign new_P1_R1117_U315 = ~new_P1_R1117_U88;
  assign new_P1_R1117_U316 = ~new_P1_U3061 | ~new_P1_R1117_U45;
  assign new_P1_R1117_U317 = ~new_P1_R1117_U315 | ~new_P1_R1117_U316;
  assign new_P1_R1117_U318 = ~new_P1_R1117_U132 | ~new_P1_R1117_U317;
  assign new_P1_R1117_U319 = ~new_P1_R1117_U88 | ~new_P1_R1117_U176;
  assign new_P1_R1117_U320 = ~new_P1_U3979 | ~new_P1_R1117_U72;
  assign new_P1_R1117_U321 = ~new_P1_R1117_U9 | ~new_P1_R1117_U320 | ~new_P1_R1117_U319;
  assign new_P1_R1117_U322 = ~new_P1_U3061 | ~new_P1_R1117_U45;
  assign new_P1_R1117_U323 = ~new_P1_R1117_U176 | ~new_P1_R1117_U322;
  assign new_P1_R1117_U324 = ~new_P1_R1117_U283 | ~new_P1_R1117_U75;
  assign new_P1_R1117_U325 = ~new_P1_R1117_U257 | ~new_P1_R1117_U167;
  assign new_P1_R1117_U326 = ~new_P1_R1117_U89;
  assign new_P1_R1117_U327 = ~new_P1_U3074 | ~new_P1_R1117_U46;
  assign new_P1_R1117_U328 = ~new_P1_R1117_U326 | ~new_P1_R1117_U327;
  assign new_P1_R1117_U329 = ~new_P1_R1117_U139 | ~new_P1_R1117_U328;
  assign new_P1_R1117_U330 = ~new_P1_R1117_U89 | ~new_P1_R1117_U175;
  assign new_P1_R1117_U331 = ~new_P1_U3500 | ~new_P1_R1117_U58;
  assign new_P1_R1117_U332 = ~new_P1_R1117_U138 | ~new_P1_R1117_U330;
  assign new_P1_R1117_U333 = ~new_P1_U3074 | ~new_P1_R1117_U46;
  assign new_P1_R1117_U334 = ~new_P1_R1117_U175 | ~new_P1_R1117_U333;
  assign new_P1_R1117_U335 = ~new_P1_R1117_U257 | ~new_P1_R1117_U61;
  assign new_P1_R1117_U336 = ~new_P1_R1117_U212 | ~new_P1_R1117_U145;
  assign new_P1_R1117_U337 = ~new_P1_R1117_U90;
  assign new_P1_R1117_U338 = ~new_P1_U3062 | ~new_P1_R1117_U47;
  assign new_P1_R1117_U339 = ~new_P1_R1117_U337 | ~new_P1_R1117_U338;
  assign new_P1_R1117_U340 = ~new_P1_R1117_U143 | ~new_P1_R1117_U339;
  assign new_P1_R1117_U341 = ~new_P1_R1117_U90 | ~new_P1_R1117_U174;
  assign new_P1_R1117_U342 = ~new_P1_U3485 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U343 = ~new_P1_R1117_U142 | ~new_P1_R1117_U341;
  assign new_P1_R1117_U344 = ~new_P1_U3062 | ~new_P1_R1117_U47;
  assign new_P1_R1117_U345 = ~new_P1_R1117_U174 | ~new_P1_R1117_U344;
  assign new_P1_R1117_U346 = ~new_P1_U3077 | ~new_P1_R1117_U22;
  assign new_P1_R1117_U347 = ~new_P1_R1117_U385 | ~new_P1_R1117_U304 | ~new_P1_R1117_U303;
  assign new_P1_R1117_U348 = ~new_P1_U3479 | ~new_P1_R1117_U40;
  assign new_P1_R1117_U349 = ~new_P1_U3083 | ~new_P1_R1117_U39;
  assign new_P1_R1117_U350 = ~new_P1_R1117_U213 | ~new_P1_R1117_U145;
  assign new_P1_R1117_U351 = ~new_P1_R1117_U211 | ~new_P1_R1117_U144;
  assign new_P1_R1117_U352 = ~new_P1_U3476 | ~new_P1_R1117_U38;
  assign new_P1_R1117_U353 = ~new_P1_U3084 | ~new_P1_R1117_U35;
  assign new_P1_R1117_U354 = ~new_P1_U3476 | ~new_P1_R1117_U38;
  assign new_P1_R1117_U355 = ~new_P1_U3084 | ~new_P1_R1117_U35;
  assign new_P1_R1117_U356 = ~new_P1_R1117_U355 | ~new_P1_R1117_U354;
  assign new_P1_R1117_U357 = ~new_P1_U3473 | ~new_P1_R1117_U36;
  assign new_P1_R1117_U358 = ~new_P1_U3070 | ~new_P1_R1117_U19;
  assign new_P1_R1117_U359 = ~new_P1_R1117_U218 | ~new_P1_R1117_U41;
  assign new_P1_R1117_U360 = ~new_P1_R1117_U146 | ~new_P1_R1117_U205;
  assign new_P1_R1117_U361 = ~new_P1_U3470 | ~new_P1_R1117_U31;
  assign new_P1_R1117_U362 = ~new_P1_U3071 | ~new_P1_R1117_U29;
  assign new_P1_R1117_U363 = ~new_P1_R1117_U362 | ~new_P1_R1117_U361;
  assign new_P1_R1117_U364 = ~new_P1_U3467 | ~new_P1_R1117_U32;
  assign new_P1_R1117_U365 = ~new_P1_U3067 | ~new_P1_R1117_U20;
  assign new_P1_R1117_U366 = ~new_P1_R1117_U228 | ~new_P1_R1117_U42;
  assign new_P1_R1117_U367 = ~new_P1_R1117_U147 | ~new_P1_R1117_U220;
  assign new_P1_R1117_U368 = ~new_P1_U3464 | ~new_P1_R1117_U33;
  assign new_P1_R1117_U369 = ~new_P1_U3060 | ~new_P1_R1117_U30;
  assign new_P1_R1117_U370 = ~new_P1_R1117_U229 | ~new_P1_R1117_U149;
  assign new_P1_R1117_U371 = ~new_P1_R1117_U195 | ~new_P1_R1117_U148;
  assign new_P1_R1117_U372 = ~new_P1_U3461 | ~new_P1_R1117_U28;
  assign new_P1_R1117_U373 = ~new_P1_U3064 | ~new_P1_R1117_U25;
  assign new_P1_R1117_U374 = ~new_P1_U3461 | ~new_P1_R1117_U28;
  assign new_P1_R1117_U375 = ~new_P1_U3064 | ~new_P1_R1117_U25;
  assign new_P1_R1117_U376 = ~new_P1_R1117_U375 | ~new_P1_R1117_U374;
  assign new_P1_R1117_U377 = ~new_P1_U3458 | ~new_P1_R1117_U26;
  assign new_P1_R1117_U378 = ~new_P1_U3068 | ~new_P1_R1117_U21;
  assign new_P1_R1117_U379 = ~new_P1_R1117_U234 | ~new_P1_R1117_U43;
  assign new_P1_R1117_U380 = ~new_P1_R1117_U150 | ~new_P1_R1117_U189;
  assign new_P1_R1117_U381 = ~new_P1_U3985 | ~new_P1_R1117_U152;
  assign new_P1_R1117_U382 = ~new_P1_U3055 | ~new_P1_R1117_U151;
  assign new_P1_R1117_U383 = ~new_P1_U3985 | ~new_P1_R1117_U152;
  assign new_P1_R1117_U384 = ~new_P1_U3055 | ~new_P1_R1117_U151;
  assign new_P1_R1117_U385 = ~new_P1_R1117_U384 | ~new_P1_R1117_U383;
  assign new_P1_R1117_U386 = ~new_P1_U3974 | ~new_P1_R1117_U85;
  assign new_P1_R1117_U387 = ~new_P1_U3054 | ~new_P1_R1117_U84;
  assign new_P1_R1117_U388 = ~new_P1_R1117_U127;
  assign new_P1_R1117_U389 = ~new_P1_R1117_U388 | ~new_P1_R1117_U301;
  assign new_P1_R1117_U390 = ~new_P1_R1117_U127 | ~new_P1_R1117_U86;
  assign new_P1_R1117_U391 = ~new_P1_U3975 | ~new_P1_R1117_U83;
  assign new_P1_R1117_U392 = ~new_P1_U3053 | ~new_P1_R1117_U80;
  assign new_P1_R1117_U393 = ~new_P1_U3975 | ~new_P1_R1117_U83;
  assign new_P1_R1117_U394 = ~new_P1_U3053 | ~new_P1_R1117_U80;
  assign new_P1_R1117_U395 = ~new_P1_R1117_U394 | ~new_P1_R1117_U393;
  assign new_P1_R1117_U396 = ~new_P1_U3976 | ~new_P1_R1117_U81;
  assign new_P1_R1117_U397 = ~new_P1_U3057 | ~new_P1_R1117_U44;
  assign new_P1_R1117_U398 = ~new_P1_R1117_U313 | ~new_P1_R1117_U87;
  assign new_P1_R1117_U399 = ~new_P1_R1117_U154 | ~new_P1_R1117_U295;
  assign new_P1_R1117_U400 = ~new_P1_U3977 | ~new_P1_R1117_U79;
  assign new_P1_R1117_U401 = ~new_P1_U3058 | ~new_P1_R1117_U78;
  assign new_P1_R1117_U402 = ~new_P1_R1117_U130;
  assign new_P1_R1117_U403 = ~new_P1_R1117_U291 | ~new_P1_R1117_U402;
  assign new_P1_R1117_U404 = ~new_P1_R1117_U130 | ~new_P1_R1117_U155;
  assign new_P1_R1117_U405 = ~new_P1_U3978 | ~new_P1_R1117_U77;
  assign new_P1_R1117_U406 = ~new_P1_U3065 | ~new_P1_R1117_U76;
  assign new_P1_R1117_U407 = ~new_P1_R1117_U131;
  assign new_P1_R1117_U408 = ~new_P1_R1117_U287 | ~new_P1_R1117_U407;
  assign new_P1_R1117_U409 = ~new_P1_R1117_U131 | ~new_P1_R1117_U156;
  assign new_P1_R1117_U410 = ~new_P1_U3979 | ~new_P1_R1117_U72;
  assign new_P1_R1117_U411 = ~new_P1_U3066 | ~new_P1_R1117_U70;
  assign new_P1_R1117_U412 = ~new_P1_R1117_U411 | ~new_P1_R1117_U410;
  assign new_P1_R1117_U413 = ~new_P1_U3980 | ~new_P1_R1117_U73;
  assign new_P1_R1117_U414 = ~new_P1_U3061 | ~new_P1_R1117_U45;
  assign new_P1_R1117_U415 = ~new_P1_R1117_U323 | ~new_P1_R1117_U88;
  assign new_P1_R1117_U416 = ~new_P1_R1117_U157 | ~new_P1_R1117_U315;
  assign new_P1_R1117_U417 = ~new_P1_U3981 | ~new_P1_R1117_U74;
  assign new_P1_R1117_U418 = ~new_P1_U3075 | ~new_P1_R1117_U71;
  assign new_P1_R1117_U419 = ~new_P1_R1117_U324 | ~new_P1_R1117_U159;
  assign new_P1_R1117_U420 = ~new_P1_R1117_U277 | ~new_P1_R1117_U158;
  assign new_P1_R1117_U421 = ~new_P1_U3982 | ~new_P1_R1117_U69;
  assign new_P1_R1117_U422 = ~new_P1_U3076 | ~new_P1_R1117_U68;
  assign new_P1_R1117_U423 = ~new_P1_R1117_U133;
  assign new_P1_R1117_U424 = ~new_P1_R1117_U273 | ~new_P1_R1117_U423;
  assign new_P1_R1117_U425 = ~new_P1_R1117_U133 | ~new_P1_R1117_U160;
  assign new_P1_R1117_U426 = ~new_P1_R1117_U185 | ~new_P1_R1117_U24;
  assign new_P1_R1117_U427 = ~new_P1_U3078 | ~new_P1_R1117_U23;
  assign new_P1_R1117_U428 = ~new_P1_R1117_U134;
  assign new_P1_R1117_U429 = ~new_P1_U3455 | ~new_P1_R1117_U428;
  assign new_P1_R1117_U430 = ~new_P1_R1117_U134 | ~new_P1_R1117_U161;
  assign new_P1_R1117_U431 = ~new_P1_U3508 | ~new_P1_R1117_U67;
  assign new_P1_R1117_U432 = ~new_P1_U3081 | ~new_P1_R1117_U66;
  assign new_P1_R1117_U433 = ~new_P1_R1117_U135;
  assign new_P1_R1117_U434 = ~new_P1_R1117_U269 | ~new_P1_R1117_U433;
  assign new_P1_R1117_U435 = ~new_P1_R1117_U135 | ~new_P1_R1117_U162;
  assign new_P1_R1117_U436 = ~new_P1_U3506 | ~new_P1_R1117_U65;
  assign new_P1_R1117_U437 = ~new_P1_U3082 | ~new_P1_R1117_U163;
  assign new_P1_R1117_U438 = ~new_P1_R1117_U136;
  assign new_P1_R1117_U439 = ~new_P1_R1117_U438 | ~new_P1_R1117_U265;
  assign new_P1_R1117_U440 = ~new_P1_R1117_U136 | ~new_P1_R1117_U64;
  assign new_P1_R1117_U441 = ~new_P1_U3503 | ~new_P1_R1117_U63;
  assign new_P1_R1117_U442 = ~new_P1_U3069 | ~new_P1_R1117_U62;
  assign new_P1_R1117_U443 = ~new_P1_R1117_U137;
  assign new_P1_R1117_U444 = ~new_P1_R1117_U261 | ~new_P1_R1117_U443;
  assign new_P1_R1117_U445 = ~new_P1_R1117_U137 | ~new_P1_R1117_U164;
  assign new_P1_R1117_U446 = ~new_P1_U3500 | ~new_P1_R1117_U58;
  assign new_P1_R1117_U447 = ~new_P1_U3073 | ~new_P1_R1117_U56;
  assign new_P1_R1117_U448 = ~new_P1_R1117_U447 | ~new_P1_R1117_U446;
  assign new_P1_R1117_U449 = ~new_P1_U3497 | ~new_P1_R1117_U59;
  assign new_P1_R1117_U450 = ~new_P1_U3074 | ~new_P1_R1117_U46;
  assign new_P1_R1117_U451 = ~new_P1_R1117_U334 | ~new_P1_R1117_U89;
  assign new_P1_R1117_U452 = ~new_P1_R1117_U165 | ~new_P1_R1117_U326;
  assign new_P1_R1117_U453 = ~new_P1_U3494 | ~new_P1_R1117_U60;
  assign new_P1_R1117_U454 = ~new_P1_U3079 | ~new_P1_R1117_U57;
  assign new_P1_R1117_U455 = ~new_P1_R1117_U335 | ~new_P1_R1117_U167;
  assign new_P1_R1117_U456 = ~new_P1_R1117_U251 | ~new_P1_R1117_U166;
  assign new_P1_R1117_U457 = ~new_P1_U3491 | ~new_P1_R1117_U55;
  assign new_P1_R1117_U458 = ~new_P1_U3080 | ~new_P1_R1117_U54;
  assign new_P1_R1117_U459 = ~new_P1_R1117_U140;
  assign new_P1_R1117_U460 = ~new_P1_R1117_U247 | ~new_P1_R1117_U459;
  assign new_P1_R1117_U461 = ~new_P1_R1117_U140 | ~new_P1_R1117_U168;
  assign new_P1_R1117_U462 = ~new_P1_U3488 | ~new_P1_R1117_U53;
  assign new_P1_R1117_U463 = ~new_P1_U3072 | ~new_P1_R1117_U52;
  assign new_P1_R1117_U464 = ~new_P1_R1117_U141;
  assign new_P1_R1117_U465 = ~new_P1_R1117_U243 | ~new_P1_R1117_U464;
  assign new_P1_R1117_U466 = ~new_P1_R1117_U141 | ~new_P1_R1117_U169;
  assign new_P1_R1117_U467 = ~new_P1_U3485 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U468 = ~new_P1_U3063 | ~new_P1_R1117_U48;
  assign new_P1_R1117_U469 = ~new_P1_R1117_U468 | ~new_P1_R1117_U467;
  assign new_P1_R1117_U470 = ~new_P1_U3482 | ~new_P1_R1117_U50;
  assign new_P1_R1117_U471 = ~new_P1_U3062 | ~new_P1_R1117_U47;
  assign new_P1_R1117_U472 = ~new_P1_R1117_U345 | ~new_P1_R1117_U90;
  assign new_P1_R1117_U473 = ~new_P1_R1117_U170 | ~new_P1_R1117_U337;
  assign new_P1_R1375_U6 = new_P1_R1375_U119 & new_P1_R1375_U120;
  assign new_P1_R1375_U7 = new_P1_R1375_U137 & new_P1_R1375_U136;
  assign new_P1_R1375_U8 = new_P1_R1375_U141 & new_P1_R1375_U142 & new_P1_R1375_U144 & new_P1_R1375_U143;
  assign new_P1_R1375_U9 = new_P1_R1375_U164 & new_P1_R1375_U163;
  assign new_P1_R1375_U10 = new_P1_R1375_U6 & new_P1_R1375_U198 & new_P1_R1375_U197 & new_P1_R1375_U196;
  assign new_P1_R1375_U11 = new_P1_U3985 & new_P1_R1375_U20;
  assign new_P1_R1375_U12 = new_P1_R1375_U117 & new_P1_R1375_U118 & new_P1_R1375_U207 & new_P1_R1375_U206;
  assign new_P1_R1375_U13 = new_P1_U3450 & new_P1_R1375_U48;
  assign new_P1_R1375_U14 = new_P1_R1375_U204 & new_P1_R1375_U205 & new_P1_R1375_U115;
  assign new_P1_R1375_U15 = ~new_P1_U3983;
  assign new_P1_R1375_U16 = ~new_P1_U3984;
  assign new_P1_R1375_U17 = ~new_P1_U3056;
  assign new_P1_R1375_U18 = ~new_P1_U3985;
  assign new_P1_R1375_U19 = ~new_P1_U3059;
  assign new_P1_R1375_U20 = ~new_P1_U3055;
  assign new_P1_R1375_U21 = ~new_P1_U3054;
  assign new_P1_R1375_U22 = ~new_P1_U3975;
  assign new_P1_R1375_U23 = ~new_P1_U3057;
  assign new_P1_R1375_U24 = ~new_P1_U3977;
  assign new_P1_R1375_U25 = ~new_P1_U3974;
  assign new_P1_R1375_U26 = ~new_P1_U3976;
  assign new_P1_R1375_U27 = ~new_P1_U3978;
  assign new_P1_R1375_U28 = ~new_P1_U3066;
  assign new_P1_R1375_U29 = ~new_P1_U3979;
  assign new_P1_R1375_U30 = ~new_P1_U3061;
  assign new_P1_R1375_U31 = ~new_P1_U3058;
  assign new_P1_R1375_U32 = ~new_P1_U3065;
  assign new_P1_R1375_U33 = ~new_P1_U3075;
  assign new_P1_R1375_U34 = ~new_P1_U3076;
  assign new_P1_R1375_U35 = ~new_P1_U3503;
  assign new_P1_R1375_U36 = ~new_P1_U3506;
  assign new_P1_R1375_U37 = ~new_P1_U3074;
  assign new_P1_R1375_U38 = ~new_P1_U3079;
  assign new_P1_R1375_U39 = ~new_P1_U3470;
  assign new_P1_R1375_U40 = ~new_P1_U3067;
  assign new_P1_R1375_U41 = ~new_P1_U3083;
  assign new_P1_R1375_U42 = ~new_P1_U3084;
  assign new_P1_R1375_U43 = ~new_P1_U3071;
  assign new_P1_R1375_U44 = ~new_P1_U3070;
  assign new_P1_R1375_U45 = ~new_P1_U3060;
  assign new_P1_R1375_U46 = ~new_P1_U3064;
  assign new_P1_R1375_U47 = ~new_P1_U3450;
  assign new_P1_R1375_U48 = ~new_P1_U3077;
  assign new_P1_R1375_U49 = ~new_P1_R1375_U147 | ~new_P1_R1375_U146;
  assign new_P1_R1375_U50 = ~new_P1_U3455;
  assign new_P1_R1375_U51 = ~new_P1_U3068;
  assign new_P1_R1375_U52 = ~new_P1_U3485;
  assign new_P1_R1375_U53 = ~new_P1_U3488;
  assign new_P1_R1375_U54 = ~new_P1_U3458;
  assign new_P1_R1375_U55 = ~new_P1_U3461;
  assign new_P1_R1375_U56 = ~new_P1_U3467;
  assign new_P1_R1375_U57 = ~new_P1_U3464;
  assign new_P1_R1375_U58 = ~new_P1_U3473;
  assign new_P1_R1375_U59 = ~new_P1_U3476;
  assign new_P1_R1375_U60 = ~new_P1_U3479;
  assign new_P1_R1375_U61 = ~new_P1_U3482;
  assign new_P1_R1375_U62 = ~new_P1_U3062;
  assign new_P1_R1375_U63 = ~new_P1_U3072;
  assign new_P1_R1375_U64 = ~new_P1_U3063;
  assign new_P1_R1375_U65 = ~new_P1_U3080;
  assign new_P1_R1375_U66 = ~new_P1_U3491;
  assign new_P1_R1375_U67 = ~new_P1_U3494;
  assign new_P1_R1375_U68 = ~new_P1_U3497;
  assign new_P1_R1375_U69 = ~new_P1_U3500;
  assign new_P1_R1375_U70 = ~new_P1_U3073;
  assign new_P1_R1375_U71 = ~new_P1_U3069;
  assign new_P1_R1375_U72 = ~new_P1_U3082;
  assign new_P1_R1375_U73 = ~new_P1_U3081;
  assign new_P1_R1375_U74 = ~new_P1_U3508;
  assign new_P1_R1375_U75 = ~new_P1_U3982;
  assign new_P1_R1375_U76 = ~new_P1_U3981;
  assign new_P1_R1375_U77 = ~new_P1_U3980;
  assign new_P1_R1375_U78 = ~new_P1_R1375_U11 | ~new_P1_R1375_U125;
  assign new_P1_R1375_U79 = ~new_P1_R1375_U12 | ~new_P1_R1375_U87 | ~new_P1_R1375_U124 | ~new_P1_R1375_U122;
  assign new_P1_R1375_U80 = ~new_P1_R1375_U109 | ~new_P1_R1375_U195;
  assign new_P1_R1375_U81 = new_P1_U3975 & new_P1_R1375_U113;
  assign new_P1_R1375_U82 = new_P1_U3977 & new_P1_R1375_U31;
  assign new_P1_R1375_U83 = new_P1_U3974 & new_P1_R1375_U21;
  assign new_P1_R1375_U84 = new_P1_U3976 & new_P1_R1375_U23;
  assign new_P1_R1375_U85 = new_P1_U3066 & new_P1_R1375_U29;
  assign new_P1_R1375_U86 = new_P1_U3061 & new_P1_R1375_U77;
  assign new_P1_R1375_U87 = new_P1_R1375_U123 & new_P1_R1375_U121;
  assign new_P1_R1375_U88 = new_P1_R1375_U129 & new_P1_R1375_U126;
  assign new_P1_R1375_U89 = new_P1_R1375_U128 & new_P1_R1375_U131 & new_P1_R1375_U201;
  assign new_P1_R1375_U90 = new_P1_U3067 & new_P1_R1375_U56;
  assign new_P1_R1375_U91 = new_P1_R1375_U145 & new_P1_R1375_U149;
  assign new_P1_R1375_U92 = new_P1_R1375_U91 & new_P1_R1375_U140;
  assign new_P1_R1375_U93 = new_P1_R1375_U8 & new_P1_R1375_U153 & new_P1_R1375_U152;
  assign new_P1_R1375_U94 = new_P1_U3458 & new_P1_R1375_U51;
  assign new_P1_R1375_U95 = new_P1_R1375_U159 & new_P1_R1375_U161 & new_P1_R1375_U160;
  assign new_P1_R1375_U96 = new_P1_U3473 & new_P1_R1375_U44;
  assign new_P1_R1375_U97 = new_P1_R1375_U171 & new_P1_R1375_U170;
  assign new_P1_R1375_U98 = new_P1_R1375_U97 & new_P1_R1375_U9;
  assign new_P1_R1375_U99 = new_P1_U3062 & new_P1_R1375_U61;
  assign new_P1_R1375_U100 = new_P1_U3063 & new_P1_R1375_U52;
  assign new_P1_R1375_U101 = new_P1_R1375_U102 & new_P1_R1375_U173 & new_P1_R1375_U174;
  assign new_P1_R1375_U102 = new_P1_R1375_U177 & new_P1_R1375_U176;
  assign new_P1_R1375_U103 = new_P1_R1375_U7 & new_P1_R1375_U104;
  assign new_P1_R1375_U104 = new_P1_R1375_U185 & new_P1_R1375_U186;
  assign new_P1_R1375_U105 = new_P1_U3073 & new_P1_R1375_U69;
  assign new_P1_R1375_U106 = new_P1_U3069 & new_P1_R1375_U35;
  assign new_P1_R1375_U107 = new_P1_R1375_U108 & new_P1_R1375_U188 & new_P1_R1375_U190;
  assign new_P1_R1375_U108 = new_P1_R1375_U192 & new_P1_R1375_U191;
  assign new_P1_R1375_U109 = new_P1_R1375_U134 & new_P1_R1375_U133;
  assign new_P1_R1375_U110 = new_P1_U3982 & new_P1_R1375_U34;
  assign new_P1_R1375_U111 = new_P1_R1375_U128 & new_P1_R1375_U127;
  assign new_P1_R1375_U112 = new_P1_R1375_U130 & new_P1_R1375_U129 & new_P1_R1375_U10 & new_P1_R1375_U131;
  assign new_P1_R1375_U113 = ~new_P1_U3053;
  assign new_P1_R1375_U114 = ~new_P1_R1375_U200 | ~new_P1_R1375_U199;
  assign new_P1_R1375_U115 = ~new_P1_U3983 | ~new_P1_R1375_U17;
  assign new_P1_R1375_U116 = ~new_P1_U3055 | ~new_P1_R1375_U18;
  assign new_P1_R1375_U117 = ~new_P1_U3054 | ~new_P1_R1375_U25;
  assign new_P1_R1375_U118 = ~new_P1_U3057 | ~new_P1_R1375_U26;
  assign new_P1_R1375_U119 = ~new_P1_U3978 | ~new_P1_R1375_U32;
  assign new_P1_R1375_U120 = ~new_P1_U3979 | ~new_P1_R1375_U28;
  assign new_P1_R1375_U121 = ~new_P1_R1375_U85 | ~new_P1_R1375_U119;
  assign new_P1_R1375_U122 = ~new_P1_R1375_U86 | ~new_P1_R1375_U6;
  assign new_P1_R1375_U123 = ~new_P1_U3058 | ~new_P1_R1375_U24;
  assign new_P1_R1375_U124 = ~new_P1_U3065 | ~new_P1_R1375_U27;
  assign new_P1_R1375_U125 = ~new_P1_U3059 | ~new_P1_R1375_U16;
  assign new_P1_R1375_U126 = ~new_P1_R1375_U115 | ~new_P1_R1375_U81 | ~new_P1_R1375_U117;
  assign new_P1_R1375_U127 = ~new_P1_R1375_U115 | ~new_P1_R1375_U82 | ~new_P1_R1375_U12;
  assign new_P1_R1375_U128 = ~new_P1_U3984 | ~new_P1_R1375_U115 | ~new_P1_R1375_U19;
  assign new_P1_R1375_U129 = ~new_P1_R1375_U83 | ~new_P1_R1375_U115;
  assign new_P1_R1375_U130 = ~new_P1_R1375_U115 | ~new_P1_R1375_U84 | ~new_P1_R1375_U12;
  assign new_P1_R1375_U131 = ~new_P1_U3056 | ~new_P1_R1375_U15;
  assign new_P1_R1375_U132 = ~new_P1_R1375_U127 | ~new_P1_R1375_U88 | ~new_P1_R1375_U79 | ~new_P1_R1375_U130;
  assign new_P1_R1375_U133 = ~new_P1_U3075 | ~new_P1_R1375_U76;
  assign new_P1_R1375_U134 = ~new_P1_U3076 | ~new_P1_R1375_U75;
  assign new_P1_R1375_U135 = ~new_P1_U3074 | ~new_P1_R1375_U68;
  assign new_P1_R1375_U136 = ~new_P1_U3503 | ~new_P1_R1375_U71;
  assign new_P1_R1375_U137 = ~new_P1_U3506 | ~new_P1_R1375_U72;
  assign new_P1_R1375_U138 = ~new_P1_U3079 | ~new_P1_R1375_U67;
  assign new_P1_R1375_U139 = ~new_P1_U3470 | ~new_P1_R1375_U43;
  assign new_P1_R1375_U140 = ~new_P1_R1375_U90 | ~new_P1_R1375_U139;
  assign new_P1_R1375_U141 = ~new_P1_U3083 | ~new_P1_R1375_U60;
  assign new_P1_R1375_U142 = ~new_P1_U3084 | ~new_P1_R1375_U59;
  assign new_P1_R1375_U143 = ~new_P1_U3071 | ~new_P1_R1375_U39;
  assign new_P1_R1375_U144 = ~new_P1_U3070 | ~new_P1_R1375_U58;
  assign new_P1_R1375_U145 = ~new_P1_U3060 | ~new_P1_R1375_U57;
  assign new_P1_R1375_U146 = new_P1_U3447 | new_P1_R1375_U13;
  assign new_P1_R1375_U147 = ~new_P1_U3077 | ~new_P1_R1375_U47;
  assign new_P1_R1375_U148 = ~new_P1_R1375_U49;
  assign new_P1_R1375_U149 = ~new_P1_U3064 | ~new_P1_R1375_U55;
  assign new_P1_R1375_U150 = ~new_P1_U3455 | ~new_P1_R1375_U148;
  assign new_P1_R1375_U151 = ~new_P1_U3078 | ~new_P1_R1375_U150;
  assign new_P1_R1375_U152 = ~new_P1_R1375_U49 | ~new_P1_R1375_U50;
  assign new_P1_R1375_U153 = ~new_P1_U3068 | ~new_P1_R1375_U54;
  assign new_P1_R1375_U154 = ~new_P1_R1375_U93 | ~new_P1_R1375_U92 | ~new_P1_R1375_U151;
  assign new_P1_R1375_U155 = ~new_P1_R1375_U94 | ~new_P1_R1375_U149;
  assign new_P1_R1375_U156 = ~new_P1_U3461 | ~new_P1_R1375_U46;
  assign new_P1_R1375_U157 = ~new_P1_R1375_U156 | ~new_P1_R1375_U155;
  assign new_P1_R1375_U158 = ~new_P1_R1375_U157 | ~new_P1_R1375_U145;
  assign new_P1_R1375_U159 = ~new_P1_U3467 | ~new_P1_R1375_U40;
  assign new_P1_R1375_U160 = ~new_P1_U3464 | ~new_P1_R1375_U45;
  assign new_P1_R1375_U161 = ~new_P1_U3470 | ~new_P1_R1375_U43;
  assign new_P1_R1375_U162 = ~new_P1_R1375_U158 | ~new_P1_R1375_U95;
  assign new_P1_R1375_U163 = ~new_P1_U3485 | ~new_P1_R1375_U64;
  assign new_P1_R1375_U164 = ~new_P1_U3488 | ~new_P1_R1375_U63;
  assign new_P1_R1375_U165 = ~new_P1_R1375_U96 | ~new_P1_R1375_U142;
  assign new_P1_R1375_U166 = ~new_P1_U3476 | ~new_P1_R1375_U42;
  assign new_P1_R1375_U167 = ~new_P1_R1375_U166 | ~new_P1_R1375_U165;
  assign new_P1_R1375_U168 = ~new_P1_R1375_U8 | ~new_P1_R1375_U162 | ~new_P1_R1375_U140;
  assign new_P1_R1375_U169 = ~new_P1_R1375_U167 | ~new_P1_R1375_U141;
  assign new_P1_R1375_U170 = ~new_P1_U3479 | ~new_P1_R1375_U41;
  assign new_P1_R1375_U171 = ~new_P1_U3482 | ~new_P1_R1375_U62;
  assign new_P1_R1375_U172 = ~new_P1_R1375_U154 | ~new_P1_R1375_U98 | ~new_P1_R1375_U168 | ~new_P1_R1375_U169;
  assign new_P1_R1375_U173 = ~new_P1_R1375_U99 | ~new_P1_R1375_U9;
  assign new_P1_R1375_U174 = ~new_P1_U3072 | ~new_P1_R1375_U53;
  assign new_P1_R1375_U175 = ~new_P1_U3488 | ~new_P1_R1375_U63;
  assign new_P1_R1375_U176 = ~new_P1_R1375_U100 | ~new_P1_R1375_U175;
  assign new_P1_R1375_U177 = ~new_P1_U3080 | ~new_P1_R1375_U66;
  assign new_P1_R1375_U178 = ~new_P1_R1375_U172 | ~new_P1_R1375_U101;
  assign new_P1_R1375_U179 = ~new_P1_U3491 | ~new_P1_R1375_U65;
  assign new_P1_R1375_U180 = ~new_P1_R1375_U179 | ~new_P1_R1375_U178;
  assign new_P1_R1375_U181 = ~new_P1_R1375_U180 | ~new_P1_R1375_U138;
  assign new_P1_R1375_U182 = ~new_P1_U3494 | ~new_P1_R1375_U38;
  assign new_P1_R1375_U183 = ~new_P1_R1375_U182 | ~new_P1_R1375_U181;
  assign new_P1_R1375_U184 = ~new_P1_R1375_U183 | ~new_P1_R1375_U135;
  assign new_P1_R1375_U185 = ~new_P1_U3497 | ~new_P1_R1375_U37;
  assign new_P1_R1375_U186 = ~new_P1_U3500 | ~new_P1_R1375_U70;
  assign new_P1_R1375_U187 = ~new_P1_R1375_U184 | ~new_P1_R1375_U103;
  assign new_P1_R1375_U188 = ~new_P1_R1375_U105 | ~new_P1_R1375_U7;
  assign new_P1_R1375_U189 = ~new_P1_U3506 | ~new_P1_R1375_U72;
  assign new_P1_R1375_U190 = ~new_P1_R1375_U106 | ~new_P1_R1375_U189;
  assign new_P1_R1375_U191 = ~new_P1_U3082 | ~new_P1_R1375_U36;
  assign new_P1_R1375_U192 = ~new_P1_U3081 | ~new_P1_R1375_U74;
  assign new_P1_R1375_U193 = ~new_P1_R1375_U187 | ~new_P1_R1375_U107;
  assign new_P1_R1375_U194 = ~new_P1_U3508 | ~new_P1_R1375_U73;
  assign new_P1_R1375_U195 = ~new_P1_R1375_U194 | ~new_P1_R1375_U193;
  assign new_P1_R1375_U196 = ~new_P1_R1375_U110 | ~new_P1_R1375_U133;
  assign new_P1_R1375_U197 = ~new_P1_U3981 | ~new_P1_R1375_U33;
  assign new_P1_R1375_U198 = ~new_P1_U3980 | ~new_P1_R1375_U30;
  assign new_P1_R1375_U199 = ~new_P1_U3984 | ~new_P1_R1375_U116;
  assign new_P1_R1375_U200 = ~new_P1_R1375_U19 | ~new_P1_R1375_U116;
  assign new_P1_R1375_U201 = ~new_P1_R1375_U11 | ~new_P1_R1375_U202;
  assign new_P1_R1375_U202 = ~new_P1_U3059 | ~new_P1_R1375_U16;
  assign new_P1_R1375_U203 = ~new_P1_R1375_U132 | ~new_P1_R1375_U114;
  assign new_P1_R1375_U204 = ~new_P1_R1375_U89 | ~new_P1_R1375_U203;
  assign new_P1_R1375_U205 = ~new_P1_R1375_U112 | ~new_P1_R1375_U111 | ~new_P1_R1375_U78 | ~new_P1_R1375_U126 | ~new_P1_R1375_U80;
  assign new_P1_R1375_U206 = ~new_P1_U3053 | ~new_P1_R1375_U22;
  assign new_P1_R1375_U207 = ~new_P1_U3975 | ~new_P1_R1375_U113;
  assign new_P1_R1352_U6 = new_P1_U3059 & new_P1_R1352_U7;
  assign new_P1_R1352_U7 = ~new_P1_U3056;
  assign new_P1_R1207_U6 = new_P1_R1207_U198 & new_P1_R1207_U197;
  assign new_P1_R1207_U7 = new_P1_R1207_U237 & new_P1_R1207_U236;
  assign new_P1_R1207_U8 = new_P1_R1207_U254 & new_P1_R1207_U253;
  assign new_P1_R1207_U9 = new_P1_R1207_U280 & new_P1_R1207_U279;
  assign new_P1_R1207_U10 = ~new_P1_R1207_U340 | ~new_P1_R1207_U343;
  assign new_P1_R1207_U11 = ~new_P1_R1207_U329 | ~new_P1_R1207_U332;
  assign new_P1_R1207_U12 = ~new_P1_R1207_U318 | ~new_P1_R1207_U321;
  assign new_P1_R1207_U13 = ~new_P1_R1207_U310 | ~new_P1_R1207_U312;
  assign new_P1_R1207_U14 = ~new_P1_R1207_U347 | ~new_P1_R1207_U308;
  assign new_P1_R1207_U15 = ~new_P1_R1207_U231 | ~new_P1_R1207_U233;
  assign new_P1_R1207_U16 = ~new_P1_R1207_U223 | ~new_P1_R1207_U226;
  assign new_P1_R1207_U17 = ~new_P1_R1207_U215 | ~new_P1_R1207_U217;
  assign new_P1_R1207_U18 = ~new_P1_R1207_U23 | ~new_P1_R1207_U346;
  assign new_P1_R1207_U19 = ~new_P1_U3473;
  assign new_P1_R1207_U20 = ~new_P1_U3467;
  assign new_P1_R1207_U21 = ~new_P1_U3458;
  assign new_P1_R1207_U22 = ~new_P1_U3450;
  assign new_P1_R1207_U23 = ~new_P1_U3450 | ~new_P1_R1207_U91;
  assign new_P1_R1207_U24 = ~new_P1_U3078;
  assign new_P1_R1207_U25 = ~new_P1_U3461;
  assign new_P1_R1207_U26 = ~new_P1_U3068;
  assign new_P1_R1207_U27 = ~new_P1_U3068 | ~new_P1_R1207_U21;
  assign new_P1_R1207_U28 = ~new_P1_U3064;
  assign new_P1_R1207_U29 = ~new_P1_U3470;
  assign new_P1_R1207_U30 = ~new_P1_U3464;
  assign new_P1_R1207_U31 = ~new_P1_U3071;
  assign new_P1_R1207_U32 = ~new_P1_U3067;
  assign new_P1_R1207_U33 = ~new_P1_U3060;
  assign new_P1_R1207_U34 = ~new_P1_U3060 | ~new_P1_R1207_U30;
  assign new_P1_R1207_U35 = ~new_P1_U3476;
  assign new_P1_R1207_U36 = ~new_P1_U3070;
  assign new_P1_R1207_U37 = ~new_P1_U3070 | ~new_P1_R1207_U19;
  assign new_P1_R1207_U38 = ~new_P1_U3084;
  assign new_P1_R1207_U39 = ~new_P1_U3479;
  assign new_P1_R1207_U40 = ~new_P1_U3083;
  assign new_P1_R1207_U41 = ~new_P1_R1207_U204 | ~new_P1_R1207_U203;
  assign new_P1_R1207_U42 = ~new_P1_R1207_U34 | ~new_P1_R1207_U219;
  assign new_P1_R1207_U43 = ~new_P1_R1207_U188 | ~new_P1_R1207_U187;
  assign new_P1_R1207_U44 = ~new_P1_U3976;
  assign new_P1_R1207_U45 = ~new_P1_U3980;
  assign new_P1_R1207_U46 = ~new_P1_U3497;
  assign new_P1_R1207_U47 = ~new_P1_U3482;
  assign new_P1_R1207_U48 = ~new_P1_U3485;
  assign new_P1_R1207_U49 = ~new_P1_U3063;
  assign new_P1_R1207_U50 = ~new_P1_U3062;
  assign new_P1_R1207_U51 = ~new_P1_U3083 | ~new_P1_R1207_U39;
  assign new_P1_R1207_U52 = ~new_P1_U3488;
  assign new_P1_R1207_U53 = ~new_P1_U3072;
  assign new_P1_R1207_U54 = ~new_P1_U3491;
  assign new_P1_R1207_U55 = ~new_P1_U3080;
  assign new_P1_R1207_U56 = ~new_P1_U3500;
  assign new_P1_R1207_U57 = ~new_P1_U3494;
  assign new_P1_R1207_U58 = ~new_P1_U3073;
  assign new_P1_R1207_U59 = ~new_P1_U3074;
  assign new_P1_R1207_U60 = ~new_P1_U3079;
  assign new_P1_R1207_U61 = ~new_P1_U3079 | ~new_P1_R1207_U57;
  assign new_P1_R1207_U62 = ~new_P1_U3503;
  assign new_P1_R1207_U63 = ~new_P1_U3069;
  assign new_P1_R1207_U64 = ~new_P1_R1207_U264 | ~new_P1_R1207_U263;
  assign new_P1_R1207_U65 = ~new_P1_U3082;
  assign new_P1_R1207_U66 = ~new_P1_U3508;
  assign new_P1_R1207_U67 = ~new_P1_U3081;
  assign new_P1_R1207_U68 = ~new_P1_U3982;
  assign new_P1_R1207_U69 = ~new_P1_U3076;
  assign new_P1_R1207_U70 = ~new_P1_U3979;
  assign new_P1_R1207_U71 = ~new_P1_U3981;
  assign new_P1_R1207_U72 = ~new_P1_U3066;
  assign new_P1_R1207_U73 = ~new_P1_U3061;
  assign new_P1_R1207_U74 = ~new_P1_U3075;
  assign new_P1_R1207_U75 = ~new_P1_U3075 | ~new_P1_R1207_U71;
  assign new_P1_R1207_U76 = ~new_P1_U3978;
  assign new_P1_R1207_U77 = ~new_P1_U3065;
  assign new_P1_R1207_U78 = ~new_P1_U3977;
  assign new_P1_R1207_U79 = ~new_P1_U3058;
  assign new_P1_R1207_U80 = ~new_P1_U3975;
  assign new_P1_R1207_U81 = ~new_P1_U3057;
  assign new_P1_R1207_U82 = ~new_P1_U3057 | ~new_P1_R1207_U44;
  assign new_P1_R1207_U83 = ~new_P1_U3053;
  assign new_P1_R1207_U84 = ~new_P1_U3974;
  assign new_P1_R1207_U85 = ~new_P1_U3054;
  assign new_P1_R1207_U86 = ~new_P1_R1207_U126 | ~new_P1_R1207_U297;
  assign new_P1_R1207_U87 = ~new_P1_R1207_U294 | ~new_P1_R1207_U293;
  assign new_P1_R1207_U88 = ~new_P1_R1207_U75 | ~new_P1_R1207_U314;
  assign new_P1_R1207_U89 = ~new_P1_R1207_U61 | ~new_P1_R1207_U325;
  assign new_P1_R1207_U90 = ~new_P1_R1207_U51 | ~new_P1_R1207_U336;
  assign new_P1_R1207_U91 = ~new_P1_U3077;
  assign new_P1_R1207_U92 = ~new_P1_R1207_U390 | ~new_P1_R1207_U389;
  assign new_P1_R1207_U93 = ~new_P1_R1207_U404 | ~new_P1_R1207_U403;
  assign new_P1_R1207_U94 = ~new_P1_R1207_U409 | ~new_P1_R1207_U408;
  assign new_P1_R1207_U95 = ~new_P1_R1207_U425 | ~new_P1_R1207_U424;
  assign new_P1_R1207_U96 = ~new_P1_R1207_U430 | ~new_P1_R1207_U429;
  assign new_P1_R1207_U97 = ~new_P1_R1207_U435 | ~new_P1_R1207_U434;
  assign new_P1_R1207_U98 = ~new_P1_R1207_U440 | ~new_P1_R1207_U439;
  assign new_P1_R1207_U99 = ~new_P1_R1207_U445 | ~new_P1_R1207_U444;
  assign new_P1_R1207_U100 = ~new_P1_R1207_U461 | ~new_P1_R1207_U460;
  assign new_P1_R1207_U101 = ~new_P1_R1207_U466 | ~new_P1_R1207_U465;
  assign new_P1_R1207_U102 = ~new_P1_R1207_U351 | ~new_P1_R1207_U350;
  assign new_P1_R1207_U103 = ~new_P1_R1207_U360 | ~new_P1_R1207_U359;
  assign new_P1_R1207_U104 = ~new_P1_R1207_U367 | ~new_P1_R1207_U366;
  assign new_P1_R1207_U105 = ~new_P1_R1207_U371 | ~new_P1_R1207_U370;
  assign new_P1_R1207_U106 = ~new_P1_R1207_U380 | ~new_P1_R1207_U379;
  assign new_P1_R1207_U107 = ~new_P1_R1207_U399 | ~new_P1_R1207_U398;
  assign new_P1_R1207_U108 = ~new_P1_R1207_U416 | ~new_P1_R1207_U415;
  assign new_P1_R1207_U109 = ~new_P1_R1207_U420 | ~new_P1_R1207_U419;
  assign new_P1_R1207_U110 = ~new_P1_R1207_U452 | ~new_P1_R1207_U451;
  assign new_P1_R1207_U111 = ~new_P1_R1207_U456 | ~new_P1_R1207_U455;
  assign new_P1_R1207_U112 = ~new_P1_R1207_U473 | ~new_P1_R1207_U472;
  assign new_P1_R1207_U113 = new_P1_R1207_U193 & new_P1_R1207_U194;
  assign new_P1_R1207_U114 = new_P1_R1207_U201 & new_P1_R1207_U196;
  assign new_P1_R1207_U115 = new_P1_R1207_U206 & new_P1_R1207_U180;
  assign new_P1_R1207_U116 = new_P1_R1207_U209 & new_P1_R1207_U210;
  assign new_P1_R1207_U117 = new_P1_R1207_U37 & new_P1_R1207_U353 & new_P1_R1207_U352;
  assign new_P1_R1207_U118 = new_P1_R1207_U356 & new_P1_R1207_U180;
  assign new_P1_R1207_U119 = new_P1_R1207_U225 & new_P1_R1207_U6;
  assign new_P1_R1207_U120 = new_P1_R1207_U363 & new_P1_R1207_U179;
  assign new_P1_R1207_U121 = new_P1_R1207_U27 & new_P1_R1207_U373 & new_P1_R1207_U372;
  assign new_P1_R1207_U122 = new_P1_R1207_U376 & new_P1_R1207_U178;
  assign new_P1_R1207_U123 = new_P1_R1207_U174 & new_P1_R1207_U235 & new_P1_R1207_U212;
  assign new_P1_R1207_U124 = new_P1_R1207_U252 & new_P1_R1207_U257 & new_P1_R1207_U175;
  assign new_P1_R1207_U125 = new_P1_R1207_U283 & new_P1_R1207_U176;
  assign new_P1_R1207_U126 = new_P1_R1207_U299 & new_P1_R1207_U300;
  assign new_P1_R1207_U127 = ~new_P1_R1207_U387 | ~new_P1_R1207_U386;
  assign new_P1_R1207_U128 = new_P1_R1207_U82 & new_P1_R1207_U392 & new_P1_R1207_U391;
  assign new_P1_R1207_U129 = new_P1_R1207_U395 & new_P1_R1207_U177;
  assign new_P1_R1207_U130 = ~new_P1_R1207_U401 | ~new_P1_R1207_U400;
  assign new_P1_R1207_U131 = ~new_P1_R1207_U406 | ~new_P1_R1207_U405;
  assign new_P1_R1207_U132 = new_P1_R1207_U412 & new_P1_R1207_U176;
  assign new_P1_R1207_U133 = ~new_P1_R1207_U422 | ~new_P1_R1207_U421;
  assign new_P1_R1207_U134 = ~new_P1_R1207_U427 | ~new_P1_R1207_U426;
  assign new_P1_R1207_U135 = ~new_P1_R1207_U432 | ~new_P1_R1207_U431;
  assign new_P1_R1207_U136 = ~new_P1_R1207_U437 | ~new_P1_R1207_U436;
  assign new_P1_R1207_U137 = ~new_P1_R1207_U442 | ~new_P1_R1207_U441;
  assign new_P1_R1207_U138 = new_P1_R1207_U331 & new_P1_R1207_U8;
  assign new_P1_R1207_U139 = new_P1_R1207_U448 & new_P1_R1207_U175;
  assign new_P1_R1207_U140 = ~new_P1_R1207_U458 | ~new_P1_R1207_U457;
  assign new_P1_R1207_U141 = ~new_P1_R1207_U463 | ~new_P1_R1207_U462;
  assign new_P1_R1207_U142 = new_P1_R1207_U342 & new_P1_R1207_U7;
  assign new_P1_R1207_U143 = new_P1_R1207_U469 & new_P1_R1207_U174;
  assign new_P1_R1207_U144 = new_P1_R1207_U349 & new_P1_R1207_U348;
  assign new_P1_R1207_U145 = ~new_P1_R1207_U116 | ~new_P1_R1207_U207;
  assign new_P1_R1207_U146 = new_P1_R1207_U358 & new_P1_R1207_U357;
  assign new_P1_R1207_U147 = new_P1_R1207_U365 & new_P1_R1207_U364;
  assign new_P1_R1207_U148 = new_P1_R1207_U369 & new_P1_R1207_U368;
  assign new_P1_R1207_U149 = ~new_P1_R1207_U113 | ~new_P1_R1207_U191;
  assign new_P1_R1207_U150 = new_P1_R1207_U378 & new_P1_R1207_U377;
  assign new_P1_R1207_U151 = ~new_P1_U3985;
  assign new_P1_R1207_U152 = ~new_P1_U3055;
  assign new_P1_R1207_U153 = new_P1_R1207_U382 & new_P1_R1207_U381;
  assign new_P1_R1207_U154 = new_P1_R1207_U397 & new_P1_R1207_U396;
  assign new_P1_R1207_U155 = ~new_P1_R1207_U290 | ~new_P1_R1207_U289;
  assign new_P1_R1207_U156 = ~new_P1_R1207_U286 | ~new_P1_R1207_U285;
  assign new_P1_R1207_U157 = new_P1_R1207_U414 & new_P1_R1207_U413;
  assign new_P1_R1207_U158 = new_P1_R1207_U418 & new_P1_R1207_U417;
  assign new_P1_R1207_U159 = ~new_P1_R1207_U276 | ~new_P1_R1207_U275;
  assign new_P1_R1207_U160 = ~new_P1_R1207_U272 | ~new_P1_R1207_U271;
  assign new_P1_R1207_U161 = ~new_P1_U3455;
  assign new_P1_R1207_U162 = ~new_P1_R1207_U268 | ~new_P1_R1207_U267;
  assign new_P1_R1207_U163 = ~new_P1_U3506;
  assign new_P1_R1207_U164 = ~new_P1_R1207_U260 | ~new_P1_R1207_U259;
  assign new_P1_R1207_U165 = new_P1_R1207_U450 & new_P1_R1207_U449;
  assign new_P1_R1207_U166 = new_P1_R1207_U454 & new_P1_R1207_U453;
  assign new_P1_R1207_U167 = ~new_P1_R1207_U250 | ~new_P1_R1207_U249;
  assign new_P1_R1207_U168 = ~new_P1_R1207_U246 | ~new_P1_R1207_U245;
  assign new_P1_R1207_U169 = ~new_P1_R1207_U242 | ~new_P1_R1207_U241;
  assign new_P1_R1207_U170 = new_P1_R1207_U471 & new_P1_R1207_U470;
  assign new_P1_R1207_U171 = ~new_P1_R1207_U82;
  assign new_P1_R1207_U172 = ~new_P1_R1207_U27;
  assign new_P1_R1207_U173 = ~new_P1_R1207_U37;
  assign new_P1_R1207_U174 = ~new_P1_U3482 | ~new_P1_R1207_U50;
  assign new_P1_R1207_U175 = ~new_P1_U3497 | ~new_P1_R1207_U59;
  assign new_P1_R1207_U176 = ~new_P1_U3980 | ~new_P1_R1207_U73;
  assign new_P1_R1207_U177 = ~new_P1_U3976 | ~new_P1_R1207_U81;
  assign new_P1_R1207_U178 = ~new_P1_U3458 | ~new_P1_R1207_U26;
  assign new_P1_R1207_U179 = ~new_P1_U3467 | ~new_P1_R1207_U32;
  assign new_P1_R1207_U180 = ~new_P1_U3473 | ~new_P1_R1207_U36;
  assign new_P1_R1207_U181 = ~new_P1_R1207_U61;
  assign new_P1_R1207_U182 = ~new_P1_R1207_U75;
  assign new_P1_R1207_U183 = ~new_P1_R1207_U34;
  assign new_P1_R1207_U184 = ~new_P1_R1207_U51;
  assign new_P1_R1207_U185 = ~new_P1_R1207_U23;
  assign new_P1_R1207_U186 = ~new_P1_R1207_U185 | ~new_P1_R1207_U24;
  assign new_P1_R1207_U187 = ~new_P1_R1207_U186 | ~new_P1_R1207_U161;
  assign new_P1_R1207_U188 = ~new_P1_U3078 | ~new_P1_R1207_U23;
  assign new_P1_R1207_U189 = ~new_P1_R1207_U43;
  assign new_P1_R1207_U190 = ~new_P1_U3461 | ~new_P1_R1207_U28;
  assign new_P1_R1207_U191 = ~new_P1_R1207_U190 | ~new_P1_R1207_U43 | ~new_P1_R1207_U178;
  assign new_P1_R1207_U192 = ~new_P1_R1207_U28 | ~new_P1_R1207_U27;
  assign new_P1_R1207_U193 = ~new_P1_R1207_U192 | ~new_P1_R1207_U25;
  assign new_P1_R1207_U194 = ~new_P1_U3064 | ~new_P1_R1207_U172;
  assign new_P1_R1207_U195 = ~new_P1_R1207_U149;
  assign new_P1_R1207_U196 = ~new_P1_U3470 | ~new_P1_R1207_U31;
  assign new_P1_R1207_U197 = ~new_P1_U3071 | ~new_P1_R1207_U29;
  assign new_P1_R1207_U198 = ~new_P1_U3067 | ~new_P1_R1207_U20;
  assign new_P1_R1207_U199 = ~new_P1_R1207_U183 | ~new_P1_R1207_U179;
  assign new_P1_R1207_U200 = ~new_P1_R1207_U6 | ~new_P1_R1207_U199;
  assign new_P1_R1207_U201 = ~new_P1_U3464 | ~new_P1_R1207_U33;
  assign new_P1_R1207_U202 = ~new_P1_U3470 | ~new_P1_R1207_U31;
  assign new_P1_R1207_U203 = ~new_P1_R1207_U114 | ~new_P1_R1207_U149 | ~new_P1_R1207_U179;
  assign new_P1_R1207_U204 = ~new_P1_R1207_U202 | ~new_P1_R1207_U200;
  assign new_P1_R1207_U205 = ~new_P1_R1207_U41;
  assign new_P1_R1207_U206 = ~new_P1_U3476 | ~new_P1_R1207_U38;
  assign new_P1_R1207_U207 = ~new_P1_R1207_U115 | ~new_P1_R1207_U41;
  assign new_P1_R1207_U208 = ~new_P1_R1207_U38 | ~new_P1_R1207_U37;
  assign new_P1_R1207_U209 = ~new_P1_R1207_U208 | ~new_P1_R1207_U35;
  assign new_P1_R1207_U210 = ~new_P1_U3084 | ~new_P1_R1207_U173;
  assign new_P1_R1207_U211 = ~new_P1_R1207_U145;
  assign new_P1_R1207_U212 = ~new_P1_U3479 | ~new_P1_R1207_U40;
  assign new_P1_R1207_U213 = ~new_P1_R1207_U212 | ~new_P1_R1207_U51;
  assign new_P1_R1207_U214 = ~new_P1_R1207_U205 | ~new_P1_R1207_U37;
  assign new_P1_R1207_U215 = ~new_P1_R1207_U118 | ~new_P1_R1207_U214;
  assign new_P1_R1207_U216 = ~new_P1_R1207_U41 | ~new_P1_R1207_U180;
  assign new_P1_R1207_U217 = ~new_P1_R1207_U117 | ~new_P1_R1207_U216;
  assign new_P1_R1207_U218 = ~new_P1_R1207_U37 | ~new_P1_R1207_U180;
  assign new_P1_R1207_U219 = ~new_P1_R1207_U201 | ~new_P1_R1207_U149;
  assign new_P1_R1207_U220 = ~new_P1_R1207_U42;
  assign new_P1_R1207_U221 = ~new_P1_U3067 | ~new_P1_R1207_U20;
  assign new_P1_R1207_U222 = ~new_P1_R1207_U220 | ~new_P1_R1207_U221;
  assign new_P1_R1207_U223 = ~new_P1_R1207_U120 | ~new_P1_R1207_U222;
  assign new_P1_R1207_U224 = ~new_P1_R1207_U42 | ~new_P1_R1207_U179;
  assign new_P1_R1207_U225 = ~new_P1_U3470 | ~new_P1_R1207_U31;
  assign new_P1_R1207_U226 = ~new_P1_R1207_U119 | ~new_P1_R1207_U224;
  assign new_P1_R1207_U227 = ~new_P1_U3067 | ~new_P1_R1207_U20;
  assign new_P1_R1207_U228 = ~new_P1_R1207_U179 | ~new_P1_R1207_U227;
  assign new_P1_R1207_U229 = ~new_P1_R1207_U201 | ~new_P1_R1207_U34;
  assign new_P1_R1207_U230 = ~new_P1_R1207_U189 | ~new_P1_R1207_U27;
  assign new_P1_R1207_U231 = ~new_P1_R1207_U122 | ~new_P1_R1207_U230;
  assign new_P1_R1207_U232 = ~new_P1_R1207_U43 | ~new_P1_R1207_U178;
  assign new_P1_R1207_U233 = ~new_P1_R1207_U121 | ~new_P1_R1207_U232;
  assign new_P1_R1207_U234 = ~new_P1_R1207_U27 | ~new_P1_R1207_U178;
  assign new_P1_R1207_U235 = ~new_P1_U3485 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U236 = ~new_P1_U3063 | ~new_P1_R1207_U48;
  assign new_P1_R1207_U237 = ~new_P1_U3062 | ~new_P1_R1207_U47;
  assign new_P1_R1207_U238 = ~new_P1_R1207_U184 | ~new_P1_R1207_U174;
  assign new_P1_R1207_U239 = ~new_P1_R1207_U7 | ~new_P1_R1207_U238;
  assign new_P1_R1207_U240 = ~new_P1_U3485 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U241 = ~new_P1_R1207_U145 | ~new_P1_R1207_U123;
  assign new_P1_R1207_U242 = ~new_P1_R1207_U240 | ~new_P1_R1207_U239;
  assign new_P1_R1207_U243 = ~new_P1_R1207_U169;
  assign new_P1_R1207_U244 = ~new_P1_U3488 | ~new_P1_R1207_U53;
  assign new_P1_R1207_U245 = ~new_P1_R1207_U244 | ~new_P1_R1207_U169;
  assign new_P1_R1207_U246 = ~new_P1_U3072 | ~new_P1_R1207_U52;
  assign new_P1_R1207_U247 = ~new_P1_R1207_U168;
  assign new_P1_R1207_U248 = ~new_P1_U3491 | ~new_P1_R1207_U55;
  assign new_P1_R1207_U249 = ~new_P1_R1207_U248 | ~new_P1_R1207_U168;
  assign new_P1_R1207_U250 = ~new_P1_U3080 | ~new_P1_R1207_U54;
  assign new_P1_R1207_U251 = ~new_P1_R1207_U167;
  assign new_P1_R1207_U252 = ~new_P1_U3500 | ~new_P1_R1207_U58;
  assign new_P1_R1207_U253 = ~new_P1_U3073 | ~new_P1_R1207_U56;
  assign new_P1_R1207_U254 = ~new_P1_U3074 | ~new_P1_R1207_U46;
  assign new_P1_R1207_U255 = ~new_P1_R1207_U181 | ~new_P1_R1207_U175;
  assign new_P1_R1207_U256 = ~new_P1_R1207_U8 | ~new_P1_R1207_U255;
  assign new_P1_R1207_U257 = ~new_P1_U3494 | ~new_P1_R1207_U60;
  assign new_P1_R1207_U258 = ~new_P1_U3500 | ~new_P1_R1207_U58;
  assign new_P1_R1207_U259 = ~new_P1_R1207_U167 | ~new_P1_R1207_U124;
  assign new_P1_R1207_U260 = ~new_P1_R1207_U258 | ~new_P1_R1207_U256;
  assign new_P1_R1207_U261 = ~new_P1_R1207_U164;
  assign new_P1_R1207_U262 = ~new_P1_U3503 | ~new_P1_R1207_U63;
  assign new_P1_R1207_U263 = ~new_P1_R1207_U262 | ~new_P1_R1207_U164;
  assign new_P1_R1207_U264 = ~new_P1_U3069 | ~new_P1_R1207_U62;
  assign new_P1_R1207_U265 = ~new_P1_R1207_U64;
  assign new_P1_R1207_U266 = ~new_P1_R1207_U265 | ~new_P1_R1207_U65;
  assign new_P1_R1207_U267 = ~new_P1_R1207_U266 | ~new_P1_R1207_U163;
  assign new_P1_R1207_U268 = ~new_P1_U3082 | ~new_P1_R1207_U64;
  assign new_P1_R1207_U269 = ~new_P1_R1207_U162;
  assign new_P1_R1207_U270 = ~new_P1_U3508 | ~new_P1_R1207_U67;
  assign new_P1_R1207_U271 = ~new_P1_R1207_U270 | ~new_P1_R1207_U162;
  assign new_P1_R1207_U272 = ~new_P1_U3081 | ~new_P1_R1207_U66;
  assign new_P1_R1207_U273 = ~new_P1_R1207_U160;
  assign new_P1_R1207_U274 = ~new_P1_U3982 | ~new_P1_R1207_U69;
  assign new_P1_R1207_U275 = ~new_P1_R1207_U274 | ~new_P1_R1207_U160;
  assign new_P1_R1207_U276 = ~new_P1_U3076 | ~new_P1_R1207_U68;
  assign new_P1_R1207_U277 = ~new_P1_R1207_U159;
  assign new_P1_R1207_U278 = ~new_P1_U3979 | ~new_P1_R1207_U72;
  assign new_P1_R1207_U279 = ~new_P1_U3066 | ~new_P1_R1207_U70;
  assign new_P1_R1207_U280 = ~new_P1_U3061 | ~new_P1_R1207_U45;
  assign new_P1_R1207_U281 = ~new_P1_R1207_U182 | ~new_P1_R1207_U176;
  assign new_P1_R1207_U282 = ~new_P1_R1207_U9 | ~new_P1_R1207_U281;
  assign new_P1_R1207_U283 = ~new_P1_U3981 | ~new_P1_R1207_U74;
  assign new_P1_R1207_U284 = ~new_P1_U3979 | ~new_P1_R1207_U72;
  assign new_P1_R1207_U285 = ~new_P1_R1207_U278 | ~new_P1_R1207_U159 | ~new_P1_R1207_U125;
  assign new_P1_R1207_U286 = ~new_P1_R1207_U284 | ~new_P1_R1207_U282;
  assign new_P1_R1207_U287 = ~new_P1_R1207_U156;
  assign new_P1_R1207_U288 = ~new_P1_U3978 | ~new_P1_R1207_U77;
  assign new_P1_R1207_U289 = ~new_P1_R1207_U288 | ~new_P1_R1207_U156;
  assign new_P1_R1207_U290 = ~new_P1_U3065 | ~new_P1_R1207_U76;
  assign new_P1_R1207_U291 = ~new_P1_R1207_U155;
  assign new_P1_R1207_U292 = ~new_P1_U3977 | ~new_P1_R1207_U79;
  assign new_P1_R1207_U293 = ~new_P1_R1207_U292 | ~new_P1_R1207_U155;
  assign new_P1_R1207_U294 = ~new_P1_U3058 | ~new_P1_R1207_U78;
  assign new_P1_R1207_U295 = ~new_P1_R1207_U87;
  assign new_P1_R1207_U296 = ~new_P1_U3975 | ~new_P1_R1207_U83;
  assign new_P1_R1207_U297 = ~new_P1_R1207_U296 | ~new_P1_R1207_U87 | ~new_P1_R1207_U177;
  assign new_P1_R1207_U298 = ~new_P1_R1207_U83 | ~new_P1_R1207_U82;
  assign new_P1_R1207_U299 = ~new_P1_R1207_U298 | ~new_P1_R1207_U80;
  assign new_P1_R1207_U300 = ~new_P1_U3053 | ~new_P1_R1207_U171;
  assign new_P1_R1207_U301 = ~new_P1_R1207_U86;
  assign new_P1_R1207_U302 = ~new_P1_U3054 | ~new_P1_R1207_U84;
  assign new_P1_R1207_U303 = ~new_P1_R1207_U301 | ~new_P1_R1207_U302;
  assign new_P1_R1207_U304 = ~new_P1_U3974 | ~new_P1_R1207_U85;
  assign new_P1_R1207_U305 = ~new_P1_U3974 | ~new_P1_R1207_U85;
  assign new_P1_R1207_U306 = ~new_P1_R1207_U305 | ~new_P1_R1207_U86;
  assign new_P1_R1207_U307 = ~new_P1_U3054 | ~new_P1_R1207_U84;
  assign new_P1_R1207_U308 = ~new_P1_R1207_U153 | ~new_P1_R1207_U307 | ~new_P1_R1207_U306;
  assign new_P1_R1207_U309 = ~new_P1_R1207_U295 | ~new_P1_R1207_U82;
  assign new_P1_R1207_U310 = ~new_P1_R1207_U129 | ~new_P1_R1207_U309;
  assign new_P1_R1207_U311 = ~new_P1_R1207_U87 | ~new_P1_R1207_U177;
  assign new_P1_R1207_U312 = ~new_P1_R1207_U128 | ~new_P1_R1207_U311;
  assign new_P1_R1207_U313 = ~new_P1_R1207_U82 | ~new_P1_R1207_U177;
  assign new_P1_R1207_U314 = ~new_P1_R1207_U283 | ~new_P1_R1207_U159;
  assign new_P1_R1207_U315 = ~new_P1_R1207_U88;
  assign new_P1_R1207_U316 = ~new_P1_U3061 | ~new_P1_R1207_U45;
  assign new_P1_R1207_U317 = ~new_P1_R1207_U315 | ~new_P1_R1207_U316;
  assign new_P1_R1207_U318 = ~new_P1_R1207_U132 | ~new_P1_R1207_U317;
  assign new_P1_R1207_U319 = ~new_P1_R1207_U88 | ~new_P1_R1207_U176;
  assign new_P1_R1207_U320 = ~new_P1_U3979 | ~new_P1_R1207_U72;
  assign new_P1_R1207_U321 = ~new_P1_R1207_U9 | ~new_P1_R1207_U320 | ~new_P1_R1207_U319;
  assign new_P1_R1207_U322 = ~new_P1_U3061 | ~new_P1_R1207_U45;
  assign new_P1_R1207_U323 = ~new_P1_R1207_U176 | ~new_P1_R1207_U322;
  assign new_P1_R1207_U324 = ~new_P1_R1207_U283 | ~new_P1_R1207_U75;
  assign new_P1_R1207_U325 = ~new_P1_R1207_U257 | ~new_P1_R1207_U167;
  assign new_P1_R1207_U326 = ~new_P1_R1207_U89;
  assign new_P1_R1207_U327 = ~new_P1_U3074 | ~new_P1_R1207_U46;
  assign new_P1_R1207_U328 = ~new_P1_R1207_U326 | ~new_P1_R1207_U327;
  assign new_P1_R1207_U329 = ~new_P1_R1207_U139 | ~new_P1_R1207_U328;
  assign new_P1_R1207_U330 = ~new_P1_R1207_U89 | ~new_P1_R1207_U175;
  assign new_P1_R1207_U331 = ~new_P1_U3500 | ~new_P1_R1207_U58;
  assign new_P1_R1207_U332 = ~new_P1_R1207_U138 | ~new_P1_R1207_U330;
  assign new_P1_R1207_U333 = ~new_P1_U3074 | ~new_P1_R1207_U46;
  assign new_P1_R1207_U334 = ~new_P1_R1207_U175 | ~new_P1_R1207_U333;
  assign new_P1_R1207_U335 = ~new_P1_R1207_U257 | ~new_P1_R1207_U61;
  assign new_P1_R1207_U336 = ~new_P1_R1207_U212 | ~new_P1_R1207_U145;
  assign new_P1_R1207_U337 = ~new_P1_R1207_U90;
  assign new_P1_R1207_U338 = ~new_P1_U3062 | ~new_P1_R1207_U47;
  assign new_P1_R1207_U339 = ~new_P1_R1207_U337 | ~new_P1_R1207_U338;
  assign new_P1_R1207_U340 = ~new_P1_R1207_U143 | ~new_P1_R1207_U339;
  assign new_P1_R1207_U341 = ~new_P1_R1207_U90 | ~new_P1_R1207_U174;
  assign new_P1_R1207_U342 = ~new_P1_U3485 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U343 = ~new_P1_R1207_U142 | ~new_P1_R1207_U341;
  assign new_P1_R1207_U344 = ~new_P1_U3062 | ~new_P1_R1207_U47;
  assign new_P1_R1207_U345 = ~new_P1_R1207_U174 | ~new_P1_R1207_U344;
  assign new_P1_R1207_U346 = ~new_P1_U3077 | ~new_P1_R1207_U22;
  assign new_P1_R1207_U347 = ~new_P1_R1207_U385 | ~new_P1_R1207_U304 | ~new_P1_R1207_U303;
  assign new_P1_R1207_U348 = ~new_P1_U3479 | ~new_P1_R1207_U40;
  assign new_P1_R1207_U349 = ~new_P1_U3083 | ~new_P1_R1207_U39;
  assign new_P1_R1207_U350 = ~new_P1_R1207_U213 | ~new_P1_R1207_U145;
  assign new_P1_R1207_U351 = ~new_P1_R1207_U211 | ~new_P1_R1207_U144;
  assign new_P1_R1207_U352 = ~new_P1_U3476 | ~new_P1_R1207_U38;
  assign new_P1_R1207_U353 = ~new_P1_U3084 | ~new_P1_R1207_U35;
  assign new_P1_R1207_U354 = ~new_P1_U3476 | ~new_P1_R1207_U38;
  assign new_P1_R1207_U355 = ~new_P1_U3084 | ~new_P1_R1207_U35;
  assign new_P1_R1207_U356 = ~new_P1_R1207_U355 | ~new_P1_R1207_U354;
  assign new_P1_R1207_U357 = ~new_P1_U3473 | ~new_P1_R1207_U36;
  assign new_P1_R1207_U358 = ~new_P1_U3070 | ~new_P1_R1207_U19;
  assign new_P1_R1207_U359 = ~new_P1_R1207_U218 | ~new_P1_R1207_U41;
  assign new_P1_R1207_U360 = ~new_P1_R1207_U146 | ~new_P1_R1207_U205;
  assign new_P1_R1207_U361 = ~new_P1_U3470 | ~new_P1_R1207_U31;
  assign new_P1_R1207_U362 = ~new_P1_U3071 | ~new_P1_R1207_U29;
  assign new_P1_R1207_U363 = ~new_P1_R1207_U362 | ~new_P1_R1207_U361;
  assign new_P1_R1207_U364 = ~new_P1_U3467 | ~new_P1_R1207_U32;
  assign new_P1_R1207_U365 = ~new_P1_U3067 | ~new_P1_R1207_U20;
  assign new_P1_R1207_U366 = ~new_P1_R1207_U228 | ~new_P1_R1207_U42;
  assign new_P1_R1207_U367 = ~new_P1_R1207_U147 | ~new_P1_R1207_U220;
  assign new_P1_R1207_U368 = ~new_P1_U3464 | ~new_P1_R1207_U33;
  assign new_P1_R1207_U369 = ~new_P1_U3060 | ~new_P1_R1207_U30;
  assign new_P1_R1207_U370 = ~new_P1_R1207_U229 | ~new_P1_R1207_U149;
  assign new_P1_R1207_U371 = ~new_P1_R1207_U195 | ~new_P1_R1207_U148;
  assign new_P1_R1207_U372 = ~new_P1_U3461 | ~new_P1_R1207_U28;
  assign new_P1_R1207_U373 = ~new_P1_U3064 | ~new_P1_R1207_U25;
  assign new_P1_R1207_U374 = ~new_P1_U3461 | ~new_P1_R1207_U28;
  assign new_P1_R1207_U375 = ~new_P1_U3064 | ~new_P1_R1207_U25;
  assign new_P1_R1207_U376 = ~new_P1_R1207_U375 | ~new_P1_R1207_U374;
  assign new_P1_R1207_U377 = ~new_P1_U3458 | ~new_P1_R1207_U26;
  assign new_P1_R1207_U378 = ~new_P1_U3068 | ~new_P1_R1207_U21;
  assign new_P1_R1207_U379 = ~new_P1_R1207_U234 | ~new_P1_R1207_U43;
  assign new_P1_R1207_U380 = ~new_P1_R1207_U150 | ~new_P1_R1207_U189;
  assign new_P1_R1207_U381 = ~new_P1_U3985 | ~new_P1_R1207_U152;
  assign new_P1_R1207_U382 = ~new_P1_U3055 | ~new_P1_R1207_U151;
  assign new_P1_R1207_U383 = ~new_P1_U3985 | ~new_P1_R1207_U152;
  assign new_P1_R1207_U384 = ~new_P1_U3055 | ~new_P1_R1207_U151;
  assign new_P1_R1207_U385 = ~new_P1_R1207_U384 | ~new_P1_R1207_U383;
  assign new_P1_R1207_U386 = ~new_P1_U3974 | ~new_P1_R1207_U85;
  assign new_P1_R1207_U387 = ~new_P1_U3054 | ~new_P1_R1207_U84;
  assign new_P1_R1207_U388 = ~new_P1_R1207_U127;
  assign new_P1_R1207_U389 = ~new_P1_R1207_U388 | ~new_P1_R1207_U301;
  assign new_P1_R1207_U390 = ~new_P1_R1207_U127 | ~new_P1_R1207_U86;
  assign new_P1_R1207_U391 = ~new_P1_U3975 | ~new_P1_R1207_U83;
  assign new_P1_R1207_U392 = ~new_P1_U3053 | ~new_P1_R1207_U80;
  assign new_P1_R1207_U393 = ~new_P1_U3975 | ~new_P1_R1207_U83;
  assign new_P1_R1207_U394 = ~new_P1_U3053 | ~new_P1_R1207_U80;
  assign new_P1_R1207_U395 = ~new_P1_R1207_U394 | ~new_P1_R1207_U393;
  assign new_P1_R1207_U396 = ~new_P1_U3976 | ~new_P1_R1207_U81;
  assign new_P1_R1207_U397 = ~new_P1_U3057 | ~new_P1_R1207_U44;
  assign new_P1_R1207_U398 = ~new_P1_R1207_U313 | ~new_P1_R1207_U87;
  assign new_P1_R1207_U399 = ~new_P1_R1207_U154 | ~new_P1_R1207_U295;
  assign new_P1_R1207_U400 = ~new_P1_U3977 | ~new_P1_R1207_U79;
  assign new_P1_R1207_U401 = ~new_P1_U3058 | ~new_P1_R1207_U78;
  assign new_P1_R1207_U402 = ~new_P1_R1207_U130;
  assign new_P1_R1207_U403 = ~new_P1_R1207_U291 | ~new_P1_R1207_U402;
  assign new_P1_R1207_U404 = ~new_P1_R1207_U130 | ~new_P1_R1207_U155;
  assign new_P1_R1207_U405 = ~new_P1_U3978 | ~new_P1_R1207_U77;
  assign new_P1_R1207_U406 = ~new_P1_U3065 | ~new_P1_R1207_U76;
  assign new_P1_R1207_U407 = ~new_P1_R1207_U131;
  assign new_P1_R1207_U408 = ~new_P1_R1207_U287 | ~new_P1_R1207_U407;
  assign new_P1_R1207_U409 = ~new_P1_R1207_U131 | ~new_P1_R1207_U156;
  assign new_P1_R1207_U410 = ~new_P1_U3979 | ~new_P1_R1207_U72;
  assign new_P1_R1207_U411 = ~new_P1_U3066 | ~new_P1_R1207_U70;
  assign new_P1_R1207_U412 = ~new_P1_R1207_U411 | ~new_P1_R1207_U410;
  assign new_P1_R1207_U413 = ~new_P1_U3980 | ~new_P1_R1207_U73;
  assign new_P1_R1207_U414 = ~new_P1_U3061 | ~new_P1_R1207_U45;
  assign new_P1_R1207_U415 = ~new_P1_R1207_U323 | ~new_P1_R1207_U88;
  assign new_P1_R1207_U416 = ~new_P1_R1207_U157 | ~new_P1_R1207_U315;
  assign new_P1_R1207_U417 = ~new_P1_U3981 | ~new_P1_R1207_U74;
  assign new_P1_R1207_U418 = ~new_P1_U3075 | ~new_P1_R1207_U71;
  assign new_P1_R1207_U419 = ~new_P1_R1207_U324 | ~new_P1_R1207_U159;
  assign new_P1_R1207_U420 = ~new_P1_R1207_U277 | ~new_P1_R1207_U158;
  assign new_P1_R1207_U421 = ~new_P1_U3982 | ~new_P1_R1207_U69;
  assign new_P1_R1207_U422 = ~new_P1_U3076 | ~new_P1_R1207_U68;
  assign new_P1_R1207_U423 = ~new_P1_R1207_U133;
  assign new_P1_R1207_U424 = ~new_P1_R1207_U273 | ~new_P1_R1207_U423;
  assign new_P1_R1207_U425 = ~new_P1_R1207_U133 | ~new_P1_R1207_U160;
  assign new_P1_R1207_U426 = ~new_P1_R1207_U185 | ~new_P1_R1207_U24;
  assign new_P1_R1207_U427 = ~new_P1_U3078 | ~new_P1_R1207_U23;
  assign new_P1_R1207_U428 = ~new_P1_R1207_U134;
  assign new_P1_R1207_U429 = ~new_P1_U3455 | ~new_P1_R1207_U428;
  assign new_P1_R1207_U430 = ~new_P1_R1207_U134 | ~new_P1_R1207_U161;
  assign new_P1_R1207_U431 = ~new_P1_U3508 | ~new_P1_R1207_U67;
  assign new_P1_R1207_U432 = ~new_P1_U3081 | ~new_P1_R1207_U66;
  assign new_P1_R1207_U433 = ~new_P1_R1207_U135;
  assign new_P1_R1207_U434 = ~new_P1_R1207_U269 | ~new_P1_R1207_U433;
  assign new_P1_R1207_U435 = ~new_P1_R1207_U135 | ~new_P1_R1207_U162;
  assign new_P1_R1207_U436 = ~new_P1_U3506 | ~new_P1_R1207_U65;
  assign new_P1_R1207_U437 = ~new_P1_U3082 | ~new_P1_R1207_U163;
  assign new_P1_R1207_U438 = ~new_P1_R1207_U136;
  assign new_P1_R1207_U439 = ~new_P1_R1207_U438 | ~new_P1_R1207_U265;
  assign new_P1_R1207_U440 = ~new_P1_R1207_U136 | ~new_P1_R1207_U64;
  assign new_P1_R1207_U441 = ~new_P1_U3503 | ~new_P1_R1207_U63;
  assign new_P1_R1207_U442 = ~new_P1_U3069 | ~new_P1_R1207_U62;
  assign new_P1_R1207_U443 = ~new_P1_R1207_U137;
  assign new_P1_R1207_U444 = ~new_P1_R1207_U261 | ~new_P1_R1207_U443;
  assign new_P1_R1207_U445 = ~new_P1_R1207_U137 | ~new_P1_R1207_U164;
  assign new_P1_R1207_U446 = ~new_P1_U3500 | ~new_P1_R1207_U58;
  assign new_P1_R1207_U447 = ~new_P1_U3073 | ~new_P1_R1207_U56;
  assign new_P1_R1207_U448 = ~new_P1_R1207_U447 | ~new_P1_R1207_U446;
  assign new_P1_R1207_U449 = ~new_P1_U3497 | ~new_P1_R1207_U59;
  assign new_P1_R1207_U450 = ~new_P1_U3074 | ~new_P1_R1207_U46;
  assign new_P1_R1207_U451 = ~new_P1_R1207_U334 | ~new_P1_R1207_U89;
  assign new_P1_R1207_U452 = ~new_P1_R1207_U165 | ~new_P1_R1207_U326;
  assign new_P1_R1207_U453 = ~new_P1_U3494 | ~new_P1_R1207_U60;
  assign new_P1_R1207_U454 = ~new_P1_U3079 | ~new_P1_R1207_U57;
  assign new_P1_R1207_U455 = ~new_P1_R1207_U335 | ~new_P1_R1207_U167;
  assign new_P1_R1207_U456 = ~new_P1_R1207_U251 | ~new_P1_R1207_U166;
  assign new_P1_R1207_U457 = ~new_P1_U3491 | ~new_P1_R1207_U55;
  assign new_P1_R1207_U458 = ~new_P1_U3080 | ~new_P1_R1207_U54;
  assign new_P1_R1207_U459 = ~new_P1_R1207_U140;
  assign new_P1_R1207_U460 = ~new_P1_R1207_U247 | ~new_P1_R1207_U459;
  assign new_P1_R1207_U461 = ~new_P1_R1207_U140 | ~new_P1_R1207_U168;
  assign new_P1_R1207_U462 = ~new_P1_U3488 | ~new_P1_R1207_U53;
  assign new_P1_R1207_U463 = ~new_P1_U3072 | ~new_P1_R1207_U52;
  assign new_P1_R1207_U464 = ~new_P1_R1207_U141;
  assign new_P1_R1207_U465 = ~new_P1_R1207_U243 | ~new_P1_R1207_U464;
  assign new_P1_R1207_U466 = ~new_P1_R1207_U141 | ~new_P1_R1207_U169;
  assign new_P1_R1207_U467 = ~new_P1_U3485 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U468 = ~new_P1_U3063 | ~new_P1_R1207_U48;
  assign new_P1_R1207_U469 = ~new_P1_R1207_U468 | ~new_P1_R1207_U467;
  assign new_P1_R1207_U470 = ~new_P1_U3482 | ~new_P1_R1207_U50;
  assign new_P1_R1207_U471 = ~new_P1_U3062 | ~new_P1_R1207_U47;
  assign new_P1_R1207_U472 = ~new_P1_R1207_U345 | ~new_P1_R1207_U90;
  assign new_P1_R1207_U473 = ~new_P1_R1207_U170 | ~new_P1_R1207_U337;
  assign new_P1_R1165_U4 = new_P1_R1165_U210 & new_P1_R1165_U209;
  assign new_P1_R1165_U5 = new_P1_R1165_U222 & new_P1_R1165_U221;
  assign new_P1_R1165_U6 = new_P1_R1165_U253 & new_P1_R1165_U252;
  assign new_P1_R1165_U7 = new_P1_R1165_U271 & new_P1_R1165_U270;
  assign new_P1_R1165_U8 = new_P1_R1165_U283 & new_P1_R1165_U282;
  assign new_P1_R1165_U9 = new_P1_R1165_U507 & new_P1_R1165_U506;
  assign new_P1_R1165_U10 = new_P1_R1165_U339 & new_P1_R1165_U336;
  assign new_P1_R1165_U11 = new_P1_R1165_U330 & new_P1_R1165_U327;
  assign new_P1_R1165_U12 = new_P1_R1165_U323 & new_P1_R1165_U320;
  assign new_P1_R1165_U13 = new_P1_R1165_U314 & new_P1_R1165_U360 & new_P1_R1165_U311;
  assign new_P1_R1165_U14 = new_P1_R1165_U245 & new_P1_R1165_U242;
  assign new_P1_R1165_U15 = new_P1_R1165_U238 & new_P1_R1165_U235;
  assign new_P1_R1165_U16 = ~new_P1_U3211;
  assign new_P1_R1165_U17 = ~new_P1_U3175;
  assign new_P1_R1165_U18 = ~new_P1_U3175 | ~new_P1_R1165_U58;
  assign new_P1_R1165_U19 = ~new_P1_U3174;
  assign new_P1_R1165_U20 = ~new_P1_U3177;
  assign new_P1_R1165_U21 = ~new_P1_U3179;
  assign new_P1_R1165_U22 = ~new_P1_U3179 | ~new_P1_R1165_U61;
  assign new_P1_R1165_U23 = ~new_P1_U3178;
  assign new_P1_R1165_U24 = ~new_P1_U3181;
  assign new_P1_R1165_U25 = ~new_P1_U3180;
  assign new_P1_R1165_U26 = ~new_P1_U3176;
  assign new_P1_R1165_U27 = ~new_P1_U3173;
  assign new_P1_R1165_U28 = ~new_P1_U3172;
  assign new_P1_R1165_U29 = ~new_P1_R1165_U219 | ~new_P1_R1165_U218;
  assign new_P1_R1165_U30 = ~new_P1_R1165_U207 | ~new_P1_R1165_U206;
  assign new_P1_R1165_U31 = ~new_P1_U3154;
  assign new_P1_R1165_U32 = ~new_P1_U3155;
  assign new_P1_R1165_U33 = ~new_P1_U3156;
  assign new_P1_R1165_U34 = ~new_P1_U3157;
  assign new_P1_R1165_U35 = ~new_P1_U3165;
  assign new_P1_R1165_U36 = ~new_P1_U3165 | ~new_P1_R1165_U71;
  assign new_P1_R1165_U37 = ~new_P1_U3164;
  assign new_P1_R1165_U38 = ~new_P1_U3171;
  assign new_P1_R1165_U39 = ~new_P1_U3169;
  assign new_P1_R1165_U40 = ~new_P1_U3170;
  assign new_P1_R1165_U41 = ~new_P1_U3170 | ~new_P1_R1165_U74;
  assign new_P1_R1165_U42 = ~new_P1_U3168;
  assign new_P1_R1165_U43 = ~new_P1_U3167;
  assign new_P1_R1165_U44 = ~new_P1_U3166;
  assign new_P1_R1165_U45 = ~new_P1_U3163;
  assign new_P1_R1165_U46 = ~new_P1_U3161;
  assign new_P1_R1165_U47 = ~new_P1_U3162;
  assign new_P1_R1165_U48 = ~new_P1_U3162 | ~new_P1_R1165_U80;
  assign new_P1_R1165_U49 = ~new_P1_U3160;
  assign new_P1_R1165_U50 = ~new_P1_U3159;
  assign new_P1_R1165_U51 = ~new_P1_U3158;
  assign new_P1_R1165_U52 = ~new_P1_U3155 | ~new_P1_R1165_U69;
  assign new_P1_R1165_U53 = ~new_P1_R1165_U200 | ~new_P1_R1165_U309;
  assign new_P1_R1165_U54 = ~new_P1_R1165_U48 | ~new_P1_R1165_U316;
  assign new_P1_R1165_U55 = ~new_P1_R1165_U268 | ~new_P1_R1165_U267;
  assign new_P1_R1165_U56 = ~new_P1_R1165_U41 | ~new_P1_R1165_U332;
  assign new_P1_R1165_U57 = ~new_P1_R1165_U366 | ~new_P1_R1165_U365;
  assign new_P1_R1165_U58 = ~new_P1_R1165_U395 | ~new_P1_R1165_U394;
  assign new_P1_R1165_U59 = ~new_P1_R1165_U392 | ~new_P1_R1165_U391;
  assign new_P1_R1165_U60 = ~new_P1_R1165_U374 | ~new_P1_R1165_U373;
  assign new_P1_R1165_U61 = ~new_P1_R1165_U386 | ~new_P1_R1165_U385;
  assign new_P1_R1165_U62 = ~new_P1_R1165_U383 | ~new_P1_R1165_U382;
  assign new_P1_R1165_U63 = ~new_P1_R1165_U377 | ~new_P1_R1165_U376;
  assign new_P1_R1165_U64 = ~new_P1_R1165_U380 | ~new_P1_R1165_U379;
  assign new_P1_R1165_U65 = ~new_P1_R1165_U389 | ~new_P1_R1165_U388;
  assign new_P1_R1165_U66 = ~new_P1_R1165_U398 | ~new_P1_R1165_U397;
  assign new_P1_R1165_U67 = ~new_P1_R1165_U438 | ~new_P1_R1165_U437;
  assign new_P1_R1165_U68 = ~new_P1_R1165_U441 | ~new_P1_R1165_U440;
  assign new_P1_R1165_U69 = ~new_P1_R1165_U444 | ~new_P1_R1165_U443;
  assign new_P1_R1165_U70 = ~new_P1_R1165_U447 | ~new_P1_R1165_U446;
  assign new_P1_R1165_U71 = ~new_P1_R1165_U471 | ~new_P1_R1165_U470;
  assign new_P1_R1165_U72 = ~new_P1_R1165_U468 | ~new_P1_R1165_U467;
  assign new_P1_R1165_U73 = ~new_P1_R1165_U450 | ~new_P1_R1165_U449;
  assign new_P1_R1165_U74 = ~new_P1_R1165_U459 | ~new_P1_R1165_U458;
  assign new_P1_R1165_U75 = ~new_P1_R1165_U453 | ~new_P1_R1165_U452;
  assign new_P1_R1165_U76 = ~new_P1_R1165_U456 | ~new_P1_R1165_U455;
  assign new_P1_R1165_U77 = ~new_P1_R1165_U462 | ~new_P1_R1165_U461;
  assign new_P1_R1165_U78 = ~new_P1_R1165_U465 | ~new_P1_R1165_U464;
  assign new_P1_R1165_U79 = ~new_P1_R1165_U474 | ~new_P1_R1165_U473;
  assign new_P1_R1165_U80 = ~new_P1_R1165_U483 | ~new_P1_R1165_U482;
  assign new_P1_R1165_U81 = ~new_P1_R1165_U477 | ~new_P1_R1165_U476;
  assign new_P1_R1165_U82 = ~new_P1_R1165_U480 | ~new_P1_R1165_U479;
  assign new_P1_R1165_U83 = ~new_P1_R1165_U486 | ~new_P1_R1165_U485;
  assign new_P1_R1165_U84 = ~new_P1_R1165_U489 | ~new_P1_R1165_U488;
  assign new_P1_R1165_U85 = ~new_P1_R1165_U495 | ~new_P1_R1165_U494;
  assign new_P1_R1165_U86 = ~new_P1_R1165_U602 | ~new_P1_R1165_U601;
  assign new_P1_R1165_U87 = ~new_P1_R1165_U401 | ~new_P1_R1165_U400;
  assign new_P1_R1165_U88 = ~new_P1_R1165_U408 | ~new_P1_R1165_U407;
  assign new_P1_R1165_U89 = ~new_P1_R1165_U415 | ~new_P1_R1165_U414;
  assign new_P1_R1165_U90 = ~new_P1_R1165_U422 | ~new_P1_R1165_U421;
  assign new_P1_R1165_U91 = ~new_P1_R1165_U429 | ~new_P1_R1165_U428;
  assign new_P1_R1165_U92 = ~new_P1_R1165_U436 | ~new_P1_R1165_U435;
  assign new_P1_R1165_U93 = ~new_P1_R1165_U498 | ~new_P1_R1165_U497;
  assign new_P1_R1165_U94 = ~new_P1_R1165_U505 | ~new_P1_R1165_U504;
  assign new_P1_R1165_U95 = ~new_P1_R1165_U512 | ~new_P1_R1165_U511;
  assign new_P1_R1165_U96 = ~new_P1_R1165_U517 | ~new_P1_R1165_U516;
  assign new_P1_R1165_U97 = ~new_P1_R1165_U524 | ~new_P1_R1165_U523;
  assign new_P1_R1165_U98 = ~new_P1_R1165_U531 | ~new_P1_R1165_U530;
  assign new_P1_R1165_U99 = ~new_P1_R1165_U538 | ~new_P1_R1165_U537;
  assign new_P1_R1165_U100 = ~new_P1_R1165_U545 | ~new_P1_R1165_U544;
  assign new_P1_R1165_U101 = ~new_P1_R1165_U550 | ~new_P1_R1165_U549;
  assign new_P1_R1165_U102 = ~new_P1_R1165_U557 | ~new_P1_R1165_U556;
  assign new_P1_R1165_U103 = ~new_P1_R1165_U564 | ~new_P1_R1165_U563;
  assign new_P1_R1165_U104 = ~new_P1_R1165_U571 | ~new_P1_R1165_U570;
  assign new_P1_R1165_U105 = ~new_P1_R1165_U578 | ~new_P1_R1165_U577;
  assign new_P1_R1165_U106 = ~new_P1_R1165_U585 | ~new_P1_R1165_U584;
  assign new_P1_R1165_U107 = ~new_P1_R1165_U590 | ~new_P1_R1165_U589;
  assign new_P1_R1165_U108 = ~new_P1_R1165_U597 | ~new_P1_R1165_U596;
  assign new_P1_R1165_U109 = new_P1_R1165_U213 & new_P1_R1165_U212;
  assign new_P1_R1165_U110 = new_P1_R1165_U226 & new_P1_R1165_U225;
  assign new_P1_R1165_U111 = new_P1_R1165_U18 & new_P1_R1165_U410 & new_P1_R1165_U409;
  assign new_P1_R1165_U112 = new_P1_R1165_U237 & new_P1_R1165_U5;
  assign new_P1_R1165_U113 = new_P1_R1165_U22 & new_P1_R1165_U431 & new_P1_R1165_U430;
  assign new_P1_R1165_U114 = new_P1_R1165_U244 & new_P1_R1165_U4;
  assign new_P1_R1165_U115 = new_P1_R1165_U257 & new_P1_R1165_U6;
  assign new_P1_R1165_U116 = new_P1_R1165_U255 & new_P1_R1165_U195;
  assign new_P1_R1165_U117 = new_P1_R1165_U275 & new_P1_R1165_U274;
  assign new_P1_R1165_U118 = new_P1_R1165_U287 & new_P1_R1165_U8;
  assign new_P1_R1165_U119 = new_P1_R1165_U285 & new_P1_R1165_U196;
  assign new_P1_R1165_U120 = new_P1_R1165_U359 & new_P1_R1165_U52;
  assign new_P1_R1165_U121 = new_P1_R1165_U308 & new_P1_R1165_U303;
  assign new_P1_R1165_U122 = new_P1_R1165_U356 & new_P1_R1165_U307;
  assign new_P1_R1165_U123 = ~new_P1_R1165_U492 | ~new_P1_R1165_U491;
  assign new_P1_R1165_U124 = new_P1_R1165_U352 & new_P1_R1165_U52;
  assign new_P1_R1165_U125 = new_P1_R1165_U442 & new_P1_R1165_U33;
  assign new_P1_R1165_U126 = new_P1_R1165_U200 & new_P1_R1165_U197;
  assign new_P1_R1165_U127 = new_P1_R1165_U313 & new_P1_R1165_U193;
  assign new_P1_R1165_U128 = new_P1_R1165_U9 & new_P1_R1165_U197;
  assign new_P1_R1165_U129 = new_P1_R1165_U196 & new_P1_R1165_U533 & new_P1_R1165_U532;
  assign new_P1_R1165_U130 = new_P1_R1165_U322 & new_P1_R1165_U8;
  assign new_P1_R1165_U131 = new_P1_R1165_U36 & new_P1_R1165_U559 & new_P1_R1165_U558;
  assign new_P1_R1165_U132 = new_P1_R1165_U329 & new_P1_R1165_U7;
  assign new_P1_R1165_U133 = new_P1_R1165_U195 & new_P1_R1165_U580 & new_P1_R1165_U579;
  assign new_P1_R1165_U134 = new_P1_R1165_U338 & new_P1_R1165_U6;
  assign new_P1_R1165_U135 = ~new_P1_R1165_U599 | ~new_P1_R1165_U598;
  assign new_P1_R1165_U136 = ~new_P1_U3201;
  assign new_P1_R1165_U137 = new_P1_R1165_U369 & new_P1_R1165_U368;
  assign new_P1_R1165_U138 = ~new_P1_U3206;
  assign new_P1_R1165_U139 = ~new_P1_U3210;
  assign new_P1_R1165_U140 = ~new_P1_U3209;
  assign new_P1_R1165_U141 = ~new_P1_U3207;
  assign new_P1_R1165_U142 = ~new_P1_U3208;
  assign new_P1_R1165_U143 = ~new_P1_U3205;
  assign new_P1_R1165_U144 = ~new_P1_U3203;
  assign new_P1_R1165_U145 = ~new_P1_U3204;
  assign new_P1_R1165_U146 = ~new_P1_U3202;
  assign new_P1_R1165_U147 = ~new_P1_R1165_U231 | ~new_P1_R1165_U230;
  assign new_P1_R1165_U148 = new_P1_R1165_U403 & new_P1_R1165_U402;
  assign new_P1_R1165_U149 = ~new_P1_R1165_U110 | ~new_P1_R1165_U227;
  assign new_P1_R1165_U150 = new_P1_R1165_U417 & new_P1_R1165_U416;
  assign new_P1_R1165_U151 = ~new_P1_R1165_U361 | ~new_P1_R1165_U350;
  assign new_P1_R1165_U152 = new_P1_R1165_U424 & new_P1_R1165_U423;
  assign new_P1_R1165_U153 = ~new_P1_R1165_U109 | ~new_P1_R1165_U214;
  assign new_P1_R1165_U154 = ~new_P1_U3183;
  assign new_P1_R1165_U155 = ~new_P1_U3185;
  assign new_P1_R1165_U156 = ~new_P1_U3184;
  assign new_P1_R1165_U157 = ~new_P1_U3186;
  assign new_P1_R1165_U158 = ~new_P1_U3200;
  assign new_P1_R1165_U159 = ~new_P1_U3197;
  assign new_P1_R1165_U160 = ~new_P1_U3198;
  assign new_P1_R1165_U161 = ~new_P1_U3199;
  assign new_P1_R1165_U162 = ~new_P1_U3196;
  assign new_P1_R1165_U163 = ~new_P1_U3195;
  assign new_P1_R1165_U164 = ~new_P1_U3193;
  assign new_P1_R1165_U165 = ~new_P1_U3194;
  assign new_P1_R1165_U166 = ~new_P1_U3192;
  assign new_P1_R1165_U167 = ~new_P1_U3189;
  assign new_P1_R1165_U168 = ~new_P1_U3190;
  assign new_P1_R1165_U169 = ~new_P1_U3191;
  assign new_P1_R1165_U170 = ~new_P1_U3188;
  assign new_P1_R1165_U171 = ~new_P1_U3187;
  assign new_P1_R1165_U172 = ~new_P1_U3153;
  assign new_P1_R1165_U173 = ~new_P1_U3182;
  assign new_P1_R1165_U174 = new_P1_R1165_U500 & new_P1_R1165_U499;
  assign new_P1_R1165_U175 = ~new_P1_R1165_U124 | ~new_P1_R1165_U304;
  assign new_P1_R1165_U176 = ~new_P1_R1165_U298 | ~new_P1_R1165_U297;
  assign new_P1_R1165_U177 = new_P1_R1165_U519 & new_P1_R1165_U518;
  assign new_P1_R1165_U178 = ~new_P1_R1165_U294 | ~new_P1_R1165_U293;
  assign new_P1_R1165_U179 = new_P1_R1165_U526 & new_P1_R1165_U525;
  assign new_P1_R1165_U180 = ~new_P1_R1165_U290 | ~new_P1_R1165_U289;
  assign new_P1_R1165_U181 = new_P1_R1165_U540 & new_P1_R1165_U539;
  assign new_P1_R1165_U182 = ~new_P1_R1165_U203 | ~new_P1_R1165_U202;
  assign new_P1_R1165_U183 = ~new_P1_R1165_U280 | ~new_P1_R1165_U279;
  assign new_P1_R1165_U184 = new_P1_R1165_U552 & new_P1_R1165_U551;
  assign new_P1_R1165_U185 = ~new_P1_R1165_U117 | ~new_P1_R1165_U276;
  assign new_P1_R1165_U186 = new_P1_R1165_U566 & new_P1_R1165_U565;
  assign new_P1_R1165_U187 = ~new_P1_R1165_U264 | ~new_P1_R1165_U263;
  assign new_P1_R1165_U188 = new_P1_R1165_U573 & new_P1_R1165_U572;
  assign new_P1_R1165_U189 = ~new_P1_R1165_U260 | ~new_P1_R1165_U259;
  assign new_P1_R1165_U190 = ~new_P1_R1165_U250 | ~new_P1_R1165_U249;
  assign new_P1_R1165_U191 = new_P1_R1165_U592 & new_P1_R1165_U591;
  assign new_P1_R1165_U192 = ~new_P1_R1165_U363 | ~new_P1_R1165_U353;
  assign new_P1_R1165_U193 = ~new_P1_R1165_U355 | ~new_P1_R1165_U354;
  assign new_P1_R1165_U194 = ~new_P1_R1165_U22;
  assign new_P1_R1165_U195 = ~new_P1_U3169 | ~new_P1_R1165_U76;
  assign new_P1_R1165_U196 = ~new_P1_U3161 | ~new_P1_R1165_U82;
  assign new_P1_R1165_U197 = ~new_P1_U3156 | ~new_P1_R1165_U68;
  assign new_P1_R1165_U198 = ~new_P1_R1165_U41;
  assign new_P1_R1165_U199 = ~new_P1_R1165_U48;
  assign new_P1_R1165_U200 = ~new_P1_U3157 | ~new_P1_R1165_U70;
  assign new_P1_R1165_U201 = new_P1_U3211 | new_P1_U3181;
  assign new_P1_R1165_U202 = ~new_P1_R1165_U63 | ~new_P1_R1165_U201;
  assign new_P1_R1165_U203 = ~new_P1_U3181 | ~new_P1_U3211;
  assign new_P1_R1165_U204 = ~new_P1_R1165_U182;
  assign new_P1_R1165_U205 = ~new_P1_R1165_U381 | ~new_P1_R1165_U25;
  assign new_P1_R1165_U206 = ~new_P1_R1165_U205 | ~new_P1_R1165_U182;
  assign new_P1_R1165_U207 = ~new_P1_U3180 | ~new_P1_R1165_U64;
  assign new_P1_R1165_U208 = ~new_P1_R1165_U30;
  assign new_P1_R1165_U209 = ~new_P1_R1165_U384 | ~new_P1_R1165_U23;
  assign new_P1_R1165_U210 = ~new_P1_R1165_U387 | ~new_P1_R1165_U21;
  assign new_P1_R1165_U211 = ~new_P1_R1165_U23 | ~new_P1_R1165_U22;
  assign new_P1_R1165_U212 = ~new_P1_R1165_U62 | ~new_P1_R1165_U211;
  assign new_P1_R1165_U213 = ~new_P1_U3178 | ~new_P1_R1165_U194;
  assign new_P1_R1165_U214 = ~new_P1_R1165_U4 | ~new_P1_R1165_U30;
  assign new_P1_R1165_U215 = ~new_P1_R1165_U153;
  assign new_P1_R1165_U216 = ~new_P1_R1165_U375 | ~new_P1_R1165_U20;
  assign new_P1_R1165_U217 = ~new_P1_R1165_U390 | ~new_P1_R1165_U26;
  assign new_P1_R1165_U218 = ~new_P1_R1165_U217 | ~new_P1_R1165_U151;
  assign new_P1_R1165_U219 = ~new_P1_U3176 | ~new_P1_R1165_U65;
  assign new_P1_R1165_U220 = ~new_P1_R1165_U29;
  assign new_P1_R1165_U221 = ~new_P1_R1165_U393 | ~new_P1_R1165_U19;
  assign new_P1_R1165_U222 = ~new_P1_R1165_U396 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U223 = ~new_P1_R1165_U18;
  assign new_P1_R1165_U224 = ~new_P1_R1165_U19 | ~new_P1_R1165_U18;
  assign new_P1_R1165_U225 = ~new_P1_R1165_U59 | ~new_P1_R1165_U224;
  assign new_P1_R1165_U226 = ~new_P1_U3174 | ~new_P1_R1165_U223;
  assign new_P1_R1165_U227 = ~new_P1_R1165_U5 | ~new_P1_R1165_U29;
  assign new_P1_R1165_U228 = ~new_P1_R1165_U149;
  assign new_P1_R1165_U229 = ~new_P1_R1165_U399 | ~new_P1_R1165_U27;
  assign new_P1_R1165_U230 = ~new_P1_R1165_U229 | ~new_P1_R1165_U149;
  assign new_P1_R1165_U231 = ~new_P1_U3173 | ~new_P1_R1165_U66;
  assign new_P1_R1165_U232 = ~new_P1_R1165_U147;
  assign new_P1_R1165_U233 = ~new_P1_R1165_U396 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U234 = ~new_P1_R1165_U233 | ~new_P1_R1165_U29;
  assign new_P1_R1165_U235 = ~new_P1_R1165_U111 | ~new_P1_R1165_U234;
  assign new_P1_R1165_U236 = ~new_P1_R1165_U220 | ~new_P1_R1165_U18;
  assign new_P1_R1165_U237 = ~new_P1_U3174 | ~new_P1_R1165_U59;
  assign new_P1_R1165_U238 = ~new_P1_R1165_U112 | ~new_P1_R1165_U236;
  assign new_P1_R1165_U239 = ~new_P1_R1165_U396 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U240 = ~new_P1_R1165_U387 | ~new_P1_R1165_U21;
  assign new_P1_R1165_U241 = ~new_P1_R1165_U240 | ~new_P1_R1165_U30;
  assign new_P1_R1165_U242 = ~new_P1_R1165_U113 | ~new_P1_R1165_U241;
  assign new_P1_R1165_U243 = ~new_P1_R1165_U208 | ~new_P1_R1165_U22;
  assign new_P1_R1165_U244 = ~new_P1_U3178 | ~new_P1_R1165_U62;
  assign new_P1_R1165_U245 = ~new_P1_R1165_U114 | ~new_P1_R1165_U243;
  assign new_P1_R1165_U246 = ~new_P1_R1165_U387 | ~new_P1_R1165_U21;
  assign new_P1_R1165_U247 = ~new_P1_R1165_U367 | ~new_P1_R1165_U28;
  assign new_P1_R1165_U248 = ~new_P1_R1165_U451 | ~new_P1_R1165_U38;
  assign new_P1_R1165_U249 = ~new_P1_R1165_U248 | ~new_P1_R1165_U192;
  assign new_P1_R1165_U250 = ~new_P1_U3171 | ~new_P1_R1165_U73;
  assign new_P1_R1165_U251 = ~new_P1_R1165_U190;
  assign new_P1_R1165_U252 = ~new_P1_R1165_U454 | ~new_P1_R1165_U42;
  assign new_P1_R1165_U253 = ~new_P1_R1165_U457 | ~new_P1_R1165_U39;
  assign new_P1_R1165_U254 = ~new_P1_R1165_U198 | ~new_P1_R1165_U6;
  assign new_P1_R1165_U255 = ~new_P1_U3168 | ~new_P1_R1165_U75;
  assign new_P1_R1165_U256 = ~new_P1_R1165_U116 | ~new_P1_R1165_U254;
  assign new_P1_R1165_U257 = ~new_P1_R1165_U460 | ~new_P1_R1165_U40;
  assign new_P1_R1165_U258 = ~new_P1_R1165_U454 | ~new_P1_R1165_U42;
  assign new_P1_R1165_U259 = ~new_P1_R1165_U115 | ~new_P1_R1165_U190;
  assign new_P1_R1165_U260 = ~new_P1_R1165_U258 | ~new_P1_R1165_U256;
  assign new_P1_R1165_U261 = ~new_P1_R1165_U189;
  assign new_P1_R1165_U262 = ~new_P1_R1165_U463 | ~new_P1_R1165_U43;
  assign new_P1_R1165_U263 = ~new_P1_R1165_U262 | ~new_P1_R1165_U189;
  assign new_P1_R1165_U264 = ~new_P1_U3167 | ~new_P1_R1165_U77;
  assign new_P1_R1165_U265 = ~new_P1_R1165_U187;
  assign new_P1_R1165_U266 = ~new_P1_R1165_U466 | ~new_P1_R1165_U44;
  assign new_P1_R1165_U267 = ~new_P1_R1165_U266 | ~new_P1_R1165_U187;
  assign new_P1_R1165_U268 = ~new_P1_U3166 | ~new_P1_R1165_U78;
  assign new_P1_R1165_U269 = ~new_P1_R1165_U55;
  assign new_P1_R1165_U270 = ~new_P1_R1165_U469 | ~new_P1_R1165_U37;
  assign new_P1_R1165_U271 = ~new_P1_R1165_U472 | ~new_P1_R1165_U35;
  assign new_P1_R1165_U272 = ~new_P1_R1165_U36;
  assign new_P1_R1165_U273 = ~new_P1_R1165_U37 | ~new_P1_R1165_U36;
  assign new_P1_R1165_U274 = ~new_P1_R1165_U72 | ~new_P1_R1165_U273;
  assign new_P1_R1165_U275 = ~new_P1_U3164 | ~new_P1_R1165_U272;
  assign new_P1_R1165_U276 = ~new_P1_R1165_U7 | ~new_P1_R1165_U55;
  assign new_P1_R1165_U277 = ~new_P1_R1165_U185;
  assign new_P1_R1165_U278 = ~new_P1_R1165_U475 | ~new_P1_R1165_U45;
  assign new_P1_R1165_U279 = ~new_P1_R1165_U278 | ~new_P1_R1165_U185;
  assign new_P1_R1165_U280 = ~new_P1_U3163 | ~new_P1_R1165_U79;
  assign new_P1_R1165_U281 = ~new_P1_R1165_U183;
  assign new_P1_R1165_U282 = ~new_P1_R1165_U478 | ~new_P1_R1165_U49;
  assign new_P1_R1165_U283 = ~new_P1_R1165_U481 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U284 = ~new_P1_R1165_U199 | ~new_P1_R1165_U8;
  assign new_P1_R1165_U285 = ~new_P1_U3160 | ~new_P1_R1165_U81;
  assign new_P1_R1165_U286 = ~new_P1_R1165_U119 | ~new_P1_R1165_U284;
  assign new_P1_R1165_U287 = ~new_P1_R1165_U484 | ~new_P1_R1165_U47;
  assign new_P1_R1165_U288 = ~new_P1_R1165_U478 | ~new_P1_R1165_U49;
  assign new_P1_R1165_U289 = ~new_P1_R1165_U118 | ~new_P1_R1165_U183;
  assign new_P1_R1165_U290 = ~new_P1_R1165_U288 | ~new_P1_R1165_U286;
  assign new_P1_R1165_U291 = ~new_P1_R1165_U180;
  assign new_P1_R1165_U292 = ~new_P1_R1165_U487 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U293 = ~new_P1_R1165_U292 | ~new_P1_R1165_U180;
  assign new_P1_R1165_U294 = ~new_P1_U3159 | ~new_P1_R1165_U83;
  assign new_P1_R1165_U295 = ~new_P1_R1165_U178;
  assign new_P1_R1165_U296 = ~new_P1_R1165_U490 | ~new_P1_R1165_U51;
  assign new_P1_R1165_U297 = ~new_P1_R1165_U296 | ~new_P1_R1165_U178;
  assign new_P1_R1165_U298 = ~new_P1_U3158 | ~new_P1_R1165_U84;
  assign new_P1_R1165_U299 = ~new_P1_R1165_U176;
  assign new_P1_R1165_U300 = ~new_P1_R1165_U442 | ~new_P1_R1165_U33;
  assign new_P1_R1165_U301 = ~new_P1_R1165_U200 | ~new_P1_R1165_U197;
  assign new_P1_R1165_U302 = ~new_P1_R1165_U52;
  assign new_P1_R1165_U303 = ~new_P1_R1165_U448 | ~new_P1_R1165_U34;
  assign new_P1_R1165_U304 = ~new_P1_R1165_U193 | ~new_P1_R1165_U176 | ~new_P1_R1165_U303;
  assign new_P1_R1165_U305 = ~new_P1_R1165_U175;
  assign new_P1_R1165_U306 = ~new_P1_R1165_U439 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U307 = ~new_P1_U3154 | ~new_P1_R1165_U67;
  assign new_P1_R1165_U308 = ~new_P1_R1165_U439 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U309 = ~new_P1_R1165_U303 | ~new_P1_R1165_U176;
  assign new_P1_R1165_U310 = ~new_P1_R1165_U53;
  assign new_P1_R1165_U311 = ~new_P1_R1165_U125 | ~new_P1_R1165_U9;
  assign new_P1_R1165_U312 = ~new_P1_R1165_U126 | ~new_P1_R1165_U309;
  assign new_P1_R1165_U313 = ~new_P1_U3155 | ~new_P1_R1165_U69;
  assign new_P1_R1165_U314 = ~new_P1_R1165_U127 | ~new_P1_R1165_U312;
  assign new_P1_R1165_U315 = ~new_P1_R1165_U442 | ~new_P1_R1165_U33;
  assign new_P1_R1165_U316 = ~new_P1_R1165_U287 | ~new_P1_R1165_U183;
  assign new_P1_R1165_U317 = ~new_P1_R1165_U54;
  assign new_P1_R1165_U318 = ~new_P1_R1165_U481 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U319 = ~new_P1_R1165_U318 | ~new_P1_R1165_U54;
  assign new_P1_R1165_U320 = ~new_P1_R1165_U129 | ~new_P1_R1165_U319;
  assign new_P1_R1165_U321 = ~new_P1_R1165_U317 | ~new_P1_R1165_U196;
  assign new_P1_R1165_U322 = ~new_P1_U3160 | ~new_P1_R1165_U81;
  assign new_P1_R1165_U323 = ~new_P1_R1165_U130 | ~new_P1_R1165_U321;
  assign new_P1_R1165_U324 = ~new_P1_R1165_U481 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U325 = ~new_P1_R1165_U472 | ~new_P1_R1165_U35;
  assign new_P1_R1165_U326 = ~new_P1_R1165_U325 | ~new_P1_R1165_U55;
  assign new_P1_R1165_U327 = ~new_P1_R1165_U131 | ~new_P1_R1165_U326;
  assign new_P1_R1165_U328 = ~new_P1_R1165_U269 | ~new_P1_R1165_U36;
  assign new_P1_R1165_U329 = ~new_P1_U3164 | ~new_P1_R1165_U72;
  assign new_P1_R1165_U330 = ~new_P1_R1165_U132 | ~new_P1_R1165_U328;
  assign new_P1_R1165_U331 = ~new_P1_R1165_U472 | ~new_P1_R1165_U35;
  assign new_P1_R1165_U332 = ~new_P1_R1165_U257 | ~new_P1_R1165_U190;
  assign new_P1_R1165_U333 = ~new_P1_R1165_U56;
  assign new_P1_R1165_U334 = ~new_P1_R1165_U457 | ~new_P1_R1165_U39;
  assign new_P1_R1165_U335 = ~new_P1_R1165_U334 | ~new_P1_R1165_U56;
  assign new_P1_R1165_U336 = ~new_P1_R1165_U133 | ~new_P1_R1165_U335;
  assign new_P1_R1165_U337 = ~new_P1_R1165_U333 | ~new_P1_R1165_U195;
  assign new_P1_R1165_U338 = ~new_P1_U3168 | ~new_P1_R1165_U75;
  assign new_P1_R1165_U339 = ~new_P1_R1165_U134 | ~new_P1_R1165_U337;
  assign new_P1_R1165_U340 = ~new_P1_R1165_U457 | ~new_P1_R1165_U39;
  assign new_P1_R1165_U341 = ~new_P1_R1165_U239 | ~new_P1_R1165_U18;
  assign new_P1_R1165_U342 = ~new_P1_R1165_U246 | ~new_P1_R1165_U22;
  assign new_P1_R1165_U343 = ~new_P1_R1165_U315 | ~new_P1_R1165_U197;
  assign new_P1_R1165_U344 = ~new_P1_R1165_U303 | ~new_P1_R1165_U200;
  assign new_P1_R1165_U345 = ~new_P1_R1165_U324 | ~new_P1_R1165_U196;
  assign new_P1_R1165_U346 = ~new_P1_R1165_U287 | ~new_P1_R1165_U48;
  assign new_P1_R1165_U347 = ~new_P1_R1165_U331 | ~new_P1_R1165_U36;
  assign new_P1_R1165_U348 = ~new_P1_R1165_U340 | ~new_P1_R1165_U195;
  assign new_P1_R1165_U349 = ~new_P1_R1165_U257 | ~new_P1_R1165_U41;
  assign new_P1_R1165_U350 = ~new_P1_U3177 | ~new_P1_R1165_U60;
  assign new_P1_R1165_U351 = ~new_P1_R1165_U120 | ~new_P1_R1165_U352 | ~new_P1_R1165_U304;
  assign new_P1_R1165_U352 = ~new_P1_R1165_U301 | ~new_P1_R1165_U193;
  assign new_P1_R1165_U353 = ~new_P1_U3172 | ~new_P1_R1165_U57;
  assign new_P1_R1165_U354 = ~new_P1_R1165_U69 | ~new_P1_R1165_U300;
  assign new_P1_R1165_U355 = ~new_P1_U3155 | ~new_P1_R1165_U300;
  assign new_P1_R1165_U356 = ~new_P1_R1165_U308 | ~new_P1_R1165_U301 | ~new_P1_R1165_U193;
  assign new_P1_R1165_U357 = ~new_P1_R1165_U121 | ~new_P1_R1165_U176 | ~new_P1_R1165_U193;
  assign new_P1_R1165_U358 = ~new_P1_R1165_U302 | ~new_P1_R1165_U308;
  assign new_P1_R1165_U359 = ~new_P1_U3154 | ~new_P1_R1165_U67;
  assign new_P1_R1165_U360 = ~new_P1_R1165_U128 | ~new_P1_R1165_U310;
  assign new_P1_R1165_U361 = ~new_P1_R1165_U216 | ~new_P1_R1165_U153;
  assign new_P1_R1165_U362 = ~new_P1_R1165_U151;
  assign new_P1_R1165_U363 = ~new_P1_R1165_U247 | ~new_P1_R1165_U147;
  assign new_P1_R1165_U364 = ~new_P1_R1165_U192;
  assign new_P1_R1165_U365 = ~new_P1_U3211 | ~new_P1_R1165_U136;
  assign new_P1_R1165_U366 = ~new_P1_U3201 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U367 = ~new_P1_R1165_U57;
  assign new_P1_R1165_U368 = ~new_P1_R1165_U367 | ~new_P1_U3172;
  assign new_P1_R1165_U369 = ~new_P1_R1165_U57 | ~new_P1_R1165_U28;
  assign new_P1_R1165_U370 = ~new_P1_R1165_U367 | ~new_P1_U3172;
  assign new_P1_R1165_U371 = ~new_P1_R1165_U57 | ~new_P1_R1165_U28;
  assign new_P1_R1165_U372 = ~new_P1_R1165_U371 | ~new_P1_R1165_U370;
  assign new_P1_R1165_U373 = ~new_P1_U3211 | ~new_P1_R1165_U138;
  assign new_P1_R1165_U374 = ~new_P1_U3206 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U375 = ~new_P1_R1165_U60;
  assign new_P1_R1165_U376 = ~new_P1_U3211 | ~new_P1_R1165_U139;
  assign new_P1_R1165_U377 = ~new_P1_U3210 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U378 = ~new_P1_R1165_U63;
  assign new_P1_R1165_U379 = ~new_P1_U3211 | ~new_P1_R1165_U140;
  assign new_P1_R1165_U380 = ~new_P1_U3209 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U381 = ~new_P1_R1165_U64;
  assign new_P1_R1165_U382 = ~new_P1_U3211 | ~new_P1_R1165_U141;
  assign new_P1_R1165_U383 = ~new_P1_U3207 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U384 = ~new_P1_R1165_U62;
  assign new_P1_R1165_U385 = ~new_P1_U3211 | ~new_P1_R1165_U142;
  assign new_P1_R1165_U386 = ~new_P1_U3208 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U387 = ~new_P1_R1165_U61;
  assign new_P1_R1165_U388 = ~new_P1_U3211 | ~new_P1_R1165_U143;
  assign new_P1_R1165_U389 = ~new_P1_U3205 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U390 = ~new_P1_R1165_U65;
  assign new_P1_R1165_U391 = ~new_P1_U3211 | ~new_P1_R1165_U144;
  assign new_P1_R1165_U392 = ~new_P1_U3203 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U393 = ~new_P1_R1165_U59;
  assign new_P1_R1165_U394 = ~new_P1_U3211 | ~new_P1_R1165_U145;
  assign new_P1_R1165_U395 = ~new_P1_U3204 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U396 = ~new_P1_R1165_U58;
  assign new_P1_R1165_U397 = ~new_P1_U3211 | ~new_P1_R1165_U146;
  assign new_P1_R1165_U398 = ~new_P1_U3202 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U399 = ~new_P1_R1165_U66;
  assign new_P1_R1165_U400 = ~new_P1_R1165_U137 | ~new_P1_R1165_U147;
  assign new_P1_R1165_U401 = ~new_P1_R1165_U232 | ~new_P1_R1165_U372;
  assign new_P1_R1165_U402 = ~new_P1_R1165_U399 | ~new_P1_U3173;
  assign new_P1_R1165_U403 = ~new_P1_R1165_U66 | ~new_P1_R1165_U27;
  assign new_P1_R1165_U404 = ~new_P1_R1165_U399 | ~new_P1_U3173;
  assign new_P1_R1165_U405 = ~new_P1_R1165_U66 | ~new_P1_R1165_U27;
  assign new_P1_R1165_U406 = ~new_P1_R1165_U405 | ~new_P1_R1165_U404;
  assign new_P1_R1165_U407 = ~new_P1_R1165_U148 | ~new_P1_R1165_U149;
  assign new_P1_R1165_U408 = ~new_P1_R1165_U228 | ~new_P1_R1165_U406;
  assign new_P1_R1165_U409 = ~new_P1_R1165_U393 | ~new_P1_U3174;
  assign new_P1_R1165_U410 = ~new_P1_R1165_U59 | ~new_P1_R1165_U19;
  assign new_P1_R1165_U411 = ~new_P1_R1165_U396 | ~new_P1_U3175;
  assign new_P1_R1165_U412 = ~new_P1_R1165_U58 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U413 = ~new_P1_R1165_U412 | ~new_P1_R1165_U411;
  assign new_P1_R1165_U414 = ~new_P1_R1165_U341 | ~new_P1_R1165_U29;
  assign new_P1_R1165_U415 = ~new_P1_R1165_U413 | ~new_P1_R1165_U220;
  assign new_P1_R1165_U416 = ~new_P1_R1165_U390 | ~new_P1_U3176;
  assign new_P1_R1165_U417 = ~new_P1_R1165_U65 | ~new_P1_R1165_U26;
  assign new_P1_R1165_U418 = ~new_P1_R1165_U390 | ~new_P1_U3176;
  assign new_P1_R1165_U419 = ~new_P1_R1165_U65 | ~new_P1_R1165_U26;
  assign new_P1_R1165_U420 = ~new_P1_R1165_U419 | ~new_P1_R1165_U418;
  assign new_P1_R1165_U421 = ~new_P1_R1165_U150 | ~new_P1_R1165_U151;
  assign new_P1_R1165_U422 = ~new_P1_R1165_U362 | ~new_P1_R1165_U420;
  assign new_P1_R1165_U423 = ~new_P1_R1165_U375 | ~new_P1_U3177;
  assign new_P1_R1165_U424 = ~new_P1_R1165_U60 | ~new_P1_R1165_U20;
  assign new_P1_R1165_U425 = ~new_P1_R1165_U375 | ~new_P1_U3177;
  assign new_P1_R1165_U426 = ~new_P1_R1165_U60 | ~new_P1_R1165_U20;
  assign new_P1_R1165_U427 = ~new_P1_R1165_U426 | ~new_P1_R1165_U425;
  assign new_P1_R1165_U428 = ~new_P1_R1165_U152 | ~new_P1_R1165_U153;
  assign new_P1_R1165_U429 = ~new_P1_R1165_U215 | ~new_P1_R1165_U427;
  assign new_P1_R1165_U430 = ~new_P1_R1165_U384 | ~new_P1_U3178;
  assign new_P1_R1165_U431 = ~new_P1_R1165_U62 | ~new_P1_R1165_U23;
  assign new_P1_R1165_U432 = ~new_P1_R1165_U387 | ~new_P1_U3179;
  assign new_P1_R1165_U433 = ~new_P1_R1165_U61 | ~new_P1_R1165_U21;
  assign new_P1_R1165_U434 = ~new_P1_R1165_U433 | ~new_P1_R1165_U432;
  assign new_P1_R1165_U435 = ~new_P1_R1165_U342 | ~new_P1_R1165_U30;
  assign new_P1_R1165_U436 = ~new_P1_R1165_U434 | ~new_P1_R1165_U208;
  assign new_P1_R1165_U437 = ~new_P1_U3211 | ~new_P1_R1165_U154;
  assign new_P1_R1165_U438 = ~new_P1_U3183 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U439 = ~new_P1_R1165_U67;
  assign new_P1_R1165_U440 = ~new_P1_U3211 | ~new_P1_R1165_U155;
  assign new_P1_R1165_U441 = ~new_P1_U3185 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U442 = ~new_P1_R1165_U68;
  assign new_P1_R1165_U443 = ~new_P1_U3211 | ~new_P1_R1165_U156;
  assign new_P1_R1165_U444 = ~new_P1_U3184 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U445 = ~new_P1_R1165_U69;
  assign new_P1_R1165_U446 = ~new_P1_U3211 | ~new_P1_R1165_U157;
  assign new_P1_R1165_U447 = ~new_P1_U3186 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U448 = ~new_P1_R1165_U70;
  assign new_P1_R1165_U449 = ~new_P1_U3211 | ~new_P1_R1165_U158;
  assign new_P1_R1165_U450 = ~new_P1_U3200 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U451 = ~new_P1_R1165_U73;
  assign new_P1_R1165_U452 = ~new_P1_U3211 | ~new_P1_R1165_U159;
  assign new_P1_R1165_U453 = ~new_P1_U3197 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U454 = ~new_P1_R1165_U75;
  assign new_P1_R1165_U455 = ~new_P1_U3211 | ~new_P1_R1165_U160;
  assign new_P1_R1165_U456 = ~new_P1_U3198 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U457 = ~new_P1_R1165_U76;
  assign new_P1_R1165_U458 = ~new_P1_U3211 | ~new_P1_R1165_U161;
  assign new_P1_R1165_U459 = ~new_P1_U3199 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U460 = ~new_P1_R1165_U74;
  assign new_P1_R1165_U461 = ~new_P1_U3211 | ~new_P1_R1165_U162;
  assign new_P1_R1165_U462 = ~new_P1_U3196 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U463 = ~new_P1_R1165_U77;
  assign new_P1_R1165_U464 = ~new_P1_U3211 | ~new_P1_R1165_U163;
  assign new_P1_R1165_U465 = ~new_P1_U3195 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U466 = ~new_P1_R1165_U78;
  assign new_P1_R1165_U467 = ~new_P1_U3211 | ~new_P1_R1165_U164;
  assign new_P1_R1165_U468 = ~new_P1_U3193 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U469 = ~new_P1_R1165_U72;
  assign new_P1_R1165_U470 = ~new_P1_U3211 | ~new_P1_R1165_U165;
  assign new_P1_R1165_U471 = ~new_P1_U3194 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U472 = ~new_P1_R1165_U71;
  assign new_P1_R1165_U473 = ~new_P1_U3211 | ~new_P1_R1165_U166;
  assign new_P1_R1165_U474 = ~new_P1_U3192 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U475 = ~new_P1_R1165_U79;
  assign new_P1_R1165_U476 = ~new_P1_U3211 | ~new_P1_R1165_U167;
  assign new_P1_R1165_U477 = ~new_P1_U3189 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U478 = ~new_P1_R1165_U81;
  assign new_P1_R1165_U479 = ~new_P1_U3211 | ~new_P1_R1165_U168;
  assign new_P1_R1165_U480 = ~new_P1_U3190 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U481 = ~new_P1_R1165_U82;
  assign new_P1_R1165_U482 = ~new_P1_U3211 | ~new_P1_R1165_U169;
  assign new_P1_R1165_U483 = ~new_P1_U3191 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U484 = ~new_P1_R1165_U80;
  assign new_P1_R1165_U485 = ~new_P1_U3211 | ~new_P1_R1165_U170;
  assign new_P1_R1165_U486 = ~new_P1_U3188 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U487 = ~new_P1_R1165_U83;
  assign new_P1_R1165_U488 = ~new_P1_U3211 | ~new_P1_R1165_U171;
  assign new_P1_R1165_U489 = ~new_P1_U3187 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U490 = ~new_P1_R1165_U84;
  assign new_P1_R1165_U491 = ~new_P1_U3211 | ~new_P1_R1165_U172;
  assign new_P1_R1165_U492 = ~new_P1_U3153 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U493 = ~new_P1_R1165_U123;
  assign new_P1_R1165_U494 = ~new_P1_U3182 | ~new_P1_R1165_U493;
  assign new_P1_R1165_U495 = ~new_P1_R1165_U123 | ~new_P1_R1165_U173;
  assign new_P1_R1165_U496 = ~new_P1_R1165_U85;
  assign new_P1_R1165_U497 = ~new_P1_R1165_U496 | ~new_P1_R1165_U351 | ~new_P1_R1165_U306;
  assign new_P1_R1165_U498 = ~new_P1_R1165_U85 | ~new_P1_R1165_U122 | ~new_P1_R1165_U358 | ~new_P1_R1165_U357;
  assign new_P1_R1165_U499 = ~new_P1_R1165_U439 | ~new_P1_U3154;
  assign new_P1_R1165_U500 = ~new_P1_R1165_U67 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U501 = ~new_P1_R1165_U439 | ~new_P1_U3154;
  assign new_P1_R1165_U502 = ~new_P1_R1165_U67 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U503 = ~new_P1_R1165_U502 | ~new_P1_R1165_U501;
  assign new_P1_R1165_U504 = ~new_P1_R1165_U174 | ~new_P1_R1165_U175;
  assign new_P1_R1165_U505 = ~new_P1_R1165_U305 | ~new_P1_R1165_U503;
  assign new_P1_R1165_U506 = ~new_P1_R1165_U445 | ~new_P1_U3155;
  assign new_P1_R1165_U507 = ~new_P1_R1165_U69 | ~new_P1_R1165_U32;
  assign new_P1_R1165_U508 = ~new_P1_R1165_U442 | ~new_P1_U3156;
  assign new_P1_R1165_U509 = ~new_P1_R1165_U68 | ~new_P1_R1165_U33;
  assign new_P1_R1165_U510 = ~new_P1_R1165_U509 | ~new_P1_R1165_U508;
  assign new_P1_R1165_U511 = ~new_P1_R1165_U343 | ~new_P1_R1165_U53;
  assign new_P1_R1165_U512 = ~new_P1_R1165_U510 | ~new_P1_R1165_U310;
  assign new_P1_R1165_U513 = ~new_P1_R1165_U448 | ~new_P1_U3157;
  assign new_P1_R1165_U514 = ~new_P1_R1165_U70 | ~new_P1_R1165_U34;
  assign new_P1_R1165_U515 = ~new_P1_R1165_U514 | ~new_P1_R1165_U513;
  assign new_P1_R1165_U516 = ~new_P1_R1165_U344 | ~new_P1_R1165_U176;
  assign new_P1_R1165_U517 = ~new_P1_R1165_U299 | ~new_P1_R1165_U515;
  assign new_P1_R1165_U518 = ~new_P1_R1165_U490 | ~new_P1_U3158;
  assign new_P1_R1165_U519 = ~new_P1_R1165_U84 | ~new_P1_R1165_U51;
  assign new_P1_R1165_U520 = ~new_P1_R1165_U490 | ~new_P1_U3158;
  assign new_P1_R1165_U521 = ~new_P1_R1165_U84 | ~new_P1_R1165_U51;
  assign new_P1_R1165_U522 = ~new_P1_R1165_U521 | ~new_P1_R1165_U520;
  assign new_P1_R1165_U523 = ~new_P1_R1165_U177 | ~new_P1_R1165_U178;
  assign new_P1_R1165_U524 = ~new_P1_R1165_U295 | ~new_P1_R1165_U522;
  assign new_P1_R1165_U525 = ~new_P1_R1165_U487 | ~new_P1_U3159;
  assign new_P1_R1165_U526 = ~new_P1_R1165_U83 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U527 = ~new_P1_R1165_U487 | ~new_P1_U3159;
  assign new_P1_R1165_U528 = ~new_P1_R1165_U83 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U529 = ~new_P1_R1165_U528 | ~new_P1_R1165_U527;
  assign new_P1_R1165_U530 = ~new_P1_R1165_U179 | ~new_P1_R1165_U180;
  assign new_P1_R1165_U531 = ~new_P1_R1165_U291 | ~new_P1_R1165_U529;
  assign new_P1_R1165_U532 = ~new_P1_R1165_U478 | ~new_P1_U3160;
  assign new_P1_R1165_U533 = ~new_P1_R1165_U81 | ~new_P1_R1165_U49;
  assign new_P1_R1165_U534 = ~new_P1_R1165_U481 | ~new_P1_U3161;
  assign new_P1_R1165_U535 = ~new_P1_R1165_U82 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U536 = ~new_P1_R1165_U535 | ~new_P1_R1165_U534;
  assign new_P1_R1165_U537 = ~new_P1_R1165_U345 | ~new_P1_R1165_U54;
  assign new_P1_R1165_U538 = ~new_P1_R1165_U536 | ~new_P1_R1165_U317;
  assign new_P1_R1165_U539 = ~new_P1_R1165_U381 | ~new_P1_U3180;
  assign new_P1_R1165_U540 = ~new_P1_R1165_U64 | ~new_P1_R1165_U25;
  assign new_P1_R1165_U541 = ~new_P1_R1165_U381 | ~new_P1_U3180;
  assign new_P1_R1165_U542 = ~new_P1_R1165_U64 | ~new_P1_R1165_U25;
  assign new_P1_R1165_U543 = ~new_P1_R1165_U542 | ~new_P1_R1165_U541;
  assign new_P1_R1165_U544 = ~new_P1_R1165_U181 | ~new_P1_R1165_U182;
  assign new_P1_R1165_U545 = ~new_P1_R1165_U204 | ~new_P1_R1165_U543;
  assign new_P1_R1165_U546 = ~new_P1_R1165_U484 | ~new_P1_U3162;
  assign new_P1_R1165_U547 = ~new_P1_R1165_U80 | ~new_P1_R1165_U47;
  assign new_P1_R1165_U548 = ~new_P1_R1165_U547 | ~new_P1_R1165_U546;
  assign new_P1_R1165_U549 = ~new_P1_R1165_U346 | ~new_P1_R1165_U183;
  assign new_P1_R1165_U550 = ~new_P1_R1165_U281 | ~new_P1_R1165_U548;
  assign new_P1_R1165_U551 = ~new_P1_R1165_U475 | ~new_P1_U3163;
  assign new_P1_R1165_U552 = ~new_P1_R1165_U79 | ~new_P1_R1165_U45;
  assign new_P1_R1165_U553 = ~new_P1_R1165_U475 | ~new_P1_U3163;
  assign new_P1_R1165_U554 = ~new_P1_R1165_U79 | ~new_P1_R1165_U45;
  assign new_P1_R1165_U555 = ~new_P1_R1165_U554 | ~new_P1_R1165_U553;
  assign new_P1_R1165_U556 = ~new_P1_R1165_U184 | ~new_P1_R1165_U185;
  assign new_P1_R1165_U557 = ~new_P1_R1165_U277 | ~new_P1_R1165_U555;
  assign new_P1_R1165_U558 = ~new_P1_R1165_U469 | ~new_P1_U3164;
  assign new_P1_R1165_U559 = ~new_P1_R1165_U72 | ~new_P1_R1165_U37;
  assign new_P1_R1165_U560 = ~new_P1_R1165_U472 | ~new_P1_U3165;
  assign new_P1_R1165_U561 = ~new_P1_R1165_U71 | ~new_P1_R1165_U35;
  assign new_P1_R1165_U562 = ~new_P1_R1165_U561 | ~new_P1_R1165_U560;
  assign new_P1_R1165_U563 = ~new_P1_R1165_U347 | ~new_P1_R1165_U55;
  assign new_P1_R1165_U564 = ~new_P1_R1165_U562 | ~new_P1_R1165_U269;
  assign new_P1_R1165_U565 = ~new_P1_R1165_U466 | ~new_P1_U3166;
  assign new_P1_R1165_U566 = ~new_P1_R1165_U78 | ~new_P1_R1165_U44;
  assign new_P1_R1165_U567 = ~new_P1_R1165_U466 | ~new_P1_U3166;
  assign new_P1_R1165_U568 = ~new_P1_R1165_U78 | ~new_P1_R1165_U44;
  assign new_P1_R1165_U569 = ~new_P1_R1165_U568 | ~new_P1_R1165_U567;
  assign new_P1_R1165_U570 = ~new_P1_R1165_U186 | ~new_P1_R1165_U187;
  assign new_P1_R1165_U571 = ~new_P1_R1165_U265 | ~new_P1_R1165_U569;
  assign new_P1_R1165_U572 = ~new_P1_R1165_U463 | ~new_P1_U3167;
  assign new_P1_R1165_U573 = ~new_P1_R1165_U77 | ~new_P1_R1165_U43;
  assign new_P1_R1165_U574 = ~new_P1_R1165_U463 | ~new_P1_U3167;
  assign new_P1_R1165_U575 = ~new_P1_R1165_U77 | ~new_P1_R1165_U43;
  assign new_P1_R1165_U576 = ~new_P1_R1165_U575 | ~new_P1_R1165_U574;
  assign new_P1_R1165_U577 = ~new_P1_R1165_U188 | ~new_P1_R1165_U189;
  assign new_P1_R1165_U578 = ~new_P1_R1165_U261 | ~new_P1_R1165_U576;
  assign new_P1_R1165_U579 = ~new_P1_R1165_U454 | ~new_P1_U3168;
  assign new_P1_R1165_U580 = ~new_P1_R1165_U75 | ~new_P1_R1165_U42;
  assign new_P1_R1165_U581 = ~new_P1_R1165_U457 | ~new_P1_U3169;
  assign new_P1_R1165_U582 = ~new_P1_R1165_U76 | ~new_P1_R1165_U39;
  assign new_P1_R1165_U583 = ~new_P1_R1165_U582 | ~new_P1_R1165_U581;
  assign new_P1_R1165_U584 = ~new_P1_R1165_U348 | ~new_P1_R1165_U56;
  assign new_P1_R1165_U585 = ~new_P1_R1165_U583 | ~new_P1_R1165_U333;
  assign new_P1_R1165_U586 = ~new_P1_R1165_U460 | ~new_P1_U3170;
  assign new_P1_R1165_U587 = ~new_P1_R1165_U74 | ~new_P1_R1165_U40;
  assign new_P1_R1165_U588 = ~new_P1_R1165_U587 | ~new_P1_R1165_U586;
  assign new_P1_R1165_U589 = ~new_P1_R1165_U349 | ~new_P1_R1165_U190;
  assign new_P1_R1165_U590 = ~new_P1_R1165_U251 | ~new_P1_R1165_U588;
  assign new_P1_R1165_U591 = ~new_P1_R1165_U451 | ~new_P1_U3171;
  assign new_P1_R1165_U592 = ~new_P1_R1165_U73 | ~new_P1_R1165_U38;
  assign new_P1_R1165_U593 = ~new_P1_R1165_U451 | ~new_P1_U3171;
  assign new_P1_R1165_U594 = ~new_P1_R1165_U73 | ~new_P1_R1165_U38;
  assign new_P1_R1165_U595 = ~new_P1_R1165_U594 | ~new_P1_R1165_U593;
  assign new_P1_R1165_U596 = ~new_P1_R1165_U191 | ~new_P1_R1165_U192;
  assign new_P1_R1165_U597 = ~new_P1_R1165_U364 | ~new_P1_R1165_U595;
  assign new_P1_R1165_U598 = ~new_P1_U3181 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U599 = ~new_P1_U3211 | ~new_P1_R1165_U24;
  assign new_P1_R1165_U600 = ~new_P1_R1165_U135;
  assign new_P1_R1165_U601 = ~new_P1_R1165_U63 | ~new_P1_R1165_U600;
  assign new_P1_R1165_U602 = ~new_P1_R1165_U135 | ~new_P1_R1165_U378;
  assign new_P1_R1150_U6 = new_P1_R1150_U198 & new_P1_R1150_U197;
  assign new_P1_R1150_U7 = new_P1_R1150_U237 & new_P1_R1150_U236;
  assign new_P1_R1150_U8 = new_P1_R1150_U254 & new_P1_R1150_U253;
  assign new_P1_R1150_U9 = new_P1_R1150_U280 & new_P1_R1150_U279;
  assign new_P1_R1150_U10 = ~new_P1_R1150_U340 | ~new_P1_R1150_U343;
  assign new_P1_R1150_U11 = ~new_P1_R1150_U329 | ~new_P1_R1150_U332;
  assign new_P1_R1150_U12 = ~new_P1_R1150_U318 | ~new_P1_R1150_U321;
  assign new_P1_R1150_U13 = ~new_P1_R1150_U310 | ~new_P1_R1150_U312;
  assign new_P1_R1150_U14 = ~new_P1_R1150_U347 | ~new_P1_R1150_U308;
  assign new_P1_R1150_U15 = ~new_P1_R1150_U231 | ~new_P1_R1150_U233;
  assign new_P1_R1150_U16 = ~new_P1_R1150_U223 | ~new_P1_R1150_U226;
  assign new_P1_R1150_U17 = ~new_P1_R1150_U215 | ~new_P1_R1150_U217;
  assign new_P1_R1150_U18 = ~new_P1_R1150_U23 | ~new_P1_R1150_U346;
  assign new_P1_R1150_U19 = ~new_P1_U3473;
  assign new_P1_R1150_U20 = ~new_P1_U3467;
  assign new_P1_R1150_U21 = ~new_P1_U3458;
  assign new_P1_R1150_U22 = ~new_P1_U3450;
  assign new_P1_R1150_U23 = ~new_P1_U3450 | ~new_P1_R1150_U91;
  assign new_P1_R1150_U24 = ~new_P1_U3078;
  assign new_P1_R1150_U25 = ~new_P1_U3461;
  assign new_P1_R1150_U26 = ~new_P1_U3068;
  assign new_P1_R1150_U27 = ~new_P1_U3068 | ~new_P1_R1150_U21;
  assign new_P1_R1150_U28 = ~new_P1_U3064;
  assign new_P1_R1150_U29 = ~new_P1_U3470;
  assign new_P1_R1150_U30 = ~new_P1_U3464;
  assign new_P1_R1150_U31 = ~new_P1_U3071;
  assign new_P1_R1150_U32 = ~new_P1_U3067;
  assign new_P1_R1150_U33 = ~new_P1_U3060;
  assign new_P1_R1150_U34 = ~new_P1_U3060 | ~new_P1_R1150_U30;
  assign new_P1_R1150_U35 = ~new_P1_U3476;
  assign new_P1_R1150_U36 = ~new_P1_U3070;
  assign new_P1_R1150_U37 = ~new_P1_U3070 | ~new_P1_R1150_U19;
  assign new_P1_R1150_U38 = ~new_P1_U3084;
  assign new_P1_R1150_U39 = ~new_P1_U3479;
  assign new_P1_R1150_U40 = ~new_P1_U3083;
  assign new_P1_R1150_U41 = ~new_P1_R1150_U204 | ~new_P1_R1150_U203;
  assign new_P1_R1150_U42 = ~new_P1_R1150_U34 | ~new_P1_R1150_U219;
  assign new_P1_R1150_U43 = ~new_P1_R1150_U188 | ~new_P1_R1150_U187;
  assign new_P1_R1150_U44 = ~new_P1_U3976;
  assign new_P1_R1150_U45 = ~new_P1_U3980;
  assign new_P1_R1150_U46 = ~new_P1_U3497;
  assign new_P1_R1150_U47 = ~new_P1_U3482;
  assign new_P1_R1150_U48 = ~new_P1_U3485;
  assign new_P1_R1150_U49 = ~new_P1_U3063;
  assign new_P1_R1150_U50 = ~new_P1_U3062;
  assign new_P1_R1150_U51 = ~new_P1_U3083 | ~new_P1_R1150_U39;
  assign new_P1_R1150_U52 = ~new_P1_U3488;
  assign new_P1_R1150_U53 = ~new_P1_U3072;
  assign new_P1_R1150_U54 = ~new_P1_U3491;
  assign new_P1_R1150_U55 = ~new_P1_U3080;
  assign new_P1_R1150_U56 = ~new_P1_U3500;
  assign new_P1_R1150_U57 = ~new_P1_U3494;
  assign new_P1_R1150_U58 = ~new_P1_U3073;
  assign new_P1_R1150_U59 = ~new_P1_U3074;
  assign new_P1_R1150_U60 = ~new_P1_U3079;
  assign new_P1_R1150_U61 = ~new_P1_U3079 | ~new_P1_R1150_U57;
  assign new_P1_R1150_U62 = ~new_P1_U3503;
  assign new_P1_R1150_U63 = ~new_P1_U3069;
  assign new_P1_R1150_U64 = ~new_P1_R1150_U264 | ~new_P1_R1150_U263;
  assign new_P1_R1150_U65 = ~new_P1_U3082;
  assign new_P1_R1150_U66 = ~new_P1_U3508;
  assign new_P1_R1150_U67 = ~new_P1_U3081;
  assign new_P1_R1150_U68 = ~new_P1_U3982;
  assign new_P1_R1150_U69 = ~new_P1_U3076;
  assign new_P1_R1150_U70 = ~new_P1_U3979;
  assign new_P1_R1150_U71 = ~new_P1_U3981;
  assign new_P1_R1150_U72 = ~new_P1_U3066;
  assign new_P1_R1150_U73 = ~new_P1_U3061;
  assign new_P1_R1150_U74 = ~new_P1_U3075;
  assign new_P1_R1150_U75 = ~new_P1_U3075 | ~new_P1_R1150_U71;
  assign new_P1_R1150_U76 = ~new_P1_U3978;
  assign new_P1_R1150_U77 = ~new_P1_U3065;
  assign new_P1_R1150_U78 = ~new_P1_U3977;
  assign new_P1_R1150_U79 = ~new_P1_U3058;
  assign new_P1_R1150_U80 = ~new_P1_U3975;
  assign new_P1_R1150_U81 = ~new_P1_U3057;
  assign new_P1_R1150_U82 = ~new_P1_U3057 | ~new_P1_R1150_U44;
  assign new_P1_R1150_U83 = ~new_P1_U3053;
  assign new_P1_R1150_U84 = ~new_P1_U3974;
  assign new_P1_R1150_U85 = ~new_P1_U3054;
  assign new_P1_R1150_U86 = ~new_P1_R1150_U126 | ~new_P1_R1150_U297;
  assign new_P1_R1150_U87 = ~new_P1_R1150_U294 | ~new_P1_R1150_U293;
  assign new_P1_R1150_U88 = ~new_P1_R1150_U75 | ~new_P1_R1150_U314;
  assign new_P1_R1150_U89 = ~new_P1_R1150_U61 | ~new_P1_R1150_U325;
  assign new_P1_R1150_U90 = ~new_P1_R1150_U51 | ~new_P1_R1150_U336;
  assign new_P1_R1150_U91 = ~new_P1_U3077;
  assign new_P1_R1150_U92 = ~new_P1_R1150_U390 | ~new_P1_R1150_U389;
  assign new_P1_R1150_U93 = ~new_P1_R1150_U404 | ~new_P1_R1150_U403;
  assign new_P1_R1150_U94 = ~new_P1_R1150_U409 | ~new_P1_R1150_U408;
  assign new_P1_R1150_U95 = ~new_P1_R1150_U425 | ~new_P1_R1150_U424;
  assign new_P1_R1150_U96 = ~new_P1_R1150_U430 | ~new_P1_R1150_U429;
  assign new_P1_R1150_U97 = ~new_P1_R1150_U435 | ~new_P1_R1150_U434;
  assign new_P1_R1150_U98 = ~new_P1_R1150_U440 | ~new_P1_R1150_U439;
  assign new_P1_R1150_U99 = ~new_P1_R1150_U445 | ~new_P1_R1150_U444;
  assign new_P1_R1150_U100 = ~new_P1_R1150_U461 | ~new_P1_R1150_U460;
  assign new_P1_R1150_U101 = ~new_P1_R1150_U466 | ~new_P1_R1150_U465;
  assign new_P1_R1150_U102 = ~new_P1_R1150_U351 | ~new_P1_R1150_U350;
  assign new_P1_R1150_U103 = ~new_P1_R1150_U360 | ~new_P1_R1150_U359;
  assign new_P1_R1150_U104 = ~new_P1_R1150_U367 | ~new_P1_R1150_U366;
  assign new_P1_R1150_U105 = ~new_P1_R1150_U371 | ~new_P1_R1150_U370;
  assign new_P1_R1150_U106 = ~new_P1_R1150_U380 | ~new_P1_R1150_U379;
  assign new_P1_R1150_U107 = ~new_P1_R1150_U399 | ~new_P1_R1150_U398;
  assign new_P1_R1150_U108 = ~new_P1_R1150_U416 | ~new_P1_R1150_U415;
  assign new_P1_R1150_U109 = ~new_P1_R1150_U420 | ~new_P1_R1150_U419;
  assign new_P1_R1150_U110 = ~new_P1_R1150_U452 | ~new_P1_R1150_U451;
  assign new_P1_R1150_U111 = ~new_P1_R1150_U456 | ~new_P1_R1150_U455;
  assign new_P1_R1150_U112 = ~new_P1_R1150_U473 | ~new_P1_R1150_U472;
  assign new_P1_R1150_U113 = new_P1_R1150_U193 & new_P1_R1150_U194;
  assign new_P1_R1150_U114 = new_P1_R1150_U201 & new_P1_R1150_U196;
  assign new_P1_R1150_U115 = new_P1_R1150_U206 & new_P1_R1150_U180;
  assign new_P1_R1150_U116 = new_P1_R1150_U209 & new_P1_R1150_U210;
  assign new_P1_R1150_U117 = new_P1_R1150_U37 & new_P1_R1150_U353 & new_P1_R1150_U352;
  assign new_P1_R1150_U118 = new_P1_R1150_U356 & new_P1_R1150_U180;
  assign new_P1_R1150_U119 = new_P1_R1150_U225 & new_P1_R1150_U6;
  assign new_P1_R1150_U120 = new_P1_R1150_U363 & new_P1_R1150_U179;
  assign new_P1_R1150_U121 = new_P1_R1150_U27 & new_P1_R1150_U373 & new_P1_R1150_U372;
  assign new_P1_R1150_U122 = new_P1_R1150_U376 & new_P1_R1150_U178;
  assign new_P1_R1150_U123 = new_P1_R1150_U174 & new_P1_R1150_U235 & new_P1_R1150_U212;
  assign new_P1_R1150_U124 = new_P1_R1150_U252 & new_P1_R1150_U257 & new_P1_R1150_U175;
  assign new_P1_R1150_U125 = new_P1_R1150_U283 & new_P1_R1150_U176;
  assign new_P1_R1150_U126 = new_P1_R1150_U299 & new_P1_R1150_U300;
  assign new_P1_R1150_U127 = ~new_P1_R1150_U387 | ~new_P1_R1150_U386;
  assign new_P1_R1150_U128 = new_P1_R1150_U82 & new_P1_R1150_U392 & new_P1_R1150_U391;
  assign new_P1_R1150_U129 = new_P1_R1150_U395 & new_P1_R1150_U177;
  assign new_P1_R1150_U130 = ~new_P1_R1150_U401 | ~new_P1_R1150_U400;
  assign new_P1_R1150_U131 = ~new_P1_R1150_U406 | ~new_P1_R1150_U405;
  assign new_P1_R1150_U132 = new_P1_R1150_U412 & new_P1_R1150_U176;
  assign new_P1_R1150_U133 = ~new_P1_R1150_U422 | ~new_P1_R1150_U421;
  assign new_P1_R1150_U134 = ~new_P1_R1150_U427 | ~new_P1_R1150_U426;
  assign new_P1_R1150_U135 = ~new_P1_R1150_U432 | ~new_P1_R1150_U431;
  assign new_P1_R1150_U136 = ~new_P1_R1150_U437 | ~new_P1_R1150_U436;
  assign new_P1_R1150_U137 = ~new_P1_R1150_U442 | ~new_P1_R1150_U441;
  assign new_P1_R1150_U138 = new_P1_R1150_U331 & new_P1_R1150_U8;
  assign new_P1_R1150_U139 = new_P1_R1150_U448 & new_P1_R1150_U175;
  assign new_P1_R1150_U140 = ~new_P1_R1150_U458 | ~new_P1_R1150_U457;
  assign new_P1_R1150_U141 = ~new_P1_R1150_U463 | ~new_P1_R1150_U462;
  assign new_P1_R1150_U142 = new_P1_R1150_U342 & new_P1_R1150_U7;
  assign new_P1_R1150_U143 = new_P1_R1150_U469 & new_P1_R1150_U174;
  assign new_P1_R1150_U144 = new_P1_R1150_U349 & new_P1_R1150_U348;
  assign new_P1_R1150_U145 = ~new_P1_R1150_U116 | ~new_P1_R1150_U207;
  assign new_P1_R1150_U146 = new_P1_R1150_U358 & new_P1_R1150_U357;
  assign new_P1_R1150_U147 = new_P1_R1150_U365 & new_P1_R1150_U364;
  assign new_P1_R1150_U148 = new_P1_R1150_U369 & new_P1_R1150_U368;
  assign new_P1_R1150_U149 = ~new_P1_R1150_U113 | ~new_P1_R1150_U191;
  assign new_P1_R1150_U150 = new_P1_R1150_U378 & new_P1_R1150_U377;
  assign new_P1_R1150_U151 = ~new_P1_U3985;
  assign new_P1_R1150_U152 = ~new_P1_U3055;
  assign new_P1_R1150_U153 = new_P1_R1150_U382 & new_P1_R1150_U381;
  assign new_P1_R1150_U154 = new_P1_R1150_U397 & new_P1_R1150_U396;
  assign new_P1_R1150_U155 = ~new_P1_R1150_U290 | ~new_P1_R1150_U289;
  assign new_P1_R1150_U156 = ~new_P1_R1150_U286 | ~new_P1_R1150_U285;
  assign new_P1_R1150_U157 = new_P1_R1150_U414 & new_P1_R1150_U413;
  assign new_P1_R1150_U158 = new_P1_R1150_U418 & new_P1_R1150_U417;
  assign new_P1_R1150_U159 = ~new_P1_R1150_U276 | ~new_P1_R1150_U275;
  assign new_P1_R1150_U160 = ~new_P1_R1150_U272 | ~new_P1_R1150_U271;
  assign new_P1_R1150_U161 = ~new_P1_U3455;
  assign new_P1_R1150_U162 = ~new_P1_R1150_U268 | ~new_P1_R1150_U267;
  assign new_P1_R1150_U163 = ~new_P1_U3506;
  assign new_P1_R1150_U164 = ~new_P1_R1150_U260 | ~new_P1_R1150_U259;
  assign new_P1_R1150_U165 = new_P1_R1150_U450 & new_P1_R1150_U449;
  assign new_P1_R1150_U166 = new_P1_R1150_U454 & new_P1_R1150_U453;
  assign new_P1_R1150_U167 = ~new_P1_R1150_U250 | ~new_P1_R1150_U249;
  assign new_P1_R1150_U168 = ~new_P1_R1150_U246 | ~new_P1_R1150_U245;
  assign new_P1_R1150_U169 = ~new_P1_R1150_U242 | ~new_P1_R1150_U241;
  assign new_P1_R1150_U170 = new_P1_R1150_U471 & new_P1_R1150_U470;
  assign new_P1_R1150_U171 = ~new_P1_R1150_U82;
  assign new_P1_R1150_U172 = ~new_P1_R1150_U27;
  assign new_P1_R1150_U173 = ~new_P1_R1150_U37;
  assign new_P1_R1150_U174 = ~new_P1_U3482 | ~new_P1_R1150_U50;
  assign new_P1_R1150_U175 = ~new_P1_U3497 | ~new_P1_R1150_U59;
  assign new_P1_R1150_U176 = ~new_P1_U3980 | ~new_P1_R1150_U73;
  assign new_P1_R1150_U177 = ~new_P1_U3976 | ~new_P1_R1150_U81;
  assign new_P1_R1150_U178 = ~new_P1_U3458 | ~new_P1_R1150_U26;
  assign new_P1_R1150_U179 = ~new_P1_U3467 | ~new_P1_R1150_U32;
  assign new_P1_R1150_U180 = ~new_P1_U3473 | ~new_P1_R1150_U36;
  assign new_P1_R1150_U181 = ~new_P1_R1150_U61;
  assign new_P1_R1150_U182 = ~new_P1_R1150_U75;
  assign new_P1_R1150_U183 = ~new_P1_R1150_U34;
  assign new_P1_R1150_U184 = ~new_P1_R1150_U51;
  assign new_P1_R1150_U185 = ~new_P1_R1150_U23;
  assign new_P1_R1150_U186 = ~new_P1_R1150_U185 | ~new_P1_R1150_U24;
  assign new_P1_R1150_U187 = ~new_P1_R1150_U186 | ~new_P1_R1150_U161;
  assign new_P1_R1150_U188 = ~new_P1_U3078 | ~new_P1_R1150_U23;
  assign new_P1_R1150_U189 = ~new_P1_R1150_U43;
  assign new_P1_R1150_U190 = ~new_P1_U3461 | ~new_P1_R1150_U28;
  assign new_P1_R1150_U191 = ~new_P1_R1150_U190 | ~new_P1_R1150_U43 | ~new_P1_R1150_U178;
  assign new_P1_R1150_U192 = ~new_P1_R1150_U28 | ~new_P1_R1150_U27;
  assign new_P1_R1150_U193 = ~new_P1_R1150_U192 | ~new_P1_R1150_U25;
  assign new_P1_R1150_U194 = ~new_P1_U3064 | ~new_P1_R1150_U172;
  assign new_P1_R1150_U195 = ~new_P1_R1150_U149;
  assign new_P1_R1150_U196 = ~new_P1_U3470 | ~new_P1_R1150_U31;
  assign new_P1_R1150_U197 = ~new_P1_U3071 | ~new_P1_R1150_U29;
  assign new_P1_R1150_U198 = ~new_P1_U3067 | ~new_P1_R1150_U20;
  assign new_P1_R1150_U199 = ~new_P1_R1150_U183 | ~new_P1_R1150_U179;
  assign new_P1_R1150_U200 = ~new_P1_R1150_U6 | ~new_P1_R1150_U199;
  assign new_P1_R1150_U201 = ~new_P1_U3464 | ~new_P1_R1150_U33;
  assign new_P1_R1150_U202 = ~new_P1_U3470 | ~new_P1_R1150_U31;
  assign new_P1_R1150_U203 = ~new_P1_R1150_U114 | ~new_P1_R1150_U149 | ~new_P1_R1150_U179;
  assign new_P1_R1150_U204 = ~new_P1_R1150_U202 | ~new_P1_R1150_U200;
  assign new_P1_R1150_U205 = ~new_P1_R1150_U41;
  assign new_P1_R1150_U206 = ~new_P1_U3476 | ~new_P1_R1150_U38;
  assign new_P1_R1150_U207 = ~new_P1_R1150_U115 | ~new_P1_R1150_U41;
  assign new_P1_R1150_U208 = ~new_P1_R1150_U38 | ~new_P1_R1150_U37;
  assign new_P1_R1150_U209 = ~new_P1_R1150_U208 | ~new_P1_R1150_U35;
  assign new_P1_R1150_U210 = ~new_P1_U3084 | ~new_P1_R1150_U173;
  assign new_P1_R1150_U211 = ~new_P1_R1150_U145;
  assign new_P1_R1150_U212 = ~new_P1_U3479 | ~new_P1_R1150_U40;
  assign new_P1_R1150_U213 = ~new_P1_R1150_U212 | ~new_P1_R1150_U51;
  assign new_P1_R1150_U214 = ~new_P1_R1150_U205 | ~new_P1_R1150_U37;
  assign new_P1_R1150_U215 = ~new_P1_R1150_U118 | ~new_P1_R1150_U214;
  assign new_P1_R1150_U216 = ~new_P1_R1150_U41 | ~new_P1_R1150_U180;
  assign new_P1_R1150_U217 = ~new_P1_R1150_U117 | ~new_P1_R1150_U216;
  assign new_P1_R1150_U218 = ~new_P1_R1150_U37 | ~new_P1_R1150_U180;
  assign new_P1_R1150_U219 = ~new_P1_R1150_U201 | ~new_P1_R1150_U149;
  assign new_P1_R1150_U220 = ~new_P1_R1150_U42;
  assign new_P1_R1150_U221 = ~new_P1_U3067 | ~new_P1_R1150_U20;
  assign new_P1_R1150_U222 = ~new_P1_R1150_U220 | ~new_P1_R1150_U221;
  assign new_P1_R1150_U223 = ~new_P1_R1150_U120 | ~new_P1_R1150_U222;
  assign new_P1_R1150_U224 = ~new_P1_R1150_U42 | ~new_P1_R1150_U179;
  assign new_P1_R1150_U225 = ~new_P1_U3470 | ~new_P1_R1150_U31;
  assign new_P1_R1150_U226 = ~new_P1_R1150_U119 | ~new_P1_R1150_U224;
  assign new_P1_R1150_U227 = ~new_P1_U3067 | ~new_P1_R1150_U20;
  assign new_P1_R1150_U228 = ~new_P1_R1150_U179 | ~new_P1_R1150_U227;
  assign new_P1_R1150_U229 = ~new_P1_R1150_U201 | ~new_P1_R1150_U34;
  assign new_P1_R1150_U230 = ~new_P1_R1150_U189 | ~new_P1_R1150_U27;
  assign new_P1_R1150_U231 = ~new_P1_R1150_U122 | ~new_P1_R1150_U230;
  assign new_P1_R1150_U232 = ~new_P1_R1150_U43 | ~new_P1_R1150_U178;
  assign new_P1_R1150_U233 = ~new_P1_R1150_U121 | ~new_P1_R1150_U232;
  assign new_P1_R1150_U234 = ~new_P1_R1150_U27 | ~new_P1_R1150_U178;
  assign new_P1_R1150_U235 = ~new_P1_U3485 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U236 = ~new_P1_U3063 | ~new_P1_R1150_U48;
  assign new_P1_R1150_U237 = ~new_P1_U3062 | ~new_P1_R1150_U47;
  assign new_P1_R1150_U238 = ~new_P1_R1150_U184 | ~new_P1_R1150_U174;
  assign new_P1_R1150_U239 = ~new_P1_R1150_U7 | ~new_P1_R1150_U238;
  assign new_P1_R1150_U240 = ~new_P1_U3485 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U241 = ~new_P1_R1150_U145 | ~new_P1_R1150_U123;
  assign new_P1_R1150_U242 = ~new_P1_R1150_U240 | ~new_P1_R1150_U239;
  assign new_P1_R1150_U243 = ~new_P1_R1150_U169;
  assign new_P1_R1150_U244 = ~new_P1_U3488 | ~new_P1_R1150_U53;
  assign new_P1_R1150_U245 = ~new_P1_R1150_U244 | ~new_P1_R1150_U169;
  assign new_P1_R1150_U246 = ~new_P1_U3072 | ~new_P1_R1150_U52;
  assign new_P1_R1150_U247 = ~new_P1_R1150_U168;
  assign new_P1_R1150_U248 = ~new_P1_U3491 | ~new_P1_R1150_U55;
  assign new_P1_R1150_U249 = ~new_P1_R1150_U248 | ~new_P1_R1150_U168;
  assign new_P1_R1150_U250 = ~new_P1_U3080 | ~new_P1_R1150_U54;
  assign new_P1_R1150_U251 = ~new_P1_R1150_U167;
  assign new_P1_R1150_U252 = ~new_P1_U3500 | ~new_P1_R1150_U58;
  assign new_P1_R1150_U253 = ~new_P1_U3073 | ~new_P1_R1150_U56;
  assign new_P1_R1150_U254 = ~new_P1_U3074 | ~new_P1_R1150_U46;
  assign new_P1_R1150_U255 = ~new_P1_R1150_U181 | ~new_P1_R1150_U175;
  assign new_P1_R1150_U256 = ~new_P1_R1150_U8 | ~new_P1_R1150_U255;
  assign new_P1_R1150_U257 = ~new_P1_U3494 | ~new_P1_R1150_U60;
  assign new_P1_R1150_U258 = ~new_P1_U3500 | ~new_P1_R1150_U58;
  assign new_P1_R1150_U259 = ~new_P1_R1150_U167 | ~new_P1_R1150_U124;
  assign new_P1_R1150_U260 = ~new_P1_R1150_U258 | ~new_P1_R1150_U256;
  assign new_P1_R1150_U261 = ~new_P1_R1150_U164;
  assign new_P1_R1150_U262 = ~new_P1_U3503 | ~new_P1_R1150_U63;
  assign new_P1_R1150_U263 = ~new_P1_R1150_U262 | ~new_P1_R1150_U164;
  assign new_P1_R1150_U264 = ~new_P1_U3069 | ~new_P1_R1150_U62;
  assign new_P1_R1150_U265 = ~new_P1_R1150_U64;
  assign new_P1_R1150_U266 = ~new_P1_R1150_U265 | ~new_P1_R1150_U65;
  assign new_P1_R1150_U267 = ~new_P1_R1150_U266 | ~new_P1_R1150_U163;
  assign new_P1_R1150_U268 = ~new_P1_U3082 | ~new_P1_R1150_U64;
  assign new_P1_R1150_U269 = ~new_P1_R1150_U162;
  assign new_P1_R1150_U270 = ~new_P1_U3508 | ~new_P1_R1150_U67;
  assign new_P1_R1150_U271 = ~new_P1_R1150_U270 | ~new_P1_R1150_U162;
  assign new_P1_R1150_U272 = ~new_P1_U3081 | ~new_P1_R1150_U66;
  assign new_P1_R1150_U273 = ~new_P1_R1150_U160;
  assign new_P1_R1150_U274 = ~new_P1_U3982 | ~new_P1_R1150_U69;
  assign new_P1_R1150_U275 = ~new_P1_R1150_U274 | ~new_P1_R1150_U160;
  assign new_P1_R1150_U276 = ~new_P1_U3076 | ~new_P1_R1150_U68;
  assign new_P1_R1150_U277 = ~new_P1_R1150_U159;
  assign new_P1_R1150_U278 = ~new_P1_U3979 | ~new_P1_R1150_U72;
  assign new_P1_R1150_U279 = ~new_P1_U3066 | ~new_P1_R1150_U70;
  assign new_P1_R1150_U280 = ~new_P1_U3061 | ~new_P1_R1150_U45;
  assign new_P1_R1150_U281 = ~new_P1_R1150_U182 | ~new_P1_R1150_U176;
  assign new_P1_R1150_U282 = ~new_P1_R1150_U9 | ~new_P1_R1150_U281;
  assign new_P1_R1150_U283 = ~new_P1_U3981 | ~new_P1_R1150_U74;
  assign new_P1_R1150_U284 = ~new_P1_U3979 | ~new_P1_R1150_U72;
  assign new_P1_R1150_U285 = ~new_P1_R1150_U278 | ~new_P1_R1150_U159 | ~new_P1_R1150_U125;
  assign new_P1_R1150_U286 = ~new_P1_R1150_U284 | ~new_P1_R1150_U282;
  assign new_P1_R1150_U287 = ~new_P1_R1150_U156;
  assign new_P1_R1150_U288 = ~new_P1_U3978 | ~new_P1_R1150_U77;
  assign new_P1_R1150_U289 = ~new_P1_R1150_U288 | ~new_P1_R1150_U156;
  assign new_P1_R1150_U290 = ~new_P1_U3065 | ~new_P1_R1150_U76;
  assign new_P1_R1150_U291 = ~new_P1_R1150_U155;
  assign new_P1_R1150_U292 = ~new_P1_U3977 | ~new_P1_R1150_U79;
  assign new_P1_R1150_U293 = ~new_P1_R1150_U292 | ~new_P1_R1150_U155;
  assign new_P1_R1150_U294 = ~new_P1_U3058 | ~new_P1_R1150_U78;
  assign new_P1_R1150_U295 = ~new_P1_R1150_U87;
  assign new_P1_R1150_U296 = ~new_P1_U3975 | ~new_P1_R1150_U83;
  assign new_P1_R1150_U297 = ~new_P1_R1150_U296 | ~new_P1_R1150_U87 | ~new_P1_R1150_U177;
  assign new_P1_R1150_U298 = ~new_P1_R1150_U83 | ~new_P1_R1150_U82;
  assign new_P1_R1150_U299 = ~new_P1_R1150_U298 | ~new_P1_R1150_U80;
  assign new_P1_R1150_U300 = ~new_P1_U3053 | ~new_P1_R1150_U171;
  assign new_P1_R1150_U301 = ~new_P1_R1150_U86;
  assign new_P1_R1150_U302 = ~new_P1_U3054 | ~new_P1_R1150_U84;
  assign new_P1_R1150_U303 = ~new_P1_R1150_U301 | ~new_P1_R1150_U302;
  assign new_P1_R1150_U304 = ~new_P1_U3974 | ~new_P1_R1150_U85;
  assign new_P1_R1150_U305 = ~new_P1_U3974 | ~new_P1_R1150_U85;
  assign new_P1_R1150_U306 = ~new_P1_R1150_U305 | ~new_P1_R1150_U86;
  assign new_P1_R1150_U307 = ~new_P1_U3054 | ~new_P1_R1150_U84;
  assign new_P1_R1150_U308 = ~new_P1_R1150_U153 | ~new_P1_R1150_U307 | ~new_P1_R1150_U306;
  assign new_P1_R1150_U309 = ~new_P1_R1150_U295 | ~new_P1_R1150_U82;
  assign new_P1_R1150_U310 = ~new_P1_R1150_U129 | ~new_P1_R1150_U309;
  assign new_P1_R1150_U311 = ~new_P1_R1150_U87 | ~new_P1_R1150_U177;
  assign new_P1_R1150_U312 = ~new_P1_R1150_U128 | ~new_P1_R1150_U311;
  assign new_P1_R1150_U313 = ~new_P1_R1150_U82 | ~new_P1_R1150_U177;
  assign new_P1_R1150_U314 = ~new_P1_R1150_U283 | ~new_P1_R1150_U159;
  assign new_P1_R1150_U315 = ~new_P1_R1150_U88;
  assign new_P1_R1150_U316 = ~new_P1_U3061 | ~new_P1_R1150_U45;
  assign new_P1_R1150_U317 = ~new_P1_R1150_U315 | ~new_P1_R1150_U316;
  assign new_P1_R1150_U318 = ~new_P1_R1150_U132 | ~new_P1_R1150_U317;
  assign new_P1_R1150_U319 = ~new_P1_R1150_U88 | ~new_P1_R1150_U176;
  assign new_P1_R1150_U320 = ~new_P1_U3979 | ~new_P1_R1150_U72;
  assign new_P1_R1150_U321 = ~new_P1_R1150_U9 | ~new_P1_R1150_U320 | ~new_P1_R1150_U319;
  assign new_P1_R1150_U322 = ~new_P1_U3061 | ~new_P1_R1150_U45;
  assign new_P1_R1150_U323 = ~new_P1_R1150_U176 | ~new_P1_R1150_U322;
  assign new_P1_R1150_U324 = ~new_P1_R1150_U283 | ~new_P1_R1150_U75;
  assign new_P1_R1150_U325 = ~new_P1_R1150_U257 | ~new_P1_R1150_U167;
  assign new_P1_R1150_U326 = ~new_P1_R1150_U89;
  assign new_P1_R1150_U327 = ~new_P1_U3074 | ~new_P1_R1150_U46;
  assign new_P1_R1150_U328 = ~new_P1_R1150_U326 | ~new_P1_R1150_U327;
  assign new_P1_R1150_U329 = ~new_P1_R1150_U139 | ~new_P1_R1150_U328;
  assign new_P1_R1150_U330 = ~new_P1_R1150_U89 | ~new_P1_R1150_U175;
  assign new_P1_R1150_U331 = ~new_P1_U3500 | ~new_P1_R1150_U58;
  assign new_P1_R1150_U332 = ~new_P1_R1150_U138 | ~new_P1_R1150_U330;
  assign new_P1_R1150_U333 = ~new_P1_U3074 | ~new_P1_R1150_U46;
  assign new_P1_R1150_U334 = ~new_P1_R1150_U175 | ~new_P1_R1150_U333;
  assign new_P1_R1150_U335 = ~new_P1_R1150_U257 | ~new_P1_R1150_U61;
  assign new_P1_R1150_U336 = ~new_P1_R1150_U212 | ~new_P1_R1150_U145;
  assign new_P1_R1150_U337 = ~new_P1_R1150_U90;
  assign new_P1_R1150_U338 = ~new_P1_U3062 | ~new_P1_R1150_U47;
  assign new_P1_R1150_U339 = ~new_P1_R1150_U337 | ~new_P1_R1150_U338;
  assign new_P1_R1150_U340 = ~new_P1_R1150_U143 | ~new_P1_R1150_U339;
  assign new_P1_R1150_U341 = ~new_P1_R1150_U90 | ~new_P1_R1150_U174;
  assign new_P1_R1150_U342 = ~new_P1_U3485 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U343 = ~new_P1_R1150_U142 | ~new_P1_R1150_U341;
  assign new_P1_R1150_U344 = ~new_P1_U3062 | ~new_P1_R1150_U47;
  assign new_P1_R1150_U345 = ~new_P1_R1150_U174 | ~new_P1_R1150_U344;
  assign new_P1_R1150_U346 = ~new_P1_U3077 | ~new_P1_R1150_U22;
  assign new_P1_R1150_U347 = ~new_P1_R1150_U385 | ~new_P1_R1150_U304 | ~new_P1_R1150_U303;
  assign new_P1_R1150_U348 = ~new_P1_U3479 | ~new_P1_R1150_U40;
  assign new_P1_R1150_U349 = ~new_P1_U3083 | ~new_P1_R1150_U39;
  assign new_P1_R1150_U350 = ~new_P1_R1150_U213 | ~new_P1_R1150_U145;
  assign new_P1_R1150_U351 = ~new_P1_R1150_U211 | ~new_P1_R1150_U144;
  assign new_P1_R1150_U352 = ~new_P1_U3476 | ~new_P1_R1150_U38;
  assign new_P1_R1150_U353 = ~new_P1_U3084 | ~new_P1_R1150_U35;
  assign new_P1_R1150_U354 = ~new_P1_U3476 | ~new_P1_R1150_U38;
  assign new_P1_R1150_U355 = ~new_P1_U3084 | ~new_P1_R1150_U35;
  assign new_P1_R1150_U356 = ~new_P1_R1150_U355 | ~new_P1_R1150_U354;
  assign new_P1_R1150_U357 = ~new_P1_U3473 | ~new_P1_R1150_U36;
  assign new_P1_R1150_U358 = ~new_P1_U3070 | ~new_P1_R1150_U19;
  assign new_P1_R1150_U359 = ~new_P1_R1150_U218 | ~new_P1_R1150_U41;
  assign new_P1_R1150_U360 = ~new_P1_R1150_U146 | ~new_P1_R1150_U205;
  assign new_P1_R1150_U361 = ~new_P1_U3470 | ~new_P1_R1150_U31;
  assign new_P1_R1150_U362 = ~new_P1_U3071 | ~new_P1_R1150_U29;
  assign new_P1_R1150_U363 = ~new_P1_R1150_U362 | ~new_P1_R1150_U361;
  assign new_P1_R1150_U364 = ~new_P1_U3467 | ~new_P1_R1150_U32;
  assign new_P1_R1150_U365 = ~new_P1_U3067 | ~new_P1_R1150_U20;
  assign new_P1_R1150_U366 = ~new_P1_R1150_U228 | ~new_P1_R1150_U42;
  assign new_P1_R1150_U367 = ~new_P1_R1150_U147 | ~new_P1_R1150_U220;
  assign new_P1_R1150_U368 = ~new_P1_U3464 | ~new_P1_R1150_U33;
  assign new_P1_R1150_U369 = ~new_P1_U3060 | ~new_P1_R1150_U30;
  assign new_P1_R1150_U370 = ~new_P1_R1150_U229 | ~new_P1_R1150_U149;
  assign new_P1_R1150_U371 = ~new_P1_R1150_U195 | ~new_P1_R1150_U148;
  assign new_P1_R1150_U372 = ~new_P1_U3461 | ~new_P1_R1150_U28;
  assign new_P1_R1150_U373 = ~new_P1_U3064 | ~new_P1_R1150_U25;
  assign new_P1_R1150_U374 = ~new_P1_U3461 | ~new_P1_R1150_U28;
  assign new_P1_R1150_U375 = ~new_P1_U3064 | ~new_P1_R1150_U25;
  assign new_P1_R1150_U376 = ~new_P1_R1150_U375 | ~new_P1_R1150_U374;
  assign new_P1_R1150_U377 = ~new_P1_U3458 | ~new_P1_R1150_U26;
  assign new_P1_R1150_U378 = ~new_P1_U3068 | ~new_P1_R1150_U21;
  assign new_P1_R1150_U379 = ~new_P1_R1150_U234 | ~new_P1_R1150_U43;
  assign new_P1_R1150_U380 = ~new_P1_R1150_U150 | ~new_P1_R1150_U189;
  assign new_P1_R1150_U381 = ~new_P1_U3985 | ~new_P1_R1150_U152;
  assign new_P1_R1150_U382 = ~new_P1_U3055 | ~new_P1_R1150_U151;
  assign new_P1_R1150_U383 = ~new_P1_U3985 | ~new_P1_R1150_U152;
  assign new_P1_R1150_U384 = ~new_P1_U3055 | ~new_P1_R1150_U151;
  assign new_P1_R1150_U385 = ~new_P1_R1150_U384 | ~new_P1_R1150_U383;
  assign new_P1_R1150_U386 = ~new_P1_U3974 | ~new_P1_R1150_U85;
  assign new_P1_R1150_U387 = ~new_P1_U3054 | ~new_P1_R1150_U84;
  assign new_P1_R1150_U388 = ~new_P1_R1150_U127;
  assign new_P1_R1150_U389 = ~new_P1_R1150_U388 | ~new_P1_R1150_U301;
  assign new_P1_R1150_U390 = ~new_P1_R1150_U127 | ~new_P1_R1150_U86;
  assign new_P1_R1150_U391 = ~new_P1_U3975 | ~new_P1_R1150_U83;
  assign new_P1_R1150_U392 = ~new_P1_U3053 | ~new_P1_R1150_U80;
  assign new_P1_R1150_U393 = ~new_P1_U3975 | ~new_P1_R1150_U83;
  assign new_P1_R1150_U394 = ~new_P1_U3053 | ~new_P1_R1150_U80;
  assign new_P1_R1150_U395 = ~new_P1_R1150_U394 | ~new_P1_R1150_U393;
  assign new_P1_R1150_U396 = ~new_P1_U3976 | ~new_P1_R1150_U81;
  assign new_P1_R1150_U397 = ~new_P1_U3057 | ~new_P1_R1150_U44;
  assign new_P1_R1150_U398 = ~new_P1_R1150_U313 | ~new_P1_R1150_U87;
  assign new_P1_R1150_U399 = ~new_P1_R1150_U154 | ~new_P1_R1150_U295;
  assign new_P1_R1150_U400 = ~new_P1_U3977 | ~new_P1_R1150_U79;
  assign new_P1_R1150_U401 = ~new_P1_U3058 | ~new_P1_R1150_U78;
  assign new_P1_R1150_U402 = ~new_P1_R1150_U130;
  assign new_P1_R1150_U403 = ~new_P1_R1150_U291 | ~new_P1_R1150_U402;
  assign new_P1_R1150_U404 = ~new_P1_R1150_U130 | ~new_P1_R1150_U155;
  assign new_P1_R1150_U405 = ~new_P1_U3978 | ~new_P1_R1150_U77;
  assign new_P1_R1150_U406 = ~new_P1_U3065 | ~new_P1_R1150_U76;
  assign new_P1_R1150_U407 = ~new_P1_R1150_U131;
  assign new_P1_R1150_U408 = ~new_P1_R1150_U287 | ~new_P1_R1150_U407;
  assign new_P1_R1150_U409 = ~new_P1_R1150_U131 | ~new_P1_R1150_U156;
  assign new_P1_R1150_U410 = ~new_P1_U3979 | ~new_P1_R1150_U72;
  assign new_P1_R1150_U411 = ~new_P1_U3066 | ~new_P1_R1150_U70;
  assign new_P1_R1150_U412 = ~new_P1_R1150_U411 | ~new_P1_R1150_U410;
  assign new_P1_R1150_U413 = ~new_P1_U3980 | ~new_P1_R1150_U73;
  assign new_P1_R1150_U414 = ~new_P1_U3061 | ~new_P1_R1150_U45;
  assign new_P1_R1150_U415 = ~new_P1_R1150_U323 | ~new_P1_R1150_U88;
  assign new_P1_R1150_U416 = ~new_P1_R1150_U157 | ~new_P1_R1150_U315;
  assign new_P1_R1150_U417 = ~new_P1_U3981 | ~new_P1_R1150_U74;
  assign new_P1_R1150_U418 = ~new_P1_U3075 | ~new_P1_R1150_U71;
  assign new_P1_R1150_U419 = ~new_P1_R1150_U324 | ~new_P1_R1150_U159;
  assign new_P1_R1150_U420 = ~new_P1_R1150_U277 | ~new_P1_R1150_U158;
  assign new_P1_R1150_U421 = ~new_P1_U3982 | ~new_P1_R1150_U69;
  assign new_P1_R1150_U422 = ~new_P1_U3076 | ~new_P1_R1150_U68;
  assign new_P1_R1150_U423 = ~new_P1_R1150_U133;
  assign new_P1_R1150_U424 = ~new_P1_R1150_U273 | ~new_P1_R1150_U423;
  assign new_P1_R1150_U425 = ~new_P1_R1150_U133 | ~new_P1_R1150_U160;
  assign new_P1_R1150_U426 = ~new_P1_R1150_U185 | ~new_P1_R1150_U24;
  assign new_P1_R1150_U427 = ~new_P1_U3078 | ~new_P1_R1150_U23;
  assign new_P1_R1150_U428 = ~new_P1_R1150_U134;
  assign new_P1_R1150_U429 = ~new_P1_U3455 | ~new_P1_R1150_U428;
  assign new_P1_R1150_U430 = ~new_P1_R1150_U134 | ~new_P1_R1150_U161;
  assign new_P1_R1150_U431 = ~new_P1_U3508 | ~new_P1_R1150_U67;
  assign new_P1_R1150_U432 = ~new_P1_U3081 | ~new_P1_R1150_U66;
  assign new_P1_R1150_U433 = ~new_P1_R1150_U135;
  assign new_P1_R1150_U434 = ~new_P1_R1150_U269 | ~new_P1_R1150_U433;
  assign new_P1_R1150_U435 = ~new_P1_R1150_U135 | ~new_P1_R1150_U162;
  assign new_P1_R1150_U436 = ~new_P1_U3506 | ~new_P1_R1150_U65;
  assign new_P1_R1150_U437 = ~new_P1_U3082 | ~new_P1_R1150_U163;
  assign new_P1_R1150_U438 = ~new_P1_R1150_U136;
  assign new_P1_R1150_U439 = ~new_P1_R1150_U438 | ~new_P1_R1150_U265;
  assign new_P1_R1150_U440 = ~new_P1_R1150_U136 | ~new_P1_R1150_U64;
  assign new_P1_R1150_U441 = ~new_P1_U3503 | ~new_P1_R1150_U63;
  assign new_P1_R1150_U442 = ~new_P1_U3069 | ~new_P1_R1150_U62;
  assign new_P1_R1150_U443 = ~new_P1_R1150_U137;
  assign new_P1_R1150_U444 = ~new_P1_R1150_U261 | ~new_P1_R1150_U443;
  assign new_P1_R1150_U445 = ~new_P1_R1150_U137 | ~new_P1_R1150_U164;
  assign new_P1_R1150_U446 = ~new_P1_U3500 | ~new_P1_R1150_U58;
  assign new_P1_R1150_U447 = ~new_P1_U3073 | ~new_P1_R1150_U56;
  assign new_P1_R1150_U448 = ~new_P1_R1150_U447 | ~new_P1_R1150_U446;
  assign new_P1_R1150_U449 = ~new_P1_U3497 | ~new_P1_R1150_U59;
  assign new_P1_R1150_U450 = ~new_P1_U3074 | ~new_P1_R1150_U46;
  assign new_P1_R1150_U451 = ~new_P1_R1150_U334 | ~new_P1_R1150_U89;
  assign new_P1_R1150_U452 = ~new_P1_R1150_U165 | ~new_P1_R1150_U326;
  assign new_P1_R1150_U453 = ~new_P1_U3494 | ~new_P1_R1150_U60;
  assign new_P1_R1150_U454 = ~new_P1_U3079 | ~new_P1_R1150_U57;
  assign new_P1_R1150_U455 = ~new_P1_R1150_U335 | ~new_P1_R1150_U167;
  assign new_P1_R1150_U456 = ~new_P1_R1150_U251 | ~new_P1_R1150_U166;
  assign new_P1_R1150_U457 = ~new_P1_U3491 | ~new_P1_R1150_U55;
  assign new_P1_R1150_U458 = ~new_P1_U3080 | ~new_P1_R1150_U54;
  assign new_P1_R1150_U459 = ~new_P1_R1150_U140;
  assign new_P1_R1150_U460 = ~new_P1_R1150_U247 | ~new_P1_R1150_U459;
  assign new_P1_R1150_U461 = ~new_P1_R1150_U140 | ~new_P1_R1150_U168;
  assign new_P1_R1150_U462 = ~new_P1_U3488 | ~new_P1_R1150_U53;
  assign new_P1_R1150_U463 = ~new_P1_U3072 | ~new_P1_R1150_U52;
  assign new_P1_R1150_U464 = ~new_P1_R1150_U141;
  assign new_P1_R1150_U465 = ~new_P1_R1150_U243 | ~new_P1_R1150_U464;
  assign new_P1_R1150_U466 = ~new_P1_R1150_U141 | ~new_P1_R1150_U169;
  assign new_P1_R1150_U467 = ~new_P1_U3485 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U468 = ~new_P1_U3063 | ~new_P1_R1150_U48;
  assign new_P1_R1150_U469 = ~new_P1_R1150_U468 | ~new_P1_R1150_U467;
  assign new_P1_R1150_U470 = ~new_P1_U3482 | ~new_P1_R1150_U50;
  assign new_P1_R1150_U471 = ~new_P1_U3062 | ~new_P1_R1150_U47;
  assign new_P1_R1150_U472 = ~new_P1_R1150_U345 | ~new_P1_R1150_U90;
  assign new_P1_R1150_U473 = ~new_P1_R1150_U170 | ~new_P1_R1150_U337;
  assign new_P1_R1192_U6 = new_P1_R1192_U198 & new_P1_R1192_U197;
  assign new_P1_R1192_U7 = new_P1_R1192_U237 & new_P1_R1192_U236;
  assign new_P1_R1192_U8 = new_P1_R1192_U254 & new_P1_R1192_U253;
  assign new_P1_R1192_U9 = new_P1_R1192_U280 & new_P1_R1192_U279;
  assign new_P1_R1192_U10 = ~new_P1_R1192_U340 | ~new_P1_R1192_U343;
  assign new_P1_R1192_U11 = ~new_P1_R1192_U329 | ~new_P1_R1192_U332;
  assign new_P1_R1192_U12 = ~new_P1_R1192_U318 | ~new_P1_R1192_U321;
  assign new_P1_R1192_U13 = ~new_P1_R1192_U310 | ~new_P1_R1192_U312;
  assign new_P1_R1192_U14 = ~new_P1_R1192_U347 | ~new_P1_R1192_U308;
  assign new_P1_R1192_U15 = ~new_P1_R1192_U231 | ~new_P1_R1192_U233;
  assign new_P1_R1192_U16 = ~new_P1_R1192_U223 | ~new_P1_R1192_U226;
  assign new_P1_R1192_U17 = ~new_P1_R1192_U215 | ~new_P1_R1192_U217;
  assign new_P1_R1192_U18 = ~new_P1_R1192_U23 | ~new_P1_R1192_U346;
  assign new_P1_R1192_U19 = ~new_P1_U3473;
  assign new_P1_R1192_U20 = ~new_P1_U3467;
  assign new_P1_R1192_U21 = ~new_P1_U3458;
  assign new_P1_R1192_U22 = ~new_P1_U3450;
  assign new_P1_R1192_U23 = ~new_P1_U3450 | ~new_P1_R1192_U91;
  assign new_P1_R1192_U24 = ~new_P1_U3078;
  assign new_P1_R1192_U25 = ~new_P1_U3461;
  assign new_P1_R1192_U26 = ~new_P1_U3068;
  assign new_P1_R1192_U27 = ~new_P1_U3068 | ~new_P1_R1192_U21;
  assign new_P1_R1192_U28 = ~new_P1_U3064;
  assign new_P1_R1192_U29 = ~new_P1_U3470;
  assign new_P1_R1192_U30 = ~new_P1_U3464;
  assign new_P1_R1192_U31 = ~new_P1_U3071;
  assign new_P1_R1192_U32 = ~new_P1_U3067;
  assign new_P1_R1192_U33 = ~new_P1_U3060;
  assign new_P1_R1192_U34 = ~new_P1_U3060 | ~new_P1_R1192_U30;
  assign new_P1_R1192_U35 = ~new_P1_U3476;
  assign new_P1_R1192_U36 = ~new_P1_U3070;
  assign new_P1_R1192_U37 = ~new_P1_U3070 | ~new_P1_R1192_U19;
  assign new_P1_R1192_U38 = ~new_P1_U3084;
  assign new_P1_R1192_U39 = ~new_P1_U3479;
  assign new_P1_R1192_U40 = ~new_P1_U3083;
  assign new_P1_R1192_U41 = ~new_P1_R1192_U204 | ~new_P1_R1192_U203;
  assign new_P1_R1192_U42 = ~new_P1_R1192_U34 | ~new_P1_R1192_U219;
  assign new_P1_R1192_U43 = ~new_P1_R1192_U188 | ~new_P1_R1192_U187;
  assign new_P1_R1192_U44 = ~new_P1_U3976;
  assign new_P1_R1192_U45 = ~new_P1_U3980;
  assign new_P1_R1192_U46 = ~new_P1_U3497;
  assign new_P1_R1192_U47 = ~new_P1_U3482;
  assign new_P1_R1192_U48 = ~new_P1_U3485;
  assign new_P1_R1192_U49 = ~new_P1_U3063;
  assign new_P1_R1192_U50 = ~new_P1_U3062;
  assign new_P1_R1192_U51 = ~new_P1_U3083 | ~new_P1_R1192_U39;
  assign new_P1_R1192_U52 = ~new_P1_U3488;
  assign new_P1_R1192_U53 = ~new_P1_U3072;
  assign new_P1_R1192_U54 = ~new_P1_U3491;
  assign new_P1_R1192_U55 = ~new_P1_U3080;
  assign new_P1_R1192_U56 = ~new_P1_U3500;
  assign new_P1_R1192_U57 = ~new_P1_U3494;
  assign new_P1_R1192_U58 = ~new_P1_U3073;
  assign new_P1_R1192_U59 = ~new_P1_U3074;
  assign new_P1_R1192_U60 = ~new_P1_U3079;
  assign new_P1_R1192_U61 = ~new_P1_U3079 | ~new_P1_R1192_U57;
  assign new_P1_R1192_U62 = ~new_P1_U3503;
  assign new_P1_R1192_U63 = ~new_P1_U3069;
  assign new_P1_R1192_U64 = ~new_P1_R1192_U264 | ~new_P1_R1192_U263;
  assign new_P1_R1192_U65 = ~new_P1_U3082;
  assign new_P1_R1192_U66 = ~new_P1_U3508;
  assign new_P1_R1192_U67 = ~new_P1_U3081;
  assign new_P1_R1192_U68 = ~new_P1_U3982;
  assign new_P1_R1192_U69 = ~new_P1_U3076;
  assign new_P1_R1192_U70 = ~new_P1_U3979;
  assign new_P1_R1192_U71 = ~new_P1_U3981;
  assign new_P1_R1192_U72 = ~new_P1_U3066;
  assign new_P1_R1192_U73 = ~new_P1_U3061;
  assign new_P1_R1192_U74 = ~new_P1_U3075;
  assign new_P1_R1192_U75 = ~new_P1_U3075 | ~new_P1_R1192_U71;
  assign new_P1_R1192_U76 = ~new_P1_U3978;
  assign new_P1_R1192_U77 = ~new_P1_U3065;
  assign new_P1_R1192_U78 = ~new_P1_U3977;
  assign new_P1_R1192_U79 = ~new_P1_U3058;
  assign new_P1_R1192_U80 = ~new_P1_U3975;
  assign new_P1_R1192_U81 = ~new_P1_U3057;
  assign new_P1_R1192_U82 = ~new_P1_U3057 | ~new_P1_R1192_U44;
  assign new_P1_R1192_U83 = ~new_P1_U3053;
  assign new_P1_R1192_U84 = ~new_P1_U3974;
  assign new_P1_R1192_U85 = ~new_P1_U3054;
  assign new_P1_R1192_U86 = ~new_P1_R1192_U126 | ~new_P1_R1192_U297;
  assign new_P1_R1192_U87 = ~new_P1_R1192_U294 | ~new_P1_R1192_U293;
  assign new_P1_R1192_U88 = ~new_P1_R1192_U75 | ~new_P1_R1192_U314;
  assign new_P1_R1192_U89 = ~new_P1_R1192_U61 | ~new_P1_R1192_U325;
  assign new_P1_R1192_U90 = ~new_P1_R1192_U51 | ~new_P1_R1192_U336;
  assign new_P1_R1192_U91 = ~new_P1_U3077;
  assign new_P1_R1192_U92 = ~new_P1_R1192_U390 | ~new_P1_R1192_U389;
  assign new_P1_R1192_U93 = ~new_P1_R1192_U404 | ~new_P1_R1192_U403;
  assign new_P1_R1192_U94 = ~new_P1_R1192_U409 | ~new_P1_R1192_U408;
  assign new_P1_R1192_U95 = ~new_P1_R1192_U425 | ~new_P1_R1192_U424;
  assign new_P1_R1192_U96 = ~new_P1_R1192_U430 | ~new_P1_R1192_U429;
  assign new_P1_R1192_U97 = ~new_P1_R1192_U435 | ~new_P1_R1192_U434;
  assign new_P1_R1192_U98 = ~new_P1_R1192_U440 | ~new_P1_R1192_U439;
  assign new_P1_R1192_U99 = ~new_P1_R1192_U445 | ~new_P1_R1192_U444;
  assign new_P1_R1192_U100 = ~new_P1_R1192_U461 | ~new_P1_R1192_U460;
  assign new_P1_R1192_U101 = ~new_P1_R1192_U466 | ~new_P1_R1192_U465;
  assign new_P1_R1192_U102 = ~new_P1_R1192_U351 | ~new_P1_R1192_U350;
  assign new_P1_R1192_U103 = ~new_P1_R1192_U360 | ~new_P1_R1192_U359;
  assign new_P1_R1192_U104 = ~new_P1_R1192_U367 | ~new_P1_R1192_U366;
  assign new_P1_R1192_U105 = ~new_P1_R1192_U371 | ~new_P1_R1192_U370;
  assign new_P1_R1192_U106 = ~new_P1_R1192_U380 | ~new_P1_R1192_U379;
  assign new_P1_R1192_U107 = ~new_P1_R1192_U399 | ~new_P1_R1192_U398;
  assign new_P1_R1192_U108 = ~new_P1_R1192_U416 | ~new_P1_R1192_U415;
  assign new_P1_R1192_U109 = ~new_P1_R1192_U420 | ~new_P1_R1192_U419;
  assign new_P1_R1192_U110 = ~new_P1_R1192_U452 | ~new_P1_R1192_U451;
  assign new_P1_R1192_U111 = ~new_P1_R1192_U456 | ~new_P1_R1192_U455;
  assign new_P1_R1192_U112 = ~new_P1_R1192_U473 | ~new_P1_R1192_U472;
  assign new_P1_R1192_U113 = new_P1_R1192_U193 & new_P1_R1192_U194;
  assign new_P1_R1192_U114 = new_P1_R1192_U201 & new_P1_R1192_U196;
  assign new_P1_R1192_U115 = new_P1_R1192_U206 & new_P1_R1192_U180;
  assign new_P1_R1192_U116 = new_P1_R1192_U209 & new_P1_R1192_U210;
  assign new_P1_R1192_U117 = new_P1_R1192_U37 & new_P1_R1192_U353 & new_P1_R1192_U352;
  assign new_P1_R1192_U118 = new_P1_R1192_U356 & new_P1_R1192_U180;
  assign new_P1_R1192_U119 = new_P1_R1192_U225 & new_P1_R1192_U6;
  assign new_P1_R1192_U120 = new_P1_R1192_U363 & new_P1_R1192_U179;
  assign new_P1_R1192_U121 = new_P1_R1192_U27 & new_P1_R1192_U373 & new_P1_R1192_U372;
  assign new_P1_R1192_U122 = new_P1_R1192_U376 & new_P1_R1192_U178;
  assign new_P1_R1192_U123 = new_P1_R1192_U174 & new_P1_R1192_U235 & new_P1_R1192_U212;
  assign new_P1_R1192_U124 = new_P1_R1192_U252 & new_P1_R1192_U257 & new_P1_R1192_U175;
  assign new_P1_R1192_U125 = new_P1_R1192_U283 & new_P1_R1192_U176;
  assign new_P1_R1192_U126 = new_P1_R1192_U299 & new_P1_R1192_U300;
  assign new_P1_R1192_U127 = ~new_P1_R1192_U387 | ~new_P1_R1192_U386;
  assign new_P1_R1192_U128 = new_P1_R1192_U82 & new_P1_R1192_U392 & new_P1_R1192_U391;
  assign new_P1_R1192_U129 = new_P1_R1192_U395 & new_P1_R1192_U177;
  assign new_P1_R1192_U130 = ~new_P1_R1192_U401 | ~new_P1_R1192_U400;
  assign new_P1_R1192_U131 = ~new_P1_R1192_U406 | ~new_P1_R1192_U405;
  assign new_P1_R1192_U132 = new_P1_R1192_U412 & new_P1_R1192_U176;
  assign new_P1_R1192_U133 = ~new_P1_R1192_U422 | ~new_P1_R1192_U421;
  assign new_P1_R1192_U134 = ~new_P1_R1192_U427 | ~new_P1_R1192_U426;
  assign new_P1_R1192_U135 = ~new_P1_R1192_U432 | ~new_P1_R1192_U431;
  assign new_P1_R1192_U136 = ~new_P1_R1192_U437 | ~new_P1_R1192_U436;
  assign new_P1_R1192_U137 = ~new_P1_R1192_U442 | ~new_P1_R1192_U441;
  assign new_P1_R1192_U138 = new_P1_R1192_U331 & new_P1_R1192_U8;
  assign new_P1_R1192_U139 = new_P1_R1192_U448 & new_P1_R1192_U175;
  assign new_P1_R1192_U140 = ~new_P1_R1192_U458 | ~new_P1_R1192_U457;
  assign new_P1_R1192_U141 = ~new_P1_R1192_U463 | ~new_P1_R1192_U462;
  assign new_P1_R1192_U142 = new_P1_R1192_U342 & new_P1_R1192_U7;
  assign new_P1_R1192_U143 = new_P1_R1192_U469 & new_P1_R1192_U174;
  assign new_P1_R1192_U144 = new_P1_R1192_U349 & new_P1_R1192_U348;
  assign new_P1_R1192_U145 = ~new_P1_R1192_U116 | ~new_P1_R1192_U207;
  assign new_P1_R1192_U146 = new_P1_R1192_U358 & new_P1_R1192_U357;
  assign new_P1_R1192_U147 = new_P1_R1192_U365 & new_P1_R1192_U364;
  assign new_P1_R1192_U148 = new_P1_R1192_U369 & new_P1_R1192_U368;
  assign new_P1_R1192_U149 = ~new_P1_R1192_U113 | ~new_P1_R1192_U191;
  assign new_P1_R1192_U150 = new_P1_R1192_U378 & new_P1_R1192_U377;
  assign new_P1_R1192_U151 = ~new_P1_U3985;
  assign new_P1_R1192_U152 = ~new_P1_U3055;
  assign new_P1_R1192_U153 = new_P1_R1192_U382 & new_P1_R1192_U381;
  assign new_P1_R1192_U154 = new_P1_R1192_U397 & new_P1_R1192_U396;
  assign new_P1_R1192_U155 = ~new_P1_R1192_U290 | ~new_P1_R1192_U289;
  assign new_P1_R1192_U156 = ~new_P1_R1192_U286 | ~new_P1_R1192_U285;
  assign new_P1_R1192_U157 = new_P1_R1192_U414 & new_P1_R1192_U413;
  assign new_P1_R1192_U158 = new_P1_R1192_U418 & new_P1_R1192_U417;
  assign new_P1_R1192_U159 = ~new_P1_R1192_U276 | ~new_P1_R1192_U275;
  assign new_P1_R1192_U160 = ~new_P1_R1192_U272 | ~new_P1_R1192_U271;
  assign new_P1_R1192_U161 = ~new_P1_U3455;
  assign new_P1_R1192_U162 = ~new_P1_R1192_U268 | ~new_P1_R1192_U267;
  assign new_P1_R1192_U163 = ~new_P1_U3506;
  assign new_P1_R1192_U164 = ~new_P1_R1192_U260 | ~new_P1_R1192_U259;
  assign new_P1_R1192_U165 = new_P1_R1192_U450 & new_P1_R1192_U449;
  assign new_P1_R1192_U166 = new_P1_R1192_U454 & new_P1_R1192_U453;
  assign new_P1_R1192_U167 = ~new_P1_R1192_U250 | ~new_P1_R1192_U249;
  assign new_P1_R1192_U168 = ~new_P1_R1192_U246 | ~new_P1_R1192_U245;
  assign new_P1_R1192_U169 = ~new_P1_R1192_U242 | ~new_P1_R1192_U241;
  assign new_P1_R1192_U170 = new_P1_R1192_U471 & new_P1_R1192_U470;
  assign new_P1_R1192_U171 = ~new_P1_R1192_U82;
  assign new_P1_R1192_U172 = ~new_P1_R1192_U27;
  assign new_P1_R1192_U173 = ~new_P1_R1192_U37;
  assign new_P1_R1192_U174 = ~new_P1_U3482 | ~new_P1_R1192_U50;
  assign new_P1_R1192_U175 = ~new_P1_U3497 | ~new_P1_R1192_U59;
  assign new_P1_R1192_U176 = ~new_P1_U3980 | ~new_P1_R1192_U73;
  assign new_P1_R1192_U177 = ~new_P1_U3976 | ~new_P1_R1192_U81;
  assign new_P1_R1192_U178 = ~new_P1_U3458 | ~new_P1_R1192_U26;
  assign new_P1_R1192_U179 = ~new_P1_U3467 | ~new_P1_R1192_U32;
  assign new_P1_R1192_U180 = ~new_P1_U3473 | ~new_P1_R1192_U36;
  assign new_P1_R1192_U181 = ~new_P1_R1192_U61;
  assign new_P1_R1192_U182 = ~new_P1_R1192_U75;
  assign new_P1_R1192_U183 = ~new_P1_R1192_U34;
  assign new_P1_R1192_U184 = ~new_P1_R1192_U51;
  assign new_P1_R1192_U185 = ~new_P1_R1192_U23;
  assign new_P1_R1192_U186 = ~new_P1_R1192_U185 | ~new_P1_R1192_U24;
  assign new_P1_R1192_U187 = ~new_P1_R1192_U186 | ~new_P1_R1192_U161;
  assign new_P1_R1192_U188 = ~new_P1_U3078 | ~new_P1_R1192_U23;
  assign new_P1_R1192_U189 = ~new_P1_R1192_U43;
  assign new_P1_R1192_U190 = ~new_P1_U3461 | ~new_P1_R1192_U28;
  assign new_P1_R1192_U191 = ~new_P1_R1192_U190 | ~new_P1_R1192_U43 | ~new_P1_R1192_U178;
  assign new_P1_R1192_U192 = ~new_P1_R1192_U28 | ~new_P1_R1192_U27;
  assign new_P1_R1192_U193 = ~new_P1_R1192_U192 | ~new_P1_R1192_U25;
  assign new_P1_R1192_U194 = ~new_P1_U3064 | ~new_P1_R1192_U172;
  assign new_P1_R1192_U195 = ~new_P1_R1192_U149;
  assign new_P1_R1192_U196 = ~new_P1_U3470 | ~new_P1_R1192_U31;
  assign new_P1_R1192_U197 = ~new_P1_U3071 | ~new_P1_R1192_U29;
  assign new_P1_R1192_U198 = ~new_P1_U3067 | ~new_P1_R1192_U20;
  assign new_P1_R1192_U199 = ~new_P1_R1192_U183 | ~new_P1_R1192_U179;
  assign new_P1_R1192_U200 = ~new_P1_R1192_U6 | ~new_P1_R1192_U199;
  assign new_P1_R1192_U201 = ~new_P1_U3464 | ~new_P1_R1192_U33;
  assign new_P1_R1192_U202 = ~new_P1_U3470 | ~new_P1_R1192_U31;
  assign new_P1_R1192_U203 = ~new_P1_R1192_U114 | ~new_P1_R1192_U149 | ~new_P1_R1192_U179;
  assign new_P1_R1192_U204 = ~new_P1_R1192_U202 | ~new_P1_R1192_U200;
  assign new_P1_R1192_U205 = ~new_P1_R1192_U41;
  assign new_P1_R1192_U206 = ~new_P1_U3476 | ~new_P1_R1192_U38;
  assign new_P1_R1192_U207 = ~new_P1_R1192_U115 | ~new_P1_R1192_U41;
  assign new_P1_R1192_U208 = ~new_P1_R1192_U38 | ~new_P1_R1192_U37;
  assign new_P1_R1192_U209 = ~new_P1_R1192_U208 | ~new_P1_R1192_U35;
  assign new_P1_R1192_U210 = ~new_P1_U3084 | ~new_P1_R1192_U173;
  assign new_P1_R1192_U211 = ~new_P1_R1192_U145;
  assign new_P1_R1192_U212 = ~new_P1_U3479 | ~new_P1_R1192_U40;
  assign new_P1_R1192_U213 = ~new_P1_R1192_U212 | ~new_P1_R1192_U51;
  assign new_P1_R1192_U214 = ~new_P1_R1192_U205 | ~new_P1_R1192_U37;
  assign new_P1_R1192_U215 = ~new_P1_R1192_U118 | ~new_P1_R1192_U214;
  assign new_P1_R1192_U216 = ~new_P1_R1192_U41 | ~new_P1_R1192_U180;
  assign new_P1_R1192_U217 = ~new_P1_R1192_U117 | ~new_P1_R1192_U216;
  assign new_P1_R1192_U218 = ~new_P1_R1192_U37 | ~new_P1_R1192_U180;
  assign new_P1_R1192_U219 = ~new_P1_R1192_U201 | ~new_P1_R1192_U149;
  assign new_P1_R1192_U220 = ~new_P1_R1192_U42;
  assign new_P1_R1192_U221 = ~new_P1_U3067 | ~new_P1_R1192_U20;
  assign new_P1_R1192_U222 = ~new_P1_R1192_U220 | ~new_P1_R1192_U221;
  assign new_P1_R1192_U223 = ~new_P1_R1192_U120 | ~new_P1_R1192_U222;
  assign new_P1_R1192_U224 = ~new_P1_R1192_U42 | ~new_P1_R1192_U179;
  assign new_P1_R1192_U225 = ~new_P1_U3470 | ~new_P1_R1192_U31;
  assign new_P1_R1192_U226 = ~new_P1_R1192_U119 | ~new_P1_R1192_U224;
  assign new_P1_R1192_U227 = ~new_P1_U3067 | ~new_P1_R1192_U20;
  assign new_P1_R1192_U228 = ~new_P1_R1192_U179 | ~new_P1_R1192_U227;
  assign new_P1_R1192_U229 = ~new_P1_R1192_U201 | ~new_P1_R1192_U34;
  assign new_P1_R1192_U230 = ~new_P1_R1192_U189 | ~new_P1_R1192_U27;
  assign new_P1_R1192_U231 = ~new_P1_R1192_U122 | ~new_P1_R1192_U230;
  assign new_P1_R1192_U232 = ~new_P1_R1192_U43 | ~new_P1_R1192_U178;
  assign new_P1_R1192_U233 = ~new_P1_R1192_U121 | ~new_P1_R1192_U232;
  assign new_P1_R1192_U234 = ~new_P1_R1192_U27 | ~new_P1_R1192_U178;
  assign new_P1_R1192_U235 = ~new_P1_U3485 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U236 = ~new_P1_U3063 | ~new_P1_R1192_U48;
  assign new_P1_R1192_U237 = ~new_P1_U3062 | ~new_P1_R1192_U47;
  assign new_P1_R1192_U238 = ~new_P1_R1192_U184 | ~new_P1_R1192_U174;
  assign new_P1_R1192_U239 = ~new_P1_R1192_U7 | ~new_P1_R1192_U238;
  assign new_P1_R1192_U240 = ~new_P1_U3485 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U241 = ~new_P1_R1192_U145 | ~new_P1_R1192_U123;
  assign new_P1_R1192_U242 = ~new_P1_R1192_U240 | ~new_P1_R1192_U239;
  assign new_P1_R1192_U243 = ~new_P1_R1192_U169;
  assign new_P1_R1192_U244 = ~new_P1_U3488 | ~new_P1_R1192_U53;
  assign new_P1_R1192_U245 = ~new_P1_R1192_U244 | ~new_P1_R1192_U169;
  assign new_P1_R1192_U246 = ~new_P1_U3072 | ~new_P1_R1192_U52;
  assign new_P1_R1192_U247 = ~new_P1_R1192_U168;
  assign new_P1_R1192_U248 = ~new_P1_U3491 | ~new_P1_R1192_U55;
  assign new_P1_R1192_U249 = ~new_P1_R1192_U248 | ~new_P1_R1192_U168;
  assign new_P1_R1192_U250 = ~new_P1_U3080 | ~new_P1_R1192_U54;
  assign new_P1_R1192_U251 = ~new_P1_R1192_U167;
  assign new_P1_R1192_U252 = ~new_P1_U3500 | ~new_P1_R1192_U58;
  assign new_P1_R1192_U253 = ~new_P1_U3073 | ~new_P1_R1192_U56;
  assign new_P1_R1192_U254 = ~new_P1_U3074 | ~new_P1_R1192_U46;
  assign new_P1_R1192_U255 = ~new_P1_R1192_U181 | ~new_P1_R1192_U175;
  assign new_P1_R1192_U256 = ~new_P1_R1192_U8 | ~new_P1_R1192_U255;
  assign new_P1_R1192_U257 = ~new_P1_U3494 | ~new_P1_R1192_U60;
  assign new_P1_R1192_U258 = ~new_P1_U3500 | ~new_P1_R1192_U58;
  assign new_P1_R1192_U259 = ~new_P1_R1192_U167 | ~new_P1_R1192_U124;
  assign new_P1_R1192_U260 = ~new_P1_R1192_U258 | ~new_P1_R1192_U256;
  assign new_P1_R1192_U261 = ~new_P1_R1192_U164;
  assign new_P1_R1192_U262 = ~new_P1_U3503 | ~new_P1_R1192_U63;
  assign new_P1_R1192_U263 = ~new_P1_R1192_U262 | ~new_P1_R1192_U164;
  assign new_P1_R1192_U264 = ~new_P1_U3069 | ~new_P1_R1192_U62;
  assign new_P1_R1192_U265 = ~new_P1_R1192_U64;
  assign new_P1_R1192_U266 = ~new_P1_R1192_U265 | ~new_P1_R1192_U65;
  assign new_P1_R1192_U267 = ~new_P1_R1192_U266 | ~new_P1_R1192_U163;
  assign new_P1_R1192_U268 = ~new_P1_U3082 | ~new_P1_R1192_U64;
  assign new_P1_R1192_U269 = ~new_P1_R1192_U162;
  assign new_P1_R1192_U270 = ~new_P1_U3508 | ~new_P1_R1192_U67;
  assign new_P1_R1192_U271 = ~new_P1_R1192_U270 | ~new_P1_R1192_U162;
  assign new_P1_R1192_U272 = ~new_P1_U3081 | ~new_P1_R1192_U66;
  assign new_P1_R1192_U273 = ~new_P1_R1192_U160;
  assign new_P1_R1192_U274 = ~new_P1_U3982 | ~new_P1_R1192_U69;
  assign new_P1_R1192_U275 = ~new_P1_R1192_U274 | ~new_P1_R1192_U160;
  assign new_P1_R1192_U276 = ~new_P1_U3076 | ~new_P1_R1192_U68;
  assign new_P1_R1192_U277 = ~new_P1_R1192_U159;
  assign new_P1_R1192_U278 = ~new_P1_U3979 | ~new_P1_R1192_U72;
  assign new_P1_R1192_U279 = ~new_P1_U3066 | ~new_P1_R1192_U70;
  assign new_P1_R1192_U280 = ~new_P1_U3061 | ~new_P1_R1192_U45;
  assign new_P1_R1192_U281 = ~new_P1_R1192_U182 | ~new_P1_R1192_U176;
  assign new_P1_R1192_U282 = ~new_P1_R1192_U9 | ~new_P1_R1192_U281;
  assign new_P1_R1192_U283 = ~new_P1_U3981 | ~new_P1_R1192_U74;
  assign new_P1_R1192_U284 = ~new_P1_U3979 | ~new_P1_R1192_U72;
  assign new_P1_R1192_U285 = ~new_P1_R1192_U278 | ~new_P1_R1192_U159 | ~new_P1_R1192_U125;
  assign new_P1_R1192_U286 = ~new_P1_R1192_U284 | ~new_P1_R1192_U282;
  assign new_P1_R1192_U287 = ~new_P1_R1192_U156;
  assign new_P1_R1192_U288 = ~new_P1_U3978 | ~new_P1_R1192_U77;
  assign new_P1_R1192_U289 = ~new_P1_R1192_U288 | ~new_P1_R1192_U156;
  assign new_P1_R1192_U290 = ~new_P1_U3065 | ~new_P1_R1192_U76;
  assign new_P1_R1192_U291 = ~new_P1_R1192_U155;
  assign new_P1_R1192_U292 = ~new_P1_U3977 | ~new_P1_R1192_U79;
  assign new_P1_R1192_U293 = ~new_P1_R1192_U292 | ~new_P1_R1192_U155;
  assign new_P1_R1192_U294 = ~new_P1_U3058 | ~new_P1_R1192_U78;
  assign new_P1_R1192_U295 = ~new_P1_R1192_U87;
  assign new_P1_R1192_U296 = ~new_P1_U3975 | ~new_P1_R1192_U83;
  assign new_P1_R1192_U297 = ~new_P1_R1192_U296 | ~new_P1_R1192_U87 | ~new_P1_R1192_U177;
  assign new_P1_R1192_U298 = ~new_P1_R1192_U83 | ~new_P1_R1192_U82;
  assign new_P1_R1192_U299 = ~new_P1_R1192_U298 | ~new_P1_R1192_U80;
  assign new_P1_R1192_U300 = ~new_P1_U3053 | ~new_P1_R1192_U171;
  assign new_P1_R1192_U301 = ~new_P1_R1192_U86;
  assign new_P1_R1192_U302 = ~new_P1_U3054 | ~new_P1_R1192_U84;
  assign new_P1_R1192_U303 = ~new_P1_R1192_U301 | ~new_P1_R1192_U302;
  assign new_P1_R1192_U304 = ~new_P1_U3974 | ~new_P1_R1192_U85;
  assign new_P1_R1192_U305 = ~new_P1_U3974 | ~new_P1_R1192_U85;
  assign new_P1_R1192_U306 = ~new_P1_R1192_U305 | ~new_P1_R1192_U86;
  assign new_P1_R1192_U307 = ~new_P1_U3054 | ~new_P1_R1192_U84;
  assign new_P1_R1192_U308 = ~new_P1_R1192_U153 | ~new_P1_R1192_U307 | ~new_P1_R1192_U306;
  assign new_P1_R1192_U309 = ~new_P1_R1192_U295 | ~new_P1_R1192_U82;
  assign new_P1_R1192_U310 = ~new_P1_R1192_U129 | ~new_P1_R1192_U309;
  assign new_P1_R1192_U311 = ~new_P1_R1192_U87 | ~new_P1_R1192_U177;
  assign new_P1_R1192_U312 = ~new_P1_R1192_U128 | ~new_P1_R1192_U311;
  assign new_P1_R1192_U313 = ~new_P1_R1192_U82 | ~new_P1_R1192_U177;
  assign new_P1_R1192_U314 = ~new_P1_R1192_U283 | ~new_P1_R1192_U159;
  assign new_P1_R1192_U315 = ~new_P1_R1192_U88;
  assign new_P1_R1192_U316 = ~new_P1_U3061 | ~new_P1_R1192_U45;
  assign new_P1_R1192_U317 = ~new_P1_R1192_U315 | ~new_P1_R1192_U316;
  assign new_P1_R1192_U318 = ~new_P1_R1192_U132 | ~new_P1_R1192_U317;
  assign new_P1_R1192_U319 = ~new_P1_R1192_U88 | ~new_P1_R1192_U176;
  assign new_P1_R1192_U320 = ~new_P1_U3979 | ~new_P1_R1192_U72;
  assign new_P1_R1192_U321 = ~new_P1_R1192_U9 | ~new_P1_R1192_U320 | ~new_P1_R1192_U319;
  assign new_P1_R1192_U322 = ~new_P1_U3061 | ~new_P1_R1192_U45;
  assign new_P1_R1192_U323 = ~new_P1_R1192_U176 | ~new_P1_R1192_U322;
  assign new_P1_R1192_U324 = ~new_P1_R1192_U283 | ~new_P1_R1192_U75;
  assign new_P1_R1192_U325 = ~new_P1_R1192_U257 | ~new_P1_R1192_U167;
  assign new_P1_R1192_U326 = ~new_P1_R1192_U89;
  assign new_P1_R1192_U327 = ~new_P1_U3074 | ~new_P1_R1192_U46;
  assign new_P1_R1192_U328 = ~new_P1_R1192_U326 | ~new_P1_R1192_U327;
  assign new_P1_R1192_U329 = ~new_P1_R1192_U139 | ~new_P1_R1192_U328;
  assign new_P1_R1192_U330 = ~new_P1_R1192_U89 | ~new_P1_R1192_U175;
  assign new_P1_R1192_U331 = ~new_P1_U3500 | ~new_P1_R1192_U58;
  assign new_P1_R1192_U332 = ~new_P1_R1192_U138 | ~new_P1_R1192_U330;
  assign new_P1_R1192_U333 = ~new_P1_U3074 | ~new_P1_R1192_U46;
  assign new_P1_R1192_U334 = ~new_P1_R1192_U175 | ~new_P1_R1192_U333;
  assign new_P1_R1192_U335 = ~new_P1_R1192_U257 | ~new_P1_R1192_U61;
  assign new_P1_R1192_U336 = ~new_P1_R1192_U212 | ~new_P1_R1192_U145;
  assign new_P1_R1192_U337 = ~new_P1_R1192_U90;
  assign new_P1_R1192_U338 = ~new_P1_U3062 | ~new_P1_R1192_U47;
  assign new_P1_R1192_U339 = ~new_P1_R1192_U337 | ~new_P1_R1192_U338;
  assign new_P1_R1192_U340 = ~new_P1_R1192_U143 | ~new_P1_R1192_U339;
  assign new_P1_R1192_U341 = ~new_P1_R1192_U90 | ~new_P1_R1192_U174;
  assign new_P1_R1192_U342 = ~new_P1_U3485 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U343 = ~new_P1_R1192_U142 | ~new_P1_R1192_U341;
  assign new_P1_R1192_U344 = ~new_P1_U3062 | ~new_P1_R1192_U47;
  assign new_P1_R1192_U345 = ~new_P1_R1192_U174 | ~new_P1_R1192_U344;
  assign new_P1_R1192_U346 = ~new_P1_U3077 | ~new_P1_R1192_U22;
  assign new_P1_R1192_U347 = ~new_P1_R1192_U385 | ~new_P1_R1192_U304 | ~new_P1_R1192_U303;
  assign new_P1_R1192_U348 = ~new_P1_U3479 | ~new_P1_R1192_U40;
  assign new_P1_R1192_U349 = ~new_P1_U3083 | ~new_P1_R1192_U39;
  assign new_P1_R1192_U350 = ~new_P1_R1192_U213 | ~new_P1_R1192_U145;
  assign new_P1_R1192_U351 = ~new_P1_R1192_U211 | ~new_P1_R1192_U144;
  assign new_P1_R1192_U352 = ~new_P1_U3476 | ~new_P1_R1192_U38;
  assign new_P1_R1192_U353 = ~new_P1_U3084 | ~new_P1_R1192_U35;
  assign new_P1_R1192_U354 = ~new_P1_U3476 | ~new_P1_R1192_U38;
  assign new_P1_R1192_U355 = ~new_P1_U3084 | ~new_P1_R1192_U35;
  assign new_P1_R1192_U356 = ~new_P1_R1192_U355 | ~new_P1_R1192_U354;
  assign new_P1_R1192_U357 = ~new_P1_U3473 | ~new_P1_R1192_U36;
  assign new_P1_R1192_U358 = ~new_P1_U3070 | ~new_P1_R1192_U19;
  assign new_P1_R1192_U359 = ~new_P1_R1192_U218 | ~new_P1_R1192_U41;
  assign new_P1_R1192_U360 = ~new_P1_R1192_U146 | ~new_P1_R1192_U205;
  assign new_P1_R1192_U361 = ~new_P1_U3470 | ~new_P1_R1192_U31;
  assign new_P1_R1192_U362 = ~new_P1_U3071 | ~new_P1_R1192_U29;
  assign new_P1_R1192_U363 = ~new_P1_R1192_U362 | ~new_P1_R1192_U361;
  assign new_P1_R1192_U364 = ~new_P1_U3467 | ~new_P1_R1192_U32;
  assign new_P1_R1192_U365 = ~new_P1_U3067 | ~new_P1_R1192_U20;
  assign new_P1_R1192_U366 = ~new_P1_R1192_U228 | ~new_P1_R1192_U42;
  assign new_P1_R1192_U367 = ~new_P1_R1192_U147 | ~new_P1_R1192_U220;
  assign new_P1_R1192_U368 = ~new_P1_U3464 | ~new_P1_R1192_U33;
  assign new_P1_R1192_U369 = ~new_P1_U3060 | ~new_P1_R1192_U30;
  assign new_P1_R1192_U370 = ~new_P1_R1192_U229 | ~new_P1_R1192_U149;
  assign new_P1_R1192_U371 = ~new_P1_R1192_U195 | ~new_P1_R1192_U148;
  assign new_P1_R1192_U372 = ~new_P1_U3461 | ~new_P1_R1192_U28;
  assign new_P1_R1192_U373 = ~new_P1_U3064 | ~new_P1_R1192_U25;
  assign new_P1_R1192_U374 = ~new_P1_U3461 | ~new_P1_R1192_U28;
  assign new_P1_R1192_U375 = ~new_P1_U3064 | ~new_P1_R1192_U25;
  assign new_P1_R1192_U376 = ~new_P1_R1192_U375 | ~new_P1_R1192_U374;
  assign new_P1_R1192_U377 = ~new_P1_U3458 | ~new_P1_R1192_U26;
  assign new_P1_R1192_U378 = ~new_P1_U3068 | ~new_P1_R1192_U21;
  assign new_P1_R1192_U379 = ~new_P1_R1192_U234 | ~new_P1_R1192_U43;
  assign new_P1_R1192_U380 = ~new_P1_R1192_U150 | ~new_P1_R1192_U189;
  assign new_P1_R1192_U381 = ~new_P1_U3985 | ~new_P1_R1192_U152;
  assign new_P1_R1192_U382 = ~new_P1_U3055 | ~new_P1_R1192_U151;
  assign new_P1_R1192_U383 = ~new_P1_U3985 | ~new_P1_R1192_U152;
  assign new_P1_R1192_U384 = ~new_P1_U3055 | ~new_P1_R1192_U151;
  assign new_P1_R1192_U385 = ~new_P1_R1192_U384 | ~new_P1_R1192_U383;
  assign new_P1_R1192_U386 = ~new_P1_U3974 | ~new_P1_R1192_U85;
  assign new_P1_R1192_U387 = ~new_P1_U3054 | ~new_P1_R1192_U84;
  assign new_P1_R1192_U388 = ~new_P1_R1192_U127;
  assign new_P1_R1192_U389 = ~new_P1_R1192_U388 | ~new_P1_R1192_U301;
  assign new_P1_R1192_U390 = ~new_P1_R1192_U127 | ~new_P1_R1192_U86;
  assign new_P1_R1192_U391 = ~new_P1_U3975 | ~new_P1_R1192_U83;
  assign new_P1_R1192_U392 = ~new_P1_U3053 | ~new_P1_R1192_U80;
  assign new_P1_R1192_U393 = ~new_P1_U3975 | ~new_P1_R1192_U83;
  assign new_P1_R1192_U394 = ~new_P1_U3053 | ~new_P1_R1192_U80;
  assign new_P1_R1192_U395 = ~new_P1_R1192_U394 | ~new_P1_R1192_U393;
  assign new_P1_R1192_U396 = ~new_P1_U3976 | ~new_P1_R1192_U81;
  assign new_P1_R1192_U397 = ~new_P1_U3057 | ~new_P1_R1192_U44;
  assign new_P1_R1192_U398 = ~new_P1_R1192_U313 | ~new_P1_R1192_U87;
  assign new_P1_R1192_U399 = ~new_P1_R1192_U154 | ~new_P1_R1192_U295;
  assign new_P1_R1192_U400 = ~new_P1_U3977 | ~new_P1_R1192_U79;
  assign new_P1_R1192_U401 = ~new_P1_U3058 | ~new_P1_R1192_U78;
  assign new_P1_R1192_U402 = ~new_P1_R1192_U130;
  assign new_P1_R1192_U403 = ~new_P1_R1192_U291 | ~new_P1_R1192_U402;
  assign new_P1_R1192_U404 = ~new_P1_R1192_U130 | ~new_P1_R1192_U155;
  assign new_P1_R1192_U405 = ~new_P1_U3978 | ~new_P1_R1192_U77;
  assign new_P1_R1192_U406 = ~new_P1_U3065 | ~new_P1_R1192_U76;
  assign new_P1_R1192_U407 = ~new_P1_R1192_U131;
  assign new_P1_R1192_U408 = ~new_P1_R1192_U287 | ~new_P1_R1192_U407;
  assign new_P1_R1192_U409 = ~new_P1_R1192_U131 | ~new_P1_R1192_U156;
  assign new_P1_R1192_U410 = ~new_P1_U3979 | ~new_P1_R1192_U72;
  assign new_P1_R1192_U411 = ~new_P1_U3066 | ~new_P1_R1192_U70;
  assign new_P1_R1192_U412 = ~new_P1_R1192_U411 | ~new_P1_R1192_U410;
  assign new_P1_R1192_U413 = ~new_P1_U3980 | ~new_P1_R1192_U73;
  assign new_P1_R1192_U414 = ~new_P1_U3061 | ~new_P1_R1192_U45;
  assign new_P1_R1192_U415 = ~new_P1_R1192_U323 | ~new_P1_R1192_U88;
  assign new_P1_R1192_U416 = ~new_P1_R1192_U157 | ~new_P1_R1192_U315;
  assign new_P1_R1192_U417 = ~new_P1_U3981 | ~new_P1_R1192_U74;
  assign new_P1_R1192_U418 = ~new_P1_U3075 | ~new_P1_R1192_U71;
  assign new_P1_R1192_U419 = ~new_P1_R1192_U324 | ~new_P1_R1192_U159;
  assign new_P1_R1192_U420 = ~new_P1_R1192_U277 | ~new_P1_R1192_U158;
  assign new_P1_R1192_U421 = ~new_P1_U3982 | ~new_P1_R1192_U69;
  assign new_P1_R1192_U422 = ~new_P1_U3076 | ~new_P1_R1192_U68;
  assign new_P1_R1192_U423 = ~new_P1_R1192_U133;
  assign new_P1_R1192_U424 = ~new_P1_R1192_U273 | ~new_P1_R1192_U423;
  assign new_P1_R1192_U425 = ~new_P1_R1192_U133 | ~new_P1_R1192_U160;
  assign new_P1_R1192_U426 = ~new_P1_R1192_U185 | ~new_P1_R1192_U24;
  assign new_P1_R1192_U427 = ~new_P1_U3078 | ~new_P1_R1192_U23;
  assign new_P1_R1192_U428 = ~new_P1_R1192_U134;
  assign new_P1_R1192_U429 = ~new_P1_U3455 | ~new_P1_R1192_U428;
  assign new_P1_R1192_U430 = ~new_P1_R1192_U134 | ~new_P1_R1192_U161;
  assign new_P1_R1192_U431 = ~new_P1_U3508 | ~new_P1_R1192_U67;
  assign new_P1_R1192_U432 = ~new_P1_U3081 | ~new_P1_R1192_U66;
  assign new_P1_R1192_U433 = ~new_P1_R1192_U135;
  assign new_P1_R1192_U434 = ~new_P1_R1192_U269 | ~new_P1_R1192_U433;
  assign new_P1_R1192_U435 = ~new_P1_R1192_U135 | ~new_P1_R1192_U162;
  assign new_P1_R1192_U436 = ~new_P1_U3506 | ~new_P1_R1192_U65;
  assign new_P1_R1192_U437 = ~new_P1_U3082 | ~new_P1_R1192_U163;
  assign new_P1_R1192_U438 = ~new_P1_R1192_U136;
  assign new_P1_R1192_U439 = ~new_P1_R1192_U438 | ~new_P1_R1192_U265;
  assign new_P1_R1192_U440 = ~new_P1_R1192_U136 | ~new_P1_R1192_U64;
  assign new_P1_R1192_U441 = ~new_P1_U3503 | ~new_P1_R1192_U63;
  assign new_P1_R1192_U442 = ~new_P1_U3069 | ~new_P1_R1192_U62;
  assign new_P1_R1192_U443 = ~new_P1_R1192_U137;
  assign new_P1_R1192_U444 = ~new_P1_R1192_U261 | ~new_P1_R1192_U443;
  assign new_P1_R1192_U445 = ~new_P1_R1192_U137 | ~new_P1_R1192_U164;
  assign new_P1_R1192_U446 = ~new_P1_U3500 | ~new_P1_R1192_U58;
  assign new_P1_R1192_U447 = ~new_P1_U3073 | ~new_P1_R1192_U56;
  assign new_P1_R1192_U448 = ~new_P1_R1192_U447 | ~new_P1_R1192_U446;
  assign new_P1_R1192_U449 = ~new_P1_U3497 | ~new_P1_R1192_U59;
  assign new_P1_R1192_U450 = ~new_P1_U3074 | ~new_P1_R1192_U46;
  assign new_P1_R1192_U451 = ~new_P1_R1192_U334 | ~new_P1_R1192_U89;
  assign new_P1_R1192_U452 = ~new_P1_R1192_U165 | ~new_P1_R1192_U326;
  assign new_P1_R1192_U453 = ~new_P1_U3494 | ~new_P1_R1192_U60;
  assign new_P1_R1192_U454 = ~new_P1_U3079 | ~new_P1_R1192_U57;
  assign new_P1_R1192_U455 = ~new_P1_R1192_U335 | ~new_P1_R1192_U167;
  assign new_P1_R1192_U456 = ~new_P1_R1192_U251 | ~new_P1_R1192_U166;
  assign new_P1_R1192_U457 = ~new_P1_U3491 | ~new_P1_R1192_U55;
  assign new_P1_R1192_U458 = ~new_P1_U3080 | ~new_P1_R1192_U54;
  assign new_P1_R1192_U459 = ~new_P1_R1192_U140;
  assign new_P1_R1192_U460 = ~new_P1_R1192_U247 | ~new_P1_R1192_U459;
  assign new_P1_R1192_U461 = ~new_P1_R1192_U140 | ~new_P1_R1192_U168;
  assign new_P1_R1192_U462 = ~new_P1_U3488 | ~new_P1_R1192_U53;
  assign new_P1_R1192_U463 = ~new_P1_U3072 | ~new_P1_R1192_U52;
  assign new_P1_R1192_U464 = ~new_P1_R1192_U141;
  assign new_P1_R1192_U465 = ~new_P1_R1192_U243 | ~new_P1_R1192_U464;
  assign new_P1_R1192_U466 = ~new_P1_R1192_U141 | ~new_P1_R1192_U169;
  assign new_P1_R1192_U467 = ~new_P1_U3485 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U468 = ~new_P1_U3063 | ~new_P1_R1192_U48;
  assign new_P1_R1192_U469 = ~new_P1_R1192_U468 | ~new_P1_R1192_U467;
  assign new_P1_R1192_U470 = ~new_P1_U3482 | ~new_P1_R1192_U50;
  assign new_P1_R1192_U471 = ~new_P1_U3062 | ~new_P1_R1192_U47;
  assign new_P1_R1192_U472 = ~new_P1_R1192_U345 | ~new_P1_R1192_U90;
  assign new_P1_R1192_U473 = ~new_P1_R1192_U170 | ~new_P1_R1192_U337;
  assign new_P1_LT_197_U6 = new_P1_LT_197_U115 & new_P1_LT_197_U116;
  assign new_P1_LT_197_U7 = new_P1_LT_197_U117 & new_P1_LT_197_U118;
  assign new_P1_LT_197_U8 = new_P1_LT_197_U7 & new_P1_LT_197_U122 & new_P1_LT_197_U81 & new_P1_LT_197_U120;
  assign new_P1_LT_197_U9 = new_P1_LT_197_U130 & new_P1_LT_197_U129;
  assign new_P1_LT_197_U10 = new_P1_LT_197_U85 & new_P1_LT_197_U84 & new_P1_LT_197_U131 & new_P1_LT_197_U128;
  assign new_P1_LT_197_U11 = new_P1_LT_197_U145 & new_P1_LT_197_U144;
  assign new_P1_LT_197_U12 = new_P1_LT_197_U193 & new_P1_LT_197_U72;
  assign new_P1_LT_197_U13 = new_P1_LT_197_U200 & new_P1_LT_197_U199;
  assign new_P1_LT_197_U14 = ~new_P1_U3983;
  assign new_P1_LT_197_U15 = ~new_P1_U3593;
  assign new_P1_LT_197_U16 = ~new_P1_U3594;
  assign new_P1_LT_197_U17 = ~new_P1_U3598;
  assign new_P1_LT_197_U18 = ~new_P1_U3599;
  assign new_P1_LT_197_U19 = ~new_P1_U3977;
  assign new_P1_LT_197_U20 = ~new_P1_U3978;
  assign new_P1_LT_197_U21 = ~new_P1_U3603;
  assign new_P1_LT_197_U22 = ~new_P1_U3981;
  assign new_P1_LT_197_U23 = ~new_P1_U3604;
  assign new_P1_LT_197_U24 = ~new_P1_U3982;
  assign new_P1_LT_197_U25 = ~new_P1_U3508;
  assign new_P1_LT_197_U26 = ~new_P1_U3608;
  assign new_P1_LT_197_U27 = ~new_P1_U3506;
  assign new_P1_LT_197_U28 = ~new_P1_U3609;
  assign new_P1_LT_197_U29 = ~new_P1_U3607;
  assign new_P1_LT_197_U30 = ~new_P1_U3605;
  assign new_P1_LT_197_U31 = ~new_P1_U3503;
  assign new_P1_LT_197_U32 = ~new_P1_U3500;
  assign new_P1_LT_197_U33 = ~new_P1_U3610;
  assign new_P1_LT_197_U34 = ~new_P1_U3611;
  assign new_P1_LT_197_U35 = ~new_P1_U3473;
  assign new_P1_LT_197_U36 = ~new_P1_U3589;
  assign new_P1_LT_197_U37 = ~new_P1_U3470;
  assign new_P1_LT_197_U38 = ~new_P1_U3590;
  assign new_P1_LT_197_U39 = ~new_P1_U3586;
  assign new_P1_LT_197_U40 = ~new_P1_U3616;
  assign new_P1_LT_197_U41 = ~new_P1_U3587;
  assign new_P1_LT_197_U42 = ~new_P1_U3588;
  assign new_P1_LT_197_U43 = ~new_P1_U3591;
  assign new_P1_LT_197_U44 = ~new_P1_U3592;
  assign new_P1_LT_197_U45 = ~new_P1_U3450 | ~new_P1_LT_197_U108;
  assign new_P1_LT_197_U46 = ~new_P1_U3455;
  assign new_P1_LT_197_U47 = ~new_P1_U3595;
  assign new_P1_LT_197_U48 = ~new_P1_U3488;
  assign new_P1_LT_197_U49 = ~new_P1_U3491;
  assign new_P1_LT_197_U50 = ~new_P1_U3458;
  assign new_P1_LT_197_U51 = ~new_P1_U3461;
  assign new_P1_LT_197_U52 = ~new_P1_U3464;
  assign new_P1_LT_197_U53 = ~new_P1_U3467;
  assign new_P1_LT_197_U54 = ~new_P1_U3476;
  assign new_P1_LT_197_U55 = ~new_P1_U3479;
  assign new_P1_LT_197_U56 = ~new_P1_U3482;
  assign new_P1_LT_197_U57 = ~new_P1_U3485;
  assign new_P1_LT_197_U58 = ~new_P1_U3614;
  assign new_P1_LT_197_U59 = ~new_P1_U3615;
  assign new_P1_LT_197_U60 = ~new_P1_U3612;
  assign new_P1_LT_197_U61 = ~new_P1_U3613;
  assign new_P1_LT_197_U62 = ~new_P1_U3494;
  assign new_P1_LT_197_U63 = ~new_P1_U3497;
  assign new_P1_LT_197_U64 = ~new_P1_U3980;
  assign new_P1_LT_197_U65 = ~new_P1_U3979;
  assign new_P1_LT_197_U66 = ~new_P1_U3602;
  assign new_P1_LT_197_U67 = ~new_P1_U3601;
  assign new_P1_LT_197_U68 = ~new_P1_U3600;
  assign new_P1_LT_197_U69 = ~new_P1_U3976;
  assign new_P1_LT_197_U70 = ~new_P1_U3975;
  assign new_P1_LT_197_U71 = ~new_P1_LT_197_U192 | ~new_P1_LT_197_U191;
  assign new_P1_LT_197_U72 = ~new_P1_U3974;
  assign new_P1_LT_197_U73 = ~new_P1_U3985;
  assign new_P1_LT_197_U74 = ~new_P1_U3596;
  assign new_P1_LT_197_U75 = ~new_P1_U3984;
  assign new_P1_LT_197_U76 = new_P1_U3981 & new_P1_LT_197_U23;
  assign new_P1_LT_197_U77 = new_P1_U3982 & new_P1_LT_197_U30;
  assign new_P1_LT_197_U78 = new_P1_LT_197_U175 & new_P1_LT_197_U174;
  assign new_P1_LT_197_U79 = new_P1_U3608 & new_P1_LT_197_U27;
  assign new_P1_LT_197_U80 = new_P1_U3609 & new_P1_LT_197_U31;
  assign new_P1_LT_197_U81 = new_P1_LT_197_U121 & new_P1_LT_197_U119;
  assign new_P1_LT_197_U82 = new_P1_U3589 & new_P1_LT_197_U37;
  assign new_P1_LT_197_U83 = new_P1_U3590 & new_P1_LT_197_U53;
  assign new_P1_LT_197_U84 = new_P1_LT_197_U133 & new_P1_LT_197_U132;
  assign new_P1_LT_197_U85 = new_P1_LT_197_U134 & new_P1_LT_197_U135 & new_P1_LT_197_U137 & new_P1_LT_197_U136;
  assign new_P1_LT_197_U86 = new_P1_LT_197_U141 & new_P1_LT_197_U142;
  assign new_P1_LT_197_U87 = new_P1_LT_197_U86 & new_P1_LT_197_U140;
  assign new_P1_LT_197_U88 = new_P1_U3458 & new_P1_LT_197_U47;
  assign new_P1_LT_197_U89 = new_P1_U3461 & new_P1_LT_197_U44;
  assign new_P1_LT_197_U90 = new_P1_LT_197_U134 & new_P1_LT_197_U135 & new_P1_LT_197_U128;
  assign new_P1_LT_197_U91 = new_P1_LT_197_U93 & new_P1_LT_197_U158 & new_P1_LT_197_U143;
  assign new_P1_LT_197_U92 = new_P1_LT_197_U161 & new_P1_LT_197_U160;
  assign new_P1_LT_197_U93 = new_P1_LT_197_U92 & new_P1_LT_197_U11;
  assign new_P1_LT_197_U94 = new_P1_U3614 & new_P1_LT_197_U48;
  assign new_P1_LT_197_U95 = new_P1_U3615 & new_P1_LT_197_U57;
  assign new_P1_LT_197_U96 = new_P1_LT_197_U164 & new_P1_LT_197_U98;
  assign new_P1_LT_197_U97 = new_P1_LT_197_U96 & new_P1_LT_197_U165;
  assign new_P1_LT_197_U98 = new_P1_LT_197_U167 & new_P1_LT_197_U166;
  assign new_P1_LT_197_U99 = new_P1_LT_197_U177 & new_P1_LT_197_U124;
  assign new_P1_LT_197_U100 = new_P1_LT_197_U179 & new_P1_LT_197_U178;
  assign new_P1_LT_197_U101 = new_P1_LT_197_U181 & new_P1_LT_197_U182;
  assign new_P1_LT_197_U102 = new_P1_U3602 & new_P1_LT_197_U65;
  assign new_P1_LT_197_U103 = new_P1_LT_197_U186 & new_P1_LT_197_U185;
  assign new_P1_LT_197_U104 = new_P1_LT_197_U189 & new_P1_LT_197_U125;
  assign new_P1_LT_197_U105 = new_P1_LT_197_U196 & new_P1_LT_197_U195;
  assign new_P1_LT_197_U106 = new_P1_U3596 & new_P1_LT_197_U73;
  assign new_P1_LT_197_U107 = new_P1_LT_197_U198 & new_P1_LT_197_U112;
  assign new_P1_LT_197_U108 = ~new_P1_U3617;
  assign new_P1_LT_197_U109 = ~new_P1_LT_197_U107 | ~new_P1_LT_197_U197;
  assign new_P1_LT_197_U110 = ~new_P1_U3984 | ~new_P1_LT_197_U16;
  assign new_P1_LT_197_U111 = ~new_P1_U3593 | ~new_P1_LT_197_U14;
  assign new_P1_LT_197_U112 = ~new_P1_LT_197_U75 | ~new_P1_LT_197_U111 | ~new_P1_U3594;
  assign new_P1_LT_197_U113 = ~new_P1_U3593 | ~new_P1_LT_197_U14;
  assign new_P1_LT_197_U114 = ~new_P1_U3598 | ~new_P1_LT_197_U70;
  assign new_P1_LT_197_U115 = ~new_P1_U3508 | ~new_P1_LT_197_U29;
  assign new_P1_LT_197_U116 = ~new_P1_U3506 | ~new_P1_LT_197_U26;
  assign new_P1_LT_197_U117 = ~new_P1_U3603 | ~new_P1_LT_197_U64;
  assign new_P1_LT_197_U118 = ~new_P1_U3604 | ~new_P1_LT_197_U22;
  assign new_P1_LT_197_U119 = ~new_P1_LT_197_U79 | ~new_P1_LT_197_U115;
  assign new_P1_LT_197_U120 = ~new_P1_LT_197_U80 | ~new_P1_LT_197_U6;
  assign new_P1_LT_197_U121 = ~new_P1_U3607 | ~new_P1_LT_197_U25;
  assign new_P1_LT_197_U122 = ~new_P1_U3605 | ~new_P1_LT_197_U24;
  assign new_P1_LT_197_U123 = ~new_P1_U3610 | ~new_P1_LT_197_U32;
  assign new_P1_LT_197_U124 = ~new_P1_U3978 | ~new_P1_LT_197_U67;
  assign new_P1_LT_197_U125 = ~new_P1_U3977 | ~new_P1_LT_197_U68;
  assign new_P1_LT_197_U126 = ~new_P1_U3611 | ~new_P1_LT_197_U63;
  assign new_P1_LT_197_U127 = ~new_P1_U3473 | ~new_P1_LT_197_U42;
  assign new_P1_LT_197_U128 = ~new_P1_LT_197_U82 | ~new_P1_LT_197_U127;
  assign new_P1_LT_197_U129 = ~new_P1_U3470 | ~new_P1_LT_197_U36;
  assign new_P1_LT_197_U130 = ~new_P1_U3473 | ~new_P1_LT_197_U42;
  assign new_P1_LT_197_U131 = ~new_P1_LT_197_U83 | ~new_P1_LT_197_U9;
  assign new_P1_LT_197_U132 = ~new_P1_U3586 | ~new_P1_LT_197_U55;
  assign new_P1_LT_197_U133 = ~new_P1_U3616 | ~new_P1_LT_197_U56;
  assign new_P1_LT_197_U134 = ~new_P1_U3587 | ~new_P1_LT_197_U54;
  assign new_P1_LT_197_U135 = ~new_P1_U3588 | ~new_P1_LT_197_U35;
  assign new_P1_LT_197_U136 = ~new_P1_U3591 | ~new_P1_LT_197_U52;
  assign new_P1_LT_197_U137 = ~new_P1_U3592 | ~new_P1_LT_197_U51;
  assign new_P1_LT_197_U138 = ~new_P1_LT_197_U45;
  assign new_P1_LT_197_U139 = ~new_P1_U3455 | ~new_P1_LT_197_U138;
  assign new_P1_LT_197_U140 = ~new_P1_U3606 | ~new_P1_LT_197_U139;
  assign new_P1_LT_197_U141 = ~new_P1_LT_197_U45 | ~new_P1_LT_197_U46;
  assign new_P1_LT_197_U142 = ~new_P1_U3595 | ~new_P1_LT_197_U50;
  assign new_P1_LT_197_U143 = ~new_P1_LT_197_U87 | ~new_P1_LT_197_U10;
  assign new_P1_LT_197_U144 = ~new_P1_U3488 | ~new_P1_LT_197_U58;
  assign new_P1_LT_197_U145 = ~new_P1_U3491 | ~new_P1_LT_197_U61;
  assign new_P1_LT_197_U146 = ~new_P1_LT_197_U89 | ~new_P1_LT_197_U136;
  assign new_P1_LT_197_U147 = ~new_P1_U3464 | ~new_P1_LT_197_U43;
  assign new_P1_LT_197_U148 = ~new_P1_LT_197_U9 | ~new_P1_LT_197_U147 | ~new_P1_LT_197_U146;
  assign new_P1_LT_197_U149 = ~new_P1_LT_197_U148 | ~new_P1_LT_197_U131;
  assign new_P1_LT_197_U150 = ~new_P1_U3467 | ~new_P1_LT_197_U38;
  assign new_P1_LT_197_U151 = ~new_P1_LT_197_U150 | ~new_P1_LT_197_U149;
  assign new_P1_LT_197_U152 = ~new_P1_LT_197_U90 | ~new_P1_LT_197_U151;
  assign new_P1_LT_197_U153 = ~new_P1_U3476 | ~new_P1_LT_197_U41;
  assign new_P1_LT_197_U154 = ~new_P1_LT_197_U153 | ~new_P1_LT_197_U152;
  assign new_P1_LT_197_U155 = ~new_P1_LT_197_U154 | ~new_P1_LT_197_U132;
  assign new_P1_LT_197_U156 = ~new_P1_U3479 | ~new_P1_LT_197_U39;
  assign new_P1_LT_197_U157 = ~new_P1_LT_197_U156 | ~new_P1_LT_197_U155;
  assign new_P1_LT_197_U158 = ~new_P1_LT_197_U88 | ~new_P1_LT_197_U10;
  assign new_P1_LT_197_U159 = ~new_P1_LT_197_U157 | ~new_P1_LT_197_U133;
  assign new_P1_LT_197_U160 = ~new_P1_U3482 | ~new_P1_LT_197_U40;
  assign new_P1_LT_197_U161 = ~new_P1_U3485 | ~new_P1_LT_197_U59;
  assign new_P1_LT_197_U162 = ~new_P1_LT_197_U159 | ~new_P1_LT_197_U91;
  assign new_P1_LT_197_U163 = ~new_P1_U3491 | ~new_P1_LT_197_U61;
  assign new_P1_LT_197_U164 = ~new_P1_LT_197_U94 | ~new_P1_LT_197_U163;
  assign new_P1_LT_197_U165 = ~new_P1_LT_197_U95 | ~new_P1_LT_197_U11;
  assign new_P1_LT_197_U166 = ~new_P1_U3612 | ~new_P1_LT_197_U62;
  assign new_P1_LT_197_U167 = ~new_P1_U3613 | ~new_P1_LT_197_U49;
  assign new_P1_LT_197_U168 = ~new_P1_LT_197_U162 | ~new_P1_LT_197_U97;
  assign new_P1_LT_197_U169 = ~new_P1_U3494 | ~new_P1_LT_197_U60;
  assign new_P1_LT_197_U170 = ~new_P1_LT_197_U169 | ~new_P1_LT_197_U168;
  assign new_P1_LT_197_U171 = ~new_P1_LT_197_U170 | ~new_P1_LT_197_U126;
  assign new_P1_LT_197_U172 = ~new_P1_U3497 | ~new_P1_LT_197_U34;
  assign new_P1_LT_197_U173 = ~new_P1_LT_197_U172 | ~new_P1_LT_197_U171;
  assign new_P1_LT_197_U174 = ~new_P1_U3503 | ~new_P1_LT_197_U28;
  assign new_P1_LT_197_U175 = ~new_P1_U3500 | ~new_P1_LT_197_U33;
  assign new_P1_LT_197_U176 = ~new_P1_LT_197_U78 | ~new_P1_LT_197_U6;
  assign new_P1_LT_197_U177 = ~new_P1_LT_197_U76 | ~new_P1_LT_197_U117;
  assign new_P1_LT_197_U178 = ~new_P1_LT_197_U77 | ~new_P1_LT_197_U7;
  assign new_P1_LT_197_U179 = ~new_P1_LT_197_U8 | ~new_P1_LT_197_U176;
  assign new_P1_LT_197_U180 = ~new_P1_LT_197_U8 | ~new_P1_LT_197_U173 | ~new_P1_LT_197_U123;
  assign new_P1_LT_197_U181 = ~new_P1_U3980 | ~new_P1_LT_197_U21;
  assign new_P1_LT_197_U182 = ~new_P1_U3979 | ~new_P1_LT_197_U66;
  assign new_P1_LT_197_U183 = ~new_P1_LT_197_U99 | ~new_P1_LT_197_U100 | ~new_P1_LT_197_U101 | ~new_P1_LT_197_U180;
  assign new_P1_LT_197_U184 = ~new_P1_LT_197_U102 | ~new_P1_LT_197_U124;
  assign new_P1_LT_197_U185 = ~new_P1_U3601 | ~new_P1_LT_197_U20;
  assign new_P1_LT_197_U186 = ~new_P1_U3600 | ~new_P1_LT_197_U19;
  assign new_P1_LT_197_U187 = ~new_P1_U3599 | ~new_P1_LT_197_U69;
  assign new_P1_LT_197_U188 = ~new_P1_LT_197_U103 | ~new_P1_LT_197_U184 | ~new_P1_LT_197_U183;
  assign new_P1_LT_197_U189 = ~new_P1_U3976 | ~new_P1_LT_197_U18;
  assign new_P1_LT_197_U190 = ~new_P1_LT_197_U104 | ~new_P1_LT_197_U188;
  assign new_P1_LT_197_U191 = ~new_P1_LT_197_U114 | ~new_P1_LT_197_U187 | ~new_P1_LT_197_U190;
  assign new_P1_LT_197_U192 = ~new_P1_U3975 | ~new_P1_LT_197_U17;
  assign new_P1_LT_197_U193 = ~new_P1_LT_197_U71;
  assign new_P1_LT_197_U194 = new_P1_U3597 | new_P1_LT_197_U12;
  assign new_P1_LT_197_U195 = ~new_P1_U3974 | ~new_P1_LT_197_U71;
  assign new_P1_LT_197_U196 = ~new_P1_U3985 | ~new_P1_LT_197_U74;
  assign new_P1_LT_197_U197 = ~new_P1_LT_197_U105 | ~new_P1_LT_197_U194 | ~new_P1_LT_197_U113;
  assign new_P1_LT_197_U198 = ~new_P1_LT_197_U106 | ~new_P1_LT_197_U113;
  assign new_P1_LT_197_U199 = ~new_P1_U3983 | ~new_P1_LT_197_U15;
  assign new_P1_LT_197_U200 = ~new_P1_LT_197_U110 | ~new_P1_LT_197_U109;
  assign new_P1_R1360_U6 = new_P1_R1360_U111 & new_P1_R1360_U112;
  assign new_P1_R1360_U7 = new_P1_R1360_U116 & new_P1_R1360_U115;
  assign new_P1_R1360_U8 = new_P1_R1360_U118 & new_P1_R1360_U119;
  assign new_P1_R1360_U9 = new_P1_R1360_U123 & new_P1_R1360_U122;
  assign new_P1_R1360_U10 = new_P1_R1360_U183 & new_P1_R1360_U184 & new_P1_R1360_U186 & new_P1_R1360_U199 & new_P1_R1360_U185;
  assign new_P1_R1360_U11 = new_P1_R1360_U183 & new_P1_R1360_U104;
  assign new_P1_R1360_U12 = new_P1_R1360_U203 & new_P1_R1360_U202;
  assign new_P1_R1360_U13 = new_P1_R1360_U205 & new_P1_R1360_U204;
  assign new_P1_R1360_U14 = ~new_P1_R1360_U107 | ~new_P1_R1360_U108 | ~new_P1_R1360_U200;
  assign new_P1_R1360_U15 = ~new_P1_U3088;
  assign new_P1_R1360_U16 = ~new_P1_U3087;
  assign new_P1_R1360_U17 = ~new_P1_U3121;
  assign new_P1_R1360_U18 = ~new_P1_U3089;
  assign new_P1_R1360_U19 = ~new_P1_U3090;
  assign new_P1_R1360_U20 = ~new_P1_U3123;
  assign new_P1_R1360_U21 = ~new_P1_U3122;
  assign new_P1_R1360_U22 = ~new_P1_U3120;
  assign new_P1_R1360_U23 = ~new_P1_U3127;
  assign new_P1_R1360_U24 = ~new_P1_U3126;
  assign new_P1_R1360_U25 = ~new_P1_U3097;
  assign new_P1_R1360_U26 = ~new_P1_U3098;
  assign new_P1_R1360_U27 = ~new_P1_U3133;
  assign new_P1_R1360_U28 = ~new_P1_U3132;
  assign new_P1_R1360_U29 = ~new_P1_U3103;
  assign new_P1_R1360_U30 = ~new_P1_U3104;
  assign new_P1_R1360_U31 = ~new_P1_U3139;
  assign new_P1_R1360_U32 = ~new_P1_U3138;
  assign new_P1_R1360_U33 = ~new_P1_U3109;
  assign new_P1_R1360_U34 = ~new_P1_U3142;
  assign new_P1_R1360_U35 = ~new_P1_U3110;
  assign new_P1_R1360_U36 = ~new_P1_U3143;
  assign new_P1_R1360_U37 = ~new_P1_U3112;
  assign new_P1_R1360_U38 = ~new_P1_U3111;
  assign new_P1_R1360_U39 = ~new_P1_U3114;
  assign new_P1_R1360_U40 = ~new_P1_U3113;
  assign new_P1_R1360_U41 = ~new_P1_U3116;
  assign new_P1_R1360_U42 = ~new_P1_U3115;
  assign new_P1_R1360_U43 = ~new_P1_U3117;
  assign new_P1_R1360_U44 = ~new_P1_U3149;
  assign new_P1_R1360_U45 = ~new_P1_U3148;
  assign new_P1_R1360_U46 = ~new_P1_U3147;
  assign new_P1_R1360_U47 = ~new_P1_U3146;
  assign new_P1_R1360_U48 = ~new_P1_U3145;
  assign new_P1_R1360_U49 = ~new_P1_U3144;
  assign new_P1_R1360_U50 = ~new_P1_U3141;
  assign new_P1_R1360_U51 = ~new_P1_U3140;
  assign new_P1_R1360_U52 = ~new_P1_U3108;
  assign new_P1_R1360_U53 = ~new_P1_U3106;
  assign new_P1_R1360_U54 = ~new_P1_U3107;
  assign new_P1_R1360_U55 = ~new_P1_U3105;
  assign new_P1_R1360_U56 = ~new_P1_U3137;
  assign new_P1_R1360_U57 = ~new_P1_U3136;
  assign new_P1_R1360_U58 = ~new_P1_U3135;
  assign new_P1_R1360_U59 = ~new_P1_U3134;
  assign new_P1_R1360_U60 = ~new_P1_U3102;
  assign new_P1_R1360_U61 = ~new_P1_U3101;
  assign new_P1_R1360_U62 = ~new_P1_U3100;
  assign new_P1_R1360_U63 = ~new_P1_U3099;
  assign new_P1_R1360_U64 = ~new_P1_U3131;
  assign new_P1_R1360_U65 = ~new_P1_U3130;
  assign new_P1_R1360_U66 = ~new_P1_U3129;
  assign new_P1_R1360_U67 = ~new_P1_U3128;
  assign new_P1_R1360_U68 = ~new_P1_U3092;
  assign new_P1_R1360_U69 = ~new_P1_U3091;
  assign new_P1_R1360_U70 = ~new_P1_U3095;
  assign new_P1_R1360_U71 = ~new_P1_U3096;
  assign new_P1_R1360_U72 = ~new_P1_U3093;
  assign new_P1_R1360_U73 = ~new_P1_U3094;
  assign new_P1_R1360_U74 = ~new_P1_U3124;
  assign new_P1_R1360_U75 = ~new_P1_U3125;
  assign new_P1_R1360_U76 = ~new_P1_U3152;
  assign new_P1_R1360_U77 = new_P1_R1360_U18 & new_P1_U3121;
  assign new_P1_R1360_U78 = new_P1_R1360_U183 & new_P1_R1360_U184;
  assign new_P1_R1360_U79 = new_P1_U3142 & new_P1_R1360_U35;
  assign new_P1_R1360_U80 = new_P1_U3143 & new_P1_R1360_U38;
  assign new_P1_R1360_U81 = new_P1_R1360_U124 & new_P1_R1360_U125 & new_P1_R1360_U127 & new_P1_R1360_U126;
  assign new_P1_R1360_U82 = new_P1_R1360_U129 & new_P1_R1360_U130 & new_P1_R1360_U131;
  assign new_P1_R1360_U83 = new_P1_U3149 & new_P1_R1360_U43;
  assign new_P1_R1360_U84 = new_P1_R1360_U85 & new_P1_R1360_U132;
  assign new_P1_R1360_U85 = new_P1_R1360_U144 & new_P1_R1360_U143;
  assign new_P1_R1360_U86 = new_P1_R1360_U121 & new_P1_R1360_U120;
  assign new_P1_R1360_U87 = new_P1_R1360_U8 & new_P1_R1360_U86;
  assign new_P1_R1360_U88 = new_P1_R1360_U90 & new_P1_R1360_U147 & new_P1_R1360_U146;
  assign new_P1_R1360_U89 = new_P1_R1360_U150 & new_P1_R1360_U149;
  assign new_P1_R1360_U90 = new_P1_R1360_U89 & new_P1_R1360_U9;
  assign new_P1_R1360_U91 = new_P1_U3108 & new_P1_R1360_U51;
  assign new_P1_R1360_U92 = new_P1_U3107 & new_P1_R1360_U31;
  assign new_P1_R1360_U93 = new_P1_R1360_U94 & new_P1_R1360_U152 & new_P1_R1360_U153;
  assign new_P1_R1360_U94 = new_P1_R1360_U156 & new_P1_R1360_U155;
  assign new_P1_R1360_U95 = new_P1_R1360_U7 & new_P1_R1360_U96;
  assign new_P1_R1360_U96 = new_P1_R1360_U164 & new_P1_R1360_U165;
  assign new_P1_R1360_U97 = new_P1_U3102 & new_P1_R1360_U59;
  assign new_P1_R1360_U98 = new_P1_U3101 & new_P1_R1360_U27;
  assign new_P1_R1360_U99 = new_P1_R1360_U100 & new_P1_R1360_U167 & new_P1_R1360_U169;
  assign new_P1_R1360_U100 = new_P1_R1360_U171 & new_P1_R1360_U170;
  assign new_P1_R1360_U101 = new_P1_R1360_U179 & new_P1_R1360_U180;
  assign new_P1_R1360_U102 = new_P1_U3095 & new_P1_R1360_U23;
  assign new_P1_R1360_U103 = new_P1_U3096 & new_P1_R1360_U67;
  assign new_P1_R1360_U104 = new_P1_R1360_U184 & new_P1_R1360_U106 & new_P1_R1360_U186 & new_P1_R1360_U181 & new_P1_R1360_U185;
  assign new_P1_R1360_U105 = new_P1_R1360_U190 & new_P1_R1360_U189;
  assign new_P1_R1360_U106 = new_P1_R1360_U105 & new_P1_R1360_U188 & new_P1_R1360_U187;
  assign new_P1_R1360_U107 = new_P1_R1360_U195 & new_P1_R1360_U196 & new_P1_R1360_U194;
  assign new_P1_R1360_U108 = new_P1_R1360_U201 & new_P1_R1360_U13;
  assign new_P1_R1360_U109 = ~new_P1_U3119;
  assign new_P1_R1360_U110 = ~new_P1_U3097 | ~new_P1_R1360_U66;
  assign new_P1_R1360_U111 = ~new_P1_U3126 | ~new_P1_R1360_U73;
  assign new_P1_R1360_U112 = ~new_P1_U3127 | ~new_P1_R1360_U70;
  assign new_P1_R1360_U113 = ~new_P1_U3098 | ~new_P1_R1360_U65;
  assign new_P1_R1360_U114 = ~new_P1_U3103 | ~new_P1_R1360_U58;
  assign new_P1_R1360_U115 = ~new_P1_U3133 | ~new_P1_R1360_U61;
  assign new_P1_R1360_U116 = ~new_P1_U3132 | ~new_P1_R1360_U62;
  assign new_P1_R1360_U117 = ~new_P1_U3104 | ~new_P1_R1360_U57;
  assign new_P1_R1360_U118 = ~new_P1_U3109 | ~new_P1_R1360_U50;
  assign new_P1_R1360_U119 = ~new_P1_U3110 | ~new_P1_R1360_U34;
  assign new_P1_R1360_U120 = ~new_P1_U3112 | ~new_P1_R1360_U49;
  assign new_P1_R1360_U121 = ~new_P1_U3111 | ~new_P1_R1360_U36;
  assign new_P1_R1360_U122 = ~new_P1_U3139 | ~new_P1_R1360_U54;
  assign new_P1_R1360_U123 = ~new_P1_U3138 | ~new_P1_R1360_U53;
  assign new_P1_R1360_U124 = ~new_P1_U3114 | ~new_P1_R1360_U47;
  assign new_P1_R1360_U125 = ~new_P1_U3113 | ~new_P1_R1360_U48;
  assign new_P1_R1360_U126 = ~new_P1_U3116 | ~new_P1_R1360_U45;
  assign new_P1_R1360_U127 = ~new_P1_U3115 | ~new_P1_R1360_U46;
  assign new_P1_R1360_U128 = ~new_P1_U3150 | ~new_P1_U3151;
  assign new_P1_R1360_U129 = ~new_P1_U3118 | ~new_P1_R1360_U128;
  assign new_P1_R1360_U130 = new_P1_U3150 | new_P1_U3151;
  assign new_P1_R1360_U131 = ~new_P1_U3117 | ~new_P1_R1360_U44;
  assign new_P1_R1360_U132 = ~new_P1_R1360_U82 | ~new_P1_R1360_U81;
  assign new_P1_R1360_U133 = ~new_P1_R1360_U83 | ~new_P1_R1360_U126;
  assign new_P1_R1360_U134 = ~new_P1_U3148 | ~new_P1_R1360_U41;
  assign new_P1_R1360_U135 = ~new_P1_R1360_U134 | ~new_P1_R1360_U133;
  assign new_P1_R1360_U136 = ~new_P1_R1360_U135 | ~new_P1_R1360_U127;
  assign new_P1_R1360_U137 = ~new_P1_U3147 | ~new_P1_R1360_U42;
  assign new_P1_R1360_U138 = ~new_P1_R1360_U137 | ~new_P1_R1360_U136;
  assign new_P1_R1360_U139 = ~new_P1_R1360_U138 | ~new_P1_R1360_U124;
  assign new_P1_R1360_U140 = ~new_P1_U3146 | ~new_P1_R1360_U39;
  assign new_P1_R1360_U141 = ~new_P1_R1360_U140 | ~new_P1_R1360_U139;
  assign new_P1_R1360_U142 = ~new_P1_R1360_U141 | ~new_P1_R1360_U125;
  assign new_P1_R1360_U143 = ~new_P1_U3145 | ~new_P1_R1360_U40;
  assign new_P1_R1360_U144 = ~new_P1_U3144 | ~new_P1_R1360_U37;
  assign new_P1_R1360_U145 = ~new_P1_R1360_U142 | ~new_P1_R1360_U84;
  assign new_P1_R1360_U146 = ~new_P1_R1360_U79 | ~new_P1_R1360_U118;
  assign new_P1_R1360_U147 = ~new_P1_R1360_U80 | ~new_P1_R1360_U8;
  assign new_P1_R1360_U148 = ~new_P1_R1360_U87 | ~new_P1_R1360_U145;
  assign new_P1_R1360_U149 = ~new_P1_U3141 | ~new_P1_R1360_U33;
  assign new_P1_R1360_U150 = ~new_P1_U3140 | ~new_P1_R1360_U52;
  assign new_P1_R1360_U151 = ~new_P1_R1360_U148 | ~new_P1_R1360_U88;
  assign new_P1_R1360_U152 = ~new_P1_R1360_U91 | ~new_P1_R1360_U9;
  assign new_P1_R1360_U153 = ~new_P1_U3106 | ~new_P1_R1360_U32;
  assign new_P1_R1360_U154 = ~new_P1_U3138 | ~new_P1_R1360_U53;
  assign new_P1_R1360_U155 = ~new_P1_R1360_U92 | ~new_P1_R1360_U154;
  assign new_P1_R1360_U156 = ~new_P1_U3105 | ~new_P1_R1360_U56;
  assign new_P1_R1360_U157 = ~new_P1_R1360_U151 | ~new_P1_R1360_U93;
  assign new_P1_R1360_U158 = ~new_P1_U3137 | ~new_P1_R1360_U55;
  assign new_P1_R1360_U159 = ~new_P1_R1360_U158 | ~new_P1_R1360_U157;
  assign new_P1_R1360_U160 = ~new_P1_R1360_U159 | ~new_P1_R1360_U117;
  assign new_P1_R1360_U161 = ~new_P1_U3136 | ~new_P1_R1360_U30;
  assign new_P1_R1360_U162 = ~new_P1_R1360_U161 | ~new_P1_R1360_U160;
  assign new_P1_R1360_U163 = ~new_P1_R1360_U162 | ~new_P1_R1360_U114;
  assign new_P1_R1360_U164 = ~new_P1_U3135 | ~new_P1_R1360_U29;
  assign new_P1_R1360_U165 = ~new_P1_U3134 | ~new_P1_R1360_U60;
  assign new_P1_R1360_U166 = ~new_P1_R1360_U163 | ~new_P1_R1360_U95;
  assign new_P1_R1360_U167 = ~new_P1_R1360_U97 | ~new_P1_R1360_U7;
  assign new_P1_R1360_U168 = ~new_P1_U3132 | ~new_P1_R1360_U62;
  assign new_P1_R1360_U169 = ~new_P1_R1360_U98 | ~new_P1_R1360_U168;
  assign new_P1_R1360_U170 = ~new_P1_U3100 | ~new_P1_R1360_U28;
  assign new_P1_R1360_U171 = ~new_P1_U3099 | ~new_P1_R1360_U64;
  assign new_P1_R1360_U172 = ~new_P1_R1360_U166 | ~new_P1_R1360_U99;
  assign new_P1_R1360_U173 = ~new_P1_U3131 | ~new_P1_R1360_U63;
  assign new_P1_R1360_U174 = ~new_P1_R1360_U173 | ~new_P1_R1360_U172;
  assign new_P1_R1360_U175 = ~new_P1_R1360_U174 | ~new_P1_R1360_U113;
  assign new_P1_R1360_U176 = ~new_P1_U3130 | ~new_P1_R1360_U26;
  assign new_P1_R1360_U177 = ~new_P1_R1360_U176 | ~new_P1_R1360_U175;
  assign new_P1_R1360_U178 = ~new_P1_R1360_U177 | ~new_P1_R1360_U110;
  assign new_P1_R1360_U179 = ~new_P1_U3129 | ~new_P1_R1360_U25;
  assign new_P1_R1360_U180 = ~new_P1_U3128 | ~new_P1_R1360_U71;
  assign new_P1_R1360_U181 = ~new_P1_R1360_U6 | ~new_P1_R1360_U101 | ~new_P1_R1360_U178;
  assign new_P1_R1360_U182 = ~new_P1_U3088 | ~new_P1_R1360_U22;
  assign new_P1_R1360_U183 = ~new_P1_U3089 | ~new_P1_R1360_U17;
  assign new_P1_R1360_U184 = ~new_P1_U3090 | ~new_P1_R1360_U21;
  assign new_P1_R1360_U185 = ~new_P1_U3092 | ~new_P1_R1360_U74;
  assign new_P1_R1360_U186 = ~new_P1_U3091 | ~new_P1_R1360_U20;
  assign new_P1_R1360_U187 = ~new_P1_R1360_U102 | ~new_P1_R1360_U111;
  assign new_P1_R1360_U188 = ~new_P1_R1360_U103 | ~new_P1_R1360_U6;
  assign new_P1_R1360_U189 = ~new_P1_U3093 | ~new_P1_R1360_U75;
  assign new_P1_R1360_U190 = ~new_P1_U3094 | ~new_P1_R1360_U24;
  assign new_P1_R1360_U191 = ~new_P1_U3123 | ~new_P1_R1360_U69;
  assign new_P1_R1360_U192 = ~new_P1_U3122 | ~new_P1_R1360_U19;
  assign new_P1_R1360_U193 = ~new_P1_R1360_U192 | ~new_P1_R1360_U191;
  assign new_P1_R1360_U194 = ~new_P1_R1360_U182 | ~new_P1_R1360_U77 | ~new_P1_R1360_U12;
  assign new_P1_R1360_U195 = ~new_P1_R1360_U182 | ~new_P1_R1360_U78 | ~new_P1_R1360_U12 | ~new_P1_R1360_U193;
  assign new_P1_R1360_U196 = ~new_P1_U3120 | ~new_P1_R1360_U12 | ~new_P1_R1360_U15;
  assign new_P1_R1360_U197 = ~new_P1_U3124 | ~new_P1_R1360_U68;
  assign new_P1_R1360_U198 = ~new_P1_U3125 | ~new_P1_R1360_U72;
  assign new_P1_R1360_U199 = ~new_P1_R1360_U198 | ~new_P1_R1360_U197;
  assign new_P1_R1360_U200 = ~new_P1_R1360_U182 | ~new_P1_R1360_U12 | ~new_P1_R1360_U11;
  assign new_P1_R1360_U201 = ~new_P1_R1360_U182 | ~new_P1_R1360_U12 | ~new_P1_R1360_U10;
  assign new_P1_R1360_U202 = ~new_P1_U3087 | ~new_P1_R1360_U109;
  assign new_P1_R1360_U203 = ~new_P1_U3119 | ~new_P1_R1360_U16;
  assign new_P1_R1360_U204 = ~new_P1_R1360_U109 | ~new_P1_U3152 | ~new_P1_U3087;
  assign new_P1_R1360_U205 = ~new_P1_U3119 | ~new_P1_R1360_U76 | ~new_P1_R1360_U16;
  assign new_P1_R1171_U4 = new_P1_R1171_U178 & new_P1_R1171_U177;
  assign new_P1_R1171_U5 = new_P1_R1171_U179 & new_P1_R1171_U180;
  assign new_P1_R1171_U6 = new_P1_R1171_U196 & new_P1_R1171_U195;
  assign new_P1_R1171_U7 = new_P1_R1171_U236 & new_P1_R1171_U235;
  assign new_P1_R1171_U8 = new_P1_R1171_U245 & new_P1_R1171_U244;
  assign new_P1_R1171_U9 = new_P1_R1171_U263 & new_P1_R1171_U262;
  assign new_P1_R1171_U10 = new_P1_R1171_U271 & new_P1_R1171_U270;
  assign new_P1_R1171_U11 = new_P1_R1171_U350 & new_P1_R1171_U347;
  assign new_P1_R1171_U12 = new_P1_R1171_U343 & new_P1_R1171_U340;
  assign new_P1_R1171_U13 = new_P1_R1171_U334 & new_P1_R1171_U331;
  assign new_P1_R1171_U14 = new_P1_R1171_U325 & new_P1_R1171_U322;
  assign new_P1_R1171_U15 = new_P1_R1171_U319 & new_P1_R1171_U317;
  assign new_P1_R1171_U16 = new_P1_R1171_U312 & new_P1_R1171_U309;
  assign new_P1_R1171_U17 = new_P1_R1171_U234 & new_P1_R1171_U231;
  assign new_P1_R1171_U18 = new_P1_R1171_U226 & new_P1_R1171_U223;
  assign new_P1_R1171_U19 = new_P1_R1171_U212 & new_P1_R1171_U209;
  assign new_P1_R1171_U20 = ~new_P1_U3470;
  assign new_P1_R1171_U21 = ~new_P1_U3071;
  assign new_P1_R1171_U22 = ~new_P1_U3070;
  assign new_P1_R1171_U23 = ~new_P1_U3071 | ~new_P1_U3470;
  assign new_P1_R1171_U24 = ~new_P1_U3473;
  assign new_P1_R1171_U25 = ~new_P1_U3464;
  assign new_P1_R1171_U26 = ~new_P1_U3060;
  assign new_P1_R1171_U27 = ~new_P1_U3067;
  assign new_P1_R1171_U28 = ~new_P1_U3458;
  assign new_P1_R1171_U29 = ~new_P1_U3068;
  assign new_P1_R1171_U30 = ~new_P1_U3450;
  assign new_P1_R1171_U31 = ~new_P1_U3077;
  assign new_P1_R1171_U32 = ~new_P1_U3077 | ~new_P1_U3450;
  assign new_P1_R1171_U33 = ~new_P1_U3461;
  assign new_P1_R1171_U34 = ~new_P1_U3064;
  assign new_P1_R1171_U35 = ~new_P1_U3060 | ~new_P1_U3464;
  assign new_P1_R1171_U36 = ~new_P1_U3467;
  assign new_P1_R1171_U37 = ~new_P1_U3476;
  assign new_P1_R1171_U38 = ~new_P1_U3084;
  assign new_P1_R1171_U39 = ~new_P1_U3083;
  assign new_P1_R1171_U40 = ~new_P1_U3479;
  assign new_P1_R1171_U41 = ~new_P1_R1171_U62 | ~new_P1_R1171_U204;
  assign new_P1_R1171_U42 = ~new_P1_R1171_U118 | ~new_P1_R1171_U192;
  assign new_P1_R1171_U43 = ~new_P1_R1171_U181 | ~new_P1_R1171_U182;
  assign new_P1_R1171_U44 = ~new_P1_U3455 | ~new_P1_U3078;
  assign new_P1_R1171_U45 = ~new_P1_R1171_U122 | ~new_P1_R1171_U218;
  assign new_P1_R1171_U46 = ~new_P1_R1171_U215 | ~new_P1_R1171_U214;
  assign new_P1_R1171_U47 = ~new_P1_U3975;
  assign new_P1_R1171_U48 = ~new_P1_U3053;
  assign new_P1_R1171_U49 = ~new_P1_U3057;
  assign new_P1_R1171_U50 = ~new_P1_U3976;
  assign new_P1_R1171_U51 = ~new_P1_U3977;
  assign new_P1_R1171_U52 = ~new_P1_U3058;
  assign new_P1_R1171_U53 = ~new_P1_U3978;
  assign new_P1_R1171_U54 = ~new_P1_U3065;
  assign new_P1_R1171_U55 = ~new_P1_U3981;
  assign new_P1_R1171_U56 = ~new_P1_U3075;
  assign new_P1_R1171_U57 = ~new_P1_U3500;
  assign new_P1_R1171_U58 = ~new_P1_U3073;
  assign new_P1_R1171_U59 = ~new_P1_U3069;
  assign new_P1_R1171_U60 = ~new_P1_U3073 | ~new_P1_U3500;
  assign new_P1_R1171_U61 = ~new_P1_U3503;
  assign new_P1_R1171_U62 = ~new_P1_U3084 | ~new_P1_U3476;
  assign new_P1_R1171_U63 = ~new_P1_U3482;
  assign new_P1_R1171_U64 = ~new_P1_U3062;
  assign new_P1_R1171_U65 = ~new_P1_U3488;
  assign new_P1_R1171_U66 = ~new_P1_U3072;
  assign new_P1_R1171_U67 = ~new_P1_U3485;
  assign new_P1_R1171_U68 = ~new_P1_U3063;
  assign new_P1_R1171_U69 = ~new_P1_U3063 | ~new_P1_U3485;
  assign new_P1_R1171_U70 = ~new_P1_U3491;
  assign new_P1_R1171_U71 = ~new_P1_U3080;
  assign new_P1_R1171_U72 = ~new_P1_U3494;
  assign new_P1_R1171_U73 = ~new_P1_U3079;
  assign new_P1_R1171_U74 = ~new_P1_U3497;
  assign new_P1_R1171_U75 = ~new_P1_U3074;
  assign new_P1_R1171_U76 = ~new_P1_U3506;
  assign new_P1_R1171_U77 = ~new_P1_U3082;
  assign new_P1_R1171_U78 = ~new_P1_U3082 | ~new_P1_U3506;
  assign new_P1_R1171_U79 = ~new_P1_U3508;
  assign new_P1_R1171_U80 = ~new_P1_U3081;
  assign new_P1_R1171_U81 = ~new_P1_U3081 | ~new_P1_U3508;
  assign new_P1_R1171_U82 = ~new_P1_U3982;
  assign new_P1_R1171_U83 = ~new_P1_U3980;
  assign new_P1_R1171_U84 = ~new_P1_U3061;
  assign new_P1_R1171_U85 = ~new_P1_U3979;
  assign new_P1_R1171_U86 = ~new_P1_U3066;
  assign new_P1_R1171_U87 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1171_U88 = ~new_P1_U3054;
  assign new_P1_R1171_U89 = ~new_P1_U3974;
  assign new_P1_R1171_U90 = ~new_P1_R1171_U305 | ~new_P1_R1171_U175;
  assign new_P1_R1171_U91 = ~new_P1_U3076;
  assign new_P1_R1171_U92 = ~new_P1_R1171_U78 | ~new_P1_R1171_U314;
  assign new_P1_R1171_U93 = ~new_P1_R1171_U260 | ~new_P1_R1171_U259;
  assign new_P1_R1171_U94 = ~new_P1_R1171_U69 | ~new_P1_R1171_U336;
  assign new_P1_R1171_U95 = ~new_P1_R1171_U456 | ~new_P1_R1171_U455;
  assign new_P1_R1171_U96 = ~new_P1_R1171_U503 | ~new_P1_R1171_U502;
  assign new_P1_R1171_U97 = ~new_P1_R1171_U374 | ~new_P1_R1171_U373;
  assign new_P1_R1171_U98 = ~new_P1_R1171_U379 | ~new_P1_R1171_U378;
  assign new_P1_R1171_U99 = ~new_P1_R1171_U386 | ~new_P1_R1171_U385;
  assign new_P1_R1171_U100 = ~new_P1_R1171_U393 | ~new_P1_R1171_U392;
  assign new_P1_R1171_U101 = ~new_P1_R1171_U398 | ~new_P1_R1171_U397;
  assign new_P1_R1171_U102 = ~new_P1_R1171_U407 | ~new_P1_R1171_U406;
  assign new_P1_R1171_U103 = ~new_P1_R1171_U414 | ~new_P1_R1171_U413;
  assign new_P1_R1171_U104 = ~new_P1_R1171_U421 | ~new_P1_R1171_U420;
  assign new_P1_R1171_U105 = ~new_P1_R1171_U428 | ~new_P1_R1171_U427;
  assign new_P1_R1171_U106 = ~new_P1_R1171_U433 | ~new_P1_R1171_U432;
  assign new_P1_R1171_U107 = ~new_P1_R1171_U440 | ~new_P1_R1171_U439;
  assign new_P1_R1171_U108 = ~new_P1_R1171_U447 | ~new_P1_R1171_U446;
  assign new_P1_R1171_U109 = ~new_P1_R1171_U461 | ~new_P1_R1171_U460;
  assign new_P1_R1171_U110 = ~new_P1_R1171_U466 | ~new_P1_R1171_U465;
  assign new_P1_R1171_U111 = ~new_P1_R1171_U473 | ~new_P1_R1171_U472;
  assign new_P1_R1171_U112 = ~new_P1_R1171_U480 | ~new_P1_R1171_U479;
  assign new_P1_R1171_U113 = ~new_P1_R1171_U487 | ~new_P1_R1171_U486;
  assign new_P1_R1171_U114 = ~new_P1_R1171_U494 | ~new_P1_R1171_U493;
  assign new_P1_R1171_U115 = ~new_P1_R1171_U499 | ~new_P1_R1171_U498;
  assign new_P1_R1171_U116 = new_P1_U3458 & new_P1_U3068;
  assign new_P1_R1171_U117 = new_P1_R1171_U188 & new_P1_R1171_U186;
  assign new_P1_R1171_U118 = new_P1_R1171_U193 & new_P1_R1171_U191;
  assign new_P1_R1171_U119 = new_P1_R1171_U200 & new_P1_R1171_U199;
  assign new_P1_R1171_U120 = new_P1_R1171_U23 & new_P1_R1171_U381 & new_P1_R1171_U380;
  assign new_P1_R1171_U121 = new_P1_R1171_U211 & new_P1_R1171_U6;
  assign new_P1_R1171_U122 = new_P1_R1171_U219 & new_P1_R1171_U217;
  assign new_P1_R1171_U123 = new_P1_R1171_U35 & new_P1_R1171_U388 & new_P1_R1171_U387;
  assign new_P1_R1171_U124 = new_P1_R1171_U225 & new_P1_R1171_U4;
  assign new_P1_R1171_U125 = new_P1_R1171_U233 & new_P1_R1171_U180;
  assign new_P1_R1171_U126 = new_P1_R1171_U203 & new_P1_R1171_U7;
  assign new_P1_R1171_U127 = new_P1_R1171_U238 & new_P1_R1171_U170;
  assign new_P1_R1171_U128 = new_P1_R1171_U249 & new_P1_R1171_U8;
  assign new_P1_R1171_U129 = new_P1_R1171_U247 & new_P1_R1171_U171;
  assign new_P1_R1171_U130 = new_P1_R1171_U267 & new_P1_R1171_U266;
  assign new_P1_R1171_U131 = new_P1_R1171_U10 & new_P1_R1171_U281;
  assign new_P1_R1171_U132 = new_P1_R1171_U284 & new_P1_R1171_U279;
  assign new_P1_R1171_U133 = new_P1_R1171_U300 & new_P1_R1171_U297;
  assign new_P1_R1171_U134 = new_P1_R1171_U367 & new_P1_R1171_U301;
  assign new_P1_R1171_U135 = new_P1_R1171_U159 & new_P1_R1171_U277;
  assign new_P1_R1171_U136 = new_P1_R1171_U81 & new_P1_R1171_U454 & new_P1_R1171_U453;
  assign new_P1_R1171_U137 = new_P1_R1171_U60 & new_P1_R1171_U468 & new_P1_R1171_U467;
  assign new_P1_R1171_U138 = new_P1_R1171_U333 & new_P1_R1171_U9;
  assign new_P1_R1171_U139 = new_P1_R1171_U171 & new_P1_R1171_U489 & new_P1_R1171_U488;
  assign new_P1_R1171_U140 = new_P1_R1171_U342 & new_P1_R1171_U8;
  assign new_P1_R1171_U141 = new_P1_R1171_U170 & new_P1_R1171_U501 & new_P1_R1171_U500;
  assign new_P1_R1171_U142 = new_P1_R1171_U349 & new_P1_R1171_U7;
  assign new_P1_R1171_U143 = ~new_P1_R1171_U119 | ~new_P1_R1171_U201;
  assign new_P1_R1171_U144 = ~new_P1_R1171_U216 | ~new_P1_R1171_U228;
  assign new_P1_R1171_U145 = ~new_P1_U3055;
  assign new_P1_R1171_U146 = ~new_P1_U3985;
  assign new_P1_R1171_U147 = new_P1_R1171_U402 & new_P1_R1171_U401;
  assign new_P1_R1171_U148 = ~new_P1_R1171_U363 | ~new_P1_R1171_U303 | ~new_P1_R1171_U168;
  assign new_P1_R1171_U149 = new_P1_R1171_U409 & new_P1_R1171_U408;
  assign new_P1_R1171_U150 = ~new_P1_R1171_U134 | ~new_P1_R1171_U369 | ~new_P1_R1171_U368;
  assign new_P1_R1171_U151 = new_P1_R1171_U416 & new_P1_R1171_U415;
  assign new_P1_R1171_U152 = ~new_P1_R1171_U87 | ~new_P1_R1171_U364 | ~new_P1_R1171_U298;
  assign new_P1_R1171_U153 = new_P1_R1171_U423 & new_P1_R1171_U422;
  assign new_P1_R1171_U154 = ~new_P1_R1171_U292 | ~new_P1_R1171_U291;
  assign new_P1_R1171_U155 = new_P1_R1171_U435 & new_P1_R1171_U434;
  assign new_P1_R1171_U156 = ~new_P1_R1171_U288 | ~new_P1_R1171_U287;
  assign new_P1_R1171_U157 = new_P1_R1171_U442 & new_P1_R1171_U441;
  assign new_P1_R1171_U158 = ~new_P1_R1171_U132 | ~new_P1_R1171_U283;
  assign new_P1_R1171_U159 = new_P1_R1171_U449 & new_P1_R1171_U448;
  assign new_P1_R1171_U160 = ~new_P1_R1171_U44 | ~new_P1_R1171_U326;
  assign new_P1_R1171_U161 = ~new_P1_R1171_U130 | ~new_P1_R1171_U268;
  assign new_P1_R1171_U162 = new_P1_R1171_U475 & new_P1_R1171_U474;
  assign new_P1_R1171_U163 = ~new_P1_R1171_U256 | ~new_P1_R1171_U255;
  assign new_P1_R1171_U164 = new_P1_R1171_U482 & new_P1_R1171_U481;
  assign new_P1_R1171_U165 = ~new_P1_R1171_U252 | ~new_P1_R1171_U251;
  assign new_P1_R1171_U166 = ~new_P1_R1171_U242 | ~new_P1_R1171_U241;
  assign new_P1_R1171_U167 = ~new_P1_R1171_U366 | ~new_P1_R1171_U365;
  assign new_P1_R1171_U168 = ~new_P1_U3054 | ~new_P1_R1171_U150;
  assign new_P1_R1171_U169 = ~new_P1_R1171_U35;
  assign new_P1_R1171_U170 = ~new_P1_U3479 | ~new_P1_U3083;
  assign new_P1_R1171_U171 = ~new_P1_U3072 | ~new_P1_U3488;
  assign new_P1_R1171_U172 = ~new_P1_U3058 | ~new_P1_U3977;
  assign new_P1_R1171_U173 = ~new_P1_R1171_U69;
  assign new_P1_R1171_U174 = ~new_P1_R1171_U78;
  assign new_P1_R1171_U175 = ~new_P1_U3065 | ~new_P1_U3978;
  assign new_P1_R1171_U176 = ~new_P1_R1171_U62;
  assign new_P1_R1171_U177 = new_P1_U3067 | new_P1_U3467;
  assign new_P1_R1171_U178 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1171_U179 = new_P1_U3461 | new_P1_U3064;
  assign new_P1_R1171_U180 = new_P1_U3458 | new_P1_U3068;
  assign new_P1_R1171_U181 = ~new_P1_R1171_U32;
  assign new_P1_R1171_U182 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1171_U183 = ~new_P1_R1171_U43;
  assign new_P1_R1171_U184 = ~new_P1_R1171_U44;
  assign new_P1_R1171_U185 = ~new_P1_R1171_U43 | ~new_P1_R1171_U44;
  assign new_P1_R1171_U186 = ~new_P1_R1171_U116 | ~new_P1_R1171_U179;
  assign new_P1_R1171_U187 = ~new_P1_R1171_U5 | ~new_P1_R1171_U185;
  assign new_P1_R1171_U188 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1171_U189 = ~new_P1_R1171_U117 | ~new_P1_R1171_U187;
  assign new_P1_R1171_U190 = ~new_P1_R1171_U36 | ~new_P1_R1171_U35;
  assign new_P1_R1171_U191 = ~new_P1_U3067 | ~new_P1_R1171_U190;
  assign new_P1_R1171_U192 = ~new_P1_R1171_U4 | ~new_P1_R1171_U189;
  assign new_P1_R1171_U193 = ~new_P1_U3467 | ~new_P1_R1171_U169;
  assign new_P1_R1171_U194 = ~new_P1_R1171_U42;
  assign new_P1_R1171_U195 = new_P1_U3070 | new_P1_U3473;
  assign new_P1_R1171_U196 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1171_U197 = ~new_P1_R1171_U23;
  assign new_P1_R1171_U198 = ~new_P1_R1171_U24 | ~new_P1_R1171_U23;
  assign new_P1_R1171_U199 = ~new_P1_U3070 | ~new_P1_R1171_U198;
  assign new_P1_R1171_U200 = ~new_P1_U3473 | ~new_P1_R1171_U197;
  assign new_P1_R1171_U201 = ~new_P1_R1171_U6 | ~new_P1_R1171_U42;
  assign new_P1_R1171_U202 = ~new_P1_R1171_U143;
  assign new_P1_R1171_U203 = new_P1_U3476 | new_P1_U3084;
  assign new_P1_R1171_U204 = ~new_P1_R1171_U203 | ~new_P1_R1171_U143;
  assign new_P1_R1171_U205 = ~new_P1_R1171_U41;
  assign new_P1_R1171_U206 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1171_U207 = new_P1_U3470 | new_P1_U3071;
  assign new_P1_R1171_U208 = ~new_P1_R1171_U207 | ~new_P1_R1171_U42;
  assign new_P1_R1171_U209 = ~new_P1_R1171_U120 | ~new_P1_R1171_U208;
  assign new_P1_R1171_U210 = ~new_P1_R1171_U194 | ~new_P1_R1171_U23;
  assign new_P1_R1171_U211 = ~new_P1_U3473 | ~new_P1_U3070;
  assign new_P1_R1171_U212 = ~new_P1_R1171_U121 | ~new_P1_R1171_U210;
  assign new_P1_R1171_U213 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1171_U214 = ~new_P1_R1171_U184 | ~new_P1_R1171_U180;
  assign new_P1_R1171_U215 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1171_U216 = ~new_P1_R1171_U46;
  assign new_P1_R1171_U217 = ~new_P1_R1171_U183 | ~new_P1_R1171_U5;
  assign new_P1_R1171_U218 = ~new_P1_R1171_U46 | ~new_P1_R1171_U179;
  assign new_P1_R1171_U219 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1171_U220 = ~new_P1_R1171_U45;
  assign new_P1_R1171_U221 = new_P1_U3464 | new_P1_U3060;
  assign new_P1_R1171_U222 = ~new_P1_R1171_U221 | ~new_P1_R1171_U45;
  assign new_P1_R1171_U223 = ~new_P1_R1171_U123 | ~new_P1_R1171_U222;
  assign new_P1_R1171_U224 = ~new_P1_R1171_U220 | ~new_P1_R1171_U35;
  assign new_P1_R1171_U225 = ~new_P1_U3467 | ~new_P1_U3067;
  assign new_P1_R1171_U226 = ~new_P1_R1171_U124 | ~new_P1_R1171_U224;
  assign new_P1_R1171_U227 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1171_U228 = ~new_P1_R1171_U183 | ~new_P1_R1171_U180;
  assign new_P1_R1171_U229 = ~new_P1_R1171_U144;
  assign new_P1_R1171_U230 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1171_U231 = ~new_P1_R1171_U43 | ~new_P1_R1171_U44 | ~new_P1_R1171_U400 | ~new_P1_R1171_U399;
  assign new_P1_R1171_U232 = ~new_P1_R1171_U44 | ~new_P1_R1171_U43;
  assign new_P1_R1171_U233 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1171_U234 = ~new_P1_R1171_U125 | ~new_P1_R1171_U232;
  assign new_P1_R1171_U235 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1171_U236 = new_P1_U3062 | new_P1_U3482;
  assign new_P1_R1171_U237 = ~new_P1_R1171_U176 | ~new_P1_R1171_U7;
  assign new_P1_R1171_U238 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1171_U239 = ~new_P1_R1171_U127 | ~new_P1_R1171_U237;
  assign new_P1_R1171_U240 = new_P1_U3482 | new_P1_U3062;
  assign new_P1_R1171_U241 = ~new_P1_R1171_U126 | ~new_P1_R1171_U143;
  assign new_P1_R1171_U242 = ~new_P1_R1171_U240 | ~new_P1_R1171_U239;
  assign new_P1_R1171_U243 = ~new_P1_R1171_U166;
  assign new_P1_R1171_U244 = new_P1_U3080 | new_P1_U3491;
  assign new_P1_R1171_U245 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1171_U246 = ~new_P1_R1171_U173 | ~new_P1_R1171_U8;
  assign new_P1_R1171_U247 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1171_U248 = ~new_P1_R1171_U129 | ~new_P1_R1171_U246;
  assign new_P1_R1171_U249 = new_P1_U3485 | new_P1_U3063;
  assign new_P1_R1171_U250 = new_P1_U3491 | new_P1_U3080;
  assign new_P1_R1171_U251 = ~new_P1_R1171_U128 | ~new_P1_R1171_U166;
  assign new_P1_R1171_U252 = ~new_P1_R1171_U250 | ~new_P1_R1171_U248;
  assign new_P1_R1171_U253 = ~new_P1_R1171_U165;
  assign new_P1_R1171_U254 = new_P1_U3494 | new_P1_U3079;
  assign new_P1_R1171_U255 = ~new_P1_R1171_U254 | ~new_P1_R1171_U165;
  assign new_P1_R1171_U256 = ~new_P1_U3079 | ~new_P1_U3494;
  assign new_P1_R1171_U257 = ~new_P1_R1171_U163;
  assign new_P1_R1171_U258 = new_P1_U3497 | new_P1_U3074;
  assign new_P1_R1171_U259 = ~new_P1_R1171_U258 | ~new_P1_R1171_U163;
  assign new_P1_R1171_U260 = ~new_P1_U3074 | ~new_P1_U3497;
  assign new_P1_R1171_U261 = ~new_P1_R1171_U93;
  assign new_P1_R1171_U262 = new_P1_U3069 | new_P1_U3503;
  assign new_P1_R1171_U263 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1171_U264 = ~new_P1_R1171_U60;
  assign new_P1_R1171_U265 = ~new_P1_R1171_U61 | ~new_P1_R1171_U60;
  assign new_P1_R1171_U266 = ~new_P1_U3069 | ~new_P1_R1171_U265;
  assign new_P1_R1171_U267 = ~new_P1_U3503 | ~new_P1_R1171_U264;
  assign new_P1_R1171_U268 = ~new_P1_R1171_U9 | ~new_P1_R1171_U93;
  assign new_P1_R1171_U269 = ~new_P1_R1171_U161;
  assign new_P1_R1171_U270 = new_P1_U3076 | new_P1_U3982;
  assign new_P1_R1171_U271 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1171_U272 = new_P1_U3075 | new_P1_U3981;
  assign new_P1_R1171_U273 = ~new_P1_R1171_U81;
  assign new_P1_R1171_U274 = ~new_P1_U3982 | ~new_P1_R1171_U273;
  assign new_P1_R1171_U275 = ~new_P1_R1171_U274 | ~new_P1_R1171_U91;
  assign new_P1_R1171_U276 = ~new_P1_R1171_U81 | ~new_P1_R1171_U82;
  assign new_P1_R1171_U277 = ~new_P1_R1171_U276 | ~new_P1_R1171_U275;
  assign new_P1_R1171_U278 = ~new_P1_R1171_U174 | ~new_P1_R1171_U10;
  assign new_P1_R1171_U279 = ~new_P1_U3075 | ~new_P1_U3981;
  assign new_P1_R1171_U280 = ~new_P1_R1171_U277 | ~new_P1_R1171_U278;
  assign new_P1_R1171_U281 = new_P1_U3506 | new_P1_U3082;
  assign new_P1_R1171_U282 = new_P1_U3981 | new_P1_U3075;
  assign new_P1_R1171_U283 = ~new_P1_R1171_U131 | ~new_P1_R1171_U272 | ~new_P1_R1171_U161;
  assign new_P1_R1171_U284 = ~new_P1_R1171_U282 | ~new_P1_R1171_U280;
  assign new_P1_R1171_U285 = ~new_P1_R1171_U158;
  assign new_P1_R1171_U286 = new_P1_U3980 | new_P1_U3061;
  assign new_P1_R1171_U287 = ~new_P1_R1171_U286 | ~new_P1_R1171_U158;
  assign new_P1_R1171_U288 = ~new_P1_U3061 | ~new_P1_U3980;
  assign new_P1_R1171_U289 = ~new_P1_R1171_U156;
  assign new_P1_R1171_U290 = new_P1_U3979 | new_P1_U3066;
  assign new_P1_R1171_U291 = ~new_P1_R1171_U290 | ~new_P1_R1171_U156;
  assign new_P1_R1171_U292 = ~new_P1_U3066 | ~new_P1_U3979;
  assign new_P1_R1171_U293 = ~new_P1_R1171_U154;
  assign new_P1_R1171_U294 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1171_U295 = ~new_P1_R1171_U175 | ~new_P1_R1171_U172;
  assign new_P1_R1171_U296 = ~new_P1_R1171_U87;
  assign new_P1_R1171_U297 = new_P1_U3978 | new_P1_U3065;
  assign new_P1_R1171_U298 = ~new_P1_R1171_U167 | ~new_P1_R1171_U154 | ~new_P1_R1171_U297;
  assign new_P1_R1171_U299 = ~new_P1_R1171_U152;
  assign new_P1_R1171_U300 = new_P1_U3975 | new_P1_U3053;
  assign new_P1_R1171_U301 = ~new_P1_U3053 | ~new_P1_U3975;
  assign new_P1_R1171_U302 = ~new_P1_R1171_U150;
  assign new_P1_R1171_U303 = ~new_P1_U3974 | ~new_P1_R1171_U150;
  assign new_P1_R1171_U304 = ~new_P1_R1171_U148;
  assign new_P1_R1171_U305 = ~new_P1_R1171_U297 | ~new_P1_R1171_U154;
  assign new_P1_R1171_U306 = ~new_P1_R1171_U90;
  assign new_P1_R1171_U307 = new_P1_U3977 | new_P1_U3058;
  assign new_P1_R1171_U308 = ~new_P1_R1171_U307 | ~new_P1_R1171_U90;
  assign new_P1_R1171_U309 = ~new_P1_R1171_U153 | ~new_P1_R1171_U308 | ~new_P1_R1171_U172;
  assign new_P1_R1171_U310 = ~new_P1_R1171_U306 | ~new_P1_R1171_U172;
  assign new_P1_R1171_U311 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1171_U312 = ~new_P1_R1171_U167 | ~new_P1_R1171_U310 | ~new_P1_R1171_U311;
  assign new_P1_R1171_U313 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1171_U314 = ~new_P1_R1171_U281 | ~new_P1_R1171_U161;
  assign new_P1_R1171_U315 = ~new_P1_R1171_U92;
  assign new_P1_R1171_U316 = ~new_P1_R1171_U10 | ~new_P1_R1171_U92;
  assign new_P1_R1171_U317 = ~new_P1_R1171_U135 | ~new_P1_R1171_U316;
  assign new_P1_R1171_U318 = ~new_P1_R1171_U316 | ~new_P1_R1171_U277;
  assign new_P1_R1171_U319 = ~new_P1_R1171_U452 | ~new_P1_R1171_U318;
  assign new_P1_R1171_U320 = new_P1_U3508 | new_P1_U3081;
  assign new_P1_R1171_U321 = ~new_P1_R1171_U320 | ~new_P1_R1171_U92;
  assign new_P1_R1171_U322 = ~new_P1_R1171_U136 | ~new_P1_R1171_U321;
  assign new_P1_R1171_U323 = ~new_P1_R1171_U315 | ~new_P1_R1171_U81;
  assign new_P1_R1171_U324 = ~new_P1_U3076 | ~new_P1_U3982;
  assign new_P1_R1171_U325 = ~new_P1_R1171_U10 | ~new_P1_R1171_U324 | ~new_P1_R1171_U323;
  assign new_P1_R1171_U326 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1171_U327 = ~new_P1_R1171_U160;
  assign new_P1_R1171_U328 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1171_U329 = new_P1_U3500 | new_P1_U3073;
  assign new_P1_R1171_U330 = ~new_P1_R1171_U329 | ~new_P1_R1171_U93;
  assign new_P1_R1171_U331 = ~new_P1_R1171_U137 | ~new_P1_R1171_U330;
  assign new_P1_R1171_U332 = ~new_P1_R1171_U261 | ~new_P1_R1171_U60;
  assign new_P1_R1171_U333 = ~new_P1_U3503 | ~new_P1_U3069;
  assign new_P1_R1171_U334 = ~new_P1_R1171_U138 | ~new_P1_R1171_U332;
  assign new_P1_R1171_U335 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1171_U336 = ~new_P1_R1171_U249 | ~new_P1_R1171_U166;
  assign new_P1_R1171_U337 = ~new_P1_R1171_U94;
  assign new_P1_R1171_U338 = new_P1_U3488 | new_P1_U3072;
  assign new_P1_R1171_U339 = ~new_P1_R1171_U338 | ~new_P1_R1171_U94;
  assign new_P1_R1171_U340 = ~new_P1_R1171_U139 | ~new_P1_R1171_U339;
  assign new_P1_R1171_U341 = ~new_P1_R1171_U337 | ~new_P1_R1171_U171;
  assign new_P1_R1171_U342 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1171_U343 = ~new_P1_R1171_U140 | ~new_P1_R1171_U341;
  assign new_P1_R1171_U344 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1171_U345 = new_P1_U3479 | new_P1_U3083;
  assign new_P1_R1171_U346 = ~new_P1_R1171_U345 | ~new_P1_R1171_U41;
  assign new_P1_R1171_U347 = ~new_P1_R1171_U141 | ~new_P1_R1171_U346;
  assign new_P1_R1171_U348 = ~new_P1_R1171_U205 | ~new_P1_R1171_U170;
  assign new_P1_R1171_U349 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1171_U350 = ~new_P1_R1171_U142 | ~new_P1_R1171_U348;
  assign new_P1_R1171_U351 = ~new_P1_R1171_U206 | ~new_P1_R1171_U170;
  assign new_P1_R1171_U352 = ~new_P1_R1171_U203 | ~new_P1_R1171_U62;
  assign new_P1_R1171_U353 = ~new_P1_R1171_U213 | ~new_P1_R1171_U23;
  assign new_P1_R1171_U354 = ~new_P1_R1171_U227 | ~new_P1_R1171_U35;
  assign new_P1_R1171_U355 = ~new_P1_R1171_U230 | ~new_P1_R1171_U179;
  assign new_P1_R1171_U356 = ~new_P1_R1171_U313 | ~new_P1_R1171_U172;
  assign new_P1_R1171_U357 = ~new_P1_R1171_U297 | ~new_P1_R1171_U175;
  assign new_P1_R1171_U358 = ~new_P1_R1171_U328 | ~new_P1_R1171_U81;
  assign new_P1_R1171_U359 = ~new_P1_R1171_U281 | ~new_P1_R1171_U78;
  assign new_P1_R1171_U360 = ~new_P1_R1171_U335 | ~new_P1_R1171_U60;
  assign new_P1_R1171_U361 = ~new_P1_R1171_U344 | ~new_P1_R1171_U171;
  assign new_P1_R1171_U362 = ~new_P1_R1171_U249 | ~new_P1_R1171_U69;
  assign new_P1_R1171_U363 = ~new_P1_U3974 | ~new_P1_U3054;
  assign new_P1_R1171_U364 = ~new_P1_R1171_U295 | ~new_P1_R1171_U167;
  assign new_P1_R1171_U365 = ~new_P1_U3057 | ~new_P1_R1171_U294;
  assign new_P1_R1171_U366 = ~new_P1_U3976 | ~new_P1_R1171_U294;
  assign new_P1_R1171_U367 = ~new_P1_R1171_U300 | ~new_P1_R1171_U295 | ~new_P1_R1171_U167;
  assign new_P1_R1171_U368 = ~new_P1_R1171_U133 | ~new_P1_R1171_U154 | ~new_P1_R1171_U167;
  assign new_P1_R1171_U369 = ~new_P1_R1171_U296 | ~new_P1_R1171_U300;
  assign new_P1_R1171_U370 = ~new_P1_U3083 | ~new_P1_R1171_U40;
  assign new_P1_R1171_U371 = ~new_P1_U3479 | ~new_P1_R1171_U39;
  assign new_P1_R1171_U372 = ~new_P1_R1171_U371 | ~new_P1_R1171_U370;
  assign new_P1_R1171_U373 = ~new_P1_R1171_U351 | ~new_P1_R1171_U41;
  assign new_P1_R1171_U374 = ~new_P1_R1171_U372 | ~new_P1_R1171_U205;
  assign new_P1_R1171_U375 = ~new_P1_U3084 | ~new_P1_R1171_U37;
  assign new_P1_R1171_U376 = ~new_P1_U3476 | ~new_P1_R1171_U38;
  assign new_P1_R1171_U377 = ~new_P1_R1171_U376 | ~new_P1_R1171_U375;
  assign new_P1_R1171_U378 = ~new_P1_R1171_U352 | ~new_P1_R1171_U143;
  assign new_P1_R1171_U379 = ~new_P1_R1171_U202 | ~new_P1_R1171_U377;
  assign new_P1_R1171_U380 = ~new_P1_U3070 | ~new_P1_R1171_U24;
  assign new_P1_R1171_U381 = ~new_P1_U3473 | ~new_P1_R1171_U22;
  assign new_P1_R1171_U382 = ~new_P1_U3071 | ~new_P1_R1171_U20;
  assign new_P1_R1171_U383 = ~new_P1_U3470 | ~new_P1_R1171_U21;
  assign new_P1_R1171_U384 = ~new_P1_R1171_U383 | ~new_P1_R1171_U382;
  assign new_P1_R1171_U385 = ~new_P1_R1171_U353 | ~new_P1_R1171_U42;
  assign new_P1_R1171_U386 = ~new_P1_R1171_U384 | ~new_P1_R1171_U194;
  assign new_P1_R1171_U387 = ~new_P1_U3067 | ~new_P1_R1171_U36;
  assign new_P1_R1171_U388 = ~new_P1_U3467 | ~new_P1_R1171_U27;
  assign new_P1_R1171_U389 = ~new_P1_U3060 | ~new_P1_R1171_U25;
  assign new_P1_R1171_U390 = ~new_P1_U3464 | ~new_P1_R1171_U26;
  assign new_P1_R1171_U391 = ~new_P1_R1171_U390 | ~new_P1_R1171_U389;
  assign new_P1_R1171_U392 = ~new_P1_R1171_U354 | ~new_P1_R1171_U45;
  assign new_P1_R1171_U393 = ~new_P1_R1171_U391 | ~new_P1_R1171_U220;
  assign new_P1_R1171_U394 = ~new_P1_U3064 | ~new_P1_R1171_U33;
  assign new_P1_R1171_U395 = ~new_P1_U3461 | ~new_P1_R1171_U34;
  assign new_P1_R1171_U396 = ~new_P1_R1171_U395 | ~new_P1_R1171_U394;
  assign new_P1_R1171_U397 = ~new_P1_R1171_U355 | ~new_P1_R1171_U144;
  assign new_P1_R1171_U398 = ~new_P1_R1171_U229 | ~new_P1_R1171_U396;
  assign new_P1_R1171_U399 = ~new_P1_U3068 | ~new_P1_R1171_U28;
  assign new_P1_R1171_U400 = ~new_P1_U3458 | ~new_P1_R1171_U29;
  assign new_P1_R1171_U401 = ~new_P1_U3055 | ~new_P1_R1171_U146;
  assign new_P1_R1171_U402 = ~new_P1_U3985 | ~new_P1_R1171_U145;
  assign new_P1_R1171_U403 = ~new_P1_U3055 | ~new_P1_R1171_U146;
  assign new_P1_R1171_U404 = ~new_P1_U3985 | ~new_P1_R1171_U145;
  assign new_P1_R1171_U405 = ~new_P1_R1171_U404 | ~new_P1_R1171_U403;
  assign new_P1_R1171_U406 = ~new_P1_R1171_U147 | ~new_P1_R1171_U148;
  assign new_P1_R1171_U407 = ~new_P1_R1171_U304 | ~new_P1_R1171_U405;
  assign new_P1_R1171_U408 = ~new_P1_U3054 | ~new_P1_R1171_U89;
  assign new_P1_R1171_U409 = ~new_P1_U3974 | ~new_P1_R1171_U88;
  assign new_P1_R1171_U410 = ~new_P1_U3054 | ~new_P1_R1171_U89;
  assign new_P1_R1171_U411 = ~new_P1_U3974 | ~new_P1_R1171_U88;
  assign new_P1_R1171_U412 = ~new_P1_R1171_U411 | ~new_P1_R1171_U410;
  assign new_P1_R1171_U413 = ~new_P1_R1171_U149 | ~new_P1_R1171_U150;
  assign new_P1_R1171_U414 = ~new_P1_R1171_U302 | ~new_P1_R1171_U412;
  assign new_P1_R1171_U415 = ~new_P1_U3053 | ~new_P1_R1171_U47;
  assign new_P1_R1171_U416 = ~new_P1_U3975 | ~new_P1_R1171_U48;
  assign new_P1_R1171_U417 = ~new_P1_U3053 | ~new_P1_R1171_U47;
  assign new_P1_R1171_U418 = ~new_P1_U3975 | ~new_P1_R1171_U48;
  assign new_P1_R1171_U419 = ~new_P1_R1171_U418 | ~new_P1_R1171_U417;
  assign new_P1_R1171_U420 = ~new_P1_R1171_U151 | ~new_P1_R1171_U152;
  assign new_P1_R1171_U421 = ~new_P1_R1171_U299 | ~new_P1_R1171_U419;
  assign new_P1_R1171_U422 = ~new_P1_U3057 | ~new_P1_R1171_U50;
  assign new_P1_R1171_U423 = ~new_P1_U3976 | ~new_P1_R1171_U49;
  assign new_P1_R1171_U424 = ~new_P1_U3058 | ~new_P1_R1171_U51;
  assign new_P1_R1171_U425 = ~new_P1_U3977 | ~new_P1_R1171_U52;
  assign new_P1_R1171_U426 = ~new_P1_R1171_U425 | ~new_P1_R1171_U424;
  assign new_P1_R1171_U427 = ~new_P1_R1171_U356 | ~new_P1_R1171_U90;
  assign new_P1_R1171_U428 = ~new_P1_R1171_U426 | ~new_P1_R1171_U306;
  assign new_P1_R1171_U429 = ~new_P1_U3065 | ~new_P1_R1171_U53;
  assign new_P1_R1171_U430 = ~new_P1_U3978 | ~new_P1_R1171_U54;
  assign new_P1_R1171_U431 = ~new_P1_R1171_U430 | ~new_P1_R1171_U429;
  assign new_P1_R1171_U432 = ~new_P1_R1171_U357 | ~new_P1_R1171_U154;
  assign new_P1_R1171_U433 = ~new_P1_R1171_U293 | ~new_P1_R1171_U431;
  assign new_P1_R1171_U434 = ~new_P1_U3066 | ~new_P1_R1171_U85;
  assign new_P1_R1171_U435 = ~new_P1_U3979 | ~new_P1_R1171_U86;
  assign new_P1_R1171_U436 = ~new_P1_U3066 | ~new_P1_R1171_U85;
  assign new_P1_R1171_U437 = ~new_P1_U3979 | ~new_P1_R1171_U86;
  assign new_P1_R1171_U438 = ~new_P1_R1171_U437 | ~new_P1_R1171_U436;
  assign new_P1_R1171_U439 = ~new_P1_R1171_U155 | ~new_P1_R1171_U156;
  assign new_P1_R1171_U440 = ~new_P1_R1171_U289 | ~new_P1_R1171_U438;
  assign new_P1_R1171_U441 = ~new_P1_U3061 | ~new_P1_R1171_U83;
  assign new_P1_R1171_U442 = ~new_P1_U3980 | ~new_P1_R1171_U84;
  assign new_P1_R1171_U443 = ~new_P1_U3061 | ~new_P1_R1171_U83;
  assign new_P1_R1171_U444 = ~new_P1_U3980 | ~new_P1_R1171_U84;
  assign new_P1_R1171_U445 = ~new_P1_R1171_U444 | ~new_P1_R1171_U443;
  assign new_P1_R1171_U446 = ~new_P1_R1171_U157 | ~new_P1_R1171_U158;
  assign new_P1_R1171_U447 = ~new_P1_R1171_U285 | ~new_P1_R1171_U445;
  assign new_P1_R1171_U448 = ~new_P1_U3075 | ~new_P1_R1171_U55;
  assign new_P1_R1171_U449 = ~new_P1_U3981 | ~new_P1_R1171_U56;
  assign new_P1_R1171_U450 = ~new_P1_U3075 | ~new_P1_R1171_U55;
  assign new_P1_R1171_U451 = ~new_P1_U3981 | ~new_P1_R1171_U56;
  assign new_P1_R1171_U452 = ~new_P1_R1171_U451 | ~new_P1_R1171_U450;
  assign new_P1_R1171_U453 = ~new_P1_U3076 | ~new_P1_R1171_U82;
  assign new_P1_R1171_U454 = ~new_P1_U3982 | ~new_P1_R1171_U91;
  assign new_P1_R1171_U455 = ~new_P1_R1171_U181 | ~new_P1_R1171_U160;
  assign new_P1_R1171_U456 = ~new_P1_R1171_U327 | ~new_P1_R1171_U32;
  assign new_P1_R1171_U457 = ~new_P1_U3081 | ~new_P1_R1171_U79;
  assign new_P1_R1171_U458 = ~new_P1_U3508 | ~new_P1_R1171_U80;
  assign new_P1_R1171_U459 = ~new_P1_R1171_U458 | ~new_P1_R1171_U457;
  assign new_P1_R1171_U460 = ~new_P1_R1171_U358 | ~new_P1_R1171_U92;
  assign new_P1_R1171_U461 = ~new_P1_R1171_U459 | ~new_P1_R1171_U315;
  assign new_P1_R1171_U462 = ~new_P1_U3082 | ~new_P1_R1171_U76;
  assign new_P1_R1171_U463 = ~new_P1_U3506 | ~new_P1_R1171_U77;
  assign new_P1_R1171_U464 = ~new_P1_R1171_U463 | ~new_P1_R1171_U462;
  assign new_P1_R1171_U465 = ~new_P1_R1171_U359 | ~new_P1_R1171_U161;
  assign new_P1_R1171_U466 = ~new_P1_R1171_U269 | ~new_P1_R1171_U464;
  assign new_P1_R1171_U467 = ~new_P1_U3069 | ~new_P1_R1171_U61;
  assign new_P1_R1171_U468 = ~new_P1_U3503 | ~new_P1_R1171_U59;
  assign new_P1_R1171_U469 = ~new_P1_U3073 | ~new_P1_R1171_U57;
  assign new_P1_R1171_U470 = ~new_P1_U3500 | ~new_P1_R1171_U58;
  assign new_P1_R1171_U471 = ~new_P1_R1171_U470 | ~new_P1_R1171_U469;
  assign new_P1_R1171_U472 = ~new_P1_R1171_U360 | ~new_P1_R1171_U93;
  assign new_P1_R1171_U473 = ~new_P1_R1171_U471 | ~new_P1_R1171_U261;
  assign new_P1_R1171_U474 = ~new_P1_U3074 | ~new_P1_R1171_U74;
  assign new_P1_R1171_U475 = ~new_P1_U3497 | ~new_P1_R1171_U75;
  assign new_P1_R1171_U476 = ~new_P1_U3074 | ~new_P1_R1171_U74;
  assign new_P1_R1171_U477 = ~new_P1_U3497 | ~new_P1_R1171_U75;
  assign new_P1_R1171_U478 = ~new_P1_R1171_U477 | ~new_P1_R1171_U476;
  assign new_P1_R1171_U479 = ~new_P1_R1171_U162 | ~new_P1_R1171_U163;
  assign new_P1_R1171_U480 = ~new_P1_R1171_U257 | ~new_P1_R1171_U478;
  assign new_P1_R1171_U481 = ~new_P1_U3079 | ~new_P1_R1171_U72;
  assign new_P1_R1171_U482 = ~new_P1_U3494 | ~new_P1_R1171_U73;
  assign new_P1_R1171_U483 = ~new_P1_U3079 | ~new_P1_R1171_U72;
  assign new_P1_R1171_U484 = ~new_P1_U3494 | ~new_P1_R1171_U73;
  assign new_P1_R1171_U485 = ~new_P1_R1171_U484 | ~new_P1_R1171_U483;
  assign new_P1_R1171_U486 = ~new_P1_R1171_U164 | ~new_P1_R1171_U165;
  assign new_P1_R1171_U487 = ~new_P1_R1171_U253 | ~new_P1_R1171_U485;
  assign new_P1_R1171_U488 = ~new_P1_U3080 | ~new_P1_R1171_U70;
  assign new_P1_R1171_U489 = ~new_P1_U3491 | ~new_P1_R1171_U71;
  assign new_P1_R1171_U490 = ~new_P1_U3072 | ~new_P1_R1171_U65;
  assign new_P1_R1171_U491 = ~new_P1_U3488 | ~new_P1_R1171_U66;
  assign new_P1_R1171_U492 = ~new_P1_R1171_U491 | ~new_P1_R1171_U490;
  assign new_P1_R1171_U493 = ~new_P1_R1171_U361 | ~new_P1_R1171_U94;
  assign new_P1_R1171_U494 = ~new_P1_R1171_U492 | ~new_P1_R1171_U337;
  assign new_P1_R1171_U495 = ~new_P1_U3063 | ~new_P1_R1171_U67;
  assign new_P1_R1171_U496 = ~new_P1_U3485 | ~new_P1_R1171_U68;
  assign new_P1_R1171_U497 = ~new_P1_R1171_U496 | ~new_P1_R1171_U495;
  assign new_P1_R1171_U498 = ~new_P1_R1171_U362 | ~new_P1_R1171_U166;
  assign new_P1_R1171_U499 = ~new_P1_R1171_U243 | ~new_P1_R1171_U497;
  assign new_P1_R1171_U500 = ~new_P1_U3062 | ~new_P1_R1171_U63;
  assign new_P1_R1171_U501 = ~new_P1_U3482 | ~new_P1_R1171_U64;
  assign new_P1_R1171_U502 = ~new_P1_U3077 | ~new_P1_R1171_U30;
  assign new_P1_R1171_U503 = ~new_P1_U3450 | ~new_P1_R1171_U31;
  assign new_P1_R1138_U4 = new_P1_R1138_U178 & new_P1_R1138_U177;
  assign new_P1_R1138_U5 = new_P1_R1138_U179 & new_P1_R1138_U180;
  assign new_P1_R1138_U6 = new_P1_R1138_U196 & new_P1_R1138_U195;
  assign new_P1_R1138_U7 = new_P1_R1138_U236 & new_P1_R1138_U235;
  assign new_P1_R1138_U8 = new_P1_R1138_U245 & new_P1_R1138_U244;
  assign new_P1_R1138_U9 = new_P1_R1138_U263 & new_P1_R1138_U262;
  assign new_P1_R1138_U10 = new_P1_R1138_U271 & new_P1_R1138_U270;
  assign new_P1_R1138_U11 = new_P1_R1138_U350 & new_P1_R1138_U347;
  assign new_P1_R1138_U12 = new_P1_R1138_U343 & new_P1_R1138_U340;
  assign new_P1_R1138_U13 = new_P1_R1138_U334 & new_P1_R1138_U331;
  assign new_P1_R1138_U14 = new_P1_R1138_U325 & new_P1_R1138_U322;
  assign new_P1_R1138_U15 = new_P1_R1138_U319 & new_P1_R1138_U317;
  assign new_P1_R1138_U16 = new_P1_R1138_U312 & new_P1_R1138_U309;
  assign new_P1_R1138_U17 = new_P1_R1138_U234 & new_P1_R1138_U231;
  assign new_P1_R1138_U18 = new_P1_R1138_U226 & new_P1_R1138_U223;
  assign new_P1_R1138_U19 = new_P1_R1138_U212 & new_P1_R1138_U209;
  assign new_P1_R1138_U20 = ~new_P1_U3470;
  assign new_P1_R1138_U21 = ~new_P1_U3071;
  assign new_P1_R1138_U22 = ~new_P1_U3070;
  assign new_P1_R1138_U23 = ~new_P1_U3071 | ~new_P1_U3470;
  assign new_P1_R1138_U24 = ~new_P1_U3473;
  assign new_P1_R1138_U25 = ~new_P1_U3464;
  assign new_P1_R1138_U26 = ~new_P1_U3060;
  assign new_P1_R1138_U27 = ~new_P1_U3067;
  assign new_P1_R1138_U28 = ~new_P1_U3458;
  assign new_P1_R1138_U29 = ~new_P1_U3068;
  assign new_P1_R1138_U30 = ~new_P1_U3450;
  assign new_P1_R1138_U31 = ~new_P1_U3077;
  assign new_P1_R1138_U32 = ~new_P1_U3077 | ~new_P1_U3450;
  assign new_P1_R1138_U33 = ~new_P1_U3461;
  assign new_P1_R1138_U34 = ~new_P1_U3064;
  assign new_P1_R1138_U35 = ~new_P1_U3060 | ~new_P1_U3464;
  assign new_P1_R1138_U36 = ~new_P1_U3467;
  assign new_P1_R1138_U37 = ~new_P1_U3476;
  assign new_P1_R1138_U38 = ~new_P1_U3084;
  assign new_P1_R1138_U39 = ~new_P1_U3083;
  assign new_P1_R1138_U40 = ~new_P1_U3479;
  assign new_P1_R1138_U41 = ~new_P1_R1138_U62 | ~new_P1_R1138_U204;
  assign new_P1_R1138_U42 = ~new_P1_R1138_U118 | ~new_P1_R1138_U192;
  assign new_P1_R1138_U43 = ~new_P1_R1138_U181 | ~new_P1_R1138_U182;
  assign new_P1_R1138_U44 = ~new_P1_U3455 | ~new_P1_U3078;
  assign new_P1_R1138_U45 = ~new_P1_R1138_U122 | ~new_P1_R1138_U218;
  assign new_P1_R1138_U46 = ~new_P1_R1138_U215 | ~new_P1_R1138_U214;
  assign new_P1_R1138_U47 = ~new_P1_U3975;
  assign new_P1_R1138_U48 = ~new_P1_U3053;
  assign new_P1_R1138_U49 = ~new_P1_U3057;
  assign new_P1_R1138_U50 = ~new_P1_U3976;
  assign new_P1_R1138_U51 = ~new_P1_U3977;
  assign new_P1_R1138_U52 = ~new_P1_U3058;
  assign new_P1_R1138_U53 = ~new_P1_U3978;
  assign new_P1_R1138_U54 = ~new_P1_U3065;
  assign new_P1_R1138_U55 = ~new_P1_U3981;
  assign new_P1_R1138_U56 = ~new_P1_U3075;
  assign new_P1_R1138_U57 = ~new_P1_U3500;
  assign new_P1_R1138_U58 = ~new_P1_U3073;
  assign new_P1_R1138_U59 = ~new_P1_U3069;
  assign new_P1_R1138_U60 = ~new_P1_U3073 | ~new_P1_U3500;
  assign new_P1_R1138_U61 = ~new_P1_U3503;
  assign new_P1_R1138_U62 = ~new_P1_U3084 | ~new_P1_U3476;
  assign new_P1_R1138_U63 = ~new_P1_U3482;
  assign new_P1_R1138_U64 = ~new_P1_U3062;
  assign new_P1_R1138_U65 = ~new_P1_U3488;
  assign new_P1_R1138_U66 = ~new_P1_U3072;
  assign new_P1_R1138_U67 = ~new_P1_U3485;
  assign new_P1_R1138_U68 = ~new_P1_U3063;
  assign new_P1_R1138_U69 = ~new_P1_U3063 | ~new_P1_U3485;
  assign new_P1_R1138_U70 = ~new_P1_U3491;
  assign new_P1_R1138_U71 = ~new_P1_U3080;
  assign new_P1_R1138_U72 = ~new_P1_U3494;
  assign new_P1_R1138_U73 = ~new_P1_U3079;
  assign new_P1_R1138_U74 = ~new_P1_U3497;
  assign new_P1_R1138_U75 = ~new_P1_U3074;
  assign new_P1_R1138_U76 = ~new_P1_U3506;
  assign new_P1_R1138_U77 = ~new_P1_U3082;
  assign new_P1_R1138_U78 = ~new_P1_U3082 | ~new_P1_U3506;
  assign new_P1_R1138_U79 = ~new_P1_U3508;
  assign new_P1_R1138_U80 = ~new_P1_U3081;
  assign new_P1_R1138_U81 = ~new_P1_U3081 | ~new_P1_U3508;
  assign new_P1_R1138_U82 = ~new_P1_U3982;
  assign new_P1_R1138_U83 = ~new_P1_U3980;
  assign new_P1_R1138_U84 = ~new_P1_U3061;
  assign new_P1_R1138_U85 = ~new_P1_U3979;
  assign new_P1_R1138_U86 = ~new_P1_U3066;
  assign new_P1_R1138_U87 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1138_U88 = ~new_P1_U3054;
  assign new_P1_R1138_U89 = ~new_P1_U3974;
  assign new_P1_R1138_U90 = ~new_P1_R1138_U305 | ~new_P1_R1138_U175;
  assign new_P1_R1138_U91 = ~new_P1_U3076;
  assign new_P1_R1138_U92 = ~new_P1_R1138_U78 | ~new_P1_R1138_U314;
  assign new_P1_R1138_U93 = ~new_P1_R1138_U260 | ~new_P1_R1138_U259;
  assign new_P1_R1138_U94 = ~new_P1_R1138_U69 | ~new_P1_R1138_U336;
  assign new_P1_R1138_U95 = ~new_P1_R1138_U456 | ~new_P1_R1138_U455;
  assign new_P1_R1138_U96 = ~new_P1_R1138_U503 | ~new_P1_R1138_U502;
  assign new_P1_R1138_U97 = ~new_P1_R1138_U374 | ~new_P1_R1138_U373;
  assign new_P1_R1138_U98 = ~new_P1_R1138_U379 | ~new_P1_R1138_U378;
  assign new_P1_R1138_U99 = ~new_P1_R1138_U386 | ~new_P1_R1138_U385;
  assign new_P1_R1138_U100 = ~new_P1_R1138_U393 | ~new_P1_R1138_U392;
  assign new_P1_R1138_U101 = ~new_P1_R1138_U398 | ~new_P1_R1138_U397;
  assign new_P1_R1138_U102 = ~new_P1_R1138_U407 | ~new_P1_R1138_U406;
  assign new_P1_R1138_U103 = ~new_P1_R1138_U414 | ~new_P1_R1138_U413;
  assign new_P1_R1138_U104 = ~new_P1_R1138_U421 | ~new_P1_R1138_U420;
  assign new_P1_R1138_U105 = ~new_P1_R1138_U428 | ~new_P1_R1138_U427;
  assign new_P1_R1138_U106 = ~new_P1_R1138_U433 | ~new_P1_R1138_U432;
  assign new_P1_R1138_U107 = ~new_P1_R1138_U440 | ~new_P1_R1138_U439;
  assign new_P1_R1138_U108 = ~new_P1_R1138_U447 | ~new_P1_R1138_U446;
  assign new_P1_R1138_U109 = ~new_P1_R1138_U461 | ~new_P1_R1138_U460;
  assign new_P1_R1138_U110 = ~new_P1_R1138_U466 | ~new_P1_R1138_U465;
  assign new_P1_R1138_U111 = ~new_P1_R1138_U473 | ~new_P1_R1138_U472;
  assign new_P1_R1138_U112 = ~new_P1_R1138_U480 | ~new_P1_R1138_U479;
  assign new_P1_R1138_U113 = ~new_P1_R1138_U487 | ~new_P1_R1138_U486;
  assign new_P1_R1138_U114 = ~new_P1_R1138_U494 | ~new_P1_R1138_U493;
  assign new_P1_R1138_U115 = ~new_P1_R1138_U499 | ~new_P1_R1138_U498;
  assign new_P1_R1138_U116 = new_P1_U3458 & new_P1_U3068;
  assign new_P1_R1138_U117 = new_P1_R1138_U188 & new_P1_R1138_U186;
  assign new_P1_R1138_U118 = new_P1_R1138_U193 & new_P1_R1138_U191;
  assign new_P1_R1138_U119 = new_P1_R1138_U200 & new_P1_R1138_U199;
  assign new_P1_R1138_U120 = new_P1_R1138_U23 & new_P1_R1138_U381 & new_P1_R1138_U380;
  assign new_P1_R1138_U121 = new_P1_R1138_U211 & new_P1_R1138_U6;
  assign new_P1_R1138_U122 = new_P1_R1138_U219 & new_P1_R1138_U217;
  assign new_P1_R1138_U123 = new_P1_R1138_U35 & new_P1_R1138_U388 & new_P1_R1138_U387;
  assign new_P1_R1138_U124 = new_P1_R1138_U225 & new_P1_R1138_U4;
  assign new_P1_R1138_U125 = new_P1_R1138_U233 & new_P1_R1138_U180;
  assign new_P1_R1138_U126 = new_P1_R1138_U203 & new_P1_R1138_U7;
  assign new_P1_R1138_U127 = new_P1_R1138_U238 & new_P1_R1138_U170;
  assign new_P1_R1138_U128 = new_P1_R1138_U249 & new_P1_R1138_U8;
  assign new_P1_R1138_U129 = new_P1_R1138_U247 & new_P1_R1138_U171;
  assign new_P1_R1138_U130 = new_P1_R1138_U267 & new_P1_R1138_U266;
  assign new_P1_R1138_U131 = new_P1_R1138_U10 & new_P1_R1138_U281;
  assign new_P1_R1138_U132 = new_P1_R1138_U284 & new_P1_R1138_U279;
  assign new_P1_R1138_U133 = new_P1_R1138_U300 & new_P1_R1138_U297;
  assign new_P1_R1138_U134 = new_P1_R1138_U367 & new_P1_R1138_U301;
  assign new_P1_R1138_U135 = new_P1_R1138_U159 & new_P1_R1138_U277;
  assign new_P1_R1138_U136 = new_P1_R1138_U81 & new_P1_R1138_U454 & new_P1_R1138_U453;
  assign new_P1_R1138_U137 = new_P1_R1138_U60 & new_P1_R1138_U468 & new_P1_R1138_U467;
  assign new_P1_R1138_U138 = new_P1_R1138_U333 & new_P1_R1138_U9;
  assign new_P1_R1138_U139 = new_P1_R1138_U171 & new_P1_R1138_U489 & new_P1_R1138_U488;
  assign new_P1_R1138_U140 = new_P1_R1138_U342 & new_P1_R1138_U8;
  assign new_P1_R1138_U141 = new_P1_R1138_U170 & new_P1_R1138_U501 & new_P1_R1138_U500;
  assign new_P1_R1138_U142 = new_P1_R1138_U349 & new_P1_R1138_U7;
  assign new_P1_R1138_U143 = ~new_P1_R1138_U119 | ~new_P1_R1138_U201;
  assign new_P1_R1138_U144 = ~new_P1_R1138_U216 | ~new_P1_R1138_U228;
  assign new_P1_R1138_U145 = ~new_P1_U3055;
  assign new_P1_R1138_U146 = ~new_P1_U3985;
  assign new_P1_R1138_U147 = new_P1_R1138_U402 & new_P1_R1138_U401;
  assign new_P1_R1138_U148 = ~new_P1_R1138_U363 | ~new_P1_R1138_U303 | ~new_P1_R1138_U168;
  assign new_P1_R1138_U149 = new_P1_R1138_U409 & new_P1_R1138_U408;
  assign new_P1_R1138_U150 = ~new_P1_R1138_U134 | ~new_P1_R1138_U369 | ~new_P1_R1138_U368;
  assign new_P1_R1138_U151 = new_P1_R1138_U416 & new_P1_R1138_U415;
  assign new_P1_R1138_U152 = ~new_P1_R1138_U87 | ~new_P1_R1138_U364 | ~new_P1_R1138_U298;
  assign new_P1_R1138_U153 = new_P1_R1138_U423 & new_P1_R1138_U422;
  assign new_P1_R1138_U154 = ~new_P1_R1138_U292 | ~new_P1_R1138_U291;
  assign new_P1_R1138_U155 = new_P1_R1138_U435 & new_P1_R1138_U434;
  assign new_P1_R1138_U156 = ~new_P1_R1138_U288 | ~new_P1_R1138_U287;
  assign new_P1_R1138_U157 = new_P1_R1138_U442 & new_P1_R1138_U441;
  assign new_P1_R1138_U158 = ~new_P1_R1138_U132 | ~new_P1_R1138_U283;
  assign new_P1_R1138_U159 = new_P1_R1138_U449 & new_P1_R1138_U448;
  assign new_P1_R1138_U160 = ~new_P1_R1138_U44 | ~new_P1_R1138_U326;
  assign new_P1_R1138_U161 = ~new_P1_R1138_U130 | ~new_P1_R1138_U268;
  assign new_P1_R1138_U162 = new_P1_R1138_U475 & new_P1_R1138_U474;
  assign new_P1_R1138_U163 = ~new_P1_R1138_U256 | ~new_P1_R1138_U255;
  assign new_P1_R1138_U164 = new_P1_R1138_U482 & new_P1_R1138_U481;
  assign new_P1_R1138_U165 = ~new_P1_R1138_U252 | ~new_P1_R1138_U251;
  assign new_P1_R1138_U166 = ~new_P1_R1138_U242 | ~new_P1_R1138_U241;
  assign new_P1_R1138_U167 = ~new_P1_R1138_U366 | ~new_P1_R1138_U365;
  assign new_P1_R1138_U168 = ~new_P1_U3054 | ~new_P1_R1138_U150;
  assign new_P1_R1138_U169 = ~new_P1_R1138_U35;
  assign new_P1_R1138_U170 = ~new_P1_U3479 | ~new_P1_U3083;
  assign new_P1_R1138_U171 = ~new_P1_U3072 | ~new_P1_U3488;
  assign new_P1_R1138_U172 = ~new_P1_U3058 | ~new_P1_U3977;
  assign new_P1_R1138_U173 = ~new_P1_R1138_U69;
  assign new_P1_R1138_U174 = ~new_P1_R1138_U78;
  assign new_P1_R1138_U175 = ~new_P1_U3065 | ~new_P1_U3978;
  assign new_P1_R1138_U176 = ~new_P1_R1138_U62;
  assign new_P1_R1138_U177 = new_P1_U3067 | new_P1_U3467;
  assign new_P1_R1138_U178 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1138_U179 = new_P1_U3461 | new_P1_U3064;
  assign new_P1_R1138_U180 = new_P1_U3458 | new_P1_U3068;
  assign new_P1_R1138_U181 = ~new_P1_R1138_U32;
  assign new_P1_R1138_U182 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1138_U183 = ~new_P1_R1138_U43;
  assign new_P1_R1138_U184 = ~new_P1_R1138_U44;
  assign new_P1_R1138_U185 = ~new_P1_R1138_U43 | ~new_P1_R1138_U44;
  assign new_P1_R1138_U186 = ~new_P1_R1138_U116 | ~new_P1_R1138_U179;
  assign new_P1_R1138_U187 = ~new_P1_R1138_U5 | ~new_P1_R1138_U185;
  assign new_P1_R1138_U188 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1138_U189 = ~new_P1_R1138_U117 | ~new_P1_R1138_U187;
  assign new_P1_R1138_U190 = ~new_P1_R1138_U36 | ~new_P1_R1138_U35;
  assign new_P1_R1138_U191 = ~new_P1_U3067 | ~new_P1_R1138_U190;
  assign new_P1_R1138_U192 = ~new_P1_R1138_U4 | ~new_P1_R1138_U189;
  assign new_P1_R1138_U193 = ~new_P1_U3467 | ~new_P1_R1138_U169;
  assign new_P1_R1138_U194 = ~new_P1_R1138_U42;
  assign new_P1_R1138_U195 = new_P1_U3070 | new_P1_U3473;
  assign new_P1_R1138_U196 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1138_U197 = ~new_P1_R1138_U23;
  assign new_P1_R1138_U198 = ~new_P1_R1138_U24 | ~new_P1_R1138_U23;
  assign new_P1_R1138_U199 = ~new_P1_U3070 | ~new_P1_R1138_U198;
  assign new_P1_R1138_U200 = ~new_P1_U3473 | ~new_P1_R1138_U197;
  assign new_P1_R1138_U201 = ~new_P1_R1138_U6 | ~new_P1_R1138_U42;
  assign new_P1_R1138_U202 = ~new_P1_R1138_U143;
  assign new_P1_R1138_U203 = new_P1_U3476 | new_P1_U3084;
  assign new_P1_R1138_U204 = ~new_P1_R1138_U203 | ~new_P1_R1138_U143;
  assign new_P1_R1138_U205 = ~new_P1_R1138_U41;
  assign new_P1_R1138_U206 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1138_U207 = new_P1_U3470 | new_P1_U3071;
  assign new_P1_R1138_U208 = ~new_P1_R1138_U207 | ~new_P1_R1138_U42;
  assign new_P1_R1138_U209 = ~new_P1_R1138_U120 | ~new_P1_R1138_U208;
  assign new_P1_R1138_U210 = ~new_P1_R1138_U194 | ~new_P1_R1138_U23;
  assign new_P1_R1138_U211 = ~new_P1_U3473 | ~new_P1_U3070;
  assign new_P1_R1138_U212 = ~new_P1_R1138_U121 | ~new_P1_R1138_U210;
  assign new_P1_R1138_U213 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1138_U214 = ~new_P1_R1138_U184 | ~new_P1_R1138_U180;
  assign new_P1_R1138_U215 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1138_U216 = ~new_P1_R1138_U46;
  assign new_P1_R1138_U217 = ~new_P1_R1138_U183 | ~new_P1_R1138_U5;
  assign new_P1_R1138_U218 = ~new_P1_R1138_U46 | ~new_P1_R1138_U179;
  assign new_P1_R1138_U219 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1138_U220 = ~new_P1_R1138_U45;
  assign new_P1_R1138_U221 = new_P1_U3464 | new_P1_U3060;
  assign new_P1_R1138_U222 = ~new_P1_R1138_U221 | ~new_P1_R1138_U45;
  assign new_P1_R1138_U223 = ~new_P1_R1138_U123 | ~new_P1_R1138_U222;
  assign new_P1_R1138_U224 = ~new_P1_R1138_U220 | ~new_P1_R1138_U35;
  assign new_P1_R1138_U225 = ~new_P1_U3467 | ~new_P1_U3067;
  assign new_P1_R1138_U226 = ~new_P1_R1138_U124 | ~new_P1_R1138_U224;
  assign new_P1_R1138_U227 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1138_U228 = ~new_P1_R1138_U183 | ~new_P1_R1138_U180;
  assign new_P1_R1138_U229 = ~new_P1_R1138_U144;
  assign new_P1_R1138_U230 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1138_U231 = ~new_P1_R1138_U43 | ~new_P1_R1138_U44 | ~new_P1_R1138_U400 | ~new_P1_R1138_U399;
  assign new_P1_R1138_U232 = ~new_P1_R1138_U44 | ~new_P1_R1138_U43;
  assign new_P1_R1138_U233 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1138_U234 = ~new_P1_R1138_U125 | ~new_P1_R1138_U232;
  assign new_P1_R1138_U235 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1138_U236 = new_P1_U3062 | new_P1_U3482;
  assign new_P1_R1138_U237 = ~new_P1_R1138_U176 | ~new_P1_R1138_U7;
  assign new_P1_R1138_U238 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1138_U239 = ~new_P1_R1138_U127 | ~new_P1_R1138_U237;
  assign new_P1_R1138_U240 = new_P1_U3482 | new_P1_U3062;
  assign new_P1_R1138_U241 = ~new_P1_R1138_U126 | ~new_P1_R1138_U143;
  assign new_P1_R1138_U242 = ~new_P1_R1138_U240 | ~new_P1_R1138_U239;
  assign new_P1_R1138_U243 = ~new_P1_R1138_U166;
  assign new_P1_R1138_U244 = new_P1_U3080 | new_P1_U3491;
  assign new_P1_R1138_U245 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1138_U246 = ~new_P1_R1138_U173 | ~new_P1_R1138_U8;
  assign new_P1_R1138_U247 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1138_U248 = ~new_P1_R1138_U129 | ~new_P1_R1138_U246;
  assign new_P1_R1138_U249 = new_P1_U3485 | new_P1_U3063;
  assign new_P1_R1138_U250 = new_P1_U3491 | new_P1_U3080;
  assign new_P1_R1138_U251 = ~new_P1_R1138_U128 | ~new_P1_R1138_U166;
  assign new_P1_R1138_U252 = ~new_P1_R1138_U250 | ~new_P1_R1138_U248;
  assign new_P1_R1138_U253 = ~new_P1_R1138_U165;
  assign new_P1_R1138_U254 = new_P1_U3494 | new_P1_U3079;
  assign new_P1_R1138_U255 = ~new_P1_R1138_U254 | ~new_P1_R1138_U165;
  assign new_P1_R1138_U256 = ~new_P1_U3079 | ~new_P1_U3494;
  assign new_P1_R1138_U257 = ~new_P1_R1138_U163;
  assign new_P1_R1138_U258 = new_P1_U3497 | new_P1_U3074;
  assign new_P1_R1138_U259 = ~new_P1_R1138_U258 | ~new_P1_R1138_U163;
  assign new_P1_R1138_U260 = ~new_P1_U3074 | ~new_P1_U3497;
  assign new_P1_R1138_U261 = ~new_P1_R1138_U93;
  assign new_P1_R1138_U262 = new_P1_U3069 | new_P1_U3503;
  assign new_P1_R1138_U263 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1138_U264 = ~new_P1_R1138_U60;
  assign new_P1_R1138_U265 = ~new_P1_R1138_U61 | ~new_P1_R1138_U60;
  assign new_P1_R1138_U266 = ~new_P1_U3069 | ~new_P1_R1138_U265;
  assign new_P1_R1138_U267 = ~new_P1_U3503 | ~new_P1_R1138_U264;
  assign new_P1_R1138_U268 = ~new_P1_R1138_U9 | ~new_P1_R1138_U93;
  assign new_P1_R1138_U269 = ~new_P1_R1138_U161;
  assign new_P1_R1138_U270 = new_P1_U3076 | new_P1_U3982;
  assign new_P1_R1138_U271 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1138_U272 = new_P1_U3075 | new_P1_U3981;
  assign new_P1_R1138_U273 = ~new_P1_R1138_U81;
  assign new_P1_R1138_U274 = ~new_P1_U3982 | ~new_P1_R1138_U273;
  assign new_P1_R1138_U275 = ~new_P1_R1138_U274 | ~new_P1_R1138_U91;
  assign new_P1_R1138_U276 = ~new_P1_R1138_U81 | ~new_P1_R1138_U82;
  assign new_P1_R1138_U277 = ~new_P1_R1138_U276 | ~new_P1_R1138_U275;
  assign new_P1_R1138_U278 = ~new_P1_R1138_U174 | ~new_P1_R1138_U10;
  assign new_P1_R1138_U279 = ~new_P1_U3075 | ~new_P1_U3981;
  assign new_P1_R1138_U280 = ~new_P1_R1138_U277 | ~new_P1_R1138_U278;
  assign new_P1_R1138_U281 = new_P1_U3506 | new_P1_U3082;
  assign new_P1_R1138_U282 = new_P1_U3981 | new_P1_U3075;
  assign new_P1_R1138_U283 = ~new_P1_R1138_U131 | ~new_P1_R1138_U272 | ~new_P1_R1138_U161;
  assign new_P1_R1138_U284 = ~new_P1_R1138_U282 | ~new_P1_R1138_U280;
  assign new_P1_R1138_U285 = ~new_P1_R1138_U158;
  assign new_P1_R1138_U286 = new_P1_U3980 | new_P1_U3061;
  assign new_P1_R1138_U287 = ~new_P1_R1138_U286 | ~new_P1_R1138_U158;
  assign new_P1_R1138_U288 = ~new_P1_U3061 | ~new_P1_U3980;
  assign new_P1_R1138_U289 = ~new_P1_R1138_U156;
  assign new_P1_R1138_U290 = new_P1_U3979 | new_P1_U3066;
  assign new_P1_R1138_U291 = ~new_P1_R1138_U290 | ~new_P1_R1138_U156;
  assign new_P1_R1138_U292 = ~new_P1_U3066 | ~new_P1_U3979;
  assign new_P1_R1138_U293 = ~new_P1_R1138_U154;
  assign new_P1_R1138_U294 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1138_U295 = ~new_P1_R1138_U175 | ~new_P1_R1138_U172;
  assign new_P1_R1138_U296 = ~new_P1_R1138_U87;
  assign new_P1_R1138_U297 = new_P1_U3978 | new_P1_U3065;
  assign new_P1_R1138_U298 = ~new_P1_R1138_U167 | ~new_P1_R1138_U154 | ~new_P1_R1138_U297;
  assign new_P1_R1138_U299 = ~new_P1_R1138_U152;
  assign new_P1_R1138_U300 = new_P1_U3975 | new_P1_U3053;
  assign new_P1_R1138_U301 = ~new_P1_U3053 | ~new_P1_U3975;
  assign new_P1_R1138_U302 = ~new_P1_R1138_U150;
  assign new_P1_R1138_U303 = ~new_P1_U3974 | ~new_P1_R1138_U150;
  assign new_P1_R1138_U304 = ~new_P1_R1138_U148;
  assign new_P1_R1138_U305 = ~new_P1_R1138_U297 | ~new_P1_R1138_U154;
  assign new_P1_R1138_U306 = ~new_P1_R1138_U90;
  assign new_P1_R1138_U307 = new_P1_U3977 | new_P1_U3058;
  assign new_P1_R1138_U308 = ~new_P1_R1138_U307 | ~new_P1_R1138_U90;
  assign new_P1_R1138_U309 = ~new_P1_R1138_U153 | ~new_P1_R1138_U308 | ~new_P1_R1138_U172;
  assign new_P1_R1138_U310 = ~new_P1_R1138_U306 | ~new_P1_R1138_U172;
  assign new_P1_R1138_U311 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1138_U312 = ~new_P1_R1138_U167 | ~new_P1_R1138_U310 | ~new_P1_R1138_U311;
  assign new_P1_R1138_U313 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1138_U314 = ~new_P1_R1138_U281 | ~new_P1_R1138_U161;
  assign new_P1_R1138_U315 = ~new_P1_R1138_U92;
  assign new_P1_R1138_U316 = ~new_P1_R1138_U10 | ~new_P1_R1138_U92;
  assign new_P1_R1138_U317 = ~new_P1_R1138_U135 | ~new_P1_R1138_U316;
  assign new_P1_R1138_U318 = ~new_P1_R1138_U316 | ~new_P1_R1138_U277;
  assign new_P1_R1138_U319 = ~new_P1_R1138_U452 | ~new_P1_R1138_U318;
  assign new_P1_R1138_U320 = new_P1_U3508 | new_P1_U3081;
  assign new_P1_R1138_U321 = ~new_P1_R1138_U320 | ~new_P1_R1138_U92;
  assign new_P1_R1138_U322 = ~new_P1_R1138_U136 | ~new_P1_R1138_U321;
  assign new_P1_R1138_U323 = ~new_P1_R1138_U315 | ~new_P1_R1138_U81;
  assign new_P1_R1138_U324 = ~new_P1_U3076 | ~new_P1_U3982;
  assign new_P1_R1138_U325 = ~new_P1_R1138_U10 | ~new_P1_R1138_U324 | ~new_P1_R1138_U323;
  assign new_P1_R1138_U326 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1138_U327 = ~new_P1_R1138_U160;
  assign new_P1_R1138_U328 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1138_U329 = new_P1_U3500 | new_P1_U3073;
  assign new_P1_R1138_U330 = ~new_P1_R1138_U329 | ~new_P1_R1138_U93;
  assign new_P1_R1138_U331 = ~new_P1_R1138_U137 | ~new_P1_R1138_U330;
  assign new_P1_R1138_U332 = ~new_P1_R1138_U261 | ~new_P1_R1138_U60;
  assign new_P1_R1138_U333 = ~new_P1_U3503 | ~new_P1_U3069;
  assign new_P1_R1138_U334 = ~new_P1_R1138_U138 | ~new_P1_R1138_U332;
  assign new_P1_R1138_U335 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1138_U336 = ~new_P1_R1138_U249 | ~new_P1_R1138_U166;
  assign new_P1_R1138_U337 = ~new_P1_R1138_U94;
  assign new_P1_R1138_U338 = new_P1_U3488 | new_P1_U3072;
  assign new_P1_R1138_U339 = ~new_P1_R1138_U338 | ~new_P1_R1138_U94;
  assign new_P1_R1138_U340 = ~new_P1_R1138_U139 | ~new_P1_R1138_U339;
  assign new_P1_R1138_U341 = ~new_P1_R1138_U337 | ~new_P1_R1138_U171;
  assign new_P1_R1138_U342 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1138_U343 = ~new_P1_R1138_U140 | ~new_P1_R1138_U341;
  assign new_P1_R1138_U344 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1138_U345 = new_P1_U3479 | new_P1_U3083;
  assign new_P1_R1138_U346 = ~new_P1_R1138_U345 | ~new_P1_R1138_U41;
  assign new_P1_R1138_U347 = ~new_P1_R1138_U141 | ~new_P1_R1138_U346;
  assign new_P1_R1138_U348 = ~new_P1_R1138_U205 | ~new_P1_R1138_U170;
  assign new_P1_R1138_U349 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1138_U350 = ~new_P1_R1138_U142 | ~new_P1_R1138_U348;
  assign new_P1_R1138_U351 = ~new_P1_R1138_U206 | ~new_P1_R1138_U170;
  assign new_P1_R1138_U352 = ~new_P1_R1138_U203 | ~new_P1_R1138_U62;
  assign new_P1_R1138_U353 = ~new_P1_R1138_U213 | ~new_P1_R1138_U23;
  assign new_P1_R1138_U354 = ~new_P1_R1138_U227 | ~new_P1_R1138_U35;
  assign new_P1_R1138_U355 = ~new_P1_R1138_U230 | ~new_P1_R1138_U179;
  assign new_P1_R1138_U356 = ~new_P1_R1138_U313 | ~new_P1_R1138_U172;
  assign new_P1_R1138_U357 = ~new_P1_R1138_U297 | ~new_P1_R1138_U175;
  assign new_P1_R1138_U358 = ~new_P1_R1138_U328 | ~new_P1_R1138_U81;
  assign new_P1_R1138_U359 = ~new_P1_R1138_U281 | ~new_P1_R1138_U78;
  assign new_P1_R1138_U360 = ~new_P1_R1138_U335 | ~new_P1_R1138_U60;
  assign new_P1_R1138_U361 = ~new_P1_R1138_U344 | ~new_P1_R1138_U171;
  assign new_P1_R1138_U362 = ~new_P1_R1138_U249 | ~new_P1_R1138_U69;
  assign new_P1_R1138_U363 = ~new_P1_U3974 | ~new_P1_U3054;
  assign new_P1_R1138_U364 = ~new_P1_R1138_U295 | ~new_P1_R1138_U167;
  assign new_P1_R1138_U365 = ~new_P1_U3057 | ~new_P1_R1138_U294;
  assign new_P1_R1138_U366 = ~new_P1_U3976 | ~new_P1_R1138_U294;
  assign new_P1_R1138_U367 = ~new_P1_R1138_U300 | ~new_P1_R1138_U295 | ~new_P1_R1138_U167;
  assign new_P1_R1138_U368 = ~new_P1_R1138_U133 | ~new_P1_R1138_U154 | ~new_P1_R1138_U167;
  assign new_P1_R1138_U369 = ~new_P1_R1138_U296 | ~new_P1_R1138_U300;
  assign new_P1_R1138_U370 = ~new_P1_U3083 | ~new_P1_R1138_U40;
  assign new_P1_R1138_U371 = ~new_P1_U3479 | ~new_P1_R1138_U39;
  assign new_P1_R1138_U372 = ~new_P1_R1138_U371 | ~new_P1_R1138_U370;
  assign new_P1_R1138_U373 = ~new_P1_R1138_U351 | ~new_P1_R1138_U41;
  assign new_P1_R1138_U374 = ~new_P1_R1138_U372 | ~new_P1_R1138_U205;
  assign new_P1_R1138_U375 = ~new_P1_U3084 | ~new_P1_R1138_U37;
  assign new_P1_R1138_U376 = ~new_P1_U3476 | ~new_P1_R1138_U38;
  assign new_P1_R1138_U377 = ~new_P1_R1138_U376 | ~new_P1_R1138_U375;
  assign new_P1_R1138_U378 = ~new_P1_R1138_U352 | ~new_P1_R1138_U143;
  assign new_P1_R1138_U379 = ~new_P1_R1138_U202 | ~new_P1_R1138_U377;
  assign new_P1_R1138_U380 = ~new_P1_U3070 | ~new_P1_R1138_U24;
  assign new_P1_R1138_U381 = ~new_P1_U3473 | ~new_P1_R1138_U22;
  assign new_P1_R1138_U382 = ~new_P1_U3071 | ~new_P1_R1138_U20;
  assign new_P1_R1138_U383 = ~new_P1_U3470 | ~new_P1_R1138_U21;
  assign new_P1_R1138_U384 = ~new_P1_R1138_U383 | ~new_P1_R1138_U382;
  assign new_P1_R1138_U385 = ~new_P1_R1138_U353 | ~new_P1_R1138_U42;
  assign new_P1_R1138_U386 = ~new_P1_R1138_U384 | ~new_P1_R1138_U194;
  assign new_P1_R1138_U387 = ~new_P1_U3067 | ~new_P1_R1138_U36;
  assign new_P1_R1138_U388 = ~new_P1_U3467 | ~new_P1_R1138_U27;
  assign new_P1_R1138_U389 = ~new_P1_U3060 | ~new_P1_R1138_U25;
  assign new_P1_R1138_U390 = ~new_P1_U3464 | ~new_P1_R1138_U26;
  assign new_P1_R1138_U391 = ~new_P1_R1138_U390 | ~new_P1_R1138_U389;
  assign new_P1_R1138_U392 = ~new_P1_R1138_U354 | ~new_P1_R1138_U45;
  assign new_P1_R1138_U393 = ~new_P1_R1138_U391 | ~new_P1_R1138_U220;
  assign new_P1_R1138_U394 = ~new_P1_U3064 | ~new_P1_R1138_U33;
  assign new_P1_R1138_U395 = ~new_P1_U3461 | ~new_P1_R1138_U34;
  assign new_P1_R1138_U396 = ~new_P1_R1138_U395 | ~new_P1_R1138_U394;
  assign new_P1_R1138_U397 = ~new_P1_R1138_U355 | ~new_P1_R1138_U144;
  assign new_P1_R1138_U398 = ~new_P1_R1138_U229 | ~new_P1_R1138_U396;
  assign new_P1_R1138_U399 = ~new_P1_U3068 | ~new_P1_R1138_U28;
  assign new_P1_R1138_U400 = ~new_P1_U3458 | ~new_P1_R1138_U29;
  assign new_P1_R1138_U401 = ~new_P1_U3055 | ~new_P1_R1138_U146;
  assign new_P1_R1138_U402 = ~new_P1_U3985 | ~new_P1_R1138_U145;
  assign new_P1_R1138_U403 = ~new_P1_U3055 | ~new_P1_R1138_U146;
  assign new_P1_R1138_U404 = ~new_P1_U3985 | ~new_P1_R1138_U145;
  assign new_P1_R1138_U405 = ~new_P1_R1138_U404 | ~new_P1_R1138_U403;
  assign new_P1_R1138_U406 = ~new_P1_R1138_U147 | ~new_P1_R1138_U148;
  assign new_P1_R1138_U407 = ~new_P1_R1138_U304 | ~new_P1_R1138_U405;
  assign new_P1_R1138_U408 = ~new_P1_U3054 | ~new_P1_R1138_U89;
  assign new_P1_R1138_U409 = ~new_P1_U3974 | ~new_P1_R1138_U88;
  assign new_P1_R1138_U410 = ~new_P1_U3054 | ~new_P1_R1138_U89;
  assign new_P1_R1138_U411 = ~new_P1_U3974 | ~new_P1_R1138_U88;
  assign new_P1_R1138_U412 = ~new_P1_R1138_U411 | ~new_P1_R1138_U410;
  assign new_P1_R1138_U413 = ~new_P1_R1138_U149 | ~new_P1_R1138_U150;
  assign new_P1_R1138_U414 = ~new_P1_R1138_U302 | ~new_P1_R1138_U412;
  assign new_P1_R1138_U415 = ~new_P1_U3053 | ~new_P1_R1138_U47;
  assign new_P1_R1138_U416 = ~new_P1_U3975 | ~new_P1_R1138_U48;
  assign new_P1_R1138_U417 = ~new_P1_U3053 | ~new_P1_R1138_U47;
  assign new_P1_R1138_U418 = ~new_P1_U3975 | ~new_P1_R1138_U48;
  assign new_P1_R1138_U419 = ~new_P1_R1138_U418 | ~new_P1_R1138_U417;
  assign new_P1_R1138_U420 = ~new_P1_R1138_U151 | ~new_P1_R1138_U152;
  assign new_P1_R1138_U421 = ~new_P1_R1138_U299 | ~new_P1_R1138_U419;
  assign new_P1_R1138_U422 = ~new_P1_U3057 | ~new_P1_R1138_U50;
  assign new_P1_R1138_U423 = ~new_P1_U3976 | ~new_P1_R1138_U49;
  assign new_P1_R1138_U424 = ~new_P1_U3058 | ~new_P1_R1138_U51;
  assign new_P1_R1138_U425 = ~new_P1_U3977 | ~new_P1_R1138_U52;
  assign new_P1_R1138_U426 = ~new_P1_R1138_U425 | ~new_P1_R1138_U424;
  assign new_P1_R1138_U427 = ~new_P1_R1138_U356 | ~new_P1_R1138_U90;
  assign new_P1_R1138_U428 = ~new_P1_R1138_U426 | ~new_P1_R1138_U306;
  assign new_P1_R1138_U429 = ~new_P1_U3065 | ~new_P1_R1138_U53;
  assign new_P1_R1138_U430 = ~new_P1_U3978 | ~new_P1_R1138_U54;
  assign new_P1_R1138_U431 = ~new_P1_R1138_U430 | ~new_P1_R1138_U429;
  assign new_P1_R1138_U432 = ~new_P1_R1138_U357 | ~new_P1_R1138_U154;
  assign new_P1_R1138_U433 = ~new_P1_R1138_U293 | ~new_P1_R1138_U431;
  assign new_P1_R1138_U434 = ~new_P1_U3066 | ~new_P1_R1138_U85;
  assign new_P1_R1138_U435 = ~new_P1_U3979 | ~new_P1_R1138_U86;
  assign new_P1_R1138_U436 = ~new_P1_U3066 | ~new_P1_R1138_U85;
  assign new_P1_R1138_U437 = ~new_P1_U3979 | ~new_P1_R1138_U86;
  assign new_P1_R1138_U438 = ~new_P1_R1138_U437 | ~new_P1_R1138_U436;
  assign new_P1_R1138_U439 = ~new_P1_R1138_U155 | ~new_P1_R1138_U156;
  assign new_P1_R1138_U440 = ~new_P1_R1138_U289 | ~new_P1_R1138_U438;
  assign new_P1_R1138_U441 = ~new_P1_U3061 | ~new_P1_R1138_U83;
  assign new_P1_R1138_U442 = ~new_P1_U3980 | ~new_P1_R1138_U84;
  assign new_P1_R1138_U443 = ~new_P1_U3061 | ~new_P1_R1138_U83;
  assign new_P1_R1138_U444 = ~new_P1_U3980 | ~new_P1_R1138_U84;
  assign new_P1_R1138_U445 = ~new_P1_R1138_U444 | ~new_P1_R1138_U443;
  assign new_P1_R1138_U446 = ~new_P1_R1138_U157 | ~new_P1_R1138_U158;
  assign new_P1_R1138_U447 = ~new_P1_R1138_U285 | ~new_P1_R1138_U445;
  assign new_P1_R1138_U448 = ~new_P1_U3075 | ~new_P1_R1138_U55;
  assign new_P1_R1138_U449 = ~new_P1_U3981 | ~new_P1_R1138_U56;
  assign new_P1_R1138_U450 = ~new_P1_U3075 | ~new_P1_R1138_U55;
  assign new_P1_R1138_U451 = ~new_P1_U3981 | ~new_P1_R1138_U56;
  assign new_P1_R1138_U452 = ~new_P1_R1138_U451 | ~new_P1_R1138_U450;
  assign new_P1_R1138_U453 = ~new_P1_U3076 | ~new_P1_R1138_U82;
  assign new_P1_R1138_U454 = ~new_P1_U3982 | ~new_P1_R1138_U91;
  assign new_P1_R1138_U455 = ~new_P1_R1138_U181 | ~new_P1_R1138_U160;
  assign new_P1_R1138_U456 = ~new_P1_R1138_U327 | ~new_P1_R1138_U32;
  assign new_P1_R1138_U457 = ~new_P1_U3081 | ~new_P1_R1138_U79;
  assign new_P1_R1138_U458 = ~new_P1_U3508 | ~new_P1_R1138_U80;
  assign new_P1_R1138_U459 = ~new_P1_R1138_U458 | ~new_P1_R1138_U457;
  assign new_P1_R1138_U460 = ~new_P1_R1138_U358 | ~new_P1_R1138_U92;
  assign new_P1_R1138_U461 = ~new_P1_R1138_U459 | ~new_P1_R1138_U315;
  assign new_P1_R1138_U462 = ~new_P1_U3082 | ~new_P1_R1138_U76;
  assign new_P1_R1138_U463 = ~new_P1_U3506 | ~new_P1_R1138_U77;
  assign new_P1_R1138_U464 = ~new_P1_R1138_U463 | ~new_P1_R1138_U462;
  assign new_P1_R1138_U465 = ~new_P1_R1138_U359 | ~new_P1_R1138_U161;
  assign new_P1_R1138_U466 = ~new_P1_R1138_U269 | ~new_P1_R1138_U464;
  assign new_P1_R1138_U467 = ~new_P1_U3069 | ~new_P1_R1138_U61;
  assign new_P1_R1138_U468 = ~new_P1_U3503 | ~new_P1_R1138_U59;
  assign new_P1_R1138_U469 = ~new_P1_U3073 | ~new_P1_R1138_U57;
  assign new_P1_R1138_U470 = ~new_P1_U3500 | ~new_P1_R1138_U58;
  assign new_P1_R1138_U471 = ~new_P1_R1138_U470 | ~new_P1_R1138_U469;
  assign new_P1_R1138_U472 = ~new_P1_R1138_U360 | ~new_P1_R1138_U93;
  assign new_P1_R1138_U473 = ~new_P1_R1138_U471 | ~new_P1_R1138_U261;
  assign new_P1_R1138_U474 = ~new_P1_U3074 | ~new_P1_R1138_U74;
  assign new_P1_R1138_U475 = ~new_P1_U3497 | ~new_P1_R1138_U75;
  assign new_P1_R1138_U476 = ~new_P1_U3074 | ~new_P1_R1138_U74;
  assign new_P1_R1138_U477 = ~new_P1_U3497 | ~new_P1_R1138_U75;
  assign new_P1_R1138_U478 = ~new_P1_R1138_U477 | ~new_P1_R1138_U476;
  assign new_P1_R1138_U479 = ~new_P1_R1138_U162 | ~new_P1_R1138_U163;
  assign new_P1_R1138_U480 = ~new_P1_R1138_U257 | ~new_P1_R1138_U478;
  assign new_P1_R1138_U481 = ~new_P1_U3079 | ~new_P1_R1138_U72;
  assign new_P1_R1138_U482 = ~new_P1_U3494 | ~new_P1_R1138_U73;
  assign new_P1_R1138_U483 = ~new_P1_U3079 | ~new_P1_R1138_U72;
  assign new_P1_R1138_U484 = ~new_P1_U3494 | ~new_P1_R1138_U73;
  assign new_P1_R1138_U485 = ~new_P1_R1138_U484 | ~new_P1_R1138_U483;
  assign new_P1_R1138_U486 = ~new_P1_R1138_U164 | ~new_P1_R1138_U165;
  assign new_P1_R1138_U487 = ~new_P1_R1138_U253 | ~new_P1_R1138_U485;
  assign new_P1_R1138_U488 = ~new_P1_U3080 | ~new_P1_R1138_U70;
  assign new_P1_R1138_U489 = ~new_P1_U3491 | ~new_P1_R1138_U71;
  assign new_P1_R1138_U490 = ~new_P1_U3072 | ~new_P1_R1138_U65;
  assign new_P1_R1138_U491 = ~new_P1_U3488 | ~new_P1_R1138_U66;
  assign new_P1_R1138_U492 = ~new_P1_R1138_U491 | ~new_P1_R1138_U490;
  assign new_P1_R1138_U493 = ~new_P1_R1138_U361 | ~new_P1_R1138_U94;
  assign new_P1_R1138_U494 = ~new_P1_R1138_U492 | ~new_P1_R1138_U337;
  assign new_P1_R1138_U495 = ~new_P1_U3063 | ~new_P1_R1138_U67;
  assign new_P1_R1138_U496 = ~new_P1_U3485 | ~new_P1_R1138_U68;
  assign new_P1_R1138_U497 = ~new_P1_R1138_U496 | ~new_P1_R1138_U495;
  assign new_P1_R1138_U498 = ~new_P1_R1138_U362 | ~new_P1_R1138_U166;
  assign new_P1_R1138_U499 = ~new_P1_R1138_U243 | ~new_P1_R1138_U497;
  assign new_P1_R1138_U500 = ~new_P1_U3062 | ~new_P1_R1138_U63;
  assign new_P1_R1138_U501 = ~new_P1_U3482 | ~new_P1_R1138_U64;
  assign new_P1_R1138_U502 = ~new_P1_U3077 | ~new_P1_R1138_U30;
  assign new_P1_R1138_U503 = ~new_P1_U3450 | ~new_P1_R1138_U31;
  assign new_P1_R1222_U4 = new_P1_R1222_U178 & new_P1_R1222_U177;
  assign new_P1_R1222_U5 = new_P1_R1222_U179 & new_P1_R1222_U180;
  assign new_P1_R1222_U6 = new_P1_R1222_U196 & new_P1_R1222_U195;
  assign new_P1_R1222_U7 = new_P1_R1222_U236 & new_P1_R1222_U235;
  assign new_P1_R1222_U8 = new_P1_R1222_U245 & new_P1_R1222_U244;
  assign new_P1_R1222_U9 = new_P1_R1222_U263 & new_P1_R1222_U262;
  assign new_P1_R1222_U10 = new_P1_R1222_U271 & new_P1_R1222_U270;
  assign new_P1_R1222_U11 = new_P1_R1222_U350 & new_P1_R1222_U347;
  assign new_P1_R1222_U12 = new_P1_R1222_U343 & new_P1_R1222_U340;
  assign new_P1_R1222_U13 = new_P1_R1222_U334 & new_P1_R1222_U331;
  assign new_P1_R1222_U14 = new_P1_R1222_U325 & new_P1_R1222_U322;
  assign new_P1_R1222_U15 = new_P1_R1222_U319 & new_P1_R1222_U317;
  assign new_P1_R1222_U16 = new_P1_R1222_U312 & new_P1_R1222_U309;
  assign new_P1_R1222_U17 = new_P1_R1222_U234 & new_P1_R1222_U231;
  assign new_P1_R1222_U18 = new_P1_R1222_U226 & new_P1_R1222_U223;
  assign new_P1_R1222_U19 = new_P1_R1222_U212 & new_P1_R1222_U209;
  assign new_P1_R1222_U20 = ~new_P1_U3470;
  assign new_P1_R1222_U21 = ~new_P1_U3071;
  assign new_P1_R1222_U22 = ~new_P1_U3070;
  assign new_P1_R1222_U23 = ~new_P1_U3071 | ~new_P1_U3470;
  assign new_P1_R1222_U24 = ~new_P1_U3473;
  assign new_P1_R1222_U25 = ~new_P1_U3464;
  assign new_P1_R1222_U26 = ~new_P1_U3060;
  assign new_P1_R1222_U27 = ~new_P1_U3067;
  assign new_P1_R1222_U28 = ~new_P1_U3458;
  assign new_P1_R1222_U29 = ~new_P1_U3068;
  assign new_P1_R1222_U30 = ~new_P1_U3450;
  assign new_P1_R1222_U31 = ~new_P1_U3077;
  assign new_P1_R1222_U32 = ~new_P1_U3077 | ~new_P1_U3450;
  assign new_P1_R1222_U33 = ~new_P1_U3461;
  assign new_P1_R1222_U34 = ~new_P1_U3064;
  assign new_P1_R1222_U35 = ~new_P1_U3060 | ~new_P1_U3464;
  assign new_P1_R1222_U36 = ~new_P1_U3467;
  assign new_P1_R1222_U37 = ~new_P1_U3476;
  assign new_P1_R1222_U38 = ~new_P1_U3084;
  assign new_P1_R1222_U39 = ~new_P1_U3083;
  assign new_P1_R1222_U40 = ~new_P1_U3479;
  assign new_P1_R1222_U41 = ~new_P1_R1222_U62 | ~new_P1_R1222_U204;
  assign new_P1_R1222_U42 = ~new_P1_R1222_U118 | ~new_P1_R1222_U192;
  assign new_P1_R1222_U43 = ~new_P1_R1222_U181 | ~new_P1_R1222_U182;
  assign new_P1_R1222_U44 = ~new_P1_U3455 | ~new_P1_U3078;
  assign new_P1_R1222_U45 = ~new_P1_R1222_U122 | ~new_P1_R1222_U218;
  assign new_P1_R1222_U46 = ~new_P1_R1222_U215 | ~new_P1_R1222_U214;
  assign new_P1_R1222_U47 = ~new_P1_U3975;
  assign new_P1_R1222_U48 = ~new_P1_U3053;
  assign new_P1_R1222_U49 = ~new_P1_U3057;
  assign new_P1_R1222_U50 = ~new_P1_U3976;
  assign new_P1_R1222_U51 = ~new_P1_U3977;
  assign new_P1_R1222_U52 = ~new_P1_U3058;
  assign new_P1_R1222_U53 = ~new_P1_U3978;
  assign new_P1_R1222_U54 = ~new_P1_U3065;
  assign new_P1_R1222_U55 = ~new_P1_U3981;
  assign new_P1_R1222_U56 = ~new_P1_U3075;
  assign new_P1_R1222_U57 = ~new_P1_U3500;
  assign new_P1_R1222_U58 = ~new_P1_U3073;
  assign new_P1_R1222_U59 = ~new_P1_U3069;
  assign new_P1_R1222_U60 = ~new_P1_U3073 | ~new_P1_U3500;
  assign new_P1_R1222_U61 = ~new_P1_U3503;
  assign new_P1_R1222_U62 = ~new_P1_U3084 | ~new_P1_U3476;
  assign new_P1_R1222_U63 = ~new_P1_U3482;
  assign new_P1_R1222_U64 = ~new_P1_U3062;
  assign new_P1_R1222_U65 = ~new_P1_U3488;
  assign new_P1_R1222_U66 = ~new_P1_U3072;
  assign new_P1_R1222_U67 = ~new_P1_U3485;
  assign new_P1_R1222_U68 = ~new_P1_U3063;
  assign new_P1_R1222_U69 = ~new_P1_U3063 | ~new_P1_U3485;
  assign new_P1_R1222_U70 = ~new_P1_U3491;
  assign new_P1_R1222_U71 = ~new_P1_U3080;
  assign new_P1_R1222_U72 = ~new_P1_U3494;
  assign new_P1_R1222_U73 = ~new_P1_U3079;
  assign new_P1_R1222_U74 = ~new_P1_U3497;
  assign new_P1_R1222_U75 = ~new_P1_U3074;
  assign new_P1_R1222_U76 = ~new_P1_U3506;
  assign new_P1_R1222_U77 = ~new_P1_U3082;
  assign new_P1_R1222_U78 = ~new_P1_U3082 | ~new_P1_U3506;
  assign new_P1_R1222_U79 = ~new_P1_U3508;
  assign new_P1_R1222_U80 = ~new_P1_U3081;
  assign new_P1_R1222_U81 = ~new_P1_U3081 | ~new_P1_U3508;
  assign new_P1_R1222_U82 = ~new_P1_U3982;
  assign new_P1_R1222_U83 = ~new_P1_U3980;
  assign new_P1_R1222_U84 = ~new_P1_U3061;
  assign new_P1_R1222_U85 = ~new_P1_U3979;
  assign new_P1_R1222_U86 = ~new_P1_U3066;
  assign new_P1_R1222_U87 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1222_U88 = ~new_P1_U3054;
  assign new_P1_R1222_U89 = ~new_P1_U3974;
  assign new_P1_R1222_U90 = ~new_P1_R1222_U305 | ~new_P1_R1222_U175;
  assign new_P1_R1222_U91 = ~new_P1_U3076;
  assign new_P1_R1222_U92 = ~new_P1_R1222_U78 | ~new_P1_R1222_U314;
  assign new_P1_R1222_U93 = ~new_P1_R1222_U260 | ~new_P1_R1222_U259;
  assign new_P1_R1222_U94 = ~new_P1_R1222_U69 | ~new_P1_R1222_U336;
  assign new_P1_R1222_U95 = ~new_P1_R1222_U456 | ~new_P1_R1222_U455;
  assign new_P1_R1222_U96 = ~new_P1_R1222_U503 | ~new_P1_R1222_U502;
  assign new_P1_R1222_U97 = ~new_P1_R1222_U374 | ~new_P1_R1222_U373;
  assign new_P1_R1222_U98 = ~new_P1_R1222_U379 | ~new_P1_R1222_U378;
  assign new_P1_R1222_U99 = ~new_P1_R1222_U386 | ~new_P1_R1222_U385;
  assign new_P1_R1222_U100 = ~new_P1_R1222_U393 | ~new_P1_R1222_U392;
  assign new_P1_R1222_U101 = ~new_P1_R1222_U398 | ~new_P1_R1222_U397;
  assign new_P1_R1222_U102 = ~new_P1_R1222_U407 | ~new_P1_R1222_U406;
  assign new_P1_R1222_U103 = ~new_P1_R1222_U414 | ~new_P1_R1222_U413;
  assign new_P1_R1222_U104 = ~new_P1_R1222_U421 | ~new_P1_R1222_U420;
  assign new_P1_R1222_U105 = ~new_P1_R1222_U428 | ~new_P1_R1222_U427;
  assign new_P1_R1222_U106 = ~new_P1_R1222_U433 | ~new_P1_R1222_U432;
  assign new_P1_R1222_U107 = ~new_P1_R1222_U440 | ~new_P1_R1222_U439;
  assign new_P1_R1222_U108 = ~new_P1_R1222_U447 | ~new_P1_R1222_U446;
  assign new_P1_R1222_U109 = ~new_P1_R1222_U461 | ~new_P1_R1222_U460;
  assign new_P1_R1222_U110 = ~new_P1_R1222_U466 | ~new_P1_R1222_U465;
  assign new_P1_R1222_U111 = ~new_P1_R1222_U473 | ~new_P1_R1222_U472;
  assign new_P1_R1222_U112 = ~new_P1_R1222_U480 | ~new_P1_R1222_U479;
  assign new_P1_R1222_U113 = ~new_P1_R1222_U487 | ~new_P1_R1222_U486;
  assign new_P1_R1222_U114 = ~new_P1_R1222_U494 | ~new_P1_R1222_U493;
  assign new_P1_R1222_U115 = ~new_P1_R1222_U499 | ~new_P1_R1222_U498;
  assign new_P1_R1222_U116 = new_P1_U3458 & new_P1_U3068;
  assign new_P1_R1222_U117 = new_P1_R1222_U188 & new_P1_R1222_U186;
  assign new_P1_R1222_U118 = new_P1_R1222_U193 & new_P1_R1222_U191;
  assign new_P1_R1222_U119 = new_P1_R1222_U200 & new_P1_R1222_U199;
  assign new_P1_R1222_U120 = new_P1_R1222_U23 & new_P1_R1222_U381 & new_P1_R1222_U380;
  assign new_P1_R1222_U121 = new_P1_R1222_U211 & new_P1_R1222_U6;
  assign new_P1_R1222_U122 = new_P1_R1222_U219 & new_P1_R1222_U217;
  assign new_P1_R1222_U123 = new_P1_R1222_U35 & new_P1_R1222_U388 & new_P1_R1222_U387;
  assign new_P1_R1222_U124 = new_P1_R1222_U225 & new_P1_R1222_U4;
  assign new_P1_R1222_U125 = new_P1_R1222_U233 & new_P1_R1222_U180;
  assign new_P1_R1222_U126 = new_P1_R1222_U203 & new_P1_R1222_U7;
  assign new_P1_R1222_U127 = new_P1_R1222_U238 & new_P1_R1222_U170;
  assign new_P1_R1222_U128 = new_P1_R1222_U249 & new_P1_R1222_U8;
  assign new_P1_R1222_U129 = new_P1_R1222_U247 & new_P1_R1222_U171;
  assign new_P1_R1222_U130 = new_P1_R1222_U267 & new_P1_R1222_U266;
  assign new_P1_R1222_U131 = new_P1_R1222_U10 & new_P1_R1222_U281;
  assign new_P1_R1222_U132 = new_P1_R1222_U284 & new_P1_R1222_U279;
  assign new_P1_R1222_U133 = new_P1_R1222_U300 & new_P1_R1222_U297;
  assign new_P1_R1222_U134 = new_P1_R1222_U367 & new_P1_R1222_U301;
  assign new_P1_R1222_U135 = new_P1_R1222_U159 & new_P1_R1222_U277;
  assign new_P1_R1222_U136 = new_P1_R1222_U81 & new_P1_R1222_U454 & new_P1_R1222_U453;
  assign new_P1_R1222_U137 = new_P1_R1222_U60 & new_P1_R1222_U468 & new_P1_R1222_U467;
  assign new_P1_R1222_U138 = new_P1_R1222_U333 & new_P1_R1222_U9;
  assign new_P1_R1222_U139 = new_P1_R1222_U171 & new_P1_R1222_U489 & new_P1_R1222_U488;
  assign new_P1_R1222_U140 = new_P1_R1222_U342 & new_P1_R1222_U8;
  assign new_P1_R1222_U141 = new_P1_R1222_U170 & new_P1_R1222_U501 & new_P1_R1222_U500;
  assign new_P1_R1222_U142 = new_P1_R1222_U349 & new_P1_R1222_U7;
  assign new_P1_R1222_U143 = ~new_P1_R1222_U119 | ~new_P1_R1222_U201;
  assign new_P1_R1222_U144 = ~new_P1_R1222_U216 | ~new_P1_R1222_U228;
  assign new_P1_R1222_U145 = ~new_P1_U3055;
  assign new_P1_R1222_U146 = ~new_P1_U3985;
  assign new_P1_R1222_U147 = new_P1_R1222_U402 & new_P1_R1222_U401;
  assign new_P1_R1222_U148 = ~new_P1_R1222_U363 | ~new_P1_R1222_U303 | ~new_P1_R1222_U168;
  assign new_P1_R1222_U149 = new_P1_R1222_U409 & new_P1_R1222_U408;
  assign new_P1_R1222_U150 = ~new_P1_R1222_U134 | ~new_P1_R1222_U369 | ~new_P1_R1222_U368;
  assign new_P1_R1222_U151 = new_P1_R1222_U416 & new_P1_R1222_U415;
  assign new_P1_R1222_U152 = ~new_P1_R1222_U87 | ~new_P1_R1222_U364 | ~new_P1_R1222_U298;
  assign new_P1_R1222_U153 = new_P1_R1222_U423 & new_P1_R1222_U422;
  assign new_P1_R1222_U154 = ~new_P1_R1222_U292 | ~new_P1_R1222_U291;
  assign new_P1_R1222_U155 = new_P1_R1222_U435 & new_P1_R1222_U434;
  assign new_P1_R1222_U156 = ~new_P1_R1222_U288 | ~new_P1_R1222_U287;
  assign new_P1_R1222_U157 = new_P1_R1222_U442 & new_P1_R1222_U441;
  assign new_P1_R1222_U158 = ~new_P1_R1222_U132 | ~new_P1_R1222_U283;
  assign new_P1_R1222_U159 = new_P1_R1222_U449 & new_P1_R1222_U448;
  assign new_P1_R1222_U160 = ~new_P1_R1222_U44 | ~new_P1_R1222_U326;
  assign new_P1_R1222_U161 = ~new_P1_R1222_U130 | ~new_P1_R1222_U268;
  assign new_P1_R1222_U162 = new_P1_R1222_U475 & new_P1_R1222_U474;
  assign new_P1_R1222_U163 = ~new_P1_R1222_U256 | ~new_P1_R1222_U255;
  assign new_P1_R1222_U164 = new_P1_R1222_U482 & new_P1_R1222_U481;
  assign new_P1_R1222_U165 = ~new_P1_R1222_U252 | ~new_P1_R1222_U251;
  assign new_P1_R1222_U166 = ~new_P1_R1222_U242 | ~new_P1_R1222_U241;
  assign new_P1_R1222_U167 = ~new_P1_R1222_U366 | ~new_P1_R1222_U365;
  assign new_P1_R1222_U168 = ~new_P1_U3054 | ~new_P1_R1222_U150;
  assign new_P1_R1222_U169 = ~new_P1_R1222_U35;
  assign new_P1_R1222_U170 = ~new_P1_U3479 | ~new_P1_U3083;
  assign new_P1_R1222_U171 = ~new_P1_U3072 | ~new_P1_U3488;
  assign new_P1_R1222_U172 = ~new_P1_U3058 | ~new_P1_U3977;
  assign new_P1_R1222_U173 = ~new_P1_R1222_U69;
  assign new_P1_R1222_U174 = ~new_P1_R1222_U78;
  assign new_P1_R1222_U175 = ~new_P1_U3065 | ~new_P1_U3978;
  assign new_P1_R1222_U176 = ~new_P1_R1222_U62;
  assign new_P1_R1222_U177 = new_P1_U3067 | new_P1_U3467;
  assign new_P1_R1222_U178 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1222_U179 = new_P1_U3461 | new_P1_U3064;
  assign new_P1_R1222_U180 = new_P1_U3458 | new_P1_U3068;
  assign new_P1_R1222_U181 = ~new_P1_R1222_U32;
  assign new_P1_R1222_U182 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1222_U183 = ~new_P1_R1222_U43;
  assign new_P1_R1222_U184 = ~new_P1_R1222_U44;
  assign new_P1_R1222_U185 = ~new_P1_R1222_U43 | ~new_P1_R1222_U44;
  assign new_P1_R1222_U186 = ~new_P1_R1222_U116 | ~new_P1_R1222_U179;
  assign new_P1_R1222_U187 = ~new_P1_R1222_U5 | ~new_P1_R1222_U185;
  assign new_P1_R1222_U188 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1222_U189 = ~new_P1_R1222_U117 | ~new_P1_R1222_U187;
  assign new_P1_R1222_U190 = ~new_P1_R1222_U36 | ~new_P1_R1222_U35;
  assign new_P1_R1222_U191 = ~new_P1_U3067 | ~new_P1_R1222_U190;
  assign new_P1_R1222_U192 = ~new_P1_R1222_U4 | ~new_P1_R1222_U189;
  assign new_P1_R1222_U193 = ~new_P1_U3467 | ~new_P1_R1222_U169;
  assign new_P1_R1222_U194 = ~new_P1_R1222_U42;
  assign new_P1_R1222_U195 = new_P1_U3070 | new_P1_U3473;
  assign new_P1_R1222_U196 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1222_U197 = ~new_P1_R1222_U23;
  assign new_P1_R1222_U198 = ~new_P1_R1222_U24 | ~new_P1_R1222_U23;
  assign new_P1_R1222_U199 = ~new_P1_U3070 | ~new_P1_R1222_U198;
  assign new_P1_R1222_U200 = ~new_P1_U3473 | ~new_P1_R1222_U197;
  assign new_P1_R1222_U201 = ~new_P1_R1222_U6 | ~new_P1_R1222_U42;
  assign new_P1_R1222_U202 = ~new_P1_R1222_U143;
  assign new_P1_R1222_U203 = new_P1_U3476 | new_P1_U3084;
  assign new_P1_R1222_U204 = ~new_P1_R1222_U203 | ~new_P1_R1222_U143;
  assign new_P1_R1222_U205 = ~new_P1_R1222_U41;
  assign new_P1_R1222_U206 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1222_U207 = new_P1_U3470 | new_P1_U3071;
  assign new_P1_R1222_U208 = ~new_P1_R1222_U207 | ~new_P1_R1222_U42;
  assign new_P1_R1222_U209 = ~new_P1_R1222_U120 | ~new_P1_R1222_U208;
  assign new_P1_R1222_U210 = ~new_P1_R1222_U194 | ~new_P1_R1222_U23;
  assign new_P1_R1222_U211 = ~new_P1_U3473 | ~new_P1_U3070;
  assign new_P1_R1222_U212 = ~new_P1_R1222_U121 | ~new_P1_R1222_U210;
  assign new_P1_R1222_U213 = new_P1_U3071 | new_P1_U3470;
  assign new_P1_R1222_U214 = ~new_P1_R1222_U184 | ~new_P1_R1222_U180;
  assign new_P1_R1222_U215 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1222_U216 = ~new_P1_R1222_U46;
  assign new_P1_R1222_U217 = ~new_P1_R1222_U183 | ~new_P1_R1222_U5;
  assign new_P1_R1222_U218 = ~new_P1_R1222_U46 | ~new_P1_R1222_U179;
  assign new_P1_R1222_U219 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1222_U220 = ~new_P1_R1222_U45;
  assign new_P1_R1222_U221 = new_P1_U3464 | new_P1_U3060;
  assign new_P1_R1222_U222 = ~new_P1_R1222_U221 | ~new_P1_R1222_U45;
  assign new_P1_R1222_U223 = ~new_P1_R1222_U123 | ~new_P1_R1222_U222;
  assign new_P1_R1222_U224 = ~new_P1_R1222_U220 | ~new_P1_R1222_U35;
  assign new_P1_R1222_U225 = ~new_P1_U3467 | ~new_P1_U3067;
  assign new_P1_R1222_U226 = ~new_P1_R1222_U124 | ~new_P1_R1222_U224;
  assign new_P1_R1222_U227 = new_P1_U3060 | new_P1_U3464;
  assign new_P1_R1222_U228 = ~new_P1_R1222_U183 | ~new_P1_R1222_U180;
  assign new_P1_R1222_U229 = ~new_P1_R1222_U144;
  assign new_P1_R1222_U230 = ~new_P1_U3064 | ~new_P1_U3461;
  assign new_P1_R1222_U231 = ~new_P1_R1222_U43 | ~new_P1_R1222_U44 | ~new_P1_R1222_U400 | ~new_P1_R1222_U399;
  assign new_P1_R1222_U232 = ~new_P1_R1222_U44 | ~new_P1_R1222_U43;
  assign new_P1_R1222_U233 = ~new_P1_U3068 | ~new_P1_U3458;
  assign new_P1_R1222_U234 = ~new_P1_R1222_U125 | ~new_P1_R1222_U232;
  assign new_P1_R1222_U235 = new_P1_U3083 | new_P1_U3479;
  assign new_P1_R1222_U236 = new_P1_U3062 | new_P1_U3482;
  assign new_P1_R1222_U237 = ~new_P1_R1222_U176 | ~new_P1_R1222_U7;
  assign new_P1_R1222_U238 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1222_U239 = ~new_P1_R1222_U127 | ~new_P1_R1222_U237;
  assign new_P1_R1222_U240 = new_P1_U3482 | new_P1_U3062;
  assign new_P1_R1222_U241 = ~new_P1_R1222_U126 | ~new_P1_R1222_U143;
  assign new_P1_R1222_U242 = ~new_P1_R1222_U240 | ~new_P1_R1222_U239;
  assign new_P1_R1222_U243 = ~new_P1_R1222_U166;
  assign new_P1_R1222_U244 = new_P1_U3080 | new_P1_U3491;
  assign new_P1_R1222_U245 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1222_U246 = ~new_P1_R1222_U173 | ~new_P1_R1222_U8;
  assign new_P1_R1222_U247 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1222_U248 = ~new_P1_R1222_U129 | ~new_P1_R1222_U246;
  assign new_P1_R1222_U249 = new_P1_U3485 | new_P1_U3063;
  assign new_P1_R1222_U250 = new_P1_U3491 | new_P1_U3080;
  assign new_P1_R1222_U251 = ~new_P1_R1222_U128 | ~new_P1_R1222_U166;
  assign new_P1_R1222_U252 = ~new_P1_R1222_U250 | ~new_P1_R1222_U248;
  assign new_P1_R1222_U253 = ~new_P1_R1222_U165;
  assign new_P1_R1222_U254 = new_P1_U3494 | new_P1_U3079;
  assign new_P1_R1222_U255 = ~new_P1_R1222_U254 | ~new_P1_R1222_U165;
  assign new_P1_R1222_U256 = ~new_P1_U3079 | ~new_P1_U3494;
  assign new_P1_R1222_U257 = ~new_P1_R1222_U163;
  assign new_P1_R1222_U258 = new_P1_U3497 | new_P1_U3074;
  assign new_P1_R1222_U259 = ~new_P1_R1222_U258 | ~new_P1_R1222_U163;
  assign new_P1_R1222_U260 = ~new_P1_U3074 | ~new_P1_U3497;
  assign new_P1_R1222_U261 = ~new_P1_R1222_U93;
  assign new_P1_R1222_U262 = new_P1_U3069 | new_P1_U3503;
  assign new_P1_R1222_U263 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1222_U264 = ~new_P1_R1222_U60;
  assign new_P1_R1222_U265 = ~new_P1_R1222_U61 | ~new_P1_R1222_U60;
  assign new_P1_R1222_U266 = ~new_P1_U3069 | ~new_P1_R1222_U265;
  assign new_P1_R1222_U267 = ~new_P1_U3503 | ~new_P1_R1222_U264;
  assign new_P1_R1222_U268 = ~new_P1_R1222_U9 | ~new_P1_R1222_U93;
  assign new_P1_R1222_U269 = ~new_P1_R1222_U161;
  assign new_P1_R1222_U270 = new_P1_U3076 | new_P1_U3982;
  assign new_P1_R1222_U271 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1222_U272 = new_P1_U3075 | new_P1_U3981;
  assign new_P1_R1222_U273 = ~new_P1_R1222_U81;
  assign new_P1_R1222_U274 = ~new_P1_U3982 | ~new_P1_R1222_U273;
  assign new_P1_R1222_U275 = ~new_P1_R1222_U274 | ~new_P1_R1222_U91;
  assign new_P1_R1222_U276 = ~new_P1_R1222_U81 | ~new_P1_R1222_U82;
  assign new_P1_R1222_U277 = ~new_P1_R1222_U276 | ~new_P1_R1222_U275;
  assign new_P1_R1222_U278 = ~new_P1_R1222_U174 | ~new_P1_R1222_U10;
  assign new_P1_R1222_U279 = ~new_P1_U3075 | ~new_P1_U3981;
  assign new_P1_R1222_U280 = ~new_P1_R1222_U277 | ~new_P1_R1222_U278;
  assign new_P1_R1222_U281 = new_P1_U3506 | new_P1_U3082;
  assign new_P1_R1222_U282 = new_P1_U3981 | new_P1_U3075;
  assign new_P1_R1222_U283 = ~new_P1_R1222_U131 | ~new_P1_R1222_U272 | ~new_P1_R1222_U161;
  assign new_P1_R1222_U284 = ~new_P1_R1222_U282 | ~new_P1_R1222_U280;
  assign new_P1_R1222_U285 = ~new_P1_R1222_U158;
  assign new_P1_R1222_U286 = new_P1_U3980 | new_P1_U3061;
  assign new_P1_R1222_U287 = ~new_P1_R1222_U286 | ~new_P1_R1222_U158;
  assign new_P1_R1222_U288 = ~new_P1_U3061 | ~new_P1_U3980;
  assign new_P1_R1222_U289 = ~new_P1_R1222_U156;
  assign new_P1_R1222_U290 = new_P1_U3979 | new_P1_U3066;
  assign new_P1_R1222_U291 = ~new_P1_R1222_U290 | ~new_P1_R1222_U156;
  assign new_P1_R1222_U292 = ~new_P1_U3066 | ~new_P1_U3979;
  assign new_P1_R1222_U293 = ~new_P1_R1222_U154;
  assign new_P1_R1222_U294 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1222_U295 = ~new_P1_R1222_U175 | ~new_P1_R1222_U172;
  assign new_P1_R1222_U296 = ~new_P1_R1222_U87;
  assign new_P1_R1222_U297 = new_P1_U3978 | new_P1_U3065;
  assign new_P1_R1222_U298 = ~new_P1_R1222_U167 | ~new_P1_R1222_U154 | ~new_P1_R1222_U297;
  assign new_P1_R1222_U299 = ~new_P1_R1222_U152;
  assign new_P1_R1222_U300 = new_P1_U3975 | new_P1_U3053;
  assign new_P1_R1222_U301 = ~new_P1_U3053 | ~new_P1_U3975;
  assign new_P1_R1222_U302 = ~new_P1_R1222_U150;
  assign new_P1_R1222_U303 = ~new_P1_U3974 | ~new_P1_R1222_U150;
  assign new_P1_R1222_U304 = ~new_P1_R1222_U148;
  assign new_P1_R1222_U305 = ~new_P1_R1222_U297 | ~new_P1_R1222_U154;
  assign new_P1_R1222_U306 = ~new_P1_R1222_U90;
  assign new_P1_R1222_U307 = new_P1_U3977 | new_P1_U3058;
  assign new_P1_R1222_U308 = ~new_P1_R1222_U307 | ~new_P1_R1222_U90;
  assign new_P1_R1222_U309 = ~new_P1_R1222_U153 | ~new_P1_R1222_U308 | ~new_P1_R1222_U172;
  assign new_P1_R1222_U310 = ~new_P1_R1222_U306 | ~new_P1_R1222_U172;
  assign new_P1_R1222_U311 = ~new_P1_U3976 | ~new_P1_U3057;
  assign new_P1_R1222_U312 = ~new_P1_R1222_U167 | ~new_P1_R1222_U310 | ~new_P1_R1222_U311;
  assign new_P1_R1222_U313 = new_P1_U3058 | new_P1_U3977;
  assign new_P1_R1222_U314 = ~new_P1_R1222_U281 | ~new_P1_R1222_U161;
  assign new_P1_R1222_U315 = ~new_P1_R1222_U92;
  assign new_P1_R1222_U316 = ~new_P1_R1222_U10 | ~new_P1_R1222_U92;
  assign new_P1_R1222_U317 = ~new_P1_R1222_U135 | ~new_P1_R1222_U316;
  assign new_P1_R1222_U318 = ~new_P1_R1222_U316 | ~new_P1_R1222_U277;
  assign new_P1_R1222_U319 = ~new_P1_R1222_U452 | ~new_P1_R1222_U318;
  assign new_P1_R1222_U320 = new_P1_U3508 | new_P1_U3081;
  assign new_P1_R1222_U321 = ~new_P1_R1222_U320 | ~new_P1_R1222_U92;
  assign new_P1_R1222_U322 = ~new_P1_R1222_U136 | ~new_P1_R1222_U321;
  assign new_P1_R1222_U323 = ~new_P1_R1222_U315 | ~new_P1_R1222_U81;
  assign new_P1_R1222_U324 = ~new_P1_U3076 | ~new_P1_U3982;
  assign new_P1_R1222_U325 = ~new_P1_R1222_U10 | ~new_P1_R1222_U324 | ~new_P1_R1222_U323;
  assign new_P1_R1222_U326 = new_P1_U3455 | new_P1_U3078;
  assign new_P1_R1222_U327 = ~new_P1_R1222_U160;
  assign new_P1_R1222_U328 = new_P1_U3081 | new_P1_U3508;
  assign new_P1_R1222_U329 = new_P1_U3500 | new_P1_U3073;
  assign new_P1_R1222_U330 = ~new_P1_R1222_U329 | ~new_P1_R1222_U93;
  assign new_P1_R1222_U331 = ~new_P1_R1222_U137 | ~new_P1_R1222_U330;
  assign new_P1_R1222_U332 = ~new_P1_R1222_U261 | ~new_P1_R1222_U60;
  assign new_P1_R1222_U333 = ~new_P1_U3503 | ~new_P1_U3069;
  assign new_P1_R1222_U334 = ~new_P1_R1222_U138 | ~new_P1_R1222_U332;
  assign new_P1_R1222_U335 = new_P1_U3073 | new_P1_U3500;
  assign new_P1_R1222_U336 = ~new_P1_R1222_U249 | ~new_P1_R1222_U166;
  assign new_P1_R1222_U337 = ~new_P1_R1222_U94;
  assign new_P1_R1222_U338 = new_P1_U3488 | new_P1_U3072;
  assign new_P1_R1222_U339 = ~new_P1_R1222_U338 | ~new_P1_R1222_U94;
  assign new_P1_R1222_U340 = ~new_P1_R1222_U139 | ~new_P1_R1222_U339;
  assign new_P1_R1222_U341 = ~new_P1_R1222_U337 | ~new_P1_R1222_U171;
  assign new_P1_R1222_U342 = ~new_P1_U3080 | ~new_P1_U3491;
  assign new_P1_R1222_U343 = ~new_P1_R1222_U140 | ~new_P1_R1222_U341;
  assign new_P1_R1222_U344 = new_P1_U3072 | new_P1_U3488;
  assign new_P1_R1222_U345 = new_P1_U3479 | new_P1_U3083;
  assign new_P1_R1222_U346 = ~new_P1_R1222_U345 | ~new_P1_R1222_U41;
  assign new_P1_R1222_U347 = ~new_P1_R1222_U141 | ~new_P1_R1222_U346;
  assign new_P1_R1222_U348 = ~new_P1_R1222_U205 | ~new_P1_R1222_U170;
  assign new_P1_R1222_U349 = ~new_P1_U3062 | ~new_P1_U3482;
  assign new_P1_R1222_U350 = ~new_P1_R1222_U142 | ~new_P1_R1222_U348;
  assign new_P1_R1222_U351 = ~new_P1_R1222_U206 | ~new_P1_R1222_U170;
  assign new_P1_R1222_U352 = ~new_P1_R1222_U203 | ~new_P1_R1222_U62;
  assign new_P1_R1222_U353 = ~new_P1_R1222_U213 | ~new_P1_R1222_U23;
  assign new_P1_R1222_U354 = ~new_P1_R1222_U227 | ~new_P1_R1222_U35;
  assign new_P1_R1222_U355 = ~new_P1_R1222_U230 | ~new_P1_R1222_U179;
  assign new_P1_R1222_U356 = ~new_P1_R1222_U313 | ~new_P1_R1222_U172;
  assign new_P1_R1222_U357 = ~new_P1_R1222_U297 | ~new_P1_R1222_U175;
  assign new_P1_R1222_U358 = ~new_P1_R1222_U328 | ~new_P1_R1222_U81;
  assign new_P1_R1222_U359 = ~new_P1_R1222_U281 | ~new_P1_R1222_U78;
  assign new_P1_R1222_U360 = ~new_P1_R1222_U335 | ~new_P1_R1222_U60;
  assign new_P1_R1222_U361 = ~new_P1_R1222_U344 | ~new_P1_R1222_U171;
  assign new_P1_R1222_U362 = ~new_P1_R1222_U249 | ~new_P1_R1222_U69;
  assign new_P1_R1222_U363 = ~new_P1_U3974 | ~new_P1_U3054;
  assign new_P1_R1222_U364 = ~new_P1_R1222_U295 | ~new_P1_R1222_U167;
  assign new_P1_R1222_U365 = ~new_P1_U3057 | ~new_P1_R1222_U294;
  assign new_P1_R1222_U366 = ~new_P1_U3976 | ~new_P1_R1222_U294;
  assign new_P1_R1222_U367 = ~new_P1_R1222_U300 | ~new_P1_R1222_U295 | ~new_P1_R1222_U167;
  assign new_P1_R1222_U368 = ~new_P1_R1222_U133 | ~new_P1_R1222_U154 | ~new_P1_R1222_U167;
  assign new_P1_R1222_U369 = ~new_P1_R1222_U296 | ~new_P1_R1222_U300;
  assign new_P1_R1222_U370 = ~new_P1_U3083 | ~new_P1_R1222_U40;
  assign new_P1_R1222_U371 = ~new_P1_U3479 | ~new_P1_R1222_U39;
  assign new_P1_R1222_U372 = ~new_P1_R1222_U371 | ~new_P1_R1222_U370;
  assign new_P1_R1222_U373 = ~new_P1_R1222_U351 | ~new_P1_R1222_U41;
  assign new_P1_R1222_U374 = ~new_P1_R1222_U372 | ~new_P1_R1222_U205;
  assign new_P1_R1222_U375 = ~new_P1_U3084 | ~new_P1_R1222_U37;
  assign new_P1_R1222_U376 = ~new_P1_U3476 | ~new_P1_R1222_U38;
  assign new_P1_R1222_U377 = ~new_P1_R1222_U376 | ~new_P1_R1222_U375;
  assign new_P1_R1222_U378 = ~new_P1_R1222_U352 | ~new_P1_R1222_U143;
  assign new_P1_R1222_U379 = ~new_P1_R1222_U202 | ~new_P1_R1222_U377;
  assign new_P1_R1222_U380 = ~new_P1_U3070 | ~new_P1_R1222_U24;
  assign new_P1_R1222_U381 = ~new_P1_U3473 | ~new_P1_R1222_U22;
  assign new_P1_R1222_U382 = ~new_P1_U3071 | ~new_P1_R1222_U20;
  assign new_P1_R1222_U383 = ~new_P1_U3470 | ~new_P1_R1222_U21;
  assign new_P1_R1222_U384 = ~new_P1_R1222_U383 | ~new_P1_R1222_U382;
  assign new_P1_R1222_U385 = ~new_P1_R1222_U353 | ~new_P1_R1222_U42;
  assign new_P1_R1222_U386 = ~new_P1_R1222_U384 | ~new_P1_R1222_U194;
  assign new_P1_R1222_U387 = ~new_P1_U3067 | ~new_P1_R1222_U36;
  assign new_P1_R1222_U388 = ~new_P1_U3467 | ~new_P1_R1222_U27;
  assign new_P1_R1222_U389 = ~new_P1_U3060 | ~new_P1_R1222_U25;
  assign new_P1_R1222_U390 = ~new_P1_U3464 | ~new_P1_R1222_U26;
  assign new_P1_R1222_U391 = ~new_P1_R1222_U390 | ~new_P1_R1222_U389;
  assign new_P1_R1222_U392 = ~new_P1_R1222_U354 | ~new_P1_R1222_U45;
  assign new_P1_R1222_U393 = ~new_P1_R1222_U391 | ~new_P1_R1222_U220;
  assign new_P1_R1222_U394 = ~new_P1_U3064 | ~new_P1_R1222_U33;
  assign new_P1_R1222_U395 = ~new_P1_U3461 | ~new_P1_R1222_U34;
  assign new_P1_R1222_U396 = ~new_P1_R1222_U395 | ~new_P1_R1222_U394;
  assign new_P1_R1222_U397 = ~new_P1_R1222_U355 | ~new_P1_R1222_U144;
  assign new_P1_R1222_U398 = ~new_P1_R1222_U229 | ~new_P1_R1222_U396;
  assign new_P1_R1222_U399 = ~new_P1_U3068 | ~new_P1_R1222_U28;
  assign new_P1_R1222_U400 = ~new_P1_U3458 | ~new_P1_R1222_U29;
  assign new_P1_R1222_U401 = ~new_P1_U3055 | ~new_P1_R1222_U146;
  assign new_P1_R1222_U402 = ~new_P1_U3985 | ~new_P1_R1222_U145;
  assign new_P1_R1222_U403 = ~new_P1_U3055 | ~new_P1_R1222_U146;
  assign new_P1_R1222_U404 = ~new_P1_U3985 | ~new_P1_R1222_U145;
  assign new_P1_R1222_U405 = ~new_P1_R1222_U404 | ~new_P1_R1222_U403;
  assign new_P1_R1222_U406 = ~new_P1_R1222_U147 | ~new_P1_R1222_U148;
  assign new_P1_R1222_U407 = ~new_P1_R1222_U304 | ~new_P1_R1222_U405;
  assign new_P1_R1222_U408 = ~new_P1_U3054 | ~new_P1_R1222_U89;
  assign new_P1_R1222_U409 = ~new_P1_U3974 | ~new_P1_R1222_U88;
  assign new_P1_R1222_U410 = ~new_P1_U3054 | ~new_P1_R1222_U89;
  assign new_P1_R1222_U411 = ~new_P1_U3974 | ~new_P1_R1222_U88;
  assign new_P1_R1222_U412 = ~new_P1_R1222_U411 | ~new_P1_R1222_U410;
  assign new_P1_R1222_U413 = ~new_P1_R1222_U149 | ~new_P1_R1222_U150;
  assign new_P1_R1222_U414 = ~new_P1_R1222_U302 | ~new_P1_R1222_U412;
  assign new_P1_R1222_U415 = ~new_P1_U3053 | ~new_P1_R1222_U47;
  assign new_P1_R1222_U416 = ~new_P1_U3975 | ~new_P1_R1222_U48;
  assign new_P1_R1222_U417 = ~new_P1_U3053 | ~new_P1_R1222_U47;
  assign new_P1_R1222_U418 = ~new_P1_U3975 | ~new_P1_R1222_U48;
  assign new_P1_R1222_U419 = ~new_P1_R1222_U418 | ~new_P1_R1222_U417;
  assign new_P1_R1222_U420 = ~new_P1_R1222_U151 | ~new_P1_R1222_U152;
  assign new_P1_R1222_U421 = ~new_P1_R1222_U299 | ~new_P1_R1222_U419;
  assign new_P1_R1222_U422 = ~new_P1_U3057 | ~new_P1_R1222_U50;
  assign new_P1_R1222_U423 = ~new_P1_U3976 | ~new_P1_R1222_U49;
  assign new_P1_R1222_U424 = ~new_P1_U3058 | ~new_P1_R1222_U51;
  assign new_P1_R1222_U425 = ~new_P1_U3977 | ~new_P1_R1222_U52;
  assign new_P1_R1222_U426 = ~new_P1_R1222_U425 | ~new_P1_R1222_U424;
  assign new_P1_R1222_U427 = ~new_P1_R1222_U356 | ~new_P1_R1222_U90;
  assign new_P1_R1222_U428 = ~new_P1_R1222_U426 | ~new_P1_R1222_U306;
  assign new_P1_R1222_U429 = ~new_P1_U3065 | ~new_P1_R1222_U53;
  assign new_P1_R1222_U430 = ~new_P1_U3978 | ~new_P1_R1222_U54;
  assign new_P1_R1222_U431 = ~new_P1_R1222_U430 | ~new_P1_R1222_U429;
  assign new_P1_R1222_U432 = ~new_P1_R1222_U357 | ~new_P1_R1222_U154;
  assign new_P1_R1222_U433 = ~new_P1_R1222_U293 | ~new_P1_R1222_U431;
  assign new_P1_R1222_U434 = ~new_P1_U3066 | ~new_P1_R1222_U85;
  assign new_P1_R1222_U435 = ~new_P1_U3979 | ~new_P1_R1222_U86;
  assign new_P1_R1222_U436 = ~new_P1_U3066 | ~new_P1_R1222_U85;
  assign new_P1_R1222_U437 = ~new_P1_U3979 | ~new_P1_R1222_U86;
  assign new_P1_R1222_U438 = ~new_P1_R1222_U437 | ~new_P1_R1222_U436;
  assign new_P1_R1222_U439 = ~new_P1_R1222_U155 | ~new_P1_R1222_U156;
  assign new_P1_R1222_U440 = ~new_P1_R1222_U289 | ~new_P1_R1222_U438;
  assign new_P1_R1222_U441 = ~new_P1_U3061 | ~new_P1_R1222_U83;
  assign new_P1_R1222_U442 = ~new_P1_U3980 | ~new_P1_R1222_U84;
  assign new_P1_R1222_U443 = ~new_P1_U3061 | ~new_P1_R1222_U83;
  assign new_P1_R1222_U444 = ~new_P1_U3980 | ~new_P1_R1222_U84;
  assign new_P1_R1222_U445 = ~new_P1_R1222_U444 | ~new_P1_R1222_U443;
  assign new_P1_R1222_U446 = ~new_P1_R1222_U157 | ~new_P1_R1222_U158;
  assign new_P1_R1222_U447 = ~new_P1_R1222_U285 | ~new_P1_R1222_U445;
  assign new_P1_R1222_U448 = ~new_P1_U3075 | ~new_P1_R1222_U55;
  assign new_P1_R1222_U449 = ~new_P1_U3981 | ~new_P1_R1222_U56;
  assign new_P1_R1222_U450 = ~new_P1_U3075 | ~new_P1_R1222_U55;
  assign new_P1_R1222_U451 = ~new_P1_U3981 | ~new_P1_R1222_U56;
  assign new_P1_R1222_U452 = ~new_P1_R1222_U451 | ~new_P1_R1222_U450;
  assign new_P1_R1222_U453 = ~new_P1_U3076 | ~new_P1_R1222_U82;
  assign new_P1_R1222_U454 = ~new_P1_U3982 | ~new_P1_R1222_U91;
  assign new_P1_R1222_U455 = ~new_P1_R1222_U181 | ~new_P1_R1222_U160;
  assign new_P1_R1222_U456 = ~new_P1_R1222_U327 | ~new_P1_R1222_U32;
  assign new_P1_R1222_U457 = ~new_P1_U3081 | ~new_P1_R1222_U79;
  assign new_P1_R1222_U458 = ~new_P1_U3508 | ~new_P1_R1222_U80;
  assign new_P1_R1222_U459 = ~new_P1_R1222_U458 | ~new_P1_R1222_U457;
  assign new_P1_R1222_U460 = ~new_P1_R1222_U358 | ~new_P1_R1222_U92;
  assign new_P1_R1222_U461 = ~new_P1_R1222_U459 | ~new_P1_R1222_U315;
  assign new_P1_R1222_U462 = ~new_P1_U3082 | ~new_P1_R1222_U76;
  assign new_P1_R1222_U463 = ~new_P1_U3506 | ~new_P1_R1222_U77;
  assign new_P1_R1222_U464 = ~new_P1_R1222_U463 | ~new_P1_R1222_U462;
  assign new_P1_R1222_U465 = ~new_P1_R1222_U359 | ~new_P1_R1222_U161;
  assign new_P1_R1222_U466 = ~new_P1_R1222_U269 | ~new_P1_R1222_U464;
  assign new_P1_R1222_U467 = ~new_P1_U3069 | ~new_P1_R1222_U61;
  assign new_P1_R1222_U468 = ~new_P1_U3503 | ~new_P1_R1222_U59;
  assign new_P1_R1222_U469 = ~new_P1_U3073 | ~new_P1_R1222_U57;
  assign new_P1_R1222_U470 = ~new_P1_U3500 | ~new_P1_R1222_U58;
  assign new_P1_R1222_U471 = ~new_P1_R1222_U470 | ~new_P1_R1222_U469;
  assign new_P1_R1222_U472 = ~new_P1_R1222_U360 | ~new_P1_R1222_U93;
  assign new_P1_R1222_U473 = ~new_P1_R1222_U471 | ~new_P1_R1222_U261;
  assign new_P1_R1222_U474 = ~new_P1_U3074 | ~new_P1_R1222_U74;
  assign new_P1_R1222_U475 = ~new_P1_U3497 | ~new_P1_R1222_U75;
  assign new_P1_R1222_U476 = ~new_P1_U3074 | ~new_P1_R1222_U74;
  assign new_P1_R1222_U477 = ~new_P1_U3497 | ~new_P1_R1222_U75;
  assign new_P1_R1222_U478 = ~new_P1_R1222_U477 | ~new_P1_R1222_U476;
  assign new_P1_R1222_U479 = ~new_P1_R1222_U162 | ~new_P1_R1222_U163;
  assign new_P1_R1222_U480 = ~new_P1_R1222_U257 | ~new_P1_R1222_U478;
  assign new_P1_R1222_U481 = ~new_P1_U3079 | ~new_P1_R1222_U72;
  assign new_P1_R1222_U482 = ~new_P1_U3494 | ~new_P1_R1222_U73;
  assign new_P1_R1222_U483 = ~new_P1_U3079 | ~new_P1_R1222_U72;
  assign new_P1_R1222_U484 = ~new_P1_U3494 | ~new_P1_R1222_U73;
  assign new_P1_R1222_U485 = ~new_P1_R1222_U484 | ~new_P1_R1222_U483;
  assign new_P1_R1222_U486 = ~new_P1_R1222_U164 | ~new_P1_R1222_U165;
  assign new_P1_R1222_U487 = ~new_P1_R1222_U253 | ~new_P1_R1222_U485;
  assign new_P1_R1222_U488 = ~new_P1_U3080 | ~new_P1_R1222_U70;
  assign new_P1_R1222_U489 = ~new_P1_U3491 | ~new_P1_R1222_U71;
  assign new_P1_R1222_U490 = ~new_P1_U3072 | ~new_P1_R1222_U65;
  assign new_P1_R1222_U491 = ~new_P1_U3488 | ~new_P1_R1222_U66;
  assign new_P1_R1222_U492 = ~new_P1_R1222_U491 | ~new_P1_R1222_U490;
  assign new_P1_R1222_U493 = ~new_P1_R1222_U361 | ~new_P1_R1222_U94;
  assign new_P1_R1222_U494 = ~new_P1_R1222_U492 | ~new_P1_R1222_U337;
  assign new_P1_R1222_U495 = ~new_P1_U3063 | ~new_P1_R1222_U67;
  assign new_P1_R1222_U496 = ~new_P1_U3485 | ~new_P1_R1222_U68;
  assign new_P1_R1222_U497 = ~new_P1_R1222_U496 | ~new_P1_R1222_U495;
  assign new_P1_R1222_U498 = ~new_P1_R1222_U362 | ~new_P1_R1222_U166;
  assign new_P1_R1222_U499 = ~new_P1_R1222_U243 | ~new_P1_R1222_U497;
  assign new_P1_R1222_U500 = ~new_P1_U3062 | ~new_P1_R1222_U63;
  assign new_P1_R1222_U501 = ~new_P1_U3482 | ~new_P1_R1222_U64;
  assign new_P1_R1222_U502 = ~new_P1_U3077 | ~new_P1_R1222_U30;
  assign new_P1_R1222_U503 = ~new_P1_U3450 | ~new_P1_R1222_U31;
  assign new_P2_SUB_594_U6 = ~P2_IR_REG_11_ & ~P2_IR_REG_10_ & ~P2_IR_REG_12_ & ~P2_IR_REG_9_;
  assign new_P2_SUB_594_U7 = ~P2_IR_REG_18_ & ~P2_IR_REG_17_ & ~P2_IR_REG_19_ & ~P2_IR_REG_20_;
  assign new_P2_SUB_594_U8 = new_P2_SUB_594_U135 & new_P2_SUB_594_U51;
  assign new_P2_SUB_594_U9 = new_P2_SUB_594_U133 & new_P2_SUB_594_U101;
  assign new_P2_SUB_594_U10 = new_P2_SUB_594_U132 & new_P2_SUB_594_U47;
  assign new_P2_SUB_594_U11 = new_P2_SUB_594_U131 & new_P2_SUB_594_U48;
  assign new_P2_SUB_594_U12 = new_P2_SUB_594_U129 & new_P2_SUB_594_U104;
  assign new_P2_SUB_594_U13 = new_P2_SUB_594_U128 & new_P2_SUB_594_U35;
  assign new_P2_SUB_594_U14 = new_P2_SUB_594_U127 & new_P2_SUB_594_U45;
  assign new_P2_SUB_594_U15 = new_P2_SUB_594_U125 & new_P2_SUB_594_U107;
  assign new_P2_SUB_594_U16 = new_P2_SUB_594_U124 & new_P2_SUB_594_U41;
  assign new_P2_SUB_594_U17 = new_P2_SUB_594_U123 & new_P2_SUB_594_U42;
  assign new_P2_SUB_594_U18 = new_P2_SUB_594_U121 & new_P2_SUB_594_U110;
  assign new_P2_SUB_594_U19 = new_P2_SUB_594_U120 & new_P2_SUB_594_U36;
  assign new_P2_SUB_594_U20 = new_P2_SUB_594_U119 & new_P2_SUB_594_U76;
  assign new_P2_SUB_594_U21 = new_P2_SUB_594_U64 & new_P2_SUB_594_U138;
  assign new_P2_SUB_594_U22 = new_P2_SUB_594_U117 & new_P2_SUB_594_U38;
  assign new_P2_SUB_594_U23 = new_P2_SUB_594_U116 & new_P2_SUB_594_U33;
  assign new_P2_SUB_594_U24 = new_P2_SUB_594_U99 & new_P2_SUB_594_U89;
  assign new_P2_SUB_594_U25 = new_P2_SUB_594_U98 & new_P2_SUB_594_U30;
  assign new_P2_SUB_594_U26 = new_P2_SUB_594_U97 & new_P2_SUB_594_U31;
  assign new_P2_SUB_594_U27 = new_P2_SUB_594_U95 & new_P2_SUB_594_U92;
  assign new_P2_SUB_594_U28 = new_P2_SUB_594_U94 & new_P2_SUB_594_U29;
  assign new_P2_SUB_594_U29 = ~new_P2_SUB_594_U56 | ~new_P2_SUB_594_U55;
  assign new_P2_SUB_594_U30 = P2_IR_REG_4_ | P2_IR_REG_3_ | P2_IR_REG_2_ | P2_IR_REG_1_ | P2_IR_REG_0_;
  assign new_P2_SUB_594_U31 = ~new_P2_SUB_594_U57 | ~new_P2_SUB_594_U90;
  assign new_P2_SUB_594_U32 = ~P2_IR_REG_7_;
  assign new_P2_SUB_594_U33 = P2_IR_REG_2_ | P2_IR_REG_1_ | P2_IR_REG_0_;
  assign new_P2_SUB_594_U34 = ~P2_IR_REG_3_;
  assign new_P2_SUB_594_U35 = ~new_P2_SUB_594_U59 | ~new_P2_SUB_594_U93;
  assign new_P2_SUB_594_U36 = ~new_P2_SUB_594_U61 | ~new_P2_SUB_594_U105;
  assign new_P2_SUB_594_U37 = ~new_P2_SUB_594_U62 | ~new_P2_SUB_594_U111;
  assign new_P2_SUB_594_U38 = ~new_P2_SUB_594_U113 | ~new_P2_SUB_594_U39;
  assign new_P2_SUB_594_U39 = ~P2_IR_REG_29_;
  assign new_P2_SUB_594_U40 = ~P2_IR_REG_27_;
  assign new_P2_SUB_594_U41 = ~new_P2_SUB_594_U105 | ~new_P2_SUB_594_U7;
  assign new_P2_SUB_594_U42 = ~new_P2_SUB_594_U65 | ~new_P2_SUB_594_U108;
  assign new_P2_SUB_594_U43 = ~P2_IR_REG_24_;
  assign new_P2_SUB_594_U44 = ~P2_IR_REG_23_;
  assign new_P2_SUB_594_U45 = ~new_P2_SUB_594_U66 | ~new_P2_SUB_594_U105;
  assign new_P2_SUB_594_U46 = ~P2_IR_REG_19_;
  assign new_P2_SUB_594_U47 = ~new_P2_SUB_594_U6 | ~new_P2_SUB_594_U93;
  assign new_P2_SUB_594_U48 = ~new_P2_SUB_594_U67 | ~new_P2_SUB_594_U102;
  assign new_P2_SUB_594_U49 = ~P2_IR_REG_16_;
  assign new_P2_SUB_594_U50 = ~P2_IR_REG_15_;
  assign new_P2_SUB_594_U51 = ~new_P2_SUB_594_U68 | ~new_P2_SUB_594_U93;
  assign new_P2_SUB_594_U52 = ~P2_IR_REG_11_;
  assign new_P2_SUB_594_U53 = ~new_P2_SUB_594_U154 | ~new_P2_SUB_594_U153;
  assign new_P2_SUB_594_U54 = ~new_P2_SUB_594_U144 | ~new_P2_SUB_594_U143;
  assign new_P2_SUB_594_U55 = ~P2_IR_REG_0_ & ~P2_IR_REG_1_ & ~P2_IR_REG_2_ & ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_594_U56 = ~P2_IR_REG_8_ & ~P2_IR_REG_7_ & ~P2_IR_REG_5_ & ~P2_IR_REG_6_;
  assign new_P2_SUB_594_U57 = ~P2_IR_REG_5_ & ~P2_IR_REG_6_;
  assign new_P2_SUB_594_U58 = ~P2_IR_REG_14_ & ~P2_IR_REG_15_ & ~P2_IR_REG_13_;
  assign new_P2_SUB_594_U59 = new_P2_SUB_594_U58 & new_P2_SUB_594_U6 & new_P2_SUB_594_U49;
  assign new_P2_SUB_594_U60 = ~P2_IR_REG_22_ & ~P2_IR_REG_23_ & ~P2_IR_REG_21_;
  assign new_P2_SUB_594_U61 = new_P2_SUB_594_U60 & new_P2_SUB_594_U7 & new_P2_SUB_594_U43;
  assign new_P2_SUB_594_U62 = ~P2_IR_REG_28_ & ~P2_IR_REG_27_ & ~P2_IR_REG_25_ & ~P2_IR_REG_26_;
  assign new_P2_SUB_594_U63 = ~P2_IR_REG_25_ & ~P2_IR_REG_26_;
  assign new_P2_SUB_594_U64 = new_P2_SUB_594_U137 & new_P2_SUB_594_U37;
  assign new_P2_SUB_594_U65 = ~P2_IR_REG_21_ & ~P2_IR_REG_22_;
  assign new_P2_SUB_594_U66 = ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign new_P2_SUB_594_U67 = ~P2_IR_REG_13_ & ~P2_IR_REG_14_;
  assign new_P2_SUB_594_U68 = ~P2_IR_REG_10_ & ~P2_IR_REG_9_;
  assign new_P2_SUB_594_U69 = ~P2_IR_REG_9_;
  assign new_P2_SUB_594_U70 = new_P2_SUB_594_U140 & new_P2_SUB_594_U139;
  assign new_P2_SUB_594_U71 = ~P2_IR_REG_5_;
  assign new_P2_SUB_594_U72 = new_P2_SUB_594_U142 & new_P2_SUB_594_U141;
  assign new_P2_SUB_594_U73 = ~P2_IR_REG_31_;
  assign new_P2_SUB_594_U74 = ~P2_IR_REG_30_;
  assign new_P2_SUB_594_U75 = new_P2_SUB_594_U146 & new_P2_SUB_594_U145;
  assign new_P2_SUB_594_U76 = ~new_P2_SUB_594_U63 | ~new_P2_SUB_594_U111;
  assign new_P2_SUB_594_U77 = new_P2_SUB_594_U148 & new_P2_SUB_594_U147;
  assign new_P2_SUB_594_U78 = ~P2_IR_REG_25_;
  assign new_P2_SUB_594_U79 = new_P2_SUB_594_U150 & new_P2_SUB_594_U149;
  assign new_P2_SUB_594_U80 = ~P2_IR_REG_21_;
  assign new_P2_SUB_594_U81 = new_P2_SUB_594_U152 & new_P2_SUB_594_U151;
  assign new_P2_SUB_594_U82 = ~P2_IR_REG_1_;
  assign new_P2_SUB_594_U83 = ~P2_IR_REG_0_;
  assign new_P2_SUB_594_U84 = ~P2_IR_REG_17_;
  assign new_P2_SUB_594_U85 = new_P2_SUB_594_U156 & new_P2_SUB_594_U155;
  assign new_P2_SUB_594_U86 = ~P2_IR_REG_13_;
  assign new_P2_SUB_594_U87 = new_P2_SUB_594_U158 & new_P2_SUB_594_U157;
  assign new_P2_SUB_594_U88 = ~new_P2_SUB_594_U33;
  assign new_P2_SUB_594_U89 = ~new_P2_SUB_594_U88 | ~new_P2_SUB_594_U34;
  assign new_P2_SUB_594_U90 = ~new_P2_SUB_594_U30;
  assign new_P2_SUB_594_U91 = ~new_P2_SUB_594_U31;
  assign new_P2_SUB_594_U92 = ~new_P2_SUB_594_U91 | ~new_P2_SUB_594_U32;
  assign new_P2_SUB_594_U93 = ~new_P2_SUB_594_U29;
  assign new_P2_SUB_594_U94 = ~P2_IR_REG_8_ | ~new_P2_SUB_594_U92;
  assign new_P2_SUB_594_U95 = ~P2_IR_REG_7_ | ~new_P2_SUB_594_U31;
  assign new_P2_SUB_594_U96 = ~new_P2_SUB_594_U90 | ~new_P2_SUB_594_U71;
  assign new_P2_SUB_594_U97 = ~P2_IR_REG_6_ | ~new_P2_SUB_594_U96;
  assign new_P2_SUB_594_U98 = ~P2_IR_REG_4_ | ~new_P2_SUB_594_U89;
  assign new_P2_SUB_594_U99 = ~P2_IR_REG_3_ | ~new_P2_SUB_594_U33;
  assign new_P2_SUB_594_U100 = ~new_P2_SUB_594_U51;
  assign new_P2_SUB_594_U101 = ~new_P2_SUB_594_U100 | ~new_P2_SUB_594_U52;
  assign new_P2_SUB_594_U102 = ~new_P2_SUB_594_U47;
  assign new_P2_SUB_594_U103 = ~new_P2_SUB_594_U48;
  assign new_P2_SUB_594_U104 = ~new_P2_SUB_594_U103 | ~new_P2_SUB_594_U50;
  assign new_P2_SUB_594_U105 = ~new_P2_SUB_594_U35;
  assign new_P2_SUB_594_U106 = ~new_P2_SUB_594_U45;
  assign new_P2_SUB_594_U107 = ~new_P2_SUB_594_U106 | ~new_P2_SUB_594_U46;
  assign new_P2_SUB_594_U108 = ~new_P2_SUB_594_U41;
  assign new_P2_SUB_594_U109 = ~new_P2_SUB_594_U42;
  assign new_P2_SUB_594_U110 = ~new_P2_SUB_594_U109 | ~new_P2_SUB_594_U44;
  assign new_P2_SUB_594_U111 = ~new_P2_SUB_594_U36;
  assign new_P2_SUB_594_U112 = ~new_P2_SUB_594_U76;
  assign new_P2_SUB_594_U113 = ~new_P2_SUB_594_U37;
  assign new_P2_SUB_594_U114 = ~new_P2_SUB_594_U38;
  assign new_P2_SUB_594_U115 = P2_IR_REG_1_ | P2_IR_REG_0_;
  assign new_P2_SUB_594_U116 = ~P2_IR_REG_2_ | ~new_P2_SUB_594_U115;
  assign new_P2_SUB_594_U117 = ~P2_IR_REG_29_ | ~new_P2_SUB_594_U37;
  assign new_P2_SUB_594_U118 = ~new_P2_SUB_594_U111 | ~new_P2_SUB_594_U78;
  assign new_P2_SUB_594_U119 = ~P2_IR_REG_26_ | ~new_P2_SUB_594_U118;
  assign new_P2_SUB_594_U120 = ~P2_IR_REG_24_ | ~new_P2_SUB_594_U110;
  assign new_P2_SUB_594_U121 = ~P2_IR_REG_23_ | ~new_P2_SUB_594_U42;
  assign new_P2_SUB_594_U122 = ~new_P2_SUB_594_U108 | ~new_P2_SUB_594_U80;
  assign new_P2_SUB_594_U123 = ~P2_IR_REG_22_ | ~new_P2_SUB_594_U122;
  assign new_P2_SUB_594_U124 = ~P2_IR_REG_20_ | ~new_P2_SUB_594_U107;
  assign new_P2_SUB_594_U125 = ~P2_IR_REG_19_ | ~new_P2_SUB_594_U45;
  assign new_P2_SUB_594_U126 = ~new_P2_SUB_594_U105 | ~new_P2_SUB_594_U84;
  assign new_P2_SUB_594_U127 = ~P2_IR_REG_18_ | ~new_P2_SUB_594_U126;
  assign new_P2_SUB_594_U128 = ~P2_IR_REG_16_ | ~new_P2_SUB_594_U104;
  assign new_P2_SUB_594_U129 = ~P2_IR_REG_15_ | ~new_P2_SUB_594_U48;
  assign new_P2_SUB_594_U130 = ~new_P2_SUB_594_U102 | ~new_P2_SUB_594_U86;
  assign new_P2_SUB_594_U131 = ~P2_IR_REG_14_ | ~new_P2_SUB_594_U130;
  assign new_P2_SUB_594_U132 = ~P2_IR_REG_12_ | ~new_P2_SUB_594_U101;
  assign new_P2_SUB_594_U133 = ~P2_IR_REG_11_ | ~new_P2_SUB_594_U51;
  assign new_P2_SUB_594_U134 = ~new_P2_SUB_594_U93 | ~new_P2_SUB_594_U69;
  assign new_P2_SUB_594_U135 = ~P2_IR_REG_10_ | ~new_P2_SUB_594_U134;
  assign new_P2_SUB_594_U136 = ~new_P2_SUB_594_U114 | ~new_P2_SUB_594_U74;
  assign new_P2_SUB_594_U137 = ~P2_IR_REG_27_ | ~P2_IR_REG_28_;
  assign new_P2_SUB_594_U138 = ~P2_IR_REG_28_ | ~new_P2_SUB_594_U76;
  assign new_P2_SUB_594_U139 = ~P2_IR_REG_9_ | ~new_P2_SUB_594_U29;
  assign new_P2_SUB_594_U140 = ~new_P2_SUB_594_U93 | ~new_P2_SUB_594_U69;
  assign new_P2_SUB_594_U141 = ~P2_IR_REG_5_ | ~new_P2_SUB_594_U30;
  assign new_P2_SUB_594_U142 = ~new_P2_SUB_594_U90 | ~new_P2_SUB_594_U71;
  assign new_P2_SUB_594_U143 = ~new_P2_SUB_594_U136 | ~new_P2_SUB_594_U73;
  assign new_P2_SUB_594_U144 = ~P2_IR_REG_31_ | ~new_P2_SUB_594_U114 | ~new_P2_SUB_594_U74;
  assign new_P2_SUB_594_U145 = ~P2_IR_REG_30_ | ~new_P2_SUB_594_U38;
  assign new_P2_SUB_594_U146 = ~new_P2_SUB_594_U114 | ~new_P2_SUB_594_U74;
  assign new_P2_SUB_594_U147 = ~P2_IR_REG_27_ | ~new_P2_SUB_594_U76;
  assign new_P2_SUB_594_U148 = ~new_P2_SUB_594_U112 | ~new_P2_SUB_594_U40;
  assign new_P2_SUB_594_U149 = ~P2_IR_REG_25_ | ~new_P2_SUB_594_U36;
  assign new_P2_SUB_594_U150 = ~new_P2_SUB_594_U111 | ~new_P2_SUB_594_U78;
  assign new_P2_SUB_594_U151 = ~P2_IR_REG_21_ | ~new_P2_SUB_594_U41;
  assign new_P2_SUB_594_U152 = ~new_P2_SUB_594_U108 | ~new_P2_SUB_594_U80;
  assign new_P2_SUB_594_U153 = ~P2_IR_REG_1_ | ~new_P2_SUB_594_U83;
  assign new_P2_SUB_594_U154 = ~P2_IR_REG_0_ | ~new_P2_SUB_594_U82;
  assign new_P2_SUB_594_U155 = ~P2_IR_REG_17_ | ~new_P2_SUB_594_U35;
  assign new_P2_SUB_594_U156 = ~new_P2_SUB_594_U105 | ~new_P2_SUB_594_U84;
  assign new_P2_SUB_594_U157 = ~P2_IR_REG_13_ | ~new_P2_SUB_594_U47;
  assign new_P2_SUB_594_U158 = ~new_P2_SUB_594_U102 | ~new_P2_SUB_594_U86;
  assign new_P2_R693_U6 = new_P2_R693_U109 & new_P2_R693_U110 & new_P2_R693_U111;
  assign new_P2_R693_U7 = new_P2_R693_U118 & new_P2_R693_U119;
  assign new_P2_R693_U8 = new_P2_R693_U120 & new_P2_R693_U121;
  assign new_P2_R693_U9 = new_P2_R693_U8 & new_P2_R693_U125 & new_P2_R693_U81 & new_P2_R693_U123;
  assign new_P2_R693_U10 = new_P2_R693_U130 & new_P2_R693_U132 & new_P2_R693_U134 & new_P2_R693_U133;
  assign new_P2_R693_U11 = new_P2_R693_U83 & new_P2_R693_U10;
  assign new_P2_R693_U12 = new_P2_R693_U11 & new_P2_R693_U138;
  assign new_P2_R693_U13 = new_P2_R693_U144 & new_P2_R693_U143;
  assign new_P2_R693_U14 = new_P2_R693_U104 & new_P2_R693_U105 & new_P2_R693_U189;
  assign new_P2_R693_U15 = ~new_P2_U3529;
  assign new_P2_R693_U16 = ~new_P2_U3904;
  assign new_P2_R693_U17 = ~new_P2_U3896;
  assign new_P2_R693_U18 = ~new_P2_U3895;
  assign new_P2_R693_U19 = ~new_P2_U3535;
  assign new_P2_R693_U20 = ~new_P2_U3532;
  assign new_P2_R693_U21 = ~new_P2_U3534;
  assign new_P2_R693_U22 = ~new_P2_U3537;
  assign new_P2_R693_U23 = ~new_P2_U3536;
  assign new_P2_R693_U24 = ~new_P2_U3901;
  assign new_P2_R693_U25 = ~new_P2_U3540;
  assign new_P2_R693_U26 = ~new_P2_U3902;
  assign new_P2_R693_U27 = ~new_P2_U3541;
  assign new_P2_R693_U28 = ~new_P2_U3543;
  assign new_P2_R693_U29 = ~new_P2_U3443;
  assign new_P2_R693_U30 = ~new_P2_U3544;
  assign new_P2_R693_U31 = ~new_P2_U3440;
  assign new_P2_R693_U32 = ~new_P2_U3445;
  assign new_P2_R693_U33 = ~new_P2_U3903;
  assign new_P2_R693_U34 = ~new_P2_U3545;
  assign new_P2_R693_U35 = ~new_P2_U3546;
  assign new_P2_R693_U36 = ~new_P2_U3437;
  assign new_P2_R693_U37 = ~new_P2_U3434;
  assign new_P2_R693_U38 = ~new_P2_U3419;
  assign new_P2_R693_U39 = ~new_P2_U3416;
  assign new_P2_R693_U40 = ~new_P2_U3410;
  assign new_P2_R693_U41 = ~new_P2_U3413;
  assign new_P2_R693_U42 = ~new_P2_U3407;
  assign new_P2_R693_U43 = ~new_P2_U3404;
  assign new_P2_R693_U44 = ~new_P2_U3401;
  assign new_P2_R693_U45 = ~new_P2_U3398;
  assign new_P2_R693_U46 = ~new_P2_U3553;
  assign new_P2_R693_U47 = ~new_P2_U3395;
  assign new_P2_R693_U48 = ~new_P2_U3392;
  assign new_P2_R693_U49 = ~new_P2_U3550;
  assign new_P2_R693_U50 = ~new_P2_U3549;
  assign new_P2_R693_U51 = ~new_P2_U3542;
  assign new_P2_R693_U52 = ~new_P2_U3531;
  assign new_P2_R693_U53 = ~new_P2_U3528;
  assign new_P2_R693_U54 = ~new_P2_U3527;
  assign new_P2_R693_U55 = ~new_P2_U3526;
  assign new_P2_R693_U56 = ~new_P2_U3525;
  assign new_P2_R693_U57 = ~new_P2_U3524;
  assign new_P2_R693_U58 = ~new_P2_U3523;
  assign new_P2_R693_U59 = ~new_P2_U3552;
  assign new_P2_R693_U60 = ~new_P2_U3551;
  assign new_P2_R693_U61 = ~new_P2_U3425;
  assign new_P2_R693_U62 = ~new_P2_U3422;
  assign new_P2_R693_U63 = ~new_P2_U3431;
  assign new_P2_R693_U64 = ~new_P2_U3428;
  assign new_P2_R693_U65 = ~new_P2_U3548;
  assign new_P2_R693_U66 = ~new_P2_U3547;
  assign new_P2_R693_U67 = ~new_P2_U3539;
  assign new_P2_R693_U68 = ~new_P2_U3538;
  assign new_P2_R693_U69 = ~new_P2_U3900;
  assign new_P2_R693_U70 = ~new_P2_U3899;
  assign new_P2_R693_U71 = ~new_P2_U3898;
  assign new_P2_R693_U72 = ~new_P2_U3897;
  assign new_P2_R693_U73 = ~new_P2_U3868;
  assign new_P2_R693_U74 = ~new_P2_U3533;
  assign new_P2_R693_U75 = new_P2_U3532 & new_P2_R693_U16;
  assign new_P2_R693_U76 = new_P2_U3540 & new_P2_R693_U26;
  assign new_P2_R693_U77 = new_P2_U3541 & new_P2_R693_U33;
  assign new_P2_R693_U78 = new_P2_R693_U174 & new_P2_R693_U173;
  assign new_P2_R693_U79 = new_P2_U3443 & new_P2_R693_U30;
  assign new_P2_R693_U80 = new_P2_U3440 & new_P2_R693_U34;
  assign new_P2_R693_U81 = new_P2_R693_U124 & new_P2_R693_U122;
  assign new_P2_R693_U82 = new_P2_U3387 & new_P2_R693_U107;
  assign new_P2_R693_U83 = new_P2_R693_U137 & new_P2_R693_U136 & new_P2_R693_U135;
  assign new_P2_R693_U84 = new_P2_R693_U140 & new_P2_R693_U141;
  assign new_P2_R693_U85 = new_P2_R693_U84 & new_P2_R693_U139;
  assign new_P2_R693_U86 = new_P2_U3542 & new_P2_R693_U47;
  assign new_P2_R693_U87 = new_P2_U3531 & new_P2_R693_U45;
  assign new_P2_R693_U88 = new_P2_R693_U136 & new_P2_R693_U135;
  assign new_P2_R693_U89 = new_P2_R693_U152 & new_P2_R693_U153;
  assign new_P2_R693_U90 = new_P2_R693_U132 & new_P2_R693_U130;
  assign new_P2_R693_U91 = new_P2_R693_U13 & new_P2_R693_U160;
  assign new_P2_R693_U92 = new_P2_R693_U91 & new_P2_R693_U159 & new_P2_R693_U158;
  assign new_P2_R693_U93 = new_P2_U3425 & new_P2_R693_U49;
  assign new_P2_R693_U94 = new_P2_U3422 & new_P2_R693_U60;
  assign new_P2_R693_U95 = new_P2_R693_U163 & new_P2_R693_U97;
  assign new_P2_R693_U96 = new_P2_R693_U95 & new_P2_R693_U164;
  assign new_P2_R693_U97 = new_P2_R693_U166 & new_P2_R693_U165;
  assign new_P2_R693_U98 = new_P2_R693_U128 & new_P2_R693_U127 & new_P2_R693_U177 & new_P2_R693_U176;
  assign new_P2_R693_U99 = new_P2_R693_U181 & new_P2_R693_U180;
  assign new_P2_R693_U100 = new_P2_R693_U188 & new_P2_R693_U187;
  assign new_P2_R693_U101 = new_P2_R693_U100 & new_P2_R693_U6;
  assign new_P2_R693_U102 = new_P2_R693_U103 & new_P2_R693_U191;
  assign new_P2_R693_U103 = new_P2_U3533 & new_P2_R693_U18;
  assign new_P2_R693_U104 = new_P2_R693_U114 & new_P2_R693_U115 & new_P2_R693_U117 & new_P2_R693_U116;
  assign new_P2_R693_U105 = new_P2_R693_U190 & new_P2_R693_U192;
  assign new_P2_R693_U106 = ~new_P2_U3869;
  assign new_P2_R693_U107 = ~new_P2_U3554;
  assign new_P2_R693_U108 = ~new_P2_R693_U113 | ~new_P2_R693_U193;
  assign new_P2_R693_U109 = ~new_P2_U3904 | ~new_P2_R693_U20;
  assign new_P2_R693_U110 = ~new_P2_U3896 | ~new_P2_R693_U21;
  assign new_P2_R693_U111 = ~new_P2_U3895 | ~new_P2_R693_U74;
  assign new_P2_R693_U112 = ~new_P2_U3529 | ~new_P2_R693_U73;
  assign new_P2_R693_U113 = ~new_P2_R693_U112 | ~new_P2_R693_U106;
  assign new_P2_R693_U114 = ~new_P2_R693_U72 | ~new_P2_R693_U108 | ~new_P2_U3535 | ~new_P2_R693_U6;
  assign new_P2_R693_U115 = ~new_P2_R693_U106 | ~new_P2_R693_U112 | ~new_P2_U3530;
  assign new_P2_R693_U116 = ~new_P2_R693_U75 | ~new_P2_R693_U108;
  assign new_P2_R693_U117 = ~new_P2_R693_U17 | ~new_P2_R693_U108 | ~new_P2_U3534 | ~new_P2_R693_U6;
  assign new_P2_R693_U118 = ~new_P2_U3543 | ~new_P2_R693_U32;
  assign new_P2_R693_U119 = ~new_P2_U3544 | ~new_P2_R693_U29;
  assign new_P2_R693_U120 = ~new_P2_U3901 | ~new_P2_R693_U67;
  assign new_P2_R693_U121 = ~new_P2_U3902 | ~new_P2_R693_U25;
  assign new_P2_R693_U122 = ~new_P2_R693_U79 | ~new_P2_R693_U118;
  assign new_P2_R693_U123 = ~new_P2_R693_U80 | ~new_P2_R693_U7;
  assign new_P2_R693_U124 = ~new_P2_U3445 | ~new_P2_R693_U28;
  assign new_P2_R693_U125 = ~new_P2_U3903 | ~new_P2_R693_U27;
  assign new_P2_R693_U126 = ~new_P2_U3437 | ~new_P2_R693_U35;
  assign new_P2_R693_U127 = ~new_P2_U3537 | ~new_P2_R693_U70;
  assign new_P2_R693_U128 = ~new_P2_U3536 | ~new_P2_R693_U71;
  assign new_P2_R693_U129 = ~new_P2_U3434 | ~new_P2_R693_U66;
  assign new_P2_R693_U130 = ~new_P2_U3419 | ~new_P2_R693_U59;
  assign new_P2_R693_U131 = ~new_P2_U3553 | ~new_P2_R693_U48;
  assign new_P2_R693_U132 = ~new_P2_U3416 | ~new_P2_R693_U58;
  assign new_P2_R693_U133 = ~new_P2_U3410 | ~new_P2_R693_U56;
  assign new_P2_R693_U134 = ~new_P2_U3413 | ~new_P2_R693_U57;
  assign new_P2_R693_U135 = ~new_P2_U3407 | ~new_P2_R693_U55;
  assign new_P2_R693_U136 = ~new_P2_U3404 | ~new_P2_R693_U54;
  assign new_P2_R693_U137 = ~new_P2_U3401 | ~new_P2_R693_U53;
  assign new_P2_R693_U138 = ~new_P2_U3398 | ~new_P2_R693_U52;
  assign new_P2_R693_U139 = ~new_P2_R693_U82 | ~new_P2_R693_U131;
  assign new_P2_R693_U140 = ~new_P2_U3395 | ~new_P2_R693_U51;
  assign new_P2_R693_U141 = ~new_P2_U3392 | ~new_P2_R693_U46;
  assign new_P2_R693_U142 = ~new_P2_R693_U85 | ~new_P2_R693_U12;
  assign new_P2_R693_U143 = ~new_P2_U3550 | ~new_P2_R693_U61;
  assign new_P2_R693_U144 = ~new_P2_U3549 | ~new_P2_R693_U64;
  assign new_P2_R693_U145 = ~new_P2_U3524 | ~new_P2_R693_U41;
  assign new_P2_R693_U146 = ~new_P2_U3523 | ~new_P2_R693_U39;
  assign new_P2_R693_U147 = ~new_P2_R693_U146 | ~new_P2_R693_U145;
  assign new_P2_R693_U148 = ~new_P2_U3528 | ~new_P2_R693_U44;
  assign new_P2_R693_U149 = ~new_P2_U3527 | ~new_P2_R693_U43;
  assign new_P2_R693_U150 = ~new_P2_R693_U149 | ~new_P2_R693_U148;
  assign new_P2_R693_U151 = ~new_P2_R693_U88 | ~new_P2_R693_U150;
  assign new_P2_R693_U152 = ~new_P2_U3526 | ~new_P2_R693_U42;
  assign new_P2_R693_U153 = ~new_P2_U3525 | ~new_P2_R693_U40;
  assign new_P2_R693_U154 = ~new_P2_R693_U89 | ~new_P2_R693_U151;
  assign new_P2_R693_U155 = ~new_P2_R693_U86 | ~new_P2_R693_U12;
  assign new_P2_R693_U156 = ~new_P2_R693_U87 | ~new_P2_R693_U11;
  assign new_P2_R693_U157 = ~new_P2_R693_U10 | ~new_P2_R693_U154;
  assign new_P2_R693_U158 = ~new_P2_R693_U90 | ~new_P2_R693_U147;
  assign new_P2_R693_U159 = ~new_P2_U3552 | ~new_P2_R693_U38;
  assign new_P2_R693_U160 = ~new_P2_U3551 | ~new_P2_R693_U62;
  assign new_P2_R693_U161 = ~new_P2_R693_U142 | ~new_P2_R693_U155 | ~new_P2_R693_U92 | ~new_P2_R693_U157 | ~new_P2_R693_U156;
  assign new_P2_R693_U162 = ~new_P2_U3549 | ~new_P2_R693_U64;
  assign new_P2_R693_U163 = ~new_P2_R693_U93 | ~new_P2_R693_U162;
  assign new_P2_R693_U164 = ~new_P2_R693_U94 | ~new_P2_R693_U13;
  assign new_P2_R693_U165 = ~new_P2_U3431 | ~new_P2_R693_U65;
  assign new_P2_R693_U166 = ~new_P2_U3428 | ~new_P2_R693_U50;
  assign new_P2_R693_U167 = ~new_P2_R693_U161 | ~new_P2_R693_U96;
  assign new_P2_R693_U168 = ~new_P2_U3548 | ~new_P2_R693_U63;
  assign new_P2_R693_U169 = ~new_P2_R693_U168 | ~new_P2_R693_U167;
  assign new_P2_R693_U170 = ~new_P2_R693_U169 | ~new_P2_R693_U129;
  assign new_P2_R693_U171 = ~new_P2_U3547 | ~new_P2_R693_U37;
  assign new_P2_R693_U172 = ~new_P2_R693_U171 | ~new_P2_R693_U170;
  assign new_P2_R693_U173 = ~new_P2_U3545 | ~new_P2_R693_U31;
  assign new_P2_R693_U174 = ~new_P2_U3546 | ~new_P2_R693_U36;
  assign new_P2_R693_U175 = ~new_P2_R693_U78 | ~new_P2_R693_U7;
  assign new_P2_R693_U176 = ~new_P2_R693_U76 | ~new_P2_R693_U120;
  assign new_P2_R693_U177 = ~new_P2_R693_U77 | ~new_P2_R693_U8;
  assign new_P2_R693_U178 = ~new_P2_R693_U9 | ~new_P2_R693_U175;
  assign new_P2_R693_U179 = ~new_P2_R693_U9 | ~new_P2_R693_U172 | ~new_P2_R693_U126;
  assign new_P2_R693_U180 = ~new_P2_U3539 | ~new_P2_R693_U24;
  assign new_P2_R693_U181 = ~new_P2_U3538 | ~new_P2_R693_U69;
  assign new_P2_R693_U182 = ~new_P2_R693_U98 | ~new_P2_R693_U99 | ~new_P2_R693_U179 | ~new_P2_R693_U178;
  assign new_P2_R693_U183 = ~new_P2_U3900 | ~new_P2_R693_U68;
  assign new_P2_R693_U184 = ~new_P2_U3899 | ~new_P2_R693_U22;
  assign new_P2_R693_U185 = ~new_P2_R693_U184 | ~new_P2_R693_U183;
  assign new_P2_R693_U186 = ~new_P2_R693_U128 | ~new_P2_R693_U185 | ~new_P2_R693_U127;
  assign new_P2_R693_U187 = ~new_P2_U3898 | ~new_P2_R693_U23;
  assign new_P2_R693_U188 = ~new_P2_U3897 | ~new_P2_R693_U19;
  assign new_P2_R693_U189 = ~new_P2_R693_U101 | ~new_P2_R693_U108 | ~new_P2_R693_U182 | ~new_P2_R693_U186;
  assign new_P2_R693_U190 = ~new_P2_U3868 | ~new_P2_R693_U15;
  assign new_P2_R693_U191 = ~new_P2_U3904 | ~new_P2_R693_U20;
  assign new_P2_R693_U192 = ~new_P2_R693_U108 | ~new_P2_R693_U102;
  assign new_P2_R693_U193 = ~new_P2_U3530 | ~new_P2_R693_U112;
  assign new_P2_SUB_605_U6 = ~new_P2_SUB_605_U39 | ~new_P2_SUB_605_U100;
  assign new_P2_SUB_605_U7 = ~new_P2_SUB_605_U81 | ~new_P2_SUB_605_U107;
  assign new_P2_SUB_605_U8 = ~new_P2_SUB_605_U65 | ~new_P2_SUB_605_U72;
  assign new_P2_SUB_605_U9 = ~new_P2_SUB_605_U34 | ~new_P2_SUB_605_U112;
  assign new_P2_SUB_605_U10 = ~new_P2_SUB_605_U89 | ~new_P2_SUB_605_U99;
  assign new_P2_SUB_605_U11 = ~new_P2_SUB_605_U83 | ~new_P2_SUB_605_U105;
  assign new_P2_SUB_605_U12 = ~new_P2_SUB_605_U67 | ~new_P2_SUB_605_U70;
  assign new_P2_SUB_605_U13 = ~new_P2_SUB_605_U75 | ~new_P2_SUB_605_U113;
  assign new_P2_SUB_605_U14 = ~new_P2_SUB_605_U68 | ~new_P2_SUB_605_U69;
  assign new_P2_SUB_605_U15 = ~new_P2_SUB_605_U37 | ~new_P2_SUB_605_U104;
  assign new_P2_SUB_605_U16 = ~new_P2_SUB_605_U40 | ~new_P2_SUB_605_U98;
  assign new_P2_SUB_605_U17 = ~new_P2_SUB_605_U87 | ~new_P2_SUB_605_U101;
  assign new_P2_SUB_605_U18 = ~new_P2_SUB_605_U32 | ~new_P2_SUB_605_U71;
  assign new_P2_SUB_605_U19 = ~new_P2_SUB_605_U36 | ~new_P2_SUB_605_U106;
  assign new_P2_SUB_605_U20 = ~new_P2_SUB_605_U85 | ~new_P2_SUB_605_U103;
  assign new_P2_SUB_605_U21 = ~new_P2_SUB_605_U35 | ~new_P2_SUB_605_U108;
  assign new_P2_SUB_605_U22 = ~new_P2_SUB_605_U64 | ~new_P2_SUB_605_U73;
  assign new_P2_SUB_605_U23 = ~new_P2_SUB_605_U41 | ~new_P2_SUB_605_U96;
  assign new_P2_SUB_605_U24 = ~new_P2_SUB_605_U77 | ~new_P2_SUB_605_U111;
  assign new_P2_SUB_605_U25 = ~new_P2_SUB_605_U49 | ~new_P2_SUB_605_U110;
  assign new_P2_SUB_605_U26 = ~P2_REG3_REG_3_;
  assign new_P2_SUB_605_U27 = ~new_P2_SUB_605_U91 | ~new_P2_SUB_605_U97;
  assign new_P2_SUB_605_U28 = ~new_P2_SUB_605_U38 | ~new_P2_SUB_605_U102;
  assign new_P2_SUB_605_U29 = ~new_P2_SUB_605_U93 | ~new_P2_SUB_605_U95;
  assign new_P2_SUB_605_U30 = ~new_P2_SUB_605_U63 | ~new_P2_SUB_605_U74;
  assign new_P2_SUB_605_U31 = ~new_P2_SUB_605_U79 | ~new_P2_SUB_605_U109;
  assign new_P2_SUB_605_U32 = P2_REG3_REG_7_ | P2_REG3_REG_6_ | P2_REG3_REG_5_ | P2_REG3_REG_4_ | P2_REG3_REG_3_;
  assign new_P2_SUB_605_U33 = ~P2_REG3_REG_8_;
  assign new_P2_SUB_605_U34 = ~new_P2_SUB_605_U53 | ~new_P2_SUB_605_U66;
  assign new_P2_SUB_605_U35 = ~new_P2_SUB_605_U54 | ~new_P2_SUB_605_U76;
  assign new_P2_SUB_605_U36 = ~new_P2_SUB_605_U55 | ~new_P2_SUB_605_U80;
  assign new_P2_SUB_605_U37 = ~new_P2_SUB_605_U56 | ~new_P2_SUB_605_U82;
  assign new_P2_SUB_605_U38 = ~new_P2_SUB_605_U57 | ~new_P2_SUB_605_U84;
  assign new_P2_SUB_605_U39 = ~new_P2_SUB_605_U58 | ~new_P2_SUB_605_U86;
  assign new_P2_SUB_605_U40 = ~new_P2_SUB_605_U59 | ~new_P2_SUB_605_U88;
  assign new_P2_SUB_605_U41 = ~new_P2_SUB_605_U60 | ~new_P2_SUB_605_U90;
  assign new_P2_SUB_605_U42 = ~P2_REG3_REG_28_;
  assign new_P2_SUB_605_U43 = ~P2_REG3_REG_26_;
  assign new_P2_SUB_605_U44 = ~P2_REG3_REG_24_;
  assign new_P2_SUB_605_U45 = ~P2_REG3_REG_22_;
  assign new_P2_SUB_605_U46 = ~P2_REG3_REG_20_;
  assign new_P2_SUB_605_U47 = ~P2_REG3_REG_18_;
  assign new_P2_SUB_605_U48 = ~P2_REG3_REG_16_;
  assign new_P2_SUB_605_U49 = ~new_P2_SUB_605_U61 | ~new_P2_SUB_605_U76;
  assign new_P2_SUB_605_U50 = ~P2_REG3_REG_14_;
  assign new_P2_SUB_605_U51 = ~P2_REG3_REG_12_;
  assign new_P2_SUB_605_U52 = ~P2_REG3_REG_8_ & ~P2_REG3_REG_9_;
  assign new_P2_SUB_605_U53 = ~P2_REG3_REG_9_ & ~P2_REG3_REG_8_ & ~P2_REG3_REG_10_ & ~P2_REG3_REG_11_;
  assign new_P2_SUB_605_U54 = ~P2_REG3_REG_15_ & ~P2_REG3_REG_14_ & ~P2_REG3_REG_12_ & ~P2_REG3_REG_13_;
  assign new_P2_SUB_605_U55 = ~P2_REG3_REG_16_ & ~P2_REG3_REG_17_;
  assign new_P2_SUB_605_U56 = ~P2_REG3_REG_18_ & ~P2_REG3_REG_19_;
  assign new_P2_SUB_605_U57 = ~P2_REG3_REG_20_ & ~P2_REG3_REG_21_;
  assign new_P2_SUB_605_U58 = ~P2_REG3_REG_22_ & ~P2_REG3_REG_23_;
  assign new_P2_SUB_605_U59 = ~P2_REG3_REG_24_ & ~P2_REG3_REG_25_;
  assign new_P2_SUB_605_U60 = ~P2_REG3_REG_26_ & ~P2_REG3_REG_27_;
  assign new_P2_SUB_605_U61 = ~P2_REG3_REG_12_ & ~P2_REG3_REG_13_;
  assign new_P2_SUB_605_U62 = ~P2_REG3_REG_8_ & ~P2_REG3_REG_9_ & ~P2_REG3_REG_10_;
  assign new_P2_SUB_605_U63 = P2_REG3_REG_3_ | P2_REG3_REG_4_;
  assign new_P2_SUB_605_U64 = P2_REG3_REG_5_ | P2_REG3_REG_4_ | P2_REG3_REG_3_;
  assign new_P2_SUB_605_U65 = P2_REG3_REG_3_ | P2_REG3_REG_4_ | P2_REG3_REG_5_ | P2_REG3_REG_6_;
  assign new_P2_SUB_605_U66 = ~new_P2_SUB_605_U32;
  assign new_P2_SUB_605_U67 = ~new_P2_SUB_605_U66 | ~new_P2_SUB_605_U33;
  assign new_P2_SUB_605_U68 = ~new_P2_SUB_605_U52 | ~new_P2_SUB_605_U66;
  assign new_P2_SUB_605_U69 = ~P2_REG3_REG_9_ | ~new_P2_SUB_605_U67;
  assign new_P2_SUB_605_U70 = ~P2_REG3_REG_8_ | ~new_P2_SUB_605_U32;
  assign new_P2_SUB_605_U71 = ~P2_REG3_REG_7_ | ~new_P2_SUB_605_U65;
  assign new_P2_SUB_605_U72 = ~P2_REG3_REG_6_ | ~new_P2_SUB_605_U64;
  assign new_P2_SUB_605_U73 = ~P2_REG3_REG_5_ | ~new_P2_SUB_605_U63;
  assign new_P2_SUB_605_U74 = ~P2_REG3_REG_4_ | ~P2_REG3_REG_3_;
  assign new_P2_SUB_605_U75 = ~new_P2_SUB_605_U62 | ~new_P2_SUB_605_U66;
  assign new_P2_SUB_605_U76 = ~new_P2_SUB_605_U34;
  assign new_P2_SUB_605_U77 = ~new_P2_SUB_605_U76 | ~new_P2_SUB_605_U51;
  assign new_P2_SUB_605_U78 = ~new_P2_SUB_605_U49;
  assign new_P2_SUB_605_U79 = ~new_P2_SUB_605_U78 | ~new_P2_SUB_605_U50;
  assign new_P2_SUB_605_U80 = ~new_P2_SUB_605_U35;
  assign new_P2_SUB_605_U81 = ~new_P2_SUB_605_U80 | ~new_P2_SUB_605_U48;
  assign new_P2_SUB_605_U82 = ~new_P2_SUB_605_U36;
  assign new_P2_SUB_605_U83 = ~new_P2_SUB_605_U82 | ~new_P2_SUB_605_U47;
  assign new_P2_SUB_605_U84 = ~new_P2_SUB_605_U37;
  assign new_P2_SUB_605_U85 = ~new_P2_SUB_605_U84 | ~new_P2_SUB_605_U46;
  assign new_P2_SUB_605_U86 = ~new_P2_SUB_605_U38;
  assign new_P2_SUB_605_U87 = ~new_P2_SUB_605_U86 | ~new_P2_SUB_605_U45;
  assign new_P2_SUB_605_U88 = ~new_P2_SUB_605_U39;
  assign new_P2_SUB_605_U89 = ~new_P2_SUB_605_U88 | ~new_P2_SUB_605_U44;
  assign new_P2_SUB_605_U90 = ~new_P2_SUB_605_U40;
  assign new_P2_SUB_605_U91 = ~new_P2_SUB_605_U90 | ~new_P2_SUB_605_U43;
  assign new_P2_SUB_605_U92 = ~new_P2_SUB_605_U41;
  assign new_P2_SUB_605_U93 = ~new_P2_SUB_605_U92 | ~new_P2_SUB_605_U42;
  assign new_P2_SUB_605_U94 = ~new_P2_SUB_605_U93;
  assign new_P2_SUB_605_U95 = ~P2_REG3_REG_28_ | ~new_P2_SUB_605_U41;
  assign new_P2_SUB_605_U96 = ~P2_REG3_REG_27_ | ~new_P2_SUB_605_U91;
  assign new_P2_SUB_605_U97 = ~P2_REG3_REG_26_ | ~new_P2_SUB_605_U40;
  assign new_P2_SUB_605_U98 = ~P2_REG3_REG_25_ | ~new_P2_SUB_605_U89;
  assign new_P2_SUB_605_U99 = ~P2_REG3_REG_24_ | ~new_P2_SUB_605_U39;
  assign new_P2_SUB_605_U100 = ~P2_REG3_REG_23_ | ~new_P2_SUB_605_U87;
  assign new_P2_SUB_605_U101 = ~P2_REG3_REG_22_ | ~new_P2_SUB_605_U38;
  assign new_P2_SUB_605_U102 = ~P2_REG3_REG_21_ | ~new_P2_SUB_605_U85;
  assign new_P2_SUB_605_U103 = ~P2_REG3_REG_20_ | ~new_P2_SUB_605_U37;
  assign new_P2_SUB_605_U104 = ~P2_REG3_REG_19_ | ~new_P2_SUB_605_U83;
  assign new_P2_SUB_605_U105 = ~P2_REG3_REG_18_ | ~new_P2_SUB_605_U36;
  assign new_P2_SUB_605_U106 = ~P2_REG3_REG_17_ | ~new_P2_SUB_605_U81;
  assign new_P2_SUB_605_U107 = ~P2_REG3_REG_16_ | ~new_P2_SUB_605_U35;
  assign new_P2_SUB_605_U108 = ~P2_REG3_REG_15_ | ~new_P2_SUB_605_U79;
  assign new_P2_SUB_605_U109 = ~P2_REG3_REG_14_ | ~new_P2_SUB_605_U49;
  assign new_P2_SUB_605_U110 = ~P2_REG3_REG_13_ | ~new_P2_SUB_605_U77;
  assign new_P2_SUB_605_U111 = ~P2_REG3_REG_12_ | ~new_P2_SUB_605_U34;
  assign new_P2_SUB_605_U112 = ~P2_REG3_REG_11_ | ~new_P2_SUB_605_U75;
  assign new_P2_SUB_605_U113 = ~P2_REG3_REG_10_ | ~new_P2_SUB_605_U68;
  assign new_P2_R1095_U6 = new_P2_R1095_U212 & new_P2_R1095_U211;
  assign new_P2_R1095_U7 = new_P2_R1095_U246 & new_P2_R1095_U245;
  assign new_P2_R1095_U8 = new_P2_R1095_U193 & new_P2_R1095_U257;
  assign new_P2_R1095_U9 = new_P2_R1095_U259 & new_P2_R1095_U258;
  assign new_P2_R1095_U10 = new_P2_R1095_U194 & new_P2_R1095_U281;
  assign new_P2_R1095_U11 = new_P2_R1095_U283 & new_P2_R1095_U282;
  assign new_P2_R1095_U12 = new_P2_R1095_U299 & new_P2_R1095_U195;
  assign new_P2_R1095_U13 = new_P2_R1095_U215 & new_P2_R1095_U210 & new_P2_R1095_U197;
  assign new_P2_R1095_U14 = new_P2_R1095_U220 & new_P2_R1095_U198;
  assign new_P2_R1095_U15 = new_P2_R1095_U244 & new_P2_R1095_U224 & new_P2_R1095_U192;
  assign new_P2_R1095_U16 = new_P2_R1095_U399 & new_P2_R1095_U398;
  assign new_P2_R1095_U17 = ~new_P2_R1095_U331 | ~new_P2_R1095_U334;
  assign new_P2_R1095_U18 = ~new_P2_R1095_U322 | ~new_P2_R1095_U325;
  assign new_P2_R1095_U19 = ~new_P2_R1095_U311 | ~new_P2_R1095_U314;
  assign new_P2_R1095_U20 = ~new_P2_R1095_U305 | ~new_P2_R1095_U357;
  assign new_P2_R1095_U21 = ~new_P2_R1095_U137 | ~new_P2_R1095_U186;
  assign new_P2_R1095_U22 = ~new_P2_R1095_U242 | ~new_P2_R1095_U347;
  assign new_P2_R1095_U23 = ~new_P2_R1095_U235 | ~new_P2_R1095_U238;
  assign new_P2_R1095_U24 = ~new_P2_R1095_U227 | ~new_P2_R1095_U229;
  assign new_P2_R1095_U25 = ~new_P2_R1095_U175 | ~new_P2_R1095_U337;
  assign new_P2_R1095_U26 = ~new_P2_U3069;
  assign new_P2_R1095_U27 = ~new_P2_U3069 | ~new_P2_R1095_U32;
  assign new_P2_R1095_U28 = ~new_P2_U3083;
  assign new_P2_R1095_U29 = ~new_P2_U3404;
  assign new_P2_R1095_U30 = ~new_P2_U3407;
  assign new_P2_R1095_U31 = ~new_P2_U3401;
  assign new_P2_R1095_U32 = ~new_P2_U3410;
  assign new_P2_R1095_U33 = ~new_P2_U3413;
  assign new_P2_R1095_U34 = ~new_P2_U3067;
  assign new_P2_R1095_U35 = ~new_P2_U3067 | ~new_P2_R1095_U37;
  assign new_P2_R1095_U36 = ~new_P2_U3063;
  assign new_P2_R1095_U37 = ~new_P2_U3395;
  assign new_P2_R1095_U38 = ~new_P2_U3387;
  assign new_P2_R1095_U39 = ~new_P2_U3077;
  assign new_P2_R1095_U40 = ~new_P2_U3398;
  assign new_P2_R1095_U41 = ~new_P2_U3070;
  assign new_P2_R1095_U42 = ~new_P2_U3066;
  assign new_P2_R1095_U43 = ~new_P2_U3059;
  assign new_P2_R1095_U44 = ~new_P2_U3059 | ~new_P2_R1095_U31;
  assign new_P2_R1095_U45 = ~new_P2_R1095_U216 | ~new_P2_R1095_U214;
  assign new_P2_R1095_U46 = ~new_P2_U3416;
  assign new_P2_R1095_U47 = ~new_P2_U3082;
  assign new_P2_R1095_U48 = ~new_P2_R1095_U45 | ~new_P2_R1095_U217;
  assign new_P2_R1095_U49 = ~new_P2_R1095_U44 | ~new_P2_R1095_U231;
  assign new_P2_R1095_U50 = ~new_P2_R1095_U338 | ~new_P2_R1095_U204 | ~new_P2_R1095_U188;
  assign new_P2_R1095_U51 = ~new_P2_U3895;
  assign new_P2_R1095_U52 = ~new_P2_U3056;
  assign new_P2_R1095_U53 = ~new_P2_U3056 | ~new_P2_R1095_U90;
  assign new_P2_R1095_U54 = ~new_P2_U3052;
  assign new_P2_R1095_U55 = ~new_P2_U3071;
  assign new_P2_R1095_U56 = ~new_P2_U3062;
  assign new_P2_R1095_U57 = ~new_P2_U3061;
  assign new_P2_R1095_U58 = ~new_P2_U3419;
  assign new_P2_R1095_U59 = ~new_P2_U3082 | ~new_P2_R1095_U46;
  assign new_P2_R1095_U60 = ~new_P2_U3422;
  assign new_P2_R1095_U61 = ~new_P2_U3425;
  assign new_P2_R1095_U62 = ~new_P2_R1095_U249 | ~new_P2_R1095_U248;
  assign new_P2_R1095_U63 = ~new_P2_U3428;
  assign new_P2_R1095_U64 = ~new_P2_U3079;
  assign new_P2_R1095_U65 = ~new_P2_U3437;
  assign new_P2_R1095_U66 = ~new_P2_U3434;
  assign new_P2_R1095_U67 = ~new_P2_U3431;
  assign new_P2_R1095_U68 = ~new_P2_U3072;
  assign new_P2_R1095_U69 = ~new_P2_U3073;
  assign new_P2_R1095_U70 = ~new_P2_U3078;
  assign new_P2_R1095_U71 = ~new_P2_U3078 | ~new_P2_R1095_U67;
  assign new_P2_R1095_U72 = ~new_P2_U3440;
  assign new_P2_R1095_U73 = ~new_P2_U3068;
  assign new_P2_R1095_U74 = ~new_P2_U3081;
  assign new_P2_R1095_U75 = ~new_P2_U3445;
  assign new_P2_R1095_U76 = ~new_P2_U3080;
  assign new_P2_R1095_U77 = ~new_P2_U3903;
  assign new_P2_R1095_U78 = ~new_P2_U3075;
  assign new_P2_R1095_U79 = ~new_P2_U3900;
  assign new_P2_R1095_U80 = ~new_P2_U3901;
  assign new_P2_R1095_U81 = ~new_P2_U3902;
  assign new_P2_R1095_U82 = ~new_P2_U3065;
  assign new_P2_R1095_U83 = ~new_P2_U3060;
  assign new_P2_R1095_U84 = ~new_P2_U3074;
  assign new_P2_R1095_U85 = ~new_P2_U3074 | ~new_P2_R1095_U81;
  assign new_P2_R1095_U86 = ~new_P2_U3899;
  assign new_P2_R1095_U87 = ~new_P2_U3064;
  assign new_P2_R1095_U88 = ~new_P2_U3898;
  assign new_P2_R1095_U89 = ~new_P2_U3057;
  assign new_P2_R1095_U90 = ~new_P2_U3897;
  assign new_P2_R1095_U91 = ~new_P2_U3896;
  assign new_P2_R1095_U92 = ~new_P2_U3053;
  assign new_P2_R1095_U93 = ~new_P2_R1095_U297 | ~new_P2_R1095_U296;
  assign new_P2_R1095_U94 = ~new_P2_R1095_U85 | ~new_P2_R1095_U307;
  assign new_P2_R1095_U95 = ~new_P2_R1095_U71 | ~new_P2_R1095_U318;
  assign new_P2_R1095_U96 = ~new_P2_R1095_U349 | ~new_P2_R1095_U59;
  assign new_P2_R1095_U97 = ~new_P2_U3076;
  assign new_P2_R1095_U98 = ~new_P2_R1095_U406 | ~new_P2_R1095_U405;
  assign new_P2_R1095_U99 = ~new_P2_R1095_U420 | ~new_P2_R1095_U419;
  assign new_P2_R1095_U100 = ~new_P2_R1095_U425 | ~new_P2_R1095_U424;
  assign new_P2_R1095_U101 = ~new_P2_R1095_U441 | ~new_P2_R1095_U440;
  assign new_P2_R1095_U102 = ~new_P2_R1095_U446 | ~new_P2_R1095_U445;
  assign new_P2_R1095_U103 = ~new_P2_R1095_U451 | ~new_P2_R1095_U450;
  assign new_P2_R1095_U104 = ~new_P2_R1095_U456 | ~new_P2_R1095_U455;
  assign new_P2_R1095_U105 = ~new_P2_R1095_U461 | ~new_P2_R1095_U460;
  assign new_P2_R1095_U106 = ~new_P2_R1095_U477 | ~new_P2_R1095_U476;
  assign new_P2_R1095_U107 = ~new_P2_R1095_U482 | ~new_P2_R1095_U481;
  assign new_P2_R1095_U108 = ~new_P2_R1095_U365 | ~new_P2_R1095_U364;
  assign new_P2_R1095_U109 = ~new_P2_R1095_U374 | ~new_P2_R1095_U373;
  assign new_P2_R1095_U110 = ~new_P2_R1095_U381 | ~new_P2_R1095_U380;
  assign new_P2_R1095_U111 = ~new_P2_R1095_U385 | ~new_P2_R1095_U384;
  assign new_P2_R1095_U112 = ~new_P2_R1095_U394 | ~new_P2_R1095_U393;
  assign new_P2_R1095_U113 = ~new_P2_R1095_U415 | ~new_P2_R1095_U414;
  assign new_P2_R1095_U114 = ~new_P2_R1095_U432 | ~new_P2_R1095_U431;
  assign new_P2_R1095_U115 = ~new_P2_R1095_U436 | ~new_P2_R1095_U435;
  assign new_P2_R1095_U116 = ~new_P2_R1095_U468 | ~new_P2_R1095_U467;
  assign new_P2_R1095_U117 = ~new_P2_R1095_U472 | ~new_P2_R1095_U471;
  assign new_P2_R1095_U118 = ~new_P2_R1095_U489 | ~new_P2_R1095_U488;
  assign new_P2_R1095_U119 = new_P2_R1095_U206 & new_P2_R1095_U196;
  assign new_P2_R1095_U120 = new_P2_R1095_U209 & new_P2_R1095_U208;
  assign new_P2_R1095_U121 = new_P2_R1095_U14 & new_P2_R1095_U13;
  assign new_P2_R1095_U122 = new_P2_R1095_U340 & new_P2_R1095_U222;
  assign new_P2_R1095_U123 = new_P2_R1095_U342 & new_P2_R1095_U122;
  assign new_P2_R1095_U124 = new_P2_R1095_U27 & new_P2_R1095_U367 & new_P2_R1095_U366;
  assign new_P2_R1095_U125 = new_P2_R1095_U370 & new_P2_R1095_U198;
  assign new_P2_R1095_U126 = new_P2_R1095_U237 & new_P2_R1095_U6;
  assign new_P2_R1095_U127 = new_P2_R1095_U377 & new_P2_R1095_U197;
  assign new_P2_R1095_U128 = new_P2_R1095_U35 & new_P2_R1095_U387 & new_P2_R1095_U386;
  assign new_P2_R1095_U129 = new_P2_R1095_U390 & new_P2_R1095_U196;
  assign new_P2_R1095_U130 = new_P2_R1095_U251 & new_P2_R1095_U15;
  assign new_P2_R1095_U131 = new_P2_R1095_U343 & new_P2_R1095_U252;
  assign new_P2_R1095_U132 = new_P2_R1095_U262 & new_P2_R1095_U8;
  assign new_P2_R1095_U133 = new_P2_R1095_U286 & new_P2_R1095_U10;
  assign new_P2_R1095_U134 = new_P2_R1095_U302 & new_P2_R1095_U301;
  assign new_P2_R1095_U135 = new_P2_R1095_U397 & new_P2_R1095_U303;
  assign new_P2_R1095_U136 = new_P2_R1095_U16 & new_P2_R1095_U304 & new_P2_R1095_U302 & new_P2_R1095_U301;
  assign new_P2_R1095_U137 = new_P2_R1095_U359 & new_P2_R1095_U165;
  assign new_P2_R1095_U138 = ~new_P2_R1095_U403 | ~new_P2_R1095_U402;
  assign new_P2_R1095_U139 = new_P2_R1095_U53 & new_P2_R1095_U408 & new_P2_R1095_U407;
  assign new_P2_R1095_U140 = new_P2_R1095_U411 & new_P2_R1095_U195;
  assign new_P2_R1095_U141 = ~new_P2_R1095_U417 | ~new_P2_R1095_U416;
  assign new_P2_R1095_U142 = ~new_P2_R1095_U422 | ~new_P2_R1095_U421;
  assign new_P2_R1095_U143 = new_P2_R1095_U313 & new_P2_R1095_U11;
  assign new_P2_R1095_U144 = new_P2_R1095_U428 & new_P2_R1095_U194;
  assign new_P2_R1095_U145 = ~new_P2_R1095_U438 | ~new_P2_R1095_U437;
  assign new_P2_R1095_U146 = ~new_P2_R1095_U443 | ~new_P2_R1095_U442;
  assign new_P2_R1095_U147 = ~new_P2_R1095_U448 | ~new_P2_R1095_U447;
  assign new_P2_R1095_U148 = ~new_P2_R1095_U453 | ~new_P2_R1095_U452;
  assign new_P2_R1095_U149 = ~new_P2_R1095_U458 | ~new_P2_R1095_U457;
  assign new_P2_R1095_U150 = new_P2_R1095_U324 & new_P2_R1095_U9;
  assign new_P2_R1095_U151 = new_P2_R1095_U464 & new_P2_R1095_U193;
  assign new_P2_R1095_U152 = ~new_P2_R1095_U474 | ~new_P2_R1095_U473;
  assign new_P2_R1095_U153 = ~new_P2_R1095_U479 | ~new_P2_R1095_U478;
  assign new_P2_R1095_U154 = new_P2_R1095_U333 & new_P2_R1095_U7;
  assign new_P2_R1095_U155 = new_P2_R1095_U485 & new_P2_R1095_U192;
  assign new_P2_R1095_U156 = new_P2_R1095_U363 & new_P2_R1095_U362;
  assign new_P2_R1095_U157 = ~new_P2_R1095_U123 | ~new_P2_R1095_U341;
  assign new_P2_R1095_U158 = new_P2_R1095_U372 & new_P2_R1095_U371;
  assign new_P2_R1095_U159 = new_P2_R1095_U379 & new_P2_R1095_U378;
  assign new_P2_R1095_U160 = new_P2_R1095_U383 & new_P2_R1095_U382;
  assign new_P2_R1095_U161 = ~new_P2_R1095_U120 | ~new_P2_R1095_U344;
  assign new_P2_R1095_U162 = new_P2_R1095_U392 & new_P2_R1095_U391;
  assign new_P2_R1095_U163 = ~new_P2_U3904;
  assign new_P2_R1095_U164 = ~new_P2_U3054;
  assign new_P2_R1095_U165 = new_P2_R1095_U401 & new_P2_R1095_U400;
  assign new_P2_R1095_U166 = ~new_P2_R1095_U134 | ~new_P2_R1095_U360;
  assign new_P2_R1095_U167 = new_P2_R1095_U413 & new_P2_R1095_U412;
  assign new_P2_R1095_U168 = ~new_P2_R1095_U293 | ~new_P2_R1095_U292;
  assign new_P2_R1095_U169 = ~new_P2_R1095_U289 | ~new_P2_R1095_U288;
  assign new_P2_R1095_U170 = new_P2_R1095_U430 & new_P2_R1095_U429;
  assign new_P2_R1095_U171 = new_P2_R1095_U434 & new_P2_R1095_U433;
  assign new_P2_R1095_U172 = ~new_P2_R1095_U279 | ~new_P2_R1095_U278;
  assign new_P2_R1095_U173 = ~new_P2_R1095_U275 | ~new_P2_R1095_U274;
  assign new_P2_R1095_U174 = ~new_P2_U3392;
  assign new_P2_R1095_U175 = ~new_P2_U3387 | ~new_P2_R1095_U97;
  assign new_P2_R1095_U176 = ~new_P2_R1095_U339 | ~new_P2_R1095_U271 | ~new_P2_R1095_U187;
  assign new_P2_R1095_U177 = ~new_P2_U3443;
  assign new_P2_R1095_U178 = ~new_P2_R1095_U269 | ~new_P2_R1095_U268;
  assign new_P2_R1095_U179 = ~new_P2_R1095_U265 | ~new_P2_R1095_U264;
  assign new_P2_R1095_U180 = new_P2_R1095_U466 & new_P2_R1095_U465;
  assign new_P2_R1095_U181 = new_P2_R1095_U470 & new_P2_R1095_U469;
  assign new_P2_R1095_U182 = ~new_P2_R1095_U255 | ~new_P2_R1095_U254;
  assign new_P2_R1095_U183 = ~new_P2_R1095_U131 | ~new_P2_R1095_U353;
  assign new_P2_R1095_U184 = ~new_P2_R1095_U351 | ~new_P2_R1095_U62;
  assign new_P2_R1095_U185 = new_P2_R1095_U487 & new_P2_R1095_U486;
  assign new_P2_R1095_U186 = ~new_P2_R1095_U135 | ~new_P2_R1095_U166;
  assign new_P2_R1095_U187 = ~new_P2_R1095_U178 | ~new_P2_R1095_U177;
  assign new_P2_R1095_U188 = ~new_P2_R1095_U175 | ~new_P2_R1095_U174;
  assign new_P2_R1095_U189 = ~new_P2_R1095_U53;
  assign new_P2_R1095_U190 = ~new_P2_R1095_U35;
  assign new_P2_R1095_U191 = ~new_P2_R1095_U27;
  assign new_P2_R1095_U192 = ~new_P2_U3419 | ~new_P2_R1095_U57;
  assign new_P2_R1095_U193 = ~new_P2_U3434 | ~new_P2_R1095_U69;
  assign new_P2_R1095_U194 = ~new_P2_U3901 | ~new_P2_R1095_U83;
  assign new_P2_R1095_U195 = ~new_P2_U3897 | ~new_P2_R1095_U52;
  assign new_P2_R1095_U196 = ~new_P2_U3395 | ~new_P2_R1095_U34;
  assign new_P2_R1095_U197 = ~new_P2_U3404 | ~new_P2_R1095_U42;
  assign new_P2_R1095_U198 = ~new_P2_U3410 | ~new_P2_R1095_U26;
  assign new_P2_R1095_U199 = ~new_P2_R1095_U71;
  assign new_P2_R1095_U200 = ~new_P2_R1095_U85;
  assign new_P2_R1095_U201 = ~new_P2_R1095_U44;
  assign new_P2_R1095_U202 = ~new_P2_R1095_U59;
  assign new_P2_R1095_U203 = ~new_P2_R1095_U175;
  assign new_P2_R1095_U204 = ~new_P2_U3077 | ~new_P2_R1095_U175;
  assign new_P2_R1095_U205 = ~new_P2_R1095_U50;
  assign new_P2_R1095_U206 = ~new_P2_U3398 | ~new_P2_R1095_U36;
  assign new_P2_R1095_U207 = ~new_P2_R1095_U36 | ~new_P2_R1095_U35;
  assign new_P2_R1095_U208 = ~new_P2_R1095_U207 | ~new_P2_R1095_U40;
  assign new_P2_R1095_U209 = ~new_P2_U3063 | ~new_P2_R1095_U190;
  assign new_P2_R1095_U210 = ~new_P2_U3407 | ~new_P2_R1095_U41;
  assign new_P2_R1095_U211 = ~new_P2_U3070 | ~new_P2_R1095_U30;
  assign new_P2_R1095_U212 = ~new_P2_U3066 | ~new_P2_R1095_U29;
  assign new_P2_R1095_U213 = ~new_P2_R1095_U201 | ~new_P2_R1095_U197;
  assign new_P2_R1095_U214 = ~new_P2_R1095_U6 | ~new_P2_R1095_U213;
  assign new_P2_R1095_U215 = ~new_P2_U3401 | ~new_P2_R1095_U43;
  assign new_P2_R1095_U216 = ~new_P2_U3407 | ~new_P2_R1095_U41;
  assign new_P2_R1095_U217 = ~new_P2_R1095_U13 | ~new_P2_R1095_U161;
  assign new_P2_R1095_U218 = ~new_P2_R1095_U45;
  assign new_P2_R1095_U219 = ~new_P2_R1095_U48;
  assign new_P2_R1095_U220 = ~new_P2_U3413 | ~new_P2_R1095_U28;
  assign new_P2_R1095_U221 = ~new_P2_R1095_U28 | ~new_P2_R1095_U27;
  assign new_P2_R1095_U222 = ~new_P2_U3083 | ~new_P2_R1095_U191;
  assign new_P2_R1095_U223 = ~new_P2_R1095_U157;
  assign new_P2_R1095_U224 = ~new_P2_U3416 | ~new_P2_R1095_U47;
  assign new_P2_R1095_U225 = ~new_P2_R1095_U224 | ~new_P2_R1095_U59;
  assign new_P2_R1095_U226 = ~new_P2_R1095_U219 | ~new_P2_R1095_U27;
  assign new_P2_R1095_U227 = ~new_P2_R1095_U125 | ~new_P2_R1095_U226;
  assign new_P2_R1095_U228 = ~new_P2_R1095_U48 | ~new_P2_R1095_U198;
  assign new_P2_R1095_U229 = ~new_P2_R1095_U124 | ~new_P2_R1095_U228;
  assign new_P2_R1095_U230 = ~new_P2_R1095_U27 | ~new_P2_R1095_U198;
  assign new_P2_R1095_U231 = ~new_P2_R1095_U215 | ~new_P2_R1095_U161;
  assign new_P2_R1095_U232 = ~new_P2_R1095_U49;
  assign new_P2_R1095_U233 = ~new_P2_U3066 | ~new_P2_R1095_U29;
  assign new_P2_R1095_U234 = ~new_P2_R1095_U232 | ~new_P2_R1095_U233;
  assign new_P2_R1095_U235 = ~new_P2_R1095_U127 | ~new_P2_R1095_U234;
  assign new_P2_R1095_U236 = ~new_P2_R1095_U49 | ~new_P2_R1095_U197;
  assign new_P2_R1095_U237 = ~new_P2_U3407 | ~new_P2_R1095_U41;
  assign new_P2_R1095_U238 = ~new_P2_R1095_U126 | ~new_P2_R1095_U236;
  assign new_P2_R1095_U239 = ~new_P2_U3066 | ~new_P2_R1095_U29;
  assign new_P2_R1095_U240 = ~new_P2_R1095_U239 | ~new_P2_R1095_U197;
  assign new_P2_R1095_U241 = ~new_P2_R1095_U215 | ~new_P2_R1095_U44;
  assign new_P2_R1095_U242 = ~new_P2_R1095_U129 | ~new_P2_R1095_U348;
  assign new_P2_R1095_U243 = ~new_P2_R1095_U35 | ~new_P2_R1095_U196;
  assign new_P2_R1095_U244 = ~new_P2_U3422 | ~new_P2_R1095_U56;
  assign new_P2_R1095_U245 = ~new_P2_U3062 | ~new_P2_R1095_U60;
  assign new_P2_R1095_U246 = ~new_P2_U3061 | ~new_P2_R1095_U58;
  assign new_P2_R1095_U247 = ~new_P2_R1095_U202 | ~new_P2_R1095_U192;
  assign new_P2_R1095_U248 = ~new_P2_R1095_U7 | ~new_P2_R1095_U247;
  assign new_P2_R1095_U249 = ~new_P2_U3422 | ~new_P2_R1095_U56;
  assign new_P2_R1095_U250 = ~new_P2_R1095_U62;
  assign new_P2_R1095_U251 = ~new_P2_U3425 | ~new_P2_R1095_U55;
  assign new_P2_R1095_U252 = ~new_P2_U3071 | ~new_P2_R1095_U61;
  assign new_P2_R1095_U253 = ~new_P2_U3428 | ~new_P2_R1095_U64;
  assign new_P2_R1095_U254 = ~new_P2_R1095_U253 | ~new_P2_R1095_U183;
  assign new_P2_R1095_U255 = ~new_P2_U3079 | ~new_P2_R1095_U63;
  assign new_P2_R1095_U256 = ~new_P2_R1095_U182;
  assign new_P2_R1095_U257 = ~new_P2_U3437 | ~new_P2_R1095_U68;
  assign new_P2_R1095_U258 = ~new_P2_U3072 | ~new_P2_R1095_U65;
  assign new_P2_R1095_U259 = ~new_P2_U3073 | ~new_P2_R1095_U66;
  assign new_P2_R1095_U260 = ~new_P2_R1095_U199 | ~new_P2_R1095_U8;
  assign new_P2_R1095_U261 = ~new_P2_R1095_U9 | ~new_P2_R1095_U260;
  assign new_P2_R1095_U262 = ~new_P2_U3431 | ~new_P2_R1095_U70;
  assign new_P2_R1095_U263 = ~new_P2_U3437 | ~new_P2_R1095_U68;
  assign new_P2_R1095_U264 = ~new_P2_R1095_U132 | ~new_P2_R1095_U182;
  assign new_P2_R1095_U265 = ~new_P2_R1095_U263 | ~new_P2_R1095_U261;
  assign new_P2_R1095_U266 = ~new_P2_R1095_U179;
  assign new_P2_R1095_U267 = ~new_P2_U3440 | ~new_P2_R1095_U73;
  assign new_P2_R1095_U268 = ~new_P2_R1095_U267 | ~new_P2_R1095_U179;
  assign new_P2_R1095_U269 = ~new_P2_U3068 | ~new_P2_R1095_U72;
  assign new_P2_R1095_U270 = ~new_P2_R1095_U178;
  assign new_P2_R1095_U271 = ~new_P2_U3081 | ~new_P2_R1095_U178;
  assign new_P2_R1095_U272 = ~new_P2_R1095_U176;
  assign new_P2_R1095_U273 = ~new_P2_U3445 | ~new_P2_R1095_U76;
  assign new_P2_R1095_U274 = ~new_P2_R1095_U273 | ~new_P2_R1095_U176;
  assign new_P2_R1095_U275 = ~new_P2_U3080 | ~new_P2_R1095_U75;
  assign new_P2_R1095_U276 = ~new_P2_R1095_U173;
  assign new_P2_R1095_U277 = ~new_P2_U3903 | ~new_P2_R1095_U78;
  assign new_P2_R1095_U278 = ~new_P2_R1095_U277 | ~new_P2_R1095_U173;
  assign new_P2_R1095_U279 = ~new_P2_U3075 | ~new_P2_R1095_U77;
  assign new_P2_R1095_U280 = ~new_P2_R1095_U172;
  assign new_P2_R1095_U281 = ~new_P2_U3900 | ~new_P2_R1095_U82;
  assign new_P2_R1095_U282 = ~new_P2_U3065 | ~new_P2_R1095_U79;
  assign new_P2_R1095_U283 = ~new_P2_U3060 | ~new_P2_R1095_U80;
  assign new_P2_R1095_U284 = ~new_P2_R1095_U200 | ~new_P2_R1095_U10;
  assign new_P2_R1095_U285 = ~new_P2_R1095_U11 | ~new_P2_R1095_U284;
  assign new_P2_R1095_U286 = ~new_P2_U3902 | ~new_P2_R1095_U84;
  assign new_P2_R1095_U287 = ~new_P2_U3900 | ~new_P2_R1095_U82;
  assign new_P2_R1095_U288 = ~new_P2_R1095_U133 | ~new_P2_R1095_U172;
  assign new_P2_R1095_U289 = ~new_P2_R1095_U287 | ~new_P2_R1095_U285;
  assign new_P2_R1095_U290 = ~new_P2_R1095_U169;
  assign new_P2_R1095_U291 = ~new_P2_U3899 | ~new_P2_R1095_U87;
  assign new_P2_R1095_U292 = ~new_P2_R1095_U291 | ~new_P2_R1095_U169;
  assign new_P2_R1095_U293 = ~new_P2_U3064 | ~new_P2_R1095_U86;
  assign new_P2_R1095_U294 = ~new_P2_R1095_U168;
  assign new_P2_R1095_U295 = ~new_P2_U3898 | ~new_P2_R1095_U89;
  assign new_P2_R1095_U296 = ~new_P2_R1095_U295 | ~new_P2_R1095_U168;
  assign new_P2_R1095_U297 = ~new_P2_U3057 | ~new_P2_R1095_U88;
  assign new_P2_R1095_U298 = ~new_P2_R1095_U93;
  assign new_P2_R1095_U299 = ~new_P2_U3896 | ~new_P2_R1095_U54;
  assign new_P2_R1095_U300 = ~new_P2_R1095_U54 | ~new_P2_R1095_U53;
  assign new_P2_R1095_U301 = ~new_P2_R1095_U300 | ~new_P2_R1095_U91;
  assign new_P2_R1095_U302 = ~new_P2_U3052 | ~new_P2_R1095_U189;
  assign new_P2_R1095_U303 = ~new_P2_U3895 | ~new_P2_R1095_U92;
  assign new_P2_R1095_U304 = ~new_P2_U3053 | ~new_P2_R1095_U51;
  assign new_P2_R1095_U305 = ~new_P2_R1095_U140 | ~new_P2_R1095_U355;
  assign new_P2_R1095_U306 = ~new_P2_R1095_U53 | ~new_P2_R1095_U195;
  assign new_P2_R1095_U307 = ~new_P2_R1095_U286 | ~new_P2_R1095_U172;
  assign new_P2_R1095_U308 = ~new_P2_R1095_U94;
  assign new_P2_R1095_U309 = ~new_P2_U3060 | ~new_P2_R1095_U80;
  assign new_P2_R1095_U310 = ~new_P2_R1095_U308 | ~new_P2_R1095_U309;
  assign new_P2_R1095_U311 = ~new_P2_R1095_U144 | ~new_P2_R1095_U310;
  assign new_P2_R1095_U312 = ~new_P2_R1095_U94 | ~new_P2_R1095_U194;
  assign new_P2_R1095_U313 = ~new_P2_U3900 | ~new_P2_R1095_U82;
  assign new_P2_R1095_U314 = ~new_P2_R1095_U143 | ~new_P2_R1095_U312;
  assign new_P2_R1095_U315 = ~new_P2_U3060 | ~new_P2_R1095_U80;
  assign new_P2_R1095_U316 = ~new_P2_R1095_U194 | ~new_P2_R1095_U315;
  assign new_P2_R1095_U317 = ~new_P2_R1095_U286 | ~new_P2_R1095_U85;
  assign new_P2_R1095_U318 = ~new_P2_R1095_U262 | ~new_P2_R1095_U182;
  assign new_P2_R1095_U319 = ~new_P2_R1095_U95;
  assign new_P2_R1095_U320 = ~new_P2_U3073 | ~new_P2_R1095_U66;
  assign new_P2_R1095_U321 = ~new_P2_R1095_U319 | ~new_P2_R1095_U320;
  assign new_P2_R1095_U322 = ~new_P2_R1095_U151 | ~new_P2_R1095_U321;
  assign new_P2_R1095_U323 = ~new_P2_R1095_U95 | ~new_P2_R1095_U193;
  assign new_P2_R1095_U324 = ~new_P2_U3437 | ~new_P2_R1095_U68;
  assign new_P2_R1095_U325 = ~new_P2_R1095_U150 | ~new_P2_R1095_U323;
  assign new_P2_R1095_U326 = ~new_P2_U3073 | ~new_P2_R1095_U66;
  assign new_P2_R1095_U327 = ~new_P2_R1095_U193 | ~new_P2_R1095_U326;
  assign new_P2_R1095_U328 = ~new_P2_R1095_U262 | ~new_P2_R1095_U71;
  assign new_P2_R1095_U329 = ~new_P2_U3061 | ~new_P2_R1095_U58;
  assign new_P2_R1095_U330 = ~new_P2_R1095_U350 | ~new_P2_R1095_U329;
  assign new_P2_R1095_U331 = ~new_P2_R1095_U155 | ~new_P2_R1095_U330;
  assign new_P2_R1095_U332 = ~new_P2_R1095_U96 | ~new_P2_R1095_U192;
  assign new_P2_R1095_U333 = ~new_P2_U3422 | ~new_P2_R1095_U56;
  assign new_P2_R1095_U334 = ~new_P2_R1095_U154 | ~new_P2_R1095_U332;
  assign new_P2_R1095_U335 = ~new_P2_U3061 | ~new_P2_R1095_U58;
  assign new_P2_R1095_U336 = ~new_P2_R1095_U192 | ~new_P2_R1095_U335;
  assign new_P2_R1095_U337 = ~new_P2_U3076 | ~new_P2_R1095_U38;
  assign new_P2_R1095_U338 = ~new_P2_U3077 | ~new_P2_R1095_U174;
  assign new_P2_R1095_U339 = ~new_P2_U3081 | ~new_P2_R1095_U177;
  assign new_P2_R1095_U340 = ~new_P2_R1095_U33 | ~new_P2_R1095_U221;
  assign new_P2_R1095_U341 = ~new_P2_R1095_U121 | ~new_P2_R1095_U161;
  assign new_P2_R1095_U342 = ~new_P2_R1095_U218 | ~new_P2_R1095_U14;
  assign new_P2_R1095_U343 = ~new_P2_R1095_U250 | ~new_P2_R1095_U251;
  assign new_P2_R1095_U344 = ~new_P2_R1095_U119 | ~new_P2_R1095_U50;
  assign new_P2_R1095_U345 = ~new_P2_R1095_U161;
  assign new_P2_R1095_U346 = ~new_P2_R1095_U196 | ~new_P2_R1095_U50;
  assign new_P2_R1095_U347 = ~new_P2_R1095_U128 | ~new_P2_R1095_U346;
  assign new_P2_R1095_U348 = ~new_P2_R1095_U205 | ~new_P2_R1095_U35;
  assign new_P2_R1095_U349 = ~new_P2_R1095_U224 | ~new_P2_R1095_U157;
  assign new_P2_R1095_U350 = ~new_P2_R1095_U96;
  assign new_P2_R1095_U351 = ~new_P2_R1095_U15 | ~new_P2_R1095_U157;
  assign new_P2_R1095_U352 = ~new_P2_R1095_U184;
  assign new_P2_R1095_U353 = ~new_P2_R1095_U130 | ~new_P2_R1095_U157;
  assign new_P2_R1095_U354 = ~new_P2_R1095_U183;
  assign new_P2_R1095_U355 = ~new_P2_R1095_U298 | ~new_P2_R1095_U53;
  assign new_P2_R1095_U356 = ~new_P2_R1095_U195 | ~new_P2_R1095_U93;
  assign new_P2_R1095_U357 = ~new_P2_R1095_U139 | ~new_P2_R1095_U356;
  assign new_P2_R1095_U358 = ~new_P2_R1095_U12 | ~new_P2_R1095_U93;
  assign new_P2_R1095_U359 = ~new_P2_R1095_U136 | ~new_P2_R1095_U358;
  assign new_P2_R1095_U360 = ~new_P2_R1095_U12 | ~new_P2_R1095_U93;
  assign new_P2_R1095_U361 = ~new_P2_R1095_U166;
  assign new_P2_R1095_U362 = ~new_P2_U3416 | ~new_P2_R1095_U47;
  assign new_P2_R1095_U363 = ~new_P2_U3082 | ~new_P2_R1095_U46;
  assign new_P2_R1095_U364 = ~new_P2_R1095_U225 | ~new_P2_R1095_U157;
  assign new_P2_R1095_U365 = ~new_P2_R1095_U223 | ~new_P2_R1095_U156;
  assign new_P2_R1095_U366 = ~new_P2_U3413 | ~new_P2_R1095_U28;
  assign new_P2_R1095_U367 = ~new_P2_U3083 | ~new_P2_R1095_U33;
  assign new_P2_R1095_U368 = ~new_P2_U3413 | ~new_P2_R1095_U28;
  assign new_P2_R1095_U369 = ~new_P2_U3083 | ~new_P2_R1095_U33;
  assign new_P2_R1095_U370 = ~new_P2_R1095_U369 | ~new_P2_R1095_U368;
  assign new_P2_R1095_U371 = ~new_P2_U3410 | ~new_P2_R1095_U26;
  assign new_P2_R1095_U372 = ~new_P2_U3069 | ~new_P2_R1095_U32;
  assign new_P2_R1095_U373 = ~new_P2_R1095_U230 | ~new_P2_R1095_U48;
  assign new_P2_R1095_U374 = ~new_P2_R1095_U158 | ~new_P2_R1095_U219;
  assign new_P2_R1095_U375 = ~new_P2_U3407 | ~new_P2_R1095_U41;
  assign new_P2_R1095_U376 = ~new_P2_U3070 | ~new_P2_R1095_U30;
  assign new_P2_R1095_U377 = ~new_P2_R1095_U376 | ~new_P2_R1095_U375;
  assign new_P2_R1095_U378 = ~new_P2_U3404 | ~new_P2_R1095_U42;
  assign new_P2_R1095_U379 = ~new_P2_U3066 | ~new_P2_R1095_U29;
  assign new_P2_R1095_U380 = ~new_P2_R1095_U240 | ~new_P2_R1095_U49;
  assign new_P2_R1095_U381 = ~new_P2_R1095_U159 | ~new_P2_R1095_U232;
  assign new_P2_R1095_U382 = ~new_P2_U3401 | ~new_P2_R1095_U43;
  assign new_P2_R1095_U383 = ~new_P2_U3059 | ~new_P2_R1095_U31;
  assign new_P2_R1095_U384 = ~new_P2_R1095_U161 | ~new_P2_R1095_U241;
  assign new_P2_R1095_U385 = ~new_P2_R1095_U345 | ~new_P2_R1095_U160;
  assign new_P2_R1095_U386 = ~new_P2_U3398 | ~new_P2_R1095_U36;
  assign new_P2_R1095_U387 = ~new_P2_U3063 | ~new_P2_R1095_U40;
  assign new_P2_R1095_U388 = ~new_P2_U3398 | ~new_P2_R1095_U36;
  assign new_P2_R1095_U389 = ~new_P2_U3063 | ~new_P2_R1095_U40;
  assign new_P2_R1095_U390 = ~new_P2_R1095_U389 | ~new_P2_R1095_U388;
  assign new_P2_R1095_U391 = ~new_P2_U3395 | ~new_P2_R1095_U34;
  assign new_P2_R1095_U392 = ~new_P2_U3067 | ~new_P2_R1095_U37;
  assign new_P2_R1095_U393 = ~new_P2_R1095_U243 | ~new_P2_R1095_U50;
  assign new_P2_R1095_U394 = ~new_P2_R1095_U162 | ~new_P2_R1095_U205;
  assign new_P2_R1095_U395 = ~new_P2_U3904 | ~new_P2_R1095_U164;
  assign new_P2_R1095_U396 = ~new_P2_U3054 | ~new_P2_R1095_U163;
  assign new_P2_R1095_U397 = ~new_P2_R1095_U396 | ~new_P2_R1095_U395;
  assign new_P2_R1095_U398 = ~new_P2_U3904 | ~new_P2_R1095_U164;
  assign new_P2_R1095_U399 = ~new_P2_U3054 | ~new_P2_R1095_U163;
  assign new_P2_R1095_U400 = ~new_P2_R1095_U51 | ~new_P2_U3053 | ~new_P2_R1095_U397;
  assign new_P2_R1095_U401 = ~new_P2_U3895 | ~new_P2_R1095_U16 | ~new_P2_R1095_U92;
  assign new_P2_R1095_U402 = ~new_P2_U3895 | ~new_P2_R1095_U92;
  assign new_P2_R1095_U403 = ~new_P2_U3053 | ~new_P2_R1095_U51;
  assign new_P2_R1095_U404 = ~new_P2_R1095_U138;
  assign new_P2_R1095_U405 = ~new_P2_R1095_U361 | ~new_P2_R1095_U404;
  assign new_P2_R1095_U406 = ~new_P2_R1095_U138 | ~new_P2_R1095_U166;
  assign new_P2_R1095_U407 = ~new_P2_U3896 | ~new_P2_R1095_U54;
  assign new_P2_R1095_U408 = ~new_P2_U3052 | ~new_P2_R1095_U91;
  assign new_P2_R1095_U409 = ~new_P2_U3896 | ~new_P2_R1095_U54;
  assign new_P2_R1095_U410 = ~new_P2_U3052 | ~new_P2_R1095_U91;
  assign new_P2_R1095_U411 = ~new_P2_R1095_U410 | ~new_P2_R1095_U409;
  assign new_P2_R1095_U412 = ~new_P2_U3897 | ~new_P2_R1095_U52;
  assign new_P2_R1095_U413 = ~new_P2_U3056 | ~new_P2_R1095_U90;
  assign new_P2_R1095_U414 = ~new_P2_R1095_U306 | ~new_P2_R1095_U93;
  assign new_P2_R1095_U415 = ~new_P2_R1095_U167 | ~new_P2_R1095_U298;
  assign new_P2_R1095_U416 = ~new_P2_U3898 | ~new_P2_R1095_U89;
  assign new_P2_R1095_U417 = ~new_P2_U3057 | ~new_P2_R1095_U88;
  assign new_P2_R1095_U418 = ~new_P2_R1095_U141;
  assign new_P2_R1095_U419 = ~new_P2_R1095_U294 | ~new_P2_R1095_U418;
  assign new_P2_R1095_U420 = ~new_P2_R1095_U141 | ~new_P2_R1095_U168;
  assign new_P2_R1095_U421 = ~new_P2_U3899 | ~new_P2_R1095_U87;
  assign new_P2_R1095_U422 = ~new_P2_U3064 | ~new_P2_R1095_U86;
  assign new_P2_R1095_U423 = ~new_P2_R1095_U142;
  assign new_P2_R1095_U424 = ~new_P2_R1095_U290 | ~new_P2_R1095_U423;
  assign new_P2_R1095_U425 = ~new_P2_R1095_U142 | ~new_P2_R1095_U169;
  assign new_P2_R1095_U426 = ~new_P2_U3900 | ~new_P2_R1095_U82;
  assign new_P2_R1095_U427 = ~new_P2_U3065 | ~new_P2_R1095_U79;
  assign new_P2_R1095_U428 = ~new_P2_R1095_U427 | ~new_P2_R1095_U426;
  assign new_P2_R1095_U429 = ~new_P2_U3901 | ~new_P2_R1095_U83;
  assign new_P2_R1095_U430 = ~new_P2_U3060 | ~new_P2_R1095_U80;
  assign new_P2_R1095_U431 = ~new_P2_R1095_U316 | ~new_P2_R1095_U94;
  assign new_P2_R1095_U432 = ~new_P2_R1095_U170 | ~new_P2_R1095_U308;
  assign new_P2_R1095_U433 = ~new_P2_U3902 | ~new_P2_R1095_U84;
  assign new_P2_R1095_U434 = ~new_P2_U3074 | ~new_P2_R1095_U81;
  assign new_P2_R1095_U435 = ~new_P2_R1095_U317 | ~new_P2_R1095_U172;
  assign new_P2_R1095_U436 = ~new_P2_R1095_U280 | ~new_P2_R1095_U171;
  assign new_P2_R1095_U437 = ~new_P2_U3903 | ~new_P2_R1095_U78;
  assign new_P2_R1095_U438 = ~new_P2_U3075 | ~new_P2_R1095_U77;
  assign new_P2_R1095_U439 = ~new_P2_R1095_U145;
  assign new_P2_R1095_U440 = ~new_P2_R1095_U276 | ~new_P2_R1095_U439;
  assign new_P2_R1095_U441 = ~new_P2_R1095_U145 | ~new_P2_R1095_U173;
  assign new_P2_R1095_U442 = ~new_P2_U3392 | ~new_P2_R1095_U39;
  assign new_P2_R1095_U443 = ~new_P2_U3077 | ~new_P2_R1095_U174;
  assign new_P2_R1095_U444 = ~new_P2_R1095_U146;
  assign new_P2_R1095_U445 = ~new_P2_R1095_U203 | ~new_P2_R1095_U444;
  assign new_P2_R1095_U446 = ~new_P2_R1095_U146 | ~new_P2_R1095_U175;
  assign new_P2_R1095_U447 = ~new_P2_U3445 | ~new_P2_R1095_U76;
  assign new_P2_R1095_U448 = ~new_P2_U3080 | ~new_P2_R1095_U75;
  assign new_P2_R1095_U449 = ~new_P2_R1095_U147;
  assign new_P2_R1095_U450 = ~new_P2_R1095_U272 | ~new_P2_R1095_U449;
  assign new_P2_R1095_U451 = ~new_P2_R1095_U147 | ~new_P2_R1095_U176;
  assign new_P2_R1095_U452 = ~new_P2_U3443 | ~new_P2_R1095_U74;
  assign new_P2_R1095_U453 = ~new_P2_U3081 | ~new_P2_R1095_U177;
  assign new_P2_R1095_U454 = ~new_P2_R1095_U148;
  assign new_P2_R1095_U455 = ~new_P2_R1095_U270 | ~new_P2_R1095_U454;
  assign new_P2_R1095_U456 = ~new_P2_R1095_U148 | ~new_P2_R1095_U178;
  assign new_P2_R1095_U457 = ~new_P2_U3440 | ~new_P2_R1095_U73;
  assign new_P2_R1095_U458 = ~new_P2_U3068 | ~new_P2_R1095_U72;
  assign new_P2_R1095_U459 = ~new_P2_R1095_U149;
  assign new_P2_R1095_U460 = ~new_P2_R1095_U266 | ~new_P2_R1095_U459;
  assign new_P2_R1095_U461 = ~new_P2_R1095_U149 | ~new_P2_R1095_U179;
  assign new_P2_R1095_U462 = ~new_P2_U3437 | ~new_P2_R1095_U68;
  assign new_P2_R1095_U463 = ~new_P2_U3072 | ~new_P2_R1095_U65;
  assign new_P2_R1095_U464 = ~new_P2_R1095_U463 | ~new_P2_R1095_U462;
  assign new_P2_R1095_U465 = ~new_P2_U3434 | ~new_P2_R1095_U69;
  assign new_P2_R1095_U466 = ~new_P2_U3073 | ~new_P2_R1095_U66;
  assign new_P2_R1095_U467 = ~new_P2_R1095_U327 | ~new_P2_R1095_U95;
  assign new_P2_R1095_U468 = ~new_P2_R1095_U180 | ~new_P2_R1095_U319;
  assign new_P2_R1095_U469 = ~new_P2_U3431 | ~new_P2_R1095_U70;
  assign new_P2_R1095_U470 = ~new_P2_U3078 | ~new_P2_R1095_U67;
  assign new_P2_R1095_U471 = ~new_P2_R1095_U328 | ~new_P2_R1095_U182;
  assign new_P2_R1095_U472 = ~new_P2_R1095_U256 | ~new_P2_R1095_U181;
  assign new_P2_R1095_U473 = ~new_P2_U3428 | ~new_P2_R1095_U64;
  assign new_P2_R1095_U474 = ~new_P2_U3079 | ~new_P2_R1095_U63;
  assign new_P2_R1095_U475 = ~new_P2_R1095_U152;
  assign new_P2_R1095_U476 = ~new_P2_R1095_U354 | ~new_P2_R1095_U475;
  assign new_P2_R1095_U477 = ~new_P2_R1095_U152 | ~new_P2_R1095_U183;
  assign new_P2_R1095_U478 = ~new_P2_U3425 | ~new_P2_R1095_U55;
  assign new_P2_R1095_U479 = ~new_P2_U3071 | ~new_P2_R1095_U61;
  assign new_P2_R1095_U480 = ~new_P2_R1095_U153;
  assign new_P2_R1095_U481 = ~new_P2_R1095_U352 | ~new_P2_R1095_U480;
  assign new_P2_R1095_U482 = ~new_P2_R1095_U153 | ~new_P2_R1095_U184;
  assign new_P2_R1095_U483 = ~new_P2_U3422 | ~new_P2_R1095_U56;
  assign new_P2_R1095_U484 = ~new_P2_U3062 | ~new_P2_R1095_U60;
  assign new_P2_R1095_U485 = ~new_P2_R1095_U484 | ~new_P2_R1095_U483;
  assign new_P2_R1095_U486 = ~new_P2_U3419 | ~new_P2_R1095_U57;
  assign new_P2_R1095_U487 = ~new_P2_U3061 | ~new_P2_R1095_U58;
  assign new_P2_R1095_U488 = ~new_P2_R1095_U96 | ~new_P2_R1095_U336;
  assign new_P2_R1095_U489 = ~new_P2_R1095_U185 | ~new_P2_R1095_U350;
  assign new_P2_R1212_U6 = ~new_P2_R1212_U176 | ~new_P2_R1212_U180;
  assign new_P2_R1212_U7 = ~new_P2_R1212_U9 | ~new_P2_R1212_U181;
  assign new_P2_R1212_U8 = ~P2_REG2_REG_0_;
  assign new_P2_R1212_U9 = ~P2_REG2_REG_0_ | ~new_P2_R1212_U48;
  assign new_P2_R1212_U10 = ~P2_REG2_REG_1_;
  assign new_P2_R1212_U11 = ~new_P2_U3391;
  assign new_P2_R1212_U12 = ~P2_REG2_REG_2_;
  assign new_P2_R1212_U13 = ~new_P2_U3394;
  assign new_P2_R1212_U14 = ~P2_REG2_REG_3_;
  assign new_P2_R1212_U15 = ~new_P2_U3397;
  assign new_P2_R1212_U16 = ~P2_REG2_REG_4_;
  assign new_P2_R1212_U17 = ~new_P2_U3400;
  assign new_P2_R1212_U18 = ~P2_REG2_REG_5_;
  assign new_P2_R1212_U19 = ~new_P2_U3403;
  assign new_P2_R1212_U20 = ~P2_REG2_REG_6_;
  assign new_P2_R1212_U21 = ~new_P2_U3406;
  assign new_P2_R1212_U22 = ~P2_REG2_REG_7_;
  assign new_P2_R1212_U23 = ~new_P2_U3409;
  assign new_P2_R1212_U24 = ~P2_REG2_REG_8_;
  assign new_P2_R1212_U25 = ~new_P2_U3412;
  assign new_P2_R1212_U26 = ~P2_REG2_REG_9_;
  assign new_P2_R1212_U27 = ~new_P2_U3415;
  assign new_P2_R1212_U28 = ~P2_REG2_REG_10_;
  assign new_P2_R1212_U29 = ~new_P2_U3418;
  assign new_P2_R1212_U30 = ~P2_REG2_REG_11_;
  assign new_P2_R1212_U31 = ~new_P2_U3421;
  assign new_P2_R1212_U32 = ~P2_REG2_REG_12_;
  assign new_P2_R1212_U33 = ~new_P2_U3424;
  assign new_P2_R1212_U34 = ~P2_REG2_REG_13_;
  assign new_P2_R1212_U35 = ~new_P2_U3427;
  assign new_P2_R1212_U36 = ~P2_REG2_REG_14_;
  assign new_P2_R1212_U37 = ~new_P2_U3430;
  assign new_P2_R1212_U38 = ~new_P2_R1212_U159 | ~new_P2_R1212_U158;
  assign new_P2_R1212_U39 = ~P2_REG2_REG_15_;
  assign new_P2_R1212_U40 = ~new_P2_U3433;
  assign new_P2_R1212_U41 = ~P2_REG2_REG_16_;
  assign new_P2_R1212_U42 = ~new_P2_U3436;
  assign new_P2_R1212_U43 = ~P2_REG2_REG_17_;
  assign new_P2_R1212_U44 = ~new_P2_U3439;
  assign new_P2_R1212_U45 = ~P2_REG2_REG_18_;
  assign new_P2_R1212_U46 = ~new_P2_U3442;
  assign new_P2_R1212_U47 = ~new_P2_R1212_U171 | ~new_P2_R1212_U170;
  assign new_P2_R1212_U48 = ~new_P2_U3386;
  assign new_P2_R1212_U49 = ~new_P2_R1212_U186 | ~new_P2_R1212_U185;
  assign new_P2_R1212_U50 = ~new_P2_R1212_U191 | ~new_P2_R1212_U190;
  assign new_P2_R1212_U51 = ~new_P2_R1212_U196 | ~new_P2_R1212_U195;
  assign new_P2_R1212_U52 = ~new_P2_R1212_U201 | ~new_P2_R1212_U200;
  assign new_P2_R1212_U53 = ~new_P2_R1212_U206 | ~new_P2_R1212_U205;
  assign new_P2_R1212_U54 = ~new_P2_R1212_U211 | ~new_P2_R1212_U210;
  assign new_P2_R1212_U55 = ~new_P2_R1212_U216 | ~new_P2_R1212_U215;
  assign new_P2_R1212_U56 = ~new_P2_R1212_U221 | ~new_P2_R1212_U220;
  assign new_P2_R1212_U57 = ~new_P2_R1212_U226 | ~new_P2_R1212_U225;
  assign new_P2_R1212_U58 = ~new_P2_R1212_U236 | ~new_P2_R1212_U235;
  assign new_P2_R1212_U59 = ~new_P2_R1212_U241 | ~new_P2_R1212_U240;
  assign new_P2_R1212_U60 = ~new_P2_R1212_U246 | ~new_P2_R1212_U245;
  assign new_P2_R1212_U61 = ~new_P2_R1212_U251 | ~new_P2_R1212_U250;
  assign new_P2_R1212_U62 = ~new_P2_R1212_U256 | ~new_P2_R1212_U255;
  assign new_P2_R1212_U63 = ~new_P2_R1212_U261 | ~new_P2_R1212_U260;
  assign new_P2_R1212_U64 = ~new_P2_R1212_U266 | ~new_P2_R1212_U265;
  assign new_P2_R1212_U65 = ~new_P2_R1212_U271 | ~new_P2_R1212_U270;
  assign new_P2_R1212_U66 = ~new_P2_R1212_U276 | ~new_P2_R1212_U275;
  assign new_P2_R1212_U67 = ~new_P2_R1212_U183 | ~new_P2_R1212_U182;
  assign new_P2_R1212_U68 = ~new_P2_R1212_U188 | ~new_P2_R1212_U187;
  assign new_P2_R1212_U69 = ~new_P2_R1212_U193 | ~new_P2_R1212_U192;
  assign new_P2_R1212_U70 = ~new_P2_R1212_U198 | ~new_P2_R1212_U197;
  assign new_P2_R1212_U71 = ~new_P2_R1212_U203 | ~new_P2_R1212_U202;
  assign new_P2_R1212_U72 = ~new_P2_R1212_U208 | ~new_P2_R1212_U207;
  assign new_P2_R1212_U73 = ~new_P2_R1212_U213 | ~new_P2_R1212_U212;
  assign new_P2_R1212_U74 = ~new_P2_R1212_U218 | ~new_P2_R1212_U217;
  assign new_P2_R1212_U75 = ~new_P2_R1212_U223 | ~new_P2_R1212_U222;
  assign new_P2_R1212_U76 = new_P2_R1212_U179 & new_P2_R1212_U228 & new_P2_R1212_U227;
  assign new_P2_R1212_U77 = new_P2_R1212_U175 & new_P2_R1212_U231;
  assign new_P2_R1212_U78 = ~new_P2_R1212_U233 | ~new_P2_R1212_U232;
  assign new_P2_R1212_U79 = ~new_P2_R1212_U238 | ~new_P2_R1212_U237;
  assign new_P2_R1212_U80 = ~new_P2_R1212_U243 | ~new_P2_R1212_U242;
  assign new_P2_R1212_U81 = ~new_P2_R1212_U248 | ~new_P2_R1212_U247;
  assign new_P2_R1212_U82 = ~new_P2_R1212_U253 | ~new_P2_R1212_U252;
  assign new_P2_R1212_U83 = ~new_P2_R1212_U258 | ~new_P2_R1212_U257;
  assign new_P2_R1212_U84 = ~new_P2_R1212_U263 | ~new_P2_R1212_U262;
  assign new_P2_R1212_U85 = ~new_P2_R1212_U268 | ~new_P2_R1212_U267;
  assign new_P2_R1212_U86 = ~new_P2_R1212_U273 | ~new_P2_R1212_U272;
  assign new_P2_R1212_U87 = ~new_P2_R1212_U135 | ~new_P2_R1212_U134;
  assign new_P2_R1212_U88 = ~new_P2_R1212_U131 | ~new_P2_R1212_U130;
  assign new_P2_R1212_U89 = ~new_P2_R1212_U127 | ~new_P2_R1212_U126;
  assign new_P2_R1212_U90 = ~new_P2_R1212_U123 | ~new_P2_R1212_U122;
  assign new_P2_R1212_U91 = ~new_P2_R1212_U119 | ~new_P2_R1212_U118;
  assign new_P2_R1212_U92 = ~new_P2_R1212_U115 | ~new_P2_R1212_U114;
  assign new_P2_R1212_U93 = ~new_P2_R1212_U111 | ~new_P2_R1212_U110;
  assign new_P2_R1212_U94 = ~new_P2_R1212_U107 | ~new_P2_R1212_U106;
  assign new_P2_R1212_U95 = ~P2_REG2_REG_19_;
  assign new_P2_R1212_U96 = ~new_P2_U3379;
  assign new_P2_R1212_U97 = ~new_P2_R1212_U167 | ~new_P2_R1212_U166;
  assign new_P2_R1212_U98 = ~new_P2_R1212_U163 | ~new_P2_R1212_U162;
  assign new_P2_R1212_U99 = ~new_P2_R1212_U155 | ~new_P2_R1212_U154;
  assign new_P2_R1212_U100 = ~new_P2_R1212_U151 | ~new_P2_R1212_U150;
  assign new_P2_R1212_U101 = ~new_P2_R1212_U147 | ~new_P2_R1212_U146;
  assign new_P2_R1212_U102 = ~new_P2_R1212_U143 | ~new_P2_R1212_U142;
  assign new_P2_R1212_U103 = ~new_P2_R1212_U139 | ~new_P2_R1212_U138;
  assign new_P2_R1212_U104 = ~new_P2_R1212_U9;
  assign new_P2_R1212_U105 = ~P2_REG2_REG_1_ | ~new_P2_R1212_U104;
  assign new_P2_R1212_U106 = ~new_P2_U3391 | ~new_P2_R1212_U105;
  assign new_P2_R1212_U107 = ~new_P2_R1212_U9 | ~new_P2_R1212_U10;
  assign new_P2_R1212_U108 = ~new_P2_R1212_U94;
  assign new_P2_R1212_U109 = ~P2_REG2_REG_2_ | ~new_P2_R1212_U13;
  assign new_P2_R1212_U110 = ~new_P2_R1212_U109 | ~new_P2_R1212_U94;
  assign new_P2_R1212_U111 = ~new_P2_U3394 | ~new_P2_R1212_U12;
  assign new_P2_R1212_U112 = ~new_P2_R1212_U93;
  assign new_P2_R1212_U113 = ~P2_REG2_REG_3_ | ~new_P2_R1212_U15;
  assign new_P2_R1212_U114 = ~new_P2_R1212_U113 | ~new_P2_R1212_U93;
  assign new_P2_R1212_U115 = ~new_P2_U3397 | ~new_P2_R1212_U14;
  assign new_P2_R1212_U116 = ~new_P2_R1212_U92;
  assign new_P2_R1212_U117 = ~P2_REG2_REG_4_ | ~new_P2_R1212_U17;
  assign new_P2_R1212_U118 = ~new_P2_R1212_U117 | ~new_P2_R1212_U92;
  assign new_P2_R1212_U119 = ~new_P2_U3400 | ~new_P2_R1212_U16;
  assign new_P2_R1212_U120 = ~new_P2_R1212_U91;
  assign new_P2_R1212_U121 = ~P2_REG2_REG_5_ | ~new_P2_R1212_U19;
  assign new_P2_R1212_U122 = ~new_P2_R1212_U121 | ~new_P2_R1212_U91;
  assign new_P2_R1212_U123 = ~new_P2_U3403 | ~new_P2_R1212_U18;
  assign new_P2_R1212_U124 = ~new_P2_R1212_U90;
  assign new_P2_R1212_U125 = ~P2_REG2_REG_6_ | ~new_P2_R1212_U21;
  assign new_P2_R1212_U126 = ~new_P2_R1212_U125 | ~new_P2_R1212_U90;
  assign new_P2_R1212_U127 = ~new_P2_U3406 | ~new_P2_R1212_U20;
  assign new_P2_R1212_U128 = ~new_P2_R1212_U89;
  assign new_P2_R1212_U129 = ~P2_REG2_REG_7_ | ~new_P2_R1212_U23;
  assign new_P2_R1212_U130 = ~new_P2_R1212_U129 | ~new_P2_R1212_U89;
  assign new_P2_R1212_U131 = ~new_P2_U3409 | ~new_P2_R1212_U22;
  assign new_P2_R1212_U132 = ~new_P2_R1212_U88;
  assign new_P2_R1212_U133 = ~P2_REG2_REG_8_ | ~new_P2_R1212_U25;
  assign new_P2_R1212_U134 = ~new_P2_R1212_U133 | ~new_P2_R1212_U88;
  assign new_P2_R1212_U135 = ~new_P2_U3412 | ~new_P2_R1212_U24;
  assign new_P2_R1212_U136 = ~new_P2_R1212_U87;
  assign new_P2_R1212_U137 = ~P2_REG2_REG_9_ | ~new_P2_R1212_U27;
  assign new_P2_R1212_U138 = ~new_P2_R1212_U137 | ~new_P2_R1212_U87;
  assign new_P2_R1212_U139 = ~new_P2_U3415 | ~new_P2_R1212_U26;
  assign new_P2_R1212_U140 = ~new_P2_R1212_U103;
  assign new_P2_R1212_U141 = ~P2_REG2_REG_10_ | ~new_P2_R1212_U29;
  assign new_P2_R1212_U142 = ~new_P2_R1212_U141 | ~new_P2_R1212_U103;
  assign new_P2_R1212_U143 = ~new_P2_U3418 | ~new_P2_R1212_U28;
  assign new_P2_R1212_U144 = ~new_P2_R1212_U102;
  assign new_P2_R1212_U145 = ~P2_REG2_REG_11_ | ~new_P2_R1212_U31;
  assign new_P2_R1212_U146 = ~new_P2_R1212_U145 | ~new_P2_R1212_U102;
  assign new_P2_R1212_U147 = ~new_P2_U3421 | ~new_P2_R1212_U30;
  assign new_P2_R1212_U148 = ~new_P2_R1212_U101;
  assign new_P2_R1212_U149 = ~P2_REG2_REG_12_ | ~new_P2_R1212_U33;
  assign new_P2_R1212_U150 = ~new_P2_R1212_U149 | ~new_P2_R1212_U101;
  assign new_P2_R1212_U151 = ~new_P2_U3424 | ~new_P2_R1212_U32;
  assign new_P2_R1212_U152 = ~new_P2_R1212_U100;
  assign new_P2_R1212_U153 = ~P2_REG2_REG_13_ | ~new_P2_R1212_U35;
  assign new_P2_R1212_U154 = ~new_P2_R1212_U153 | ~new_P2_R1212_U100;
  assign new_P2_R1212_U155 = ~new_P2_U3427 | ~new_P2_R1212_U34;
  assign new_P2_R1212_U156 = ~new_P2_R1212_U99;
  assign new_P2_R1212_U157 = ~P2_REG2_REG_14_ | ~new_P2_R1212_U37;
  assign new_P2_R1212_U158 = ~new_P2_R1212_U157 | ~new_P2_R1212_U99;
  assign new_P2_R1212_U159 = ~new_P2_U3430 | ~new_P2_R1212_U36;
  assign new_P2_R1212_U160 = ~new_P2_R1212_U38;
  assign new_P2_R1212_U161 = ~P2_REG2_REG_15_ | ~new_P2_R1212_U160;
  assign new_P2_R1212_U162 = ~new_P2_U3433 | ~new_P2_R1212_U161;
  assign new_P2_R1212_U163 = ~new_P2_R1212_U38 | ~new_P2_R1212_U39;
  assign new_P2_R1212_U164 = ~new_P2_R1212_U98;
  assign new_P2_R1212_U165 = ~P2_REG2_REG_16_ | ~new_P2_R1212_U42;
  assign new_P2_R1212_U166 = ~new_P2_R1212_U165 | ~new_P2_R1212_U98;
  assign new_P2_R1212_U167 = ~new_P2_U3436 | ~new_P2_R1212_U41;
  assign new_P2_R1212_U168 = ~new_P2_R1212_U97;
  assign new_P2_R1212_U169 = ~P2_REG2_REG_17_ | ~new_P2_R1212_U44;
  assign new_P2_R1212_U170 = ~new_P2_R1212_U169 | ~new_P2_R1212_U97;
  assign new_P2_R1212_U171 = ~new_P2_U3439 | ~new_P2_R1212_U43;
  assign new_P2_R1212_U172 = ~new_P2_R1212_U47;
  assign new_P2_R1212_U173 = ~new_P2_U3442 | ~new_P2_R1212_U45;
  assign new_P2_R1212_U174 = ~new_P2_R1212_U172 | ~new_P2_R1212_U173;
  assign new_P2_R1212_U175 = ~P2_REG2_REG_18_ | ~new_P2_R1212_U46;
  assign new_P2_R1212_U176 = ~new_P2_R1212_U77 | ~new_P2_R1212_U174;
  assign new_P2_R1212_U177 = ~P2_REG2_REG_18_ | ~new_P2_R1212_U46;
  assign new_P2_R1212_U178 = ~new_P2_R1212_U177 | ~new_P2_R1212_U47;
  assign new_P2_R1212_U179 = ~new_P2_U3442 | ~new_P2_R1212_U45;
  assign new_P2_R1212_U180 = ~new_P2_R1212_U76 | ~new_P2_R1212_U178;
  assign new_P2_R1212_U181 = ~new_P2_U3386 | ~new_P2_R1212_U8;
  assign new_P2_R1212_U182 = ~P2_REG2_REG_9_ | ~new_P2_R1212_U27;
  assign new_P2_R1212_U183 = ~new_P2_U3415 | ~new_P2_R1212_U26;
  assign new_P2_R1212_U184 = ~new_P2_R1212_U67;
  assign new_P2_R1212_U185 = ~new_P2_R1212_U136 | ~new_P2_R1212_U184;
  assign new_P2_R1212_U186 = ~new_P2_R1212_U67 | ~new_P2_R1212_U87;
  assign new_P2_R1212_U187 = ~P2_REG2_REG_8_ | ~new_P2_R1212_U25;
  assign new_P2_R1212_U188 = ~new_P2_U3412 | ~new_P2_R1212_U24;
  assign new_P2_R1212_U189 = ~new_P2_R1212_U68;
  assign new_P2_R1212_U190 = ~new_P2_R1212_U132 | ~new_P2_R1212_U189;
  assign new_P2_R1212_U191 = ~new_P2_R1212_U68 | ~new_P2_R1212_U88;
  assign new_P2_R1212_U192 = ~P2_REG2_REG_7_ | ~new_P2_R1212_U23;
  assign new_P2_R1212_U193 = ~new_P2_U3409 | ~new_P2_R1212_U22;
  assign new_P2_R1212_U194 = ~new_P2_R1212_U69;
  assign new_P2_R1212_U195 = ~new_P2_R1212_U128 | ~new_P2_R1212_U194;
  assign new_P2_R1212_U196 = ~new_P2_R1212_U69 | ~new_P2_R1212_U89;
  assign new_P2_R1212_U197 = ~P2_REG2_REG_6_ | ~new_P2_R1212_U21;
  assign new_P2_R1212_U198 = ~new_P2_U3406 | ~new_P2_R1212_U20;
  assign new_P2_R1212_U199 = ~new_P2_R1212_U70;
  assign new_P2_R1212_U200 = ~new_P2_R1212_U124 | ~new_P2_R1212_U199;
  assign new_P2_R1212_U201 = ~new_P2_R1212_U70 | ~new_P2_R1212_U90;
  assign new_P2_R1212_U202 = ~P2_REG2_REG_5_ | ~new_P2_R1212_U19;
  assign new_P2_R1212_U203 = ~new_P2_U3403 | ~new_P2_R1212_U18;
  assign new_P2_R1212_U204 = ~new_P2_R1212_U71;
  assign new_P2_R1212_U205 = ~new_P2_R1212_U120 | ~new_P2_R1212_U204;
  assign new_P2_R1212_U206 = ~new_P2_R1212_U71 | ~new_P2_R1212_U91;
  assign new_P2_R1212_U207 = ~P2_REG2_REG_4_ | ~new_P2_R1212_U17;
  assign new_P2_R1212_U208 = ~new_P2_U3400 | ~new_P2_R1212_U16;
  assign new_P2_R1212_U209 = ~new_P2_R1212_U72;
  assign new_P2_R1212_U210 = ~new_P2_R1212_U116 | ~new_P2_R1212_U209;
  assign new_P2_R1212_U211 = ~new_P2_R1212_U72 | ~new_P2_R1212_U92;
  assign new_P2_R1212_U212 = ~P2_REG2_REG_3_ | ~new_P2_R1212_U15;
  assign new_P2_R1212_U213 = ~new_P2_U3397 | ~new_P2_R1212_U14;
  assign new_P2_R1212_U214 = ~new_P2_R1212_U73;
  assign new_P2_R1212_U215 = ~new_P2_R1212_U112 | ~new_P2_R1212_U214;
  assign new_P2_R1212_U216 = ~new_P2_R1212_U73 | ~new_P2_R1212_U93;
  assign new_P2_R1212_U217 = ~P2_REG2_REG_2_ | ~new_P2_R1212_U13;
  assign new_P2_R1212_U218 = ~new_P2_U3394 | ~new_P2_R1212_U12;
  assign new_P2_R1212_U219 = ~new_P2_R1212_U74;
  assign new_P2_R1212_U220 = ~new_P2_R1212_U108 | ~new_P2_R1212_U219;
  assign new_P2_R1212_U221 = ~new_P2_R1212_U74 | ~new_P2_R1212_U94;
  assign new_P2_R1212_U222 = ~new_P2_R1212_U104 | ~new_P2_R1212_U10;
  assign new_P2_R1212_U223 = ~P2_REG2_REG_1_ | ~new_P2_R1212_U9;
  assign new_P2_R1212_U224 = ~new_P2_R1212_U75;
  assign new_P2_R1212_U225 = ~new_P2_R1212_U224 | ~new_P2_U3391;
  assign new_P2_R1212_U226 = ~new_P2_R1212_U75 | ~new_P2_R1212_U11;
  assign new_P2_R1212_U227 = ~P2_REG2_REG_19_ | ~new_P2_R1212_U96;
  assign new_P2_R1212_U228 = ~new_P2_U3379 | ~new_P2_R1212_U95;
  assign new_P2_R1212_U229 = ~P2_REG2_REG_19_ | ~new_P2_R1212_U96;
  assign new_P2_R1212_U230 = ~new_P2_U3379 | ~new_P2_R1212_U95;
  assign new_P2_R1212_U231 = ~new_P2_R1212_U230 | ~new_P2_R1212_U229;
  assign new_P2_R1212_U232 = ~P2_REG2_REG_18_ | ~new_P2_R1212_U46;
  assign new_P2_R1212_U233 = ~new_P2_U3442 | ~new_P2_R1212_U45;
  assign new_P2_R1212_U234 = ~new_P2_R1212_U78;
  assign new_P2_R1212_U235 = ~new_P2_R1212_U234 | ~new_P2_R1212_U172;
  assign new_P2_R1212_U236 = ~new_P2_R1212_U78 | ~new_P2_R1212_U47;
  assign new_P2_R1212_U237 = ~P2_REG2_REG_17_ | ~new_P2_R1212_U44;
  assign new_P2_R1212_U238 = ~new_P2_U3439 | ~new_P2_R1212_U43;
  assign new_P2_R1212_U239 = ~new_P2_R1212_U79;
  assign new_P2_R1212_U240 = ~new_P2_R1212_U168 | ~new_P2_R1212_U239;
  assign new_P2_R1212_U241 = ~new_P2_R1212_U79 | ~new_P2_R1212_U97;
  assign new_P2_R1212_U242 = ~P2_REG2_REG_16_ | ~new_P2_R1212_U42;
  assign new_P2_R1212_U243 = ~new_P2_U3436 | ~new_P2_R1212_U41;
  assign new_P2_R1212_U244 = ~new_P2_R1212_U80;
  assign new_P2_R1212_U245 = ~new_P2_R1212_U164 | ~new_P2_R1212_U244;
  assign new_P2_R1212_U246 = ~new_P2_R1212_U80 | ~new_P2_R1212_U98;
  assign new_P2_R1212_U247 = ~new_P2_U3433 | ~new_P2_R1212_U39;
  assign new_P2_R1212_U248 = ~P2_REG2_REG_15_ | ~new_P2_R1212_U40;
  assign new_P2_R1212_U249 = ~new_P2_R1212_U81;
  assign new_P2_R1212_U250 = ~new_P2_R1212_U249 | ~new_P2_R1212_U160;
  assign new_P2_R1212_U251 = ~new_P2_R1212_U81 | ~new_P2_R1212_U38;
  assign new_P2_R1212_U252 = ~P2_REG2_REG_14_ | ~new_P2_R1212_U37;
  assign new_P2_R1212_U253 = ~new_P2_U3430 | ~new_P2_R1212_U36;
  assign new_P2_R1212_U254 = ~new_P2_R1212_U82;
  assign new_P2_R1212_U255 = ~new_P2_R1212_U156 | ~new_P2_R1212_U254;
  assign new_P2_R1212_U256 = ~new_P2_R1212_U82 | ~new_P2_R1212_U99;
  assign new_P2_R1212_U257 = ~P2_REG2_REG_13_ | ~new_P2_R1212_U35;
  assign new_P2_R1212_U258 = ~new_P2_U3427 | ~new_P2_R1212_U34;
  assign new_P2_R1212_U259 = ~new_P2_R1212_U83;
  assign new_P2_R1212_U260 = ~new_P2_R1212_U152 | ~new_P2_R1212_U259;
  assign new_P2_R1212_U261 = ~new_P2_R1212_U83 | ~new_P2_R1212_U100;
  assign new_P2_R1212_U262 = ~P2_REG2_REG_12_ | ~new_P2_R1212_U33;
  assign new_P2_R1212_U263 = ~new_P2_U3424 | ~new_P2_R1212_U32;
  assign new_P2_R1212_U264 = ~new_P2_R1212_U84;
  assign new_P2_R1212_U265 = ~new_P2_R1212_U148 | ~new_P2_R1212_U264;
  assign new_P2_R1212_U266 = ~new_P2_R1212_U84 | ~new_P2_R1212_U101;
  assign new_P2_R1212_U267 = ~P2_REG2_REG_11_ | ~new_P2_R1212_U31;
  assign new_P2_R1212_U268 = ~new_P2_U3421 | ~new_P2_R1212_U30;
  assign new_P2_R1212_U269 = ~new_P2_R1212_U85;
  assign new_P2_R1212_U270 = ~new_P2_R1212_U144 | ~new_P2_R1212_U269;
  assign new_P2_R1212_U271 = ~new_P2_R1212_U85 | ~new_P2_R1212_U102;
  assign new_P2_R1212_U272 = ~P2_REG2_REG_10_ | ~new_P2_R1212_U29;
  assign new_P2_R1212_U273 = ~new_P2_U3418 | ~new_P2_R1212_U28;
  assign new_P2_R1212_U274 = ~new_P2_R1212_U86;
  assign new_P2_R1212_U275 = ~new_P2_R1212_U140 | ~new_P2_R1212_U274;
  assign new_P2_R1212_U276 = ~new_P2_R1212_U86 | ~new_P2_R1212_U103;
  assign new_P2_R1209_U6 = ~new_P2_R1209_U176 | ~new_P2_R1209_U180;
  assign new_P2_R1209_U7 = ~new_P2_R1209_U9 | ~new_P2_R1209_U181;
  assign new_P2_R1209_U8 = ~P2_REG1_REG_0_;
  assign new_P2_R1209_U9 = ~P2_REG1_REG_0_ | ~new_P2_R1209_U48;
  assign new_P2_R1209_U10 = ~P2_REG1_REG_1_;
  assign new_P2_R1209_U11 = ~new_P2_U3391;
  assign new_P2_R1209_U12 = ~P2_REG1_REG_2_;
  assign new_P2_R1209_U13 = ~new_P2_U3394;
  assign new_P2_R1209_U14 = ~P2_REG1_REG_3_;
  assign new_P2_R1209_U15 = ~new_P2_U3397;
  assign new_P2_R1209_U16 = ~P2_REG1_REG_4_;
  assign new_P2_R1209_U17 = ~new_P2_U3400;
  assign new_P2_R1209_U18 = ~P2_REG1_REG_5_;
  assign new_P2_R1209_U19 = ~new_P2_U3403;
  assign new_P2_R1209_U20 = ~P2_REG1_REG_6_;
  assign new_P2_R1209_U21 = ~new_P2_U3406;
  assign new_P2_R1209_U22 = ~P2_REG1_REG_7_;
  assign new_P2_R1209_U23 = ~new_P2_U3409;
  assign new_P2_R1209_U24 = ~P2_REG1_REG_8_;
  assign new_P2_R1209_U25 = ~new_P2_U3412;
  assign new_P2_R1209_U26 = ~P2_REG1_REG_9_;
  assign new_P2_R1209_U27 = ~new_P2_U3415;
  assign new_P2_R1209_U28 = ~P2_REG1_REG_10_;
  assign new_P2_R1209_U29 = ~new_P2_U3418;
  assign new_P2_R1209_U30 = ~P2_REG1_REG_11_;
  assign new_P2_R1209_U31 = ~new_P2_U3421;
  assign new_P2_R1209_U32 = ~P2_REG1_REG_12_;
  assign new_P2_R1209_U33 = ~new_P2_U3424;
  assign new_P2_R1209_U34 = ~P2_REG1_REG_13_;
  assign new_P2_R1209_U35 = ~new_P2_U3427;
  assign new_P2_R1209_U36 = ~P2_REG1_REG_14_;
  assign new_P2_R1209_U37 = ~new_P2_U3430;
  assign new_P2_R1209_U38 = ~new_P2_R1209_U159 | ~new_P2_R1209_U158;
  assign new_P2_R1209_U39 = ~P2_REG1_REG_15_;
  assign new_P2_R1209_U40 = ~new_P2_U3433;
  assign new_P2_R1209_U41 = ~P2_REG1_REG_16_;
  assign new_P2_R1209_U42 = ~new_P2_U3436;
  assign new_P2_R1209_U43 = ~P2_REG1_REG_17_;
  assign new_P2_R1209_U44 = ~new_P2_U3439;
  assign new_P2_R1209_U45 = ~P2_REG1_REG_18_;
  assign new_P2_R1209_U46 = ~new_P2_U3442;
  assign new_P2_R1209_U47 = ~new_P2_R1209_U171 | ~new_P2_R1209_U170;
  assign new_P2_R1209_U48 = ~new_P2_U3386;
  assign new_P2_R1209_U49 = ~new_P2_R1209_U186 | ~new_P2_R1209_U185;
  assign new_P2_R1209_U50 = ~new_P2_R1209_U191 | ~new_P2_R1209_U190;
  assign new_P2_R1209_U51 = ~new_P2_R1209_U196 | ~new_P2_R1209_U195;
  assign new_P2_R1209_U52 = ~new_P2_R1209_U201 | ~new_P2_R1209_U200;
  assign new_P2_R1209_U53 = ~new_P2_R1209_U206 | ~new_P2_R1209_U205;
  assign new_P2_R1209_U54 = ~new_P2_R1209_U211 | ~new_P2_R1209_U210;
  assign new_P2_R1209_U55 = ~new_P2_R1209_U216 | ~new_P2_R1209_U215;
  assign new_P2_R1209_U56 = ~new_P2_R1209_U221 | ~new_P2_R1209_U220;
  assign new_P2_R1209_U57 = ~new_P2_R1209_U226 | ~new_P2_R1209_U225;
  assign new_P2_R1209_U58 = ~new_P2_R1209_U236 | ~new_P2_R1209_U235;
  assign new_P2_R1209_U59 = ~new_P2_R1209_U241 | ~new_P2_R1209_U240;
  assign new_P2_R1209_U60 = ~new_P2_R1209_U246 | ~new_P2_R1209_U245;
  assign new_P2_R1209_U61 = ~new_P2_R1209_U251 | ~new_P2_R1209_U250;
  assign new_P2_R1209_U62 = ~new_P2_R1209_U256 | ~new_P2_R1209_U255;
  assign new_P2_R1209_U63 = ~new_P2_R1209_U261 | ~new_P2_R1209_U260;
  assign new_P2_R1209_U64 = ~new_P2_R1209_U266 | ~new_P2_R1209_U265;
  assign new_P2_R1209_U65 = ~new_P2_R1209_U271 | ~new_P2_R1209_U270;
  assign new_P2_R1209_U66 = ~new_P2_R1209_U276 | ~new_P2_R1209_U275;
  assign new_P2_R1209_U67 = ~new_P2_R1209_U183 | ~new_P2_R1209_U182;
  assign new_P2_R1209_U68 = ~new_P2_R1209_U188 | ~new_P2_R1209_U187;
  assign new_P2_R1209_U69 = ~new_P2_R1209_U193 | ~new_P2_R1209_U192;
  assign new_P2_R1209_U70 = ~new_P2_R1209_U198 | ~new_P2_R1209_U197;
  assign new_P2_R1209_U71 = ~new_P2_R1209_U203 | ~new_P2_R1209_U202;
  assign new_P2_R1209_U72 = ~new_P2_R1209_U208 | ~new_P2_R1209_U207;
  assign new_P2_R1209_U73 = ~new_P2_R1209_U213 | ~new_P2_R1209_U212;
  assign new_P2_R1209_U74 = ~new_P2_R1209_U218 | ~new_P2_R1209_U217;
  assign new_P2_R1209_U75 = ~new_P2_R1209_U223 | ~new_P2_R1209_U222;
  assign new_P2_R1209_U76 = new_P2_R1209_U179 & new_P2_R1209_U228 & new_P2_R1209_U227;
  assign new_P2_R1209_U77 = new_P2_R1209_U175 & new_P2_R1209_U231;
  assign new_P2_R1209_U78 = ~new_P2_R1209_U233 | ~new_P2_R1209_U232;
  assign new_P2_R1209_U79 = ~new_P2_R1209_U238 | ~new_P2_R1209_U237;
  assign new_P2_R1209_U80 = ~new_P2_R1209_U243 | ~new_P2_R1209_U242;
  assign new_P2_R1209_U81 = ~new_P2_R1209_U248 | ~new_P2_R1209_U247;
  assign new_P2_R1209_U82 = ~new_P2_R1209_U253 | ~new_P2_R1209_U252;
  assign new_P2_R1209_U83 = ~new_P2_R1209_U258 | ~new_P2_R1209_U257;
  assign new_P2_R1209_U84 = ~new_P2_R1209_U263 | ~new_P2_R1209_U262;
  assign new_P2_R1209_U85 = ~new_P2_R1209_U268 | ~new_P2_R1209_U267;
  assign new_P2_R1209_U86 = ~new_P2_R1209_U273 | ~new_P2_R1209_U272;
  assign new_P2_R1209_U87 = ~new_P2_R1209_U135 | ~new_P2_R1209_U134;
  assign new_P2_R1209_U88 = ~new_P2_R1209_U131 | ~new_P2_R1209_U130;
  assign new_P2_R1209_U89 = ~new_P2_R1209_U127 | ~new_P2_R1209_U126;
  assign new_P2_R1209_U90 = ~new_P2_R1209_U123 | ~new_P2_R1209_U122;
  assign new_P2_R1209_U91 = ~new_P2_R1209_U119 | ~new_P2_R1209_U118;
  assign new_P2_R1209_U92 = ~new_P2_R1209_U115 | ~new_P2_R1209_U114;
  assign new_P2_R1209_U93 = ~new_P2_R1209_U111 | ~new_P2_R1209_U110;
  assign new_P2_R1209_U94 = ~new_P2_R1209_U107 | ~new_P2_R1209_U106;
  assign new_P2_R1209_U95 = ~P2_REG1_REG_19_;
  assign new_P2_R1209_U96 = ~new_P2_U3379;
  assign new_P2_R1209_U97 = ~new_P2_R1209_U167 | ~new_P2_R1209_U166;
  assign new_P2_R1209_U98 = ~new_P2_R1209_U163 | ~new_P2_R1209_U162;
  assign new_P2_R1209_U99 = ~new_P2_R1209_U155 | ~new_P2_R1209_U154;
  assign new_P2_R1209_U100 = ~new_P2_R1209_U151 | ~new_P2_R1209_U150;
  assign new_P2_R1209_U101 = ~new_P2_R1209_U147 | ~new_P2_R1209_U146;
  assign new_P2_R1209_U102 = ~new_P2_R1209_U143 | ~new_P2_R1209_U142;
  assign new_P2_R1209_U103 = ~new_P2_R1209_U139 | ~new_P2_R1209_U138;
  assign new_P2_R1209_U104 = ~new_P2_R1209_U9;
  assign new_P2_R1209_U105 = ~P2_REG1_REG_1_ | ~new_P2_R1209_U104;
  assign new_P2_R1209_U106 = ~new_P2_U3391 | ~new_P2_R1209_U105;
  assign new_P2_R1209_U107 = ~new_P2_R1209_U9 | ~new_P2_R1209_U10;
  assign new_P2_R1209_U108 = ~new_P2_R1209_U94;
  assign new_P2_R1209_U109 = ~P2_REG1_REG_2_ | ~new_P2_R1209_U13;
  assign new_P2_R1209_U110 = ~new_P2_R1209_U109 | ~new_P2_R1209_U94;
  assign new_P2_R1209_U111 = ~new_P2_U3394 | ~new_P2_R1209_U12;
  assign new_P2_R1209_U112 = ~new_P2_R1209_U93;
  assign new_P2_R1209_U113 = ~P2_REG1_REG_3_ | ~new_P2_R1209_U15;
  assign new_P2_R1209_U114 = ~new_P2_R1209_U113 | ~new_P2_R1209_U93;
  assign new_P2_R1209_U115 = ~new_P2_U3397 | ~new_P2_R1209_U14;
  assign new_P2_R1209_U116 = ~new_P2_R1209_U92;
  assign new_P2_R1209_U117 = ~P2_REG1_REG_4_ | ~new_P2_R1209_U17;
  assign new_P2_R1209_U118 = ~new_P2_R1209_U117 | ~new_P2_R1209_U92;
  assign new_P2_R1209_U119 = ~new_P2_U3400 | ~new_P2_R1209_U16;
  assign new_P2_R1209_U120 = ~new_P2_R1209_U91;
  assign new_P2_R1209_U121 = ~P2_REG1_REG_5_ | ~new_P2_R1209_U19;
  assign new_P2_R1209_U122 = ~new_P2_R1209_U121 | ~new_P2_R1209_U91;
  assign new_P2_R1209_U123 = ~new_P2_U3403 | ~new_P2_R1209_U18;
  assign new_P2_R1209_U124 = ~new_P2_R1209_U90;
  assign new_P2_R1209_U125 = ~P2_REG1_REG_6_ | ~new_P2_R1209_U21;
  assign new_P2_R1209_U126 = ~new_P2_R1209_U125 | ~new_P2_R1209_U90;
  assign new_P2_R1209_U127 = ~new_P2_U3406 | ~new_P2_R1209_U20;
  assign new_P2_R1209_U128 = ~new_P2_R1209_U89;
  assign new_P2_R1209_U129 = ~P2_REG1_REG_7_ | ~new_P2_R1209_U23;
  assign new_P2_R1209_U130 = ~new_P2_R1209_U129 | ~new_P2_R1209_U89;
  assign new_P2_R1209_U131 = ~new_P2_U3409 | ~new_P2_R1209_U22;
  assign new_P2_R1209_U132 = ~new_P2_R1209_U88;
  assign new_P2_R1209_U133 = ~P2_REG1_REG_8_ | ~new_P2_R1209_U25;
  assign new_P2_R1209_U134 = ~new_P2_R1209_U133 | ~new_P2_R1209_U88;
  assign new_P2_R1209_U135 = ~new_P2_U3412 | ~new_P2_R1209_U24;
  assign new_P2_R1209_U136 = ~new_P2_R1209_U87;
  assign new_P2_R1209_U137 = ~P2_REG1_REG_9_ | ~new_P2_R1209_U27;
  assign new_P2_R1209_U138 = ~new_P2_R1209_U137 | ~new_P2_R1209_U87;
  assign new_P2_R1209_U139 = ~new_P2_U3415 | ~new_P2_R1209_U26;
  assign new_P2_R1209_U140 = ~new_P2_R1209_U103;
  assign new_P2_R1209_U141 = ~P2_REG1_REG_10_ | ~new_P2_R1209_U29;
  assign new_P2_R1209_U142 = ~new_P2_R1209_U141 | ~new_P2_R1209_U103;
  assign new_P2_R1209_U143 = ~new_P2_U3418 | ~new_P2_R1209_U28;
  assign new_P2_R1209_U144 = ~new_P2_R1209_U102;
  assign new_P2_R1209_U145 = ~P2_REG1_REG_11_ | ~new_P2_R1209_U31;
  assign new_P2_R1209_U146 = ~new_P2_R1209_U145 | ~new_P2_R1209_U102;
  assign new_P2_R1209_U147 = ~new_P2_U3421 | ~new_P2_R1209_U30;
  assign new_P2_R1209_U148 = ~new_P2_R1209_U101;
  assign new_P2_R1209_U149 = ~P2_REG1_REG_12_ | ~new_P2_R1209_U33;
  assign new_P2_R1209_U150 = ~new_P2_R1209_U149 | ~new_P2_R1209_U101;
  assign new_P2_R1209_U151 = ~new_P2_U3424 | ~new_P2_R1209_U32;
  assign new_P2_R1209_U152 = ~new_P2_R1209_U100;
  assign new_P2_R1209_U153 = ~P2_REG1_REG_13_ | ~new_P2_R1209_U35;
  assign new_P2_R1209_U154 = ~new_P2_R1209_U153 | ~new_P2_R1209_U100;
  assign new_P2_R1209_U155 = ~new_P2_U3427 | ~new_P2_R1209_U34;
  assign new_P2_R1209_U156 = ~new_P2_R1209_U99;
  assign new_P2_R1209_U157 = ~P2_REG1_REG_14_ | ~new_P2_R1209_U37;
  assign new_P2_R1209_U158 = ~new_P2_R1209_U157 | ~new_P2_R1209_U99;
  assign new_P2_R1209_U159 = ~new_P2_U3430 | ~new_P2_R1209_U36;
  assign new_P2_R1209_U160 = ~new_P2_R1209_U38;
  assign new_P2_R1209_U161 = ~P2_REG1_REG_15_ | ~new_P2_R1209_U160;
  assign new_P2_R1209_U162 = ~new_P2_U3433 | ~new_P2_R1209_U161;
  assign new_P2_R1209_U163 = ~new_P2_R1209_U38 | ~new_P2_R1209_U39;
  assign new_P2_R1209_U164 = ~new_P2_R1209_U98;
  assign new_P2_R1209_U165 = ~P2_REG1_REG_16_ | ~new_P2_R1209_U42;
  assign new_P2_R1209_U166 = ~new_P2_R1209_U165 | ~new_P2_R1209_U98;
  assign new_P2_R1209_U167 = ~new_P2_U3436 | ~new_P2_R1209_U41;
  assign new_P2_R1209_U168 = ~new_P2_R1209_U97;
  assign new_P2_R1209_U169 = ~P2_REG1_REG_17_ | ~new_P2_R1209_U44;
  assign new_P2_R1209_U170 = ~new_P2_R1209_U169 | ~new_P2_R1209_U97;
  assign new_P2_R1209_U171 = ~new_P2_U3439 | ~new_P2_R1209_U43;
  assign new_P2_R1209_U172 = ~new_P2_R1209_U47;
  assign new_P2_R1209_U173 = ~new_P2_U3442 | ~new_P2_R1209_U45;
  assign new_P2_R1209_U174 = ~new_P2_R1209_U172 | ~new_P2_R1209_U173;
  assign new_P2_R1209_U175 = ~P2_REG1_REG_18_ | ~new_P2_R1209_U46;
  assign new_P2_R1209_U176 = ~new_P2_R1209_U77 | ~new_P2_R1209_U174;
  assign new_P2_R1209_U177 = ~P2_REG1_REG_18_ | ~new_P2_R1209_U46;
  assign new_P2_R1209_U178 = ~new_P2_R1209_U177 | ~new_P2_R1209_U47;
  assign new_P2_R1209_U179 = ~new_P2_U3442 | ~new_P2_R1209_U45;
  assign new_P2_R1209_U180 = ~new_P2_R1209_U76 | ~new_P2_R1209_U178;
  assign new_P2_R1209_U181 = ~new_P2_U3386 | ~new_P2_R1209_U8;
  assign new_P2_R1209_U182 = ~P2_REG1_REG_9_ | ~new_P2_R1209_U27;
  assign new_P2_R1209_U183 = ~new_P2_U3415 | ~new_P2_R1209_U26;
  assign new_P2_R1209_U184 = ~new_P2_R1209_U67;
  assign new_P2_R1209_U185 = ~new_P2_R1209_U136 | ~new_P2_R1209_U184;
  assign new_P2_R1209_U186 = ~new_P2_R1209_U67 | ~new_P2_R1209_U87;
  assign new_P2_R1209_U187 = ~P2_REG1_REG_8_ | ~new_P2_R1209_U25;
  assign new_P2_R1209_U188 = ~new_P2_U3412 | ~new_P2_R1209_U24;
  assign new_P2_R1209_U189 = ~new_P2_R1209_U68;
  assign new_P2_R1209_U190 = ~new_P2_R1209_U132 | ~new_P2_R1209_U189;
  assign new_P2_R1209_U191 = ~new_P2_R1209_U68 | ~new_P2_R1209_U88;
  assign new_P2_R1209_U192 = ~P2_REG1_REG_7_ | ~new_P2_R1209_U23;
  assign new_P2_R1209_U193 = ~new_P2_U3409 | ~new_P2_R1209_U22;
  assign new_P2_R1209_U194 = ~new_P2_R1209_U69;
  assign new_P2_R1209_U195 = ~new_P2_R1209_U128 | ~new_P2_R1209_U194;
  assign new_P2_R1209_U196 = ~new_P2_R1209_U69 | ~new_P2_R1209_U89;
  assign new_P2_R1209_U197 = ~P2_REG1_REG_6_ | ~new_P2_R1209_U21;
  assign new_P2_R1209_U198 = ~new_P2_U3406 | ~new_P2_R1209_U20;
  assign new_P2_R1209_U199 = ~new_P2_R1209_U70;
  assign new_P2_R1209_U200 = ~new_P2_R1209_U124 | ~new_P2_R1209_U199;
  assign new_P2_R1209_U201 = ~new_P2_R1209_U70 | ~new_P2_R1209_U90;
  assign new_P2_R1209_U202 = ~P2_REG1_REG_5_ | ~new_P2_R1209_U19;
  assign new_P2_R1209_U203 = ~new_P2_U3403 | ~new_P2_R1209_U18;
  assign new_P2_R1209_U204 = ~new_P2_R1209_U71;
  assign new_P2_R1209_U205 = ~new_P2_R1209_U120 | ~new_P2_R1209_U204;
  assign new_P2_R1209_U206 = ~new_P2_R1209_U71 | ~new_P2_R1209_U91;
  assign new_P2_R1209_U207 = ~P2_REG1_REG_4_ | ~new_P2_R1209_U17;
  assign new_P2_R1209_U208 = ~new_P2_U3400 | ~new_P2_R1209_U16;
  assign new_P2_R1209_U209 = ~new_P2_R1209_U72;
  assign new_P2_R1209_U210 = ~new_P2_R1209_U116 | ~new_P2_R1209_U209;
  assign new_P2_R1209_U211 = ~new_P2_R1209_U72 | ~new_P2_R1209_U92;
  assign new_P2_R1209_U212 = ~P2_REG1_REG_3_ | ~new_P2_R1209_U15;
  assign new_P2_R1209_U213 = ~new_P2_U3397 | ~new_P2_R1209_U14;
  assign new_P2_R1209_U214 = ~new_P2_R1209_U73;
  assign new_P2_R1209_U215 = ~new_P2_R1209_U112 | ~new_P2_R1209_U214;
  assign new_P2_R1209_U216 = ~new_P2_R1209_U73 | ~new_P2_R1209_U93;
  assign new_P2_R1209_U217 = ~P2_REG1_REG_2_ | ~new_P2_R1209_U13;
  assign new_P2_R1209_U218 = ~new_P2_U3394 | ~new_P2_R1209_U12;
  assign new_P2_R1209_U219 = ~new_P2_R1209_U74;
  assign new_P2_R1209_U220 = ~new_P2_R1209_U108 | ~new_P2_R1209_U219;
  assign new_P2_R1209_U221 = ~new_P2_R1209_U74 | ~new_P2_R1209_U94;
  assign new_P2_R1209_U222 = ~new_P2_R1209_U104 | ~new_P2_R1209_U10;
  assign new_P2_R1209_U223 = ~P2_REG1_REG_1_ | ~new_P2_R1209_U9;
  assign new_P2_R1209_U224 = ~new_P2_R1209_U75;
  assign new_P2_R1209_U225 = ~new_P2_R1209_U224 | ~new_P2_U3391;
  assign new_P2_R1209_U226 = ~new_P2_R1209_U75 | ~new_P2_R1209_U11;
  assign new_P2_R1209_U227 = ~P2_REG1_REG_19_ | ~new_P2_R1209_U96;
  assign new_P2_R1209_U228 = ~new_P2_U3379 | ~new_P2_R1209_U95;
  assign new_P2_R1209_U229 = ~P2_REG1_REG_19_ | ~new_P2_R1209_U96;
  assign new_P2_R1209_U230 = ~new_P2_U3379 | ~new_P2_R1209_U95;
  assign new_P2_R1209_U231 = ~new_P2_R1209_U230 | ~new_P2_R1209_U229;
  assign new_P2_R1209_U232 = ~P2_REG1_REG_18_ | ~new_P2_R1209_U46;
  assign new_P2_R1209_U233 = ~new_P2_U3442 | ~new_P2_R1209_U45;
  assign new_P2_R1209_U234 = ~new_P2_R1209_U78;
  assign new_P2_R1209_U235 = ~new_P2_R1209_U234 | ~new_P2_R1209_U172;
  assign new_P2_R1209_U236 = ~new_P2_R1209_U78 | ~new_P2_R1209_U47;
  assign new_P2_R1209_U237 = ~P2_REG1_REG_17_ | ~new_P2_R1209_U44;
  assign new_P2_R1209_U238 = ~new_P2_U3439 | ~new_P2_R1209_U43;
  assign new_P2_R1209_U239 = ~new_P2_R1209_U79;
  assign new_P2_R1209_U240 = ~new_P2_R1209_U168 | ~new_P2_R1209_U239;
  assign new_P2_R1209_U241 = ~new_P2_R1209_U79 | ~new_P2_R1209_U97;
  assign new_P2_R1209_U242 = ~P2_REG1_REG_16_ | ~new_P2_R1209_U42;
  assign new_P2_R1209_U243 = ~new_P2_U3436 | ~new_P2_R1209_U41;
  assign new_P2_R1209_U244 = ~new_P2_R1209_U80;
  assign new_P2_R1209_U245 = ~new_P2_R1209_U164 | ~new_P2_R1209_U244;
  assign new_P2_R1209_U246 = ~new_P2_R1209_U80 | ~new_P2_R1209_U98;
  assign new_P2_R1209_U247 = ~new_P2_U3433 | ~new_P2_R1209_U39;
  assign new_P2_R1209_U248 = ~P2_REG1_REG_15_ | ~new_P2_R1209_U40;
  assign new_P2_R1209_U249 = ~new_P2_R1209_U81;
  assign new_P2_R1209_U250 = ~new_P2_R1209_U249 | ~new_P2_R1209_U160;
  assign new_P2_R1209_U251 = ~new_P2_R1209_U81 | ~new_P2_R1209_U38;
  assign new_P2_R1209_U252 = ~P2_REG1_REG_14_ | ~new_P2_R1209_U37;
  assign new_P2_R1209_U253 = ~new_P2_U3430 | ~new_P2_R1209_U36;
  assign new_P2_R1209_U254 = ~new_P2_R1209_U82;
  assign new_P2_R1209_U255 = ~new_P2_R1209_U156 | ~new_P2_R1209_U254;
  assign new_P2_R1209_U256 = ~new_P2_R1209_U82 | ~new_P2_R1209_U99;
  assign new_P2_R1209_U257 = ~P2_REG1_REG_13_ | ~new_P2_R1209_U35;
  assign new_P2_R1209_U258 = ~new_P2_U3427 | ~new_P2_R1209_U34;
  assign new_P2_R1209_U259 = ~new_P2_R1209_U83;
  assign new_P2_R1209_U260 = ~new_P2_R1209_U152 | ~new_P2_R1209_U259;
  assign new_P2_R1209_U261 = ~new_P2_R1209_U83 | ~new_P2_R1209_U100;
  assign new_P2_R1209_U262 = ~P2_REG1_REG_12_ | ~new_P2_R1209_U33;
  assign new_P2_R1209_U263 = ~new_P2_U3424 | ~new_P2_R1209_U32;
  assign new_P2_R1209_U264 = ~new_P2_R1209_U84;
  assign new_P2_R1209_U265 = ~new_P2_R1209_U148 | ~new_P2_R1209_U264;
  assign new_P2_R1209_U266 = ~new_P2_R1209_U84 | ~new_P2_R1209_U101;
  assign new_P2_R1209_U267 = ~P2_REG1_REG_11_ | ~new_P2_R1209_U31;
  assign new_P2_R1209_U268 = ~new_P2_U3421 | ~new_P2_R1209_U30;
  assign new_P2_R1209_U269 = ~new_P2_R1209_U85;
  assign new_P2_R1209_U270 = ~new_P2_R1209_U144 | ~new_P2_R1209_U269;
  assign new_P2_R1209_U271 = ~new_P2_R1209_U85 | ~new_P2_R1209_U102;
  assign new_P2_R1209_U272 = ~P2_REG1_REG_10_ | ~new_P2_R1209_U29;
  assign new_P2_R1209_U273 = ~new_P2_U3418 | ~new_P2_R1209_U28;
  assign new_P2_R1209_U274 = ~new_P2_R1209_U86;
  assign new_P2_R1209_U275 = ~new_P2_R1209_U140 | ~new_P2_R1209_U274;
  assign new_P2_R1209_U276 = ~new_P2_R1209_U86 | ~new_P2_R1209_U103;
  assign new_P2_R1300_U6 = ~new_P2_U3058;
  assign new_P2_R1300_U7 = ~new_P2_U3055;
  assign new_P2_R1300_U8 = new_P2_R1300_U10 & new_P2_R1300_U9;
  assign new_P2_R1300_U9 = ~new_P2_U3055 | ~new_P2_R1300_U6;
  assign new_P2_R1300_U10 = ~new_P2_U3058 | ~new_P2_R1300_U7;
  assign new_P2_R1200_U6 = new_P2_R1200_U212 & new_P2_R1200_U211;
  assign new_P2_R1200_U7 = new_P2_R1200_U246 & new_P2_R1200_U245;
  assign new_P2_R1200_U8 = new_P2_R1200_U193 & new_P2_R1200_U257;
  assign new_P2_R1200_U9 = new_P2_R1200_U259 & new_P2_R1200_U258;
  assign new_P2_R1200_U10 = new_P2_R1200_U194 & new_P2_R1200_U281;
  assign new_P2_R1200_U11 = new_P2_R1200_U283 & new_P2_R1200_U282;
  assign new_P2_R1200_U12 = new_P2_R1200_U299 & new_P2_R1200_U195;
  assign new_P2_R1200_U13 = new_P2_R1200_U215 & new_P2_R1200_U210 & new_P2_R1200_U197;
  assign new_P2_R1200_U14 = new_P2_R1200_U220 & new_P2_R1200_U198;
  assign new_P2_R1200_U15 = new_P2_R1200_U244 & new_P2_R1200_U224 & new_P2_R1200_U192;
  assign new_P2_R1200_U16 = new_P2_R1200_U399 & new_P2_R1200_U398;
  assign new_P2_R1200_U17 = ~new_P2_R1200_U331 | ~new_P2_R1200_U334;
  assign new_P2_R1200_U18 = ~new_P2_R1200_U322 | ~new_P2_R1200_U325;
  assign new_P2_R1200_U19 = ~new_P2_R1200_U311 | ~new_P2_R1200_U314;
  assign new_P2_R1200_U20 = ~new_P2_R1200_U305 | ~new_P2_R1200_U357;
  assign new_P2_R1200_U21 = ~new_P2_R1200_U137 | ~new_P2_R1200_U186;
  assign new_P2_R1200_U22 = ~new_P2_R1200_U242 | ~new_P2_R1200_U347;
  assign new_P2_R1200_U23 = ~new_P2_R1200_U235 | ~new_P2_R1200_U238;
  assign new_P2_R1200_U24 = ~new_P2_R1200_U227 | ~new_P2_R1200_U229;
  assign new_P2_R1200_U25 = ~new_P2_R1200_U175 | ~new_P2_R1200_U337;
  assign new_P2_R1200_U26 = ~new_P2_U3069;
  assign new_P2_R1200_U27 = ~new_P2_U3069 | ~new_P2_R1200_U32;
  assign new_P2_R1200_U28 = ~new_P2_U3083;
  assign new_P2_R1200_U29 = ~new_P2_U3404;
  assign new_P2_R1200_U30 = ~new_P2_U3407;
  assign new_P2_R1200_U31 = ~new_P2_U3401;
  assign new_P2_R1200_U32 = ~new_P2_U3410;
  assign new_P2_R1200_U33 = ~new_P2_U3413;
  assign new_P2_R1200_U34 = ~new_P2_U3067;
  assign new_P2_R1200_U35 = ~new_P2_U3067 | ~new_P2_R1200_U37;
  assign new_P2_R1200_U36 = ~new_P2_U3063;
  assign new_P2_R1200_U37 = ~new_P2_U3395;
  assign new_P2_R1200_U38 = ~new_P2_U3387;
  assign new_P2_R1200_U39 = ~new_P2_U3077;
  assign new_P2_R1200_U40 = ~new_P2_U3398;
  assign new_P2_R1200_U41 = ~new_P2_U3070;
  assign new_P2_R1200_U42 = ~new_P2_U3066;
  assign new_P2_R1200_U43 = ~new_P2_U3059;
  assign new_P2_R1200_U44 = ~new_P2_U3059 | ~new_P2_R1200_U31;
  assign new_P2_R1200_U45 = ~new_P2_R1200_U216 | ~new_P2_R1200_U214;
  assign new_P2_R1200_U46 = ~new_P2_U3416;
  assign new_P2_R1200_U47 = ~new_P2_U3082;
  assign new_P2_R1200_U48 = ~new_P2_R1200_U45 | ~new_P2_R1200_U217;
  assign new_P2_R1200_U49 = ~new_P2_R1200_U44 | ~new_P2_R1200_U231;
  assign new_P2_R1200_U50 = ~new_P2_R1200_U338 | ~new_P2_R1200_U204 | ~new_P2_R1200_U188;
  assign new_P2_R1200_U51 = ~new_P2_U3895;
  assign new_P2_R1200_U52 = ~new_P2_U3056;
  assign new_P2_R1200_U53 = ~new_P2_U3056 | ~new_P2_R1200_U90;
  assign new_P2_R1200_U54 = ~new_P2_U3052;
  assign new_P2_R1200_U55 = ~new_P2_U3071;
  assign new_P2_R1200_U56 = ~new_P2_U3062;
  assign new_P2_R1200_U57 = ~new_P2_U3061;
  assign new_P2_R1200_U58 = ~new_P2_U3419;
  assign new_P2_R1200_U59 = ~new_P2_U3082 | ~new_P2_R1200_U46;
  assign new_P2_R1200_U60 = ~new_P2_U3422;
  assign new_P2_R1200_U61 = ~new_P2_U3425;
  assign new_P2_R1200_U62 = ~new_P2_R1200_U249 | ~new_P2_R1200_U248;
  assign new_P2_R1200_U63 = ~new_P2_U3428;
  assign new_P2_R1200_U64 = ~new_P2_U3079;
  assign new_P2_R1200_U65 = ~new_P2_U3437;
  assign new_P2_R1200_U66 = ~new_P2_U3434;
  assign new_P2_R1200_U67 = ~new_P2_U3431;
  assign new_P2_R1200_U68 = ~new_P2_U3072;
  assign new_P2_R1200_U69 = ~new_P2_U3073;
  assign new_P2_R1200_U70 = ~new_P2_U3078;
  assign new_P2_R1200_U71 = ~new_P2_U3078 | ~new_P2_R1200_U67;
  assign new_P2_R1200_U72 = ~new_P2_U3440;
  assign new_P2_R1200_U73 = ~new_P2_U3068;
  assign new_P2_R1200_U74 = ~new_P2_U3081;
  assign new_P2_R1200_U75 = ~new_P2_U3445;
  assign new_P2_R1200_U76 = ~new_P2_U3080;
  assign new_P2_R1200_U77 = ~new_P2_U3903;
  assign new_P2_R1200_U78 = ~new_P2_U3075;
  assign new_P2_R1200_U79 = ~new_P2_U3900;
  assign new_P2_R1200_U80 = ~new_P2_U3901;
  assign new_P2_R1200_U81 = ~new_P2_U3902;
  assign new_P2_R1200_U82 = ~new_P2_U3065;
  assign new_P2_R1200_U83 = ~new_P2_U3060;
  assign new_P2_R1200_U84 = ~new_P2_U3074;
  assign new_P2_R1200_U85 = ~new_P2_U3074 | ~new_P2_R1200_U81;
  assign new_P2_R1200_U86 = ~new_P2_U3899;
  assign new_P2_R1200_U87 = ~new_P2_U3064;
  assign new_P2_R1200_U88 = ~new_P2_U3898;
  assign new_P2_R1200_U89 = ~new_P2_U3057;
  assign new_P2_R1200_U90 = ~new_P2_U3897;
  assign new_P2_R1200_U91 = ~new_P2_U3896;
  assign new_P2_R1200_U92 = ~new_P2_U3053;
  assign new_P2_R1200_U93 = ~new_P2_R1200_U297 | ~new_P2_R1200_U296;
  assign new_P2_R1200_U94 = ~new_P2_R1200_U85 | ~new_P2_R1200_U307;
  assign new_P2_R1200_U95 = ~new_P2_R1200_U71 | ~new_P2_R1200_U318;
  assign new_P2_R1200_U96 = ~new_P2_R1200_U349 | ~new_P2_R1200_U59;
  assign new_P2_R1200_U97 = ~new_P2_U3076;
  assign new_P2_R1200_U98 = ~new_P2_R1200_U406 | ~new_P2_R1200_U405;
  assign new_P2_R1200_U99 = ~new_P2_R1200_U420 | ~new_P2_R1200_U419;
  assign new_P2_R1200_U100 = ~new_P2_R1200_U425 | ~new_P2_R1200_U424;
  assign new_P2_R1200_U101 = ~new_P2_R1200_U441 | ~new_P2_R1200_U440;
  assign new_P2_R1200_U102 = ~new_P2_R1200_U446 | ~new_P2_R1200_U445;
  assign new_P2_R1200_U103 = ~new_P2_R1200_U451 | ~new_P2_R1200_U450;
  assign new_P2_R1200_U104 = ~new_P2_R1200_U456 | ~new_P2_R1200_U455;
  assign new_P2_R1200_U105 = ~new_P2_R1200_U461 | ~new_P2_R1200_U460;
  assign new_P2_R1200_U106 = ~new_P2_R1200_U477 | ~new_P2_R1200_U476;
  assign new_P2_R1200_U107 = ~new_P2_R1200_U482 | ~new_P2_R1200_U481;
  assign new_P2_R1200_U108 = ~new_P2_R1200_U365 | ~new_P2_R1200_U364;
  assign new_P2_R1200_U109 = ~new_P2_R1200_U374 | ~new_P2_R1200_U373;
  assign new_P2_R1200_U110 = ~new_P2_R1200_U381 | ~new_P2_R1200_U380;
  assign new_P2_R1200_U111 = ~new_P2_R1200_U385 | ~new_P2_R1200_U384;
  assign new_P2_R1200_U112 = ~new_P2_R1200_U394 | ~new_P2_R1200_U393;
  assign new_P2_R1200_U113 = ~new_P2_R1200_U415 | ~new_P2_R1200_U414;
  assign new_P2_R1200_U114 = ~new_P2_R1200_U432 | ~new_P2_R1200_U431;
  assign new_P2_R1200_U115 = ~new_P2_R1200_U436 | ~new_P2_R1200_U435;
  assign new_P2_R1200_U116 = ~new_P2_R1200_U468 | ~new_P2_R1200_U467;
  assign new_P2_R1200_U117 = ~new_P2_R1200_U472 | ~new_P2_R1200_U471;
  assign new_P2_R1200_U118 = ~new_P2_R1200_U489 | ~new_P2_R1200_U488;
  assign new_P2_R1200_U119 = new_P2_R1200_U206 & new_P2_R1200_U196;
  assign new_P2_R1200_U120 = new_P2_R1200_U209 & new_P2_R1200_U208;
  assign new_P2_R1200_U121 = new_P2_R1200_U14 & new_P2_R1200_U13;
  assign new_P2_R1200_U122 = new_P2_R1200_U340 & new_P2_R1200_U222;
  assign new_P2_R1200_U123 = new_P2_R1200_U342 & new_P2_R1200_U122;
  assign new_P2_R1200_U124 = new_P2_R1200_U27 & new_P2_R1200_U367 & new_P2_R1200_U366;
  assign new_P2_R1200_U125 = new_P2_R1200_U370 & new_P2_R1200_U198;
  assign new_P2_R1200_U126 = new_P2_R1200_U237 & new_P2_R1200_U6;
  assign new_P2_R1200_U127 = new_P2_R1200_U377 & new_P2_R1200_U197;
  assign new_P2_R1200_U128 = new_P2_R1200_U35 & new_P2_R1200_U387 & new_P2_R1200_U386;
  assign new_P2_R1200_U129 = new_P2_R1200_U390 & new_P2_R1200_U196;
  assign new_P2_R1200_U130 = new_P2_R1200_U251 & new_P2_R1200_U15;
  assign new_P2_R1200_U131 = new_P2_R1200_U343 & new_P2_R1200_U252;
  assign new_P2_R1200_U132 = new_P2_R1200_U262 & new_P2_R1200_U8;
  assign new_P2_R1200_U133 = new_P2_R1200_U286 & new_P2_R1200_U10;
  assign new_P2_R1200_U134 = new_P2_R1200_U302 & new_P2_R1200_U301;
  assign new_P2_R1200_U135 = new_P2_R1200_U397 & new_P2_R1200_U303;
  assign new_P2_R1200_U136 = new_P2_R1200_U16 & new_P2_R1200_U304 & new_P2_R1200_U302 & new_P2_R1200_U301;
  assign new_P2_R1200_U137 = new_P2_R1200_U359 & new_P2_R1200_U165;
  assign new_P2_R1200_U138 = ~new_P2_R1200_U403 | ~new_P2_R1200_U402;
  assign new_P2_R1200_U139 = new_P2_R1200_U53 & new_P2_R1200_U408 & new_P2_R1200_U407;
  assign new_P2_R1200_U140 = new_P2_R1200_U411 & new_P2_R1200_U195;
  assign new_P2_R1200_U141 = ~new_P2_R1200_U417 | ~new_P2_R1200_U416;
  assign new_P2_R1200_U142 = ~new_P2_R1200_U422 | ~new_P2_R1200_U421;
  assign new_P2_R1200_U143 = new_P2_R1200_U313 & new_P2_R1200_U11;
  assign new_P2_R1200_U144 = new_P2_R1200_U428 & new_P2_R1200_U194;
  assign new_P2_R1200_U145 = ~new_P2_R1200_U438 | ~new_P2_R1200_U437;
  assign new_P2_R1200_U146 = ~new_P2_R1200_U443 | ~new_P2_R1200_U442;
  assign new_P2_R1200_U147 = ~new_P2_R1200_U448 | ~new_P2_R1200_U447;
  assign new_P2_R1200_U148 = ~new_P2_R1200_U453 | ~new_P2_R1200_U452;
  assign new_P2_R1200_U149 = ~new_P2_R1200_U458 | ~new_P2_R1200_U457;
  assign new_P2_R1200_U150 = new_P2_R1200_U324 & new_P2_R1200_U9;
  assign new_P2_R1200_U151 = new_P2_R1200_U464 & new_P2_R1200_U193;
  assign new_P2_R1200_U152 = ~new_P2_R1200_U474 | ~new_P2_R1200_U473;
  assign new_P2_R1200_U153 = ~new_P2_R1200_U479 | ~new_P2_R1200_U478;
  assign new_P2_R1200_U154 = new_P2_R1200_U333 & new_P2_R1200_U7;
  assign new_P2_R1200_U155 = new_P2_R1200_U485 & new_P2_R1200_U192;
  assign new_P2_R1200_U156 = new_P2_R1200_U363 & new_P2_R1200_U362;
  assign new_P2_R1200_U157 = ~new_P2_R1200_U123 | ~new_P2_R1200_U341;
  assign new_P2_R1200_U158 = new_P2_R1200_U372 & new_P2_R1200_U371;
  assign new_P2_R1200_U159 = new_P2_R1200_U379 & new_P2_R1200_U378;
  assign new_P2_R1200_U160 = new_P2_R1200_U383 & new_P2_R1200_U382;
  assign new_P2_R1200_U161 = ~new_P2_R1200_U120 | ~new_P2_R1200_U344;
  assign new_P2_R1200_U162 = new_P2_R1200_U392 & new_P2_R1200_U391;
  assign new_P2_R1200_U163 = ~new_P2_U3904;
  assign new_P2_R1200_U164 = ~new_P2_U3054;
  assign new_P2_R1200_U165 = new_P2_R1200_U401 & new_P2_R1200_U400;
  assign new_P2_R1200_U166 = ~new_P2_R1200_U134 | ~new_P2_R1200_U360;
  assign new_P2_R1200_U167 = new_P2_R1200_U413 & new_P2_R1200_U412;
  assign new_P2_R1200_U168 = ~new_P2_R1200_U293 | ~new_P2_R1200_U292;
  assign new_P2_R1200_U169 = ~new_P2_R1200_U289 | ~new_P2_R1200_U288;
  assign new_P2_R1200_U170 = new_P2_R1200_U430 & new_P2_R1200_U429;
  assign new_P2_R1200_U171 = new_P2_R1200_U434 & new_P2_R1200_U433;
  assign new_P2_R1200_U172 = ~new_P2_R1200_U279 | ~new_P2_R1200_U278;
  assign new_P2_R1200_U173 = ~new_P2_R1200_U275 | ~new_P2_R1200_U274;
  assign new_P2_R1200_U174 = ~new_P2_U3392;
  assign new_P2_R1200_U175 = ~new_P2_U3387 | ~new_P2_R1200_U97;
  assign new_P2_R1200_U176 = ~new_P2_R1200_U339 | ~new_P2_R1200_U271 | ~new_P2_R1200_U187;
  assign new_P2_R1200_U177 = ~new_P2_U3443;
  assign new_P2_R1200_U178 = ~new_P2_R1200_U269 | ~new_P2_R1200_U268;
  assign new_P2_R1200_U179 = ~new_P2_R1200_U265 | ~new_P2_R1200_U264;
  assign new_P2_R1200_U180 = new_P2_R1200_U466 & new_P2_R1200_U465;
  assign new_P2_R1200_U181 = new_P2_R1200_U470 & new_P2_R1200_U469;
  assign new_P2_R1200_U182 = ~new_P2_R1200_U255 | ~new_P2_R1200_U254;
  assign new_P2_R1200_U183 = ~new_P2_R1200_U131 | ~new_P2_R1200_U353;
  assign new_P2_R1200_U184 = ~new_P2_R1200_U351 | ~new_P2_R1200_U62;
  assign new_P2_R1200_U185 = new_P2_R1200_U487 & new_P2_R1200_U486;
  assign new_P2_R1200_U186 = ~new_P2_R1200_U135 | ~new_P2_R1200_U166;
  assign new_P2_R1200_U187 = ~new_P2_R1200_U178 | ~new_P2_R1200_U177;
  assign new_P2_R1200_U188 = ~new_P2_R1200_U175 | ~new_P2_R1200_U174;
  assign new_P2_R1200_U189 = ~new_P2_R1200_U53;
  assign new_P2_R1200_U190 = ~new_P2_R1200_U35;
  assign new_P2_R1200_U191 = ~new_P2_R1200_U27;
  assign new_P2_R1200_U192 = ~new_P2_U3419 | ~new_P2_R1200_U57;
  assign new_P2_R1200_U193 = ~new_P2_U3434 | ~new_P2_R1200_U69;
  assign new_P2_R1200_U194 = ~new_P2_U3901 | ~new_P2_R1200_U83;
  assign new_P2_R1200_U195 = ~new_P2_U3897 | ~new_P2_R1200_U52;
  assign new_P2_R1200_U196 = ~new_P2_U3395 | ~new_P2_R1200_U34;
  assign new_P2_R1200_U197 = ~new_P2_U3404 | ~new_P2_R1200_U42;
  assign new_P2_R1200_U198 = ~new_P2_U3410 | ~new_P2_R1200_U26;
  assign new_P2_R1200_U199 = ~new_P2_R1200_U71;
  assign new_P2_R1200_U200 = ~new_P2_R1200_U85;
  assign new_P2_R1200_U201 = ~new_P2_R1200_U44;
  assign new_P2_R1200_U202 = ~new_P2_R1200_U59;
  assign new_P2_R1200_U203 = ~new_P2_R1200_U175;
  assign new_P2_R1200_U204 = ~new_P2_U3077 | ~new_P2_R1200_U175;
  assign new_P2_R1200_U205 = ~new_P2_R1200_U50;
  assign new_P2_R1200_U206 = ~new_P2_U3398 | ~new_P2_R1200_U36;
  assign new_P2_R1200_U207 = ~new_P2_R1200_U36 | ~new_P2_R1200_U35;
  assign new_P2_R1200_U208 = ~new_P2_R1200_U207 | ~new_P2_R1200_U40;
  assign new_P2_R1200_U209 = ~new_P2_U3063 | ~new_P2_R1200_U190;
  assign new_P2_R1200_U210 = ~new_P2_U3407 | ~new_P2_R1200_U41;
  assign new_P2_R1200_U211 = ~new_P2_U3070 | ~new_P2_R1200_U30;
  assign new_P2_R1200_U212 = ~new_P2_U3066 | ~new_P2_R1200_U29;
  assign new_P2_R1200_U213 = ~new_P2_R1200_U201 | ~new_P2_R1200_U197;
  assign new_P2_R1200_U214 = ~new_P2_R1200_U6 | ~new_P2_R1200_U213;
  assign new_P2_R1200_U215 = ~new_P2_U3401 | ~new_P2_R1200_U43;
  assign new_P2_R1200_U216 = ~new_P2_U3407 | ~new_P2_R1200_U41;
  assign new_P2_R1200_U217 = ~new_P2_R1200_U13 | ~new_P2_R1200_U161;
  assign new_P2_R1200_U218 = ~new_P2_R1200_U45;
  assign new_P2_R1200_U219 = ~new_P2_R1200_U48;
  assign new_P2_R1200_U220 = ~new_P2_U3413 | ~new_P2_R1200_U28;
  assign new_P2_R1200_U221 = ~new_P2_R1200_U28 | ~new_P2_R1200_U27;
  assign new_P2_R1200_U222 = ~new_P2_U3083 | ~new_P2_R1200_U191;
  assign new_P2_R1200_U223 = ~new_P2_R1200_U157;
  assign new_P2_R1200_U224 = ~new_P2_U3416 | ~new_P2_R1200_U47;
  assign new_P2_R1200_U225 = ~new_P2_R1200_U224 | ~new_P2_R1200_U59;
  assign new_P2_R1200_U226 = ~new_P2_R1200_U219 | ~new_P2_R1200_U27;
  assign new_P2_R1200_U227 = ~new_P2_R1200_U125 | ~new_P2_R1200_U226;
  assign new_P2_R1200_U228 = ~new_P2_R1200_U48 | ~new_P2_R1200_U198;
  assign new_P2_R1200_U229 = ~new_P2_R1200_U124 | ~new_P2_R1200_U228;
  assign new_P2_R1200_U230 = ~new_P2_R1200_U27 | ~new_P2_R1200_U198;
  assign new_P2_R1200_U231 = ~new_P2_R1200_U215 | ~new_P2_R1200_U161;
  assign new_P2_R1200_U232 = ~new_P2_R1200_U49;
  assign new_P2_R1200_U233 = ~new_P2_U3066 | ~new_P2_R1200_U29;
  assign new_P2_R1200_U234 = ~new_P2_R1200_U232 | ~new_P2_R1200_U233;
  assign new_P2_R1200_U235 = ~new_P2_R1200_U127 | ~new_P2_R1200_U234;
  assign new_P2_R1200_U236 = ~new_P2_R1200_U49 | ~new_P2_R1200_U197;
  assign new_P2_R1200_U237 = ~new_P2_U3407 | ~new_P2_R1200_U41;
  assign new_P2_R1200_U238 = ~new_P2_R1200_U126 | ~new_P2_R1200_U236;
  assign new_P2_R1200_U239 = ~new_P2_U3066 | ~new_P2_R1200_U29;
  assign new_P2_R1200_U240 = ~new_P2_R1200_U239 | ~new_P2_R1200_U197;
  assign new_P2_R1200_U241 = ~new_P2_R1200_U215 | ~new_P2_R1200_U44;
  assign new_P2_R1200_U242 = ~new_P2_R1200_U129 | ~new_P2_R1200_U348;
  assign new_P2_R1200_U243 = ~new_P2_R1200_U35 | ~new_P2_R1200_U196;
  assign new_P2_R1200_U244 = ~new_P2_U3422 | ~new_P2_R1200_U56;
  assign new_P2_R1200_U245 = ~new_P2_U3062 | ~new_P2_R1200_U60;
  assign new_P2_R1200_U246 = ~new_P2_U3061 | ~new_P2_R1200_U58;
  assign new_P2_R1200_U247 = ~new_P2_R1200_U202 | ~new_P2_R1200_U192;
  assign new_P2_R1200_U248 = ~new_P2_R1200_U7 | ~new_P2_R1200_U247;
  assign new_P2_R1200_U249 = ~new_P2_U3422 | ~new_P2_R1200_U56;
  assign new_P2_R1200_U250 = ~new_P2_R1200_U62;
  assign new_P2_R1200_U251 = ~new_P2_U3425 | ~new_P2_R1200_U55;
  assign new_P2_R1200_U252 = ~new_P2_U3071 | ~new_P2_R1200_U61;
  assign new_P2_R1200_U253 = ~new_P2_U3428 | ~new_P2_R1200_U64;
  assign new_P2_R1200_U254 = ~new_P2_R1200_U253 | ~new_P2_R1200_U183;
  assign new_P2_R1200_U255 = ~new_P2_U3079 | ~new_P2_R1200_U63;
  assign new_P2_R1200_U256 = ~new_P2_R1200_U182;
  assign new_P2_R1200_U257 = ~new_P2_U3437 | ~new_P2_R1200_U68;
  assign new_P2_R1200_U258 = ~new_P2_U3072 | ~new_P2_R1200_U65;
  assign new_P2_R1200_U259 = ~new_P2_U3073 | ~new_P2_R1200_U66;
  assign new_P2_R1200_U260 = ~new_P2_R1200_U199 | ~new_P2_R1200_U8;
  assign new_P2_R1200_U261 = ~new_P2_R1200_U9 | ~new_P2_R1200_U260;
  assign new_P2_R1200_U262 = ~new_P2_U3431 | ~new_P2_R1200_U70;
  assign new_P2_R1200_U263 = ~new_P2_U3437 | ~new_P2_R1200_U68;
  assign new_P2_R1200_U264 = ~new_P2_R1200_U132 | ~new_P2_R1200_U182;
  assign new_P2_R1200_U265 = ~new_P2_R1200_U263 | ~new_P2_R1200_U261;
  assign new_P2_R1200_U266 = ~new_P2_R1200_U179;
  assign new_P2_R1200_U267 = ~new_P2_U3440 | ~new_P2_R1200_U73;
  assign new_P2_R1200_U268 = ~new_P2_R1200_U267 | ~new_P2_R1200_U179;
  assign new_P2_R1200_U269 = ~new_P2_U3068 | ~new_P2_R1200_U72;
  assign new_P2_R1200_U270 = ~new_P2_R1200_U178;
  assign new_P2_R1200_U271 = ~new_P2_U3081 | ~new_P2_R1200_U178;
  assign new_P2_R1200_U272 = ~new_P2_R1200_U176;
  assign new_P2_R1200_U273 = ~new_P2_U3445 | ~new_P2_R1200_U76;
  assign new_P2_R1200_U274 = ~new_P2_R1200_U273 | ~new_P2_R1200_U176;
  assign new_P2_R1200_U275 = ~new_P2_U3080 | ~new_P2_R1200_U75;
  assign new_P2_R1200_U276 = ~new_P2_R1200_U173;
  assign new_P2_R1200_U277 = ~new_P2_U3903 | ~new_P2_R1200_U78;
  assign new_P2_R1200_U278 = ~new_P2_R1200_U277 | ~new_P2_R1200_U173;
  assign new_P2_R1200_U279 = ~new_P2_U3075 | ~new_P2_R1200_U77;
  assign new_P2_R1200_U280 = ~new_P2_R1200_U172;
  assign new_P2_R1200_U281 = ~new_P2_U3900 | ~new_P2_R1200_U82;
  assign new_P2_R1200_U282 = ~new_P2_U3065 | ~new_P2_R1200_U79;
  assign new_P2_R1200_U283 = ~new_P2_U3060 | ~new_P2_R1200_U80;
  assign new_P2_R1200_U284 = ~new_P2_R1200_U200 | ~new_P2_R1200_U10;
  assign new_P2_R1200_U285 = ~new_P2_R1200_U11 | ~new_P2_R1200_U284;
  assign new_P2_R1200_U286 = ~new_P2_U3902 | ~new_P2_R1200_U84;
  assign new_P2_R1200_U287 = ~new_P2_U3900 | ~new_P2_R1200_U82;
  assign new_P2_R1200_U288 = ~new_P2_R1200_U133 | ~new_P2_R1200_U172;
  assign new_P2_R1200_U289 = ~new_P2_R1200_U287 | ~new_P2_R1200_U285;
  assign new_P2_R1200_U290 = ~new_P2_R1200_U169;
  assign new_P2_R1200_U291 = ~new_P2_U3899 | ~new_P2_R1200_U87;
  assign new_P2_R1200_U292 = ~new_P2_R1200_U291 | ~new_P2_R1200_U169;
  assign new_P2_R1200_U293 = ~new_P2_U3064 | ~new_P2_R1200_U86;
  assign new_P2_R1200_U294 = ~new_P2_R1200_U168;
  assign new_P2_R1200_U295 = ~new_P2_U3898 | ~new_P2_R1200_U89;
  assign new_P2_R1200_U296 = ~new_P2_R1200_U295 | ~new_P2_R1200_U168;
  assign new_P2_R1200_U297 = ~new_P2_U3057 | ~new_P2_R1200_U88;
  assign new_P2_R1200_U298 = ~new_P2_R1200_U93;
  assign new_P2_R1200_U299 = ~new_P2_U3896 | ~new_P2_R1200_U54;
  assign new_P2_R1200_U300 = ~new_P2_R1200_U54 | ~new_P2_R1200_U53;
  assign new_P2_R1200_U301 = ~new_P2_R1200_U300 | ~new_P2_R1200_U91;
  assign new_P2_R1200_U302 = ~new_P2_U3052 | ~new_P2_R1200_U189;
  assign new_P2_R1200_U303 = ~new_P2_U3895 | ~new_P2_R1200_U92;
  assign new_P2_R1200_U304 = ~new_P2_U3053 | ~new_P2_R1200_U51;
  assign new_P2_R1200_U305 = ~new_P2_R1200_U140 | ~new_P2_R1200_U355;
  assign new_P2_R1200_U306 = ~new_P2_R1200_U53 | ~new_P2_R1200_U195;
  assign new_P2_R1200_U307 = ~new_P2_R1200_U286 | ~new_P2_R1200_U172;
  assign new_P2_R1200_U308 = ~new_P2_R1200_U94;
  assign new_P2_R1200_U309 = ~new_P2_U3060 | ~new_P2_R1200_U80;
  assign new_P2_R1200_U310 = ~new_P2_R1200_U308 | ~new_P2_R1200_U309;
  assign new_P2_R1200_U311 = ~new_P2_R1200_U144 | ~new_P2_R1200_U310;
  assign new_P2_R1200_U312 = ~new_P2_R1200_U94 | ~new_P2_R1200_U194;
  assign new_P2_R1200_U313 = ~new_P2_U3900 | ~new_P2_R1200_U82;
  assign new_P2_R1200_U314 = ~new_P2_R1200_U143 | ~new_P2_R1200_U312;
  assign new_P2_R1200_U315 = ~new_P2_U3060 | ~new_P2_R1200_U80;
  assign new_P2_R1200_U316 = ~new_P2_R1200_U194 | ~new_P2_R1200_U315;
  assign new_P2_R1200_U317 = ~new_P2_R1200_U286 | ~new_P2_R1200_U85;
  assign new_P2_R1200_U318 = ~new_P2_R1200_U262 | ~new_P2_R1200_U182;
  assign new_P2_R1200_U319 = ~new_P2_R1200_U95;
  assign new_P2_R1200_U320 = ~new_P2_U3073 | ~new_P2_R1200_U66;
  assign new_P2_R1200_U321 = ~new_P2_R1200_U319 | ~new_P2_R1200_U320;
  assign new_P2_R1200_U322 = ~new_P2_R1200_U151 | ~new_P2_R1200_U321;
  assign new_P2_R1200_U323 = ~new_P2_R1200_U95 | ~new_P2_R1200_U193;
  assign new_P2_R1200_U324 = ~new_P2_U3437 | ~new_P2_R1200_U68;
  assign new_P2_R1200_U325 = ~new_P2_R1200_U150 | ~new_P2_R1200_U323;
  assign new_P2_R1200_U326 = ~new_P2_U3073 | ~new_P2_R1200_U66;
  assign new_P2_R1200_U327 = ~new_P2_R1200_U193 | ~new_P2_R1200_U326;
  assign new_P2_R1200_U328 = ~new_P2_R1200_U262 | ~new_P2_R1200_U71;
  assign new_P2_R1200_U329 = ~new_P2_U3061 | ~new_P2_R1200_U58;
  assign new_P2_R1200_U330 = ~new_P2_R1200_U350 | ~new_P2_R1200_U329;
  assign new_P2_R1200_U331 = ~new_P2_R1200_U155 | ~new_P2_R1200_U330;
  assign new_P2_R1200_U332 = ~new_P2_R1200_U96 | ~new_P2_R1200_U192;
  assign new_P2_R1200_U333 = ~new_P2_U3422 | ~new_P2_R1200_U56;
  assign new_P2_R1200_U334 = ~new_P2_R1200_U154 | ~new_P2_R1200_U332;
  assign new_P2_R1200_U335 = ~new_P2_U3061 | ~new_P2_R1200_U58;
  assign new_P2_R1200_U336 = ~new_P2_R1200_U192 | ~new_P2_R1200_U335;
  assign new_P2_R1200_U337 = ~new_P2_U3076 | ~new_P2_R1200_U38;
  assign new_P2_R1200_U338 = ~new_P2_U3077 | ~new_P2_R1200_U174;
  assign new_P2_R1200_U339 = ~new_P2_U3081 | ~new_P2_R1200_U177;
  assign new_P2_R1200_U340 = ~new_P2_R1200_U33 | ~new_P2_R1200_U221;
  assign new_P2_R1200_U341 = ~new_P2_R1200_U121 | ~new_P2_R1200_U161;
  assign new_P2_R1200_U342 = ~new_P2_R1200_U218 | ~new_P2_R1200_U14;
  assign new_P2_R1200_U343 = ~new_P2_R1200_U250 | ~new_P2_R1200_U251;
  assign new_P2_R1200_U344 = ~new_P2_R1200_U119 | ~new_P2_R1200_U50;
  assign new_P2_R1200_U345 = ~new_P2_R1200_U161;
  assign new_P2_R1200_U346 = ~new_P2_R1200_U196 | ~new_P2_R1200_U50;
  assign new_P2_R1200_U347 = ~new_P2_R1200_U128 | ~new_P2_R1200_U346;
  assign new_P2_R1200_U348 = ~new_P2_R1200_U205 | ~new_P2_R1200_U35;
  assign new_P2_R1200_U349 = ~new_P2_R1200_U224 | ~new_P2_R1200_U157;
  assign new_P2_R1200_U350 = ~new_P2_R1200_U96;
  assign new_P2_R1200_U351 = ~new_P2_R1200_U15 | ~new_P2_R1200_U157;
  assign new_P2_R1200_U352 = ~new_P2_R1200_U184;
  assign new_P2_R1200_U353 = ~new_P2_R1200_U130 | ~new_P2_R1200_U157;
  assign new_P2_R1200_U354 = ~new_P2_R1200_U183;
  assign new_P2_R1200_U355 = ~new_P2_R1200_U298 | ~new_P2_R1200_U53;
  assign new_P2_R1200_U356 = ~new_P2_R1200_U195 | ~new_P2_R1200_U93;
  assign new_P2_R1200_U357 = ~new_P2_R1200_U139 | ~new_P2_R1200_U356;
  assign new_P2_R1200_U358 = ~new_P2_R1200_U12 | ~new_P2_R1200_U93;
  assign new_P2_R1200_U359 = ~new_P2_R1200_U136 | ~new_P2_R1200_U358;
  assign new_P2_R1200_U360 = ~new_P2_R1200_U12 | ~new_P2_R1200_U93;
  assign new_P2_R1200_U361 = ~new_P2_R1200_U166;
  assign new_P2_R1200_U362 = ~new_P2_U3416 | ~new_P2_R1200_U47;
  assign new_P2_R1200_U363 = ~new_P2_U3082 | ~new_P2_R1200_U46;
  assign new_P2_R1200_U364 = ~new_P2_R1200_U225 | ~new_P2_R1200_U157;
  assign new_P2_R1200_U365 = ~new_P2_R1200_U223 | ~new_P2_R1200_U156;
  assign new_P2_R1200_U366 = ~new_P2_U3413 | ~new_P2_R1200_U28;
  assign new_P2_R1200_U367 = ~new_P2_U3083 | ~new_P2_R1200_U33;
  assign new_P2_R1200_U368 = ~new_P2_U3413 | ~new_P2_R1200_U28;
  assign new_P2_R1200_U369 = ~new_P2_U3083 | ~new_P2_R1200_U33;
  assign new_P2_R1200_U370 = ~new_P2_R1200_U369 | ~new_P2_R1200_U368;
  assign new_P2_R1200_U371 = ~new_P2_U3410 | ~new_P2_R1200_U26;
  assign new_P2_R1200_U372 = ~new_P2_U3069 | ~new_P2_R1200_U32;
  assign new_P2_R1200_U373 = ~new_P2_R1200_U230 | ~new_P2_R1200_U48;
  assign new_P2_R1200_U374 = ~new_P2_R1200_U158 | ~new_P2_R1200_U219;
  assign new_P2_R1200_U375 = ~new_P2_U3407 | ~new_P2_R1200_U41;
  assign new_P2_R1200_U376 = ~new_P2_U3070 | ~new_P2_R1200_U30;
  assign new_P2_R1200_U377 = ~new_P2_R1200_U376 | ~new_P2_R1200_U375;
  assign new_P2_R1200_U378 = ~new_P2_U3404 | ~new_P2_R1200_U42;
  assign new_P2_R1200_U379 = ~new_P2_U3066 | ~new_P2_R1200_U29;
  assign new_P2_R1200_U380 = ~new_P2_R1200_U240 | ~new_P2_R1200_U49;
  assign new_P2_R1200_U381 = ~new_P2_R1200_U159 | ~new_P2_R1200_U232;
  assign new_P2_R1200_U382 = ~new_P2_U3401 | ~new_P2_R1200_U43;
  assign new_P2_R1200_U383 = ~new_P2_U3059 | ~new_P2_R1200_U31;
  assign new_P2_R1200_U384 = ~new_P2_R1200_U161 | ~new_P2_R1200_U241;
  assign new_P2_R1200_U385 = ~new_P2_R1200_U345 | ~new_P2_R1200_U160;
  assign new_P2_R1200_U386 = ~new_P2_U3398 | ~new_P2_R1200_U36;
  assign new_P2_R1200_U387 = ~new_P2_U3063 | ~new_P2_R1200_U40;
  assign new_P2_R1200_U388 = ~new_P2_U3398 | ~new_P2_R1200_U36;
  assign new_P2_R1200_U389 = ~new_P2_U3063 | ~new_P2_R1200_U40;
  assign new_P2_R1200_U390 = ~new_P2_R1200_U389 | ~new_P2_R1200_U388;
  assign new_P2_R1200_U391 = ~new_P2_U3395 | ~new_P2_R1200_U34;
  assign new_P2_R1200_U392 = ~new_P2_U3067 | ~new_P2_R1200_U37;
  assign new_P2_R1200_U393 = ~new_P2_R1200_U243 | ~new_P2_R1200_U50;
  assign new_P2_R1200_U394 = ~new_P2_R1200_U162 | ~new_P2_R1200_U205;
  assign new_P2_R1200_U395 = ~new_P2_U3904 | ~new_P2_R1200_U164;
  assign new_P2_R1200_U396 = ~new_P2_U3054 | ~new_P2_R1200_U163;
  assign new_P2_R1200_U397 = ~new_P2_R1200_U396 | ~new_P2_R1200_U395;
  assign new_P2_R1200_U398 = ~new_P2_U3904 | ~new_P2_R1200_U164;
  assign new_P2_R1200_U399 = ~new_P2_U3054 | ~new_P2_R1200_U163;
  assign new_P2_R1200_U400 = ~new_P2_R1200_U51 | ~new_P2_U3053 | ~new_P2_R1200_U397;
  assign new_P2_R1200_U401 = ~new_P2_U3895 | ~new_P2_R1200_U16 | ~new_P2_R1200_U92;
  assign new_P2_R1200_U402 = ~new_P2_U3895 | ~new_P2_R1200_U92;
  assign new_P2_R1200_U403 = ~new_P2_U3053 | ~new_P2_R1200_U51;
  assign new_P2_R1200_U404 = ~new_P2_R1200_U138;
  assign new_P2_R1200_U405 = ~new_P2_R1200_U361 | ~new_P2_R1200_U404;
  assign new_P2_R1200_U406 = ~new_P2_R1200_U138 | ~new_P2_R1200_U166;
  assign new_P2_R1200_U407 = ~new_P2_U3896 | ~new_P2_R1200_U54;
  assign new_P2_R1200_U408 = ~new_P2_U3052 | ~new_P2_R1200_U91;
  assign new_P2_R1200_U409 = ~new_P2_U3896 | ~new_P2_R1200_U54;
  assign new_P2_R1200_U410 = ~new_P2_U3052 | ~new_P2_R1200_U91;
  assign new_P2_R1200_U411 = ~new_P2_R1200_U410 | ~new_P2_R1200_U409;
  assign new_P2_R1200_U412 = ~new_P2_U3897 | ~new_P2_R1200_U52;
  assign new_P2_R1200_U413 = ~new_P2_U3056 | ~new_P2_R1200_U90;
  assign new_P2_R1200_U414 = ~new_P2_R1200_U306 | ~new_P2_R1200_U93;
  assign new_P2_R1200_U415 = ~new_P2_R1200_U167 | ~new_P2_R1200_U298;
  assign new_P2_R1200_U416 = ~new_P2_U3898 | ~new_P2_R1200_U89;
  assign new_P2_R1200_U417 = ~new_P2_U3057 | ~new_P2_R1200_U88;
  assign new_P2_R1200_U418 = ~new_P2_R1200_U141;
  assign new_P2_R1200_U419 = ~new_P2_R1200_U294 | ~new_P2_R1200_U418;
  assign new_P2_R1200_U420 = ~new_P2_R1200_U141 | ~new_P2_R1200_U168;
  assign new_P2_R1200_U421 = ~new_P2_U3899 | ~new_P2_R1200_U87;
  assign new_P2_R1200_U422 = ~new_P2_U3064 | ~new_P2_R1200_U86;
  assign new_P2_R1200_U423 = ~new_P2_R1200_U142;
  assign new_P2_R1200_U424 = ~new_P2_R1200_U290 | ~new_P2_R1200_U423;
  assign new_P2_R1200_U425 = ~new_P2_R1200_U142 | ~new_P2_R1200_U169;
  assign new_P2_R1200_U426 = ~new_P2_U3900 | ~new_P2_R1200_U82;
  assign new_P2_R1200_U427 = ~new_P2_U3065 | ~new_P2_R1200_U79;
  assign new_P2_R1200_U428 = ~new_P2_R1200_U427 | ~new_P2_R1200_U426;
  assign new_P2_R1200_U429 = ~new_P2_U3901 | ~new_P2_R1200_U83;
  assign new_P2_R1200_U430 = ~new_P2_U3060 | ~new_P2_R1200_U80;
  assign new_P2_R1200_U431 = ~new_P2_R1200_U316 | ~new_P2_R1200_U94;
  assign new_P2_R1200_U432 = ~new_P2_R1200_U170 | ~new_P2_R1200_U308;
  assign new_P2_R1200_U433 = ~new_P2_U3902 | ~new_P2_R1200_U84;
  assign new_P2_R1200_U434 = ~new_P2_U3074 | ~new_P2_R1200_U81;
  assign new_P2_R1200_U435 = ~new_P2_R1200_U317 | ~new_P2_R1200_U172;
  assign new_P2_R1200_U436 = ~new_P2_R1200_U280 | ~new_P2_R1200_U171;
  assign new_P2_R1200_U437 = ~new_P2_U3903 | ~new_P2_R1200_U78;
  assign new_P2_R1200_U438 = ~new_P2_U3075 | ~new_P2_R1200_U77;
  assign new_P2_R1200_U439 = ~new_P2_R1200_U145;
  assign new_P2_R1200_U440 = ~new_P2_R1200_U276 | ~new_P2_R1200_U439;
  assign new_P2_R1200_U441 = ~new_P2_R1200_U145 | ~new_P2_R1200_U173;
  assign new_P2_R1200_U442 = ~new_P2_U3392 | ~new_P2_R1200_U39;
  assign new_P2_R1200_U443 = ~new_P2_U3077 | ~new_P2_R1200_U174;
  assign new_P2_R1200_U444 = ~new_P2_R1200_U146;
  assign new_P2_R1200_U445 = ~new_P2_R1200_U203 | ~new_P2_R1200_U444;
  assign new_P2_R1200_U446 = ~new_P2_R1200_U146 | ~new_P2_R1200_U175;
  assign new_P2_R1200_U447 = ~new_P2_U3445 | ~new_P2_R1200_U76;
  assign new_P2_R1200_U448 = ~new_P2_U3080 | ~new_P2_R1200_U75;
  assign new_P2_R1200_U449 = ~new_P2_R1200_U147;
  assign new_P2_R1200_U450 = ~new_P2_R1200_U272 | ~new_P2_R1200_U449;
  assign new_P2_R1200_U451 = ~new_P2_R1200_U147 | ~new_P2_R1200_U176;
  assign new_P2_R1200_U452 = ~new_P2_U3443 | ~new_P2_R1200_U74;
  assign new_P2_R1200_U453 = ~new_P2_U3081 | ~new_P2_R1200_U177;
  assign new_P2_R1200_U454 = ~new_P2_R1200_U148;
  assign new_P2_R1200_U455 = ~new_P2_R1200_U270 | ~new_P2_R1200_U454;
  assign new_P2_R1200_U456 = ~new_P2_R1200_U148 | ~new_P2_R1200_U178;
  assign new_P2_R1200_U457 = ~new_P2_U3440 | ~new_P2_R1200_U73;
  assign new_P2_R1200_U458 = ~new_P2_U3068 | ~new_P2_R1200_U72;
  assign new_P2_R1200_U459 = ~new_P2_R1200_U149;
  assign new_P2_R1200_U460 = ~new_P2_R1200_U266 | ~new_P2_R1200_U459;
  assign new_P2_R1200_U461 = ~new_P2_R1200_U149 | ~new_P2_R1200_U179;
  assign new_P2_R1200_U462 = ~new_P2_U3437 | ~new_P2_R1200_U68;
  assign new_P2_R1200_U463 = ~new_P2_U3072 | ~new_P2_R1200_U65;
  assign new_P2_R1200_U464 = ~new_P2_R1200_U463 | ~new_P2_R1200_U462;
  assign new_P2_R1200_U465 = ~new_P2_U3434 | ~new_P2_R1200_U69;
  assign new_P2_R1200_U466 = ~new_P2_U3073 | ~new_P2_R1200_U66;
  assign new_P2_R1200_U467 = ~new_P2_R1200_U327 | ~new_P2_R1200_U95;
  assign new_P2_R1200_U468 = ~new_P2_R1200_U180 | ~new_P2_R1200_U319;
  assign new_P2_R1200_U469 = ~new_P2_U3431 | ~new_P2_R1200_U70;
  assign new_P2_R1200_U470 = ~new_P2_U3078 | ~new_P2_R1200_U67;
  assign new_P2_R1200_U471 = ~new_P2_R1200_U328 | ~new_P2_R1200_U182;
  assign new_P2_R1200_U472 = ~new_P2_R1200_U256 | ~new_P2_R1200_U181;
  assign new_P2_R1200_U473 = ~new_P2_U3428 | ~new_P2_R1200_U64;
  assign new_P2_R1200_U474 = ~new_P2_U3079 | ~new_P2_R1200_U63;
  assign new_P2_R1200_U475 = ~new_P2_R1200_U152;
  assign new_P2_R1200_U476 = ~new_P2_R1200_U354 | ~new_P2_R1200_U475;
  assign new_P2_R1200_U477 = ~new_P2_R1200_U152 | ~new_P2_R1200_U183;
  assign new_P2_R1200_U478 = ~new_P2_U3425 | ~new_P2_R1200_U55;
  assign new_P2_R1200_U479 = ~new_P2_U3071 | ~new_P2_R1200_U61;
  assign new_P2_R1200_U480 = ~new_P2_R1200_U153;
  assign new_P2_R1200_U481 = ~new_P2_R1200_U352 | ~new_P2_R1200_U480;
  assign new_P2_R1200_U482 = ~new_P2_R1200_U153 | ~new_P2_R1200_U184;
  assign new_P2_R1200_U483 = ~new_P2_U3422 | ~new_P2_R1200_U56;
  assign new_P2_R1200_U484 = ~new_P2_U3062 | ~new_P2_R1200_U60;
  assign new_P2_R1200_U485 = ~new_P2_R1200_U484 | ~new_P2_R1200_U483;
  assign new_P2_R1200_U486 = ~new_P2_U3419 | ~new_P2_R1200_U57;
  assign new_P2_R1200_U487 = ~new_P2_U3061 | ~new_P2_R1200_U58;
  assign new_P2_R1200_U488 = ~new_P2_R1200_U96 | ~new_P2_R1200_U336;
  assign new_P2_R1200_U489 = ~new_P2_R1200_U185 | ~new_P2_R1200_U350;
  assign new_P2_R1179_U6 = new_P2_R1179_U212 & new_P2_R1179_U211;
  assign new_P2_R1179_U7 = new_P2_R1179_U246 & new_P2_R1179_U245;
  assign new_P2_R1179_U8 = new_P2_R1179_U193 & new_P2_R1179_U257;
  assign new_P2_R1179_U9 = new_P2_R1179_U259 & new_P2_R1179_U258;
  assign new_P2_R1179_U10 = new_P2_R1179_U194 & new_P2_R1179_U281;
  assign new_P2_R1179_U11 = new_P2_R1179_U283 & new_P2_R1179_U282;
  assign new_P2_R1179_U12 = new_P2_R1179_U299 & new_P2_R1179_U195;
  assign new_P2_R1179_U13 = new_P2_R1179_U215 & new_P2_R1179_U210 & new_P2_R1179_U197;
  assign new_P2_R1179_U14 = new_P2_R1179_U220 & new_P2_R1179_U198;
  assign new_P2_R1179_U15 = new_P2_R1179_U244 & new_P2_R1179_U224 & new_P2_R1179_U192;
  assign new_P2_R1179_U16 = new_P2_R1179_U399 & new_P2_R1179_U398;
  assign new_P2_R1179_U17 = ~new_P2_R1179_U331 | ~new_P2_R1179_U334;
  assign new_P2_R1179_U18 = ~new_P2_R1179_U322 | ~new_P2_R1179_U325;
  assign new_P2_R1179_U19 = ~new_P2_R1179_U311 | ~new_P2_R1179_U314;
  assign new_P2_R1179_U20 = ~new_P2_R1179_U305 | ~new_P2_R1179_U357;
  assign new_P2_R1179_U21 = ~new_P2_R1179_U137 | ~new_P2_R1179_U186;
  assign new_P2_R1179_U22 = ~new_P2_R1179_U242 | ~new_P2_R1179_U347;
  assign new_P2_R1179_U23 = ~new_P2_R1179_U235 | ~new_P2_R1179_U238;
  assign new_P2_R1179_U24 = ~new_P2_R1179_U227 | ~new_P2_R1179_U229;
  assign new_P2_R1179_U25 = ~new_P2_R1179_U175 | ~new_P2_R1179_U337;
  assign new_P2_R1179_U26 = ~new_P2_U3069;
  assign new_P2_R1179_U27 = ~new_P2_U3069 | ~new_P2_R1179_U32;
  assign new_P2_R1179_U28 = ~new_P2_U3083;
  assign new_P2_R1179_U29 = ~new_P2_U3404;
  assign new_P2_R1179_U30 = ~new_P2_U3407;
  assign new_P2_R1179_U31 = ~new_P2_U3401;
  assign new_P2_R1179_U32 = ~new_P2_U3410;
  assign new_P2_R1179_U33 = ~new_P2_U3413;
  assign new_P2_R1179_U34 = ~new_P2_U3067;
  assign new_P2_R1179_U35 = ~new_P2_U3067 | ~new_P2_R1179_U37;
  assign new_P2_R1179_U36 = ~new_P2_U3063;
  assign new_P2_R1179_U37 = ~new_P2_U3395;
  assign new_P2_R1179_U38 = ~new_P2_U3387;
  assign new_P2_R1179_U39 = ~new_P2_U3077;
  assign new_P2_R1179_U40 = ~new_P2_U3398;
  assign new_P2_R1179_U41 = ~new_P2_U3070;
  assign new_P2_R1179_U42 = ~new_P2_U3066;
  assign new_P2_R1179_U43 = ~new_P2_U3059;
  assign new_P2_R1179_U44 = ~new_P2_U3059 | ~new_P2_R1179_U31;
  assign new_P2_R1179_U45 = ~new_P2_R1179_U216 | ~new_P2_R1179_U214;
  assign new_P2_R1179_U46 = ~new_P2_U3416;
  assign new_P2_R1179_U47 = ~new_P2_U3082;
  assign new_P2_R1179_U48 = ~new_P2_R1179_U45 | ~new_P2_R1179_U217;
  assign new_P2_R1179_U49 = ~new_P2_R1179_U44 | ~new_P2_R1179_U231;
  assign new_P2_R1179_U50 = ~new_P2_R1179_U338 | ~new_P2_R1179_U204 | ~new_P2_R1179_U188;
  assign new_P2_R1179_U51 = ~new_P2_U3895;
  assign new_P2_R1179_U52 = ~new_P2_U3056;
  assign new_P2_R1179_U53 = ~new_P2_U3056 | ~new_P2_R1179_U90;
  assign new_P2_R1179_U54 = ~new_P2_U3052;
  assign new_P2_R1179_U55 = ~new_P2_U3071;
  assign new_P2_R1179_U56 = ~new_P2_U3062;
  assign new_P2_R1179_U57 = ~new_P2_U3061;
  assign new_P2_R1179_U58 = ~new_P2_U3419;
  assign new_P2_R1179_U59 = ~new_P2_U3082 | ~new_P2_R1179_U46;
  assign new_P2_R1179_U60 = ~new_P2_U3422;
  assign new_P2_R1179_U61 = ~new_P2_U3425;
  assign new_P2_R1179_U62 = ~new_P2_R1179_U249 | ~new_P2_R1179_U248;
  assign new_P2_R1179_U63 = ~new_P2_U3428;
  assign new_P2_R1179_U64 = ~new_P2_U3079;
  assign new_P2_R1179_U65 = ~new_P2_U3437;
  assign new_P2_R1179_U66 = ~new_P2_U3434;
  assign new_P2_R1179_U67 = ~new_P2_U3431;
  assign new_P2_R1179_U68 = ~new_P2_U3072;
  assign new_P2_R1179_U69 = ~new_P2_U3073;
  assign new_P2_R1179_U70 = ~new_P2_U3078;
  assign new_P2_R1179_U71 = ~new_P2_U3078 | ~new_P2_R1179_U67;
  assign new_P2_R1179_U72 = ~new_P2_U3440;
  assign new_P2_R1179_U73 = ~new_P2_U3068;
  assign new_P2_R1179_U74 = ~new_P2_U3081;
  assign new_P2_R1179_U75 = ~new_P2_U3445;
  assign new_P2_R1179_U76 = ~new_P2_U3080;
  assign new_P2_R1179_U77 = ~new_P2_U3903;
  assign new_P2_R1179_U78 = ~new_P2_U3075;
  assign new_P2_R1179_U79 = ~new_P2_U3900;
  assign new_P2_R1179_U80 = ~new_P2_U3901;
  assign new_P2_R1179_U81 = ~new_P2_U3902;
  assign new_P2_R1179_U82 = ~new_P2_U3065;
  assign new_P2_R1179_U83 = ~new_P2_U3060;
  assign new_P2_R1179_U84 = ~new_P2_U3074;
  assign new_P2_R1179_U85 = ~new_P2_U3074 | ~new_P2_R1179_U81;
  assign new_P2_R1179_U86 = ~new_P2_U3899;
  assign new_P2_R1179_U87 = ~new_P2_U3064;
  assign new_P2_R1179_U88 = ~new_P2_U3898;
  assign new_P2_R1179_U89 = ~new_P2_U3057;
  assign new_P2_R1179_U90 = ~new_P2_U3897;
  assign new_P2_R1179_U91 = ~new_P2_U3896;
  assign new_P2_R1179_U92 = ~new_P2_U3053;
  assign new_P2_R1179_U93 = ~new_P2_R1179_U297 | ~new_P2_R1179_U296;
  assign new_P2_R1179_U94 = ~new_P2_R1179_U85 | ~new_P2_R1179_U307;
  assign new_P2_R1179_U95 = ~new_P2_R1179_U71 | ~new_P2_R1179_U318;
  assign new_P2_R1179_U96 = ~new_P2_R1179_U349 | ~new_P2_R1179_U59;
  assign new_P2_R1179_U97 = ~new_P2_U3076;
  assign new_P2_R1179_U98 = ~new_P2_R1179_U406 | ~new_P2_R1179_U405;
  assign new_P2_R1179_U99 = ~new_P2_R1179_U420 | ~new_P2_R1179_U419;
  assign new_P2_R1179_U100 = ~new_P2_R1179_U425 | ~new_P2_R1179_U424;
  assign new_P2_R1179_U101 = ~new_P2_R1179_U441 | ~new_P2_R1179_U440;
  assign new_P2_R1179_U102 = ~new_P2_R1179_U446 | ~new_P2_R1179_U445;
  assign new_P2_R1179_U103 = ~new_P2_R1179_U451 | ~new_P2_R1179_U450;
  assign new_P2_R1179_U104 = ~new_P2_R1179_U456 | ~new_P2_R1179_U455;
  assign new_P2_R1179_U105 = ~new_P2_R1179_U461 | ~new_P2_R1179_U460;
  assign new_P2_R1179_U106 = ~new_P2_R1179_U477 | ~new_P2_R1179_U476;
  assign new_P2_R1179_U107 = ~new_P2_R1179_U482 | ~new_P2_R1179_U481;
  assign new_P2_R1179_U108 = ~new_P2_R1179_U365 | ~new_P2_R1179_U364;
  assign new_P2_R1179_U109 = ~new_P2_R1179_U374 | ~new_P2_R1179_U373;
  assign new_P2_R1179_U110 = ~new_P2_R1179_U381 | ~new_P2_R1179_U380;
  assign new_P2_R1179_U111 = ~new_P2_R1179_U385 | ~new_P2_R1179_U384;
  assign new_P2_R1179_U112 = ~new_P2_R1179_U394 | ~new_P2_R1179_U393;
  assign new_P2_R1179_U113 = ~new_P2_R1179_U415 | ~new_P2_R1179_U414;
  assign new_P2_R1179_U114 = ~new_P2_R1179_U432 | ~new_P2_R1179_U431;
  assign new_P2_R1179_U115 = ~new_P2_R1179_U436 | ~new_P2_R1179_U435;
  assign new_P2_R1179_U116 = ~new_P2_R1179_U468 | ~new_P2_R1179_U467;
  assign new_P2_R1179_U117 = ~new_P2_R1179_U472 | ~new_P2_R1179_U471;
  assign new_P2_R1179_U118 = ~new_P2_R1179_U489 | ~new_P2_R1179_U488;
  assign new_P2_R1179_U119 = new_P2_R1179_U206 & new_P2_R1179_U196;
  assign new_P2_R1179_U120 = new_P2_R1179_U209 & new_P2_R1179_U208;
  assign new_P2_R1179_U121 = new_P2_R1179_U14 & new_P2_R1179_U13;
  assign new_P2_R1179_U122 = new_P2_R1179_U340 & new_P2_R1179_U222;
  assign new_P2_R1179_U123 = new_P2_R1179_U342 & new_P2_R1179_U122;
  assign new_P2_R1179_U124 = new_P2_R1179_U27 & new_P2_R1179_U367 & new_P2_R1179_U366;
  assign new_P2_R1179_U125 = new_P2_R1179_U370 & new_P2_R1179_U198;
  assign new_P2_R1179_U126 = new_P2_R1179_U237 & new_P2_R1179_U6;
  assign new_P2_R1179_U127 = new_P2_R1179_U377 & new_P2_R1179_U197;
  assign new_P2_R1179_U128 = new_P2_R1179_U35 & new_P2_R1179_U387 & new_P2_R1179_U386;
  assign new_P2_R1179_U129 = new_P2_R1179_U390 & new_P2_R1179_U196;
  assign new_P2_R1179_U130 = new_P2_R1179_U251 & new_P2_R1179_U15;
  assign new_P2_R1179_U131 = new_P2_R1179_U343 & new_P2_R1179_U252;
  assign new_P2_R1179_U132 = new_P2_R1179_U262 & new_P2_R1179_U8;
  assign new_P2_R1179_U133 = new_P2_R1179_U286 & new_P2_R1179_U10;
  assign new_P2_R1179_U134 = new_P2_R1179_U302 & new_P2_R1179_U301;
  assign new_P2_R1179_U135 = new_P2_R1179_U397 & new_P2_R1179_U303;
  assign new_P2_R1179_U136 = new_P2_R1179_U16 & new_P2_R1179_U304 & new_P2_R1179_U302 & new_P2_R1179_U301;
  assign new_P2_R1179_U137 = new_P2_R1179_U359 & new_P2_R1179_U165;
  assign new_P2_R1179_U138 = ~new_P2_R1179_U403 | ~new_P2_R1179_U402;
  assign new_P2_R1179_U139 = new_P2_R1179_U53 & new_P2_R1179_U408 & new_P2_R1179_U407;
  assign new_P2_R1179_U140 = new_P2_R1179_U411 & new_P2_R1179_U195;
  assign new_P2_R1179_U141 = ~new_P2_R1179_U417 | ~new_P2_R1179_U416;
  assign new_P2_R1179_U142 = ~new_P2_R1179_U422 | ~new_P2_R1179_U421;
  assign new_P2_R1179_U143 = new_P2_R1179_U313 & new_P2_R1179_U11;
  assign new_P2_R1179_U144 = new_P2_R1179_U428 & new_P2_R1179_U194;
  assign new_P2_R1179_U145 = ~new_P2_R1179_U438 | ~new_P2_R1179_U437;
  assign new_P2_R1179_U146 = ~new_P2_R1179_U443 | ~new_P2_R1179_U442;
  assign new_P2_R1179_U147 = ~new_P2_R1179_U448 | ~new_P2_R1179_U447;
  assign new_P2_R1179_U148 = ~new_P2_R1179_U453 | ~new_P2_R1179_U452;
  assign new_P2_R1179_U149 = ~new_P2_R1179_U458 | ~new_P2_R1179_U457;
  assign new_P2_R1179_U150 = new_P2_R1179_U324 & new_P2_R1179_U9;
  assign new_P2_R1179_U151 = new_P2_R1179_U464 & new_P2_R1179_U193;
  assign new_P2_R1179_U152 = ~new_P2_R1179_U474 | ~new_P2_R1179_U473;
  assign new_P2_R1179_U153 = ~new_P2_R1179_U479 | ~new_P2_R1179_U478;
  assign new_P2_R1179_U154 = new_P2_R1179_U333 & new_P2_R1179_U7;
  assign new_P2_R1179_U155 = new_P2_R1179_U485 & new_P2_R1179_U192;
  assign new_P2_R1179_U156 = new_P2_R1179_U363 & new_P2_R1179_U362;
  assign new_P2_R1179_U157 = ~new_P2_R1179_U123 | ~new_P2_R1179_U341;
  assign new_P2_R1179_U158 = new_P2_R1179_U372 & new_P2_R1179_U371;
  assign new_P2_R1179_U159 = new_P2_R1179_U379 & new_P2_R1179_U378;
  assign new_P2_R1179_U160 = new_P2_R1179_U383 & new_P2_R1179_U382;
  assign new_P2_R1179_U161 = ~new_P2_R1179_U120 | ~new_P2_R1179_U344;
  assign new_P2_R1179_U162 = new_P2_R1179_U392 & new_P2_R1179_U391;
  assign new_P2_R1179_U163 = ~new_P2_U3904;
  assign new_P2_R1179_U164 = ~new_P2_U3054;
  assign new_P2_R1179_U165 = new_P2_R1179_U401 & new_P2_R1179_U400;
  assign new_P2_R1179_U166 = ~new_P2_R1179_U134 | ~new_P2_R1179_U360;
  assign new_P2_R1179_U167 = new_P2_R1179_U413 & new_P2_R1179_U412;
  assign new_P2_R1179_U168 = ~new_P2_R1179_U293 | ~new_P2_R1179_U292;
  assign new_P2_R1179_U169 = ~new_P2_R1179_U289 | ~new_P2_R1179_U288;
  assign new_P2_R1179_U170 = new_P2_R1179_U430 & new_P2_R1179_U429;
  assign new_P2_R1179_U171 = new_P2_R1179_U434 & new_P2_R1179_U433;
  assign new_P2_R1179_U172 = ~new_P2_R1179_U279 | ~new_P2_R1179_U278;
  assign new_P2_R1179_U173 = ~new_P2_R1179_U275 | ~new_P2_R1179_U274;
  assign new_P2_R1179_U174 = ~new_P2_U3392;
  assign new_P2_R1179_U175 = ~new_P2_U3387 | ~new_P2_R1179_U97;
  assign new_P2_R1179_U176 = ~new_P2_R1179_U339 | ~new_P2_R1179_U271 | ~new_P2_R1179_U187;
  assign new_P2_R1179_U177 = ~new_P2_U3443;
  assign new_P2_R1179_U178 = ~new_P2_R1179_U269 | ~new_P2_R1179_U268;
  assign new_P2_R1179_U179 = ~new_P2_R1179_U265 | ~new_P2_R1179_U264;
  assign new_P2_R1179_U180 = new_P2_R1179_U466 & new_P2_R1179_U465;
  assign new_P2_R1179_U181 = new_P2_R1179_U470 & new_P2_R1179_U469;
  assign new_P2_R1179_U182 = ~new_P2_R1179_U255 | ~new_P2_R1179_U254;
  assign new_P2_R1179_U183 = ~new_P2_R1179_U131 | ~new_P2_R1179_U353;
  assign new_P2_R1179_U184 = ~new_P2_R1179_U351 | ~new_P2_R1179_U62;
  assign new_P2_R1179_U185 = new_P2_R1179_U487 & new_P2_R1179_U486;
  assign new_P2_R1179_U186 = ~new_P2_R1179_U135 | ~new_P2_R1179_U166;
  assign new_P2_R1179_U187 = ~new_P2_R1179_U178 | ~new_P2_R1179_U177;
  assign new_P2_R1179_U188 = ~new_P2_R1179_U175 | ~new_P2_R1179_U174;
  assign new_P2_R1179_U189 = ~new_P2_R1179_U53;
  assign new_P2_R1179_U190 = ~new_P2_R1179_U35;
  assign new_P2_R1179_U191 = ~new_P2_R1179_U27;
  assign new_P2_R1179_U192 = ~new_P2_U3419 | ~new_P2_R1179_U57;
  assign new_P2_R1179_U193 = ~new_P2_U3434 | ~new_P2_R1179_U69;
  assign new_P2_R1179_U194 = ~new_P2_U3901 | ~new_P2_R1179_U83;
  assign new_P2_R1179_U195 = ~new_P2_U3897 | ~new_P2_R1179_U52;
  assign new_P2_R1179_U196 = ~new_P2_U3395 | ~new_P2_R1179_U34;
  assign new_P2_R1179_U197 = ~new_P2_U3404 | ~new_P2_R1179_U42;
  assign new_P2_R1179_U198 = ~new_P2_U3410 | ~new_P2_R1179_U26;
  assign new_P2_R1179_U199 = ~new_P2_R1179_U71;
  assign new_P2_R1179_U200 = ~new_P2_R1179_U85;
  assign new_P2_R1179_U201 = ~new_P2_R1179_U44;
  assign new_P2_R1179_U202 = ~new_P2_R1179_U59;
  assign new_P2_R1179_U203 = ~new_P2_R1179_U175;
  assign new_P2_R1179_U204 = ~new_P2_U3077 | ~new_P2_R1179_U175;
  assign new_P2_R1179_U205 = ~new_P2_R1179_U50;
  assign new_P2_R1179_U206 = ~new_P2_U3398 | ~new_P2_R1179_U36;
  assign new_P2_R1179_U207 = ~new_P2_R1179_U36 | ~new_P2_R1179_U35;
  assign new_P2_R1179_U208 = ~new_P2_R1179_U207 | ~new_P2_R1179_U40;
  assign new_P2_R1179_U209 = ~new_P2_U3063 | ~new_P2_R1179_U190;
  assign new_P2_R1179_U210 = ~new_P2_U3407 | ~new_P2_R1179_U41;
  assign new_P2_R1179_U211 = ~new_P2_U3070 | ~new_P2_R1179_U30;
  assign new_P2_R1179_U212 = ~new_P2_U3066 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U213 = ~new_P2_R1179_U201 | ~new_P2_R1179_U197;
  assign new_P2_R1179_U214 = ~new_P2_R1179_U6 | ~new_P2_R1179_U213;
  assign new_P2_R1179_U215 = ~new_P2_U3401 | ~new_P2_R1179_U43;
  assign new_P2_R1179_U216 = ~new_P2_U3407 | ~new_P2_R1179_U41;
  assign new_P2_R1179_U217 = ~new_P2_R1179_U13 | ~new_P2_R1179_U161;
  assign new_P2_R1179_U218 = ~new_P2_R1179_U45;
  assign new_P2_R1179_U219 = ~new_P2_R1179_U48;
  assign new_P2_R1179_U220 = ~new_P2_U3413 | ~new_P2_R1179_U28;
  assign new_P2_R1179_U221 = ~new_P2_R1179_U28 | ~new_P2_R1179_U27;
  assign new_P2_R1179_U222 = ~new_P2_U3083 | ~new_P2_R1179_U191;
  assign new_P2_R1179_U223 = ~new_P2_R1179_U157;
  assign new_P2_R1179_U224 = ~new_P2_U3416 | ~new_P2_R1179_U47;
  assign new_P2_R1179_U225 = ~new_P2_R1179_U224 | ~new_P2_R1179_U59;
  assign new_P2_R1179_U226 = ~new_P2_R1179_U219 | ~new_P2_R1179_U27;
  assign new_P2_R1179_U227 = ~new_P2_R1179_U125 | ~new_P2_R1179_U226;
  assign new_P2_R1179_U228 = ~new_P2_R1179_U48 | ~new_P2_R1179_U198;
  assign new_P2_R1179_U229 = ~new_P2_R1179_U124 | ~new_P2_R1179_U228;
  assign new_P2_R1179_U230 = ~new_P2_R1179_U27 | ~new_P2_R1179_U198;
  assign new_P2_R1179_U231 = ~new_P2_R1179_U215 | ~new_P2_R1179_U161;
  assign new_P2_R1179_U232 = ~new_P2_R1179_U49;
  assign new_P2_R1179_U233 = ~new_P2_U3066 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U234 = ~new_P2_R1179_U232 | ~new_P2_R1179_U233;
  assign new_P2_R1179_U235 = ~new_P2_R1179_U127 | ~new_P2_R1179_U234;
  assign new_P2_R1179_U236 = ~new_P2_R1179_U49 | ~new_P2_R1179_U197;
  assign new_P2_R1179_U237 = ~new_P2_U3407 | ~new_P2_R1179_U41;
  assign new_P2_R1179_U238 = ~new_P2_R1179_U126 | ~new_P2_R1179_U236;
  assign new_P2_R1179_U239 = ~new_P2_U3066 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U240 = ~new_P2_R1179_U239 | ~new_P2_R1179_U197;
  assign new_P2_R1179_U241 = ~new_P2_R1179_U215 | ~new_P2_R1179_U44;
  assign new_P2_R1179_U242 = ~new_P2_R1179_U129 | ~new_P2_R1179_U348;
  assign new_P2_R1179_U243 = ~new_P2_R1179_U35 | ~new_P2_R1179_U196;
  assign new_P2_R1179_U244 = ~new_P2_U3422 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U245 = ~new_P2_U3062 | ~new_P2_R1179_U60;
  assign new_P2_R1179_U246 = ~new_P2_U3061 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U247 = ~new_P2_R1179_U202 | ~new_P2_R1179_U192;
  assign new_P2_R1179_U248 = ~new_P2_R1179_U7 | ~new_P2_R1179_U247;
  assign new_P2_R1179_U249 = ~new_P2_U3422 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U250 = ~new_P2_R1179_U62;
  assign new_P2_R1179_U251 = ~new_P2_U3425 | ~new_P2_R1179_U55;
  assign new_P2_R1179_U252 = ~new_P2_U3071 | ~new_P2_R1179_U61;
  assign new_P2_R1179_U253 = ~new_P2_U3428 | ~new_P2_R1179_U64;
  assign new_P2_R1179_U254 = ~new_P2_R1179_U253 | ~new_P2_R1179_U183;
  assign new_P2_R1179_U255 = ~new_P2_U3079 | ~new_P2_R1179_U63;
  assign new_P2_R1179_U256 = ~new_P2_R1179_U182;
  assign new_P2_R1179_U257 = ~new_P2_U3437 | ~new_P2_R1179_U68;
  assign new_P2_R1179_U258 = ~new_P2_U3072 | ~new_P2_R1179_U65;
  assign new_P2_R1179_U259 = ~new_P2_U3073 | ~new_P2_R1179_U66;
  assign new_P2_R1179_U260 = ~new_P2_R1179_U199 | ~new_P2_R1179_U8;
  assign new_P2_R1179_U261 = ~new_P2_R1179_U9 | ~new_P2_R1179_U260;
  assign new_P2_R1179_U262 = ~new_P2_U3431 | ~new_P2_R1179_U70;
  assign new_P2_R1179_U263 = ~new_P2_U3437 | ~new_P2_R1179_U68;
  assign new_P2_R1179_U264 = ~new_P2_R1179_U132 | ~new_P2_R1179_U182;
  assign new_P2_R1179_U265 = ~new_P2_R1179_U263 | ~new_P2_R1179_U261;
  assign new_P2_R1179_U266 = ~new_P2_R1179_U179;
  assign new_P2_R1179_U267 = ~new_P2_U3440 | ~new_P2_R1179_U73;
  assign new_P2_R1179_U268 = ~new_P2_R1179_U267 | ~new_P2_R1179_U179;
  assign new_P2_R1179_U269 = ~new_P2_U3068 | ~new_P2_R1179_U72;
  assign new_P2_R1179_U270 = ~new_P2_R1179_U178;
  assign new_P2_R1179_U271 = ~new_P2_U3081 | ~new_P2_R1179_U178;
  assign new_P2_R1179_U272 = ~new_P2_R1179_U176;
  assign new_P2_R1179_U273 = ~new_P2_U3445 | ~new_P2_R1179_U76;
  assign new_P2_R1179_U274 = ~new_P2_R1179_U273 | ~new_P2_R1179_U176;
  assign new_P2_R1179_U275 = ~new_P2_U3080 | ~new_P2_R1179_U75;
  assign new_P2_R1179_U276 = ~new_P2_R1179_U173;
  assign new_P2_R1179_U277 = ~new_P2_U3903 | ~new_P2_R1179_U78;
  assign new_P2_R1179_U278 = ~new_P2_R1179_U277 | ~new_P2_R1179_U173;
  assign new_P2_R1179_U279 = ~new_P2_U3075 | ~new_P2_R1179_U77;
  assign new_P2_R1179_U280 = ~new_P2_R1179_U172;
  assign new_P2_R1179_U281 = ~new_P2_U3900 | ~new_P2_R1179_U82;
  assign new_P2_R1179_U282 = ~new_P2_U3065 | ~new_P2_R1179_U79;
  assign new_P2_R1179_U283 = ~new_P2_U3060 | ~new_P2_R1179_U80;
  assign new_P2_R1179_U284 = ~new_P2_R1179_U200 | ~new_P2_R1179_U10;
  assign new_P2_R1179_U285 = ~new_P2_R1179_U11 | ~new_P2_R1179_U284;
  assign new_P2_R1179_U286 = ~new_P2_U3902 | ~new_P2_R1179_U84;
  assign new_P2_R1179_U287 = ~new_P2_U3900 | ~new_P2_R1179_U82;
  assign new_P2_R1179_U288 = ~new_P2_R1179_U133 | ~new_P2_R1179_U172;
  assign new_P2_R1179_U289 = ~new_P2_R1179_U287 | ~new_P2_R1179_U285;
  assign new_P2_R1179_U290 = ~new_P2_R1179_U169;
  assign new_P2_R1179_U291 = ~new_P2_U3899 | ~new_P2_R1179_U87;
  assign new_P2_R1179_U292 = ~new_P2_R1179_U291 | ~new_P2_R1179_U169;
  assign new_P2_R1179_U293 = ~new_P2_U3064 | ~new_P2_R1179_U86;
  assign new_P2_R1179_U294 = ~new_P2_R1179_U168;
  assign new_P2_R1179_U295 = ~new_P2_U3898 | ~new_P2_R1179_U89;
  assign new_P2_R1179_U296 = ~new_P2_R1179_U295 | ~new_P2_R1179_U168;
  assign new_P2_R1179_U297 = ~new_P2_U3057 | ~new_P2_R1179_U88;
  assign new_P2_R1179_U298 = ~new_P2_R1179_U93;
  assign new_P2_R1179_U299 = ~new_P2_U3896 | ~new_P2_R1179_U54;
  assign new_P2_R1179_U300 = ~new_P2_R1179_U54 | ~new_P2_R1179_U53;
  assign new_P2_R1179_U301 = ~new_P2_R1179_U300 | ~new_P2_R1179_U91;
  assign new_P2_R1179_U302 = ~new_P2_U3052 | ~new_P2_R1179_U189;
  assign new_P2_R1179_U303 = ~new_P2_U3895 | ~new_P2_R1179_U92;
  assign new_P2_R1179_U304 = ~new_P2_U3053 | ~new_P2_R1179_U51;
  assign new_P2_R1179_U305 = ~new_P2_R1179_U140 | ~new_P2_R1179_U355;
  assign new_P2_R1179_U306 = ~new_P2_R1179_U53 | ~new_P2_R1179_U195;
  assign new_P2_R1179_U307 = ~new_P2_R1179_U286 | ~new_P2_R1179_U172;
  assign new_P2_R1179_U308 = ~new_P2_R1179_U94;
  assign new_P2_R1179_U309 = ~new_P2_U3060 | ~new_P2_R1179_U80;
  assign new_P2_R1179_U310 = ~new_P2_R1179_U308 | ~new_P2_R1179_U309;
  assign new_P2_R1179_U311 = ~new_P2_R1179_U144 | ~new_P2_R1179_U310;
  assign new_P2_R1179_U312 = ~new_P2_R1179_U94 | ~new_P2_R1179_U194;
  assign new_P2_R1179_U313 = ~new_P2_U3900 | ~new_P2_R1179_U82;
  assign new_P2_R1179_U314 = ~new_P2_R1179_U143 | ~new_P2_R1179_U312;
  assign new_P2_R1179_U315 = ~new_P2_U3060 | ~new_P2_R1179_U80;
  assign new_P2_R1179_U316 = ~new_P2_R1179_U194 | ~new_P2_R1179_U315;
  assign new_P2_R1179_U317 = ~new_P2_R1179_U286 | ~new_P2_R1179_U85;
  assign new_P2_R1179_U318 = ~new_P2_R1179_U262 | ~new_P2_R1179_U182;
  assign new_P2_R1179_U319 = ~new_P2_R1179_U95;
  assign new_P2_R1179_U320 = ~new_P2_U3073 | ~new_P2_R1179_U66;
  assign new_P2_R1179_U321 = ~new_P2_R1179_U319 | ~new_P2_R1179_U320;
  assign new_P2_R1179_U322 = ~new_P2_R1179_U151 | ~new_P2_R1179_U321;
  assign new_P2_R1179_U323 = ~new_P2_R1179_U95 | ~new_P2_R1179_U193;
  assign new_P2_R1179_U324 = ~new_P2_U3437 | ~new_P2_R1179_U68;
  assign new_P2_R1179_U325 = ~new_P2_R1179_U150 | ~new_P2_R1179_U323;
  assign new_P2_R1179_U326 = ~new_P2_U3073 | ~new_P2_R1179_U66;
  assign new_P2_R1179_U327 = ~new_P2_R1179_U193 | ~new_P2_R1179_U326;
  assign new_P2_R1179_U328 = ~new_P2_R1179_U262 | ~new_P2_R1179_U71;
  assign new_P2_R1179_U329 = ~new_P2_U3061 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U330 = ~new_P2_R1179_U350 | ~new_P2_R1179_U329;
  assign new_P2_R1179_U331 = ~new_P2_R1179_U155 | ~new_P2_R1179_U330;
  assign new_P2_R1179_U332 = ~new_P2_R1179_U96 | ~new_P2_R1179_U192;
  assign new_P2_R1179_U333 = ~new_P2_U3422 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U334 = ~new_P2_R1179_U154 | ~new_P2_R1179_U332;
  assign new_P2_R1179_U335 = ~new_P2_U3061 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U336 = ~new_P2_R1179_U192 | ~new_P2_R1179_U335;
  assign new_P2_R1179_U337 = ~new_P2_U3076 | ~new_P2_R1179_U38;
  assign new_P2_R1179_U338 = ~new_P2_U3077 | ~new_P2_R1179_U174;
  assign new_P2_R1179_U339 = ~new_P2_U3081 | ~new_P2_R1179_U177;
  assign new_P2_R1179_U340 = ~new_P2_R1179_U33 | ~new_P2_R1179_U221;
  assign new_P2_R1179_U341 = ~new_P2_R1179_U121 | ~new_P2_R1179_U161;
  assign new_P2_R1179_U342 = ~new_P2_R1179_U218 | ~new_P2_R1179_U14;
  assign new_P2_R1179_U343 = ~new_P2_R1179_U250 | ~new_P2_R1179_U251;
  assign new_P2_R1179_U344 = ~new_P2_R1179_U119 | ~new_P2_R1179_U50;
  assign new_P2_R1179_U345 = ~new_P2_R1179_U161;
  assign new_P2_R1179_U346 = ~new_P2_R1179_U196 | ~new_P2_R1179_U50;
  assign new_P2_R1179_U347 = ~new_P2_R1179_U128 | ~new_P2_R1179_U346;
  assign new_P2_R1179_U348 = ~new_P2_R1179_U205 | ~new_P2_R1179_U35;
  assign new_P2_R1179_U349 = ~new_P2_R1179_U224 | ~new_P2_R1179_U157;
  assign new_P2_R1179_U350 = ~new_P2_R1179_U96;
  assign new_P2_R1179_U351 = ~new_P2_R1179_U15 | ~new_P2_R1179_U157;
  assign new_P2_R1179_U352 = ~new_P2_R1179_U184;
  assign new_P2_R1179_U353 = ~new_P2_R1179_U130 | ~new_P2_R1179_U157;
  assign new_P2_R1179_U354 = ~new_P2_R1179_U183;
  assign new_P2_R1179_U355 = ~new_P2_R1179_U298 | ~new_P2_R1179_U53;
  assign new_P2_R1179_U356 = ~new_P2_R1179_U195 | ~new_P2_R1179_U93;
  assign new_P2_R1179_U357 = ~new_P2_R1179_U139 | ~new_P2_R1179_U356;
  assign new_P2_R1179_U358 = ~new_P2_R1179_U12 | ~new_P2_R1179_U93;
  assign new_P2_R1179_U359 = ~new_P2_R1179_U136 | ~new_P2_R1179_U358;
  assign new_P2_R1179_U360 = ~new_P2_R1179_U12 | ~new_P2_R1179_U93;
  assign new_P2_R1179_U361 = ~new_P2_R1179_U166;
  assign new_P2_R1179_U362 = ~new_P2_U3416 | ~new_P2_R1179_U47;
  assign new_P2_R1179_U363 = ~new_P2_U3082 | ~new_P2_R1179_U46;
  assign new_P2_R1179_U364 = ~new_P2_R1179_U225 | ~new_P2_R1179_U157;
  assign new_P2_R1179_U365 = ~new_P2_R1179_U223 | ~new_P2_R1179_U156;
  assign new_P2_R1179_U366 = ~new_P2_U3413 | ~new_P2_R1179_U28;
  assign new_P2_R1179_U367 = ~new_P2_U3083 | ~new_P2_R1179_U33;
  assign new_P2_R1179_U368 = ~new_P2_U3413 | ~new_P2_R1179_U28;
  assign new_P2_R1179_U369 = ~new_P2_U3083 | ~new_P2_R1179_U33;
  assign new_P2_R1179_U370 = ~new_P2_R1179_U369 | ~new_P2_R1179_U368;
  assign new_P2_R1179_U371 = ~new_P2_U3410 | ~new_P2_R1179_U26;
  assign new_P2_R1179_U372 = ~new_P2_U3069 | ~new_P2_R1179_U32;
  assign new_P2_R1179_U373 = ~new_P2_R1179_U230 | ~new_P2_R1179_U48;
  assign new_P2_R1179_U374 = ~new_P2_R1179_U158 | ~new_P2_R1179_U219;
  assign new_P2_R1179_U375 = ~new_P2_U3407 | ~new_P2_R1179_U41;
  assign new_P2_R1179_U376 = ~new_P2_U3070 | ~new_P2_R1179_U30;
  assign new_P2_R1179_U377 = ~new_P2_R1179_U376 | ~new_P2_R1179_U375;
  assign new_P2_R1179_U378 = ~new_P2_U3404 | ~new_P2_R1179_U42;
  assign new_P2_R1179_U379 = ~new_P2_U3066 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U380 = ~new_P2_R1179_U240 | ~new_P2_R1179_U49;
  assign new_P2_R1179_U381 = ~new_P2_R1179_U159 | ~new_P2_R1179_U232;
  assign new_P2_R1179_U382 = ~new_P2_U3401 | ~new_P2_R1179_U43;
  assign new_P2_R1179_U383 = ~new_P2_U3059 | ~new_P2_R1179_U31;
  assign new_P2_R1179_U384 = ~new_P2_R1179_U161 | ~new_P2_R1179_U241;
  assign new_P2_R1179_U385 = ~new_P2_R1179_U345 | ~new_P2_R1179_U160;
  assign new_P2_R1179_U386 = ~new_P2_U3398 | ~new_P2_R1179_U36;
  assign new_P2_R1179_U387 = ~new_P2_U3063 | ~new_P2_R1179_U40;
  assign new_P2_R1179_U388 = ~new_P2_U3398 | ~new_P2_R1179_U36;
  assign new_P2_R1179_U389 = ~new_P2_U3063 | ~new_P2_R1179_U40;
  assign new_P2_R1179_U390 = ~new_P2_R1179_U389 | ~new_P2_R1179_U388;
  assign new_P2_R1179_U391 = ~new_P2_U3395 | ~new_P2_R1179_U34;
  assign new_P2_R1179_U392 = ~new_P2_U3067 | ~new_P2_R1179_U37;
  assign new_P2_R1179_U393 = ~new_P2_R1179_U243 | ~new_P2_R1179_U50;
  assign new_P2_R1179_U394 = ~new_P2_R1179_U162 | ~new_P2_R1179_U205;
  assign new_P2_R1179_U395 = ~new_P2_U3904 | ~new_P2_R1179_U164;
  assign new_P2_R1179_U396 = ~new_P2_U3054 | ~new_P2_R1179_U163;
  assign new_P2_R1179_U397 = ~new_P2_R1179_U396 | ~new_P2_R1179_U395;
  assign new_P2_R1179_U398 = ~new_P2_U3904 | ~new_P2_R1179_U164;
  assign new_P2_R1179_U399 = ~new_P2_U3054 | ~new_P2_R1179_U163;
  assign new_P2_R1179_U400 = ~new_P2_R1179_U51 | ~new_P2_U3053 | ~new_P2_R1179_U397;
  assign new_P2_R1179_U401 = ~new_P2_U3895 | ~new_P2_R1179_U16 | ~new_P2_R1179_U92;
  assign new_P2_R1179_U402 = ~new_P2_U3895 | ~new_P2_R1179_U92;
  assign new_P2_R1179_U403 = ~new_P2_U3053 | ~new_P2_R1179_U51;
  assign new_P2_R1179_U404 = ~new_P2_R1179_U138;
  assign new_P2_R1179_U405 = ~new_P2_R1179_U361 | ~new_P2_R1179_U404;
  assign new_P2_R1179_U406 = ~new_P2_R1179_U138 | ~new_P2_R1179_U166;
  assign new_P2_R1179_U407 = ~new_P2_U3896 | ~new_P2_R1179_U54;
  assign new_P2_R1179_U408 = ~new_P2_U3052 | ~new_P2_R1179_U91;
  assign new_P2_R1179_U409 = ~new_P2_U3896 | ~new_P2_R1179_U54;
  assign new_P2_R1179_U410 = ~new_P2_U3052 | ~new_P2_R1179_U91;
  assign new_P2_R1179_U411 = ~new_P2_R1179_U410 | ~new_P2_R1179_U409;
  assign new_P2_R1179_U412 = ~new_P2_U3897 | ~new_P2_R1179_U52;
  assign new_P2_R1179_U413 = ~new_P2_U3056 | ~new_P2_R1179_U90;
  assign new_P2_R1179_U414 = ~new_P2_R1179_U306 | ~new_P2_R1179_U93;
  assign new_P2_R1179_U415 = ~new_P2_R1179_U167 | ~new_P2_R1179_U298;
  assign new_P2_R1179_U416 = ~new_P2_U3898 | ~new_P2_R1179_U89;
  assign new_P2_R1179_U417 = ~new_P2_U3057 | ~new_P2_R1179_U88;
  assign new_P2_R1179_U418 = ~new_P2_R1179_U141;
  assign new_P2_R1179_U419 = ~new_P2_R1179_U294 | ~new_P2_R1179_U418;
  assign new_P2_R1179_U420 = ~new_P2_R1179_U141 | ~new_P2_R1179_U168;
  assign new_P2_R1179_U421 = ~new_P2_U3899 | ~new_P2_R1179_U87;
  assign new_P2_R1179_U422 = ~new_P2_U3064 | ~new_P2_R1179_U86;
  assign new_P2_R1179_U423 = ~new_P2_R1179_U142;
  assign new_P2_R1179_U424 = ~new_P2_R1179_U290 | ~new_P2_R1179_U423;
  assign new_P2_R1179_U425 = ~new_P2_R1179_U142 | ~new_P2_R1179_U169;
  assign new_P2_R1179_U426 = ~new_P2_U3900 | ~new_P2_R1179_U82;
  assign new_P2_R1179_U427 = ~new_P2_U3065 | ~new_P2_R1179_U79;
  assign new_P2_R1179_U428 = ~new_P2_R1179_U427 | ~new_P2_R1179_U426;
  assign new_P2_R1179_U429 = ~new_P2_U3901 | ~new_P2_R1179_U83;
  assign new_P2_R1179_U430 = ~new_P2_U3060 | ~new_P2_R1179_U80;
  assign new_P2_R1179_U431 = ~new_P2_R1179_U316 | ~new_P2_R1179_U94;
  assign new_P2_R1179_U432 = ~new_P2_R1179_U170 | ~new_P2_R1179_U308;
  assign new_P2_R1179_U433 = ~new_P2_U3902 | ~new_P2_R1179_U84;
  assign new_P2_R1179_U434 = ~new_P2_U3074 | ~new_P2_R1179_U81;
  assign new_P2_R1179_U435 = ~new_P2_R1179_U317 | ~new_P2_R1179_U172;
  assign new_P2_R1179_U436 = ~new_P2_R1179_U280 | ~new_P2_R1179_U171;
  assign new_P2_R1179_U437 = ~new_P2_U3903 | ~new_P2_R1179_U78;
  assign new_P2_R1179_U438 = ~new_P2_U3075 | ~new_P2_R1179_U77;
  assign new_P2_R1179_U439 = ~new_P2_R1179_U145;
  assign new_P2_R1179_U440 = ~new_P2_R1179_U276 | ~new_P2_R1179_U439;
  assign new_P2_R1179_U441 = ~new_P2_R1179_U145 | ~new_P2_R1179_U173;
  assign new_P2_R1179_U442 = ~new_P2_U3392 | ~new_P2_R1179_U39;
  assign new_P2_R1179_U443 = ~new_P2_U3077 | ~new_P2_R1179_U174;
  assign new_P2_R1179_U444 = ~new_P2_R1179_U146;
  assign new_P2_R1179_U445 = ~new_P2_R1179_U203 | ~new_P2_R1179_U444;
  assign new_P2_R1179_U446 = ~new_P2_R1179_U146 | ~new_P2_R1179_U175;
  assign new_P2_R1179_U447 = ~new_P2_U3445 | ~new_P2_R1179_U76;
  assign new_P2_R1179_U448 = ~new_P2_U3080 | ~new_P2_R1179_U75;
  assign new_P2_R1179_U449 = ~new_P2_R1179_U147;
  assign new_P2_R1179_U450 = ~new_P2_R1179_U272 | ~new_P2_R1179_U449;
  assign new_P2_R1179_U451 = ~new_P2_R1179_U147 | ~new_P2_R1179_U176;
  assign new_P2_R1179_U452 = ~new_P2_U3443 | ~new_P2_R1179_U74;
  assign new_P2_R1179_U453 = ~new_P2_U3081 | ~new_P2_R1179_U177;
  assign new_P2_R1179_U454 = ~new_P2_R1179_U148;
  assign new_P2_R1179_U455 = ~new_P2_R1179_U270 | ~new_P2_R1179_U454;
  assign new_P2_R1179_U456 = ~new_P2_R1179_U148 | ~new_P2_R1179_U178;
  assign new_P2_R1179_U457 = ~new_P2_U3440 | ~new_P2_R1179_U73;
  assign new_P2_R1179_U458 = ~new_P2_U3068 | ~new_P2_R1179_U72;
  assign new_P2_R1179_U459 = ~new_P2_R1179_U149;
  assign new_P2_R1179_U460 = ~new_P2_R1179_U266 | ~new_P2_R1179_U459;
  assign new_P2_R1179_U461 = ~new_P2_R1179_U149 | ~new_P2_R1179_U179;
  assign new_P2_R1179_U462 = ~new_P2_U3437 | ~new_P2_R1179_U68;
  assign new_P2_R1179_U463 = ~new_P2_U3072 | ~new_P2_R1179_U65;
  assign new_P2_R1179_U464 = ~new_P2_R1179_U463 | ~new_P2_R1179_U462;
  assign new_P2_R1179_U465 = ~new_P2_U3434 | ~new_P2_R1179_U69;
  assign new_P2_R1179_U466 = ~new_P2_U3073 | ~new_P2_R1179_U66;
  assign new_P2_R1179_U467 = ~new_P2_R1179_U327 | ~new_P2_R1179_U95;
  assign new_P2_R1179_U468 = ~new_P2_R1179_U180 | ~new_P2_R1179_U319;
  assign new_P2_R1179_U469 = ~new_P2_U3431 | ~new_P2_R1179_U70;
  assign new_P2_R1179_U470 = ~new_P2_U3078 | ~new_P2_R1179_U67;
  assign new_P2_R1179_U471 = ~new_P2_R1179_U328 | ~new_P2_R1179_U182;
  assign new_P2_R1179_U472 = ~new_P2_R1179_U256 | ~new_P2_R1179_U181;
  assign new_P2_R1179_U473 = ~new_P2_U3428 | ~new_P2_R1179_U64;
  assign new_P2_R1179_U474 = ~new_P2_U3079 | ~new_P2_R1179_U63;
  assign new_P2_R1179_U475 = ~new_P2_R1179_U152;
  assign new_P2_R1179_U476 = ~new_P2_R1179_U354 | ~new_P2_R1179_U475;
  assign new_P2_R1179_U477 = ~new_P2_R1179_U152 | ~new_P2_R1179_U183;
  assign new_P2_R1179_U478 = ~new_P2_U3425 | ~new_P2_R1179_U55;
  assign new_P2_R1179_U479 = ~new_P2_U3071 | ~new_P2_R1179_U61;
  assign new_P2_R1179_U480 = ~new_P2_R1179_U153;
  assign new_P2_R1179_U481 = ~new_P2_R1179_U352 | ~new_P2_R1179_U480;
  assign new_P2_R1179_U482 = ~new_P2_R1179_U153 | ~new_P2_R1179_U184;
  assign new_P2_R1179_U483 = ~new_P2_U3422 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U484 = ~new_P2_U3062 | ~new_P2_R1179_U60;
  assign new_P2_R1179_U485 = ~new_P2_R1179_U484 | ~new_P2_R1179_U483;
  assign new_P2_R1179_U486 = ~new_P2_U3419 | ~new_P2_R1179_U57;
  assign new_P2_R1179_U487 = ~new_P2_U3061 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U488 = ~new_P2_R1179_U96 | ~new_P2_R1179_U336;
  assign new_P2_R1179_U489 = ~new_P2_R1179_U185 | ~new_P2_R1179_U350;
  assign new_P2_R1269_U6 = new_P2_R1269_U130 & new_P2_R1269_U131;
  assign new_P2_R1269_U7 = new_P2_R1269_U132 & new_P2_R1269_U133;
  assign new_P2_R1269_U8 = new_P2_R1269_U7 & new_P2_R1269_U137 & new_P2_R1269_U91 & new_P2_R1269_U135;
  assign new_P2_R1269_U9 = new_P2_R1269_U144 & new_P2_R1269_U145;
  assign new_P2_R1269_U10 = new_P2_R1269_U147 & new_P2_R1269_U146;
  assign new_P2_R1269_U11 = new_P2_R1269_U95 & new_P2_R1269_U94 & new_P2_R1269_U148;
  assign new_P2_R1269_U12 = new_P2_R1269_U96 & new_P2_R1269_U11;
  assign new_P2_R1269_U13 = new_P2_R1269_U163 & new_P2_R1269_U162;
  assign new_P2_R1269_U14 = new_P2_R1269_U21 & new_P2_R1269_U20 & new_P2_R1269_U113 & new_P2_R1269_U195 & new_P2_R1269_U191;
  assign new_P2_R1269_U15 = new_P2_R1269_U129 & new_P2_R1269_U128;
  assign new_P2_R1269_U16 = new_P2_R1269_U21 & new_P2_R1269_U114 & new_P2_R1269_U20;
  assign new_P2_R1269_U17 = new_P2_R1269_U21 & new_P2_R1269_U115 & new_P2_R1269_U20;
  assign new_P2_R1269_U18 = new_P2_R1269_U117 & new_P2_R1269_U21;
  assign new_P2_R1269_U19 = new_P2_R1269_U118 & new_P2_R1269_U21;
  assign new_P2_R1269_U20 = new_P2_R1269_U123 & new_P2_R1269_U124 & new_P2_R1269_U125;
  assign new_P2_R1269_U21 = new_P2_R1269_U207 & new_P2_R1269_U206;
  assign new_P2_R1269_U22 = ~new_P2_R1269_U120 | ~new_P2_R1269_U119 | ~new_P2_R1269_U200 | ~new_P2_R1269_U127;
  assign new_P2_R1269_U23 = ~new_P2_U3085;
  assign new_P2_R1269_U24 = ~new_P2_U3084;
  assign new_P2_R1269_U25 = ~new_P2_U3116;
  assign new_P2_R1269_U26 = ~new_P2_U3118;
  assign new_P2_R1269_U27 = ~new_P2_U3117;
  assign new_P2_R1269_U28 = ~new_P2_U3086;
  assign new_P2_R1269_U29 = ~new_P2_U3124;
  assign new_P2_R1269_U30 = ~new_P2_U3123;
  assign new_P2_R1269_U31 = ~new_P2_U3094;
  assign new_P2_R1269_U32 = ~new_P2_U3127;
  assign new_P2_R1269_U33 = ~new_P2_U3095;
  assign new_P2_R1269_U34 = ~new_P2_U3128;
  assign new_P2_R1269_U35 = ~new_P2_U3129;
  assign new_P2_R1269_U36 = ~new_P2_U3098;
  assign new_P2_R1269_U37 = ~new_P2_U3130;
  assign new_P2_R1269_U38 = ~new_P2_U3099;
  assign new_P2_R1269_U39 = ~new_P2_U3097;
  assign new_P2_R1269_U40 = ~new_P2_U3096;
  assign new_P2_R1269_U41 = ~new_P2_U3131;
  assign new_P2_R1269_U42 = ~new_P2_U3132;
  assign new_P2_R1269_U43 = ~new_P2_U3100;
  assign new_P2_R1269_U44 = ~new_P2_U3101;
  assign new_P2_R1269_U45 = ~new_P2_U3141;
  assign new_P2_R1269_U46 = ~new_P2_U3110;
  assign new_P2_R1269_U47 = ~new_P2_U3107;
  assign new_P2_R1269_U48 = ~new_P2_U3106;
  assign new_P2_R1269_U49 = ~new_P2_U3142;
  assign new_P2_R1269_U50 = ~new_P2_U3111;
  assign new_P2_R1269_U51 = ~new_P2_U3109;
  assign new_P2_R1269_U52 = ~new_P2_U3108;
  assign new_P2_R1269_U53 = ~new_P2_U3112;
  assign new_P2_R1269_U54 = ~new_P2_U3113;
  assign new_P2_R1269_U55 = ~new_P2_U3114;
  assign new_P2_R1269_U56 = ~new_P2_U3136;
  assign new_P2_R1269_U57 = ~new_P2_U3135;
  assign new_P2_R1269_U58 = ~new_P2_U3139;
  assign new_P2_R1269_U59 = ~new_P2_U3140;
  assign new_P2_R1269_U60 = ~new_P2_U3146;
  assign new_P2_R1269_U61 = ~new_P2_U3145;
  assign new_P2_R1269_U62 = ~new_P2_U3143;
  assign new_P2_R1269_U63 = ~new_P2_U3144;
  assign new_P2_R1269_U64 = ~new_P2_U3138;
  assign new_P2_R1269_U65 = ~new_P2_U3137;
  assign new_P2_R1269_U66 = ~new_P2_U3104;
  assign new_P2_R1269_U67 = ~new_P2_U3105;
  assign new_P2_R1269_U68 = ~new_P2_U3102;
  assign new_P2_R1269_U69 = ~new_P2_U3103;
  assign new_P2_R1269_U70 = ~new_P2_U3134;
  assign new_P2_R1269_U71 = ~new_P2_U3133;
  assign new_P2_R1269_U72 = ~new_P2_U3126;
  assign new_P2_R1269_U73 = ~new_P2_U3125;
  assign new_P2_R1269_U74 = ~new_P2_U3093;
  assign new_P2_R1269_U75 = ~new_P2_U3092;
  assign new_P2_R1269_U76 = ~new_P2_U3090;
  assign new_P2_R1269_U77 = ~new_P2_U3091;
  assign new_P2_R1269_U78 = ~new_P2_U3087;
  assign new_P2_R1269_U79 = ~new_P2_U3089;
  assign new_P2_R1269_U80 = ~new_P2_U3088;
  assign new_P2_R1269_U81 = ~new_P2_U3122;
  assign new_P2_R1269_U82 = ~new_P2_U3121;
  assign new_P2_R1269_U83 = ~new_P2_U3120;
  assign new_P2_R1269_U84 = ~new_P2_U3119;
  assign new_P2_R1269_U85 = new_P2_R1269_U28 & new_P2_U3118;
  assign new_P2_R1269_U86 = new_P2_U3127 & new_P2_R1269_U33;
  assign new_P2_R1269_U87 = new_P2_U3128 & new_P2_R1269_U40;
  assign new_P2_R1269_U88 = new_P2_R1269_U183 & new_P2_R1269_U182;
  assign new_P2_R1269_U89 = new_P2_U3098 & new_P2_R1269_U37;
  assign new_P2_R1269_U90 = new_P2_U3099 & new_P2_R1269_U41;
  assign new_P2_R1269_U91 = new_P2_R1269_U136 & new_P2_R1269_U134;
  assign new_P2_R1269_U92 = new_P2_U3110 & new_P2_R1269_U49;
  assign new_P2_R1269_U93 = new_P2_U3111 & new_P2_R1269_U62;
  assign new_P2_R1269_U94 = new_P2_R1269_U149 & new_P2_R1269_U143;
  assign new_P2_R1269_U95 = new_P2_R1269_U9 & new_P2_R1269_U150;
  assign new_P2_R1269_U96 = new_P2_R1269_U152 & new_P2_R1269_U151;
  assign new_P2_R1269_U97 = new_P2_R1269_U154 & new_P2_R1269_U155 & new_P2_R1269_U156;
  assign new_P2_R1269_U98 = new_P2_U3139 & new_P2_R1269_U47;
  assign new_P2_R1269_U99 = new_P2_U3140 & new_P2_R1269_U52;
  assign new_P2_R1269_U100 = new_P2_U3146 & new_P2_R1269_U55;
  assign new_P2_R1269_U101 = new_P2_U3145 & new_P2_R1269_U54;
  assign new_P2_R1269_U102 = new_P2_R1269_U13 & new_P2_R1269_U103;
  assign new_P2_R1269_U103 = new_P2_R1269_U168 & new_P2_R1269_U169;
  assign new_P2_R1269_U104 = new_P2_R1269_U167 & new_P2_R1269_U102;
  assign new_P2_R1269_U105 = new_P2_U3104 & new_P2_R1269_U56;
  assign new_P2_R1269_U106 = new_P2_U3105 & new_P2_R1269_U65;
  assign new_P2_R1269_U107 = new_P2_R1269_U172 & new_P2_R1269_U109;
  assign new_P2_R1269_U108 = new_P2_R1269_U107 & new_P2_R1269_U173;
  assign new_P2_R1269_U109 = new_P2_R1269_U175 & new_P2_R1269_U174;
  assign new_P2_R1269_U110 = new_P2_R1269_U139 & new_P2_R1269_U186 & new_P2_R1269_U185;
  assign new_P2_R1269_U111 = new_P2_R1269_U190 & new_P2_R1269_U189;
  assign new_P2_R1269_U112 = new_P2_U3093 & new_P2_R1269_U73;
  assign new_P2_R1269_U113 = new_P2_R1269_U197 & new_P2_R1269_U196;
  assign new_P2_R1269_U114 = new_P2_U3122 & new_P2_R1269_U76;
  assign new_P2_R1269_U115 = new_P2_U3121 & new_P2_R1269_U79;
  assign new_P2_R1269_U116 = new_P2_U3120 & new_P2_R1269_U80;
  assign new_P2_R1269_U117 = new_P2_R1269_U116 & new_P2_R1269_U123;
  assign new_P2_R1269_U118 = new_P2_U3119 & new_P2_R1269_U78;
  assign new_P2_R1269_U119 = new_P2_R1269_U202 & new_P2_R1269_U201;
  assign new_P2_R1269_U120 = new_P2_R1269_U15 & new_P2_R1269_U204 & new_P2_R1269_U203;
  assign new_P2_R1269_U121 = ~new_P2_R1269_U199 | ~new_P2_R1269_U198;
  assign new_P2_R1269_U122 = ~new_P2_U3086 | ~new_P2_R1269_U26;
  assign new_P2_R1269_U123 = ~new_P2_U3087 | ~new_P2_R1269_U84;
  assign new_P2_R1269_U124 = ~new_P2_U3089 | ~new_P2_R1269_U82;
  assign new_P2_R1269_U125 = ~new_P2_U3088 | ~new_P2_R1269_U83;
  assign new_P2_R1269_U126 = ~new_P2_U3085 | ~new_P2_R1269_U27;
  assign new_P2_R1269_U127 = ~new_P2_R1269_U126 | ~new_P2_R1269_U85 | ~new_P2_R1269_U21;
  assign new_P2_R1269_U128 = ~new_P2_R1269_U205 | ~new_P2_R1269_U209 | ~new_P2_R1269_U208;
  assign new_P2_R1269_U129 = ~new_P2_U3117 | ~new_P2_R1269_U21 | ~new_P2_R1269_U23;
  assign new_P2_R1269_U130 = ~new_P2_U3129 | ~new_P2_R1269_U39;
  assign new_P2_R1269_U131 = ~new_P2_U3130 | ~new_P2_R1269_U36;
  assign new_P2_R1269_U132 = ~new_P2_U3094 | ~new_P2_R1269_U72;
  assign new_P2_R1269_U133 = ~new_P2_U3095 | ~new_P2_R1269_U32;
  assign new_P2_R1269_U134 = ~new_P2_R1269_U89 | ~new_P2_R1269_U130;
  assign new_P2_R1269_U135 = ~new_P2_R1269_U90 | ~new_P2_R1269_U6;
  assign new_P2_R1269_U136 = ~new_P2_U3097 | ~new_P2_R1269_U35;
  assign new_P2_R1269_U137 = ~new_P2_U3096 | ~new_P2_R1269_U34;
  assign new_P2_R1269_U138 = ~new_P2_U3100 | ~new_P2_R1269_U42;
  assign new_P2_R1269_U139 = ~new_P2_U3124 | ~new_P2_R1269_U75;
  assign new_P2_R1269_U140 = ~new_P2_U3123 | ~new_P2_R1269_U77;
  assign new_P2_R1269_U141 = ~new_P2_U3101 | ~new_P2_R1269_U71;
  assign new_P2_R1269_U142 = ~new_P2_U3141 | ~new_P2_R1269_U51;
  assign new_P2_R1269_U143 = ~new_P2_R1269_U92 | ~new_P2_R1269_U142;
  assign new_P2_R1269_U144 = ~new_P2_U3106 | ~new_P2_R1269_U64;
  assign new_P2_R1269_U145 = ~new_P2_U3107 | ~new_P2_R1269_U58;
  assign new_P2_R1269_U146 = ~new_P2_U3142 | ~new_P2_R1269_U46;
  assign new_P2_R1269_U147 = ~new_P2_U3141 | ~new_P2_R1269_U51;
  assign new_P2_R1269_U148 = ~new_P2_R1269_U93 | ~new_P2_R1269_U10;
  assign new_P2_R1269_U149 = ~new_P2_U3109 | ~new_P2_R1269_U45;
  assign new_P2_R1269_U150 = ~new_P2_U3108 | ~new_P2_R1269_U59;
  assign new_P2_R1269_U151 = ~new_P2_U3112 | ~new_P2_R1269_U63;
  assign new_P2_R1269_U152 = ~new_P2_U3113 | ~new_P2_R1269_U61;
  assign new_P2_R1269_U153 = ~new_P2_U3147 | ~new_P2_U3148;
  assign new_P2_R1269_U154 = ~new_P2_U3115 | ~new_P2_R1269_U153;
  assign new_P2_R1269_U155 = new_P2_U3147 | new_P2_U3148;
  assign new_P2_R1269_U156 = ~new_P2_U3114 | ~new_P2_R1269_U60;
  assign new_P2_R1269_U157 = ~new_P2_R1269_U97 | ~new_P2_R1269_U12;
  assign new_P2_R1269_U158 = ~new_P2_R1269_U101 | ~new_P2_R1269_U151;
  assign new_P2_R1269_U159 = ~new_P2_U3143 | ~new_P2_R1269_U50;
  assign new_P2_R1269_U160 = ~new_P2_U3144 | ~new_P2_R1269_U53;
  assign new_P2_R1269_U161 = ~new_P2_R1269_U158 | ~new_P2_R1269_U159 | ~new_P2_R1269_U10 | ~new_P2_R1269_U160;
  assign new_P2_R1269_U162 = ~new_P2_U3136 | ~new_P2_R1269_U66;
  assign new_P2_R1269_U163 = ~new_P2_U3135 | ~new_P2_R1269_U69;
  assign new_P2_R1269_U164 = ~new_P2_R1269_U98 | ~new_P2_R1269_U144;
  assign new_P2_R1269_U165 = ~new_P2_R1269_U99 | ~new_P2_R1269_U9;
  assign new_P2_R1269_U166 = ~new_P2_R1269_U100 | ~new_P2_R1269_U12;
  assign new_P2_R1269_U167 = ~new_P2_R1269_U11 | ~new_P2_R1269_U161;
  assign new_P2_R1269_U168 = ~new_P2_U3138 | ~new_P2_R1269_U48;
  assign new_P2_R1269_U169 = ~new_P2_U3137 | ~new_P2_R1269_U67;
  assign new_P2_R1269_U170 = ~new_P2_R1269_U104 | ~new_P2_R1269_U157 | ~new_P2_R1269_U164 | ~new_P2_R1269_U166 | ~new_P2_R1269_U165;
  assign new_P2_R1269_U171 = ~new_P2_U3135 | ~new_P2_R1269_U69;
  assign new_P2_R1269_U172 = ~new_P2_R1269_U105 | ~new_P2_R1269_U171;
  assign new_P2_R1269_U173 = ~new_P2_R1269_U106 | ~new_P2_R1269_U13;
  assign new_P2_R1269_U174 = ~new_P2_U3102 | ~new_P2_R1269_U70;
  assign new_P2_R1269_U175 = ~new_P2_U3103 | ~new_P2_R1269_U57;
  assign new_P2_R1269_U176 = ~new_P2_R1269_U170 | ~new_P2_R1269_U108;
  assign new_P2_R1269_U177 = ~new_P2_U3134 | ~new_P2_R1269_U68;
  assign new_P2_R1269_U178 = ~new_P2_R1269_U177 | ~new_P2_R1269_U176;
  assign new_P2_R1269_U179 = ~new_P2_R1269_U178 | ~new_P2_R1269_U141;
  assign new_P2_R1269_U180 = ~new_P2_U3133 | ~new_P2_R1269_U44;
  assign new_P2_R1269_U181 = ~new_P2_R1269_U180 | ~new_P2_R1269_U179;
  assign new_P2_R1269_U182 = ~new_P2_U3131 | ~new_P2_R1269_U38;
  assign new_P2_R1269_U183 = ~new_P2_U3132 | ~new_P2_R1269_U43;
  assign new_P2_R1269_U184 = ~new_P2_R1269_U88 | ~new_P2_R1269_U6;
  assign new_P2_R1269_U185 = ~new_P2_R1269_U86 | ~new_P2_R1269_U132;
  assign new_P2_R1269_U186 = ~new_P2_R1269_U87 | ~new_P2_R1269_U7;
  assign new_P2_R1269_U187 = ~new_P2_R1269_U8 | ~new_P2_R1269_U184;
  assign new_P2_R1269_U188 = ~new_P2_R1269_U8 | ~new_P2_R1269_U181 | ~new_P2_R1269_U138;
  assign new_P2_R1269_U189 = ~new_P2_U3126 | ~new_P2_R1269_U31;
  assign new_P2_R1269_U190 = ~new_P2_U3125 | ~new_P2_R1269_U74;
  assign new_P2_R1269_U191 = ~new_P2_R1269_U140 | ~new_P2_R1269_U110 | ~new_P2_R1269_U111 | ~new_P2_R1269_U188 | ~new_P2_R1269_U187;
  assign new_P2_R1269_U192 = ~new_P2_R1269_U112 | ~new_P2_R1269_U139;
  assign new_P2_R1269_U193 = ~new_P2_U3092 | ~new_P2_R1269_U29;
  assign new_P2_R1269_U194 = ~new_P2_R1269_U193 | ~new_P2_R1269_U192;
  assign new_P2_R1269_U195 = ~new_P2_R1269_U194 | ~new_P2_R1269_U140;
  assign new_P2_R1269_U196 = ~new_P2_U3090 | ~new_P2_R1269_U81;
  assign new_P2_R1269_U197 = ~new_P2_U3091 | ~new_P2_R1269_U30;
  assign new_P2_R1269_U198 = ~new_P2_U3117 | ~new_P2_R1269_U122;
  assign new_P2_R1269_U199 = ~new_P2_R1269_U122 | ~new_P2_R1269_U23;
  assign new_P2_R1269_U200 = ~new_P2_R1269_U14 | ~new_P2_R1269_U121;
  assign new_P2_R1269_U201 = ~new_P2_R1269_U16 | ~new_P2_R1269_U121;
  assign new_P2_R1269_U202 = ~new_P2_R1269_U17 | ~new_P2_R1269_U121;
  assign new_P2_R1269_U203 = ~new_P2_R1269_U18 | ~new_P2_R1269_U121;
  assign new_P2_R1269_U204 = ~new_P2_R1269_U19 | ~new_P2_R1269_U121;
  assign new_P2_R1269_U205 = ~new_P2_U3116 | ~new_P2_U3084;
  assign new_P2_R1269_U206 = ~new_P2_U3084 | ~new_P2_R1269_U25;
  assign new_P2_R1269_U207 = ~new_P2_U3116 | ~new_P2_R1269_U24;
  assign new_P2_R1269_U208 = new_P2_U3149 | new_P2_U3116;
  assign new_P2_R1269_U209 = ~new_P2_U3149 | ~new_P2_R1269_U24;
  assign new_P2_R1110_U4 = new_P2_R1110_U179 & new_P2_R1110_U178;
  assign new_P2_R1110_U5 = new_P2_R1110_U197 & new_P2_R1110_U196;
  assign new_P2_R1110_U6 = new_P2_R1110_U237 & new_P2_R1110_U236;
  assign new_P2_R1110_U7 = new_P2_R1110_U246 & new_P2_R1110_U245;
  assign new_P2_R1110_U8 = new_P2_R1110_U264 & new_P2_R1110_U263;
  assign new_P2_R1110_U9 = new_P2_R1110_U272 & new_P2_R1110_U271;
  assign new_P2_R1110_U10 = new_P2_R1110_U351 & new_P2_R1110_U348;
  assign new_P2_R1110_U11 = new_P2_R1110_U344 & new_P2_R1110_U341;
  assign new_P2_R1110_U12 = new_P2_R1110_U335 & new_P2_R1110_U332;
  assign new_P2_R1110_U13 = new_P2_R1110_U326 & new_P2_R1110_U323;
  assign new_P2_R1110_U14 = new_P2_R1110_U320 & new_P2_R1110_U318;
  assign new_P2_R1110_U15 = new_P2_R1110_U313 & new_P2_R1110_U310;
  assign new_P2_R1110_U16 = new_P2_R1110_U235 & new_P2_R1110_U232;
  assign new_P2_R1110_U17 = new_P2_R1110_U227 & new_P2_R1110_U224;
  assign new_P2_R1110_U18 = new_P2_R1110_U213 & new_P2_R1110_U210;
  assign new_P2_R1110_U19 = ~new_P2_U3407;
  assign new_P2_R1110_U20 = ~new_P2_U3070;
  assign new_P2_R1110_U21 = ~new_P2_U3069;
  assign new_P2_R1110_U22 = ~new_P2_U3070 | ~new_P2_U3407;
  assign new_P2_R1110_U23 = ~new_P2_U3410;
  assign new_P2_R1110_U24 = ~new_P2_U3401;
  assign new_P2_R1110_U25 = ~new_P2_U3059;
  assign new_P2_R1110_U26 = ~new_P2_U3066;
  assign new_P2_R1110_U27 = ~new_P2_U3395;
  assign new_P2_R1110_U28 = ~new_P2_U3067;
  assign new_P2_R1110_U29 = ~new_P2_U3387;
  assign new_P2_R1110_U30 = ~new_P2_U3076;
  assign new_P2_R1110_U31 = ~new_P2_U3076 | ~new_P2_U3387;
  assign new_P2_R1110_U32 = ~new_P2_U3398;
  assign new_P2_R1110_U33 = ~new_P2_U3063;
  assign new_P2_R1110_U34 = ~new_P2_U3059 | ~new_P2_U3401;
  assign new_P2_R1110_U35 = ~new_P2_U3404;
  assign new_P2_R1110_U36 = ~new_P2_U3413;
  assign new_P2_R1110_U37 = ~new_P2_U3083;
  assign new_P2_R1110_U38 = ~new_P2_U3082;
  assign new_P2_R1110_U39 = ~new_P2_U3416;
  assign new_P2_R1110_U40 = ~new_P2_R1110_U65 | ~new_P2_R1110_U205;
  assign new_P2_R1110_U41 = ~new_P2_R1110_U117 | ~new_P2_R1110_U193;
  assign new_P2_R1110_U42 = ~new_P2_R1110_U182 | ~new_P2_R1110_U183;
  assign new_P2_R1110_U43 = ~new_P2_U3392 | ~new_P2_U3077;
  assign new_P2_R1110_U44 = ~new_P2_R1110_U122 | ~new_P2_R1110_U219;
  assign new_P2_R1110_U45 = ~new_P2_R1110_U216 | ~new_P2_R1110_U215;
  assign new_P2_R1110_U46 = ~new_P2_U3896;
  assign new_P2_R1110_U47 = ~new_P2_U3052;
  assign new_P2_R1110_U48 = ~new_P2_U3056;
  assign new_P2_R1110_U49 = ~new_P2_U3897;
  assign new_P2_R1110_U50 = ~new_P2_U3898;
  assign new_P2_R1110_U51 = ~new_P2_U3057;
  assign new_P2_R1110_U52 = ~new_P2_U3899;
  assign new_P2_R1110_U53 = ~new_P2_U3064;
  assign new_P2_R1110_U54 = ~new_P2_U3902;
  assign new_P2_R1110_U55 = ~new_P2_U3074;
  assign new_P2_R1110_U56 = ~new_P2_U3437;
  assign new_P2_R1110_U57 = ~new_P2_U3072;
  assign new_P2_R1110_U58 = ~new_P2_U3068;
  assign new_P2_R1110_U59 = ~new_P2_U3072 | ~new_P2_U3437;
  assign new_P2_R1110_U60 = ~new_P2_U3440;
  assign new_P2_R1110_U61 = ~new_P2_U3428;
  assign new_P2_R1110_U62 = ~new_P2_U3079;
  assign new_P2_R1110_U63 = ~new_P2_U3419;
  assign new_P2_R1110_U64 = ~new_P2_U3061;
  assign new_P2_R1110_U65 = ~new_P2_U3083 | ~new_P2_U3413;
  assign new_P2_R1110_U66 = ~new_P2_U3422;
  assign new_P2_R1110_U67 = ~new_P2_U3062;
  assign new_P2_R1110_U68 = ~new_P2_U3062 | ~new_P2_U3422;
  assign new_P2_R1110_U69 = ~new_P2_U3425;
  assign new_P2_R1110_U70 = ~new_P2_U3071;
  assign new_P2_R1110_U71 = ~new_P2_U3431;
  assign new_P2_R1110_U72 = ~new_P2_U3078;
  assign new_P2_R1110_U73 = ~new_P2_U3434;
  assign new_P2_R1110_U74 = ~new_P2_U3073;
  assign new_P2_R1110_U75 = ~new_P2_U3443;
  assign new_P2_R1110_U76 = ~new_P2_U3081;
  assign new_P2_R1110_U77 = ~new_P2_U3081 | ~new_P2_U3443;
  assign new_P2_R1110_U78 = ~new_P2_U3445;
  assign new_P2_R1110_U79 = ~new_P2_U3080;
  assign new_P2_R1110_U80 = ~new_P2_U3080 | ~new_P2_U3445;
  assign new_P2_R1110_U81 = ~new_P2_U3903;
  assign new_P2_R1110_U82 = ~new_P2_U3901;
  assign new_P2_R1110_U83 = ~new_P2_U3060;
  assign new_P2_R1110_U84 = ~new_P2_U3900;
  assign new_P2_R1110_U85 = ~new_P2_U3065;
  assign new_P2_R1110_U86 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1110_U87 = ~new_P2_U3053;
  assign new_P2_R1110_U88 = ~new_P2_U3895;
  assign new_P2_R1110_U89 = ~new_P2_R1110_U306 | ~new_P2_R1110_U176;
  assign new_P2_R1110_U90 = ~new_P2_U3075;
  assign new_P2_R1110_U91 = ~new_P2_R1110_U77 | ~new_P2_R1110_U315;
  assign new_P2_R1110_U92 = ~new_P2_R1110_U261 | ~new_P2_R1110_U260;
  assign new_P2_R1110_U93 = ~new_P2_R1110_U68 | ~new_P2_R1110_U337;
  assign new_P2_R1110_U94 = ~new_P2_R1110_U457 | ~new_P2_R1110_U456;
  assign new_P2_R1110_U95 = ~new_P2_R1110_U504 | ~new_P2_R1110_U503;
  assign new_P2_R1110_U96 = ~new_P2_R1110_U375 | ~new_P2_R1110_U374;
  assign new_P2_R1110_U97 = ~new_P2_R1110_U380 | ~new_P2_R1110_U379;
  assign new_P2_R1110_U98 = ~new_P2_R1110_U387 | ~new_P2_R1110_U386;
  assign new_P2_R1110_U99 = ~new_P2_R1110_U394 | ~new_P2_R1110_U393;
  assign new_P2_R1110_U100 = ~new_P2_R1110_U399 | ~new_P2_R1110_U398;
  assign new_P2_R1110_U101 = ~new_P2_R1110_U408 | ~new_P2_R1110_U407;
  assign new_P2_R1110_U102 = ~new_P2_R1110_U415 | ~new_P2_R1110_U414;
  assign new_P2_R1110_U103 = ~new_P2_R1110_U422 | ~new_P2_R1110_U421;
  assign new_P2_R1110_U104 = ~new_P2_R1110_U429 | ~new_P2_R1110_U428;
  assign new_P2_R1110_U105 = ~new_P2_R1110_U434 | ~new_P2_R1110_U433;
  assign new_P2_R1110_U106 = ~new_P2_R1110_U441 | ~new_P2_R1110_U440;
  assign new_P2_R1110_U107 = ~new_P2_R1110_U448 | ~new_P2_R1110_U447;
  assign new_P2_R1110_U108 = ~new_P2_R1110_U462 | ~new_P2_R1110_U461;
  assign new_P2_R1110_U109 = ~new_P2_R1110_U467 | ~new_P2_R1110_U466;
  assign new_P2_R1110_U110 = ~new_P2_R1110_U474 | ~new_P2_R1110_U473;
  assign new_P2_R1110_U111 = ~new_P2_R1110_U481 | ~new_P2_R1110_U480;
  assign new_P2_R1110_U112 = ~new_P2_R1110_U488 | ~new_P2_R1110_U487;
  assign new_P2_R1110_U113 = ~new_P2_R1110_U495 | ~new_P2_R1110_U494;
  assign new_P2_R1110_U114 = ~new_P2_R1110_U500 | ~new_P2_R1110_U499;
  assign new_P2_R1110_U115 = new_P2_R1110_U189 & new_P2_R1110_U187;
  assign new_P2_R1110_U116 = new_P2_R1110_U4 & new_P2_R1110_U180;
  assign new_P2_R1110_U117 = new_P2_R1110_U194 & new_P2_R1110_U192;
  assign new_P2_R1110_U118 = new_P2_R1110_U201 & new_P2_R1110_U200;
  assign new_P2_R1110_U119 = new_P2_R1110_U22 & new_P2_R1110_U382 & new_P2_R1110_U381;
  assign new_P2_R1110_U120 = new_P2_R1110_U212 & new_P2_R1110_U5;
  assign new_P2_R1110_U121 = new_P2_R1110_U181 & new_P2_R1110_U180;
  assign new_P2_R1110_U122 = new_P2_R1110_U220 & new_P2_R1110_U218;
  assign new_P2_R1110_U123 = new_P2_R1110_U34 & new_P2_R1110_U389 & new_P2_R1110_U388;
  assign new_P2_R1110_U124 = new_P2_R1110_U226 & new_P2_R1110_U4;
  assign new_P2_R1110_U125 = new_P2_R1110_U234 & new_P2_R1110_U181;
  assign new_P2_R1110_U126 = new_P2_R1110_U204 & new_P2_R1110_U6;
  assign new_P2_R1110_U127 = new_P2_R1110_U243 & new_P2_R1110_U239;
  assign new_P2_R1110_U128 = new_P2_R1110_U250 & new_P2_R1110_U7;
  assign new_P2_R1110_U129 = new_P2_R1110_U253 & new_P2_R1110_U248;
  assign new_P2_R1110_U130 = new_P2_R1110_U268 & new_P2_R1110_U267;
  assign new_P2_R1110_U131 = new_P2_R1110_U9 & new_P2_R1110_U282;
  assign new_P2_R1110_U132 = new_P2_R1110_U285 & new_P2_R1110_U280;
  assign new_P2_R1110_U133 = new_P2_R1110_U301 & new_P2_R1110_U298;
  assign new_P2_R1110_U134 = new_P2_R1110_U368 & new_P2_R1110_U302;
  assign new_P2_R1110_U135 = new_P2_R1110_U160 & new_P2_R1110_U278;
  assign new_P2_R1110_U136 = new_P2_R1110_U80 & new_P2_R1110_U455 & new_P2_R1110_U454;
  assign new_P2_R1110_U137 = new_P2_R1110_U325 & new_P2_R1110_U9;
  assign new_P2_R1110_U138 = new_P2_R1110_U59 & new_P2_R1110_U469 & new_P2_R1110_U468;
  assign new_P2_R1110_U139 = new_P2_R1110_U334 & new_P2_R1110_U8;
  assign new_P2_R1110_U140 = new_P2_R1110_U172 & new_P2_R1110_U490 & new_P2_R1110_U489;
  assign new_P2_R1110_U141 = new_P2_R1110_U343 & new_P2_R1110_U7;
  assign new_P2_R1110_U142 = new_P2_R1110_U171 & new_P2_R1110_U502 & new_P2_R1110_U501;
  assign new_P2_R1110_U143 = new_P2_R1110_U350 & new_P2_R1110_U6;
  assign new_P2_R1110_U144 = ~new_P2_R1110_U118 | ~new_P2_R1110_U202;
  assign new_P2_R1110_U145 = ~new_P2_R1110_U217 | ~new_P2_R1110_U229;
  assign new_P2_R1110_U146 = ~new_P2_U3054;
  assign new_P2_R1110_U147 = ~new_P2_U3904;
  assign new_P2_R1110_U148 = new_P2_R1110_U403 & new_P2_R1110_U402;
  assign new_P2_R1110_U149 = ~new_P2_R1110_U364 | ~new_P2_R1110_U304 | ~new_P2_R1110_U169;
  assign new_P2_R1110_U150 = new_P2_R1110_U410 & new_P2_R1110_U409;
  assign new_P2_R1110_U151 = ~new_P2_R1110_U134 | ~new_P2_R1110_U370 | ~new_P2_R1110_U369;
  assign new_P2_R1110_U152 = new_P2_R1110_U417 & new_P2_R1110_U416;
  assign new_P2_R1110_U153 = ~new_P2_R1110_U86 | ~new_P2_R1110_U365 | ~new_P2_R1110_U299;
  assign new_P2_R1110_U154 = new_P2_R1110_U424 & new_P2_R1110_U423;
  assign new_P2_R1110_U155 = ~new_P2_R1110_U293 | ~new_P2_R1110_U292;
  assign new_P2_R1110_U156 = new_P2_R1110_U436 & new_P2_R1110_U435;
  assign new_P2_R1110_U157 = ~new_P2_R1110_U289 | ~new_P2_R1110_U288;
  assign new_P2_R1110_U158 = new_P2_R1110_U443 & new_P2_R1110_U442;
  assign new_P2_R1110_U159 = ~new_P2_R1110_U132 | ~new_P2_R1110_U284;
  assign new_P2_R1110_U160 = new_P2_R1110_U450 & new_P2_R1110_U449;
  assign new_P2_R1110_U161 = ~new_P2_R1110_U43 | ~new_P2_R1110_U327;
  assign new_P2_R1110_U162 = ~new_P2_R1110_U130 | ~new_P2_R1110_U269;
  assign new_P2_R1110_U163 = new_P2_R1110_U476 & new_P2_R1110_U475;
  assign new_P2_R1110_U164 = ~new_P2_R1110_U257 | ~new_P2_R1110_U256;
  assign new_P2_R1110_U165 = new_P2_R1110_U483 & new_P2_R1110_U482;
  assign new_P2_R1110_U166 = ~new_P2_R1110_U129 | ~new_P2_R1110_U252;
  assign new_P2_R1110_U167 = ~new_P2_R1110_U127 | ~new_P2_R1110_U242;
  assign new_P2_R1110_U168 = ~new_P2_R1110_U367 | ~new_P2_R1110_U366;
  assign new_P2_R1110_U169 = ~new_P2_U3053 | ~new_P2_R1110_U151;
  assign new_P2_R1110_U170 = ~new_P2_R1110_U34;
  assign new_P2_R1110_U171 = ~new_P2_U3416 | ~new_P2_U3082;
  assign new_P2_R1110_U172 = ~new_P2_U3071 | ~new_P2_U3425;
  assign new_P2_R1110_U173 = ~new_P2_U3057 | ~new_P2_U3898;
  assign new_P2_R1110_U174 = ~new_P2_R1110_U68;
  assign new_P2_R1110_U175 = ~new_P2_R1110_U77;
  assign new_P2_R1110_U176 = ~new_P2_U3064 | ~new_P2_U3899;
  assign new_P2_R1110_U177 = ~new_P2_R1110_U65;
  assign new_P2_R1110_U178 = new_P2_U3066 | new_P2_U3404;
  assign new_P2_R1110_U179 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1110_U180 = new_P2_U3398 | new_P2_U3063;
  assign new_P2_R1110_U181 = new_P2_U3395 | new_P2_U3067;
  assign new_P2_R1110_U182 = ~new_P2_R1110_U31;
  assign new_P2_R1110_U183 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1110_U184 = ~new_P2_R1110_U42;
  assign new_P2_R1110_U185 = ~new_P2_R1110_U43;
  assign new_P2_R1110_U186 = ~new_P2_R1110_U42 | ~new_P2_R1110_U43;
  assign new_P2_R1110_U187 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1110_U188 = ~new_P2_R1110_U186 | ~new_P2_R1110_U181;
  assign new_P2_R1110_U189 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1110_U190 = ~new_P2_R1110_U115 | ~new_P2_R1110_U188;
  assign new_P2_R1110_U191 = ~new_P2_R1110_U35 | ~new_P2_R1110_U34;
  assign new_P2_R1110_U192 = ~new_P2_U3066 | ~new_P2_R1110_U191;
  assign new_P2_R1110_U193 = ~new_P2_R1110_U116 | ~new_P2_R1110_U190;
  assign new_P2_R1110_U194 = ~new_P2_U3404 | ~new_P2_R1110_U170;
  assign new_P2_R1110_U195 = ~new_P2_R1110_U41;
  assign new_P2_R1110_U196 = new_P2_U3069 | new_P2_U3410;
  assign new_P2_R1110_U197 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1110_U198 = ~new_P2_R1110_U22;
  assign new_P2_R1110_U199 = ~new_P2_R1110_U23 | ~new_P2_R1110_U22;
  assign new_P2_R1110_U200 = ~new_P2_U3069 | ~new_P2_R1110_U199;
  assign new_P2_R1110_U201 = ~new_P2_U3410 | ~new_P2_R1110_U198;
  assign new_P2_R1110_U202 = ~new_P2_R1110_U5 | ~new_P2_R1110_U41;
  assign new_P2_R1110_U203 = ~new_P2_R1110_U144;
  assign new_P2_R1110_U204 = new_P2_U3413 | new_P2_U3083;
  assign new_P2_R1110_U205 = ~new_P2_R1110_U204 | ~new_P2_R1110_U144;
  assign new_P2_R1110_U206 = ~new_P2_R1110_U40;
  assign new_P2_R1110_U207 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1110_U208 = new_P2_U3407 | new_P2_U3070;
  assign new_P2_R1110_U209 = ~new_P2_R1110_U208 | ~new_P2_R1110_U41;
  assign new_P2_R1110_U210 = ~new_P2_R1110_U119 | ~new_P2_R1110_U209;
  assign new_P2_R1110_U211 = ~new_P2_R1110_U195 | ~new_P2_R1110_U22;
  assign new_P2_R1110_U212 = ~new_P2_U3410 | ~new_P2_U3069;
  assign new_P2_R1110_U213 = ~new_P2_R1110_U120 | ~new_P2_R1110_U211;
  assign new_P2_R1110_U214 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1110_U215 = ~new_P2_R1110_U185 | ~new_P2_R1110_U181;
  assign new_P2_R1110_U216 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1110_U217 = ~new_P2_R1110_U45;
  assign new_P2_R1110_U218 = ~new_P2_R1110_U121 | ~new_P2_R1110_U184;
  assign new_P2_R1110_U219 = ~new_P2_R1110_U45 | ~new_P2_R1110_U180;
  assign new_P2_R1110_U220 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1110_U221 = ~new_P2_R1110_U44;
  assign new_P2_R1110_U222 = new_P2_U3401 | new_P2_U3059;
  assign new_P2_R1110_U223 = ~new_P2_R1110_U222 | ~new_P2_R1110_U44;
  assign new_P2_R1110_U224 = ~new_P2_R1110_U123 | ~new_P2_R1110_U223;
  assign new_P2_R1110_U225 = ~new_P2_R1110_U221 | ~new_P2_R1110_U34;
  assign new_P2_R1110_U226 = ~new_P2_U3404 | ~new_P2_U3066;
  assign new_P2_R1110_U227 = ~new_P2_R1110_U124 | ~new_P2_R1110_U225;
  assign new_P2_R1110_U228 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1110_U229 = ~new_P2_R1110_U184 | ~new_P2_R1110_U181;
  assign new_P2_R1110_U230 = ~new_P2_R1110_U145;
  assign new_P2_R1110_U231 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1110_U232 = ~new_P2_R1110_U42 | ~new_P2_R1110_U43 | ~new_P2_R1110_U401 | ~new_P2_R1110_U400;
  assign new_P2_R1110_U233 = ~new_P2_R1110_U43 | ~new_P2_R1110_U42;
  assign new_P2_R1110_U234 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1110_U235 = ~new_P2_R1110_U125 | ~new_P2_R1110_U233;
  assign new_P2_R1110_U236 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1110_U237 = new_P2_U3061 | new_P2_U3419;
  assign new_P2_R1110_U238 = ~new_P2_R1110_U177 | ~new_P2_R1110_U6;
  assign new_P2_R1110_U239 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1110_U240 = ~new_P2_R1110_U171 | ~new_P2_R1110_U238;
  assign new_P2_R1110_U241 = new_P2_U3419 | new_P2_U3061;
  assign new_P2_R1110_U242 = ~new_P2_R1110_U126 | ~new_P2_R1110_U144;
  assign new_P2_R1110_U243 = ~new_P2_R1110_U241 | ~new_P2_R1110_U240;
  assign new_P2_R1110_U244 = ~new_P2_R1110_U167;
  assign new_P2_R1110_U245 = new_P2_U3079 | new_P2_U3428;
  assign new_P2_R1110_U246 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1110_U247 = ~new_P2_R1110_U174 | ~new_P2_R1110_U7;
  assign new_P2_R1110_U248 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1110_U249 = ~new_P2_R1110_U172 | ~new_P2_R1110_U247;
  assign new_P2_R1110_U250 = new_P2_U3422 | new_P2_U3062;
  assign new_P2_R1110_U251 = new_P2_U3428 | new_P2_U3079;
  assign new_P2_R1110_U252 = ~new_P2_R1110_U128 | ~new_P2_R1110_U167;
  assign new_P2_R1110_U253 = ~new_P2_R1110_U251 | ~new_P2_R1110_U249;
  assign new_P2_R1110_U254 = ~new_P2_R1110_U166;
  assign new_P2_R1110_U255 = new_P2_U3431 | new_P2_U3078;
  assign new_P2_R1110_U256 = ~new_P2_R1110_U255 | ~new_P2_R1110_U166;
  assign new_P2_R1110_U257 = ~new_P2_U3078 | ~new_P2_U3431;
  assign new_P2_R1110_U258 = ~new_P2_R1110_U164;
  assign new_P2_R1110_U259 = new_P2_U3434 | new_P2_U3073;
  assign new_P2_R1110_U260 = ~new_P2_R1110_U259 | ~new_P2_R1110_U164;
  assign new_P2_R1110_U261 = ~new_P2_U3073 | ~new_P2_U3434;
  assign new_P2_R1110_U262 = ~new_P2_R1110_U92;
  assign new_P2_R1110_U263 = new_P2_U3068 | new_P2_U3440;
  assign new_P2_R1110_U264 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1110_U265 = ~new_P2_R1110_U59;
  assign new_P2_R1110_U266 = ~new_P2_R1110_U60 | ~new_P2_R1110_U59;
  assign new_P2_R1110_U267 = ~new_P2_U3068 | ~new_P2_R1110_U266;
  assign new_P2_R1110_U268 = ~new_P2_U3440 | ~new_P2_R1110_U265;
  assign new_P2_R1110_U269 = ~new_P2_R1110_U8 | ~new_P2_R1110_U92;
  assign new_P2_R1110_U270 = ~new_P2_R1110_U162;
  assign new_P2_R1110_U271 = new_P2_U3075 | new_P2_U3903;
  assign new_P2_R1110_U272 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1110_U273 = new_P2_U3074 | new_P2_U3902;
  assign new_P2_R1110_U274 = ~new_P2_R1110_U80;
  assign new_P2_R1110_U275 = ~new_P2_U3903 | ~new_P2_R1110_U274;
  assign new_P2_R1110_U276 = ~new_P2_R1110_U275 | ~new_P2_R1110_U90;
  assign new_P2_R1110_U277 = ~new_P2_R1110_U80 | ~new_P2_R1110_U81;
  assign new_P2_R1110_U278 = ~new_P2_R1110_U277 | ~new_P2_R1110_U276;
  assign new_P2_R1110_U279 = ~new_P2_R1110_U175 | ~new_P2_R1110_U9;
  assign new_P2_R1110_U280 = ~new_P2_U3074 | ~new_P2_U3902;
  assign new_P2_R1110_U281 = ~new_P2_R1110_U278 | ~new_P2_R1110_U279;
  assign new_P2_R1110_U282 = new_P2_U3443 | new_P2_U3081;
  assign new_P2_R1110_U283 = new_P2_U3902 | new_P2_U3074;
  assign new_P2_R1110_U284 = ~new_P2_R1110_U131 | ~new_P2_R1110_U273 | ~new_P2_R1110_U162;
  assign new_P2_R1110_U285 = ~new_P2_R1110_U283 | ~new_P2_R1110_U281;
  assign new_P2_R1110_U286 = ~new_P2_R1110_U159;
  assign new_P2_R1110_U287 = new_P2_U3901 | new_P2_U3060;
  assign new_P2_R1110_U288 = ~new_P2_R1110_U287 | ~new_P2_R1110_U159;
  assign new_P2_R1110_U289 = ~new_P2_U3060 | ~new_P2_U3901;
  assign new_P2_R1110_U290 = ~new_P2_R1110_U157;
  assign new_P2_R1110_U291 = new_P2_U3900 | new_P2_U3065;
  assign new_P2_R1110_U292 = ~new_P2_R1110_U291 | ~new_P2_R1110_U157;
  assign new_P2_R1110_U293 = ~new_P2_U3065 | ~new_P2_U3900;
  assign new_P2_R1110_U294 = ~new_P2_R1110_U155;
  assign new_P2_R1110_U295 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1110_U296 = ~new_P2_R1110_U176 | ~new_P2_R1110_U173;
  assign new_P2_R1110_U297 = ~new_P2_R1110_U86;
  assign new_P2_R1110_U298 = new_P2_U3899 | new_P2_U3064;
  assign new_P2_R1110_U299 = ~new_P2_R1110_U168 | ~new_P2_R1110_U155 | ~new_P2_R1110_U298;
  assign new_P2_R1110_U300 = ~new_P2_R1110_U153;
  assign new_P2_R1110_U301 = new_P2_U3896 | new_P2_U3052;
  assign new_P2_R1110_U302 = ~new_P2_U3052 | ~new_P2_U3896;
  assign new_P2_R1110_U303 = ~new_P2_R1110_U151;
  assign new_P2_R1110_U304 = ~new_P2_U3895 | ~new_P2_R1110_U151;
  assign new_P2_R1110_U305 = ~new_P2_R1110_U149;
  assign new_P2_R1110_U306 = ~new_P2_R1110_U298 | ~new_P2_R1110_U155;
  assign new_P2_R1110_U307 = ~new_P2_R1110_U89;
  assign new_P2_R1110_U308 = new_P2_U3898 | new_P2_U3057;
  assign new_P2_R1110_U309 = ~new_P2_R1110_U308 | ~new_P2_R1110_U89;
  assign new_P2_R1110_U310 = ~new_P2_R1110_U154 | ~new_P2_R1110_U309 | ~new_P2_R1110_U173;
  assign new_P2_R1110_U311 = ~new_P2_R1110_U307 | ~new_P2_R1110_U173;
  assign new_P2_R1110_U312 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1110_U313 = ~new_P2_R1110_U168 | ~new_P2_R1110_U311 | ~new_P2_R1110_U312;
  assign new_P2_R1110_U314 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1110_U315 = ~new_P2_R1110_U282 | ~new_P2_R1110_U162;
  assign new_P2_R1110_U316 = ~new_P2_R1110_U91;
  assign new_P2_R1110_U317 = ~new_P2_R1110_U9 | ~new_P2_R1110_U91;
  assign new_P2_R1110_U318 = ~new_P2_R1110_U135 | ~new_P2_R1110_U317;
  assign new_P2_R1110_U319 = ~new_P2_R1110_U317 | ~new_P2_R1110_U278;
  assign new_P2_R1110_U320 = ~new_P2_R1110_U453 | ~new_P2_R1110_U319;
  assign new_P2_R1110_U321 = new_P2_U3445 | new_P2_U3080;
  assign new_P2_R1110_U322 = ~new_P2_R1110_U321 | ~new_P2_R1110_U91;
  assign new_P2_R1110_U323 = ~new_P2_R1110_U136 | ~new_P2_R1110_U322;
  assign new_P2_R1110_U324 = ~new_P2_R1110_U316 | ~new_P2_R1110_U80;
  assign new_P2_R1110_U325 = ~new_P2_U3075 | ~new_P2_U3903;
  assign new_P2_R1110_U326 = ~new_P2_R1110_U137 | ~new_P2_R1110_U324;
  assign new_P2_R1110_U327 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1110_U328 = ~new_P2_R1110_U161;
  assign new_P2_R1110_U329 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1110_U330 = new_P2_U3437 | new_P2_U3072;
  assign new_P2_R1110_U331 = ~new_P2_R1110_U330 | ~new_P2_R1110_U92;
  assign new_P2_R1110_U332 = ~new_P2_R1110_U138 | ~new_P2_R1110_U331;
  assign new_P2_R1110_U333 = ~new_P2_R1110_U262 | ~new_P2_R1110_U59;
  assign new_P2_R1110_U334 = ~new_P2_U3440 | ~new_P2_U3068;
  assign new_P2_R1110_U335 = ~new_P2_R1110_U139 | ~new_P2_R1110_U333;
  assign new_P2_R1110_U336 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1110_U337 = ~new_P2_R1110_U250 | ~new_P2_R1110_U167;
  assign new_P2_R1110_U338 = ~new_P2_R1110_U93;
  assign new_P2_R1110_U339 = new_P2_U3425 | new_P2_U3071;
  assign new_P2_R1110_U340 = ~new_P2_R1110_U339 | ~new_P2_R1110_U93;
  assign new_P2_R1110_U341 = ~new_P2_R1110_U140 | ~new_P2_R1110_U340;
  assign new_P2_R1110_U342 = ~new_P2_R1110_U338 | ~new_P2_R1110_U172;
  assign new_P2_R1110_U343 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1110_U344 = ~new_P2_R1110_U141 | ~new_P2_R1110_U342;
  assign new_P2_R1110_U345 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1110_U346 = new_P2_U3416 | new_P2_U3082;
  assign new_P2_R1110_U347 = ~new_P2_R1110_U346 | ~new_P2_R1110_U40;
  assign new_P2_R1110_U348 = ~new_P2_R1110_U142 | ~new_P2_R1110_U347;
  assign new_P2_R1110_U349 = ~new_P2_R1110_U206 | ~new_P2_R1110_U171;
  assign new_P2_R1110_U350 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1110_U351 = ~new_P2_R1110_U143 | ~new_P2_R1110_U349;
  assign new_P2_R1110_U352 = ~new_P2_R1110_U207 | ~new_P2_R1110_U171;
  assign new_P2_R1110_U353 = ~new_P2_R1110_U204 | ~new_P2_R1110_U65;
  assign new_P2_R1110_U354 = ~new_P2_R1110_U214 | ~new_P2_R1110_U22;
  assign new_P2_R1110_U355 = ~new_P2_R1110_U228 | ~new_P2_R1110_U34;
  assign new_P2_R1110_U356 = ~new_P2_R1110_U231 | ~new_P2_R1110_U180;
  assign new_P2_R1110_U357 = ~new_P2_R1110_U314 | ~new_P2_R1110_U173;
  assign new_P2_R1110_U358 = ~new_P2_R1110_U298 | ~new_P2_R1110_U176;
  assign new_P2_R1110_U359 = ~new_P2_R1110_U329 | ~new_P2_R1110_U80;
  assign new_P2_R1110_U360 = ~new_P2_R1110_U282 | ~new_P2_R1110_U77;
  assign new_P2_R1110_U361 = ~new_P2_R1110_U336 | ~new_P2_R1110_U59;
  assign new_P2_R1110_U362 = ~new_P2_R1110_U345 | ~new_P2_R1110_U172;
  assign new_P2_R1110_U363 = ~new_P2_R1110_U250 | ~new_P2_R1110_U68;
  assign new_P2_R1110_U364 = ~new_P2_U3895 | ~new_P2_U3053;
  assign new_P2_R1110_U365 = ~new_P2_R1110_U296 | ~new_P2_R1110_U168;
  assign new_P2_R1110_U366 = ~new_P2_U3056 | ~new_P2_R1110_U295;
  assign new_P2_R1110_U367 = ~new_P2_U3897 | ~new_P2_R1110_U295;
  assign new_P2_R1110_U368 = ~new_P2_R1110_U301 | ~new_P2_R1110_U296 | ~new_P2_R1110_U168;
  assign new_P2_R1110_U369 = ~new_P2_R1110_U133 | ~new_P2_R1110_U155 | ~new_P2_R1110_U168;
  assign new_P2_R1110_U370 = ~new_P2_R1110_U297 | ~new_P2_R1110_U301;
  assign new_P2_R1110_U371 = ~new_P2_U3082 | ~new_P2_R1110_U39;
  assign new_P2_R1110_U372 = ~new_P2_U3416 | ~new_P2_R1110_U38;
  assign new_P2_R1110_U373 = ~new_P2_R1110_U372 | ~new_P2_R1110_U371;
  assign new_P2_R1110_U374 = ~new_P2_R1110_U352 | ~new_P2_R1110_U40;
  assign new_P2_R1110_U375 = ~new_P2_R1110_U373 | ~new_P2_R1110_U206;
  assign new_P2_R1110_U376 = ~new_P2_U3083 | ~new_P2_R1110_U36;
  assign new_P2_R1110_U377 = ~new_P2_U3413 | ~new_P2_R1110_U37;
  assign new_P2_R1110_U378 = ~new_P2_R1110_U377 | ~new_P2_R1110_U376;
  assign new_P2_R1110_U379 = ~new_P2_R1110_U353 | ~new_P2_R1110_U144;
  assign new_P2_R1110_U380 = ~new_P2_R1110_U203 | ~new_P2_R1110_U378;
  assign new_P2_R1110_U381 = ~new_P2_U3069 | ~new_P2_R1110_U23;
  assign new_P2_R1110_U382 = ~new_P2_U3410 | ~new_P2_R1110_U21;
  assign new_P2_R1110_U383 = ~new_P2_U3070 | ~new_P2_R1110_U19;
  assign new_P2_R1110_U384 = ~new_P2_U3407 | ~new_P2_R1110_U20;
  assign new_P2_R1110_U385 = ~new_P2_R1110_U384 | ~new_P2_R1110_U383;
  assign new_P2_R1110_U386 = ~new_P2_R1110_U354 | ~new_P2_R1110_U41;
  assign new_P2_R1110_U387 = ~new_P2_R1110_U385 | ~new_P2_R1110_U195;
  assign new_P2_R1110_U388 = ~new_P2_U3066 | ~new_P2_R1110_U35;
  assign new_P2_R1110_U389 = ~new_P2_U3404 | ~new_P2_R1110_U26;
  assign new_P2_R1110_U390 = ~new_P2_U3059 | ~new_P2_R1110_U24;
  assign new_P2_R1110_U391 = ~new_P2_U3401 | ~new_P2_R1110_U25;
  assign new_P2_R1110_U392 = ~new_P2_R1110_U391 | ~new_P2_R1110_U390;
  assign new_P2_R1110_U393 = ~new_P2_R1110_U355 | ~new_P2_R1110_U44;
  assign new_P2_R1110_U394 = ~new_P2_R1110_U392 | ~new_P2_R1110_U221;
  assign new_P2_R1110_U395 = ~new_P2_U3063 | ~new_P2_R1110_U32;
  assign new_P2_R1110_U396 = ~new_P2_U3398 | ~new_P2_R1110_U33;
  assign new_P2_R1110_U397 = ~new_P2_R1110_U396 | ~new_P2_R1110_U395;
  assign new_P2_R1110_U398 = ~new_P2_R1110_U356 | ~new_P2_R1110_U145;
  assign new_P2_R1110_U399 = ~new_P2_R1110_U230 | ~new_P2_R1110_U397;
  assign new_P2_R1110_U400 = ~new_P2_U3067 | ~new_P2_R1110_U27;
  assign new_P2_R1110_U401 = ~new_P2_U3395 | ~new_P2_R1110_U28;
  assign new_P2_R1110_U402 = ~new_P2_U3054 | ~new_P2_R1110_U147;
  assign new_P2_R1110_U403 = ~new_P2_U3904 | ~new_P2_R1110_U146;
  assign new_P2_R1110_U404 = ~new_P2_U3054 | ~new_P2_R1110_U147;
  assign new_P2_R1110_U405 = ~new_P2_U3904 | ~new_P2_R1110_U146;
  assign new_P2_R1110_U406 = ~new_P2_R1110_U405 | ~new_P2_R1110_U404;
  assign new_P2_R1110_U407 = ~new_P2_R1110_U148 | ~new_P2_R1110_U149;
  assign new_P2_R1110_U408 = ~new_P2_R1110_U305 | ~new_P2_R1110_U406;
  assign new_P2_R1110_U409 = ~new_P2_U3053 | ~new_P2_R1110_U88;
  assign new_P2_R1110_U410 = ~new_P2_U3895 | ~new_P2_R1110_U87;
  assign new_P2_R1110_U411 = ~new_P2_U3053 | ~new_P2_R1110_U88;
  assign new_P2_R1110_U412 = ~new_P2_U3895 | ~new_P2_R1110_U87;
  assign new_P2_R1110_U413 = ~new_P2_R1110_U412 | ~new_P2_R1110_U411;
  assign new_P2_R1110_U414 = ~new_P2_R1110_U150 | ~new_P2_R1110_U151;
  assign new_P2_R1110_U415 = ~new_P2_R1110_U303 | ~new_P2_R1110_U413;
  assign new_P2_R1110_U416 = ~new_P2_U3052 | ~new_P2_R1110_U46;
  assign new_P2_R1110_U417 = ~new_P2_U3896 | ~new_P2_R1110_U47;
  assign new_P2_R1110_U418 = ~new_P2_U3052 | ~new_P2_R1110_U46;
  assign new_P2_R1110_U419 = ~new_P2_U3896 | ~new_P2_R1110_U47;
  assign new_P2_R1110_U420 = ~new_P2_R1110_U419 | ~new_P2_R1110_U418;
  assign new_P2_R1110_U421 = ~new_P2_R1110_U152 | ~new_P2_R1110_U153;
  assign new_P2_R1110_U422 = ~new_P2_R1110_U300 | ~new_P2_R1110_U420;
  assign new_P2_R1110_U423 = ~new_P2_U3056 | ~new_P2_R1110_U49;
  assign new_P2_R1110_U424 = ~new_P2_U3897 | ~new_P2_R1110_U48;
  assign new_P2_R1110_U425 = ~new_P2_U3057 | ~new_P2_R1110_U50;
  assign new_P2_R1110_U426 = ~new_P2_U3898 | ~new_P2_R1110_U51;
  assign new_P2_R1110_U427 = ~new_P2_R1110_U426 | ~new_P2_R1110_U425;
  assign new_P2_R1110_U428 = ~new_P2_R1110_U357 | ~new_P2_R1110_U89;
  assign new_P2_R1110_U429 = ~new_P2_R1110_U427 | ~new_P2_R1110_U307;
  assign new_P2_R1110_U430 = ~new_P2_U3064 | ~new_P2_R1110_U52;
  assign new_P2_R1110_U431 = ~new_P2_U3899 | ~new_P2_R1110_U53;
  assign new_P2_R1110_U432 = ~new_P2_R1110_U431 | ~new_P2_R1110_U430;
  assign new_P2_R1110_U433 = ~new_P2_R1110_U358 | ~new_P2_R1110_U155;
  assign new_P2_R1110_U434 = ~new_P2_R1110_U294 | ~new_P2_R1110_U432;
  assign new_P2_R1110_U435 = ~new_P2_U3065 | ~new_P2_R1110_U84;
  assign new_P2_R1110_U436 = ~new_P2_U3900 | ~new_P2_R1110_U85;
  assign new_P2_R1110_U437 = ~new_P2_U3065 | ~new_P2_R1110_U84;
  assign new_P2_R1110_U438 = ~new_P2_U3900 | ~new_P2_R1110_U85;
  assign new_P2_R1110_U439 = ~new_P2_R1110_U438 | ~new_P2_R1110_U437;
  assign new_P2_R1110_U440 = ~new_P2_R1110_U156 | ~new_P2_R1110_U157;
  assign new_P2_R1110_U441 = ~new_P2_R1110_U290 | ~new_P2_R1110_U439;
  assign new_P2_R1110_U442 = ~new_P2_U3060 | ~new_P2_R1110_U82;
  assign new_P2_R1110_U443 = ~new_P2_U3901 | ~new_P2_R1110_U83;
  assign new_P2_R1110_U444 = ~new_P2_U3060 | ~new_P2_R1110_U82;
  assign new_P2_R1110_U445 = ~new_P2_U3901 | ~new_P2_R1110_U83;
  assign new_P2_R1110_U446 = ~new_P2_R1110_U445 | ~new_P2_R1110_U444;
  assign new_P2_R1110_U447 = ~new_P2_R1110_U158 | ~new_P2_R1110_U159;
  assign new_P2_R1110_U448 = ~new_P2_R1110_U286 | ~new_P2_R1110_U446;
  assign new_P2_R1110_U449 = ~new_P2_U3074 | ~new_P2_R1110_U54;
  assign new_P2_R1110_U450 = ~new_P2_U3902 | ~new_P2_R1110_U55;
  assign new_P2_R1110_U451 = ~new_P2_U3074 | ~new_P2_R1110_U54;
  assign new_P2_R1110_U452 = ~new_P2_U3902 | ~new_P2_R1110_U55;
  assign new_P2_R1110_U453 = ~new_P2_R1110_U452 | ~new_P2_R1110_U451;
  assign new_P2_R1110_U454 = ~new_P2_U3075 | ~new_P2_R1110_U81;
  assign new_P2_R1110_U455 = ~new_P2_U3903 | ~new_P2_R1110_U90;
  assign new_P2_R1110_U456 = ~new_P2_R1110_U182 | ~new_P2_R1110_U161;
  assign new_P2_R1110_U457 = ~new_P2_R1110_U328 | ~new_P2_R1110_U31;
  assign new_P2_R1110_U458 = ~new_P2_U3080 | ~new_P2_R1110_U78;
  assign new_P2_R1110_U459 = ~new_P2_U3445 | ~new_P2_R1110_U79;
  assign new_P2_R1110_U460 = ~new_P2_R1110_U459 | ~new_P2_R1110_U458;
  assign new_P2_R1110_U461 = ~new_P2_R1110_U359 | ~new_P2_R1110_U91;
  assign new_P2_R1110_U462 = ~new_P2_R1110_U460 | ~new_P2_R1110_U316;
  assign new_P2_R1110_U463 = ~new_P2_U3081 | ~new_P2_R1110_U75;
  assign new_P2_R1110_U464 = ~new_P2_U3443 | ~new_P2_R1110_U76;
  assign new_P2_R1110_U465 = ~new_P2_R1110_U464 | ~new_P2_R1110_U463;
  assign new_P2_R1110_U466 = ~new_P2_R1110_U360 | ~new_P2_R1110_U162;
  assign new_P2_R1110_U467 = ~new_P2_R1110_U270 | ~new_P2_R1110_U465;
  assign new_P2_R1110_U468 = ~new_P2_U3068 | ~new_P2_R1110_U60;
  assign new_P2_R1110_U469 = ~new_P2_U3440 | ~new_P2_R1110_U58;
  assign new_P2_R1110_U470 = ~new_P2_U3072 | ~new_P2_R1110_U56;
  assign new_P2_R1110_U471 = ~new_P2_U3437 | ~new_P2_R1110_U57;
  assign new_P2_R1110_U472 = ~new_P2_R1110_U471 | ~new_P2_R1110_U470;
  assign new_P2_R1110_U473 = ~new_P2_R1110_U361 | ~new_P2_R1110_U92;
  assign new_P2_R1110_U474 = ~new_P2_R1110_U472 | ~new_P2_R1110_U262;
  assign new_P2_R1110_U475 = ~new_P2_U3073 | ~new_P2_R1110_U73;
  assign new_P2_R1110_U476 = ~new_P2_U3434 | ~new_P2_R1110_U74;
  assign new_P2_R1110_U477 = ~new_P2_U3073 | ~new_P2_R1110_U73;
  assign new_P2_R1110_U478 = ~new_P2_U3434 | ~new_P2_R1110_U74;
  assign new_P2_R1110_U479 = ~new_P2_R1110_U478 | ~new_P2_R1110_U477;
  assign new_P2_R1110_U480 = ~new_P2_R1110_U163 | ~new_P2_R1110_U164;
  assign new_P2_R1110_U481 = ~new_P2_R1110_U258 | ~new_P2_R1110_U479;
  assign new_P2_R1110_U482 = ~new_P2_U3078 | ~new_P2_R1110_U71;
  assign new_P2_R1110_U483 = ~new_P2_U3431 | ~new_P2_R1110_U72;
  assign new_P2_R1110_U484 = ~new_P2_U3078 | ~new_P2_R1110_U71;
  assign new_P2_R1110_U485 = ~new_P2_U3431 | ~new_P2_R1110_U72;
  assign new_P2_R1110_U486 = ~new_P2_R1110_U485 | ~new_P2_R1110_U484;
  assign new_P2_R1110_U487 = ~new_P2_R1110_U165 | ~new_P2_R1110_U166;
  assign new_P2_R1110_U488 = ~new_P2_R1110_U254 | ~new_P2_R1110_U486;
  assign new_P2_R1110_U489 = ~new_P2_U3079 | ~new_P2_R1110_U61;
  assign new_P2_R1110_U490 = ~new_P2_U3428 | ~new_P2_R1110_U62;
  assign new_P2_R1110_U491 = ~new_P2_U3071 | ~new_P2_R1110_U69;
  assign new_P2_R1110_U492 = ~new_P2_U3425 | ~new_P2_R1110_U70;
  assign new_P2_R1110_U493 = ~new_P2_R1110_U492 | ~new_P2_R1110_U491;
  assign new_P2_R1110_U494 = ~new_P2_R1110_U362 | ~new_P2_R1110_U93;
  assign new_P2_R1110_U495 = ~new_P2_R1110_U493 | ~new_P2_R1110_U338;
  assign new_P2_R1110_U496 = ~new_P2_U3062 | ~new_P2_R1110_U66;
  assign new_P2_R1110_U497 = ~new_P2_U3422 | ~new_P2_R1110_U67;
  assign new_P2_R1110_U498 = ~new_P2_R1110_U497 | ~new_P2_R1110_U496;
  assign new_P2_R1110_U499 = ~new_P2_R1110_U363 | ~new_P2_R1110_U167;
  assign new_P2_R1110_U500 = ~new_P2_R1110_U244 | ~new_P2_R1110_U498;
  assign new_P2_R1110_U501 = ~new_P2_U3061 | ~new_P2_R1110_U63;
  assign new_P2_R1110_U502 = ~new_P2_U3419 | ~new_P2_R1110_U64;
  assign new_P2_R1110_U503 = ~new_P2_U3076 | ~new_P2_R1110_U29;
  assign new_P2_R1110_U504 = ~new_P2_U3387 | ~new_P2_R1110_U30;
  assign new_P2_R1297_U6 = new_P2_U3058 & new_P2_R1297_U7;
  assign new_P2_R1297_U7 = ~new_P2_U3055;
  assign new_P2_R1077_U4 = new_P2_R1077_U179 & new_P2_R1077_U178;
  assign new_P2_R1077_U5 = new_P2_R1077_U197 & new_P2_R1077_U196;
  assign new_P2_R1077_U6 = new_P2_R1077_U237 & new_P2_R1077_U236;
  assign new_P2_R1077_U7 = new_P2_R1077_U246 & new_P2_R1077_U245;
  assign new_P2_R1077_U8 = new_P2_R1077_U264 & new_P2_R1077_U263;
  assign new_P2_R1077_U9 = new_P2_R1077_U272 & new_P2_R1077_U271;
  assign new_P2_R1077_U10 = new_P2_R1077_U351 & new_P2_R1077_U348;
  assign new_P2_R1077_U11 = new_P2_R1077_U344 & new_P2_R1077_U341;
  assign new_P2_R1077_U12 = new_P2_R1077_U335 & new_P2_R1077_U332;
  assign new_P2_R1077_U13 = new_P2_R1077_U326 & new_P2_R1077_U323;
  assign new_P2_R1077_U14 = new_P2_R1077_U320 & new_P2_R1077_U318;
  assign new_P2_R1077_U15 = new_P2_R1077_U313 & new_P2_R1077_U310;
  assign new_P2_R1077_U16 = new_P2_R1077_U235 & new_P2_R1077_U232;
  assign new_P2_R1077_U17 = new_P2_R1077_U227 & new_P2_R1077_U224;
  assign new_P2_R1077_U18 = new_P2_R1077_U213 & new_P2_R1077_U210;
  assign new_P2_R1077_U19 = ~new_P2_U3407;
  assign new_P2_R1077_U20 = ~new_P2_U3070;
  assign new_P2_R1077_U21 = ~new_P2_U3069;
  assign new_P2_R1077_U22 = ~new_P2_U3070 | ~new_P2_U3407;
  assign new_P2_R1077_U23 = ~new_P2_U3410;
  assign new_P2_R1077_U24 = ~new_P2_U3401;
  assign new_P2_R1077_U25 = ~new_P2_U3059;
  assign new_P2_R1077_U26 = ~new_P2_U3066;
  assign new_P2_R1077_U27 = ~new_P2_U3395;
  assign new_P2_R1077_U28 = ~new_P2_U3067;
  assign new_P2_R1077_U29 = ~new_P2_U3387;
  assign new_P2_R1077_U30 = ~new_P2_U3076;
  assign new_P2_R1077_U31 = ~new_P2_U3076 | ~new_P2_U3387;
  assign new_P2_R1077_U32 = ~new_P2_U3398;
  assign new_P2_R1077_U33 = ~new_P2_U3063;
  assign new_P2_R1077_U34 = ~new_P2_U3059 | ~new_P2_U3401;
  assign new_P2_R1077_U35 = ~new_P2_U3404;
  assign new_P2_R1077_U36 = ~new_P2_U3413;
  assign new_P2_R1077_U37 = ~new_P2_U3083;
  assign new_P2_R1077_U38 = ~new_P2_U3082;
  assign new_P2_R1077_U39 = ~new_P2_U3416;
  assign new_P2_R1077_U40 = ~new_P2_R1077_U65 | ~new_P2_R1077_U205;
  assign new_P2_R1077_U41 = ~new_P2_R1077_U117 | ~new_P2_R1077_U193;
  assign new_P2_R1077_U42 = ~new_P2_R1077_U182 | ~new_P2_R1077_U183;
  assign new_P2_R1077_U43 = ~new_P2_U3392 | ~new_P2_U3077;
  assign new_P2_R1077_U44 = ~new_P2_R1077_U122 | ~new_P2_R1077_U219;
  assign new_P2_R1077_U45 = ~new_P2_R1077_U216 | ~new_P2_R1077_U215;
  assign new_P2_R1077_U46 = ~new_P2_U3896;
  assign new_P2_R1077_U47 = ~new_P2_U3052;
  assign new_P2_R1077_U48 = ~new_P2_U3056;
  assign new_P2_R1077_U49 = ~new_P2_U3897;
  assign new_P2_R1077_U50 = ~new_P2_U3898;
  assign new_P2_R1077_U51 = ~new_P2_U3057;
  assign new_P2_R1077_U52 = ~new_P2_U3899;
  assign new_P2_R1077_U53 = ~new_P2_U3064;
  assign new_P2_R1077_U54 = ~new_P2_U3902;
  assign new_P2_R1077_U55 = ~new_P2_U3074;
  assign new_P2_R1077_U56 = ~new_P2_U3437;
  assign new_P2_R1077_U57 = ~new_P2_U3072;
  assign new_P2_R1077_U58 = ~new_P2_U3068;
  assign new_P2_R1077_U59 = ~new_P2_U3072 | ~new_P2_U3437;
  assign new_P2_R1077_U60 = ~new_P2_U3440;
  assign new_P2_R1077_U61 = ~new_P2_U3428;
  assign new_P2_R1077_U62 = ~new_P2_U3079;
  assign new_P2_R1077_U63 = ~new_P2_U3419;
  assign new_P2_R1077_U64 = ~new_P2_U3061;
  assign new_P2_R1077_U65 = ~new_P2_U3083 | ~new_P2_U3413;
  assign new_P2_R1077_U66 = ~new_P2_U3422;
  assign new_P2_R1077_U67 = ~new_P2_U3062;
  assign new_P2_R1077_U68 = ~new_P2_U3062 | ~new_P2_U3422;
  assign new_P2_R1077_U69 = ~new_P2_U3425;
  assign new_P2_R1077_U70 = ~new_P2_U3071;
  assign new_P2_R1077_U71 = ~new_P2_U3431;
  assign new_P2_R1077_U72 = ~new_P2_U3078;
  assign new_P2_R1077_U73 = ~new_P2_U3434;
  assign new_P2_R1077_U74 = ~new_P2_U3073;
  assign new_P2_R1077_U75 = ~new_P2_U3443;
  assign new_P2_R1077_U76 = ~new_P2_U3081;
  assign new_P2_R1077_U77 = ~new_P2_U3081 | ~new_P2_U3443;
  assign new_P2_R1077_U78 = ~new_P2_U3445;
  assign new_P2_R1077_U79 = ~new_P2_U3080;
  assign new_P2_R1077_U80 = ~new_P2_U3080 | ~new_P2_U3445;
  assign new_P2_R1077_U81 = ~new_P2_U3903;
  assign new_P2_R1077_U82 = ~new_P2_U3901;
  assign new_P2_R1077_U83 = ~new_P2_U3060;
  assign new_P2_R1077_U84 = ~new_P2_U3900;
  assign new_P2_R1077_U85 = ~new_P2_U3065;
  assign new_P2_R1077_U86 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1077_U87 = ~new_P2_U3053;
  assign new_P2_R1077_U88 = ~new_P2_U3895;
  assign new_P2_R1077_U89 = ~new_P2_R1077_U306 | ~new_P2_R1077_U176;
  assign new_P2_R1077_U90 = ~new_P2_U3075;
  assign new_P2_R1077_U91 = ~new_P2_R1077_U77 | ~new_P2_R1077_U315;
  assign new_P2_R1077_U92 = ~new_P2_R1077_U261 | ~new_P2_R1077_U260;
  assign new_P2_R1077_U93 = ~new_P2_R1077_U68 | ~new_P2_R1077_U337;
  assign new_P2_R1077_U94 = ~new_P2_R1077_U457 | ~new_P2_R1077_U456;
  assign new_P2_R1077_U95 = ~new_P2_R1077_U504 | ~new_P2_R1077_U503;
  assign new_P2_R1077_U96 = ~new_P2_R1077_U375 | ~new_P2_R1077_U374;
  assign new_P2_R1077_U97 = ~new_P2_R1077_U380 | ~new_P2_R1077_U379;
  assign new_P2_R1077_U98 = ~new_P2_R1077_U387 | ~new_P2_R1077_U386;
  assign new_P2_R1077_U99 = ~new_P2_R1077_U394 | ~new_P2_R1077_U393;
  assign new_P2_R1077_U100 = ~new_P2_R1077_U399 | ~new_P2_R1077_U398;
  assign new_P2_R1077_U101 = ~new_P2_R1077_U408 | ~new_P2_R1077_U407;
  assign new_P2_R1077_U102 = ~new_P2_R1077_U415 | ~new_P2_R1077_U414;
  assign new_P2_R1077_U103 = ~new_P2_R1077_U422 | ~new_P2_R1077_U421;
  assign new_P2_R1077_U104 = ~new_P2_R1077_U429 | ~new_P2_R1077_U428;
  assign new_P2_R1077_U105 = ~new_P2_R1077_U434 | ~new_P2_R1077_U433;
  assign new_P2_R1077_U106 = ~new_P2_R1077_U441 | ~new_P2_R1077_U440;
  assign new_P2_R1077_U107 = ~new_P2_R1077_U448 | ~new_P2_R1077_U447;
  assign new_P2_R1077_U108 = ~new_P2_R1077_U462 | ~new_P2_R1077_U461;
  assign new_P2_R1077_U109 = ~new_P2_R1077_U467 | ~new_P2_R1077_U466;
  assign new_P2_R1077_U110 = ~new_P2_R1077_U474 | ~new_P2_R1077_U473;
  assign new_P2_R1077_U111 = ~new_P2_R1077_U481 | ~new_P2_R1077_U480;
  assign new_P2_R1077_U112 = ~new_P2_R1077_U488 | ~new_P2_R1077_U487;
  assign new_P2_R1077_U113 = ~new_P2_R1077_U495 | ~new_P2_R1077_U494;
  assign new_P2_R1077_U114 = ~new_P2_R1077_U500 | ~new_P2_R1077_U499;
  assign new_P2_R1077_U115 = new_P2_R1077_U189 & new_P2_R1077_U187;
  assign new_P2_R1077_U116 = new_P2_R1077_U4 & new_P2_R1077_U180;
  assign new_P2_R1077_U117 = new_P2_R1077_U194 & new_P2_R1077_U192;
  assign new_P2_R1077_U118 = new_P2_R1077_U201 & new_P2_R1077_U200;
  assign new_P2_R1077_U119 = new_P2_R1077_U22 & new_P2_R1077_U382 & new_P2_R1077_U381;
  assign new_P2_R1077_U120 = new_P2_R1077_U212 & new_P2_R1077_U5;
  assign new_P2_R1077_U121 = new_P2_R1077_U181 & new_P2_R1077_U180;
  assign new_P2_R1077_U122 = new_P2_R1077_U220 & new_P2_R1077_U218;
  assign new_P2_R1077_U123 = new_P2_R1077_U34 & new_P2_R1077_U389 & new_P2_R1077_U388;
  assign new_P2_R1077_U124 = new_P2_R1077_U226 & new_P2_R1077_U4;
  assign new_P2_R1077_U125 = new_P2_R1077_U234 & new_P2_R1077_U181;
  assign new_P2_R1077_U126 = new_P2_R1077_U204 & new_P2_R1077_U6;
  assign new_P2_R1077_U127 = new_P2_R1077_U243 & new_P2_R1077_U239;
  assign new_P2_R1077_U128 = new_P2_R1077_U250 & new_P2_R1077_U7;
  assign new_P2_R1077_U129 = new_P2_R1077_U253 & new_P2_R1077_U248;
  assign new_P2_R1077_U130 = new_P2_R1077_U268 & new_P2_R1077_U267;
  assign new_P2_R1077_U131 = new_P2_R1077_U9 & new_P2_R1077_U282;
  assign new_P2_R1077_U132 = new_P2_R1077_U285 & new_P2_R1077_U280;
  assign new_P2_R1077_U133 = new_P2_R1077_U301 & new_P2_R1077_U298;
  assign new_P2_R1077_U134 = new_P2_R1077_U368 & new_P2_R1077_U302;
  assign new_P2_R1077_U135 = new_P2_R1077_U160 & new_P2_R1077_U278;
  assign new_P2_R1077_U136 = new_P2_R1077_U80 & new_P2_R1077_U455 & new_P2_R1077_U454;
  assign new_P2_R1077_U137 = new_P2_R1077_U325 & new_P2_R1077_U9;
  assign new_P2_R1077_U138 = new_P2_R1077_U59 & new_P2_R1077_U469 & new_P2_R1077_U468;
  assign new_P2_R1077_U139 = new_P2_R1077_U334 & new_P2_R1077_U8;
  assign new_P2_R1077_U140 = new_P2_R1077_U172 & new_P2_R1077_U490 & new_P2_R1077_U489;
  assign new_P2_R1077_U141 = new_P2_R1077_U343 & new_P2_R1077_U7;
  assign new_P2_R1077_U142 = new_P2_R1077_U171 & new_P2_R1077_U502 & new_P2_R1077_U501;
  assign new_P2_R1077_U143 = new_P2_R1077_U350 & new_P2_R1077_U6;
  assign new_P2_R1077_U144 = ~new_P2_R1077_U118 | ~new_P2_R1077_U202;
  assign new_P2_R1077_U145 = ~new_P2_R1077_U217 | ~new_P2_R1077_U229;
  assign new_P2_R1077_U146 = ~new_P2_U3054;
  assign new_P2_R1077_U147 = ~new_P2_U3904;
  assign new_P2_R1077_U148 = new_P2_R1077_U403 & new_P2_R1077_U402;
  assign new_P2_R1077_U149 = ~new_P2_R1077_U364 | ~new_P2_R1077_U304 | ~new_P2_R1077_U169;
  assign new_P2_R1077_U150 = new_P2_R1077_U410 & new_P2_R1077_U409;
  assign new_P2_R1077_U151 = ~new_P2_R1077_U134 | ~new_P2_R1077_U370 | ~new_P2_R1077_U369;
  assign new_P2_R1077_U152 = new_P2_R1077_U417 & new_P2_R1077_U416;
  assign new_P2_R1077_U153 = ~new_P2_R1077_U86 | ~new_P2_R1077_U365 | ~new_P2_R1077_U299;
  assign new_P2_R1077_U154 = new_P2_R1077_U424 & new_P2_R1077_U423;
  assign new_P2_R1077_U155 = ~new_P2_R1077_U293 | ~new_P2_R1077_U292;
  assign new_P2_R1077_U156 = new_P2_R1077_U436 & new_P2_R1077_U435;
  assign new_P2_R1077_U157 = ~new_P2_R1077_U289 | ~new_P2_R1077_U288;
  assign new_P2_R1077_U158 = new_P2_R1077_U443 & new_P2_R1077_U442;
  assign new_P2_R1077_U159 = ~new_P2_R1077_U132 | ~new_P2_R1077_U284;
  assign new_P2_R1077_U160 = new_P2_R1077_U450 & new_P2_R1077_U449;
  assign new_P2_R1077_U161 = ~new_P2_R1077_U43 | ~new_P2_R1077_U327;
  assign new_P2_R1077_U162 = ~new_P2_R1077_U130 | ~new_P2_R1077_U269;
  assign new_P2_R1077_U163 = new_P2_R1077_U476 & new_P2_R1077_U475;
  assign new_P2_R1077_U164 = ~new_P2_R1077_U257 | ~new_P2_R1077_U256;
  assign new_P2_R1077_U165 = new_P2_R1077_U483 & new_P2_R1077_U482;
  assign new_P2_R1077_U166 = ~new_P2_R1077_U129 | ~new_P2_R1077_U252;
  assign new_P2_R1077_U167 = ~new_P2_R1077_U127 | ~new_P2_R1077_U242;
  assign new_P2_R1077_U168 = ~new_P2_R1077_U367 | ~new_P2_R1077_U366;
  assign new_P2_R1077_U169 = ~new_P2_U3053 | ~new_P2_R1077_U151;
  assign new_P2_R1077_U170 = ~new_P2_R1077_U34;
  assign new_P2_R1077_U171 = ~new_P2_U3416 | ~new_P2_U3082;
  assign new_P2_R1077_U172 = ~new_P2_U3071 | ~new_P2_U3425;
  assign new_P2_R1077_U173 = ~new_P2_U3057 | ~new_P2_U3898;
  assign new_P2_R1077_U174 = ~new_P2_R1077_U68;
  assign new_P2_R1077_U175 = ~new_P2_R1077_U77;
  assign new_P2_R1077_U176 = ~new_P2_U3064 | ~new_P2_U3899;
  assign new_P2_R1077_U177 = ~new_P2_R1077_U65;
  assign new_P2_R1077_U178 = new_P2_U3066 | new_P2_U3404;
  assign new_P2_R1077_U179 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1077_U180 = new_P2_U3398 | new_P2_U3063;
  assign new_P2_R1077_U181 = new_P2_U3395 | new_P2_U3067;
  assign new_P2_R1077_U182 = ~new_P2_R1077_U31;
  assign new_P2_R1077_U183 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1077_U184 = ~new_P2_R1077_U42;
  assign new_P2_R1077_U185 = ~new_P2_R1077_U43;
  assign new_P2_R1077_U186 = ~new_P2_R1077_U42 | ~new_P2_R1077_U43;
  assign new_P2_R1077_U187 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1077_U188 = ~new_P2_R1077_U186 | ~new_P2_R1077_U181;
  assign new_P2_R1077_U189 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1077_U190 = ~new_P2_R1077_U115 | ~new_P2_R1077_U188;
  assign new_P2_R1077_U191 = ~new_P2_R1077_U35 | ~new_P2_R1077_U34;
  assign new_P2_R1077_U192 = ~new_P2_U3066 | ~new_P2_R1077_U191;
  assign new_P2_R1077_U193 = ~new_P2_R1077_U116 | ~new_P2_R1077_U190;
  assign new_P2_R1077_U194 = ~new_P2_U3404 | ~new_P2_R1077_U170;
  assign new_P2_R1077_U195 = ~new_P2_R1077_U41;
  assign new_P2_R1077_U196 = new_P2_U3069 | new_P2_U3410;
  assign new_P2_R1077_U197 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1077_U198 = ~new_P2_R1077_U22;
  assign new_P2_R1077_U199 = ~new_P2_R1077_U23 | ~new_P2_R1077_U22;
  assign new_P2_R1077_U200 = ~new_P2_U3069 | ~new_P2_R1077_U199;
  assign new_P2_R1077_U201 = ~new_P2_U3410 | ~new_P2_R1077_U198;
  assign new_P2_R1077_U202 = ~new_P2_R1077_U5 | ~new_P2_R1077_U41;
  assign new_P2_R1077_U203 = ~new_P2_R1077_U144;
  assign new_P2_R1077_U204 = new_P2_U3413 | new_P2_U3083;
  assign new_P2_R1077_U205 = ~new_P2_R1077_U204 | ~new_P2_R1077_U144;
  assign new_P2_R1077_U206 = ~new_P2_R1077_U40;
  assign new_P2_R1077_U207 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1077_U208 = new_P2_U3407 | new_P2_U3070;
  assign new_P2_R1077_U209 = ~new_P2_R1077_U208 | ~new_P2_R1077_U41;
  assign new_P2_R1077_U210 = ~new_P2_R1077_U119 | ~new_P2_R1077_U209;
  assign new_P2_R1077_U211 = ~new_P2_R1077_U195 | ~new_P2_R1077_U22;
  assign new_P2_R1077_U212 = ~new_P2_U3410 | ~new_P2_U3069;
  assign new_P2_R1077_U213 = ~new_P2_R1077_U120 | ~new_P2_R1077_U211;
  assign new_P2_R1077_U214 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1077_U215 = ~new_P2_R1077_U185 | ~new_P2_R1077_U181;
  assign new_P2_R1077_U216 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1077_U217 = ~new_P2_R1077_U45;
  assign new_P2_R1077_U218 = ~new_P2_R1077_U121 | ~new_P2_R1077_U184;
  assign new_P2_R1077_U219 = ~new_P2_R1077_U45 | ~new_P2_R1077_U180;
  assign new_P2_R1077_U220 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1077_U221 = ~new_P2_R1077_U44;
  assign new_P2_R1077_U222 = new_P2_U3401 | new_P2_U3059;
  assign new_P2_R1077_U223 = ~new_P2_R1077_U222 | ~new_P2_R1077_U44;
  assign new_P2_R1077_U224 = ~new_P2_R1077_U123 | ~new_P2_R1077_U223;
  assign new_P2_R1077_U225 = ~new_P2_R1077_U221 | ~new_P2_R1077_U34;
  assign new_P2_R1077_U226 = ~new_P2_U3404 | ~new_P2_U3066;
  assign new_P2_R1077_U227 = ~new_P2_R1077_U124 | ~new_P2_R1077_U225;
  assign new_P2_R1077_U228 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1077_U229 = ~new_P2_R1077_U184 | ~new_P2_R1077_U181;
  assign new_P2_R1077_U230 = ~new_P2_R1077_U145;
  assign new_P2_R1077_U231 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1077_U232 = ~new_P2_R1077_U42 | ~new_P2_R1077_U43 | ~new_P2_R1077_U401 | ~new_P2_R1077_U400;
  assign new_P2_R1077_U233 = ~new_P2_R1077_U43 | ~new_P2_R1077_U42;
  assign new_P2_R1077_U234 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1077_U235 = ~new_P2_R1077_U125 | ~new_P2_R1077_U233;
  assign new_P2_R1077_U236 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1077_U237 = new_P2_U3061 | new_P2_U3419;
  assign new_P2_R1077_U238 = ~new_P2_R1077_U177 | ~new_P2_R1077_U6;
  assign new_P2_R1077_U239 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1077_U240 = ~new_P2_R1077_U171 | ~new_P2_R1077_U238;
  assign new_P2_R1077_U241 = new_P2_U3419 | new_P2_U3061;
  assign new_P2_R1077_U242 = ~new_P2_R1077_U126 | ~new_P2_R1077_U144;
  assign new_P2_R1077_U243 = ~new_P2_R1077_U241 | ~new_P2_R1077_U240;
  assign new_P2_R1077_U244 = ~new_P2_R1077_U167;
  assign new_P2_R1077_U245 = new_P2_U3079 | new_P2_U3428;
  assign new_P2_R1077_U246 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1077_U247 = ~new_P2_R1077_U174 | ~new_P2_R1077_U7;
  assign new_P2_R1077_U248 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1077_U249 = ~new_P2_R1077_U172 | ~new_P2_R1077_U247;
  assign new_P2_R1077_U250 = new_P2_U3422 | new_P2_U3062;
  assign new_P2_R1077_U251 = new_P2_U3428 | new_P2_U3079;
  assign new_P2_R1077_U252 = ~new_P2_R1077_U128 | ~new_P2_R1077_U167;
  assign new_P2_R1077_U253 = ~new_P2_R1077_U251 | ~new_P2_R1077_U249;
  assign new_P2_R1077_U254 = ~new_P2_R1077_U166;
  assign new_P2_R1077_U255 = new_P2_U3431 | new_P2_U3078;
  assign new_P2_R1077_U256 = ~new_P2_R1077_U255 | ~new_P2_R1077_U166;
  assign new_P2_R1077_U257 = ~new_P2_U3078 | ~new_P2_U3431;
  assign new_P2_R1077_U258 = ~new_P2_R1077_U164;
  assign new_P2_R1077_U259 = new_P2_U3434 | new_P2_U3073;
  assign new_P2_R1077_U260 = ~new_P2_R1077_U259 | ~new_P2_R1077_U164;
  assign new_P2_R1077_U261 = ~new_P2_U3073 | ~new_P2_U3434;
  assign new_P2_R1077_U262 = ~new_P2_R1077_U92;
  assign new_P2_R1077_U263 = new_P2_U3068 | new_P2_U3440;
  assign new_P2_R1077_U264 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1077_U265 = ~new_P2_R1077_U59;
  assign new_P2_R1077_U266 = ~new_P2_R1077_U60 | ~new_P2_R1077_U59;
  assign new_P2_R1077_U267 = ~new_P2_U3068 | ~new_P2_R1077_U266;
  assign new_P2_R1077_U268 = ~new_P2_U3440 | ~new_P2_R1077_U265;
  assign new_P2_R1077_U269 = ~new_P2_R1077_U8 | ~new_P2_R1077_U92;
  assign new_P2_R1077_U270 = ~new_P2_R1077_U162;
  assign new_P2_R1077_U271 = new_P2_U3075 | new_P2_U3903;
  assign new_P2_R1077_U272 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1077_U273 = new_P2_U3074 | new_P2_U3902;
  assign new_P2_R1077_U274 = ~new_P2_R1077_U80;
  assign new_P2_R1077_U275 = ~new_P2_U3903 | ~new_P2_R1077_U274;
  assign new_P2_R1077_U276 = ~new_P2_R1077_U275 | ~new_P2_R1077_U90;
  assign new_P2_R1077_U277 = ~new_P2_R1077_U80 | ~new_P2_R1077_U81;
  assign new_P2_R1077_U278 = ~new_P2_R1077_U277 | ~new_P2_R1077_U276;
  assign new_P2_R1077_U279 = ~new_P2_R1077_U175 | ~new_P2_R1077_U9;
  assign new_P2_R1077_U280 = ~new_P2_U3074 | ~new_P2_U3902;
  assign new_P2_R1077_U281 = ~new_P2_R1077_U278 | ~new_P2_R1077_U279;
  assign new_P2_R1077_U282 = new_P2_U3443 | new_P2_U3081;
  assign new_P2_R1077_U283 = new_P2_U3902 | new_P2_U3074;
  assign new_P2_R1077_U284 = ~new_P2_R1077_U131 | ~new_P2_R1077_U273 | ~new_P2_R1077_U162;
  assign new_P2_R1077_U285 = ~new_P2_R1077_U283 | ~new_P2_R1077_U281;
  assign new_P2_R1077_U286 = ~new_P2_R1077_U159;
  assign new_P2_R1077_U287 = new_P2_U3901 | new_P2_U3060;
  assign new_P2_R1077_U288 = ~new_P2_R1077_U287 | ~new_P2_R1077_U159;
  assign new_P2_R1077_U289 = ~new_P2_U3060 | ~new_P2_U3901;
  assign new_P2_R1077_U290 = ~new_P2_R1077_U157;
  assign new_P2_R1077_U291 = new_P2_U3900 | new_P2_U3065;
  assign new_P2_R1077_U292 = ~new_P2_R1077_U291 | ~new_P2_R1077_U157;
  assign new_P2_R1077_U293 = ~new_P2_U3065 | ~new_P2_U3900;
  assign new_P2_R1077_U294 = ~new_P2_R1077_U155;
  assign new_P2_R1077_U295 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1077_U296 = ~new_P2_R1077_U176 | ~new_P2_R1077_U173;
  assign new_P2_R1077_U297 = ~new_P2_R1077_U86;
  assign new_P2_R1077_U298 = new_P2_U3899 | new_P2_U3064;
  assign new_P2_R1077_U299 = ~new_P2_R1077_U168 | ~new_P2_R1077_U155 | ~new_P2_R1077_U298;
  assign new_P2_R1077_U300 = ~new_P2_R1077_U153;
  assign new_P2_R1077_U301 = new_P2_U3896 | new_P2_U3052;
  assign new_P2_R1077_U302 = ~new_P2_U3052 | ~new_P2_U3896;
  assign new_P2_R1077_U303 = ~new_P2_R1077_U151;
  assign new_P2_R1077_U304 = ~new_P2_U3895 | ~new_P2_R1077_U151;
  assign new_P2_R1077_U305 = ~new_P2_R1077_U149;
  assign new_P2_R1077_U306 = ~new_P2_R1077_U298 | ~new_P2_R1077_U155;
  assign new_P2_R1077_U307 = ~new_P2_R1077_U89;
  assign new_P2_R1077_U308 = new_P2_U3898 | new_P2_U3057;
  assign new_P2_R1077_U309 = ~new_P2_R1077_U308 | ~new_P2_R1077_U89;
  assign new_P2_R1077_U310 = ~new_P2_R1077_U154 | ~new_P2_R1077_U309 | ~new_P2_R1077_U173;
  assign new_P2_R1077_U311 = ~new_P2_R1077_U307 | ~new_P2_R1077_U173;
  assign new_P2_R1077_U312 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1077_U313 = ~new_P2_R1077_U168 | ~new_P2_R1077_U311 | ~new_P2_R1077_U312;
  assign new_P2_R1077_U314 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1077_U315 = ~new_P2_R1077_U282 | ~new_P2_R1077_U162;
  assign new_P2_R1077_U316 = ~new_P2_R1077_U91;
  assign new_P2_R1077_U317 = ~new_P2_R1077_U9 | ~new_P2_R1077_U91;
  assign new_P2_R1077_U318 = ~new_P2_R1077_U135 | ~new_P2_R1077_U317;
  assign new_P2_R1077_U319 = ~new_P2_R1077_U317 | ~new_P2_R1077_U278;
  assign new_P2_R1077_U320 = ~new_P2_R1077_U453 | ~new_P2_R1077_U319;
  assign new_P2_R1077_U321 = new_P2_U3445 | new_P2_U3080;
  assign new_P2_R1077_U322 = ~new_P2_R1077_U321 | ~new_P2_R1077_U91;
  assign new_P2_R1077_U323 = ~new_P2_R1077_U136 | ~new_P2_R1077_U322;
  assign new_P2_R1077_U324 = ~new_P2_R1077_U316 | ~new_P2_R1077_U80;
  assign new_P2_R1077_U325 = ~new_P2_U3075 | ~new_P2_U3903;
  assign new_P2_R1077_U326 = ~new_P2_R1077_U137 | ~new_P2_R1077_U324;
  assign new_P2_R1077_U327 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1077_U328 = ~new_P2_R1077_U161;
  assign new_P2_R1077_U329 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1077_U330 = new_P2_U3437 | new_P2_U3072;
  assign new_P2_R1077_U331 = ~new_P2_R1077_U330 | ~new_P2_R1077_U92;
  assign new_P2_R1077_U332 = ~new_P2_R1077_U138 | ~new_P2_R1077_U331;
  assign new_P2_R1077_U333 = ~new_P2_R1077_U262 | ~new_P2_R1077_U59;
  assign new_P2_R1077_U334 = ~new_P2_U3440 | ~new_P2_U3068;
  assign new_P2_R1077_U335 = ~new_P2_R1077_U139 | ~new_P2_R1077_U333;
  assign new_P2_R1077_U336 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1077_U337 = ~new_P2_R1077_U250 | ~new_P2_R1077_U167;
  assign new_P2_R1077_U338 = ~new_P2_R1077_U93;
  assign new_P2_R1077_U339 = new_P2_U3425 | new_P2_U3071;
  assign new_P2_R1077_U340 = ~new_P2_R1077_U339 | ~new_P2_R1077_U93;
  assign new_P2_R1077_U341 = ~new_P2_R1077_U140 | ~new_P2_R1077_U340;
  assign new_P2_R1077_U342 = ~new_P2_R1077_U338 | ~new_P2_R1077_U172;
  assign new_P2_R1077_U343 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1077_U344 = ~new_P2_R1077_U141 | ~new_P2_R1077_U342;
  assign new_P2_R1077_U345 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1077_U346 = new_P2_U3416 | new_P2_U3082;
  assign new_P2_R1077_U347 = ~new_P2_R1077_U346 | ~new_P2_R1077_U40;
  assign new_P2_R1077_U348 = ~new_P2_R1077_U142 | ~new_P2_R1077_U347;
  assign new_P2_R1077_U349 = ~new_P2_R1077_U206 | ~new_P2_R1077_U171;
  assign new_P2_R1077_U350 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1077_U351 = ~new_P2_R1077_U143 | ~new_P2_R1077_U349;
  assign new_P2_R1077_U352 = ~new_P2_R1077_U207 | ~new_P2_R1077_U171;
  assign new_P2_R1077_U353 = ~new_P2_R1077_U204 | ~new_P2_R1077_U65;
  assign new_P2_R1077_U354 = ~new_P2_R1077_U214 | ~new_P2_R1077_U22;
  assign new_P2_R1077_U355 = ~new_P2_R1077_U228 | ~new_P2_R1077_U34;
  assign new_P2_R1077_U356 = ~new_P2_R1077_U231 | ~new_P2_R1077_U180;
  assign new_P2_R1077_U357 = ~new_P2_R1077_U314 | ~new_P2_R1077_U173;
  assign new_P2_R1077_U358 = ~new_P2_R1077_U298 | ~new_P2_R1077_U176;
  assign new_P2_R1077_U359 = ~new_P2_R1077_U329 | ~new_P2_R1077_U80;
  assign new_P2_R1077_U360 = ~new_P2_R1077_U282 | ~new_P2_R1077_U77;
  assign new_P2_R1077_U361 = ~new_P2_R1077_U336 | ~new_P2_R1077_U59;
  assign new_P2_R1077_U362 = ~new_P2_R1077_U345 | ~new_P2_R1077_U172;
  assign new_P2_R1077_U363 = ~new_P2_R1077_U250 | ~new_P2_R1077_U68;
  assign new_P2_R1077_U364 = ~new_P2_U3895 | ~new_P2_U3053;
  assign new_P2_R1077_U365 = ~new_P2_R1077_U296 | ~new_P2_R1077_U168;
  assign new_P2_R1077_U366 = ~new_P2_U3056 | ~new_P2_R1077_U295;
  assign new_P2_R1077_U367 = ~new_P2_U3897 | ~new_P2_R1077_U295;
  assign new_P2_R1077_U368 = ~new_P2_R1077_U301 | ~new_P2_R1077_U296 | ~new_P2_R1077_U168;
  assign new_P2_R1077_U369 = ~new_P2_R1077_U133 | ~new_P2_R1077_U155 | ~new_P2_R1077_U168;
  assign new_P2_R1077_U370 = ~new_P2_R1077_U297 | ~new_P2_R1077_U301;
  assign new_P2_R1077_U371 = ~new_P2_U3082 | ~new_P2_R1077_U39;
  assign new_P2_R1077_U372 = ~new_P2_U3416 | ~new_P2_R1077_U38;
  assign new_P2_R1077_U373 = ~new_P2_R1077_U372 | ~new_P2_R1077_U371;
  assign new_P2_R1077_U374 = ~new_P2_R1077_U352 | ~new_P2_R1077_U40;
  assign new_P2_R1077_U375 = ~new_P2_R1077_U373 | ~new_P2_R1077_U206;
  assign new_P2_R1077_U376 = ~new_P2_U3083 | ~new_P2_R1077_U36;
  assign new_P2_R1077_U377 = ~new_P2_U3413 | ~new_P2_R1077_U37;
  assign new_P2_R1077_U378 = ~new_P2_R1077_U377 | ~new_P2_R1077_U376;
  assign new_P2_R1077_U379 = ~new_P2_R1077_U353 | ~new_P2_R1077_U144;
  assign new_P2_R1077_U380 = ~new_P2_R1077_U203 | ~new_P2_R1077_U378;
  assign new_P2_R1077_U381 = ~new_P2_U3069 | ~new_P2_R1077_U23;
  assign new_P2_R1077_U382 = ~new_P2_U3410 | ~new_P2_R1077_U21;
  assign new_P2_R1077_U383 = ~new_P2_U3070 | ~new_P2_R1077_U19;
  assign new_P2_R1077_U384 = ~new_P2_U3407 | ~new_P2_R1077_U20;
  assign new_P2_R1077_U385 = ~new_P2_R1077_U384 | ~new_P2_R1077_U383;
  assign new_P2_R1077_U386 = ~new_P2_R1077_U354 | ~new_P2_R1077_U41;
  assign new_P2_R1077_U387 = ~new_P2_R1077_U385 | ~new_P2_R1077_U195;
  assign new_P2_R1077_U388 = ~new_P2_U3066 | ~new_P2_R1077_U35;
  assign new_P2_R1077_U389 = ~new_P2_U3404 | ~new_P2_R1077_U26;
  assign new_P2_R1077_U390 = ~new_P2_U3059 | ~new_P2_R1077_U24;
  assign new_P2_R1077_U391 = ~new_P2_U3401 | ~new_P2_R1077_U25;
  assign new_P2_R1077_U392 = ~new_P2_R1077_U391 | ~new_P2_R1077_U390;
  assign new_P2_R1077_U393 = ~new_P2_R1077_U355 | ~new_P2_R1077_U44;
  assign new_P2_R1077_U394 = ~new_P2_R1077_U392 | ~new_P2_R1077_U221;
  assign new_P2_R1077_U395 = ~new_P2_U3063 | ~new_P2_R1077_U32;
  assign new_P2_R1077_U396 = ~new_P2_U3398 | ~new_P2_R1077_U33;
  assign new_P2_R1077_U397 = ~new_P2_R1077_U396 | ~new_P2_R1077_U395;
  assign new_P2_R1077_U398 = ~new_P2_R1077_U356 | ~new_P2_R1077_U145;
  assign new_P2_R1077_U399 = ~new_P2_R1077_U230 | ~new_P2_R1077_U397;
  assign new_P2_R1077_U400 = ~new_P2_U3067 | ~new_P2_R1077_U27;
  assign new_P2_R1077_U401 = ~new_P2_U3395 | ~new_P2_R1077_U28;
  assign new_P2_R1077_U402 = ~new_P2_U3054 | ~new_P2_R1077_U147;
  assign new_P2_R1077_U403 = ~new_P2_U3904 | ~new_P2_R1077_U146;
  assign new_P2_R1077_U404 = ~new_P2_U3054 | ~new_P2_R1077_U147;
  assign new_P2_R1077_U405 = ~new_P2_U3904 | ~new_P2_R1077_U146;
  assign new_P2_R1077_U406 = ~new_P2_R1077_U405 | ~new_P2_R1077_U404;
  assign new_P2_R1077_U407 = ~new_P2_R1077_U148 | ~new_P2_R1077_U149;
  assign new_P2_R1077_U408 = ~new_P2_R1077_U305 | ~new_P2_R1077_U406;
  assign new_P2_R1077_U409 = ~new_P2_U3053 | ~new_P2_R1077_U88;
  assign new_P2_R1077_U410 = ~new_P2_U3895 | ~new_P2_R1077_U87;
  assign new_P2_R1077_U411 = ~new_P2_U3053 | ~new_P2_R1077_U88;
  assign new_P2_R1077_U412 = ~new_P2_U3895 | ~new_P2_R1077_U87;
  assign new_P2_R1077_U413 = ~new_P2_R1077_U412 | ~new_P2_R1077_U411;
  assign new_P2_R1077_U414 = ~new_P2_R1077_U150 | ~new_P2_R1077_U151;
  assign new_P2_R1077_U415 = ~new_P2_R1077_U303 | ~new_P2_R1077_U413;
  assign new_P2_R1077_U416 = ~new_P2_U3052 | ~new_P2_R1077_U46;
  assign new_P2_R1077_U417 = ~new_P2_U3896 | ~new_P2_R1077_U47;
  assign new_P2_R1077_U418 = ~new_P2_U3052 | ~new_P2_R1077_U46;
  assign new_P2_R1077_U419 = ~new_P2_U3896 | ~new_P2_R1077_U47;
  assign new_P2_R1077_U420 = ~new_P2_R1077_U419 | ~new_P2_R1077_U418;
  assign new_P2_R1077_U421 = ~new_P2_R1077_U152 | ~new_P2_R1077_U153;
  assign new_P2_R1077_U422 = ~new_P2_R1077_U300 | ~new_P2_R1077_U420;
  assign new_P2_R1077_U423 = ~new_P2_U3056 | ~new_P2_R1077_U49;
  assign new_P2_R1077_U424 = ~new_P2_U3897 | ~new_P2_R1077_U48;
  assign new_P2_R1077_U425 = ~new_P2_U3057 | ~new_P2_R1077_U50;
  assign new_P2_R1077_U426 = ~new_P2_U3898 | ~new_P2_R1077_U51;
  assign new_P2_R1077_U427 = ~new_P2_R1077_U426 | ~new_P2_R1077_U425;
  assign new_P2_R1077_U428 = ~new_P2_R1077_U357 | ~new_P2_R1077_U89;
  assign new_P2_R1077_U429 = ~new_P2_R1077_U427 | ~new_P2_R1077_U307;
  assign new_P2_R1077_U430 = ~new_P2_U3064 | ~new_P2_R1077_U52;
  assign new_P2_R1077_U431 = ~new_P2_U3899 | ~new_P2_R1077_U53;
  assign new_P2_R1077_U432 = ~new_P2_R1077_U431 | ~new_P2_R1077_U430;
  assign new_P2_R1077_U433 = ~new_P2_R1077_U358 | ~new_P2_R1077_U155;
  assign new_P2_R1077_U434 = ~new_P2_R1077_U294 | ~new_P2_R1077_U432;
  assign new_P2_R1077_U435 = ~new_P2_U3065 | ~new_P2_R1077_U84;
  assign new_P2_R1077_U436 = ~new_P2_U3900 | ~new_P2_R1077_U85;
  assign new_P2_R1077_U437 = ~new_P2_U3065 | ~new_P2_R1077_U84;
  assign new_P2_R1077_U438 = ~new_P2_U3900 | ~new_P2_R1077_U85;
  assign new_P2_R1077_U439 = ~new_P2_R1077_U438 | ~new_P2_R1077_U437;
  assign new_P2_R1077_U440 = ~new_P2_R1077_U156 | ~new_P2_R1077_U157;
  assign new_P2_R1077_U441 = ~new_P2_R1077_U290 | ~new_P2_R1077_U439;
  assign new_P2_R1077_U442 = ~new_P2_U3060 | ~new_P2_R1077_U82;
  assign new_P2_R1077_U443 = ~new_P2_U3901 | ~new_P2_R1077_U83;
  assign new_P2_R1077_U444 = ~new_P2_U3060 | ~new_P2_R1077_U82;
  assign new_P2_R1077_U445 = ~new_P2_U3901 | ~new_P2_R1077_U83;
  assign new_P2_R1077_U446 = ~new_P2_R1077_U445 | ~new_P2_R1077_U444;
  assign new_P2_R1077_U447 = ~new_P2_R1077_U158 | ~new_P2_R1077_U159;
  assign new_P2_R1077_U448 = ~new_P2_R1077_U286 | ~new_P2_R1077_U446;
  assign new_P2_R1077_U449 = ~new_P2_U3074 | ~new_P2_R1077_U54;
  assign new_P2_R1077_U450 = ~new_P2_U3902 | ~new_P2_R1077_U55;
  assign new_P2_R1077_U451 = ~new_P2_U3074 | ~new_P2_R1077_U54;
  assign new_P2_R1077_U452 = ~new_P2_U3902 | ~new_P2_R1077_U55;
  assign new_P2_R1077_U453 = ~new_P2_R1077_U452 | ~new_P2_R1077_U451;
  assign new_P2_R1077_U454 = ~new_P2_U3075 | ~new_P2_R1077_U81;
  assign new_P2_R1077_U455 = ~new_P2_U3903 | ~new_P2_R1077_U90;
  assign new_P2_R1077_U456 = ~new_P2_R1077_U182 | ~new_P2_R1077_U161;
  assign new_P2_R1077_U457 = ~new_P2_R1077_U328 | ~new_P2_R1077_U31;
  assign new_P2_R1077_U458 = ~new_P2_U3080 | ~new_P2_R1077_U78;
  assign new_P2_R1077_U459 = ~new_P2_U3445 | ~new_P2_R1077_U79;
  assign new_P2_R1077_U460 = ~new_P2_R1077_U459 | ~new_P2_R1077_U458;
  assign new_P2_R1077_U461 = ~new_P2_R1077_U359 | ~new_P2_R1077_U91;
  assign new_P2_R1077_U462 = ~new_P2_R1077_U460 | ~new_P2_R1077_U316;
  assign new_P2_R1077_U463 = ~new_P2_U3081 | ~new_P2_R1077_U75;
  assign new_P2_R1077_U464 = ~new_P2_U3443 | ~new_P2_R1077_U76;
  assign new_P2_R1077_U465 = ~new_P2_R1077_U464 | ~new_P2_R1077_U463;
  assign new_P2_R1077_U466 = ~new_P2_R1077_U360 | ~new_P2_R1077_U162;
  assign new_P2_R1077_U467 = ~new_P2_R1077_U270 | ~new_P2_R1077_U465;
  assign new_P2_R1077_U468 = ~new_P2_U3068 | ~new_P2_R1077_U60;
  assign new_P2_R1077_U469 = ~new_P2_U3440 | ~new_P2_R1077_U58;
  assign new_P2_R1077_U470 = ~new_P2_U3072 | ~new_P2_R1077_U56;
  assign new_P2_R1077_U471 = ~new_P2_U3437 | ~new_P2_R1077_U57;
  assign new_P2_R1077_U472 = ~new_P2_R1077_U471 | ~new_P2_R1077_U470;
  assign new_P2_R1077_U473 = ~new_P2_R1077_U361 | ~new_P2_R1077_U92;
  assign new_P2_R1077_U474 = ~new_P2_R1077_U472 | ~new_P2_R1077_U262;
  assign new_P2_R1077_U475 = ~new_P2_U3073 | ~new_P2_R1077_U73;
  assign new_P2_R1077_U476 = ~new_P2_U3434 | ~new_P2_R1077_U74;
  assign new_P2_R1077_U477 = ~new_P2_U3073 | ~new_P2_R1077_U73;
  assign new_P2_R1077_U478 = ~new_P2_U3434 | ~new_P2_R1077_U74;
  assign new_P2_R1077_U479 = ~new_P2_R1077_U478 | ~new_P2_R1077_U477;
  assign new_P2_R1077_U480 = ~new_P2_R1077_U163 | ~new_P2_R1077_U164;
  assign new_P2_R1077_U481 = ~new_P2_R1077_U258 | ~new_P2_R1077_U479;
  assign new_P2_R1077_U482 = ~new_P2_U3078 | ~new_P2_R1077_U71;
  assign new_P2_R1077_U483 = ~new_P2_U3431 | ~new_P2_R1077_U72;
  assign new_P2_R1077_U484 = ~new_P2_U3078 | ~new_P2_R1077_U71;
  assign new_P2_R1077_U485 = ~new_P2_U3431 | ~new_P2_R1077_U72;
  assign new_P2_R1077_U486 = ~new_P2_R1077_U485 | ~new_P2_R1077_U484;
  assign new_P2_R1077_U487 = ~new_P2_R1077_U165 | ~new_P2_R1077_U166;
  assign new_P2_R1077_U488 = ~new_P2_R1077_U254 | ~new_P2_R1077_U486;
  assign new_P2_R1077_U489 = ~new_P2_U3079 | ~new_P2_R1077_U61;
  assign new_P2_R1077_U490 = ~new_P2_U3428 | ~new_P2_R1077_U62;
  assign new_P2_R1077_U491 = ~new_P2_U3071 | ~new_P2_R1077_U69;
  assign new_P2_R1077_U492 = ~new_P2_U3425 | ~new_P2_R1077_U70;
  assign new_P2_R1077_U493 = ~new_P2_R1077_U492 | ~new_P2_R1077_U491;
  assign new_P2_R1077_U494 = ~new_P2_R1077_U362 | ~new_P2_R1077_U93;
  assign new_P2_R1077_U495 = ~new_P2_R1077_U493 | ~new_P2_R1077_U338;
  assign new_P2_R1077_U496 = ~new_P2_U3062 | ~new_P2_R1077_U66;
  assign new_P2_R1077_U497 = ~new_P2_U3422 | ~new_P2_R1077_U67;
  assign new_P2_R1077_U498 = ~new_P2_R1077_U497 | ~new_P2_R1077_U496;
  assign new_P2_R1077_U499 = ~new_P2_R1077_U363 | ~new_P2_R1077_U167;
  assign new_P2_R1077_U500 = ~new_P2_R1077_U244 | ~new_P2_R1077_U498;
  assign new_P2_R1077_U501 = ~new_P2_U3061 | ~new_P2_R1077_U63;
  assign new_P2_R1077_U502 = ~new_P2_U3419 | ~new_P2_R1077_U64;
  assign new_P2_R1077_U503 = ~new_P2_U3076 | ~new_P2_R1077_U29;
  assign new_P2_R1077_U504 = ~new_P2_U3387 | ~new_P2_R1077_U30;
  assign new_P2_R1143_U4 = new_P2_R1143_U179 & new_P2_R1143_U178;
  assign new_P2_R1143_U5 = new_P2_R1143_U197 & new_P2_R1143_U196;
  assign new_P2_R1143_U6 = new_P2_R1143_U237 & new_P2_R1143_U236;
  assign new_P2_R1143_U7 = new_P2_R1143_U246 & new_P2_R1143_U245;
  assign new_P2_R1143_U8 = new_P2_R1143_U264 & new_P2_R1143_U263;
  assign new_P2_R1143_U9 = new_P2_R1143_U272 & new_P2_R1143_U271;
  assign new_P2_R1143_U10 = new_P2_R1143_U351 & new_P2_R1143_U348;
  assign new_P2_R1143_U11 = new_P2_R1143_U344 & new_P2_R1143_U341;
  assign new_P2_R1143_U12 = new_P2_R1143_U335 & new_P2_R1143_U332;
  assign new_P2_R1143_U13 = new_P2_R1143_U326 & new_P2_R1143_U323;
  assign new_P2_R1143_U14 = new_P2_R1143_U320 & new_P2_R1143_U318;
  assign new_P2_R1143_U15 = new_P2_R1143_U313 & new_P2_R1143_U310;
  assign new_P2_R1143_U16 = new_P2_R1143_U235 & new_P2_R1143_U232;
  assign new_P2_R1143_U17 = new_P2_R1143_U227 & new_P2_R1143_U224;
  assign new_P2_R1143_U18 = new_P2_R1143_U213 & new_P2_R1143_U210;
  assign new_P2_R1143_U19 = ~new_P2_U3407;
  assign new_P2_R1143_U20 = ~new_P2_U3070;
  assign new_P2_R1143_U21 = ~new_P2_U3069;
  assign new_P2_R1143_U22 = ~new_P2_U3070 | ~new_P2_U3407;
  assign new_P2_R1143_U23 = ~new_P2_U3410;
  assign new_P2_R1143_U24 = ~new_P2_U3401;
  assign new_P2_R1143_U25 = ~new_P2_U3059;
  assign new_P2_R1143_U26 = ~new_P2_U3066;
  assign new_P2_R1143_U27 = ~new_P2_U3395;
  assign new_P2_R1143_U28 = ~new_P2_U3067;
  assign new_P2_R1143_U29 = ~new_P2_U3387;
  assign new_P2_R1143_U30 = ~new_P2_U3076;
  assign new_P2_R1143_U31 = ~new_P2_U3076 | ~new_P2_U3387;
  assign new_P2_R1143_U32 = ~new_P2_U3398;
  assign new_P2_R1143_U33 = ~new_P2_U3063;
  assign new_P2_R1143_U34 = ~new_P2_U3059 | ~new_P2_U3401;
  assign new_P2_R1143_U35 = ~new_P2_U3404;
  assign new_P2_R1143_U36 = ~new_P2_U3413;
  assign new_P2_R1143_U37 = ~new_P2_U3083;
  assign new_P2_R1143_U38 = ~new_P2_U3082;
  assign new_P2_R1143_U39 = ~new_P2_U3416;
  assign new_P2_R1143_U40 = ~new_P2_R1143_U65 | ~new_P2_R1143_U205;
  assign new_P2_R1143_U41 = ~new_P2_R1143_U117 | ~new_P2_R1143_U193;
  assign new_P2_R1143_U42 = ~new_P2_R1143_U182 | ~new_P2_R1143_U183;
  assign new_P2_R1143_U43 = ~new_P2_U3392 | ~new_P2_U3077;
  assign new_P2_R1143_U44 = ~new_P2_R1143_U122 | ~new_P2_R1143_U219;
  assign new_P2_R1143_U45 = ~new_P2_R1143_U216 | ~new_P2_R1143_U215;
  assign new_P2_R1143_U46 = ~new_P2_U3896;
  assign new_P2_R1143_U47 = ~new_P2_U3052;
  assign new_P2_R1143_U48 = ~new_P2_U3056;
  assign new_P2_R1143_U49 = ~new_P2_U3897;
  assign new_P2_R1143_U50 = ~new_P2_U3898;
  assign new_P2_R1143_U51 = ~new_P2_U3057;
  assign new_P2_R1143_U52 = ~new_P2_U3899;
  assign new_P2_R1143_U53 = ~new_P2_U3064;
  assign new_P2_R1143_U54 = ~new_P2_U3902;
  assign new_P2_R1143_U55 = ~new_P2_U3074;
  assign new_P2_R1143_U56 = ~new_P2_U3437;
  assign new_P2_R1143_U57 = ~new_P2_U3072;
  assign new_P2_R1143_U58 = ~new_P2_U3068;
  assign new_P2_R1143_U59 = ~new_P2_U3072 | ~new_P2_U3437;
  assign new_P2_R1143_U60 = ~new_P2_U3440;
  assign new_P2_R1143_U61 = ~new_P2_U3428;
  assign new_P2_R1143_U62 = ~new_P2_U3079;
  assign new_P2_R1143_U63 = ~new_P2_U3419;
  assign new_P2_R1143_U64 = ~new_P2_U3061;
  assign new_P2_R1143_U65 = ~new_P2_U3083 | ~new_P2_U3413;
  assign new_P2_R1143_U66 = ~new_P2_U3422;
  assign new_P2_R1143_U67 = ~new_P2_U3062;
  assign new_P2_R1143_U68 = ~new_P2_U3062 | ~new_P2_U3422;
  assign new_P2_R1143_U69 = ~new_P2_U3425;
  assign new_P2_R1143_U70 = ~new_P2_U3071;
  assign new_P2_R1143_U71 = ~new_P2_U3431;
  assign new_P2_R1143_U72 = ~new_P2_U3078;
  assign new_P2_R1143_U73 = ~new_P2_U3434;
  assign new_P2_R1143_U74 = ~new_P2_U3073;
  assign new_P2_R1143_U75 = ~new_P2_U3443;
  assign new_P2_R1143_U76 = ~new_P2_U3081;
  assign new_P2_R1143_U77 = ~new_P2_U3081 | ~new_P2_U3443;
  assign new_P2_R1143_U78 = ~new_P2_U3445;
  assign new_P2_R1143_U79 = ~new_P2_U3080;
  assign new_P2_R1143_U80 = ~new_P2_U3080 | ~new_P2_U3445;
  assign new_P2_R1143_U81 = ~new_P2_U3903;
  assign new_P2_R1143_U82 = ~new_P2_U3901;
  assign new_P2_R1143_U83 = ~new_P2_U3060;
  assign new_P2_R1143_U84 = ~new_P2_U3900;
  assign new_P2_R1143_U85 = ~new_P2_U3065;
  assign new_P2_R1143_U86 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1143_U87 = ~new_P2_U3053;
  assign new_P2_R1143_U88 = ~new_P2_U3895;
  assign new_P2_R1143_U89 = ~new_P2_R1143_U306 | ~new_P2_R1143_U176;
  assign new_P2_R1143_U90 = ~new_P2_U3075;
  assign new_P2_R1143_U91 = ~new_P2_R1143_U77 | ~new_P2_R1143_U315;
  assign new_P2_R1143_U92 = ~new_P2_R1143_U261 | ~new_P2_R1143_U260;
  assign new_P2_R1143_U93 = ~new_P2_R1143_U68 | ~new_P2_R1143_U337;
  assign new_P2_R1143_U94 = ~new_P2_R1143_U457 | ~new_P2_R1143_U456;
  assign new_P2_R1143_U95 = ~new_P2_R1143_U504 | ~new_P2_R1143_U503;
  assign new_P2_R1143_U96 = ~new_P2_R1143_U375 | ~new_P2_R1143_U374;
  assign new_P2_R1143_U97 = ~new_P2_R1143_U380 | ~new_P2_R1143_U379;
  assign new_P2_R1143_U98 = ~new_P2_R1143_U387 | ~new_P2_R1143_U386;
  assign new_P2_R1143_U99 = ~new_P2_R1143_U394 | ~new_P2_R1143_U393;
  assign new_P2_R1143_U100 = ~new_P2_R1143_U399 | ~new_P2_R1143_U398;
  assign new_P2_R1143_U101 = ~new_P2_R1143_U408 | ~new_P2_R1143_U407;
  assign new_P2_R1143_U102 = ~new_P2_R1143_U415 | ~new_P2_R1143_U414;
  assign new_P2_R1143_U103 = ~new_P2_R1143_U422 | ~new_P2_R1143_U421;
  assign new_P2_R1143_U104 = ~new_P2_R1143_U429 | ~new_P2_R1143_U428;
  assign new_P2_R1143_U105 = ~new_P2_R1143_U434 | ~new_P2_R1143_U433;
  assign new_P2_R1143_U106 = ~new_P2_R1143_U441 | ~new_P2_R1143_U440;
  assign new_P2_R1143_U107 = ~new_P2_R1143_U448 | ~new_P2_R1143_U447;
  assign new_P2_R1143_U108 = ~new_P2_R1143_U462 | ~new_P2_R1143_U461;
  assign new_P2_R1143_U109 = ~new_P2_R1143_U467 | ~new_P2_R1143_U466;
  assign new_P2_R1143_U110 = ~new_P2_R1143_U474 | ~new_P2_R1143_U473;
  assign new_P2_R1143_U111 = ~new_P2_R1143_U481 | ~new_P2_R1143_U480;
  assign new_P2_R1143_U112 = ~new_P2_R1143_U488 | ~new_P2_R1143_U487;
  assign new_P2_R1143_U113 = ~new_P2_R1143_U495 | ~new_P2_R1143_U494;
  assign new_P2_R1143_U114 = ~new_P2_R1143_U500 | ~new_P2_R1143_U499;
  assign new_P2_R1143_U115 = new_P2_R1143_U189 & new_P2_R1143_U187;
  assign new_P2_R1143_U116 = new_P2_R1143_U4 & new_P2_R1143_U180;
  assign new_P2_R1143_U117 = new_P2_R1143_U194 & new_P2_R1143_U192;
  assign new_P2_R1143_U118 = new_P2_R1143_U201 & new_P2_R1143_U200;
  assign new_P2_R1143_U119 = new_P2_R1143_U22 & new_P2_R1143_U382 & new_P2_R1143_U381;
  assign new_P2_R1143_U120 = new_P2_R1143_U212 & new_P2_R1143_U5;
  assign new_P2_R1143_U121 = new_P2_R1143_U181 & new_P2_R1143_U180;
  assign new_P2_R1143_U122 = new_P2_R1143_U220 & new_P2_R1143_U218;
  assign new_P2_R1143_U123 = new_P2_R1143_U34 & new_P2_R1143_U389 & new_P2_R1143_U388;
  assign new_P2_R1143_U124 = new_P2_R1143_U226 & new_P2_R1143_U4;
  assign new_P2_R1143_U125 = new_P2_R1143_U234 & new_P2_R1143_U181;
  assign new_P2_R1143_U126 = new_P2_R1143_U204 & new_P2_R1143_U6;
  assign new_P2_R1143_U127 = new_P2_R1143_U243 & new_P2_R1143_U239;
  assign new_P2_R1143_U128 = new_P2_R1143_U250 & new_P2_R1143_U7;
  assign new_P2_R1143_U129 = new_P2_R1143_U253 & new_P2_R1143_U248;
  assign new_P2_R1143_U130 = new_P2_R1143_U268 & new_P2_R1143_U267;
  assign new_P2_R1143_U131 = new_P2_R1143_U9 & new_P2_R1143_U282;
  assign new_P2_R1143_U132 = new_P2_R1143_U285 & new_P2_R1143_U280;
  assign new_P2_R1143_U133 = new_P2_R1143_U301 & new_P2_R1143_U298;
  assign new_P2_R1143_U134 = new_P2_R1143_U368 & new_P2_R1143_U302;
  assign new_P2_R1143_U135 = new_P2_R1143_U160 & new_P2_R1143_U278;
  assign new_P2_R1143_U136 = new_P2_R1143_U80 & new_P2_R1143_U455 & new_P2_R1143_U454;
  assign new_P2_R1143_U137 = new_P2_R1143_U325 & new_P2_R1143_U9;
  assign new_P2_R1143_U138 = new_P2_R1143_U59 & new_P2_R1143_U469 & new_P2_R1143_U468;
  assign new_P2_R1143_U139 = new_P2_R1143_U334 & new_P2_R1143_U8;
  assign new_P2_R1143_U140 = new_P2_R1143_U172 & new_P2_R1143_U490 & new_P2_R1143_U489;
  assign new_P2_R1143_U141 = new_P2_R1143_U343 & new_P2_R1143_U7;
  assign new_P2_R1143_U142 = new_P2_R1143_U171 & new_P2_R1143_U502 & new_P2_R1143_U501;
  assign new_P2_R1143_U143 = new_P2_R1143_U350 & new_P2_R1143_U6;
  assign new_P2_R1143_U144 = ~new_P2_R1143_U118 | ~new_P2_R1143_U202;
  assign new_P2_R1143_U145 = ~new_P2_R1143_U217 | ~new_P2_R1143_U229;
  assign new_P2_R1143_U146 = ~new_P2_U3054;
  assign new_P2_R1143_U147 = ~new_P2_U3904;
  assign new_P2_R1143_U148 = new_P2_R1143_U403 & new_P2_R1143_U402;
  assign new_P2_R1143_U149 = ~new_P2_R1143_U364 | ~new_P2_R1143_U304 | ~new_P2_R1143_U169;
  assign new_P2_R1143_U150 = new_P2_R1143_U410 & new_P2_R1143_U409;
  assign new_P2_R1143_U151 = ~new_P2_R1143_U134 | ~new_P2_R1143_U370 | ~new_P2_R1143_U369;
  assign new_P2_R1143_U152 = new_P2_R1143_U417 & new_P2_R1143_U416;
  assign new_P2_R1143_U153 = ~new_P2_R1143_U86 | ~new_P2_R1143_U365 | ~new_P2_R1143_U299;
  assign new_P2_R1143_U154 = new_P2_R1143_U424 & new_P2_R1143_U423;
  assign new_P2_R1143_U155 = ~new_P2_R1143_U293 | ~new_P2_R1143_U292;
  assign new_P2_R1143_U156 = new_P2_R1143_U436 & new_P2_R1143_U435;
  assign new_P2_R1143_U157 = ~new_P2_R1143_U289 | ~new_P2_R1143_U288;
  assign new_P2_R1143_U158 = new_P2_R1143_U443 & new_P2_R1143_U442;
  assign new_P2_R1143_U159 = ~new_P2_R1143_U132 | ~new_P2_R1143_U284;
  assign new_P2_R1143_U160 = new_P2_R1143_U450 & new_P2_R1143_U449;
  assign new_P2_R1143_U161 = ~new_P2_R1143_U43 | ~new_P2_R1143_U327;
  assign new_P2_R1143_U162 = ~new_P2_R1143_U130 | ~new_P2_R1143_U269;
  assign new_P2_R1143_U163 = new_P2_R1143_U476 & new_P2_R1143_U475;
  assign new_P2_R1143_U164 = ~new_P2_R1143_U257 | ~new_P2_R1143_U256;
  assign new_P2_R1143_U165 = new_P2_R1143_U483 & new_P2_R1143_U482;
  assign new_P2_R1143_U166 = ~new_P2_R1143_U129 | ~new_P2_R1143_U252;
  assign new_P2_R1143_U167 = ~new_P2_R1143_U127 | ~new_P2_R1143_U242;
  assign new_P2_R1143_U168 = ~new_P2_R1143_U367 | ~new_P2_R1143_U366;
  assign new_P2_R1143_U169 = ~new_P2_U3053 | ~new_P2_R1143_U151;
  assign new_P2_R1143_U170 = ~new_P2_R1143_U34;
  assign new_P2_R1143_U171 = ~new_P2_U3416 | ~new_P2_U3082;
  assign new_P2_R1143_U172 = ~new_P2_U3071 | ~new_P2_U3425;
  assign new_P2_R1143_U173 = ~new_P2_U3057 | ~new_P2_U3898;
  assign new_P2_R1143_U174 = ~new_P2_R1143_U68;
  assign new_P2_R1143_U175 = ~new_P2_R1143_U77;
  assign new_P2_R1143_U176 = ~new_P2_U3064 | ~new_P2_U3899;
  assign new_P2_R1143_U177 = ~new_P2_R1143_U65;
  assign new_P2_R1143_U178 = new_P2_U3066 | new_P2_U3404;
  assign new_P2_R1143_U179 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1143_U180 = new_P2_U3398 | new_P2_U3063;
  assign new_P2_R1143_U181 = new_P2_U3395 | new_P2_U3067;
  assign new_P2_R1143_U182 = ~new_P2_R1143_U31;
  assign new_P2_R1143_U183 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1143_U184 = ~new_P2_R1143_U42;
  assign new_P2_R1143_U185 = ~new_P2_R1143_U43;
  assign new_P2_R1143_U186 = ~new_P2_R1143_U42 | ~new_P2_R1143_U43;
  assign new_P2_R1143_U187 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1143_U188 = ~new_P2_R1143_U186 | ~new_P2_R1143_U181;
  assign new_P2_R1143_U189 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1143_U190 = ~new_P2_R1143_U115 | ~new_P2_R1143_U188;
  assign new_P2_R1143_U191 = ~new_P2_R1143_U35 | ~new_P2_R1143_U34;
  assign new_P2_R1143_U192 = ~new_P2_U3066 | ~new_P2_R1143_U191;
  assign new_P2_R1143_U193 = ~new_P2_R1143_U116 | ~new_P2_R1143_U190;
  assign new_P2_R1143_U194 = ~new_P2_U3404 | ~new_P2_R1143_U170;
  assign new_P2_R1143_U195 = ~new_P2_R1143_U41;
  assign new_P2_R1143_U196 = new_P2_U3069 | new_P2_U3410;
  assign new_P2_R1143_U197 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1143_U198 = ~new_P2_R1143_U22;
  assign new_P2_R1143_U199 = ~new_P2_R1143_U23 | ~new_P2_R1143_U22;
  assign new_P2_R1143_U200 = ~new_P2_U3069 | ~new_P2_R1143_U199;
  assign new_P2_R1143_U201 = ~new_P2_U3410 | ~new_P2_R1143_U198;
  assign new_P2_R1143_U202 = ~new_P2_R1143_U5 | ~new_P2_R1143_U41;
  assign new_P2_R1143_U203 = ~new_P2_R1143_U144;
  assign new_P2_R1143_U204 = new_P2_U3413 | new_P2_U3083;
  assign new_P2_R1143_U205 = ~new_P2_R1143_U204 | ~new_P2_R1143_U144;
  assign new_P2_R1143_U206 = ~new_P2_R1143_U40;
  assign new_P2_R1143_U207 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1143_U208 = new_P2_U3407 | new_P2_U3070;
  assign new_P2_R1143_U209 = ~new_P2_R1143_U208 | ~new_P2_R1143_U41;
  assign new_P2_R1143_U210 = ~new_P2_R1143_U119 | ~new_P2_R1143_U209;
  assign new_P2_R1143_U211 = ~new_P2_R1143_U195 | ~new_P2_R1143_U22;
  assign new_P2_R1143_U212 = ~new_P2_U3410 | ~new_P2_U3069;
  assign new_P2_R1143_U213 = ~new_P2_R1143_U120 | ~new_P2_R1143_U211;
  assign new_P2_R1143_U214 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1143_U215 = ~new_P2_R1143_U185 | ~new_P2_R1143_U181;
  assign new_P2_R1143_U216 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1143_U217 = ~new_P2_R1143_U45;
  assign new_P2_R1143_U218 = ~new_P2_R1143_U121 | ~new_P2_R1143_U184;
  assign new_P2_R1143_U219 = ~new_P2_R1143_U45 | ~new_P2_R1143_U180;
  assign new_P2_R1143_U220 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1143_U221 = ~new_P2_R1143_U44;
  assign new_P2_R1143_U222 = new_P2_U3401 | new_P2_U3059;
  assign new_P2_R1143_U223 = ~new_P2_R1143_U222 | ~new_P2_R1143_U44;
  assign new_P2_R1143_U224 = ~new_P2_R1143_U123 | ~new_P2_R1143_U223;
  assign new_P2_R1143_U225 = ~new_P2_R1143_U221 | ~new_P2_R1143_U34;
  assign new_P2_R1143_U226 = ~new_P2_U3404 | ~new_P2_U3066;
  assign new_P2_R1143_U227 = ~new_P2_R1143_U124 | ~new_P2_R1143_U225;
  assign new_P2_R1143_U228 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1143_U229 = ~new_P2_R1143_U184 | ~new_P2_R1143_U181;
  assign new_P2_R1143_U230 = ~new_P2_R1143_U145;
  assign new_P2_R1143_U231 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1143_U232 = ~new_P2_R1143_U42 | ~new_P2_R1143_U43 | ~new_P2_R1143_U401 | ~new_P2_R1143_U400;
  assign new_P2_R1143_U233 = ~new_P2_R1143_U43 | ~new_P2_R1143_U42;
  assign new_P2_R1143_U234 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1143_U235 = ~new_P2_R1143_U125 | ~new_P2_R1143_U233;
  assign new_P2_R1143_U236 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1143_U237 = new_P2_U3061 | new_P2_U3419;
  assign new_P2_R1143_U238 = ~new_P2_R1143_U177 | ~new_P2_R1143_U6;
  assign new_P2_R1143_U239 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1143_U240 = ~new_P2_R1143_U171 | ~new_P2_R1143_U238;
  assign new_P2_R1143_U241 = new_P2_U3419 | new_P2_U3061;
  assign new_P2_R1143_U242 = ~new_P2_R1143_U126 | ~new_P2_R1143_U144;
  assign new_P2_R1143_U243 = ~new_P2_R1143_U241 | ~new_P2_R1143_U240;
  assign new_P2_R1143_U244 = ~new_P2_R1143_U167;
  assign new_P2_R1143_U245 = new_P2_U3079 | new_P2_U3428;
  assign new_P2_R1143_U246 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1143_U247 = ~new_P2_R1143_U174 | ~new_P2_R1143_U7;
  assign new_P2_R1143_U248 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1143_U249 = ~new_P2_R1143_U172 | ~new_P2_R1143_U247;
  assign new_P2_R1143_U250 = new_P2_U3422 | new_P2_U3062;
  assign new_P2_R1143_U251 = new_P2_U3428 | new_P2_U3079;
  assign new_P2_R1143_U252 = ~new_P2_R1143_U128 | ~new_P2_R1143_U167;
  assign new_P2_R1143_U253 = ~new_P2_R1143_U251 | ~new_P2_R1143_U249;
  assign new_P2_R1143_U254 = ~new_P2_R1143_U166;
  assign new_P2_R1143_U255 = new_P2_U3431 | new_P2_U3078;
  assign new_P2_R1143_U256 = ~new_P2_R1143_U255 | ~new_P2_R1143_U166;
  assign new_P2_R1143_U257 = ~new_P2_U3078 | ~new_P2_U3431;
  assign new_P2_R1143_U258 = ~new_P2_R1143_U164;
  assign new_P2_R1143_U259 = new_P2_U3434 | new_P2_U3073;
  assign new_P2_R1143_U260 = ~new_P2_R1143_U259 | ~new_P2_R1143_U164;
  assign new_P2_R1143_U261 = ~new_P2_U3073 | ~new_P2_U3434;
  assign new_P2_R1143_U262 = ~new_P2_R1143_U92;
  assign new_P2_R1143_U263 = new_P2_U3068 | new_P2_U3440;
  assign new_P2_R1143_U264 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1143_U265 = ~new_P2_R1143_U59;
  assign new_P2_R1143_U266 = ~new_P2_R1143_U60 | ~new_P2_R1143_U59;
  assign new_P2_R1143_U267 = ~new_P2_U3068 | ~new_P2_R1143_U266;
  assign new_P2_R1143_U268 = ~new_P2_U3440 | ~new_P2_R1143_U265;
  assign new_P2_R1143_U269 = ~new_P2_R1143_U8 | ~new_P2_R1143_U92;
  assign new_P2_R1143_U270 = ~new_P2_R1143_U162;
  assign new_P2_R1143_U271 = new_P2_U3075 | new_P2_U3903;
  assign new_P2_R1143_U272 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1143_U273 = new_P2_U3074 | new_P2_U3902;
  assign new_P2_R1143_U274 = ~new_P2_R1143_U80;
  assign new_P2_R1143_U275 = ~new_P2_U3903 | ~new_P2_R1143_U274;
  assign new_P2_R1143_U276 = ~new_P2_R1143_U275 | ~new_P2_R1143_U90;
  assign new_P2_R1143_U277 = ~new_P2_R1143_U80 | ~new_P2_R1143_U81;
  assign new_P2_R1143_U278 = ~new_P2_R1143_U277 | ~new_P2_R1143_U276;
  assign new_P2_R1143_U279 = ~new_P2_R1143_U175 | ~new_P2_R1143_U9;
  assign new_P2_R1143_U280 = ~new_P2_U3074 | ~new_P2_U3902;
  assign new_P2_R1143_U281 = ~new_P2_R1143_U278 | ~new_P2_R1143_U279;
  assign new_P2_R1143_U282 = new_P2_U3443 | new_P2_U3081;
  assign new_P2_R1143_U283 = new_P2_U3902 | new_P2_U3074;
  assign new_P2_R1143_U284 = ~new_P2_R1143_U131 | ~new_P2_R1143_U273 | ~new_P2_R1143_U162;
  assign new_P2_R1143_U285 = ~new_P2_R1143_U283 | ~new_P2_R1143_U281;
  assign new_P2_R1143_U286 = ~new_P2_R1143_U159;
  assign new_P2_R1143_U287 = new_P2_U3901 | new_P2_U3060;
  assign new_P2_R1143_U288 = ~new_P2_R1143_U287 | ~new_P2_R1143_U159;
  assign new_P2_R1143_U289 = ~new_P2_U3060 | ~new_P2_U3901;
  assign new_P2_R1143_U290 = ~new_P2_R1143_U157;
  assign new_P2_R1143_U291 = new_P2_U3900 | new_P2_U3065;
  assign new_P2_R1143_U292 = ~new_P2_R1143_U291 | ~new_P2_R1143_U157;
  assign new_P2_R1143_U293 = ~new_P2_U3065 | ~new_P2_U3900;
  assign new_P2_R1143_U294 = ~new_P2_R1143_U155;
  assign new_P2_R1143_U295 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1143_U296 = ~new_P2_R1143_U176 | ~new_P2_R1143_U173;
  assign new_P2_R1143_U297 = ~new_P2_R1143_U86;
  assign new_P2_R1143_U298 = new_P2_U3899 | new_P2_U3064;
  assign new_P2_R1143_U299 = ~new_P2_R1143_U168 | ~new_P2_R1143_U155 | ~new_P2_R1143_U298;
  assign new_P2_R1143_U300 = ~new_P2_R1143_U153;
  assign new_P2_R1143_U301 = new_P2_U3896 | new_P2_U3052;
  assign new_P2_R1143_U302 = ~new_P2_U3052 | ~new_P2_U3896;
  assign new_P2_R1143_U303 = ~new_P2_R1143_U151;
  assign new_P2_R1143_U304 = ~new_P2_U3895 | ~new_P2_R1143_U151;
  assign new_P2_R1143_U305 = ~new_P2_R1143_U149;
  assign new_P2_R1143_U306 = ~new_P2_R1143_U298 | ~new_P2_R1143_U155;
  assign new_P2_R1143_U307 = ~new_P2_R1143_U89;
  assign new_P2_R1143_U308 = new_P2_U3898 | new_P2_U3057;
  assign new_P2_R1143_U309 = ~new_P2_R1143_U308 | ~new_P2_R1143_U89;
  assign new_P2_R1143_U310 = ~new_P2_R1143_U154 | ~new_P2_R1143_U309 | ~new_P2_R1143_U173;
  assign new_P2_R1143_U311 = ~new_P2_R1143_U307 | ~new_P2_R1143_U173;
  assign new_P2_R1143_U312 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1143_U313 = ~new_P2_R1143_U168 | ~new_P2_R1143_U311 | ~new_P2_R1143_U312;
  assign new_P2_R1143_U314 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1143_U315 = ~new_P2_R1143_U282 | ~new_P2_R1143_U162;
  assign new_P2_R1143_U316 = ~new_P2_R1143_U91;
  assign new_P2_R1143_U317 = ~new_P2_R1143_U9 | ~new_P2_R1143_U91;
  assign new_P2_R1143_U318 = ~new_P2_R1143_U135 | ~new_P2_R1143_U317;
  assign new_P2_R1143_U319 = ~new_P2_R1143_U317 | ~new_P2_R1143_U278;
  assign new_P2_R1143_U320 = ~new_P2_R1143_U453 | ~new_P2_R1143_U319;
  assign new_P2_R1143_U321 = new_P2_U3445 | new_P2_U3080;
  assign new_P2_R1143_U322 = ~new_P2_R1143_U321 | ~new_P2_R1143_U91;
  assign new_P2_R1143_U323 = ~new_P2_R1143_U136 | ~new_P2_R1143_U322;
  assign new_P2_R1143_U324 = ~new_P2_R1143_U316 | ~new_P2_R1143_U80;
  assign new_P2_R1143_U325 = ~new_P2_U3075 | ~new_P2_U3903;
  assign new_P2_R1143_U326 = ~new_P2_R1143_U137 | ~new_P2_R1143_U324;
  assign new_P2_R1143_U327 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1143_U328 = ~new_P2_R1143_U161;
  assign new_P2_R1143_U329 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1143_U330 = new_P2_U3437 | new_P2_U3072;
  assign new_P2_R1143_U331 = ~new_P2_R1143_U330 | ~new_P2_R1143_U92;
  assign new_P2_R1143_U332 = ~new_P2_R1143_U138 | ~new_P2_R1143_U331;
  assign new_P2_R1143_U333 = ~new_P2_R1143_U262 | ~new_P2_R1143_U59;
  assign new_P2_R1143_U334 = ~new_P2_U3440 | ~new_P2_U3068;
  assign new_P2_R1143_U335 = ~new_P2_R1143_U139 | ~new_P2_R1143_U333;
  assign new_P2_R1143_U336 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1143_U337 = ~new_P2_R1143_U250 | ~new_P2_R1143_U167;
  assign new_P2_R1143_U338 = ~new_P2_R1143_U93;
  assign new_P2_R1143_U339 = new_P2_U3425 | new_P2_U3071;
  assign new_P2_R1143_U340 = ~new_P2_R1143_U339 | ~new_P2_R1143_U93;
  assign new_P2_R1143_U341 = ~new_P2_R1143_U140 | ~new_P2_R1143_U340;
  assign new_P2_R1143_U342 = ~new_P2_R1143_U338 | ~new_P2_R1143_U172;
  assign new_P2_R1143_U343 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1143_U344 = ~new_P2_R1143_U141 | ~new_P2_R1143_U342;
  assign new_P2_R1143_U345 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1143_U346 = new_P2_U3416 | new_P2_U3082;
  assign new_P2_R1143_U347 = ~new_P2_R1143_U346 | ~new_P2_R1143_U40;
  assign new_P2_R1143_U348 = ~new_P2_R1143_U142 | ~new_P2_R1143_U347;
  assign new_P2_R1143_U349 = ~new_P2_R1143_U206 | ~new_P2_R1143_U171;
  assign new_P2_R1143_U350 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1143_U351 = ~new_P2_R1143_U143 | ~new_P2_R1143_U349;
  assign new_P2_R1143_U352 = ~new_P2_R1143_U207 | ~new_P2_R1143_U171;
  assign new_P2_R1143_U353 = ~new_P2_R1143_U204 | ~new_P2_R1143_U65;
  assign new_P2_R1143_U354 = ~new_P2_R1143_U214 | ~new_P2_R1143_U22;
  assign new_P2_R1143_U355 = ~new_P2_R1143_U228 | ~new_P2_R1143_U34;
  assign new_P2_R1143_U356 = ~new_P2_R1143_U231 | ~new_P2_R1143_U180;
  assign new_P2_R1143_U357 = ~new_P2_R1143_U314 | ~new_P2_R1143_U173;
  assign new_P2_R1143_U358 = ~new_P2_R1143_U298 | ~new_P2_R1143_U176;
  assign new_P2_R1143_U359 = ~new_P2_R1143_U329 | ~new_P2_R1143_U80;
  assign new_P2_R1143_U360 = ~new_P2_R1143_U282 | ~new_P2_R1143_U77;
  assign new_P2_R1143_U361 = ~new_P2_R1143_U336 | ~new_P2_R1143_U59;
  assign new_P2_R1143_U362 = ~new_P2_R1143_U345 | ~new_P2_R1143_U172;
  assign new_P2_R1143_U363 = ~new_P2_R1143_U250 | ~new_P2_R1143_U68;
  assign new_P2_R1143_U364 = ~new_P2_U3895 | ~new_P2_U3053;
  assign new_P2_R1143_U365 = ~new_P2_R1143_U296 | ~new_P2_R1143_U168;
  assign new_P2_R1143_U366 = ~new_P2_U3056 | ~new_P2_R1143_U295;
  assign new_P2_R1143_U367 = ~new_P2_U3897 | ~new_P2_R1143_U295;
  assign new_P2_R1143_U368 = ~new_P2_R1143_U301 | ~new_P2_R1143_U296 | ~new_P2_R1143_U168;
  assign new_P2_R1143_U369 = ~new_P2_R1143_U133 | ~new_P2_R1143_U155 | ~new_P2_R1143_U168;
  assign new_P2_R1143_U370 = ~new_P2_R1143_U297 | ~new_P2_R1143_U301;
  assign new_P2_R1143_U371 = ~new_P2_U3082 | ~new_P2_R1143_U39;
  assign new_P2_R1143_U372 = ~new_P2_U3416 | ~new_P2_R1143_U38;
  assign new_P2_R1143_U373 = ~new_P2_R1143_U372 | ~new_P2_R1143_U371;
  assign new_P2_R1143_U374 = ~new_P2_R1143_U352 | ~new_P2_R1143_U40;
  assign new_P2_R1143_U375 = ~new_P2_R1143_U373 | ~new_P2_R1143_U206;
  assign new_P2_R1143_U376 = ~new_P2_U3083 | ~new_P2_R1143_U36;
  assign new_P2_R1143_U377 = ~new_P2_U3413 | ~new_P2_R1143_U37;
  assign new_P2_R1143_U378 = ~new_P2_R1143_U377 | ~new_P2_R1143_U376;
  assign new_P2_R1143_U379 = ~new_P2_R1143_U353 | ~new_P2_R1143_U144;
  assign new_P2_R1143_U380 = ~new_P2_R1143_U203 | ~new_P2_R1143_U378;
  assign new_P2_R1143_U381 = ~new_P2_U3069 | ~new_P2_R1143_U23;
  assign new_P2_R1143_U382 = ~new_P2_U3410 | ~new_P2_R1143_U21;
  assign new_P2_R1143_U383 = ~new_P2_U3070 | ~new_P2_R1143_U19;
  assign new_P2_R1143_U384 = ~new_P2_U3407 | ~new_P2_R1143_U20;
  assign new_P2_R1143_U385 = ~new_P2_R1143_U384 | ~new_P2_R1143_U383;
  assign new_P2_R1143_U386 = ~new_P2_R1143_U354 | ~new_P2_R1143_U41;
  assign new_P2_R1143_U387 = ~new_P2_R1143_U385 | ~new_P2_R1143_U195;
  assign new_P2_R1143_U388 = ~new_P2_U3066 | ~new_P2_R1143_U35;
  assign new_P2_R1143_U389 = ~new_P2_U3404 | ~new_P2_R1143_U26;
  assign new_P2_R1143_U390 = ~new_P2_U3059 | ~new_P2_R1143_U24;
  assign new_P2_R1143_U391 = ~new_P2_U3401 | ~new_P2_R1143_U25;
  assign new_P2_R1143_U392 = ~new_P2_R1143_U391 | ~new_P2_R1143_U390;
  assign new_P2_R1143_U393 = ~new_P2_R1143_U355 | ~new_P2_R1143_U44;
  assign new_P2_R1143_U394 = ~new_P2_R1143_U392 | ~new_P2_R1143_U221;
  assign new_P2_R1143_U395 = ~new_P2_U3063 | ~new_P2_R1143_U32;
  assign new_P2_R1143_U396 = ~new_P2_U3398 | ~new_P2_R1143_U33;
  assign new_P2_R1143_U397 = ~new_P2_R1143_U396 | ~new_P2_R1143_U395;
  assign new_P2_R1143_U398 = ~new_P2_R1143_U356 | ~new_P2_R1143_U145;
  assign new_P2_R1143_U399 = ~new_P2_R1143_U230 | ~new_P2_R1143_U397;
  assign new_P2_R1143_U400 = ~new_P2_U3067 | ~new_P2_R1143_U27;
  assign new_P2_R1143_U401 = ~new_P2_U3395 | ~new_P2_R1143_U28;
  assign new_P2_R1143_U402 = ~new_P2_U3054 | ~new_P2_R1143_U147;
  assign new_P2_R1143_U403 = ~new_P2_U3904 | ~new_P2_R1143_U146;
  assign new_P2_R1143_U404 = ~new_P2_U3054 | ~new_P2_R1143_U147;
  assign new_P2_R1143_U405 = ~new_P2_U3904 | ~new_P2_R1143_U146;
  assign new_P2_R1143_U406 = ~new_P2_R1143_U405 | ~new_P2_R1143_U404;
  assign new_P2_R1143_U407 = ~new_P2_R1143_U148 | ~new_P2_R1143_U149;
  assign new_P2_R1143_U408 = ~new_P2_R1143_U305 | ~new_P2_R1143_U406;
  assign new_P2_R1143_U409 = ~new_P2_U3053 | ~new_P2_R1143_U88;
  assign new_P2_R1143_U410 = ~new_P2_U3895 | ~new_P2_R1143_U87;
  assign new_P2_R1143_U411 = ~new_P2_U3053 | ~new_P2_R1143_U88;
  assign new_P2_R1143_U412 = ~new_P2_U3895 | ~new_P2_R1143_U87;
  assign new_P2_R1143_U413 = ~new_P2_R1143_U412 | ~new_P2_R1143_U411;
  assign new_P2_R1143_U414 = ~new_P2_R1143_U150 | ~new_P2_R1143_U151;
  assign new_P2_R1143_U415 = ~new_P2_R1143_U303 | ~new_P2_R1143_U413;
  assign new_P2_R1143_U416 = ~new_P2_U3052 | ~new_P2_R1143_U46;
  assign new_P2_R1143_U417 = ~new_P2_U3896 | ~new_P2_R1143_U47;
  assign new_P2_R1143_U418 = ~new_P2_U3052 | ~new_P2_R1143_U46;
  assign new_P2_R1143_U419 = ~new_P2_U3896 | ~new_P2_R1143_U47;
  assign new_P2_R1143_U420 = ~new_P2_R1143_U419 | ~new_P2_R1143_U418;
  assign new_P2_R1143_U421 = ~new_P2_R1143_U152 | ~new_P2_R1143_U153;
  assign new_P2_R1143_U422 = ~new_P2_R1143_U300 | ~new_P2_R1143_U420;
  assign new_P2_R1143_U423 = ~new_P2_U3056 | ~new_P2_R1143_U49;
  assign new_P2_R1143_U424 = ~new_P2_U3897 | ~new_P2_R1143_U48;
  assign new_P2_R1143_U425 = ~new_P2_U3057 | ~new_P2_R1143_U50;
  assign new_P2_R1143_U426 = ~new_P2_U3898 | ~new_P2_R1143_U51;
  assign new_P2_R1143_U427 = ~new_P2_R1143_U426 | ~new_P2_R1143_U425;
  assign new_P2_R1143_U428 = ~new_P2_R1143_U357 | ~new_P2_R1143_U89;
  assign new_P2_R1143_U429 = ~new_P2_R1143_U427 | ~new_P2_R1143_U307;
  assign new_P2_R1143_U430 = ~new_P2_U3064 | ~new_P2_R1143_U52;
  assign new_P2_R1143_U431 = ~new_P2_U3899 | ~new_P2_R1143_U53;
  assign new_P2_R1143_U432 = ~new_P2_R1143_U431 | ~new_P2_R1143_U430;
  assign new_P2_R1143_U433 = ~new_P2_R1143_U358 | ~new_P2_R1143_U155;
  assign new_P2_R1143_U434 = ~new_P2_R1143_U294 | ~new_P2_R1143_U432;
  assign new_P2_R1143_U435 = ~new_P2_U3065 | ~new_P2_R1143_U84;
  assign new_P2_R1143_U436 = ~new_P2_U3900 | ~new_P2_R1143_U85;
  assign new_P2_R1143_U437 = ~new_P2_U3065 | ~new_P2_R1143_U84;
  assign new_P2_R1143_U438 = ~new_P2_U3900 | ~new_P2_R1143_U85;
  assign new_P2_R1143_U439 = ~new_P2_R1143_U438 | ~new_P2_R1143_U437;
  assign new_P2_R1143_U440 = ~new_P2_R1143_U156 | ~new_P2_R1143_U157;
  assign new_P2_R1143_U441 = ~new_P2_R1143_U290 | ~new_P2_R1143_U439;
  assign new_P2_R1143_U442 = ~new_P2_U3060 | ~new_P2_R1143_U82;
  assign new_P2_R1143_U443 = ~new_P2_U3901 | ~new_P2_R1143_U83;
  assign new_P2_R1143_U444 = ~new_P2_U3060 | ~new_P2_R1143_U82;
  assign new_P2_R1143_U445 = ~new_P2_U3901 | ~new_P2_R1143_U83;
  assign new_P2_R1143_U446 = ~new_P2_R1143_U445 | ~new_P2_R1143_U444;
  assign new_P2_R1143_U447 = ~new_P2_R1143_U158 | ~new_P2_R1143_U159;
  assign new_P2_R1143_U448 = ~new_P2_R1143_U286 | ~new_P2_R1143_U446;
  assign new_P2_R1143_U449 = ~new_P2_U3074 | ~new_P2_R1143_U54;
  assign new_P2_R1143_U450 = ~new_P2_U3902 | ~new_P2_R1143_U55;
  assign new_P2_R1143_U451 = ~new_P2_U3074 | ~new_P2_R1143_U54;
  assign new_P2_R1143_U452 = ~new_P2_U3902 | ~new_P2_R1143_U55;
  assign new_P2_R1143_U453 = ~new_P2_R1143_U452 | ~new_P2_R1143_U451;
  assign new_P2_R1143_U454 = ~new_P2_U3075 | ~new_P2_R1143_U81;
  assign new_P2_R1143_U455 = ~new_P2_U3903 | ~new_P2_R1143_U90;
  assign new_P2_R1143_U456 = ~new_P2_R1143_U182 | ~new_P2_R1143_U161;
  assign new_P2_R1143_U457 = ~new_P2_R1143_U328 | ~new_P2_R1143_U31;
  assign new_P2_R1143_U458 = ~new_P2_U3080 | ~new_P2_R1143_U78;
  assign new_P2_R1143_U459 = ~new_P2_U3445 | ~new_P2_R1143_U79;
  assign new_P2_R1143_U460 = ~new_P2_R1143_U459 | ~new_P2_R1143_U458;
  assign new_P2_R1143_U461 = ~new_P2_R1143_U359 | ~new_P2_R1143_U91;
  assign new_P2_R1143_U462 = ~new_P2_R1143_U460 | ~new_P2_R1143_U316;
  assign new_P2_R1143_U463 = ~new_P2_U3081 | ~new_P2_R1143_U75;
  assign new_P2_R1143_U464 = ~new_P2_U3443 | ~new_P2_R1143_U76;
  assign new_P2_R1143_U465 = ~new_P2_R1143_U464 | ~new_P2_R1143_U463;
  assign new_P2_R1143_U466 = ~new_P2_R1143_U360 | ~new_P2_R1143_U162;
  assign new_P2_R1143_U467 = ~new_P2_R1143_U270 | ~new_P2_R1143_U465;
  assign new_P2_R1143_U468 = ~new_P2_U3068 | ~new_P2_R1143_U60;
  assign new_P2_R1143_U469 = ~new_P2_U3440 | ~new_P2_R1143_U58;
  assign new_P2_R1143_U470 = ~new_P2_U3072 | ~new_P2_R1143_U56;
  assign new_P2_R1143_U471 = ~new_P2_U3437 | ~new_P2_R1143_U57;
  assign new_P2_R1143_U472 = ~new_P2_R1143_U471 | ~new_P2_R1143_U470;
  assign new_P2_R1143_U473 = ~new_P2_R1143_U361 | ~new_P2_R1143_U92;
  assign new_P2_R1143_U474 = ~new_P2_R1143_U472 | ~new_P2_R1143_U262;
  assign new_P2_R1143_U475 = ~new_P2_U3073 | ~new_P2_R1143_U73;
  assign new_P2_R1143_U476 = ~new_P2_U3434 | ~new_P2_R1143_U74;
  assign new_P2_R1143_U477 = ~new_P2_U3073 | ~new_P2_R1143_U73;
  assign new_P2_R1143_U478 = ~new_P2_U3434 | ~new_P2_R1143_U74;
  assign new_P2_R1143_U479 = ~new_P2_R1143_U478 | ~new_P2_R1143_U477;
  assign new_P2_R1143_U480 = ~new_P2_R1143_U163 | ~new_P2_R1143_U164;
  assign new_P2_R1143_U481 = ~new_P2_R1143_U258 | ~new_P2_R1143_U479;
  assign new_P2_R1143_U482 = ~new_P2_U3078 | ~new_P2_R1143_U71;
  assign new_P2_R1143_U483 = ~new_P2_U3431 | ~new_P2_R1143_U72;
  assign new_P2_R1143_U484 = ~new_P2_U3078 | ~new_P2_R1143_U71;
  assign new_P2_R1143_U485 = ~new_P2_U3431 | ~new_P2_R1143_U72;
  assign new_P2_R1143_U486 = ~new_P2_R1143_U485 | ~new_P2_R1143_U484;
  assign new_P2_R1143_U487 = ~new_P2_R1143_U165 | ~new_P2_R1143_U166;
  assign new_P2_R1143_U488 = ~new_P2_R1143_U254 | ~new_P2_R1143_U486;
  assign new_P2_R1143_U489 = ~new_P2_U3079 | ~new_P2_R1143_U61;
  assign new_P2_R1143_U490 = ~new_P2_U3428 | ~new_P2_R1143_U62;
  assign new_P2_R1143_U491 = ~new_P2_U3071 | ~new_P2_R1143_U69;
  assign new_P2_R1143_U492 = ~new_P2_U3425 | ~new_P2_R1143_U70;
  assign new_P2_R1143_U493 = ~new_P2_R1143_U492 | ~new_P2_R1143_U491;
  assign new_P2_R1143_U494 = ~new_P2_R1143_U362 | ~new_P2_R1143_U93;
  assign new_P2_R1143_U495 = ~new_P2_R1143_U493 | ~new_P2_R1143_U338;
  assign new_P2_R1143_U496 = ~new_P2_U3062 | ~new_P2_R1143_U66;
  assign new_P2_R1143_U497 = ~new_P2_U3422 | ~new_P2_R1143_U67;
  assign new_P2_R1143_U498 = ~new_P2_R1143_U497 | ~new_P2_R1143_U496;
  assign new_P2_R1143_U499 = ~new_P2_R1143_U363 | ~new_P2_R1143_U167;
  assign new_P2_R1143_U500 = ~new_P2_R1143_U244 | ~new_P2_R1143_U498;
  assign new_P2_R1143_U501 = ~new_P2_U3061 | ~new_P2_R1143_U63;
  assign new_P2_R1143_U502 = ~new_P2_U3419 | ~new_P2_R1143_U64;
  assign new_P2_R1143_U503 = ~new_P2_U3076 | ~new_P2_R1143_U29;
  assign new_P2_R1143_U504 = ~new_P2_U3387 | ~new_P2_R1143_U30;
  assign new_P2_R1158_U4 = new_P2_R1158_U227 & new_P2_R1158_U226;
  assign new_P2_R1158_U5 = new_P2_R1158_U238 & new_P2_R1158_U237;
  assign new_P2_R1158_U6 = new_P2_R1158_U264 & new_P2_R1158_U263;
  assign new_P2_R1158_U7 = new_P2_R1158_U276 & new_P2_R1158_U275;
  assign new_P2_R1158_U8 = new_P2_R1158_U288 & new_P2_R1158_U287;
  assign new_P2_R1158_U9 = new_P2_R1158_U6 & new_P2_R1158_U268;
  assign new_P2_R1158_U10 = new_P2_R1158_U5 & new_P2_R1158_U235;
  assign new_P2_R1158_U11 = new_P2_R1158_U9 & new_P2_R1158_U261;
  assign new_P2_R1158_U12 = new_P2_R1158_U11 & new_P2_R1158_U271;
  assign new_P2_R1158_U13 = new_P2_R1158_U537 & new_P2_R1158_U536;
  assign new_P2_R1158_U14 = new_P2_R1158_U343 & new_P2_R1158_U340;
  assign new_P2_R1158_U15 = new_P2_R1158_U334 & new_P2_R1158_U331;
  assign new_P2_R1158_U16 = new_P2_R1158_U327 & new_P2_R1158_U324;
  assign new_P2_R1158_U17 = new_P2_R1158_U538 & new_P2_R1158_U539 & new_P2_R1158_U142 & new_P2_R1158_U394;
  assign new_P2_R1158_U18 = new_P2_R1158_U257 & new_P2_R1158_U254;
  assign new_P2_R1158_U19 = new_P2_R1158_U250 & new_P2_R1158_U247;
  assign new_P2_R1158_U20 = ~new_P2_U3056 | ~new_P2_R1158_U305;
  assign new_P2_R1158_U21 = ~new_P2_U3152;
  assign new_P2_R1158_U22 = ~new_P2_U3083;
  assign new_P2_R1158_U23 = ~new_P2_U3070;
  assign new_P2_R1158_U24 = ~new_P2_U3070 | ~new_P2_R1158_U69;
  assign new_P2_R1158_U25 = ~new_P2_U3069;
  assign new_P2_R1158_U26 = ~new_P2_U3066;
  assign new_P2_R1158_U27 = ~new_P2_U3066 | ~new_P2_R1158_U71;
  assign new_P2_R1158_U28 = ~new_P2_U3067;
  assign new_P2_R1158_U29 = ~new_P2_U3067 | ~new_P2_R1158_U72;
  assign new_P2_R1158_U30 = ~new_P2_U3063;
  assign new_P2_R1158_U31 = ~new_P2_U3077;
  assign new_P2_R1158_U32 = ~new_P2_U3076;
  assign new_P2_R1158_U33 = ~new_P2_U3059;
  assign new_P2_R1158_U34 = ~new_P2_U3082;
  assign new_P2_R1158_U35 = ~new_P2_R1158_U359 | ~new_P2_R1158_U242 | ~new_P2_R1158_U241;
  assign new_P2_R1158_U36 = ~new_P2_R1158_U386 | ~new_P2_R1158_U27;
  assign new_P2_R1158_U37 = ~new_P2_R1158_U357 | ~new_P2_R1158_U358 | ~new_P2_R1158_U224;
  assign new_P2_R1158_U38 = ~new_P2_U3052;
  assign new_P2_R1158_U39 = ~new_P2_U3057;
  assign new_P2_R1158_U40 = ~new_P2_U3064;
  assign new_P2_R1158_U41 = ~new_P2_U3056;
  assign new_P2_R1158_U42 = ~new_P2_U3072;
  assign new_P2_R1158_U43 = ~new_P2_U3072 | ~new_P2_R1158_U81;
  assign new_P2_R1158_U44 = ~new_P2_U3068;
  assign new_P2_R1158_U45 = ~new_P2_U3073;
  assign new_P2_R1158_U46 = ~new_P2_U3078;
  assign new_P2_R1158_U47 = ~new_P2_U3071;
  assign new_P2_R1158_U48 = ~new_P2_U3062;
  assign new_P2_R1158_U49 = ~new_P2_U3062 | ~new_P2_R1158_U87;
  assign new_P2_R1158_U50 = ~new_P2_U3079;
  assign new_P2_R1158_U51 = ~new_P2_U3061;
  assign new_P2_R1158_U52 = ~new_P2_U3061 | ~new_P2_R1158_U88;
  assign new_P2_R1158_U53 = ~new_P2_U3081;
  assign new_P2_R1158_U54 = ~new_P2_U3075;
  assign new_P2_R1158_U55 = ~new_P2_U3080;
  assign new_P2_R1158_U56 = ~new_P2_U3080 | ~new_P2_R1158_U90;
  assign new_P2_R1158_U57 = ~new_P2_U3074;
  assign new_P2_R1158_U58 = ~new_P2_U3060;
  assign new_P2_R1158_U59 = ~new_P2_U3065;
  assign new_P2_R1158_U60 = ~new_P2_U3057 | ~new_P2_R1158_U78;
  assign new_P2_R1158_U61 = ~new_P2_R1158_U308 | ~new_P2_R1158_U192;
  assign new_P2_R1158_U62 = ~new_P2_R1158_U56 | ~new_P2_R1158_U320;
  assign new_P2_R1158_U63 = ~new_P2_R1158_U129 | ~new_P2_R1158_U384;
  assign new_P2_R1158_U64 = ~new_P2_R1158_U364 | ~new_P2_R1158_U272;
  assign new_P2_R1158_U65 = ~new_P2_R1158_U362 | ~new_P2_R1158_U270;
  assign new_P2_R1158_U66 = ~new_P2_R1158_U49 | ~new_P2_R1158_U336;
  assign new_P2_R1158_U67 = ~new_P2_R1158_U396 | ~new_P2_R1158_U395;
  assign new_P2_R1158_U68 = ~new_P2_R1158_U428 | ~new_P2_R1158_U427;
  assign new_P2_R1158_U69 = ~new_P2_R1158_U425 | ~new_P2_R1158_U424;
  assign new_P2_R1158_U70 = ~new_P2_R1158_U422 | ~new_P2_R1158_U421;
  assign new_P2_R1158_U71 = ~new_P2_R1158_U419 | ~new_P2_R1158_U418;
  assign new_P2_R1158_U72 = ~new_P2_R1158_U416 | ~new_P2_R1158_U415;
  assign new_P2_R1158_U73 = ~new_P2_R1158_U413 | ~new_P2_R1158_U412;
  assign new_P2_R1158_U74 = ~new_P2_R1158_U407 | ~new_P2_R1158_U406;
  assign new_P2_R1158_U75 = ~new_P2_R1158_U410 | ~new_P2_R1158_U409;
  assign new_P2_R1158_U76 = ~new_P2_R1158_U404 | ~new_P2_R1158_U403;
  assign new_P2_R1158_U77 = ~new_P2_R1158_U468 | ~new_P2_R1158_U467;
  assign new_P2_R1158_U78 = ~new_P2_R1158_U516 | ~new_P2_R1158_U515;
  assign new_P2_R1158_U79 = ~new_P2_R1158_U519 | ~new_P2_R1158_U518;
  assign new_P2_R1158_U80 = ~new_P2_R1158_U513 | ~new_P2_R1158_U512;
  assign new_P2_R1158_U81 = ~new_P2_R1158_U492 | ~new_P2_R1158_U491;
  assign new_P2_R1158_U82 = ~new_P2_R1158_U489 | ~new_P2_R1158_U488;
  assign new_P2_R1158_U83 = ~new_P2_R1158_U486 | ~new_P2_R1158_U485;
  assign new_P2_R1158_U84 = ~new_P2_R1158_U471 | ~new_P2_R1158_U470;
  assign new_P2_R1158_U85 = ~new_P2_R1158_U483 | ~new_P2_R1158_U482;
  assign new_P2_R1158_U86 = ~new_P2_R1158_U480 | ~new_P2_R1158_U479;
  assign new_P2_R1158_U87 = ~new_P2_R1158_U477 | ~new_P2_R1158_U476;
  assign new_P2_R1158_U88 = ~new_P2_R1158_U474 | ~new_P2_R1158_U473;
  assign new_P2_R1158_U89 = ~new_P2_R1158_U495 | ~new_P2_R1158_U494;
  assign new_P2_R1158_U90 = ~new_P2_R1158_U504 | ~new_P2_R1158_U503;
  assign new_P2_R1158_U91 = ~new_P2_R1158_U498 | ~new_P2_R1158_U497;
  assign new_P2_R1158_U92 = ~new_P2_R1158_U501 | ~new_P2_R1158_U500;
  assign new_P2_R1158_U93 = ~new_P2_R1158_U507 | ~new_P2_R1158_U506;
  assign new_P2_R1158_U94 = ~new_P2_R1158_U510 | ~new_P2_R1158_U509;
  assign new_P2_R1158_U95 = ~new_P2_R1158_U525 | ~new_P2_R1158_U524;
  assign new_P2_R1158_U96 = ~new_P2_R1158_U634 | ~new_P2_R1158_U633;
  assign new_P2_R1158_U97 = ~new_P2_R1158_U431 | ~new_P2_R1158_U430;
  assign new_P2_R1158_U98 = ~new_P2_R1158_U438 | ~new_P2_R1158_U437;
  assign new_P2_R1158_U99 = ~new_P2_R1158_U445 | ~new_P2_R1158_U444;
  assign new_P2_R1158_U100 = ~new_P2_R1158_U452 | ~new_P2_R1158_U451;
  assign new_P2_R1158_U101 = ~new_P2_R1158_U459 | ~new_P2_R1158_U458;
  assign new_P2_R1158_U102 = ~new_P2_R1158_U466 | ~new_P2_R1158_U465;
  assign new_P2_R1158_U103 = ~new_P2_R1158_U528 | ~new_P2_R1158_U527;
  assign new_P2_R1158_U104 = ~new_P2_R1158_U535 | ~new_P2_R1158_U534;
  assign new_P2_R1158_U105 = ~new_P2_R1158_U544 | ~new_P2_R1158_U543;
  assign new_P2_R1158_U106 = ~new_P2_R1158_U549 | ~new_P2_R1158_U548;
  assign new_P2_R1158_U107 = ~new_P2_R1158_U556 | ~new_P2_R1158_U555;
  assign new_P2_R1158_U108 = ~new_P2_R1158_U563 | ~new_P2_R1158_U562;
  assign new_P2_R1158_U109 = ~new_P2_R1158_U570 | ~new_P2_R1158_U569;
  assign new_P2_R1158_U110 = ~new_P2_R1158_U577 | ~new_P2_R1158_U576;
  assign new_P2_R1158_U111 = ~new_P2_R1158_U582 | ~new_P2_R1158_U581;
  assign new_P2_R1158_U112 = ~new_P2_R1158_U589 | ~new_P2_R1158_U588;
  assign new_P2_R1158_U113 = ~new_P2_R1158_U596 | ~new_P2_R1158_U595;
  assign new_P2_R1158_U114 = ~new_P2_R1158_U603 | ~new_P2_R1158_U602;
  assign new_P2_R1158_U115 = ~new_P2_R1158_U610 | ~new_P2_R1158_U609;
  assign new_P2_R1158_U116 = ~new_P2_R1158_U617 | ~new_P2_R1158_U616;
  assign new_P2_R1158_U117 = ~new_P2_R1158_U622 | ~new_P2_R1158_U621;
  assign new_P2_R1158_U118 = ~new_P2_R1158_U629 | ~new_P2_R1158_U628;
  assign new_P2_R1158_U119 = new_P2_R1158_U75 & new_P2_U3152;
  assign new_P2_R1158_U120 = new_P2_R1158_U230 & new_P2_R1158_U229;
  assign new_P2_R1158_U121 = new_P2_R1158_U243 & new_P2_R1158_U10;
  assign new_P2_R1158_U122 = new_P2_R1158_U361 & new_P2_R1158_U244;
  assign new_P2_R1158_U123 = new_P2_R1158_U24 & new_P2_R1158_U440 & new_P2_R1158_U439;
  assign new_P2_R1158_U124 = new_P2_R1158_U249 & new_P2_R1158_U5;
  assign new_P2_R1158_U125 = new_P2_R1158_U29 & new_P2_R1158_U461 & new_P2_R1158_U460;
  assign new_P2_R1158_U126 = new_P2_R1158_U256 & new_P2_R1158_U4;
  assign new_P2_R1158_U127 = new_P2_R1158_U266 & new_P2_R1158_U213;
  assign new_P2_R1158_U128 = new_P2_R1158_U273 & new_P2_R1158_U12;
  assign new_P2_R1158_U129 = new_P2_R1158_U372 & new_P2_R1158_U274;
  assign new_P2_R1158_U130 = new_P2_R1158_U280 & new_P2_R1158_U279;
  assign new_P2_R1158_U131 = new_P2_R1158_U292 & new_P2_R1158_U8;
  assign new_P2_R1158_U132 = new_P2_R1158_U290 & new_P2_R1158_U214;
  assign new_P2_R1158_U133 = new_P2_R1158_U313 & new_P2_R1158_U375;
  assign new_P2_R1158_U134 = new_P2_R1158_U315 & new_P2_R1158_U306;
  assign new_P2_R1158_U135 = new_P2_R1158_U315 & new_P2_R1158_U369;
  assign new_P2_R1158_U136 = new_P2_R1158_U373 & new_P2_R1158_U314;
  assign new_P2_R1158_U137 = ~new_P2_R1158_U522 | ~new_P2_R1158_U521;
  assign new_P2_R1158_U138 = new_P2_R1158_U318 & new_P2_R1158_U215;
  assign new_P2_R1158_U139 = new_P2_R1158_U517 & new_P2_R1158_U39;
  assign new_P2_R1158_U140 = new_P2_R1158_U318 & new_P2_R1158_U209;
  assign new_P2_R1158_U141 = new_P2_R1158_U13 & new_P2_R1158_U60;
  assign new_P2_R1158_U142 = new_P2_R1158_U393 & new_P2_R1158_U392;
  assign new_P2_R1158_U143 = new_P2_R1158_U214 & new_P2_R1158_U565 & new_P2_R1158_U564;
  assign new_P2_R1158_U144 = new_P2_R1158_U326 & new_P2_R1158_U8;
  assign new_P2_R1158_U145 = new_P2_R1158_U43 & new_P2_R1158_U591 & new_P2_R1158_U590;
  assign new_P2_R1158_U146 = new_P2_R1158_U333 & new_P2_R1158_U7;
  assign new_P2_R1158_U147 = new_P2_R1158_U213 & new_P2_R1158_U612 & new_P2_R1158_U611;
  assign new_P2_R1158_U148 = new_P2_R1158_U342 & new_P2_R1158_U6;
  assign new_P2_R1158_U149 = ~new_P2_R1158_U631 | ~new_P2_R1158_U630;
  assign new_P2_R1158_U150 = ~new_P2_U3416;
  assign new_P2_R1158_U151 = new_P2_R1158_U399 & new_P2_R1158_U398;
  assign new_P2_R1158_U152 = ~new_P2_U3401;
  assign new_P2_R1158_U153 = ~new_P2_U3392;
  assign new_P2_R1158_U154 = ~new_P2_U3387;
  assign new_P2_R1158_U155 = ~new_P2_U3398;
  assign new_P2_R1158_U156 = ~new_P2_U3395;
  assign new_P2_R1158_U157 = ~new_P2_U3404;
  assign new_P2_R1158_U158 = ~new_P2_U3410;
  assign new_P2_R1158_U159 = ~new_P2_U3407;
  assign new_P2_R1158_U160 = ~new_P2_U3413;
  assign new_P2_R1158_U161 = ~new_P2_R1158_U122 | ~new_P2_R1158_U390;
  assign new_P2_R1158_U162 = new_P2_R1158_U433 & new_P2_R1158_U432;
  assign new_P2_R1158_U163 = ~new_P2_R1158_U360 | ~new_P2_R1158_U388;
  assign new_P2_R1158_U164 = new_P2_R1158_U447 & new_P2_R1158_U446;
  assign new_P2_R1158_U165 = ~new_P2_R1158_U354 | ~new_P2_R1158_U233 | ~new_P2_R1158_U211;
  assign new_P2_R1158_U166 = new_P2_R1158_U454 & new_P2_R1158_U453;
  assign new_P2_R1158_U167 = ~new_P2_R1158_U120 | ~new_P2_R1158_U231;
  assign new_P2_R1158_U168 = ~new_P2_U3896;
  assign new_P2_R1158_U169 = ~new_P2_U3431;
  assign new_P2_R1158_U170 = ~new_P2_U3419;
  assign new_P2_R1158_U171 = ~new_P2_U3422;
  assign new_P2_R1158_U172 = ~new_P2_U3428;
  assign new_P2_R1158_U173 = ~new_P2_U3425;
  assign new_P2_R1158_U174 = ~new_P2_U3434;
  assign new_P2_R1158_U175 = ~new_P2_U3440;
  assign new_P2_R1158_U176 = ~new_P2_U3437;
  assign new_P2_R1158_U177 = ~new_P2_U3443;
  assign new_P2_R1158_U178 = ~new_P2_U3902;
  assign new_P2_R1158_U179 = ~new_P2_U3903;
  assign new_P2_R1158_U180 = ~new_P2_U3445;
  assign new_P2_R1158_U181 = ~new_P2_U3901;
  assign new_P2_R1158_U182 = ~new_P2_U3900;
  assign new_P2_R1158_U183 = ~new_P2_U3897;
  assign new_P2_R1158_U184 = ~new_P2_U3898;
  assign new_P2_R1158_U185 = ~new_P2_U3899;
  assign new_P2_R1158_U186 = ~new_P2_U3053;
  assign new_P2_R1158_U187 = ~new_P2_U3895;
  assign new_P2_R1158_U188 = new_P2_R1158_U530 & new_P2_R1158_U529;
  assign new_P2_R1158_U189 = ~new_P2_R1158_U310 | ~new_P2_R1158_U309;
  assign new_P2_R1158_U190 = ~new_P2_U3064 | ~new_P2_R1158_U79;
  assign new_P2_R1158_U191 = ~new_P2_R1158_U190 | ~new_P2_R1158_U61;
  assign new_P2_R1158_U192 = ~new_P2_R1158_U303 | ~new_P2_R1158_U302;
  assign new_P2_R1158_U193 = new_P2_R1158_U551 & new_P2_R1158_U550;
  assign new_P2_R1158_U194 = ~new_P2_R1158_U299 | ~new_P2_R1158_U298;
  assign new_P2_R1158_U195 = new_P2_R1158_U558 & new_P2_R1158_U557;
  assign new_P2_R1158_U196 = ~new_P2_R1158_U295 | ~new_P2_R1158_U294;
  assign new_P2_R1158_U197 = new_P2_R1158_U572 & new_P2_R1158_U571;
  assign new_P2_R1158_U198 = ~new_P2_R1158_U221 | ~new_P2_R1158_U220;
  assign new_P2_R1158_U199 = ~new_P2_R1158_U285 | ~new_P2_R1158_U284;
  assign new_P2_R1158_U200 = new_P2_R1158_U584 & new_P2_R1158_U583;
  assign new_P2_R1158_U201 = ~new_P2_R1158_U130 | ~new_P2_R1158_U281;
  assign new_P2_R1158_U202 = new_P2_R1158_U598 & new_P2_R1158_U597;
  assign new_P2_R1158_U203 = ~new_P2_R1158_U368 | ~new_P2_R1158_U382;
  assign new_P2_R1158_U204 = new_P2_R1158_U605 & new_P2_R1158_U604;
  assign new_P2_R1158_U205 = ~new_P2_R1158_U363 | ~new_P2_R1158_U380;
  assign new_P2_R1158_U206 = ~new_P2_R1158_U378 | ~new_P2_R1158_U52;
  assign new_P2_R1158_U207 = new_P2_R1158_U624 & new_P2_R1158_U623;
  assign new_P2_R1158_U208 = ~new_P2_R1158_U355 | ~new_P2_R1158_U259 | ~new_P2_R1158_U210;
  assign new_P2_R1158_U209 = ~new_P2_R1158_U20 | ~new_P2_R1158_U366;
  assign new_P2_R1158_U210 = ~new_P2_R1158_U67 | ~new_P2_R1158_U161;
  assign new_P2_R1158_U211 = ~new_P2_R1158_U76 | ~new_P2_R1158_U167;
  assign new_P2_R1158_U212 = ~new_P2_R1158_U29;
  assign new_P2_R1158_U213 = ~new_P2_U3071 | ~new_P2_R1158_U85;
  assign new_P2_R1158_U214 = ~new_P2_U3075 | ~new_P2_R1158_U92;
  assign new_P2_R1158_U215 = ~new_P2_R1158_U60;
  assign new_P2_R1158_U216 = ~new_P2_R1158_U49;
  assign new_P2_R1158_U217 = ~new_P2_R1158_U56;
  assign new_P2_R1158_U218 = ~new_P2_R1158_U190;
  assign new_P2_R1158_U219 = ~new_P2_R1158_U411 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U220 = ~new_P2_U3076 | ~new_P2_R1158_U219;
  assign new_P2_R1158_U221 = ~new_P2_U3152 | ~new_P2_R1158_U75;
  assign new_P2_R1158_U222 = ~new_P2_R1158_U198;
  assign new_P2_R1158_U223 = ~new_P2_R1158_U408 | ~new_P2_R1158_U31;
  assign new_P2_R1158_U224 = ~new_P2_U3077 | ~new_P2_R1158_U74;
  assign new_P2_R1158_U225 = ~new_P2_R1158_U37;
  assign new_P2_R1158_U226 = ~new_P2_R1158_U414 | ~new_P2_R1158_U30;
  assign new_P2_R1158_U227 = ~new_P2_R1158_U417 | ~new_P2_R1158_U28;
  assign new_P2_R1158_U228 = ~new_P2_R1158_U30 | ~new_P2_R1158_U29;
  assign new_P2_R1158_U229 = ~new_P2_R1158_U73 | ~new_P2_R1158_U228;
  assign new_P2_R1158_U230 = ~new_P2_U3063 | ~new_P2_R1158_U212;
  assign new_P2_R1158_U231 = ~new_P2_R1158_U4 | ~new_P2_R1158_U37;
  assign new_P2_R1158_U232 = ~new_P2_R1158_U167;
  assign new_P2_R1158_U233 = ~new_P2_U3059 | ~new_P2_R1158_U167;
  assign new_P2_R1158_U234 = ~new_P2_R1158_U165;
  assign new_P2_R1158_U235 = ~new_P2_R1158_U420 | ~new_P2_R1158_U26;
  assign new_P2_R1158_U236 = ~new_P2_R1158_U27;
  assign new_P2_R1158_U237 = ~new_P2_R1158_U423 | ~new_P2_R1158_U25;
  assign new_P2_R1158_U238 = ~new_P2_R1158_U426 | ~new_P2_R1158_U23;
  assign new_P2_R1158_U239 = ~new_P2_R1158_U24;
  assign new_P2_R1158_U240 = ~new_P2_R1158_U25 | ~new_P2_R1158_U24;
  assign new_P2_R1158_U241 = ~new_P2_R1158_U70 | ~new_P2_R1158_U240;
  assign new_P2_R1158_U242 = ~new_P2_U3069 | ~new_P2_R1158_U239;
  assign new_P2_R1158_U243 = ~new_P2_R1158_U429 | ~new_P2_R1158_U22;
  assign new_P2_R1158_U244 = ~new_P2_U3083 | ~new_P2_R1158_U68;
  assign new_P2_R1158_U245 = ~new_P2_R1158_U426 | ~new_P2_R1158_U23;
  assign new_P2_R1158_U246 = ~new_P2_R1158_U245 | ~new_P2_R1158_U36;
  assign new_P2_R1158_U247 = ~new_P2_R1158_U123 | ~new_P2_R1158_U246;
  assign new_P2_R1158_U248 = ~new_P2_R1158_U387 | ~new_P2_R1158_U24;
  assign new_P2_R1158_U249 = ~new_P2_U3069 | ~new_P2_R1158_U70;
  assign new_P2_R1158_U250 = ~new_P2_R1158_U124 | ~new_P2_R1158_U248;
  assign new_P2_R1158_U251 = ~new_P2_R1158_U426 | ~new_P2_R1158_U23;
  assign new_P2_R1158_U252 = ~new_P2_R1158_U417 | ~new_P2_R1158_U28;
  assign new_P2_R1158_U253 = ~new_P2_R1158_U252 | ~new_P2_R1158_U37;
  assign new_P2_R1158_U254 = ~new_P2_R1158_U125 | ~new_P2_R1158_U253;
  assign new_P2_R1158_U255 = ~new_P2_R1158_U225 | ~new_P2_R1158_U29;
  assign new_P2_R1158_U256 = ~new_P2_U3063 | ~new_P2_R1158_U73;
  assign new_P2_R1158_U257 = ~new_P2_R1158_U126 | ~new_P2_R1158_U255;
  assign new_P2_R1158_U258 = ~new_P2_R1158_U417 | ~new_P2_R1158_U28;
  assign new_P2_R1158_U259 = ~new_P2_U3082 | ~new_P2_R1158_U161;
  assign new_P2_R1158_U260 = ~new_P2_R1158_U208;
  assign new_P2_R1158_U261 = ~new_P2_R1158_U475 | ~new_P2_R1158_U51;
  assign new_P2_R1158_U262 = ~new_P2_R1158_U52;
  assign new_P2_R1158_U263 = ~new_P2_R1158_U481 | ~new_P2_R1158_U50;
  assign new_P2_R1158_U264 = ~new_P2_R1158_U484 | ~new_P2_R1158_U47;
  assign new_P2_R1158_U265 = ~new_P2_R1158_U216 | ~new_P2_R1158_U6;
  assign new_P2_R1158_U266 = ~new_P2_U3079 | ~new_P2_R1158_U86;
  assign new_P2_R1158_U267 = ~new_P2_R1158_U127 | ~new_P2_R1158_U265;
  assign new_P2_R1158_U268 = ~new_P2_R1158_U478 | ~new_P2_R1158_U48;
  assign new_P2_R1158_U269 = ~new_P2_R1158_U481 | ~new_P2_R1158_U50;
  assign new_P2_R1158_U270 = ~new_P2_R1158_U269 | ~new_P2_R1158_U267;
  assign new_P2_R1158_U271 = ~new_P2_R1158_U472 | ~new_P2_R1158_U46;
  assign new_P2_R1158_U272 = ~new_P2_U3078 | ~new_P2_R1158_U84;
  assign new_P2_R1158_U273 = ~new_P2_R1158_U487 | ~new_P2_R1158_U45;
  assign new_P2_R1158_U274 = ~new_P2_U3073 | ~new_P2_R1158_U83;
  assign new_P2_R1158_U275 = ~new_P2_R1158_U490 | ~new_P2_R1158_U44;
  assign new_P2_R1158_U276 = ~new_P2_R1158_U493 | ~new_P2_R1158_U42;
  assign new_P2_R1158_U277 = ~new_P2_R1158_U43;
  assign new_P2_R1158_U278 = ~new_P2_R1158_U44 | ~new_P2_R1158_U43;
  assign new_P2_R1158_U279 = ~new_P2_R1158_U82 | ~new_P2_R1158_U278;
  assign new_P2_R1158_U280 = ~new_P2_U3068 | ~new_P2_R1158_U277;
  assign new_P2_R1158_U281 = ~new_P2_R1158_U7 | ~new_P2_R1158_U63;
  assign new_P2_R1158_U282 = ~new_P2_R1158_U201;
  assign new_P2_R1158_U283 = ~new_P2_R1158_U496 | ~new_P2_R1158_U53;
  assign new_P2_R1158_U284 = ~new_P2_R1158_U283 | ~new_P2_R1158_U201;
  assign new_P2_R1158_U285 = ~new_P2_U3081 | ~new_P2_R1158_U89;
  assign new_P2_R1158_U286 = ~new_P2_R1158_U199;
  assign new_P2_R1158_U287 = ~new_P2_R1158_U499 | ~new_P2_R1158_U57;
  assign new_P2_R1158_U288 = ~new_P2_R1158_U502 | ~new_P2_R1158_U54;
  assign new_P2_R1158_U289 = ~new_P2_R1158_U217 | ~new_P2_R1158_U8;
  assign new_P2_R1158_U290 = ~new_P2_U3074 | ~new_P2_R1158_U91;
  assign new_P2_R1158_U291 = ~new_P2_R1158_U132 | ~new_P2_R1158_U289;
  assign new_P2_R1158_U292 = ~new_P2_R1158_U505 | ~new_P2_R1158_U55;
  assign new_P2_R1158_U293 = ~new_P2_R1158_U499 | ~new_P2_R1158_U57;
  assign new_P2_R1158_U294 = ~new_P2_R1158_U131 | ~new_P2_R1158_U199;
  assign new_P2_R1158_U295 = ~new_P2_R1158_U293 | ~new_P2_R1158_U291;
  assign new_P2_R1158_U296 = ~new_P2_R1158_U196;
  assign new_P2_R1158_U297 = ~new_P2_R1158_U508 | ~new_P2_R1158_U58;
  assign new_P2_R1158_U298 = ~new_P2_R1158_U297 | ~new_P2_R1158_U196;
  assign new_P2_R1158_U299 = ~new_P2_U3060 | ~new_P2_R1158_U93;
  assign new_P2_R1158_U300 = ~new_P2_R1158_U194;
  assign new_P2_R1158_U301 = ~new_P2_R1158_U511 | ~new_P2_R1158_U59;
  assign new_P2_R1158_U302 = ~new_P2_R1158_U301 | ~new_P2_R1158_U194;
  assign new_P2_R1158_U303 = ~new_P2_U3065 | ~new_P2_R1158_U94;
  assign new_P2_R1158_U304 = ~new_P2_R1158_U192;
  assign new_P2_R1158_U305 = ~new_P2_R1158_U517 | ~new_P2_R1158_U39;
  assign new_P2_R1158_U306 = ~new_P2_R1158_U307 | ~new_P2_R1158_U190 | ~new_P2_R1158_U60;
  assign new_P2_R1158_U307 = ~new_P2_U3056 | ~new_P2_R1158_U80;
  assign new_P2_R1158_U308 = ~new_P2_R1158_U520 | ~new_P2_R1158_U40;
  assign new_P2_R1158_U309 = ~new_P2_R1158_U369 | ~new_P2_R1158_U192;
  assign new_P2_R1158_U310 = ~new_P2_R1158_U365 | ~new_P2_R1158_U306;
  assign new_P2_R1158_U311 = ~new_P2_R1158_U189;
  assign new_P2_R1158_U312 = ~new_P2_R1158_U469 | ~new_P2_R1158_U38;
  assign new_P2_R1158_U313 = ~new_P2_U3052 | ~new_P2_R1158_U77;
  assign new_P2_R1158_U314 = ~new_P2_U3052 | ~new_P2_R1158_U77;
  assign new_P2_R1158_U315 = ~new_P2_R1158_U469 | ~new_P2_R1158_U38;
  assign new_P2_R1158_U316 = ~new_P2_R1158_U61;
  assign new_P2_R1158_U317 = ~new_P2_R1158_U191;
  assign new_P2_R1158_U318 = ~new_P2_U3056 | ~new_P2_R1158_U80;
  assign new_P2_R1158_U319 = ~new_P2_R1158_U517 | ~new_P2_R1158_U39;
  assign new_P2_R1158_U320 = ~new_P2_R1158_U292 | ~new_P2_R1158_U199;
  assign new_P2_R1158_U321 = ~new_P2_R1158_U62;
  assign new_P2_R1158_U322 = ~new_P2_R1158_U502 | ~new_P2_R1158_U54;
  assign new_P2_R1158_U323 = ~new_P2_R1158_U322 | ~new_P2_R1158_U62;
  assign new_P2_R1158_U324 = ~new_P2_R1158_U143 | ~new_P2_R1158_U323;
  assign new_P2_R1158_U325 = ~new_P2_R1158_U321 | ~new_P2_R1158_U214;
  assign new_P2_R1158_U326 = ~new_P2_U3074 | ~new_P2_R1158_U91;
  assign new_P2_R1158_U327 = ~new_P2_R1158_U144 | ~new_P2_R1158_U325;
  assign new_P2_R1158_U328 = ~new_P2_R1158_U502 | ~new_P2_R1158_U54;
  assign new_P2_R1158_U329 = ~new_P2_R1158_U493 | ~new_P2_R1158_U42;
  assign new_P2_R1158_U330 = ~new_P2_R1158_U329 | ~new_P2_R1158_U63;
  assign new_P2_R1158_U331 = ~new_P2_R1158_U145 | ~new_P2_R1158_U330;
  assign new_P2_R1158_U332 = ~new_P2_R1158_U385 | ~new_P2_R1158_U43;
  assign new_P2_R1158_U333 = ~new_P2_U3068 | ~new_P2_R1158_U82;
  assign new_P2_R1158_U334 = ~new_P2_R1158_U146 | ~new_P2_R1158_U332;
  assign new_P2_R1158_U335 = ~new_P2_R1158_U493 | ~new_P2_R1158_U42;
  assign new_P2_R1158_U336 = ~new_P2_R1158_U268 | ~new_P2_R1158_U206;
  assign new_P2_R1158_U337 = ~new_P2_R1158_U66;
  assign new_P2_R1158_U338 = ~new_P2_R1158_U484 | ~new_P2_R1158_U47;
  assign new_P2_R1158_U339 = ~new_P2_R1158_U338 | ~new_P2_R1158_U66;
  assign new_P2_R1158_U340 = ~new_P2_R1158_U147 | ~new_P2_R1158_U339;
  assign new_P2_R1158_U341 = ~new_P2_R1158_U337 | ~new_P2_R1158_U213;
  assign new_P2_R1158_U342 = ~new_P2_U3079 | ~new_P2_R1158_U86;
  assign new_P2_R1158_U343 = ~new_P2_R1158_U148 | ~new_P2_R1158_U341;
  assign new_P2_R1158_U344 = ~new_P2_R1158_U484 | ~new_P2_R1158_U47;
  assign new_P2_R1158_U345 = ~new_P2_R1158_U251 | ~new_P2_R1158_U24;
  assign new_P2_R1158_U346 = ~new_P2_R1158_U258 | ~new_P2_R1158_U29;
  assign new_P2_R1158_U347 = ~new_P2_R1158_U319 | ~new_P2_R1158_U60;
  assign new_P2_R1158_U348 = ~new_P2_R1158_U308 | ~new_P2_R1158_U190;
  assign new_P2_R1158_U349 = ~new_P2_R1158_U328 | ~new_P2_R1158_U214;
  assign new_P2_R1158_U350 = ~new_P2_R1158_U292 | ~new_P2_R1158_U56;
  assign new_P2_R1158_U351 = ~new_P2_R1158_U335 | ~new_P2_R1158_U43;
  assign new_P2_R1158_U352 = ~new_P2_R1158_U344 | ~new_P2_R1158_U213;
  assign new_P2_R1158_U353 = ~new_P2_R1158_U268 | ~new_P2_R1158_U49;
  assign new_P2_R1158_U354 = ~new_P2_U3059 | ~new_P2_R1158_U76;
  assign new_P2_R1158_U355 = ~new_P2_U3082 | ~new_P2_R1158_U67;
  assign new_P2_R1158_U356 = ~new_P2_R1158_U133 | ~new_P2_R1158_U309;
  assign new_P2_R1158_U357 = ~new_P2_R1158_U223 | ~new_P2_U3076 | ~new_P2_R1158_U219;
  assign new_P2_R1158_U358 = ~new_P2_R1158_U119 | ~new_P2_R1158_U223;
  assign new_P2_R1158_U359 = ~new_P2_R1158_U236 | ~new_P2_R1158_U5;
  assign new_P2_R1158_U360 = ~new_P2_R1158_U35;
  assign new_P2_R1158_U361 = ~new_P2_R1158_U35 | ~new_P2_R1158_U243;
  assign new_P2_R1158_U362 = ~new_P2_R1158_U262 | ~new_P2_R1158_U9;
  assign new_P2_R1158_U363 = ~new_P2_R1158_U65;
  assign new_P2_R1158_U364 = ~new_P2_R1158_U65 | ~new_P2_R1158_U271;
  assign new_P2_R1158_U365 = ~new_P2_R1158_U20 | ~new_P2_R1158_U366 | ~new_P2_R1158_U307;
  assign new_P2_R1158_U366 = ~new_P2_R1158_U80 | ~new_P2_R1158_U305;
  assign new_P2_R1158_U367 = ~new_P2_R1158_U20;
  assign new_P2_R1158_U368 = ~new_P2_R1158_U64;
  assign new_P2_R1158_U369 = ~new_P2_R1158_U371 | ~new_P2_R1158_U370;
  assign new_P2_R1158_U370 = ~new_P2_R1158_U80 | ~new_P2_R1158_U308 | ~new_P2_R1158_U305;
  assign new_P2_R1158_U371 = ~new_P2_R1158_U367 | ~new_P2_R1158_U308;
  assign new_P2_R1158_U372 = ~new_P2_R1158_U64 | ~new_P2_R1158_U273;
  assign new_P2_R1158_U373 = ~new_P2_R1158_U134 | ~new_P2_R1158_U365;
  assign new_P2_R1158_U374 = ~new_P2_R1158_U135 | ~new_P2_R1158_U192;
  assign new_P2_R1158_U375 = ~new_P2_R1158_U377 | ~new_P2_R1158_U376;
  assign new_P2_R1158_U376 = ~new_P2_R1158_U307 | ~new_P2_R1158_U190 | ~new_P2_R1158_U60;
  assign new_P2_R1158_U377 = ~new_P2_R1158_U20 | ~new_P2_R1158_U366 | ~new_P2_R1158_U307;
  assign new_P2_R1158_U378 = ~new_P2_R1158_U261 | ~new_P2_R1158_U208;
  assign new_P2_R1158_U379 = ~new_P2_R1158_U206;
  assign new_P2_R1158_U380 = ~new_P2_R1158_U11 | ~new_P2_R1158_U208;
  assign new_P2_R1158_U381 = ~new_P2_R1158_U205;
  assign new_P2_R1158_U382 = ~new_P2_R1158_U12 | ~new_P2_R1158_U208;
  assign new_P2_R1158_U383 = ~new_P2_R1158_U203;
  assign new_P2_R1158_U384 = ~new_P2_R1158_U128 | ~new_P2_R1158_U208;
  assign new_P2_R1158_U385 = ~new_P2_R1158_U63;
  assign new_P2_R1158_U386 = ~new_P2_R1158_U235 | ~new_P2_R1158_U165;
  assign new_P2_R1158_U387 = ~new_P2_R1158_U36;
  assign new_P2_R1158_U388 = ~new_P2_R1158_U10 | ~new_P2_R1158_U165;
  assign new_P2_R1158_U389 = ~new_P2_R1158_U163;
  assign new_P2_R1158_U390 = ~new_P2_R1158_U121 | ~new_P2_R1158_U165;
  assign new_P2_R1158_U391 = ~new_P2_R1158_U161;
  assign new_P2_R1158_U392 = ~new_P2_R1158_U138 | ~new_P2_R1158_U209;
  assign new_P2_R1158_U393 = ~new_P2_R1158_U139 | ~new_P2_R1158_U13;
  assign new_P2_R1158_U394 = ~new_P2_R1158_U140 | ~new_P2_R1158_U316;
  assign new_P2_R1158_U395 = ~new_P2_U3152 | ~new_P2_R1158_U150;
  assign new_P2_R1158_U396 = ~new_P2_U3416 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U397 = ~new_P2_R1158_U67;
  assign new_P2_R1158_U398 = ~new_P2_R1158_U397 | ~new_P2_U3082;
  assign new_P2_R1158_U399 = ~new_P2_R1158_U67 | ~new_P2_R1158_U34;
  assign new_P2_R1158_U400 = ~new_P2_R1158_U397 | ~new_P2_U3082;
  assign new_P2_R1158_U401 = ~new_P2_R1158_U67 | ~new_P2_R1158_U34;
  assign new_P2_R1158_U402 = ~new_P2_R1158_U401 | ~new_P2_R1158_U400;
  assign new_P2_R1158_U403 = ~new_P2_U3152 | ~new_P2_R1158_U152;
  assign new_P2_R1158_U404 = ~new_P2_U3401 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U405 = ~new_P2_R1158_U76;
  assign new_P2_R1158_U406 = ~new_P2_U3152 | ~new_P2_R1158_U153;
  assign new_P2_R1158_U407 = ~new_P2_U3392 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U408 = ~new_P2_R1158_U74;
  assign new_P2_R1158_U409 = ~new_P2_U3152 | ~new_P2_R1158_U154;
  assign new_P2_R1158_U410 = ~new_P2_U3387 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U411 = ~new_P2_R1158_U75;
  assign new_P2_R1158_U412 = ~new_P2_U3152 | ~new_P2_R1158_U155;
  assign new_P2_R1158_U413 = ~new_P2_U3398 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U414 = ~new_P2_R1158_U73;
  assign new_P2_R1158_U415 = ~new_P2_U3152 | ~new_P2_R1158_U156;
  assign new_P2_R1158_U416 = ~new_P2_U3395 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U417 = ~new_P2_R1158_U72;
  assign new_P2_R1158_U418 = ~new_P2_U3152 | ~new_P2_R1158_U157;
  assign new_P2_R1158_U419 = ~new_P2_U3404 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U420 = ~new_P2_R1158_U71;
  assign new_P2_R1158_U421 = ~new_P2_U3152 | ~new_P2_R1158_U158;
  assign new_P2_R1158_U422 = ~new_P2_U3410 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U423 = ~new_P2_R1158_U70;
  assign new_P2_R1158_U424 = ~new_P2_U3152 | ~new_P2_R1158_U159;
  assign new_P2_R1158_U425 = ~new_P2_U3407 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U426 = ~new_P2_R1158_U69;
  assign new_P2_R1158_U427 = ~new_P2_U3152 | ~new_P2_R1158_U160;
  assign new_P2_R1158_U428 = ~new_P2_U3413 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U429 = ~new_P2_R1158_U68;
  assign new_P2_R1158_U430 = ~new_P2_R1158_U151 | ~new_P2_R1158_U161;
  assign new_P2_R1158_U431 = ~new_P2_R1158_U391 | ~new_P2_R1158_U402;
  assign new_P2_R1158_U432 = ~new_P2_R1158_U429 | ~new_P2_U3083;
  assign new_P2_R1158_U433 = ~new_P2_R1158_U68 | ~new_P2_R1158_U22;
  assign new_P2_R1158_U434 = ~new_P2_R1158_U429 | ~new_P2_U3083;
  assign new_P2_R1158_U435 = ~new_P2_R1158_U68 | ~new_P2_R1158_U22;
  assign new_P2_R1158_U436 = ~new_P2_R1158_U435 | ~new_P2_R1158_U434;
  assign new_P2_R1158_U437 = ~new_P2_R1158_U162 | ~new_P2_R1158_U163;
  assign new_P2_R1158_U438 = ~new_P2_R1158_U389 | ~new_P2_R1158_U436;
  assign new_P2_R1158_U439 = ~new_P2_R1158_U423 | ~new_P2_U3069;
  assign new_P2_R1158_U440 = ~new_P2_R1158_U70 | ~new_P2_R1158_U25;
  assign new_P2_R1158_U441 = ~new_P2_R1158_U426 | ~new_P2_U3070;
  assign new_P2_R1158_U442 = ~new_P2_R1158_U69 | ~new_P2_R1158_U23;
  assign new_P2_R1158_U443 = ~new_P2_R1158_U442 | ~new_P2_R1158_U441;
  assign new_P2_R1158_U444 = ~new_P2_R1158_U36 | ~new_P2_R1158_U345;
  assign new_P2_R1158_U445 = ~new_P2_R1158_U443 | ~new_P2_R1158_U387;
  assign new_P2_R1158_U446 = ~new_P2_R1158_U420 | ~new_P2_U3066;
  assign new_P2_R1158_U447 = ~new_P2_R1158_U71 | ~new_P2_R1158_U26;
  assign new_P2_R1158_U448 = ~new_P2_R1158_U420 | ~new_P2_U3066;
  assign new_P2_R1158_U449 = ~new_P2_R1158_U71 | ~new_P2_R1158_U26;
  assign new_P2_R1158_U450 = ~new_P2_R1158_U449 | ~new_P2_R1158_U448;
  assign new_P2_R1158_U451 = ~new_P2_R1158_U164 | ~new_P2_R1158_U165;
  assign new_P2_R1158_U452 = ~new_P2_R1158_U234 | ~new_P2_R1158_U450;
  assign new_P2_R1158_U453 = ~new_P2_R1158_U405 | ~new_P2_U3059;
  assign new_P2_R1158_U454 = ~new_P2_R1158_U76 | ~new_P2_R1158_U33;
  assign new_P2_R1158_U455 = ~new_P2_R1158_U405 | ~new_P2_U3059;
  assign new_P2_R1158_U456 = ~new_P2_R1158_U76 | ~new_P2_R1158_U33;
  assign new_P2_R1158_U457 = ~new_P2_R1158_U456 | ~new_P2_R1158_U455;
  assign new_P2_R1158_U458 = ~new_P2_R1158_U166 | ~new_P2_R1158_U167;
  assign new_P2_R1158_U459 = ~new_P2_R1158_U232 | ~new_P2_R1158_U457;
  assign new_P2_R1158_U460 = ~new_P2_R1158_U414 | ~new_P2_U3063;
  assign new_P2_R1158_U461 = ~new_P2_R1158_U73 | ~new_P2_R1158_U30;
  assign new_P2_R1158_U462 = ~new_P2_R1158_U417 | ~new_P2_U3067;
  assign new_P2_R1158_U463 = ~new_P2_R1158_U72 | ~new_P2_R1158_U28;
  assign new_P2_R1158_U464 = ~new_P2_R1158_U463 | ~new_P2_R1158_U462;
  assign new_P2_R1158_U465 = ~new_P2_R1158_U346 | ~new_P2_R1158_U37;
  assign new_P2_R1158_U466 = ~new_P2_R1158_U464 | ~new_P2_R1158_U225;
  assign new_P2_R1158_U467 = ~new_P2_U3152 | ~new_P2_R1158_U168;
  assign new_P2_R1158_U468 = ~new_P2_U3896 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U469 = ~new_P2_R1158_U77;
  assign new_P2_R1158_U470 = ~new_P2_U3152 | ~new_P2_R1158_U169;
  assign new_P2_R1158_U471 = ~new_P2_U3431 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U472 = ~new_P2_R1158_U84;
  assign new_P2_R1158_U473 = ~new_P2_U3152 | ~new_P2_R1158_U170;
  assign new_P2_R1158_U474 = ~new_P2_U3419 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U475 = ~new_P2_R1158_U88;
  assign new_P2_R1158_U476 = ~new_P2_U3152 | ~new_P2_R1158_U171;
  assign new_P2_R1158_U477 = ~new_P2_U3422 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U478 = ~new_P2_R1158_U87;
  assign new_P2_R1158_U479 = ~new_P2_U3152 | ~new_P2_R1158_U172;
  assign new_P2_R1158_U480 = ~new_P2_U3428 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U481 = ~new_P2_R1158_U86;
  assign new_P2_R1158_U482 = ~new_P2_U3152 | ~new_P2_R1158_U173;
  assign new_P2_R1158_U483 = ~new_P2_U3425 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U484 = ~new_P2_R1158_U85;
  assign new_P2_R1158_U485 = ~new_P2_U3152 | ~new_P2_R1158_U174;
  assign new_P2_R1158_U486 = ~new_P2_U3434 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U487 = ~new_P2_R1158_U83;
  assign new_P2_R1158_U488 = ~new_P2_U3152 | ~new_P2_R1158_U175;
  assign new_P2_R1158_U489 = ~new_P2_U3440 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U490 = ~new_P2_R1158_U82;
  assign new_P2_R1158_U491 = ~new_P2_U3152 | ~new_P2_R1158_U176;
  assign new_P2_R1158_U492 = ~new_P2_U3437 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U493 = ~new_P2_R1158_U81;
  assign new_P2_R1158_U494 = ~new_P2_U3152 | ~new_P2_R1158_U177;
  assign new_P2_R1158_U495 = ~new_P2_U3443 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U496 = ~new_P2_R1158_U89;
  assign new_P2_R1158_U497 = ~new_P2_U3152 | ~new_P2_R1158_U178;
  assign new_P2_R1158_U498 = ~new_P2_U3902 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U499 = ~new_P2_R1158_U91;
  assign new_P2_R1158_U500 = ~new_P2_U3152 | ~new_P2_R1158_U179;
  assign new_P2_R1158_U501 = ~new_P2_U3903 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U502 = ~new_P2_R1158_U92;
  assign new_P2_R1158_U503 = ~new_P2_U3152 | ~new_P2_R1158_U180;
  assign new_P2_R1158_U504 = ~new_P2_U3445 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U505 = ~new_P2_R1158_U90;
  assign new_P2_R1158_U506 = ~new_P2_U3152 | ~new_P2_R1158_U181;
  assign new_P2_R1158_U507 = ~new_P2_U3901 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U508 = ~new_P2_R1158_U93;
  assign new_P2_R1158_U509 = ~new_P2_U3152 | ~new_P2_R1158_U182;
  assign new_P2_R1158_U510 = ~new_P2_U3900 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U511 = ~new_P2_R1158_U94;
  assign new_P2_R1158_U512 = ~new_P2_U3152 | ~new_P2_R1158_U183;
  assign new_P2_R1158_U513 = ~new_P2_U3897 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U514 = ~new_P2_R1158_U80;
  assign new_P2_R1158_U515 = ~new_P2_U3152 | ~new_P2_R1158_U184;
  assign new_P2_R1158_U516 = ~new_P2_U3898 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U517 = ~new_P2_R1158_U78;
  assign new_P2_R1158_U518 = ~new_P2_U3152 | ~new_P2_R1158_U185;
  assign new_P2_R1158_U519 = ~new_P2_U3899 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U520 = ~new_P2_R1158_U79;
  assign new_P2_R1158_U521 = ~new_P2_U3152 | ~new_P2_R1158_U186;
  assign new_P2_R1158_U522 = ~new_P2_U3053 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U523 = ~new_P2_R1158_U137;
  assign new_P2_R1158_U524 = ~new_P2_U3895 | ~new_P2_R1158_U523;
  assign new_P2_R1158_U525 = ~new_P2_R1158_U137 | ~new_P2_R1158_U187;
  assign new_P2_R1158_U526 = ~new_P2_R1158_U95;
  assign new_P2_R1158_U527 = ~new_P2_R1158_U526 | ~new_P2_R1158_U356 | ~new_P2_R1158_U312;
  assign new_P2_R1158_U528 = ~new_P2_R1158_U95 | ~new_P2_R1158_U136 | ~new_P2_R1158_U374;
  assign new_P2_R1158_U529 = ~new_P2_R1158_U469 | ~new_P2_U3052;
  assign new_P2_R1158_U530 = ~new_P2_R1158_U77 | ~new_P2_R1158_U38;
  assign new_P2_R1158_U531 = ~new_P2_R1158_U469 | ~new_P2_U3052;
  assign new_P2_R1158_U532 = ~new_P2_R1158_U77 | ~new_P2_R1158_U38;
  assign new_P2_R1158_U533 = ~new_P2_R1158_U532 | ~new_P2_R1158_U531;
  assign new_P2_R1158_U534 = ~new_P2_R1158_U188 | ~new_P2_R1158_U189;
  assign new_P2_R1158_U535 = ~new_P2_R1158_U311 | ~new_P2_R1158_U533;
  assign new_P2_R1158_U536 = ~new_P2_R1158_U514 | ~new_P2_U3056;
  assign new_P2_R1158_U537 = ~new_P2_R1158_U80 | ~new_P2_R1158_U41;
  assign new_P2_R1158_U538 = ~new_P2_R1158_U190 | ~new_P2_R1158_U141 | ~new_P2_R1158_U61;
  assign new_P2_R1158_U539 = ~new_P2_R1158_U218 | ~new_P2_R1158_U318 | ~new_P2_R1158_U209;
  assign new_P2_R1158_U540 = ~new_P2_R1158_U517 | ~new_P2_U3057;
  assign new_P2_R1158_U541 = ~new_P2_R1158_U78 | ~new_P2_R1158_U39;
  assign new_P2_R1158_U542 = ~new_P2_R1158_U541 | ~new_P2_R1158_U540;
  assign new_P2_R1158_U543 = ~new_P2_R1158_U347 | ~new_P2_R1158_U191;
  assign new_P2_R1158_U544 = ~new_P2_R1158_U317 | ~new_P2_R1158_U542;
  assign new_P2_R1158_U545 = ~new_P2_R1158_U520 | ~new_P2_U3064;
  assign new_P2_R1158_U546 = ~new_P2_R1158_U79 | ~new_P2_R1158_U40;
  assign new_P2_R1158_U547 = ~new_P2_R1158_U546 | ~new_P2_R1158_U545;
  assign new_P2_R1158_U548 = ~new_P2_R1158_U348 | ~new_P2_R1158_U192;
  assign new_P2_R1158_U549 = ~new_P2_R1158_U304 | ~new_P2_R1158_U547;
  assign new_P2_R1158_U550 = ~new_P2_R1158_U511 | ~new_P2_U3065;
  assign new_P2_R1158_U551 = ~new_P2_R1158_U94 | ~new_P2_R1158_U59;
  assign new_P2_R1158_U552 = ~new_P2_R1158_U511 | ~new_P2_U3065;
  assign new_P2_R1158_U553 = ~new_P2_R1158_U94 | ~new_P2_R1158_U59;
  assign new_P2_R1158_U554 = ~new_P2_R1158_U553 | ~new_P2_R1158_U552;
  assign new_P2_R1158_U555 = ~new_P2_R1158_U193 | ~new_P2_R1158_U194;
  assign new_P2_R1158_U556 = ~new_P2_R1158_U300 | ~new_P2_R1158_U554;
  assign new_P2_R1158_U557 = ~new_P2_R1158_U508 | ~new_P2_U3060;
  assign new_P2_R1158_U558 = ~new_P2_R1158_U93 | ~new_P2_R1158_U58;
  assign new_P2_R1158_U559 = ~new_P2_R1158_U508 | ~new_P2_U3060;
  assign new_P2_R1158_U560 = ~new_P2_R1158_U93 | ~new_P2_R1158_U58;
  assign new_P2_R1158_U561 = ~new_P2_R1158_U560 | ~new_P2_R1158_U559;
  assign new_P2_R1158_U562 = ~new_P2_R1158_U195 | ~new_P2_R1158_U196;
  assign new_P2_R1158_U563 = ~new_P2_R1158_U296 | ~new_P2_R1158_U561;
  assign new_P2_R1158_U564 = ~new_P2_R1158_U499 | ~new_P2_U3074;
  assign new_P2_R1158_U565 = ~new_P2_R1158_U91 | ~new_P2_R1158_U57;
  assign new_P2_R1158_U566 = ~new_P2_R1158_U502 | ~new_P2_U3075;
  assign new_P2_R1158_U567 = ~new_P2_R1158_U92 | ~new_P2_R1158_U54;
  assign new_P2_R1158_U568 = ~new_P2_R1158_U567 | ~new_P2_R1158_U566;
  assign new_P2_R1158_U569 = ~new_P2_R1158_U349 | ~new_P2_R1158_U62;
  assign new_P2_R1158_U570 = ~new_P2_R1158_U568 | ~new_P2_R1158_U321;
  assign new_P2_R1158_U571 = ~new_P2_R1158_U408 | ~new_P2_U3077;
  assign new_P2_R1158_U572 = ~new_P2_R1158_U74 | ~new_P2_R1158_U31;
  assign new_P2_R1158_U573 = ~new_P2_R1158_U408 | ~new_P2_U3077;
  assign new_P2_R1158_U574 = ~new_P2_R1158_U74 | ~new_P2_R1158_U31;
  assign new_P2_R1158_U575 = ~new_P2_R1158_U574 | ~new_P2_R1158_U573;
  assign new_P2_R1158_U576 = ~new_P2_R1158_U197 | ~new_P2_R1158_U198;
  assign new_P2_R1158_U577 = ~new_P2_R1158_U222 | ~new_P2_R1158_U575;
  assign new_P2_R1158_U578 = ~new_P2_R1158_U505 | ~new_P2_U3080;
  assign new_P2_R1158_U579 = ~new_P2_R1158_U90 | ~new_P2_R1158_U55;
  assign new_P2_R1158_U580 = ~new_P2_R1158_U579 | ~new_P2_R1158_U578;
  assign new_P2_R1158_U581 = ~new_P2_R1158_U350 | ~new_P2_R1158_U199;
  assign new_P2_R1158_U582 = ~new_P2_R1158_U286 | ~new_P2_R1158_U580;
  assign new_P2_R1158_U583 = ~new_P2_R1158_U496 | ~new_P2_U3081;
  assign new_P2_R1158_U584 = ~new_P2_R1158_U89 | ~new_P2_R1158_U53;
  assign new_P2_R1158_U585 = ~new_P2_R1158_U496 | ~new_P2_U3081;
  assign new_P2_R1158_U586 = ~new_P2_R1158_U89 | ~new_P2_R1158_U53;
  assign new_P2_R1158_U587 = ~new_P2_R1158_U586 | ~new_P2_R1158_U585;
  assign new_P2_R1158_U588 = ~new_P2_R1158_U200 | ~new_P2_R1158_U201;
  assign new_P2_R1158_U589 = ~new_P2_R1158_U282 | ~new_P2_R1158_U587;
  assign new_P2_R1158_U590 = ~new_P2_R1158_U490 | ~new_P2_U3068;
  assign new_P2_R1158_U591 = ~new_P2_R1158_U82 | ~new_P2_R1158_U44;
  assign new_P2_R1158_U592 = ~new_P2_R1158_U493 | ~new_P2_U3072;
  assign new_P2_R1158_U593 = ~new_P2_R1158_U81 | ~new_P2_R1158_U42;
  assign new_P2_R1158_U594 = ~new_P2_R1158_U593 | ~new_P2_R1158_U592;
  assign new_P2_R1158_U595 = ~new_P2_R1158_U63 | ~new_P2_R1158_U351;
  assign new_P2_R1158_U596 = ~new_P2_R1158_U594 | ~new_P2_R1158_U385;
  assign new_P2_R1158_U597 = ~new_P2_R1158_U487 | ~new_P2_U3073;
  assign new_P2_R1158_U598 = ~new_P2_R1158_U83 | ~new_P2_R1158_U45;
  assign new_P2_R1158_U599 = ~new_P2_R1158_U487 | ~new_P2_U3073;
  assign new_P2_R1158_U600 = ~new_P2_R1158_U83 | ~new_P2_R1158_U45;
  assign new_P2_R1158_U601 = ~new_P2_R1158_U600 | ~new_P2_R1158_U599;
  assign new_P2_R1158_U602 = ~new_P2_R1158_U202 | ~new_P2_R1158_U203;
  assign new_P2_R1158_U603 = ~new_P2_R1158_U383 | ~new_P2_R1158_U601;
  assign new_P2_R1158_U604 = ~new_P2_R1158_U472 | ~new_P2_U3078;
  assign new_P2_R1158_U605 = ~new_P2_R1158_U84 | ~new_P2_R1158_U46;
  assign new_P2_R1158_U606 = ~new_P2_R1158_U472 | ~new_P2_U3078;
  assign new_P2_R1158_U607 = ~new_P2_R1158_U84 | ~new_P2_R1158_U46;
  assign new_P2_R1158_U608 = ~new_P2_R1158_U607 | ~new_P2_R1158_U606;
  assign new_P2_R1158_U609 = ~new_P2_R1158_U204 | ~new_P2_R1158_U205;
  assign new_P2_R1158_U610 = ~new_P2_R1158_U381 | ~new_P2_R1158_U608;
  assign new_P2_R1158_U611 = ~new_P2_R1158_U481 | ~new_P2_U3079;
  assign new_P2_R1158_U612 = ~new_P2_R1158_U86 | ~new_P2_R1158_U50;
  assign new_P2_R1158_U613 = ~new_P2_R1158_U484 | ~new_P2_U3071;
  assign new_P2_R1158_U614 = ~new_P2_R1158_U85 | ~new_P2_R1158_U47;
  assign new_P2_R1158_U615 = ~new_P2_R1158_U614 | ~new_P2_R1158_U613;
  assign new_P2_R1158_U616 = ~new_P2_R1158_U352 | ~new_P2_R1158_U66;
  assign new_P2_R1158_U617 = ~new_P2_R1158_U615 | ~new_P2_R1158_U337;
  assign new_P2_R1158_U618 = ~new_P2_R1158_U478 | ~new_P2_U3062;
  assign new_P2_R1158_U619 = ~new_P2_R1158_U87 | ~new_P2_R1158_U48;
  assign new_P2_R1158_U620 = ~new_P2_R1158_U619 | ~new_P2_R1158_U618;
  assign new_P2_R1158_U621 = ~new_P2_R1158_U206 | ~new_P2_R1158_U353;
  assign new_P2_R1158_U622 = ~new_P2_R1158_U379 | ~new_P2_R1158_U620;
  assign new_P2_R1158_U623 = ~new_P2_R1158_U475 | ~new_P2_U3061;
  assign new_P2_R1158_U624 = ~new_P2_R1158_U88 | ~new_P2_R1158_U51;
  assign new_P2_R1158_U625 = ~new_P2_R1158_U475 | ~new_P2_U3061;
  assign new_P2_R1158_U626 = ~new_P2_R1158_U88 | ~new_P2_R1158_U51;
  assign new_P2_R1158_U627 = ~new_P2_R1158_U626 | ~new_P2_R1158_U625;
  assign new_P2_R1158_U628 = ~new_P2_R1158_U207 | ~new_P2_R1158_U208;
  assign new_P2_R1158_U629 = ~new_P2_R1158_U260 | ~new_P2_R1158_U627;
  assign new_P2_R1158_U630 = ~new_P2_R1158_U75 | ~new_P2_R1158_U21;
  assign new_P2_R1158_U631 = ~new_P2_R1158_U411 | ~new_P2_U3152;
  assign new_P2_R1158_U632 = ~new_P2_R1158_U149;
  assign new_P2_R1158_U633 = ~new_P2_R1158_U632 | ~new_P2_U3076;
  assign new_P2_R1158_U634 = ~new_P2_R1158_U149 | ~new_P2_R1158_U32;
  assign new_P2_R1131_U6 = new_P2_R1131_U212 & new_P2_R1131_U211;
  assign new_P2_R1131_U7 = new_P2_R1131_U246 & new_P2_R1131_U245;
  assign new_P2_R1131_U8 = new_P2_R1131_U193 & new_P2_R1131_U257;
  assign new_P2_R1131_U9 = new_P2_R1131_U259 & new_P2_R1131_U258;
  assign new_P2_R1131_U10 = new_P2_R1131_U194 & new_P2_R1131_U281;
  assign new_P2_R1131_U11 = new_P2_R1131_U283 & new_P2_R1131_U282;
  assign new_P2_R1131_U12 = new_P2_R1131_U299 & new_P2_R1131_U195;
  assign new_P2_R1131_U13 = new_P2_R1131_U215 & new_P2_R1131_U210 & new_P2_R1131_U197;
  assign new_P2_R1131_U14 = new_P2_R1131_U220 & new_P2_R1131_U198;
  assign new_P2_R1131_U15 = new_P2_R1131_U244 & new_P2_R1131_U224 & new_P2_R1131_U192;
  assign new_P2_R1131_U16 = new_P2_R1131_U399 & new_P2_R1131_U398;
  assign new_P2_R1131_U17 = ~new_P2_R1131_U331 | ~new_P2_R1131_U334;
  assign new_P2_R1131_U18 = ~new_P2_R1131_U322 | ~new_P2_R1131_U325;
  assign new_P2_R1131_U19 = ~new_P2_R1131_U311 | ~new_P2_R1131_U314;
  assign new_P2_R1131_U20 = ~new_P2_R1131_U305 | ~new_P2_R1131_U357;
  assign new_P2_R1131_U21 = ~new_P2_R1131_U137 | ~new_P2_R1131_U186;
  assign new_P2_R1131_U22 = ~new_P2_R1131_U242 | ~new_P2_R1131_U347;
  assign new_P2_R1131_U23 = ~new_P2_R1131_U235 | ~new_P2_R1131_U238;
  assign new_P2_R1131_U24 = ~new_P2_R1131_U227 | ~new_P2_R1131_U229;
  assign new_P2_R1131_U25 = ~new_P2_R1131_U175 | ~new_P2_R1131_U337;
  assign new_P2_R1131_U26 = ~new_P2_U3069;
  assign new_P2_R1131_U27 = ~new_P2_U3069 | ~new_P2_R1131_U32;
  assign new_P2_R1131_U28 = ~new_P2_U3083;
  assign new_P2_R1131_U29 = ~new_P2_U3404;
  assign new_P2_R1131_U30 = ~new_P2_U3407;
  assign new_P2_R1131_U31 = ~new_P2_U3401;
  assign new_P2_R1131_U32 = ~new_P2_U3410;
  assign new_P2_R1131_U33 = ~new_P2_U3413;
  assign new_P2_R1131_U34 = ~new_P2_U3067;
  assign new_P2_R1131_U35 = ~new_P2_U3067 | ~new_P2_R1131_U37;
  assign new_P2_R1131_U36 = ~new_P2_U3063;
  assign new_P2_R1131_U37 = ~new_P2_U3395;
  assign new_P2_R1131_U38 = ~new_P2_U3387;
  assign new_P2_R1131_U39 = ~new_P2_U3077;
  assign new_P2_R1131_U40 = ~new_P2_U3398;
  assign new_P2_R1131_U41 = ~new_P2_U3070;
  assign new_P2_R1131_U42 = ~new_P2_U3066;
  assign new_P2_R1131_U43 = ~new_P2_U3059;
  assign new_P2_R1131_U44 = ~new_P2_U3059 | ~new_P2_R1131_U31;
  assign new_P2_R1131_U45 = ~new_P2_R1131_U216 | ~new_P2_R1131_U214;
  assign new_P2_R1131_U46 = ~new_P2_U3416;
  assign new_P2_R1131_U47 = ~new_P2_U3082;
  assign new_P2_R1131_U48 = ~new_P2_R1131_U45 | ~new_P2_R1131_U217;
  assign new_P2_R1131_U49 = ~new_P2_R1131_U44 | ~new_P2_R1131_U231;
  assign new_P2_R1131_U50 = ~new_P2_R1131_U338 | ~new_P2_R1131_U204 | ~new_P2_R1131_U188;
  assign new_P2_R1131_U51 = ~new_P2_U3895;
  assign new_P2_R1131_U52 = ~new_P2_U3056;
  assign new_P2_R1131_U53 = ~new_P2_U3056 | ~new_P2_R1131_U90;
  assign new_P2_R1131_U54 = ~new_P2_U3052;
  assign new_P2_R1131_U55 = ~new_P2_U3071;
  assign new_P2_R1131_U56 = ~new_P2_U3062;
  assign new_P2_R1131_U57 = ~new_P2_U3061;
  assign new_P2_R1131_U58 = ~new_P2_U3419;
  assign new_P2_R1131_U59 = ~new_P2_U3082 | ~new_P2_R1131_U46;
  assign new_P2_R1131_U60 = ~new_P2_U3422;
  assign new_P2_R1131_U61 = ~new_P2_U3425;
  assign new_P2_R1131_U62 = ~new_P2_R1131_U249 | ~new_P2_R1131_U248;
  assign new_P2_R1131_U63 = ~new_P2_U3428;
  assign new_P2_R1131_U64 = ~new_P2_U3079;
  assign new_P2_R1131_U65 = ~new_P2_U3437;
  assign new_P2_R1131_U66 = ~new_P2_U3434;
  assign new_P2_R1131_U67 = ~new_P2_U3431;
  assign new_P2_R1131_U68 = ~new_P2_U3072;
  assign new_P2_R1131_U69 = ~new_P2_U3073;
  assign new_P2_R1131_U70 = ~new_P2_U3078;
  assign new_P2_R1131_U71 = ~new_P2_U3078 | ~new_P2_R1131_U67;
  assign new_P2_R1131_U72 = ~new_P2_U3440;
  assign new_P2_R1131_U73 = ~new_P2_U3068;
  assign new_P2_R1131_U74 = ~new_P2_U3081;
  assign new_P2_R1131_U75 = ~new_P2_U3445;
  assign new_P2_R1131_U76 = ~new_P2_U3080;
  assign new_P2_R1131_U77 = ~new_P2_U3903;
  assign new_P2_R1131_U78 = ~new_P2_U3075;
  assign new_P2_R1131_U79 = ~new_P2_U3900;
  assign new_P2_R1131_U80 = ~new_P2_U3901;
  assign new_P2_R1131_U81 = ~new_P2_U3902;
  assign new_P2_R1131_U82 = ~new_P2_U3065;
  assign new_P2_R1131_U83 = ~new_P2_U3060;
  assign new_P2_R1131_U84 = ~new_P2_U3074;
  assign new_P2_R1131_U85 = ~new_P2_U3074 | ~new_P2_R1131_U81;
  assign new_P2_R1131_U86 = ~new_P2_U3899;
  assign new_P2_R1131_U87 = ~new_P2_U3064;
  assign new_P2_R1131_U88 = ~new_P2_U3898;
  assign new_P2_R1131_U89 = ~new_P2_U3057;
  assign new_P2_R1131_U90 = ~new_P2_U3897;
  assign new_P2_R1131_U91 = ~new_P2_U3896;
  assign new_P2_R1131_U92 = ~new_P2_U3053;
  assign new_P2_R1131_U93 = ~new_P2_R1131_U297 | ~new_P2_R1131_U296;
  assign new_P2_R1131_U94 = ~new_P2_R1131_U85 | ~new_P2_R1131_U307;
  assign new_P2_R1131_U95 = ~new_P2_R1131_U71 | ~new_P2_R1131_U318;
  assign new_P2_R1131_U96 = ~new_P2_R1131_U349 | ~new_P2_R1131_U59;
  assign new_P2_R1131_U97 = ~new_P2_U3076;
  assign new_P2_R1131_U98 = ~new_P2_R1131_U406 | ~new_P2_R1131_U405;
  assign new_P2_R1131_U99 = ~new_P2_R1131_U420 | ~new_P2_R1131_U419;
  assign new_P2_R1131_U100 = ~new_P2_R1131_U425 | ~new_P2_R1131_U424;
  assign new_P2_R1131_U101 = ~new_P2_R1131_U441 | ~new_P2_R1131_U440;
  assign new_P2_R1131_U102 = ~new_P2_R1131_U446 | ~new_P2_R1131_U445;
  assign new_P2_R1131_U103 = ~new_P2_R1131_U451 | ~new_P2_R1131_U450;
  assign new_P2_R1131_U104 = ~new_P2_R1131_U456 | ~new_P2_R1131_U455;
  assign new_P2_R1131_U105 = ~new_P2_R1131_U461 | ~new_P2_R1131_U460;
  assign new_P2_R1131_U106 = ~new_P2_R1131_U477 | ~new_P2_R1131_U476;
  assign new_P2_R1131_U107 = ~new_P2_R1131_U482 | ~new_P2_R1131_U481;
  assign new_P2_R1131_U108 = ~new_P2_R1131_U365 | ~new_P2_R1131_U364;
  assign new_P2_R1131_U109 = ~new_P2_R1131_U374 | ~new_P2_R1131_U373;
  assign new_P2_R1131_U110 = ~new_P2_R1131_U381 | ~new_P2_R1131_U380;
  assign new_P2_R1131_U111 = ~new_P2_R1131_U385 | ~new_P2_R1131_U384;
  assign new_P2_R1131_U112 = ~new_P2_R1131_U394 | ~new_P2_R1131_U393;
  assign new_P2_R1131_U113 = ~new_P2_R1131_U415 | ~new_P2_R1131_U414;
  assign new_P2_R1131_U114 = ~new_P2_R1131_U432 | ~new_P2_R1131_U431;
  assign new_P2_R1131_U115 = ~new_P2_R1131_U436 | ~new_P2_R1131_U435;
  assign new_P2_R1131_U116 = ~new_P2_R1131_U468 | ~new_P2_R1131_U467;
  assign new_P2_R1131_U117 = ~new_P2_R1131_U472 | ~new_P2_R1131_U471;
  assign new_P2_R1131_U118 = ~new_P2_R1131_U489 | ~new_P2_R1131_U488;
  assign new_P2_R1131_U119 = new_P2_R1131_U206 & new_P2_R1131_U196;
  assign new_P2_R1131_U120 = new_P2_R1131_U209 & new_P2_R1131_U208;
  assign new_P2_R1131_U121 = new_P2_R1131_U14 & new_P2_R1131_U13;
  assign new_P2_R1131_U122 = new_P2_R1131_U340 & new_P2_R1131_U222;
  assign new_P2_R1131_U123 = new_P2_R1131_U342 & new_P2_R1131_U122;
  assign new_P2_R1131_U124 = new_P2_R1131_U27 & new_P2_R1131_U367 & new_P2_R1131_U366;
  assign new_P2_R1131_U125 = new_P2_R1131_U370 & new_P2_R1131_U198;
  assign new_P2_R1131_U126 = new_P2_R1131_U237 & new_P2_R1131_U6;
  assign new_P2_R1131_U127 = new_P2_R1131_U377 & new_P2_R1131_U197;
  assign new_P2_R1131_U128 = new_P2_R1131_U35 & new_P2_R1131_U387 & new_P2_R1131_U386;
  assign new_P2_R1131_U129 = new_P2_R1131_U390 & new_P2_R1131_U196;
  assign new_P2_R1131_U130 = new_P2_R1131_U251 & new_P2_R1131_U15;
  assign new_P2_R1131_U131 = new_P2_R1131_U343 & new_P2_R1131_U252;
  assign new_P2_R1131_U132 = new_P2_R1131_U262 & new_P2_R1131_U8;
  assign new_P2_R1131_U133 = new_P2_R1131_U286 & new_P2_R1131_U10;
  assign new_P2_R1131_U134 = new_P2_R1131_U302 & new_P2_R1131_U301;
  assign new_P2_R1131_U135 = new_P2_R1131_U397 & new_P2_R1131_U303;
  assign new_P2_R1131_U136 = new_P2_R1131_U16 & new_P2_R1131_U304 & new_P2_R1131_U302 & new_P2_R1131_U301;
  assign new_P2_R1131_U137 = new_P2_R1131_U359 & new_P2_R1131_U165;
  assign new_P2_R1131_U138 = ~new_P2_R1131_U403 | ~new_P2_R1131_U402;
  assign new_P2_R1131_U139 = new_P2_R1131_U53 & new_P2_R1131_U408 & new_P2_R1131_U407;
  assign new_P2_R1131_U140 = new_P2_R1131_U411 & new_P2_R1131_U195;
  assign new_P2_R1131_U141 = ~new_P2_R1131_U417 | ~new_P2_R1131_U416;
  assign new_P2_R1131_U142 = ~new_P2_R1131_U422 | ~new_P2_R1131_U421;
  assign new_P2_R1131_U143 = new_P2_R1131_U313 & new_P2_R1131_U11;
  assign new_P2_R1131_U144 = new_P2_R1131_U428 & new_P2_R1131_U194;
  assign new_P2_R1131_U145 = ~new_P2_R1131_U438 | ~new_P2_R1131_U437;
  assign new_P2_R1131_U146 = ~new_P2_R1131_U443 | ~new_P2_R1131_U442;
  assign new_P2_R1131_U147 = ~new_P2_R1131_U448 | ~new_P2_R1131_U447;
  assign new_P2_R1131_U148 = ~new_P2_R1131_U453 | ~new_P2_R1131_U452;
  assign new_P2_R1131_U149 = ~new_P2_R1131_U458 | ~new_P2_R1131_U457;
  assign new_P2_R1131_U150 = new_P2_R1131_U324 & new_P2_R1131_U9;
  assign new_P2_R1131_U151 = new_P2_R1131_U464 & new_P2_R1131_U193;
  assign new_P2_R1131_U152 = ~new_P2_R1131_U474 | ~new_P2_R1131_U473;
  assign new_P2_R1131_U153 = ~new_P2_R1131_U479 | ~new_P2_R1131_U478;
  assign new_P2_R1131_U154 = new_P2_R1131_U333 & new_P2_R1131_U7;
  assign new_P2_R1131_U155 = new_P2_R1131_U485 & new_P2_R1131_U192;
  assign new_P2_R1131_U156 = new_P2_R1131_U363 & new_P2_R1131_U362;
  assign new_P2_R1131_U157 = ~new_P2_R1131_U123 | ~new_P2_R1131_U341;
  assign new_P2_R1131_U158 = new_P2_R1131_U372 & new_P2_R1131_U371;
  assign new_P2_R1131_U159 = new_P2_R1131_U379 & new_P2_R1131_U378;
  assign new_P2_R1131_U160 = new_P2_R1131_U383 & new_P2_R1131_U382;
  assign new_P2_R1131_U161 = ~new_P2_R1131_U120 | ~new_P2_R1131_U344;
  assign new_P2_R1131_U162 = new_P2_R1131_U392 & new_P2_R1131_U391;
  assign new_P2_R1131_U163 = ~new_P2_U3904;
  assign new_P2_R1131_U164 = ~new_P2_U3054;
  assign new_P2_R1131_U165 = new_P2_R1131_U401 & new_P2_R1131_U400;
  assign new_P2_R1131_U166 = ~new_P2_R1131_U134 | ~new_P2_R1131_U360;
  assign new_P2_R1131_U167 = new_P2_R1131_U413 & new_P2_R1131_U412;
  assign new_P2_R1131_U168 = ~new_P2_R1131_U293 | ~new_P2_R1131_U292;
  assign new_P2_R1131_U169 = ~new_P2_R1131_U289 | ~new_P2_R1131_U288;
  assign new_P2_R1131_U170 = new_P2_R1131_U430 & new_P2_R1131_U429;
  assign new_P2_R1131_U171 = new_P2_R1131_U434 & new_P2_R1131_U433;
  assign new_P2_R1131_U172 = ~new_P2_R1131_U279 | ~new_P2_R1131_U278;
  assign new_P2_R1131_U173 = ~new_P2_R1131_U275 | ~new_P2_R1131_U274;
  assign new_P2_R1131_U174 = ~new_P2_U3392;
  assign new_P2_R1131_U175 = ~new_P2_U3387 | ~new_P2_R1131_U97;
  assign new_P2_R1131_U176 = ~new_P2_R1131_U339 | ~new_P2_R1131_U271 | ~new_P2_R1131_U187;
  assign new_P2_R1131_U177 = ~new_P2_U3443;
  assign new_P2_R1131_U178 = ~new_P2_R1131_U269 | ~new_P2_R1131_U268;
  assign new_P2_R1131_U179 = ~new_P2_R1131_U265 | ~new_P2_R1131_U264;
  assign new_P2_R1131_U180 = new_P2_R1131_U466 & new_P2_R1131_U465;
  assign new_P2_R1131_U181 = new_P2_R1131_U470 & new_P2_R1131_U469;
  assign new_P2_R1131_U182 = ~new_P2_R1131_U255 | ~new_P2_R1131_U254;
  assign new_P2_R1131_U183 = ~new_P2_R1131_U131 | ~new_P2_R1131_U353;
  assign new_P2_R1131_U184 = ~new_P2_R1131_U351 | ~new_P2_R1131_U62;
  assign new_P2_R1131_U185 = new_P2_R1131_U487 & new_P2_R1131_U486;
  assign new_P2_R1131_U186 = ~new_P2_R1131_U135 | ~new_P2_R1131_U166;
  assign new_P2_R1131_U187 = ~new_P2_R1131_U178 | ~new_P2_R1131_U177;
  assign new_P2_R1131_U188 = ~new_P2_R1131_U175 | ~new_P2_R1131_U174;
  assign new_P2_R1131_U189 = ~new_P2_R1131_U53;
  assign new_P2_R1131_U190 = ~new_P2_R1131_U35;
  assign new_P2_R1131_U191 = ~new_P2_R1131_U27;
  assign new_P2_R1131_U192 = ~new_P2_U3419 | ~new_P2_R1131_U57;
  assign new_P2_R1131_U193 = ~new_P2_U3434 | ~new_P2_R1131_U69;
  assign new_P2_R1131_U194 = ~new_P2_U3901 | ~new_P2_R1131_U83;
  assign new_P2_R1131_U195 = ~new_P2_U3897 | ~new_P2_R1131_U52;
  assign new_P2_R1131_U196 = ~new_P2_U3395 | ~new_P2_R1131_U34;
  assign new_P2_R1131_U197 = ~new_P2_U3404 | ~new_P2_R1131_U42;
  assign new_P2_R1131_U198 = ~new_P2_U3410 | ~new_P2_R1131_U26;
  assign new_P2_R1131_U199 = ~new_P2_R1131_U71;
  assign new_P2_R1131_U200 = ~new_P2_R1131_U85;
  assign new_P2_R1131_U201 = ~new_P2_R1131_U44;
  assign new_P2_R1131_U202 = ~new_P2_R1131_U59;
  assign new_P2_R1131_U203 = ~new_P2_R1131_U175;
  assign new_P2_R1131_U204 = ~new_P2_U3077 | ~new_P2_R1131_U175;
  assign new_P2_R1131_U205 = ~new_P2_R1131_U50;
  assign new_P2_R1131_U206 = ~new_P2_U3398 | ~new_P2_R1131_U36;
  assign new_P2_R1131_U207 = ~new_P2_R1131_U36 | ~new_P2_R1131_U35;
  assign new_P2_R1131_U208 = ~new_P2_R1131_U207 | ~new_P2_R1131_U40;
  assign new_P2_R1131_U209 = ~new_P2_U3063 | ~new_P2_R1131_U190;
  assign new_P2_R1131_U210 = ~new_P2_U3407 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U211 = ~new_P2_U3070 | ~new_P2_R1131_U30;
  assign new_P2_R1131_U212 = ~new_P2_U3066 | ~new_P2_R1131_U29;
  assign new_P2_R1131_U213 = ~new_P2_R1131_U201 | ~new_P2_R1131_U197;
  assign new_P2_R1131_U214 = ~new_P2_R1131_U6 | ~new_P2_R1131_U213;
  assign new_P2_R1131_U215 = ~new_P2_U3401 | ~new_P2_R1131_U43;
  assign new_P2_R1131_U216 = ~new_P2_U3407 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U217 = ~new_P2_R1131_U13 | ~new_P2_R1131_U161;
  assign new_P2_R1131_U218 = ~new_P2_R1131_U45;
  assign new_P2_R1131_U219 = ~new_P2_R1131_U48;
  assign new_P2_R1131_U220 = ~new_P2_U3413 | ~new_P2_R1131_U28;
  assign new_P2_R1131_U221 = ~new_P2_R1131_U28 | ~new_P2_R1131_U27;
  assign new_P2_R1131_U222 = ~new_P2_U3083 | ~new_P2_R1131_U191;
  assign new_P2_R1131_U223 = ~new_P2_R1131_U157;
  assign new_P2_R1131_U224 = ~new_P2_U3416 | ~new_P2_R1131_U47;
  assign new_P2_R1131_U225 = ~new_P2_R1131_U224 | ~new_P2_R1131_U59;
  assign new_P2_R1131_U226 = ~new_P2_R1131_U219 | ~new_P2_R1131_U27;
  assign new_P2_R1131_U227 = ~new_P2_R1131_U125 | ~new_P2_R1131_U226;
  assign new_P2_R1131_U228 = ~new_P2_R1131_U48 | ~new_P2_R1131_U198;
  assign new_P2_R1131_U229 = ~new_P2_R1131_U124 | ~new_P2_R1131_U228;
  assign new_P2_R1131_U230 = ~new_P2_R1131_U27 | ~new_P2_R1131_U198;
  assign new_P2_R1131_U231 = ~new_P2_R1131_U215 | ~new_P2_R1131_U161;
  assign new_P2_R1131_U232 = ~new_P2_R1131_U49;
  assign new_P2_R1131_U233 = ~new_P2_U3066 | ~new_P2_R1131_U29;
  assign new_P2_R1131_U234 = ~new_P2_R1131_U232 | ~new_P2_R1131_U233;
  assign new_P2_R1131_U235 = ~new_P2_R1131_U127 | ~new_P2_R1131_U234;
  assign new_P2_R1131_U236 = ~new_P2_R1131_U49 | ~new_P2_R1131_U197;
  assign new_P2_R1131_U237 = ~new_P2_U3407 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U238 = ~new_P2_R1131_U126 | ~new_P2_R1131_U236;
  assign new_P2_R1131_U239 = ~new_P2_U3066 | ~new_P2_R1131_U29;
  assign new_P2_R1131_U240 = ~new_P2_R1131_U239 | ~new_P2_R1131_U197;
  assign new_P2_R1131_U241 = ~new_P2_R1131_U215 | ~new_P2_R1131_U44;
  assign new_P2_R1131_U242 = ~new_P2_R1131_U129 | ~new_P2_R1131_U348;
  assign new_P2_R1131_U243 = ~new_P2_R1131_U35 | ~new_P2_R1131_U196;
  assign new_P2_R1131_U244 = ~new_P2_U3422 | ~new_P2_R1131_U56;
  assign new_P2_R1131_U245 = ~new_P2_U3062 | ~new_P2_R1131_U60;
  assign new_P2_R1131_U246 = ~new_P2_U3061 | ~new_P2_R1131_U58;
  assign new_P2_R1131_U247 = ~new_P2_R1131_U202 | ~new_P2_R1131_U192;
  assign new_P2_R1131_U248 = ~new_P2_R1131_U7 | ~new_P2_R1131_U247;
  assign new_P2_R1131_U249 = ~new_P2_U3422 | ~new_P2_R1131_U56;
  assign new_P2_R1131_U250 = ~new_P2_R1131_U62;
  assign new_P2_R1131_U251 = ~new_P2_U3425 | ~new_P2_R1131_U55;
  assign new_P2_R1131_U252 = ~new_P2_U3071 | ~new_P2_R1131_U61;
  assign new_P2_R1131_U253 = ~new_P2_U3428 | ~new_P2_R1131_U64;
  assign new_P2_R1131_U254 = ~new_P2_R1131_U253 | ~new_P2_R1131_U183;
  assign new_P2_R1131_U255 = ~new_P2_U3079 | ~new_P2_R1131_U63;
  assign new_P2_R1131_U256 = ~new_P2_R1131_U182;
  assign new_P2_R1131_U257 = ~new_P2_U3437 | ~new_P2_R1131_U68;
  assign new_P2_R1131_U258 = ~new_P2_U3072 | ~new_P2_R1131_U65;
  assign new_P2_R1131_U259 = ~new_P2_U3073 | ~new_P2_R1131_U66;
  assign new_P2_R1131_U260 = ~new_P2_R1131_U199 | ~new_P2_R1131_U8;
  assign new_P2_R1131_U261 = ~new_P2_R1131_U9 | ~new_P2_R1131_U260;
  assign new_P2_R1131_U262 = ~new_P2_U3431 | ~new_P2_R1131_U70;
  assign new_P2_R1131_U263 = ~new_P2_U3437 | ~new_P2_R1131_U68;
  assign new_P2_R1131_U264 = ~new_P2_R1131_U132 | ~new_P2_R1131_U182;
  assign new_P2_R1131_U265 = ~new_P2_R1131_U263 | ~new_P2_R1131_U261;
  assign new_P2_R1131_U266 = ~new_P2_R1131_U179;
  assign new_P2_R1131_U267 = ~new_P2_U3440 | ~new_P2_R1131_U73;
  assign new_P2_R1131_U268 = ~new_P2_R1131_U267 | ~new_P2_R1131_U179;
  assign new_P2_R1131_U269 = ~new_P2_U3068 | ~new_P2_R1131_U72;
  assign new_P2_R1131_U270 = ~new_P2_R1131_U178;
  assign new_P2_R1131_U271 = ~new_P2_U3081 | ~new_P2_R1131_U178;
  assign new_P2_R1131_U272 = ~new_P2_R1131_U176;
  assign new_P2_R1131_U273 = ~new_P2_U3445 | ~new_P2_R1131_U76;
  assign new_P2_R1131_U274 = ~new_P2_R1131_U273 | ~new_P2_R1131_U176;
  assign new_P2_R1131_U275 = ~new_P2_U3080 | ~new_P2_R1131_U75;
  assign new_P2_R1131_U276 = ~new_P2_R1131_U173;
  assign new_P2_R1131_U277 = ~new_P2_U3903 | ~new_P2_R1131_U78;
  assign new_P2_R1131_U278 = ~new_P2_R1131_U277 | ~new_P2_R1131_U173;
  assign new_P2_R1131_U279 = ~new_P2_U3075 | ~new_P2_R1131_U77;
  assign new_P2_R1131_U280 = ~new_P2_R1131_U172;
  assign new_P2_R1131_U281 = ~new_P2_U3900 | ~new_P2_R1131_U82;
  assign new_P2_R1131_U282 = ~new_P2_U3065 | ~new_P2_R1131_U79;
  assign new_P2_R1131_U283 = ~new_P2_U3060 | ~new_P2_R1131_U80;
  assign new_P2_R1131_U284 = ~new_P2_R1131_U200 | ~new_P2_R1131_U10;
  assign new_P2_R1131_U285 = ~new_P2_R1131_U11 | ~new_P2_R1131_U284;
  assign new_P2_R1131_U286 = ~new_P2_U3902 | ~new_P2_R1131_U84;
  assign new_P2_R1131_U287 = ~new_P2_U3900 | ~new_P2_R1131_U82;
  assign new_P2_R1131_U288 = ~new_P2_R1131_U133 | ~new_P2_R1131_U172;
  assign new_P2_R1131_U289 = ~new_P2_R1131_U287 | ~new_P2_R1131_U285;
  assign new_P2_R1131_U290 = ~new_P2_R1131_U169;
  assign new_P2_R1131_U291 = ~new_P2_U3899 | ~new_P2_R1131_U87;
  assign new_P2_R1131_U292 = ~new_P2_R1131_U291 | ~new_P2_R1131_U169;
  assign new_P2_R1131_U293 = ~new_P2_U3064 | ~new_P2_R1131_U86;
  assign new_P2_R1131_U294 = ~new_P2_R1131_U168;
  assign new_P2_R1131_U295 = ~new_P2_U3898 | ~new_P2_R1131_U89;
  assign new_P2_R1131_U296 = ~new_P2_R1131_U295 | ~new_P2_R1131_U168;
  assign new_P2_R1131_U297 = ~new_P2_U3057 | ~new_P2_R1131_U88;
  assign new_P2_R1131_U298 = ~new_P2_R1131_U93;
  assign new_P2_R1131_U299 = ~new_P2_U3896 | ~new_P2_R1131_U54;
  assign new_P2_R1131_U300 = ~new_P2_R1131_U54 | ~new_P2_R1131_U53;
  assign new_P2_R1131_U301 = ~new_P2_R1131_U300 | ~new_P2_R1131_U91;
  assign new_P2_R1131_U302 = ~new_P2_U3052 | ~new_P2_R1131_U189;
  assign new_P2_R1131_U303 = ~new_P2_U3895 | ~new_P2_R1131_U92;
  assign new_P2_R1131_U304 = ~new_P2_U3053 | ~new_P2_R1131_U51;
  assign new_P2_R1131_U305 = ~new_P2_R1131_U140 | ~new_P2_R1131_U355;
  assign new_P2_R1131_U306 = ~new_P2_R1131_U53 | ~new_P2_R1131_U195;
  assign new_P2_R1131_U307 = ~new_P2_R1131_U286 | ~new_P2_R1131_U172;
  assign new_P2_R1131_U308 = ~new_P2_R1131_U94;
  assign new_P2_R1131_U309 = ~new_P2_U3060 | ~new_P2_R1131_U80;
  assign new_P2_R1131_U310 = ~new_P2_R1131_U308 | ~new_P2_R1131_U309;
  assign new_P2_R1131_U311 = ~new_P2_R1131_U144 | ~new_P2_R1131_U310;
  assign new_P2_R1131_U312 = ~new_P2_R1131_U94 | ~new_P2_R1131_U194;
  assign new_P2_R1131_U313 = ~new_P2_U3900 | ~new_P2_R1131_U82;
  assign new_P2_R1131_U314 = ~new_P2_R1131_U143 | ~new_P2_R1131_U312;
  assign new_P2_R1131_U315 = ~new_P2_U3060 | ~new_P2_R1131_U80;
  assign new_P2_R1131_U316 = ~new_P2_R1131_U194 | ~new_P2_R1131_U315;
  assign new_P2_R1131_U317 = ~new_P2_R1131_U286 | ~new_P2_R1131_U85;
  assign new_P2_R1131_U318 = ~new_P2_R1131_U262 | ~new_P2_R1131_U182;
  assign new_P2_R1131_U319 = ~new_P2_R1131_U95;
  assign new_P2_R1131_U320 = ~new_P2_U3073 | ~new_P2_R1131_U66;
  assign new_P2_R1131_U321 = ~new_P2_R1131_U319 | ~new_P2_R1131_U320;
  assign new_P2_R1131_U322 = ~new_P2_R1131_U151 | ~new_P2_R1131_U321;
  assign new_P2_R1131_U323 = ~new_P2_R1131_U95 | ~new_P2_R1131_U193;
  assign new_P2_R1131_U324 = ~new_P2_U3437 | ~new_P2_R1131_U68;
  assign new_P2_R1131_U325 = ~new_P2_R1131_U150 | ~new_P2_R1131_U323;
  assign new_P2_R1131_U326 = ~new_P2_U3073 | ~new_P2_R1131_U66;
  assign new_P2_R1131_U327 = ~new_P2_R1131_U193 | ~new_P2_R1131_U326;
  assign new_P2_R1131_U328 = ~new_P2_R1131_U262 | ~new_P2_R1131_U71;
  assign new_P2_R1131_U329 = ~new_P2_U3061 | ~new_P2_R1131_U58;
  assign new_P2_R1131_U330 = ~new_P2_R1131_U350 | ~new_P2_R1131_U329;
  assign new_P2_R1131_U331 = ~new_P2_R1131_U155 | ~new_P2_R1131_U330;
  assign new_P2_R1131_U332 = ~new_P2_R1131_U96 | ~new_P2_R1131_U192;
  assign new_P2_R1131_U333 = ~new_P2_U3422 | ~new_P2_R1131_U56;
  assign new_P2_R1131_U334 = ~new_P2_R1131_U154 | ~new_P2_R1131_U332;
  assign new_P2_R1131_U335 = ~new_P2_U3061 | ~new_P2_R1131_U58;
  assign new_P2_R1131_U336 = ~new_P2_R1131_U192 | ~new_P2_R1131_U335;
  assign new_P2_R1131_U337 = ~new_P2_U3076 | ~new_P2_R1131_U38;
  assign new_P2_R1131_U338 = ~new_P2_U3077 | ~new_P2_R1131_U174;
  assign new_P2_R1131_U339 = ~new_P2_U3081 | ~new_P2_R1131_U177;
  assign new_P2_R1131_U340 = ~new_P2_R1131_U33 | ~new_P2_R1131_U221;
  assign new_P2_R1131_U341 = ~new_P2_R1131_U121 | ~new_P2_R1131_U161;
  assign new_P2_R1131_U342 = ~new_P2_R1131_U218 | ~new_P2_R1131_U14;
  assign new_P2_R1131_U343 = ~new_P2_R1131_U250 | ~new_P2_R1131_U251;
  assign new_P2_R1131_U344 = ~new_P2_R1131_U119 | ~new_P2_R1131_U50;
  assign new_P2_R1131_U345 = ~new_P2_R1131_U161;
  assign new_P2_R1131_U346 = ~new_P2_R1131_U196 | ~new_P2_R1131_U50;
  assign new_P2_R1131_U347 = ~new_P2_R1131_U128 | ~new_P2_R1131_U346;
  assign new_P2_R1131_U348 = ~new_P2_R1131_U205 | ~new_P2_R1131_U35;
  assign new_P2_R1131_U349 = ~new_P2_R1131_U224 | ~new_P2_R1131_U157;
  assign new_P2_R1131_U350 = ~new_P2_R1131_U96;
  assign new_P2_R1131_U351 = ~new_P2_R1131_U15 | ~new_P2_R1131_U157;
  assign new_P2_R1131_U352 = ~new_P2_R1131_U184;
  assign new_P2_R1131_U353 = ~new_P2_R1131_U130 | ~new_P2_R1131_U157;
  assign new_P2_R1131_U354 = ~new_P2_R1131_U183;
  assign new_P2_R1131_U355 = ~new_P2_R1131_U298 | ~new_P2_R1131_U53;
  assign new_P2_R1131_U356 = ~new_P2_R1131_U195 | ~new_P2_R1131_U93;
  assign new_P2_R1131_U357 = ~new_P2_R1131_U139 | ~new_P2_R1131_U356;
  assign new_P2_R1131_U358 = ~new_P2_R1131_U12 | ~new_P2_R1131_U93;
  assign new_P2_R1131_U359 = ~new_P2_R1131_U136 | ~new_P2_R1131_U358;
  assign new_P2_R1131_U360 = ~new_P2_R1131_U12 | ~new_P2_R1131_U93;
  assign new_P2_R1131_U361 = ~new_P2_R1131_U166;
  assign new_P2_R1131_U362 = ~new_P2_U3416 | ~new_P2_R1131_U47;
  assign new_P2_R1131_U363 = ~new_P2_U3082 | ~new_P2_R1131_U46;
  assign new_P2_R1131_U364 = ~new_P2_R1131_U225 | ~new_P2_R1131_U157;
  assign new_P2_R1131_U365 = ~new_P2_R1131_U223 | ~new_P2_R1131_U156;
  assign new_P2_R1131_U366 = ~new_P2_U3413 | ~new_P2_R1131_U28;
  assign new_P2_R1131_U367 = ~new_P2_U3083 | ~new_P2_R1131_U33;
  assign new_P2_R1131_U368 = ~new_P2_U3413 | ~new_P2_R1131_U28;
  assign new_P2_R1131_U369 = ~new_P2_U3083 | ~new_P2_R1131_U33;
  assign new_P2_R1131_U370 = ~new_P2_R1131_U369 | ~new_P2_R1131_U368;
  assign new_P2_R1131_U371 = ~new_P2_U3410 | ~new_P2_R1131_U26;
  assign new_P2_R1131_U372 = ~new_P2_U3069 | ~new_P2_R1131_U32;
  assign new_P2_R1131_U373 = ~new_P2_R1131_U230 | ~new_P2_R1131_U48;
  assign new_P2_R1131_U374 = ~new_P2_R1131_U158 | ~new_P2_R1131_U219;
  assign new_P2_R1131_U375 = ~new_P2_U3407 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U376 = ~new_P2_U3070 | ~new_P2_R1131_U30;
  assign new_P2_R1131_U377 = ~new_P2_R1131_U376 | ~new_P2_R1131_U375;
  assign new_P2_R1131_U378 = ~new_P2_U3404 | ~new_P2_R1131_U42;
  assign new_P2_R1131_U379 = ~new_P2_U3066 | ~new_P2_R1131_U29;
  assign new_P2_R1131_U380 = ~new_P2_R1131_U240 | ~new_P2_R1131_U49;
  assign new_P2_R1131_U381 = ~new_P2_R1131_U159 | ~new_P2_R1131_U232;
  assign new_P2_R1131_U382 = ~new_P2_U3401 | ~new_P2_R1131_U43;
  assign new_P2_R1131_U383 = ~new_P2_U3059 | ~new_P2_R1131_U31;
  assign new_P2_R1131_U384 = ~new_P2_R1131_U161 | ~new_P2_R1131_U241;
  assign new_P2_R1131_U385 = ~new_P2_R1131_U345 | ~new_P2_R1131_U160;
  assign new_P2_R1131_U386 = ~new_P2_U3398 | ~new_P2_R1131_U36;
  assign new_P2_R1131_U387 = ~new_P2_U3063 | ~new_P2_R1131_U40;
  assign new_P2_R1131_U388 = ~new_P2_U3398 | ~new_P2_R1131_U36;
  assign new_P2_R1131_U389 = ~new_P2_U3063 | ~new_P2_R1131_U40;
  assign new_P2_R1131_U390 = ~new_P2_R1131_U389 | ~new_P2_R1131_U388;
  assign new_P2_R1131_U391 = ~new_P2_U3395 | ~new_P2_R1131_U34;
  assign new_P2_R1131_U392 = ~new_P2_U3067 | ~new_P2_R1131_U37;
  assign new_P2_R1131_U393 = ~new_P2_R1131_U243 | ~new_P2_R1131_U50;
  assign new_P2_R1131_U394 = ~new_P2_R1131_U162 | ~new_P2_R1131_U205;
  assign new_P2_R1131_U395 = ~new_P2_U3904 | ~new_P2_R1131_U164;
  assign new_P2_R1131_U396 = ~new_P2_U3054 | ~new_P2_R1131_U163;
  assign new_P2_R1131_U397 = ~new_P2_R1131_U396 | ~new_P2_R1131_U395;
  assign new_P2_R1131_U398 = ~new_P2_U3904 | ~new_P2_R1131_U164;
  assign new_P2_R1131_U399 = ~new_P2_U3054 | ~new_P2_R1131_U163;
  assign new_P2_R1131_U400 = ~new_P2_R1131_U51 | ~new_P2_U3053 | ~new_P2_R1131_U397;
  assign new_P2_R1131_U401 = ~new_P2_U3895 | ~new_P2_R1131_U16 | ~new_P2_R1131_U92;
  assign new_P2_R1131_U402 = ~new_P2_U3895 | ~new_P2_R1131_U92;
  assign new_P2_R1131_U403 = ~new_P2_U3053 | ~new_P2_R1131_U51;
  assign new_P2_R1131_U404 = ~new_P2_R1131_U138;
  assign new_P2_R1131_U405 = ~new_P2_R1131_U361 | ~new_P2_R1131_U404;
  assign new_P2_R1131_U406 = ~new_P2_R1131_U138 | ~new_P2_R1131_U166;
  assign new_P2_R1131_U407 = ~new_P2_U3896 | ~new_P2_R1131_U54;
  assign new_P2_R1131_U408 = ~new_P2_U3052 | ~new_P2_R1131_U91;
  assign new_P2_R1131_U409 = ~new_P2_U3896 | ~new_P2_R1131_U54;
  assign new_P2_R1131_U410 = ~new_P2_U3052 | ~new_P2_R1131_U91;
  assign new_P2_R1131_U411 = ~new_P2_R1131_U410 | ~new_P2_R1131_U409;
  assign new_P2_R1131_U412 = ~new_P2_U3897 | ~new_P2_R1131_U52;
  assign new_P2_R1131_U413 = ~new_P2_U3056 | ~new_P2_R1131_U90;
  assign new_P2_R1131_U414 = ~new_P2_R1131_U306 | ~new_P2_R1131_U93;
  assign new_P2_R1131_U415 = ~new_P2_R1131_U167 | ~new_P2_R1131_U298;
  assign new_P2_R1131_U416 = ~new_P2_U3898 | ~new_P2_R1131_U89;
  assign new_P2_R1131_U417 = ~new_P2_U3057 | ~new_P2_R1131_U88;
  assign new_P2_R1131_U418 = ~new_P2_R1131_U141;
  assign new_P2_R1131_U419 = ~new_P2_R1131_U294 | ~new_P2_R1131_U418;
  assign new_P2_R1131_U420 = ~new_P2_R1131_U141 | ~new_P2_R1131_U168;
  assign new_P2_R1131_U421 = ~new_P2_U3899 | ~new_P2_R1131_U87;
  assign new_P2_R1131_U422 = ~new_P2_U3064 | ~new_P2_R1131_U86;
  assign new_P2_R1131_U423 = ~new_P2_R1131_U142;
  assign new_P2_R1131_U424 = ~new_P2_R1131_U290 | ~new_P2_R1131_U423;
  assign new_P2_R1131_U425 = ~new_P2_R1131_U142 | ~new_P2_R1131_U169;
  assign new_P2_R1131_U426 = ~new_P2_U3900 | ~new_P2_R1131_U82;
  assign new_P2_R1131_U427 = ~new_P2_U3065 | ~new_P2_R1131_U79;
  assign new_P2_R1131_U428 = ~new_P2_R1131_U427 | ~new_P2_R1131_U426;
  assign new_P2_R1131_U429 = ~new_P2_U3901 | ~new_P2_R1131_U83;
  assign new_P2_R1131_U430 = ~new_P2_U3060 | ~new_P2_R1131_U80;
  assign new_P2_R1131_U431 = ~new_P2_R1131_U316 | ~new_P2_R1131_U94;
  assign new_P2_R1131_U432 = ~new_P2_R1131_U170 | ~new_P2_R1131_U308;
  assign new_P2_R1131_U433 = ~new_P2_U3902 | ~new_P2_R1131_U84;
  assign new_P2_R1131_U434 = ~new_P2_U3074 | ~new_P2_R1131_U81;
  assign new_P2_R1131_U435 = ~new_P2_R1131_U317 | ~new_P2_R1131_U172;
  assign new_P2_R1131_U436 = ~new_P2_R1131_U280 | ~new_P2_R1131_U171;
  assign new_P2_R1131_U437 = ~new_P2_U3903 | ~new_P2_R1131_U78;
  assign new_P2_R1131_U438 = ~new_P2_U3075 | ~new_P2_R1131_U77;
  assign new_P2_R1131_U439 = ~new_P2_R1131_U145;
  assign new_P2_R1131_U440 = ~new_P2_R1131_U276 | ~new_P2_R1131_U439;
  assign new_P2_R1131_U441 = ~new_P2_R1131_U145 | ~new_P2_R1131_U173;
  assign new_P2_R1131_U442 = ~new_P2_U3392 | ~new_P2_R1131_U39;
  assign new_P2_R1131_U443 = ~new_P2_U3077 | ~new_P2_R1131_U174;
  assign new_P2_R1131_U444 = ~new_P2_R1131_U146;
  assign new_P2_R1131_U445 = ~new_P2_R1131_U203 | ~new_P2_R1131_U444;
  assign new_P2_R1131_U446 = ~new_P2_R1131_U146 | ~new_P2_R1131_U175;
  assign new_P2_R1131_U447 = ~new_P2_U3445 | ~new_P2_R1131_U76;
  assign new_P2_R1131_U448 = ~new_P2_U3080 | ~new_P2_R1131_U75;
  assign new_P2_R1131_U449 = ~new_P2_R1131_U147;
  assign new_P2_R1131_U450 = ~new_P2_R1131_U272 | ~new_P2_R1131_U449;
  assign new_P2_R1131_U451 = ~new_P2_R1131_U147 | ~new_P2_R1131_U176;
  assign new_P2_R1131_U452 = ~new_P2_U3443 | ~new_P2_R1131_U74;
  assign new_P2_R1131_U453 = ~new_P2_U3081 | ~new_P2_R1131_U177;
  assign new_P2_R1131_U454 = ~new_P2_R1131_U148;
  assign new_P2_R1131_U455 = ~new_P2_R1131_U270 | ~new_P2_R1131_U454;
  assign new_P2_R1131_U456 = ~new_P2_R1131_U148 | ~new_P2_R1131_U178;
  assign new_P2_R1131_U457 = ~new_P2_U3440 | ~new_P2_R1131_U73;
  assign new_P2_R1131_U458 = ~new_P2_U3068 | ~new_P2_R1131_U72;
  assign new_P2_R1131_U459 = ~new_P2_R1131_U149;
  assign new_P2_R1131_U460 = ~new_P2_R1131_U266 | ~new_P2_R1131_U459;
  assign new_P2_R1131_U461 = ~new_P2_R1131_U149 | ~new_P2_R1131_U179;
  assign new_P2_R1131_U462 = ~new_P2_U3437 | ~new_P2_R1131_U68;
  assign new_P2_R1131_U463 = ~new_P2_U3072 | ~new_P2_R1131_U65;
  assign new_P2_R1131_U464 = ~new_P2_R1131_U463 | ~new_P2_R1131_U462;
  assign new_P2_R1131_U465 = ~new_P2_U3434 | ~new_P2_R1131_U69;
  assign new_P2_R1131_U466 = ~new_P2_U3073 | ~new_P2_R1131_U66;
  assign new_P2_R1131_U467 = ~new_P2_R1131_U327 | ~new_P2_R1131_U95;
  assign new_P2_R1131_U468 = ~new_P2_R1131_U180 | ~new_P2_R1131_U319;
  assign new_P2_R1131_U469 = ~new_P2_U3431 | ~new_P2_R1131_U70;
  assign new_P2_R1131_U470 = ~new_P2_U3078 | ~new_P2_R1131_U67;
  assign new_P2_R1131_U471 = ~new_P2_R1131_U328 | ~new_P2_R1131_U182;
  assign new_P2_R1131_U472 = ~new_P2_R1131_U256 | ~new_P2_R1131_U181;
  assign new_P2_R1131_U473 = ~new_P2_U3428 | ~new_P2_R1131_U64;
  assign new_P2_R1131_U474 = ~new_P2_U3079 | ~new_P2_R1131_U63;
  assign new_P2_R1131_U475 = ~new_P2_R1131_U152;
  assign new_P2_R1131_U476 = ~new_P2_R1131_U354 | ~new_P2_R1131_U475;
  assign new_P2_R1131_U477 = ~new_P2_R1131_U152 | ~new_P2_R1131_U183;
  assign new_P2_R1131_U478 = ~new_P2_U3425 | ~new_P2_R1131_U55;
  assign new_P2_R1131_U479 = ~new_P2_U3071 | ~new_P2_R1131_U61;
  assign new_P2_R1131_U480 = ~new_P2_R1131_U153;
  assign new_P2_R1131_U481 = ~new_P2_R1131_U352 | ~new_P2_R1131_U480;
  assign new_P2_R1131_U482 = ~new_P2_R1131_U153 | ~new_P2_R1131_U184;
  assign new_P2_R1131_U483 = ~new_P2_U3422 | ~new_P2_R1131_U56;
  assign new_P2_R1131_U484 = ~new_P2_U3062 | ~new_P2_R1131_U60;
  assign new_P2_R1131_U485 = ~new_P2_R1131_U484 | ~new_P2_R1131_U483;
  assign new_P2_R1131_U486 = ~new_P2_U3419 | ~new_P2_R1131_U57;
  assign new_P2_R1131_U487 = ~new_P2_U3061 | ~new_P2_R1131_U58;
  assign new_P2_R1131_U488 = ~new_P2_R1131_U96 | ~new_P2_R1131_U336;
  assign new_P2_R1131_U489 = ~new_P2_R1131_U185 | ~new_P2_R1131_U350;
  assign new_P2_R1054_U6 = new_P2_R1054_U102 & new_P2_R1054_U118;
  assign new_P2_R1054_U7 = new_P2_R1054_U120 & new_P2_R1054_U119;
  assign new_P2_R1054_U8 = new_P2_R1054_U99 & new_P2_R1054_U157;
  assign new_P2_R1054_U9 = new_P2_R1054_U159 & new_P2_R1054_U158;
  assign new_P2_R1054_U10 = new_P2_R1054_U100 & new_P2_R1054_U174;
  assign new_P2_R1054_U11 = new_P2_R1054_U176 & new_P2_R1054_U175;
  assign new_P2_R1054_U12 = ~new_P2_R1054_U207 | ~new_P2_R1054_U210;
  assign new_P2_R1054_U13 = ~new_P2_R1054_U196 | ~new_P2_R1054_U199;
  assign new_P2_R1054_U14 = ~new_P2_R1054_U153 | ~new_P2_R1054_U155;
  assign new_P2_R1054_U15 = ~new_P2_R1054_U145 | ~new_P2_R1054_U148;
  assign new_P2_R1054_U16 = ~new_P2_R1054_U137 | ~new_P2_R1054_U139;
  assign new_P2_R1054_U17 = ~new_P2_R1054_U21 | ~new_P2_R1054_U213;
  assign new_P2_R1054_U18 = ~new_P2_U3409;
  assign new_P2_R1054_U19 = ~new_P2_U3394;
  assign new_P2_R1054_U20 = ~new_P2_U3386;
  assign new_P2_R1054_U21 = ~new_P2_U3386 | ~new_P2_R1054_U65;
  assign new_P2_R1054_U22 = ~new_P2_U3573;
  assign new_P2_R1054_U23 = ~new_P2_U3397;
  assign new_P2_R1054_U24 = ~new_P2_U3562;
  assign new_P2_R1054_U25 = ~new_P2_U3562 | ~new_P2_R1054_U19;
  assign new_P2_R1054_U26 = ~new_P2_U3561;
  assign new_P2_R1054_U27 = ~new_P2_U3406;
  assign new_P2_R1054_U28 = ~new_P2_U3403;
  assign new_P2_R1054_U29 = ~new_P2_U3400;
  assign new_P2_R1054_U30 = ~new_P2_U3558;
  assign new_P2_R1054_U31 = ~new_P2_U3559;
  assign new_P2_R1054_U32 = ~new_P2_U3560;
  assign new_P2_R1054_U33 = ~new_P2_U3560 | ~new_P2_R1054_U29;
  assign new_P2_R1054_U34 = ~new_P2_U3412;
  assign new_P2_R1054_U35 = ~new_P2_U3557;
  assign new_P2_R1054_U36 = ~new_P2_U3557 | ~new_P2_R1054_U18;
  assign new_P2_R1054_U37 = ~new_P2_U3556;
  assign new_P2_R1054_U38 = ~new_P2_U3415;
  assign new_P2_R1054_U39 = ~new_P2_U3555;
  assign new_P2_R1054_U40 = ~new_P2_R1054_U126 | ~new_P2_R1054_U125;
  assign new_P2_R1054_U41 = ~new_P2_R1054_U33 | ~new_P2_R1054_U141;
  assign new_P2_R1054_U42 = ~new_P2_R1054_U110 | ~new_P2_R1054_U109;
  assign new_P2_R1054_U43 = ~new_P2_U3421;
  assign new_P2_R1054_U44 = ~new_P2_U3418;
  assign new_P2_R1054_U45 = ~new_P2_U3571;
  assign new_P2_R1054_U46 = ~new_P2_U3572;
  assign new_P2_R1054_U47 = ~new_P2_U3555 | ~new_P2_R1054_U38;
  assign new_P2_R1054_U48 = ~new_P2_U3424;
  assign new_P2_R1054_U49 = ~new_P2_U3570;
  assign new_P2_R1054_U50 = ~new_P2_U3427;
  assign new_P2_R1054_U51 = ~new_P2_U3569;
  assign new_P2_R1054_U52 = ~new_P2_U3436;
  assign new_P2_R1054_U53 = ~new_P2_U3433;
  assign new_P2_R1054_U54 = ~new_P2_U3430;
  assign new_P2_R1054_U55 = ~new_P2_U3566;
  assign new_P2_R1054_U56 = ~new_P2_U3567;
  assign new_P2_R1054_U57 = ~new_P2_U3568;
  assign new_P2_R1054_U58 = ~new_P2_U3568 | ~new_P2_R1054_U54;
  assign new_P2_R1054_U59 = ~new_P2_U3439;
  assign new_P2_R1054_U60 = ~new_P2_U3565;
  assign new_P2_R1054_U61 = ~new_P2_R1054_U186 | ~new_P2_R1054_U185;
  assign new_P2_R1054_U62 = ~new_P2_U3564;
  assign new_P2_R1054_U63 = ~new_P2_R1054_U58 | ~new_P2_R1054_U192;
  assign new_P2_R1054_U64 = ~new_P2_R1054_U47 | ~new_P2_R1054_U203;
  assign new_P2_R1054_U65 = ~new_P2_U3574;
  assign new_P2_R1054_U66 = ~new_P2_R1054_U251 | ~new_P2_R1054_U250;
  assign new_P2_R1054_U67 = ~new_P2_R1054_U256 | ~new_P2_R1054_U255;
  assign new_P2_R1054_U68 = ~new_P2_R1054_U261 | ~new_P2_R1054_U260;
  assign new_P2_R1054_U69 = ~new_P2_R1054_U266 | ~new_P2_R1054_U265;
  assign new_P2_R1054_U70 = ~new_P2_R1054_U282 | ~new_P2_R1054_U281;
  assign new_P2_R1054_U71 = ~new_P2_R1054_U287 | ~new_P2_R1054_U286;
  assign new_P2_R1054_U72 = ~new_P2_R1054_U217 | ~new_P2_R1054_U216;
  assign new_P2_R1054_U73 = ~new_P2_R1054_U226 | ~new_P2_R1054_U225;
  assign new_P2_R1054_U74 = ~new_P2_R1054_U233 | ~new_P2_R1054_U232;
  assign new_P2_R1054_U75 = ~new_P2_R1054_U237 | ~new_P2_R1054_U236;
  assign new_P2_R1054_U76 = ~new_P2_R1054_U246 | ~new_P2_R1054_U245;
  assign new_P2_R1054_U77 = ~new_P2_R1054_U273 | ~new_P2_R1054_U272;
  assign new_P2_R1054_U78 = ~new_P2_R1054_U277 | ~new_P2_R1054_U276;
  assign new_P2_R1054_U79 = ~new_P2_R1054_U294 | ~new_P2_R1054_U293;
  assign new_P2_R1054_U80 = ~new_P2_R1054_U248 | ~new_P2_R1054_U247;
  assign new_P2_R1054_U81 = ~new_P2_R1054_U253 | ~new_P2_R1054_U252;
  assign new_P2_R1054_U82 = ~new_P2_R1054_U258 | ~new_P2_R1054_U257;
  assign new_P2_R1054_U83 = ~new_P2_R1054_U263 | ~new_P2_R1054_U262;
  assign new_P2_R1054_U84 = ~new_P2_R1054_U279 | ~new_P2_R1054_U278;
  assign new_P2_R1054_U85 = ~new_P2_R1054_U284 | ~new_P2_R1054_U283;
  assign new_P2_R1054_U86 = ~new_P2_R1054_U129 | ~new_P2_R1054_U131 | ~new_P2_R1054_U132;
  assign new_P2_R1054_U87 = ~new_P2_R1054_U113 | ~new_P2_R1054_U115 | ~new_P2_R1054_U116;
  assign new_P2_R1054_U88 = ~new_P2_U3391;
  assign new_P2_R1054_U89 = ~new_P2_U3379;
  assign new_P2_R1054_U90 = ~new_P2_U3563;
  assign new_P2_R1054_U91 = ~new_P2_R1054_U190 | ~new_P2_R1054_U189;
  assign new_P2_R1054_U92 = ~new_P2_U3442;
  assign new_P2_R1054_U93 = ~new_P2_R1054_U182 | ~new_P2_R1054_U181;
  assign new_P2_R1054_U94 = ~new_P2_R1054_U172 | ~new_P2_R1054_U171;
  assign new_P2_R1054_U95 = ~new_P2_R1054_U168 | ~new_P2_R1054_U167;
  assign new_P2_R1054_U96 = ~new_P2_R1054_U164 | ~new_P2_R1054_U163;
  assign new_P2_R1054_U97 = ~new_P2_R1054_U25;
  assign new_P2_R1054_U98 = ~new_P2_R1054_U36;
  assign new_P2_R1054_U99 = ~new_P2_U3418 | ~new_P2_R1054_U46;
  assign new_P2_R1054_U100 = ~new_P2_U3433 | ~new_P2_R1054_U56;
  assign new_P2_R1054_U101 = ~new_P2_U3394 | ~new_P2_R1054_U24;
  assign new_P2_R1054_U102 = ~new_P2_U3403 | ~new_P2_R1054_U31;
  assign new_P2_R1054_U103 = ~new_P2_U3409 | ~new_P2_R1054_U35;
  assign new_P2_R1054_U104 = ~new_P2_R1054_U58;
  assign new_P2_R1054_U105 = ~new_P2_R1054_U33;
  assign new_P2_R1054_U106 = ~new_P2_R1054_U47;
  assign new_P2_R1054_U107 = ~new_P2_R1054_U21;
  assign new_P2_R1054_U108 = ~new_P2_R1054_U107 | ~new_P2_R1054_U22;
  assign new_P2_R1054_U109 = ~new_P2_R1054_U108 | ~new_P2_R1054_U88;
  assign new_P2_R1054_U110 = ~new_P2_U3573 | ~new_P2_R1054_U21;
  assign new_P2_R1054_U111 = ~new_P2_R1054_U42;
  assign new_P2_R1054_U112 = ~new_P2_U3397 | ~new_P2_R1054_U26;
  assign new_P2_R1054_U113 = ~new_P2_R1054_U42 | ~new_P2_R1054_U112 | ~new_P2_R1054_U101;
  assign new_P2_R1054_U114 = ~new_P2_R1054_U26 | ~new_P2_R1054_U25;
  assign new_P2_R1054_U115 = ~new_P2_R1054_U114 | ~new_P2_R1054_U23;
  assign new_P2_R1054_U116 = ~new_P2_U3561 | ~new_P2_R1054_U97;
  assign new_P2_R1054_U117 = ~new_P2_R1054_U87;
  assign new_P2_R1054_U118 = ~new_P2_U3406 | ~new_P2_R1054_U30;
  assign new_P2_R1054_U119 = ~new_P2_U3558 | ~new_P2_R1054_U27;
  assign new_P2_R1054_U120 = ~new_P2_U3559 | ~new_P2_R1054_U28;
  assign new_P2_R1054_U121 = ~new_P2_R1054_U105 | ~new_P2_R1054_U6;
  assign new_P2_R1054_U122 = ~new_P2_R1054_U7 | ~new_P2_R1054_U121;
  assign new_P2_R1054_U123 = ~new_P2_U3400 | ~new_P2_R1054_U32;
  assign new_P2_R1054_U124 = ~new_P2_U3406 | ~new_P2_R1054_U30;
  assign new_P2_R1054_U125 = ~new_P2_R1054_U87 | ~new_P2_R1054_U123 | ~new_P2_R1054_U6;
  assign new_P2_R1054_U126 = ~new_P2_R1054_U124 | ~new_P2_R1054_U122;
  assign new_P2_R1054_U127 = ~new_P2_R1054_U40;
  assign new_P2_R1054_U128 = ~new_P2_U3412 | ~new_P2_R1054_U37;
  assign new_P2_R1054_U129 = ~new_P2_R1054_U40 | ~new_P2_R1054_U128 | ~new_P2_R1054_U103;
  assign new_P2_R1054_U130 = ~new_P2_R1054_U37 | ~new_P2_R1054_U36;
  assign new_P2_R1054_U131 = ~new_P2_R1054_U130 | ~new_P2_R1054_U34;
  assign new_P2_R1054_U132 = ~new_P2_U3556 | ~new_P2_R1054_U98;
  assign new_P2_R1054_U133 = ~new_P2_R1054_U86;
  assign new_P2_R1054_U134 = ~new_P2_U3415 | ~new_P2_R1054_U39;
  assign new_P2_R1054_U135 = ~new_P2_R1054_U134 | ~new_P2_R1054_U47;
  assign new_P2_R1054_U136 = ~new_P2_R1054_U127 | ~new_P2_R1054_U36;
  assign new_P2_R1054_U137 = ~new_P2_R1054_U136 | ~new_P2_R1054_U222 | ~new_P2_R1054_U103;
  assign new_P2_R1054_U138 = ~new_P2_R1054_U40 | ~new_P2_R1054_U103;
  assign new_P2_R1054_U139 = ~new_P2_R1054_U138 | ~new_P2_R1054_U36 | ~new_P2_R1054_U219 | ~new_P2_R1054_U218;
  assign new_P2_R1054_U140 = ~new_P2_R1054_U36 | ~new_P2_R1054_U103;
  assign new_P2_R1054_U141 = ~new_P2_R1054_U123 | ~new_P2_R1054_U87;
  assign new_P2_R1054_U142 = ~new_P2_R1054_U41;
  assign new_P2_R1054_U143 = ~new_P2_U3559 | ~new_P2_R1054_U28;
  assign new_P2_R1054_U144 = ~new_P2_R1054_U142 | ~new_P2_R1054_U143;
  assign new_P2_R1054_U145 = ~new_P2_R1054_U144 | ~new_P2_R1054_U229 | ~new_P2_R1054_U102;
  assign new_P2_R1054_U146 = ~new_P2_R1054_U41 | ~new_P2_R1054_U102;
  assign new_P2_R1054_U147 = ~new_P2_U3406 | ~new_P2_R1054_U30;
  assign new_P2_R1054_U148 = ~new_P2_R1054_U146 | ~new_P2_R1054_U147 | ~new_P2_R1054_U7;
  assign new_P2_R1054_U149 = ~new_P2_U3559 | ~new_P2_R1054_U28;
  assign new_P2_R1054_U150 = ~new_P2_R1054_U102 | ~new_P2_R1054_U149;
  assign new_P2_R1054_U151 = ~new_P2_R1054_U123 | ~new_P2_R1054_U33;
  assign new_P2_R1054_U152 = ~new_P2_R1054_U111 | ~new_P2_R1054_U25;
  assign new_P2_R1054_U153 = ~new_P2_R1054_U152 | ~new_P2_R1054_U242 | ~new_P2_R1054_U101;
  assign new_P2_R1054_U154 = ~new_P2_R1054_U42 | ~new_P2_R1054_U101;
  assign new_P2_R1054_U155 = ~new_P2_R1054_U154 | ~new_P2_R1054_U25 | ~new_P2_R1054_U239 | ~new_P2_R1054_U238;
  assign new_P2_R1054_U156 = ~new_P2_R1054_U25 | ~new_P2_R1054_U101;
  assign new_P2_R1054_U157 = ~new_P2_U3421 | ~new_P2_R1054_U45;
  assign new_P2_R1054_U158 = ~new_P2_U3571 | ~new_P2_R1054_U43;
  assign new_P2_R1054_U159 = ~new_P2_U3572 | ~new_P2_R1054_U44;
  assign new_P2_R1054_U160 = ~new_P2_R1054_U106 | ~new_P2_R1054_U8;
  assign new_P2_R1054_U161 = ~new_P2_R1054_U9 | ~new_P2_R1054_U160;
  assign new_P2_R1054_U162 = ~new_P2_U3421 | ~new_P2_R1054_U45;
  assign new_P2_R1054_U163 = ~new_P2_R1054_U86 | ~new_P2_R1054_U134 | ~new_P2_R1054_U8;
  assign new_P2_R1054_U164 = ~new_P2_R1054_U162 | ~new_P2_R1054_U161;
  assign new_P2_R1054_U165 = ~new_P2_R1054_U96;
  assign new_P2_R1054_U166 = ~new_P2_U3424 | ~new_P2_R1054_U49;
  assign new_P2_R1054_U167 = ~new_P2_R1054_U166 | ~new_P2_R1054_U96;
  assign new_P2_R1054_U168 = ~new_P2_U3570 | ~new_P2_R1054_U48;
  assign new_P2_R1054_U169 = ~new_P2_R1054_U95;
  assign new_P2_R1054_U170 = ~new_P2_U3427 | ~new_P2_R1054_U51;
  assign new_P2_R1054_U171 = ~new_P2_R1054_U170 | ~new_P2_R1054_U95;
  assign new_P2_R1054_U172 = ~new_P2_U3569 | ~new_P2_R1054_U50;
  assign new_P2_R1054_U173 = ~new_P2_R1054_U94;
  assign new_P2_R1054_U174 = ~new_P2_U3436 | ~new_P2_R1054_U55;
  assign new_P2_R1054_U175 = ~new_P2_U3566 | ~new_P2_R1054_U52;
  assign new_P2_R1054_U176 = ~new_P2_U3567 | ~new_P2_R1054_U53;
  assign new_P2_R1054_U177 = ~new_P2_R1054_U104 | ~new_P2_R1054_U10;
  assign new_P2_R1054_U178 = ~new_P2_R1054_U11 | ~new_P2_R1054_U177;
  assign new_P2_R1054_U179 = ~new_P2_U3430 | ~new_P2_R1054_U57;
  assign new_P2_R1054_U180 = ~new_P2_U3436 | ~new_P2_R1054_U55;
  assign new_P2_R1054_U181 = ~new_P2_R1054_U94 | ~new_P2_R1054_U179 | ~new_P2_R1054_U10;
  assign new_P2_R1054_U182 = ~new_P2_R1054_U180 | ~new_P2_R1054_U178;
  assign new_P2_R1054_U183 = ~new_P2_R1054_U93;
  assign new_P2_R1054_U184 = ~new_P2_U3439 | ~new_P2_R1054_U60;
  assign new_P2_R1054_U185 = ~new_P2_R1054_U184 | ~new_P2_R1054_U93;
  assign new_P2_R1054_U186 = ~new_P2_U3565 | ~new_P2_R1054_U59;
  assign new_P2_R1054_U187 = ~new_P2_R1054_U61;
  assign new_P2_R1054_U188 = ~new_P2_R1054_U187 | ~new_P2_R1054_U62;
  assign new_P2_R1054_U189 = ~new_P2_R1054_U188 | ~new_P2_R1054_U92;
  assign new_P2_R1054_U190 = ~new_P2_U3564 | ~new_P2_R1054_U61;
  assign new_P2_R1054_U191 = ~new_P2_R1054_U91;
  assign new_P2_R1054_U192 = ~new_P2_R1054_U179 | ~new_P2_R1054_U94;
  assign new_P2_R1054_U193 = ~new_P2_R1054_U63;
  assign new_P2_R1054_U194 = ~new_P2_U3567 | ~new_P2_R1054_U53;
  assign new_P2_R1054_U195 = ~new_P2_R1054_U193 | ~new_P2_R1054_U194;
  assign new_P2_R1054_U196 = ~new_P2_R1054_U195 | ~new_P2_R1054_U269 | ~new_P2_R1054_U100;
  assign new_P2_R1054_U197 = ~new_P2_R1054_U63 | ~new_P2_R1054_U100;
  assign new_P2_R1054_U198 = ~new_P2_U3436 | ~new_P2_R1054_U55;
  assign new_P2_R1054_U199 = ~new_P2_R1054_U197 | ~new_P2_R1054_U198 | ~new_P2_R1054_U11;
  assign new_P2_R1054_U200 = ~new_P2_U3567 | ~new_P2_R1054_U53;
  assign new_P2_R1054_U201 = ~new_P2_R1054_U100 | ~new_P2_R1054_U200;
  assign new_P2_R1054_U202 = ~new_P2_R1054_U179 | ~new_P2_R1054_U58;
  assign new_P2_R1054_U203 = ~new_P2_R1054_U134 | ~new_P2_R1054_U86;
  assign new_P2_R1054_U204 = ~new_P2_R1054_U64;
  assign new_P2_R1054_U205 = ~new_P2_U3572 | ~new_P2_R1054_U44;
  assign new_P2_R1054_U206 = ~new_P2_R1054_U204 | ~new_P2_R1054_U205;
  assign new_P2_R1054_U207 = ~new_P2_R1054_U206 | ~new_P2_R1054_U290 | ~new_P2_R1054_U99;
  assign new_P2_R1054_U208 = ~new_P2_R1054_U64 | ~new_P2_R1054_U99;
  assign new_P2_R1054_U209 = ~new_P2_U3421 | ~new_P2_R1054_U45;
  assign new_P2_R1054_U210 = ~new_P2_R1054_U208 | ~new_P2_R1054_U209 | ~new_P2_R1054_U9;
  assign new_P2_R1054_U211 = ~new_P2_U3572 | ~new_P2_R1054_U44;
  assign new_P2_R1054_U212 = ~new_P2_R1054_U99 | ~new_P2_R1054_U211;
  assign new_P2_R1054_U213 = ~new_P2_U3574 | ~new_P2_R1054_U20;
  assign new_P2_R1054_U214 = ~new_P2_U3415 | ~new_P2_R1054_U39;
  assign new_P2_R1054_U215 = ~new_P2_U3555 | ~new_P2_R1054_U38;
  assign new_P2_R1054_U216 = ~new_P2_R1054_U135 | ~new_P2_R1054_U86;
  assign new_P2_R1054_U217 = ~new_P2_R1054_U133 | ~new_P2_R1054_U215 | ~new_P2_R1054_U214;
  assign new_P2_R1054_U218 = ~new_P2_U3412 | ~new_P2_R1054_U37;
  assign new_P2_R1054_U219 = ~new_P2_U3556 | ~new_P2_R1054_U34;
  assign new_P2_R1054_U220 = ~new_P2_U3412 | ~new_P2_R1054_U37;
  assign new_P2_R1054_U221 = ~new_P2_U3556 | ~new_P2_R1054_U34;
  assign new_P2_R1054_U222 = ~new_P2_R1054_U221 | ~new_P2_R1054_U220;
  assign new_P2_R1054_U223 = ~new_P2_U3409 | ~new_P2_R1054_U35;
  assign new_P2_R1054_U224 = ~new_P2_U3557 | ~new_P2_R1054_U18;
  assign new_P2_R1054_U225 = ~new_P2_R1054_U140 | ~new_P2_R1054_U40;
  assign new_P2_R1054_U226 = ~new_P2_R1054_U127 | ~new_P2_R1054_U224 | ~new_P2_R1054_U223;
  assign new_P2_R1054_U227 = ~new_P2_U3406 | ~new_P2_R1054_U30;
  assign new_P2_R1054_U228 = ~new_P2_U3558 | ~new_P2_R1054_U27;
  assign new_P2_R1054_U229 = ~new_P2_R1054_U228 | ~new_P2_R1054_U227;
  assign new_P2_R1054_U230 = ~new_P2_U3403 | ~new_P2_R1054_U31;
  assign new_P2_R1054_U231 = ~new_P2_U3559 | ~new_P2_R1054_U28;
  assign new_P2_R1054_U232 = ~new_P2_R1054_U150 | ~new_P2_R1054_U41;
  assign new_P2_R1054_U233 = ~new_P2_R1054_U142 | ~new_P2_R1054_U231 | ~new_P2_R1054_U230;
  assign new_P2_R1054_U234 = ~new_P2_U3400 | ~new_P2_R1054_U32;
  assign new_P2_R1054_U235 = ~new_P2_U3560 | ~new_P2_R1054_U29;
  assign new_P2_R1054_U236 = ~new_P2_R1054_U151 | ~new_P2_R1054_U87;
  assign new_P2_R1054_U237 = ~new_P2_R1054_U117 | ~new_P2_R1054_U235 | ~new_P2_R1054_U234;
  assign new_P2_R1054_U238 = ~new_P2_U3397 | ~new_P2_R1054_U26;
  assign new_P2_R1054_U239 = ~new_P2_U3561 | ~new_P2_R1054_U23;
  assign new_P2_R1054_U240 = ~new_P2_U3397 | ~new_P2_R1054_U26;
  assign new_P2_R1054_U241 = ~new_P2_U3561 | ~new_P2_R1054_U23;
  assign new_P2_R1054_U242 = ~new_P2_R1054_U241 | ~new_P2_R1054_U240;
  assign new_P2_R1054_U243 = ~new_P2_U3394 | ~new_P2_R1054_U24;
  assign new_P2_R1054_U244 = ~new_P2_U3562 | ~new_P2_R1054_U19;
  assign new_P2_R1054_U245 = ~new_P2_R1054_U156 | ~new_P2_R1054_U42;
  assign new_P2_R1054_U246 = ~new_P2_R1054_U111 | ~new_P2_R1054_U244 | ~new_P2_R1054_U243;
  assign new_P2_R1054_U247 = ~new_P2_U3391 | ~new_P2_R1054_U22;
  assign new_P2_R1054_U248 = ~new_P2_U3573 | ~new_P2_R1054_U88;
  assign new_P2_R1054_U249 = ~new_P2_R1054_U80;
  assign new_P2_R1054_U250 = ~new_P2_R1054_U249 | ~new_P2_R1054_U107;
  assign new_P2_R1054_U251 = ~new_P2_R1054_U80 | ~new_P2_R1054_U21;
  assign new_P2_R1054_U252 = ~new_P2_U3379 | ~new_P2_R1054_U90;
  assign new_P2_R1054_U253 = ~new_P2_U3563 | ~new_P2_R1054_U89;
  assign new_P2_R1054_U254 = ~new_P2_R1054_U81;
  assign new_P2_R1054_U255 = ~new_P2_R1054_U191 | ~new_P2_R1054_U254;
  assign new_P2_R1054_U256 = ~new_P2_R1054_U81 | ~new_P2_R1054_U91;
  assign new_P2_R1054_U257 = ~new_P2_U3442 | ~new_P2_R1054_U62;
  assign new_P2_R1054_U258 = ~new_P2_U3564 | ~new_P2_R1054_U92;
  assign new_P2_R1054_U259 = ~new_P2_R1054_U82;
  assign new_P2_R1054_U260 = ~new_P2_R1054_U259 | ~new_P2_R1054_U187;
  assign new_P2_R1054_U261 = ~new_P2_R1054_U82 | ~new_P2_R1054_U61;
  assign new_P2_R1054_U262 = ~new_P2_U3439 | ~new_P2_R1054_U60;
  assign new_P2_R1054_U263 = ~new_P2_U3565 | ~new_P2_R1054_U59;
  assign new_P2_R1054_U264 = ~new_P2_R1054_U83;
  assign new_P2_R1054_U265 = ~new_P2_R1054_U183 | ~new_P2_R1054_U264;
  assign new_P2_R1054_U266 = ~new_P2_R1054_U83 | ~new_P2_R1054_U93;
  assign new_P2_R1054_U267 = ~new_P2_U3436 | ~new_P2_R1054_U55;
  assign new_P2_R1054_U268 = ~new_P2_U3566 | ~new_P2_R1054_U52;
  assign new_P2_R1054_U269 = ~new_P2_R1054_U268 | ~new_P2_R1054_U267;
  assign new_P2_R1054_U270 = ~new_P2_U3433 | ~new_P2_R1054_U56;
  assign new_P2_R1054_U271 = ~new_P2_U3567 | ~new_P2_R1054_U53;
  assign new_P2_R1054_U272 = ~new_P2_R1054_U201 | ~new_P2_R1054_U63;
  assign new_P2_R1054_U273 = ~new_P2_R1054_U193 | ~new_P2_R1054_U271 | ~new_P2_R1054_U270;
  assign new_P2_R1054_U274 = ~new_P2_U3430 | ~new_P2_R1054_U57;
  assign new_P2_R1054_U275 = ~new_P2_U3568 | ~new_P2_R1054_U54;
  assign new_P2_R1054_U276 = ~new_P2_R1054_U202 | ~new_P2_R1054_U94;
  assign new_P2_R1054_U277 = ~new_P2_R1054_U173 | ~new_P2_R1054_U275 | ~new_P2_R1054_U274;
  assign new_P2_R1054_U278 = ~new_P2_U3427 | ~new_P2_R1054_U51;
  assign new_P2_R1054_U279 = ~new_P2_U3569 | ~new_P2_R1054_U50;
  assign new_P2_R1054_U280 = ~new_P2_R1054_U84;
  assign new_P2_R1054_U281 = ~new_P2_R1054_U169 | ~new_P2_R1054_U280;
  assign new_P2_R1054_U282 = ~new_P2_R1054_U84 | ~new_P2_R1054_U95;
  assign new_P2_R1054_U283 = ~new_P2_U3424 | ~new_P2_R1054_U49;
  assign new_P2_R1054_U284 = ~new_P2_U3570 | ~new_P2_R1054_U48;
  assign new_P2_R1054_U285 = ~new_P2_R1054_U85;
  assign new_P2_R1054_U286 = ~new_P2_R1054_U165 | ~new_P2_R1054_U285;
  assign new_P2_R1054_U287 = ~new_P2_R1054_U85 | ~new_P2_R1054_U96;
  assign new_P2_R1054_U288 = ~new_P2_U3421 | ~new_P2_R1054_U45;
  assign new_P2_R1054_U289 = ~new_P2_U3571 | ~new_P2_R1054_U43;
  assign new_P2_R1054_U290 = ~new_P2_R1054_U289 | ~new_P2_R1054_U288;
  assign new_P2_R1054_U291 = ~new_P2_U3418 | ~new_P2_R1054_U46;
  assign new_P2_R1054_U292 = ~new_P2_U3572 | ~new_P2_R1054_U44;
  assign new_P2_R1054_U293 = ~new_P2_R1054_U212 | ~new_P2_R1054_U64;
  assign new_P2_R1054_U294 = ~new_P2_R1054_U204 | ~new_P2_R1054_U292 | ~new_P2_R1054_U291;
  assign new_P2_R1161_U4 = new_P2_R1161_U179 & new_P2_R1161_U178;
  assign new_P2_R1161_U5 = new_P2_R1161_U197 & new_P2_R1161_U196;
  assign new_P2_R1161_U6 = new_P2_R1161_U237 & new_P2_R1161_U236;
  assign new_P2_R1161_U7 = new_P2_R1161_U246 & new_P2_R1161_U245;
  assign new_P2_R1161_U8 = new_P2_R1161_U264 & new_P2_R1161_U263;
  assign new_P2_R1161_U9 = new_P2_R1161_U272 & new_P2_R1161_U271;
  assign new_P2_R1161_U10 = new_P2_R1161_U351 & new_P2_R1161_U348;
  assign new_P2_R1161_U11 = new_P2_R1161_U344 & new_P2_R1161_U341;
  assign new_P2_R1161_U12 = new_P2_R1161_U335 & new_P2_R1161_U332;
  assign new_P2_R1161_U13 = new_P2_R1161_U326 & new_P2_R1161_U323;
  assign new_P2_R1161_U14 = new_P2_R1161_U320 & new_P2_R1161_U318;
  assign new_P2_R1161_U15 = new_P2_R1161_U313 & new_P2_R1161_U310;
  assign new_P2_R1161_U16 = new_P2_R1161_U235 & new_P2_R1161_U232;
  assign new_P2_R1161_U17 = new_P2_R1161_U227 & new_P2_R1161_U224;
  assign new_P2_R1161_U18 = new_P2_R1161_U213 & new_P2_R1161_U210;
  assign new_P2_R1161_U19 = ~new_P2_U3407;
  assign new_P2_R1161_U20 = ~new_P2_U3070;
  assign new_P2_R1161_U21 = ~new_P2_U3069;
  assign new_P2_R1161_U22 = ~new_P2_U3070 | ~new_P2_U3407;
  assign new_P2_R1161_U23 = ~new_P2_U3410;
  assign new_P2_R1161_U24 = ~new_P2_U3401;
  assign new_P2_R1161_U25 = ~new_P2_U3059;
  assign new_P2_R1161_U26 = ~new_P2_U3066;
  assign new_P2_R1161_U27 = ~new_P2_U3395;
  assign new_P2_R1161_U28 = ~new_P2_U3067;
  assign new_P2_R1161_U29 = ~new_P2_U3387;
  assign new_P2_R1161_U30 = ~new_P2_U3076;
  assign new_P2_R1161_U31 = ~new_P2_U3076 | ~new_P2_U3387;
  assign new_P2_R1161_U32 = ~new_P2_U3398;
  assign new_P2_R1161_U33 = ~new_P2_U3063;
  assign new_P2_R1161_U34 = ~new_P2_U3059 | ~new_P2_U3401;
  assign new_P2_R1161_U35 = ~new_P2_U3404;
  assign new_P2_R1161_U36 = ~new_P2_U3413;
  assign new_P2_R1161_U37 = ~new_P2_U3083;
  assign new_P2_R1161_U38 = ~new_P2_U3082;
  assign new_P2_R1161_U39 = ~new_P2_U3416;
  assign new_P2_R1161_U40 = ~new_P2_R1161_U65 | ~new_P2_R1161_U205;
  assign new_P2_R1161_U41 = ~new_P2_R1161_U117 | ~new_P2_R1161_U193;
  assign new_P2_R1161_U42 = ~new_P2_R1161_U182 | ~new_P2_R1161_U183;
  assign new_P2_R1161_U43 = ~new_P2_U3392 | ~new_P2_U3077;
  assign new_P2_R1161_U44 = ~new_P2_R1161_U122 | ~new_P2_R1161_U219;
  assign new_P2_R1161_U45 = ~new_P2_R1161_U216 | ~new_P2_R1161_U215;
  assign new_P2_R1161_U46 = ~new_P2_U3896;
  assign new_P2_R1161_U47 = ~new_P2_U3052;
  assign new_P2_R1161_U48 = ~new_P2_U3056;
  assign new_P2_R1161_U49 = ~new_P2_U3897;
  assign new_P2_R1161_U50 = ~new_P2_U3898;
  assign new_P2_R1161_U51 = ~new_P2_U3057;
  assign new_P2_R1161_U52 = ~new_P2_U3899;
  assign new_P2_R1161_U53 = ~new_P2_U3064;
  assign new_P2_R1161_U54 = ~new_P2_U3902;
  assign new_P2_R1161_U55 = ~new_P2_U3074;
  assign new_P2_R1161_U56 = ~new_P2_U3437;
  assign new_P2_R1161_U57 = ~new_P2_U3072;
  assign new_P2_R1161_U58 = ~new_P2_U3068;
  assign new_P2_R1161_U59 = ~new_P2_U3072 | ~new_P2_U3437;
  assign new_P2_R1161_U60 = ~new_P2_U3440;
  assign new_P2_R1161_U61 = ~new_P2_U3428;
  assign new_P2_R1161_U62 = ~new_P2_U3079;
  assign new_P2_R1161_U63 = ~new_P2_U3419;
  assign new_P2_R1161_U64 = ~new_P2_U3061;
  assign new_P2_R1161_U65 = ~new_P2_U3083 | ~new_P2_U3413;
  assign new_P2_R1161_U66 = ~new_P2_U3422;
  assign new_P2_R1161_U67 = ~new_P2_U3062;
  assign new_P2_R1161_U68 = ~new_P2_U3062 | ~new_P2_U3422;
  assign new_P2_R1161_U69 = ~new_P2_U3425;
  assign new_P2_R1161_U70 = ~new_P2_U3071;
  assign new_P2_R1161_U71 = ~new_P2_U3431;
  assign new_P2_R1161_U72 = ~new_P2_U3078;
  assign new_P2_R1161_U73 = ~new_P2_U3434;
  assign new_P2_R1161_U74 = ~new_P2_U3073;
  assign new_P2_R1161_U75 = ~new_P2_U3443;
  assign new_P2_R1161_U76 = ~new_P2_U3081;
  assign new_P2_R1161_U77 = ~new_P2_U3081 | ~new_P2_U3443;
  assign new_P2_R1161_U78 = ~new_P2_U3445;
  assign new_P2_R1161_U79 = ~new_P2_U3080;
  assign new_P2_R1161_U80 = ~new_P2_U3080 | ~new_P2_U3445;
  assign new_P2_R1161_U81 = ~new_P2_U3903;
  assign new_P2_R1161_U82 = ~new_P2_U3901;
  assign new_P2_R1161_U83 = ~new_P2_U3060;
  assign new_P2_R1161_U84 = ~new_P2_U3900;
  assign new_P2_R1161_U85 = ~new_P2_U3065;
  assign new_P2_R1161_U86 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1161_U87 = ~new_P2_U3053;
  assign new_P2_R1161_U88 = ~new_P2_U3895;
  assign new_P2_R1161_U89 = ~new_P2_R1161_U306 | ~new_P2_R1161_U176;
  assign new_P2_R1161_U90 = ~new_P2_U3075;
  assign new_P2_R1161_U91 = ~new_P2_R1161_U77 | ~new_P2_R1161_U315;
  assign new_P2_R1161_U92 = ~new_P2_R1161_U261 | ~new_P2_R1161_U260;
  assign new_P2_R1161_U93 = ~new_P2_R1161_U68 | ~new_P2_R1161_U337;
  assign new_P2_R1161_U94 = ~new_P2_R1161_U457 | ~new_P2_R1161_U456;
  assign new_P2_R1161_U95 = ~new_P2_R1161_U504 | ~new_P2_R1161_U503;
  assign new_P2_R1161_U96 = ~new_P2_R1161_U375 | ~new_P2_R1161_U374;
  assign new_P2_R1161_U97 = ~new_P2_R1161_U380 | ~new_P2_R1161_U379;
  assign new_P2_R1161_U98 = ~new_P2_R1161_U387 | ~new_P2_R1161_U386;
  assign new_P2_R1161_U99 = ~new_P2_R1161_U394 | ~new_P2_R1161_U393;
  assign new_P2_R1161_U100 = ~new_P2_R1161_U399 | ~new_P2_R1161_U398;
  assign new_P2_R1161_U101 = ~new_P2_R1161_U408 | ~new_P2_R1161_U407;
  assign new_P2_R1161_U102 = ~new_P2_R1161_U415 | ~new_P2_R1161_U414;
  assign new_P2_R1161_U103 = ~new_P2_R1161_U422 | ~new_P2_R1161_U421;
  assign new_P2_R1161_U104 = ~new_P2_R1161_U429 | ~new_P2_R1161_U428;
  assign new_P2_R1161_U105 = ~new_P2_R1161_U434 | ~new_P2_R1161_U433;
  assign new_P2_R1161_U106 = ~new_P2_R1161_U441 | ~new_P2_R1161_U440;
  assign new_P2_R1161_U107 = ~new_P2_R1161_U448 | ~new_P2_R1161_U447;
  assign new_P2_R1161_U108 = ~new_P2_R1161_U462 | ~new_P2_R1161_U461;
  assign new_P2_R1161_U109 = ~new_P2_R1161_U467 | ~new_P2_R1161_U466;
  assign new_P2_R1161_U110 = ~new_P2_R1161_U474 | ~new_P2_R1161_U473;
  assign new_P2_R1161_U111 = ~new_P2_R1161_U481 | ~new_P2_R1161_U480;
  assign new_P2_R1161_U112 = ~new_P2_R1161_U488 | ~new_P2_R1161_U487;
  assign new_P2_R1161_U113 = ~new_P2_R1161_U495 | ~new_P2_R1161_U494;
  assign new_P2_R1161_U114 = ~new_P2_R1161_U500 | ~new_P2_R1161_U499;
  assign new_P2_R1161_U115 = new_P2_R1161_U189 & new_P2_R1161_U187;
  assign new_P2_R1161_U116 = new_P2_R1161_U4 & new_P2_R1161_U180;
  assign new_P2_R1161_U117 = new_P2_R1161_U194 & new_P2_R1161_U192;
  assign new_P2_R1161_U118 = new_P2_R1161_U201 & new_P2_R1161_U200;
  assign new_P2_R1161_U119 = new_P2_R1161_U22 & new_P2_R1161_U382 & new_P2_R1161_U381;
  assign new_P2_R1161_U120 = new_P2_R1161_U212 & new_P2_R1161_U5;
  assign new_P2_R1161_U121 = new_P2_R1161_U181 & new_P2_R1161_U180;
  assign new_P2_R1161_U122 = new_P2_R1161_U220 & new_P2_R1161_U218;
  assign new_P2_R1161_U123 = new_P2_R1161_U34 & new_P2_R1161_U389 & new_P2_R1161_U388;
  assign new_P2_R1161_U124 = new_P2_R1161_U226 & new_P2_R1161_U4;
  assign new_P2_R1161_U125 = new_P2_R1161_U234 & new_P2_R1161_U181;
  assign new_P2_R1161_U126 = new_P2_R1161_U204 & new_P2_R1161_U6;
  assign new_P2_R1161_U127 = new_P2_R1161_U243 & new_P2_R1161_U239;
  assign new_P2_R1161_U128 = new_P2_R1161_U250 & new_P2_R1161_U7;
  assign new_P2_R1161_U129 = new_P2_R1161_U253 & new_P2_R1161_U248;
  assign new_P2_R1161_U130 = new_P2_R1161_U268 & new_P2_R1161_U267;
  assign new_P2_R1161_U131 = new_P2_R1161_U9 & new_P2_R1161_U282;
  assign new_P2_R1161_U132 = new_P2_R1161_U285 & new_P2_R1161_U280;
  assign new_P2_R1161_U133 = new_P2_R1161_U301 & new_P2_R1161_U298;
  assign new_P2_R1161_U134 = new_P2_R1161_U368 & new_P2_R1161_U302;
  assign new_P2_R1161_U135 = new_P2_R1161_U160 & new_P2_R1161_U278;
  assign new_P2_R1161_U136 = new_P2_R1161_U80 & new_P2_R1161_U455 & new_P2_R1161_U454;
  assign new_P2_R1161_U137 = new_P2_R1161_U325 & new_P2_R1161_U9;
  assign new_P2_R1161_U138 = new_P2_R1161_U59 & new_P2_R1161_U469 & new_P2_R1161_U468;
  assign new_P2_R1161_U139 = new_P2_R1161_U334 & new_P2_R1161_U8;
  assign new_P2_R1161_U140 = new_P2_R1161_U172 & new_P2_R1161_U490 & new_P2_R1161_U489;
  assign new_P2_R1161_U141 = new_P2_R1161_U343 & new_P2_R1161_U7;
  assign new_P2_R1161_U142 = new_P2_R1161_U171 & new_P2_R1161_U502 & new_P2_R1161_U501;
  assign new_P2_R1161_U143 = new_P2_R1161_U350 & new_P2_R1161_U6;
  assign new_P2_R1161_U144 = ~new_P2_R1161_U118 | ~new_P2_R1161_U202;
  assign new_P2_R1161_U145 = ~new_P2_R1161_U217 | ~new_P2_R1161_U229;
  assign new_P2_R1161_U146 = ~new_P2_U3054;
  assign new_P2_R1161_U147 = ~new_P2_U3904;
  assign new_P2_R1161_U148 = new_P2_R1161_U403 & new_P2_R1161_U402;
  assign new_P2_R1161_U149 = ~new_P2_R1161_U364 | ~new_P2_R1161_U304 | ~new_P2_R1161_U169;
  assign new_P2_R1161_U150 = new_P2_R1161_U410 & new_P2_R1161_U409;
  assign new_P2_R1161_U151 = ~new_P2_R1161_U134 | ~new_P2_R1161_U370 | ~new_P2_R1161_U369;
  assign new_P2_R1161_U152 = new_P2_R1161_U417 & new_P2_R1161_U416;
  assign new_P2_R1161_U153 = ~new_P2_R1161_U86 | ~new_P2_R1161_U365 | ~new_P2_R1161_U299;
  assign new_P2_R1161_U154 = new_P2_R1161_U424 & new_P2_R1161_U423;
  assign new_P2_R1161_U155 = ~new_P2_R1161_U293 | ~new_P2_R1161_U292;
  assign new_P2_R1161_U156 = new_P2_R1161_U436 & new_P2_R1161_U435;
  assign new_P2_R1161_U157 = ~new_P2_R1161_U289 | ~new_P2_R1161_U288;
  assign new_P2_R1161_U158 = new_P2_R1161_U443 & new_P2_R1161_U442;
  assign new_P2_R1161_U159 = ~new_P2_R1161_U132 | ~new_P2_R1161_U284;
  assign new_P2_R1161_U160 = new_P2_R1161_U450 & new_P2_R1161_U449;
  assign new_P2_R1161_U161 = ~new_P2_R1161_U43 | ~new_P2_R1161_U327;
  assign new_P2_R1161_U162 = ~new_P2_R1161_U130 | ~new_P2_R1161_U269;
  assign new_P2_R1161_U163 = new_P2_R1161_U476 & new_P2_R1161_U475;
  assign new_P2_R1161_U164 = ~new_P2_R1161_U257 | ~new_P2_R1161_U256;
  assign new_P2_R1161_U165 = new_P2_R1161_U483 & new_P2_R1161_U482;
  assign new_P2_R1161_U166 = ~new_P2_R1161_U129 | ~new_P2_R1161_U252;
  assign new_P2_R1161_U167 = ~new_P2_R1161_U127 | ~new_P2_R1161_U242;
  assign new_P2_R1161_U168 = ~new_P2_R1161_U367 | ~new_P2_R1161_U366;
  assign new_P2_R1161_U169 = ~new_P2_U3053 | ~new_P2_R1161_U151;
  assign new_P2_R1161_U170 = ~new_P2_R1161_U34;
  assign new_P2_R1161_U171 = ~new_P2_U3416 | ~new_P2_U3082;
  assign new_P2_R1161_U172 = ~new_P2_U3071 | ~new_P2_U3425;
  assign new_P2_R1161_U173 = ~new_P2_U3057 | ~new_P2_U3898;
  assign new_P2_R1161_U174 = ~new_P2_R1161_U68;
  assign new_P2_R1161_U175 = ~new_P2_R1161_U77;
  assign new_P2_R1161_U176 = ~new_P2_U3064 | ~new_P2_U3899;
  assign new_P2_R1161_U177 = ~new_P2_R1161_U65;
  assign new_P2_R1161_U178 = new_P2_U3066 | new_P2_U3404;
  assign new_P2_R1161_U179 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1161_U180 = new_P2_U3398 | new_P2_U3063;
  assign new_P2_R1161_U181 = new_P2_U3395 | new_P2_U3067;
  assign new_P2_R1161_U182 = ~new_P2_R1161_U31;
  assign new_P2_R1161_U183 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1161_U184 = ~new_P2_R1161_U42;
  assign new_P2_R1161_U185 = ~new_P2_R1161_U43;
  assign new_P2_R1161_U186 = ~new_P2_R1161_U42 | ~new_P2_R1161_U43;
  assign new_P2_R1161_U187 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1161_U188 = ~new_P2_R1161_U186 | ~new_P2_R1161_U181;
  assign new_P2_R1161_U189 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1161_U190 = ~new_P2_R1161_U115 | ~new_P2_R1161_U188;
  assign new_P2_R1161_U191 = ~new_P2_R1161_U35 | ~new_P2_R1161_U34;
  assign new_P2_R1161_U192 = ~new_P2_U3066 | ~new_P2_R1161_U191;
  assign new_P2_R1161_U193 = ~new_P2_R1161_U116 | ~new_P2_R1161_U190;
  assign new_P2_R1161_U194 = ~new_P2_U3404 | ~new_P2_R1161_U170;
  assign new_P2_R1161_U195 = ~new_P2_R1161_U41;
  assign new_P2_R1161_U196 = new_P2_U3069 | new_P2_U3410;
  assign new_P2_R1161_U197 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1161_U198 = ~new_P2_R1161_U22;
  assign new_P2_R1161_U199 = ~new_P2_R1161_U23 | ~new_P2_R1161_U22;
  assign new_P2_R1161_U200 = ~new_P2_U3069 | ~new_P2_R1161_U199;
  assign new_P2_R1161_U201 = ~new_P2_U3410 | ~new_P2_R1161_U198;
  assign new_P2_R1161_U202 = ~new_P2_R1161_U5 | ~new_P2_R1161_U41;
  assign new_P2_R1161_U203 = ~new_P2_R1161_U144;
  assign new_P2_R1161_U204 = new_P2_U3413 | new_P2_U3083;
  assign new_P2_R1161_U205 = ~new_P2_R1161_U204 | ~new_P2_R1161_U144;
  assign new_P2_R1161_U206 = ~new_P2_R1161_U40;
  assign new_P2_R1161_U207 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1161_U208 = new_P2_U3407 | new_P2_U3070;
  assign new_P2_R1161_U209 = ~new_P2_R1161_U208 | ~new_P2_R1161_U41;
  assign new_P2_R1161_U210 = ~new_P2_R1161_U119 | ~new_P2_R1161_U209;
  assign new_P2_R1161_U211 = ~new_P2_R1161_U195 | ~new_P2_R1161_U22;
  assign new_P2_R1161_U212 = ~new_P2_U3410 | ~new_P2_U3069;
  assign new_P2_R1161_U213 = ~new_P2_R1161_U120 | ~new_P2_R1161_U211;
  assign new_P2_R1161_U214 = new_P2_U3070 | new_P2_U3407;
  assign new_P2_R1161_U215 = ~new_P2_R1161_U185 | ~new_P2_R1161_U181;
  assign new_P2_R1161_U216 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1161_U217 = ~new_P2_R1161_U45;
  assign new_P2_R1161_U218 = ~new_P2_R1161_U121 | ~new_P2_R1161_U184;
  assign new_P2_R1161_U219 = ~new_P2_R1161_U45 | ~new_P2_R1161_U180;
  assign new_P2_R1161_U220 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1161_U221 = ~new_P2_R1161_U44;
  assign new_P2_R1161_U222 = new_P2_U3401 | new_P2_U3059;
  assign new_P2_R1161_U223 = ~new_P2_R1161_U222 | ~new_P2_R1161_U44;
  assign new_P2_R1161_U224 = ~new_P2_R1161_U123 | ~new_P2_R1161_U223;
  assign new_P2_R1161_U225 = ~new_P2_R1161_U221 | ~new_P2_R1161_U34;
  assign new_P2_R1161_U226 = ~new_P2_U3404 | ~new_P2_U3066;
  assign new_P2_R1161_U227 = ~new_P2_R1161_U124 | ~new_P2_R1161_U225;
  assign new_P2_R1161_U228 = new_P2_U3059 | new_P2_U3401;
  assign new_P2_R1161_U229 = ~new_P2_R1161_U184 | ~new_P2_R1161_U181;
  assign new_P2_R1161_U230 = ~new_P2_R1161_U145;
  assign new_P2_R1161_U231 = ~new_P2_U3063 | ~new_P2_U3398;
  assign new_P2_R1161_U232 = ~new_P2_R1161_U42 | ~new_P2_R1161_U43 | ~new_P2_R1161_U401 | ~new_P2_R1161_U400;
  assign new_P2_R1161_U233 = ~new_P2_R1161_U43 | ~new_P2_R1161_U42;
  assign new_P2_R1161_U234 = ~new_P2_U3067 | ~new_P2_U3395;
  assign new_P2_R1161_U235 = ~new_P2_R1161_U125 | ~new_P2_R1161_U233;
  assign new_P2_R1161_U236 = new_P2_U3082 | new_P2_U3416;
  assign new_P2_R1161_U237 = new_P2_U3061 | new_P2_U3419;
  assign new_P2_R1161_U238 = ~new_P2_R1161_U177 | ~new_P2_R1161_U6;
  assign new_P2_R1161_U239 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1161_U240 = ~new_P2_R1161_U171 | ~new_P2_R1161_U238;
  assign new_P2_R1161_U241 = new_P2_U3419 | new_P2_U3061;
  assign new_P2_R1161_U242 = ~new_P2_R1161_U126 | ~new_P2_R1161_U144;
  assign new_P2_R1161_U243 = ~new_P2_R1161_U241 | ~new_P2_R1161_U240;
  assign new_P2_R1161_U244 = ~new_P2_R1161_U167;
  assign new_P2_R1161_U245 = new_P2_U3079 | new_P2_U3428;
  assign new_P2_R1161_U246 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1161_U247 = ~new_P2_R1161_U174 | ~new_P2_R1161_U7;
  assign new_P2_R1161_U248 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1161_U249 = ~new_P2_R1161_U172 | ~new_P2_R1161_U247;
  assign new_P2_R1161_U250 = new_P2_U3422 | new_P2_U3062;
  assign new_P2_R1161_U251 = new_P2_U3428 | new_P2_U3079;
  assign new_P2_R1161_U252 = ~new_P2_R1161_U128 | ~new_P2_R1161_U167;
  assign new_P2_R1161_U253 = ~new_P2_R1161_U251 | ~new_P2_R1161_U249;
  assign new_P2_R1161_U254 = ~new_P2_R1161_U166;
  assign new_P2_R1161_U255 = new_P2_U3431 | new_P2_U3078;
  assign new_P2_R1161_U256 = ~new_P2_R1161_U255 | ~new_P2_R1161_U166;
  assign new_P2_R1161_U257 = ~new_P2_U3078 | ~new_P2_U3431;
  assign new_P2_R1161_U258 = ~new_P2_R1161_U164;
  assign new_P2_R1161_U259 = new_P2_U3434 | new_P2_U3073;
  assign new_P2_R1161_U260 = ~new_P2_R1161_U259 | ~new_P2_R1161_U164;
  assign new_P2_R1161_U261 = ~new_P2_U3073 | ~new_P2_U3434;
  assign new_P2_R1161_U262 = ~new_P2_R1161_U92;
  assign new_P2_R1161_U263 = new_P2_U3068 | new_P2_U3440;
  assign new_P2_R1161_U264 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1161_U265 = ~new_P2_R1161_U59;
  assign new_P2_R1161_U266 = ~new_P2_R1161_U60 | ~new_P2_R1161_U59;
  assign new_P2_R1161_U267 = ~new_P2_U3068 | ~new_P2_R1161_U266;
  assign new_P2_R1161_U268 = ~new_P2_U3440 | ~new_P2_R1161_U265;
  assign new_P2_R1161_U269 = ~new_P2_R1161_U8 | ~new_P2_R1161_U92;
  assign new_P2_R1161_U270 = ~new_P2_R1161_U162;
  assign new_P2_R1161_U271 = new_P2_U3075 | new_P2_U3903;
  assign new_P2_R1161_U272 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1161_U273 = new_P2_U3074 | new_P2_U3902;
  assign new_P2_R1161_U274 = ~new_P2_R1161_U80;
  assign new_P2_R1161_U275 = ~new_P2_U3903 | ~new_P2_R1161_U274;
  assign new_P2_R1161_U276 = ~new_P2_R1161_U275 | ~new_P2_R1161_U90;
  assign new_P2_R1161_U277 = ~new_P2_R1161_U80 | ~new_P2_R1161_U81;
  assign new_P2_R1161_U278 = ~new_P2_R1161_U277 | ~new_P2_R1161_U276;
  assign new_P2_R1161_U279 = ~new_P2_R1161_U175 | ~new_P2_R1161_U9;
  assign new_P2_R1161_U280 = ~new_P2_U3074 | ~new_P2_U3902;
  assign new_P2_R1161_U281 = ~new_P2_R1161_U278 | ~new_P2_R1161_U279;
  assign new_P2_R1161_U282 = new_P2_U3443 | new_P2_U3081;
  assign new_P2_R1161_U283 = new_P2_U3902 | new_P2_U3074;
  assign new_P2_R1161_U284 = ~new_P2_R1161_U131 | ~new_P2_R1161_U273 | ~new_P2_R1161_U162;
  assign new_P2_R1161_U285 = ~new_P2_R1161_U283 | ~new_P2_R1161_U281;
  assign new_P2_R1161_U286 = ~new_P2_R1161_U159;
  assign new_P2_R1161_U287 = new_P2_U3901 | new_P2_U3060;
  assign new_P2_R1161_U288 = ~new_P2_R1161_U287 | ~new_P2_R1161_U159;
  assign new_P2_R1161_U289 = ~new_P2_U3060 | ~new_P2_U3901;
  assign new_P2_R1161_U290 = ~new_P2_R1161_U157;
  assign new_P2_R1161_U291 = new_P2_U3900 | new_P2_U3065;
  assign new_P2_R1161_U292 = ~new_P2_R1161_U291 | ~new_P2_R1161_U157;
  assign new_P2_R1161_U293 = ~new_P2_U3065 | ~new_P2_U3900;
  assign new_P2_R1161_U294 = ~new_P2_R1161_U155;
  assign new_P2_R1161_U295 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1161_U296 = ~new_P2_R1161_U176 | ~new_P2_R1161_U173;
  assign new_P2_R1161_U297 = ~new_P2_R1161_U86;
  assign new_P2_R1161_U298 = new_P2_U3899 | new_P2_U3064;
  assign new_P2_R1161_U299 = ~new_P2_R1161_U168 | ~new_P2_R1161_U155 | ~new_P2_R1161_U298;
  assign new_P2_R1161_U300 = ~new_P2_R1161_U153;
  assign new_P2_R1161_U301 = new_P2_U3896 | new_P2_U3052;
  assign new_P2_R1161_U302 = ~new_P2_U3052 | ~new_P2_U3896;
  assign new_P2_R1161_U303 = ~new_P2_R1161_U151;
  assign new_P2_R1161_U304 = ~new_P2_U3895 | ~new_P2_R1161_U151;
  assign new_P2_R1161_U305 = ~new_P2_R1161_U149;
  assign new_P2_R1161_U306 = ~new_P2_R1161_U298 | ~new_P2_R1161_U155;
  assign new_P2_R1161_U307 = ~new_P2_R1161_U89;
  assign new_P2_R1161_U308 = new_P2_U3898 | new_P2_U3057;
  assign new_P2_R1161_U309 = ~new_P2_R1161_U308 | ~new_P2_R1161_U89;
  assign new_P2_R1161_U310 = ~new_P2_R1161_U154 | ~new_P2_R1161_U309 | ~new_P2_R1161_U173;
  assign new_P2_R1161_U311 = ~new_P2_R1161_U307 | ~new_P2_R1161_U173;
  assign new_P2_R1161_U312 = ~new_P2_U3897 | ~new_P2_U3056;
  assign new_P2_R1161_U313 = ~new_P2_R1161_U168 | ~new_P2_R1161_U311 | ~new_P2_R1161_U312;
  assign new_P2_R1161_U314 = new_P2_U3057 | new_P2_U3898;
  assign new_P2_R1161_U315 = ~new_P2_R1161_U282 | ~new_P2_R1161_U162;
  assign new_P2_R1161_U316 = ~new_P2_R1161_U91;
  assign new_P2_R1161_U317 = ~new_P2_R1161_U9 | ~new_P2_R1161_U91;
  assign new_P2_R1161_U318 = ~new_P2_R1161_U135 | ~new_P2_R1161_U317;
  assign new_P2_R1161_U319 = ~new_P2_R1161_U317 | ~new_P2_R1161_U278;
  assign new_P2_R1161_U320 = ~new_P2_R1161_U453 | ~new_P2_R1161_U319;
  assign new_P2_R1161_U321 = new_P2_U3445 | new_P2_U3080;
  assign new_P2_R1161_U322 = ~new_P2_R1161_U321 | ~new_P2_R1161_U91;
  assign new_P2_R1161_U323 = ~new_P2_R1161_U136 | ~new_P2_R1161_U322;
  assign new_P2_R1161_U324 = ~new_P2_R1161_U316 | ~new_P2_R1161_U80;
  assign new_P2_R1161_U325 = ~new_P2_U3075 | ~new_P2_U3903;
  assign new_P2_R1161_U326 = ~new_P2_R1161_U137 | ~new_P2_R1161_U324;
  assign new_P2_R1161_U327 = new_P2_U3392 | new_P2_U3077;
  assign new_P2_R1161_U328 = ~new_P2_R1161_U161;
  assign new_P2_R1161_U329 = new_P2_U3080 | new_P2_U3445;
  assign new_P2_R1161_U330 = new_P2_U3437 | new_P2_U3072;
  assign new_P2_R1161_U331 = ~new_P2_R1161_U330 | ~new_P2_R1161_U92;
  assign new_P2_R1161_U332 = ~new_P2_R1161_U138 | ~new_P2_R1161_U331;
  assign new_P2_R1161_U333 = ~new_P2_R1161_U262 | ~new_P2_R1161_U59;
  assign new_P2_R1161_U334 = ~new_P2_U3440 | ~new_P2_U3068;
  assign new_P2_R1161_U335 = ~new_P2_R1161_U139 | ~new_P2_R1161_U333;
  assign new_P2_R1161_U336 = new_P2_U3072 | new_P2_U3437;
  assign new_P2_R1161_U337 = ~new_P2_R1161_U250 | ~new_P2_R1161_U167;
  assign new_P2_R1161_U338 = ~new_P2_R1161_U93;
  assign new_P2_R1161_U339 = new_P2_U3425 | new_P2_U3071;
  assign new_P2_R1161_U340 = ~new_P2_R1161_U339 | ~new_P2_R1161_U93;
  assign new_P2_R1161_U341 = ~new_P2_R1161_U140 | ~new_P2_R1161_U340;
  assign new_P2_R1161_U342 = ~new_P2_R1161_U338 | ~new_P2_R1161_U172;
  assign new_P2_R1161_U343 = ~new_P2_U3079 | ~new_P2_U3428;
  assign new_P2_R1161_U344 = ~new_P2_R1161_U141 | ~new_P2_R1161_U342;
  assign new_P2_R1161_U345 = new_P2_U3071 | new_P2_U3425;
  assign new_P2_R1161_U346 = new_P2_U3416 | new_P2_U3082;
  assign new_P2_R1161_U347 = ~new_P2_R1161_U346 | ~new_P2_R1161_U40;
  assign new_P2_R1161_U348 = ~new_P2_R1161_U142 | ~new_P2_R1161_U347;
  assign new_P2_R1161_U349 = ~new_P2_R1161_U206 | ~new_P2_R1161_U171;
  assign new_P2_R1161_U350 = ~new_P2_U3061 | ~new_P2_U3419;
  assign new_P2_R1161_U351 = ~new_P2_R1161_U143 | ~new_P2_R1161_U349;
  assign new_P2_R1161_U352 = ~new_P2_R1161_U207 | ~new_P2_R1161_U171;
  assign new_P2_R1161_U353 = ~new_P2_R1161_U204 | ~new_P2_R1161_U65;
  assign new_P2_R1161_U354 = ~new_P2_R1161_U214 | ~new_P2_R1161_U22;
  assign new_P2_R1161_U355 = ~new_P2_R1161_U228 | ~new_P2_R1161_U34;
  assign new_P2_R1161_U356 = ~new_P2_R1161_U231 | ~new_P2_R1161_U180;
  assign new_P2_R1161_U357 = ~new_P2_R1161_U314 | ~new_P2_R1161_U173;
  assign new_P2_R1161_U358 = ~new_P2_R1161_U298 | ~new_P2_R1161_U176;
  assign new_P2_R1161_U359 = ~new_P2_R1161_U329 | ~new_P2_R1161_U80;
  assign new_P2_R1161_U360 = ~new_P2_R1161_U282 | ~new_P2_R1161_U77;
  assign new_P2_R1161_U361 = ~new_P2_R1161_U336 | ~new_P2_R1161_U59;
  assign new_P2_R1161_U362 = ~new_P2_R1161_U345 | ~new_P2_R1161_U172;
  assign new_P2_R1161_U363 = ~new_P2_R1161_U250 | ~new_P2_R1161_U68;
  assign new_P2_R1161_U364 = ~new_P2_U3895 | ~new_P2_U3053;
  assign new_P2_R1161_U365 = ~new_P2_R1161_U296 | ~new_P2_R1161_U168;
  assign new_P2_R1161_U366 = ~new_P2_U3056 | ~new_P2_R1161_U295;
  assign new_P2_R1161_U367 = ~new_P2_U3897 | ~new_P2_R1161_U295;
  assign new_P2_R1161_U368 = ~new_P2_R1161_U301 | ~new_P2_R1161_U296 | ~new_P2_R1161_U168;
  assign new_P2_R1161_U369 = ~new_P2_R1161_U133 | ~new_P2_R1161_U155 | ~new_P2_R1161_U168;
  assign new_P2_R1161_U370 = ~new_P2_R1161_U297 | ~new_P2_R1161_U301;
  assign new_P2_R1161_U371 = ~new_P2_U3082 | ~new_P2_R1161_U39;
  assign new_P2_R1161_U372 = ~new_P2_U3416 | ~new_P2_R1161_U38;
  assign new_P2_R1161_U373 = ~new_P2_R1161_U372 | ~new_P2_R1161_U371;
  assign new_P2_R1161_U374 = ~new_P2_R1161_U352 | ~new_P2_R1161_U40;
  assign new_P2_R1161_U375 = ~new_P2_R1161_U373 | ~new_P2_R1161_U206;
  assign new_P2_R1161_U376 = ~new_P2_U3083 | ~new_P2_R1161_U36;
  assign new_P2_R1161_U377 = ~new_P2_U3413 | ~new_P2_R1161_U37;
  assign new_P2_R1161_U378 = ~new_P2_R1161_U377 | ~new_P2_R1161_U376;
  assign new_P2_R1161_U379 = ~new_P2_R1161_U353 | ~new_P2_R1161_U144;
  assign new_P2_R1161_U380 = ~new_P2_R1161_U203 | ~new_P2_R1161_U378;
  assign new_P2_R1161_U381 = ~new_P2_U3069 | ~new_P2_R1161_U23;
  assign new_P2_R1161_U382 = ~new_P2_U3410 | ~new_P2_R1161_U21;
  assign new_P2_R1161_U383 = ~new_P2_U3070 | ~new_P2_R1161_U19;
  assign new_P2_R1161_U384 = ~new_P2_U3407 | ~new_P2_R1161_U20;
  assign new_P2_R1161_U385 = ~new_P2_R1161_U384 | ~new_P2_R1161_U383;
  assign new_P2_R1161_U386 = ~new_P2_R1161_U354 | ~new_P2_R1161_U41;
  assign new_P2_R1161_U387 = ~new_P2_R1161_U385 | ~new_P2_R1161_U195;
  assign new_P2_R1161_U388 = ~new_P2_U3066 | ~new_P2_R1161_U35;
  assign new_P2_R1161_U389 = ~new_P2_U3404 | ~new_P2_R1161_U26;
  assign new_P2_R1161_U390 = ~new_P2_U3059 | ~new_P2_R1161_U24;
  assign new_P2_R1161_U391 = ~new_P2_U3401 | ~new_P2_R1161_U25;
  assign new_P2_R1161_U392 = ~new_P2_R1161_U391 | ~new_P2_R1161_U390;
  assign new_P2_R1161_U393 = ~new_P2_R1161_U355 | ~new_P2_R1161_U44;
  assign new_P2_R1161_U394 = ~new_P2_R1161_U392 | ~new_P2_R1161_U221;
  assign new_P2_R1161_U395 = ~new_P2_U3063 | ~new_P2_R1161_U32;
  assign new_P2_R1161_U396 = ~new_P2_U3398 | ~new_P2_R1161_U33;
  assign new_P2_R1161_U397 = ~new_P2_R1161_U396 | ~new_P2_R1161_U395;
  assign new_P2_R1161_U398 = ~new_P2_R1161_U356 | ~new_P2_R1161_U145;
  assign new_P2_R1161_U399 = ~new_P2_R1161_U230 | ~new_P2_R1161_U397;
  assign new_P2_R1161_U400 = ~new_P2_U3067 | ~new_P2_R1161_U27;
  assign new_P2_R1161_U401 = ~new_P2_U3395 | ~new_P2_R1161_U28;
  assign new_P2_R1161_U402 = ~new_P2_U3054 | ~new_P2_R1161_U147;
  assign new_P2_R1161_U403 = ~new_P2_U3904 | ~new_P2_R1161_U146;
  assign new_P2_R1161_U404 = ~new_P2_U3054 | ~new_P2_R1161_U147;
  assign new_P2_R1161_U405 = ~new_P2_U3904 | ~new_P2_R1161_U146;
  assign new_P2_R1161_U406 = ~new_P2_R1161_U405 | ~new_P2_R1161_U404;
  assign new_P2_R1161_U407 = ~new_P2_R1161_U148 | ~new_P2_R1161_U149;
  assign new_P2_R1161_U408 = ~new_P2_R1161_U305 | ~new_P2_R1161_U406;
  assign new_P2_R1161_U409 = ~new_P2_U3053 | ~new_P2_R1161_U88;
  assign new_P2_R1161_U410 = ~new_P2_U3895 | ~new_P2_R1161_U87;
  assign new_P2_R1161_U411 = ~new_P2_U3053 | ~new_P2_R1161_U88;
  assign new_P2_R1161_U412 = ~new_P2_U3895 | ~new_P2_R1161_U87;
  assign new_P2_R1161_U413 = ~new_P2_R1161_U412 | ~new_P2_R1161_U411;
  assign new_P2_R1161_U414 = ~new_P2_R1161_U150 | ~new_P2_R1161_U151;
  assign new_P2_R1161_U415 = ~new_P2_R1161_U303 | ~new_P2_R1161_U413;
  assign new_P2_R1161_U416 = ~new_P2_U3052 | ~new_P2_R1161_U46;
  assign new_P2_R1161_U417 = ~new_P2_U3896 | ~new_P2_R1161_U47;
  assign new_P2_R1161_U418 = ~new_P2_U3052 | ~new_P2_R1161_U46;
  assign new_P2_R1161_U419 = ~new_P2_U3896 | ~new_P2_R1161_U47;
  assign new_P2_R1161_U420 = ~new_P2_R1161_U419 | ~new_P2_R1161_U418;
  assign new_P2_R1161_U421 = ~new_P2_R1161_U152 | ~new_P2_R1161_U153;
  assign new_P2_R1161_U422 = ~new_P2_R1161_U300 | ~new_P2_R1161_U420;
  assign new_P2_R1161_U423 = ~new_P2_U3056 | ~new_P2_R1161_U49;
  assign new_P2_R1161_U424 = ~new_P2_U3897 | ~new_P2_R1161_U48;
  assign new_P2_R1161_U425 = ~new_P2_U3057 | ~new_P2_R1161_U50;
  assign new_P2_R1161_U426 = ~new_P2_U3898 | ~new_P2_R1161_U51;
  assign new_P2_R1161_U427 = ~new_P2_R1161_U426 | ~new_P2_R1161_U425;
  assign new_P2_R1161_U428 = ~new_P2_R1161_U357 | ~new_P2_R1161_U89;
  assign new_P2_R1161_U429 = ~new_P2_R1161_U427 | ~new_P2_R1161_U307;
  assign new_P2_R1161_U430 = ~new_P2_U3064 | ~new_P2_R1161_U52;
  assign new_P2_R1161_U431 = ~new_P2_U3899 | ~new_P2_R1161_U53;
  assign new_P2_R1161_U432 = ~new_P2_R1161_U431 | ~new_P2_R1161_U430;
  assign new_P2_R1161_U433 = ~new_P2_R1161_U358 | ~new_P2_R1161_U155;
  assign new_P2_R1161_U434 = ~new_P2_R1161_U294 | ~new_P2_R1161_U432;
  assign new_P2_R1161_U435 = ~new_P2_U3065 | ~new_P2_R1161_U84;
  assign new_P2_R1161_U436 = ~new_P2_U3900 | ~new_P2_R1161_U85;
  assign new_P2_R1161_U437 = ~new_P2_U3065 | ~new_P2_R1161_U84;
  assign new_P2_R1161_U438 = ~new_P2_U3900 | ~new_P2_R1161_U85;
  assign new_P2_R1161_U439 = ~new_P2_R1161_U438 | ~new_P2_R1161_U437;
  assign new_P2_R1161_U440 = ~new_P2_R1161_U156 | ~new_P2_R1161_U157;
  assign new_P2_R1161_U441 = ~new_P2_R1161_U290 | ~new_P2_R1161_U439;
  assign new_P2_R1161_U442 = ~new_P2_U3060 | ~new_P2_R1161_U82;
  assign new_P2_R1161_U443 = ~new_P2_U3901 | ~new_P2_R1161_U83;
  assign new_P2_R1161_U444 = ~new_P2_U3060 | ~new_P2_R1161_U82;
  assign new_P2_R1161_U445 = ~new_P2_U3901 | ~new_P2_R1161_U83;
  assign new_P2_R1161_U446 = ~new_P2_R1161_U445 | ~new_P2_R1161_U444;
  assign new_not_keyinput0 = ~keyinput0;
  assign new_not_keyinput1 = ~keyinput1;
  assign new_not_keyinput2 = ~keyinput2;
  assign new_not_keyinput3 = ~keyinput3;
  assign new_not_keyinput4 = ~keyinput4;
  assign new_not_0 = ~Q_1;
  assign new_and_1 = new_not_0 & Q_3;
  assign new_not_2 = ~Q_2;
  assign new_and_3 = new_not_2 & Q_3;
  assign new_not_4 = ~Q_0;
  assign new_and_5 = new_not_4 & Q_3;
  assign new_not_6 = ~Q_3;
  assign new_and_7 = new_not_6 & Q_2 & Q_0 & Q_1;
  assign n41489 = new_and_7 | new_and_5 | new_and_1 | new_and_3;
  assign new_not_9 = ~Q_2;
  assign new_and_10 = new_not_9 & Q_0 & Q_1;
  assign new_not_11 = ~Q_0;
  assign new_and_12 = new_not_11 & Q_2;
  assign new_not_13 = ~Q_1;
  assign new_and_14 = new_not_13 & Q_2;
  assign n41486 = new_and_14 | new_and_10 | new_and_12;
  assign new_not_16 = ~Q_1;
  assign new_and_17 = Q_0 & new_not_16;
  assign new_not_18 = ~Q_0;
  assign new_and_19 = new_not_18 & Q_1;
  assign n41483 = new_and_17 | new_and_19;
  assign n41480 = ~Q_0;
  assign new_not_Q_0 = ~Q_0;
  assign new_not_Q_1 = ~Q_1;
  assign new_not_Q_2 = ~Q_2;
  assign new_not_Q_3 = ~Q_3;
  assign new_count_state_1 = Q_0 & new_not_Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_2 = new_not_Q_0 & Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_3 = Q_0 & Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_4 = new_not_Q_0 & new_not_Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_5 = Q_0 & new_not_Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_6 = new_not_Q_0 & Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_7 = Q_0 & Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_8 = new_not_Q_0 & new_not_Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_9 = Q_0 & new_not_Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_10 = new_not_Q_0 & Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_11 = Q_0 & Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_12 = new_not_Q_0 & new_not_Q_1 & Q_3 & Q_2;
  assign new_count_state_13 = Q_0 & new_not_Q_1 & Q_3 & Q_2;
  assign new_count_state_14 = new_not_Q_0 & Q_1 & Q_3 & Q_2;
  assign new_count_state_15 = Q_0 & Q_1 & Q_3 & Q_2;
  assign new_y_mux_key0_and_0 = n130 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_1 = new_P1_U3355 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0 = new_y_mux_key0_and_0 | new_y_mux_key0_and_1;
  assign new_y_mux_key1_and_0 = n130 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key1_and_1 = new_P1_U3355 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1 = new_y_mux_key1_and_0 | new_y_mux_key1_and_1;
  assign new_y_mux_key2_and_0 = n130 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key2_and_1 = new_P1_U3355 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2 = new_y_mux_key2_and_0 | new_y_mux_key2_and_1;
  assign new_y_mux_key3_and_0 = n130 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_1 = new_P1_U3355 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3 = new_y_mux_key3_and_0 | new_y_mux_key3_and_1;
  assign new_y_mux_key4_and_0 = n130 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key4_and_1 = new_P1_U3355 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4 = new_y_mux_key4_and_0 | new_y_mux_key4_and_1;
  assign new_y_mux_key5_and_0 = n130 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_1 = new_P1_U3355 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5 = new_y_mux_key5_and_0 | new_y_mux_key5_and_1;
  assign new_y_mux_key6_and_0 = n130 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6_and_1 = new_P1_U3355 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6 = new_y_mux_key6_and_0 | new_y_mux_key6_and_1;
  assign new_y_mux_key7_and_0 = n130 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_1 = new_P1_U3355 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7 = new_y_mux_key7_and_0 | new_y_mux_key7_and_1;
  assign new_y_mux_key8_and_0 = n130 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_1 = new_P1_U3355 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8 = new_y_mux_key8_and_0 | new_y_mux_key8_and_1;
  assign new_y_mux_key9_and_0 = n130 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9_and_1 = new_P1_U3355 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9 = new_y_mux_key9_and_0 | new_y_mux_key9_and_1;
  assign new_y_mux_key10_and_0 = n130 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_1 = new_P1_U3355 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10 = new_y_mux_key10_and_0 | new_y_mux_key10_and_1;
  assign new_y_mux_key11_and_0 = n130 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11_and_1 = new_P1_U3355 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11 = new_y_mux_key11_and_0 | new_y_mux_key11_and_1;
  assign new_y_mux_key12_and_0 = n130 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key12_and_1 = new_P1_U3355 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12 = new_y_mux_key12_and_0 | new_y_mux_key12_and_1;
  assign new_y_mux_key13_and_0 = n130 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_1 = new_P1_U3355 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key13 = new_y_mux_key13_and_0 | new_y_mux_key13_and_1;
  assign new_y_mux_key14_and_0 = n130 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_1 = new_P1_U3355 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14 = new_y_mux_key14_and_0 | new_y_mux_key14_and_1;
  assign new_y_mux_key15_and_0 = n130 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_1 = new_P1_U3355 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15 = new_y_mux_key15_and_0 | new_y_mux_key15_and_1;
  assign new__state_1 = new_count_state_1;
  assign new__state_2 = new_count_state_2;
  assign new__state_3 = new_count_state_3;
  assign new__state_4 = new_count_state_4;
  assign new__state_5 = new_count_state_5;
  assign new__state_6 = new_count_state_6;
  assign new__state_7 = new_count_state_7;
  assign new__state_8 = new_count_state_8;
  assign new__state_9 = new_count_state_9;
  assign new__state_10 = new_count_state_10;
  assign new__state_11 = new_count_state_11;
  assign new__state_12 = new_count_state_12;
  assign new__state_13 = new_count_state_13;
  assign new__state_14 = new_count_state_14;
  assign new__state_15 = new_count_state_15;
  assign new__state_17 = new__state_2 | new__state_3;
  assign new__state_18 = new__state_4 | new__state_5;
  assign new__state_19 = new__state_6 | new__state_7;
  assign new__state_20 = new__state_8 | new__state_9;
  assign new__state_21 = new__state_10 | new__state_11;
  assign new__state_22 = new__state_12 | new__state_13;
  assign new__state_23 = new__state_14 | new__state_15;
  assign new__state_25 = new__state_18 | new__state_19;
  assign new__state_26 = new__state_20 | new__state_21;
  assign new__state_27 = new__state_22 | new__state_23;
  assign new__state_29 = new__state_26 | new__state_27;
  assign new_s__state_1 = new__state_1;
  assign new_not_s__state_1 = ~new_s__state_1;
  assign new_I0__state_1 = new_y_mux_key0;
  assign new_I1__state_1 = new_y_mux_key1;
  assign new_and_mux__state_1 = new_not_s__state_1 & new_I0__state_1;
  assign new_and_mux__state_1_2 = new_s__state_1 & new_I1__state_1;
  assign new_y_mux_16 = new_and_mux__state_1 | new_and_mux__state_1_2;
  assign new_s__state_3 = new__state_3;
  assign new_not_s__state_3 = ~new_s__state_3;
  assign new_I0__state_3 = new_y_mux_key2;
  assign new_I1__state_3 = new_y_mux_key3;
  assign new_and_mux__state_3 = new_not_s__state_3 & new_I0__state_3;
  assign new_and_mux__state_3_2 = new_s__state_3 & new_I1__state_3;
  assign new_y_mux_17 = new_and_mux__state_3 | new_and_mux__state_3_2;
  assign new_s__state_5 = new__state_5;
  assign new_not_s__state_5 = ~new_s__state_5;
  assign new_I0__state_5 = new_y_mux_key4;
  assign new_I1__state_5 = new_y_mux_key5;
  assign new_and_mux__state_5 = new_not_s__state_5 & new_I0__state_5;
  assign new_and_mux__state_5_2 = new_s__state_5 & new_I1__state_5;
  assign new_y_mux_18 = new_and_mux__state_5 | new_and_mux__state_5_2;
  assign new_s__state_7 = new__state_7;
  assign new_not_s__state_7 = ~new_s__state_7;
  assign new_I0__state_7 = new_y_mux_key6;
  assign new_I1__state_7 = new_y_mux_key7;
  assign new_and_mux__state_7 = new_not_s__state_7 & new_I0__state_7;
  assign new_and_mux__state_7_2 = new_s__state_7 & new_I1__state_7;
  assign new_y_mux_19 = new_and_mux__state_7 | new_and_mux__state_7_2;
  assign new_s__state_9 = new__state_9;
  assign new_not_s__state_9 = ~new_s__state_9;
  assign new_I0__state_9 = new_y_mux_key8;
  assign new_I1__state_9 = new_y_mux_key9;
  assign new_and_mux__state_9 = new_not_s__state_9 & new_I0__state_9;
  assign new_and_mux__state_9_2 = new_s__state_9 & new_I1__state_9;
  assign new_y_mux_20 = new_and_mux__state_9 | new_and_mux__state_9_2;
  assign new_s__state_11 = new__state_11;
  assign new_not_s__state_11 = ~new_s__state_11;
  assign new_I0__state_11 = new_y_mux_key10;
  assign new_I1__state_11 = new_y_mux_key11;
  assign new_and_mux__state_11 = new_not_s__state_11 & new_I0__state_11;
  assign new_and_mux__state_11_2 = new_s__state_11 & new_I1__state_11;
  assign new_y_mux_21 = new_and_mux__state_11 | new_and_mux__state_11_2;
  assign new_s__state_13 = new__state_13;
  assign new_not_s__state_13 = ~new_s__state_13;
  assign new_I0__state_13 = new_y_mux_key12;
  assign new_I1__state_13 = new_y_mux_key13;
  assign new_and_mux__state_13 = new_not_s__state_13 & new_I0__state_13;
  assign new_and_mux__state_13_2 = new_s__state_13 & new_I1__state_13;
  assign new_y_mux_22 = new_and_mux__state_13 | new_and_mux__state_13_2;
  assign new_s__state_15 = new__state_15;
  assign new_not_s__state_15 = ~new_s__state_15;
  assign new_I0__state_15 = new_y_mux_key14;
  assign new_I1__state_15 = new_y_mux_key15;
  assign new_and_mux__state_15 = new_not_s__state_15 & new_I0__state_15;
  assign new_and_mux__state_15_2 = new_s__state_15 & new_I1__state_15;
  assign new_y_mux_23 = new_and_mux__state_15 | new_and_mux__state_15_2;
  assign new_s__state_17 = new__state_17;
  assign new_not_s__state_17 = ~new_s__state_17;
  assign new_I0__state_17 = new_y_mux_16;
  assign new_I1__state_17 = new_y_mux_17;
  assign new_and_mux__state_17 = new_not_s__state_17 & new_I0__state_17;
  assign new_and_mux__state_17_2 = new_s__state_17 & new_I1__state_17;
  assign new_y_mux_24 = new_and_mux__state_17 | new_and_mux__state_17_2;
  assign new_s__state_19 = new__state_19;
  assign new_not_s__state_19 = ~new_s__state_19;
  assign new_I0__state_19 = new_y_mux_18;
  assign new_I1__state_19 = new_y_mux_19;
  assign new_and_mux__state_19 = new_not_s__state_19 & new_I0__state_19;
  assign new_and_mux__state_19_2 = new_s__state_19 & new_I1__state_19;
  assign new_y_mux_25 = new_and_mux__state_19 | new_and_mux__state_19_2;
  assign new_s__state_21 = new__state_21;
  assign new_not_s__state_21 = ~new_s__state_21;
  assign new_I0__state_21 = new_y_mux_20;
  assign new_I1__state_21 = new_y_mux_21;
  assign new_and_mux__state_21 = new_not_s__state_21 & new_I0__state_21;
  assign new_and_mux__state_21_2 = new_s__state_21 & new_I1__state_21;
  assign new_y_mux_26 = new_and_mux__state_21 | new_and_mux__state_21_2;
  assign new_s__state_23 = new__state_23;
  assign new_not_s__state_23 = ~new_s__state_23;
  assign new_I0__state_23 = new_y_mux_22;
  assign new_I1__state_23 = new_y_mux_23;
  assign new_and_mux__state_23 = new_not_s__state_23 & new_I0__state_23;
  assign new_and_mux__state_23_2 = new_s__state_23 & new_I1__state_23;
  assign new_y_mux_27 = new_and_mux__state_23 | new_and_mux__state_23_2;
  assign new_s__state_25 = new__state_25;
  assign new_not_s__state_25 = ~new_s__state_25;
  assign new_I0__state_25 = new_y_mux_24;
  assign new_I1__state_25 = new_y_mux_25;
  assign new_and_mux__state_25 = new_not_s__state_25 & new_I0__state_25;
  assign new_and_mux__state_25_2 = new_s__state_25 & new_I1__state_25;
  assign new_y_mux_28 = new_and_mux__state_25 | new_and_mux__state_25_2;
  assign new_s__state_27 = new__state_27;
  assign new_not_s__state_27 = ~new_s__state_27;
  assign new_I0__state_27 = new_y_mux_26;
  assign new_I1__state_27 = new_y_mux_27;
  assign new_and_mux__state_27 = new_not_s__state_27 & new_I0__state_27;
  assign new_and_mux__state_27_2 = new_s__state_27 & new_I1__state_27;
  assign new_y_mux_29 = new_and_mux__state_27 | new_and_mux__state_27_2;
  assign new_s__state_29 = new__state_29;
  assign new_not_s__state_29 = ~new_s__state_29;
  assign new_I0__state_29 = new_y_mux_28;
  assign new_I1__state_29 = new_y_mux_29;
  assign new_and_mux__state_29 = new_not_s__state_29 & new_I0__state_29;
  assign new_and_mux__state_29_2 = new_s__state_29 & new_I1__state_29;
  assign n120 = new_and_mux__state_29 | new_and_mux__state_29_2;
  always @ (posedge clock) begin
    P1_IR_REG_0_ <= n120;
    P1_IR_REG_1_ <= n125;
    P1_IR_REG_2_ <= n130;
    P1_IR_REG_3_ <= n135;
    P1_IR_REG_4_ <= n140;
    P1_IR_REG_5_ <= n145;
    P1_IR_REG_6_ <= n150;
    P1_IR_REG_7_ <= n155;
    P1_IR_REG_8_ <= n160;
    P1_IR_REG_9_ <= n165;
    P1_IR_REG_10_ <= n170;
    P1_IR_REG_11_ <= n175;
    P1_IR_REG_12_ <= n180;
    P1_IR_REG_13_ <= n185;
    P1_IR_REG_14_ <= n190;
    P1_IR_REG_15_ <= n195;
    P1_IR_REG_16_ <= n200;
    P1_IR_REG_17_ <= n205;
    P1_IR_REG_18_ <= n210;
    P1_IR_REG_19_ <= n215;
    P1_IR_REG_20_ <= n220;
    P1_IR_REG_21_ <= n225;
    P1_IR_REG_22_ <= n230;
    P1_IR_REG_23_ <= n235;
    P1_IR_REG_24_ <= n240;
    P1_IR_REG_25_ <= n245;
    P1_IR_REG_26_ <= n250;
    P1_IR_REG_27_ <= n255;
    P1_IR_REG_28_ <= n260;
    P1_IR_REG_29_ <= n265;
    P1_IR_REG_30_ <= n270;
    P1_IR_REG_31_ <= n275;
    P1_D_REG_0_ <= n280;
    P1_D_REG_1_ <= n285;
    P1_D_REG_2_ <= n290;
    P1_D_REG_3_ <= n295;
    P1_D_REG_4_ <= n300;
    P1_D_REG_5_ <= n305;
    P1_D_REG_6_ <= n310;
    P1_D_REG_7_ <= n315;
    P1_D_REG_8_ <= n320;
    P1_D_REG_9_ <= n325;
    P1_D_REG_10_ <= n330;
    P1_D_REG_11_ <= n335;
    P1_D_REG_12_ <= n340;
    P1_D_REG_13_ <= n345;
    P1_D_REG_14_ <= n350;
    P1_D_REG_15_ <= n355;
    P1_D_REG_16_ <= n360;
    P1_D_REG_17_ <= n365;
    P1_D_REG_18_ <= n370;
    P1_D_REG_19_ <= n375;
    P1_D_REG_20_ <= n380;
    P1_D_REG_21_ <= n385;
    P1_D_REG_22_ <= n390;
    P1_D_REG_23_ <= n395;
    P1_D_REG_24_ <= n400;
    P1_D_REG_25_ <= n405;
    P1_D_REG_26_ <= n410;
    P1_D_REG_27_ <= n415;
    P1_D_REG_28_ <= n420;
    P1_D_REG_29_ <= n425;
    P1_D_REG_30_ <= n430;
    P1_D_REG_31_ <= n435;
    P1_REG0_REG_0_ <= n440;
    P1_REG0_REG_1_ <= n445;
    P1_REG0_REG_2_ <= n450;
    P1_REG0_REG_3_ <= n455;
    P1_REG0_REG_4_ <= n460;
    P1_REG0_REG_5_ <= n465;
    P1_REG0_REG_6_ <= n470;
    P1_REG0_REG_7_ <= n475;
    P1_REG0_REG_8_ <= n480;
    P1_REG0_REG_9_ <= n485;
    P1_REG0_REG_10_ <= n490;
    P1_REG0_REG_11_ <= n495;
    P1_REG0_REG_12_ <= n500;
    P1_REG0_REG_13_ <= n505;
    P1_REG0_REG_14_ <= n510;
    P1_REG0_REG_15_ <= n515;
    P1_REG0_REG_16_ <= n520;
    P1_REG0_REG_17_ <= n525;
    P1_REG0_REG_18_ <= n530;
    P1_REG0_REG_19_ <= n535;
    P1_REG0_REG_20_ <= n540;
    P1_REG0_REG_21_ <= n545;
    P1_REG0_REG_22_ <= n550;
    P1_REG0_REG_23_ <= n555;
    P1_REG0_REG_24_ <= n560;
    P1_REG0_REG_25_ <= n565;
    P1_REG0_REG_26_ <= n570;
    P1_REG0_REG_27_ <= n575;
    P1_REG0_REG_28_ <= n580;
    P1_REG0_REG_29_ <= n585;
    P1_REG0_REG_30_ <= n590;
    P1_REG0_REG_31_ <= n595;
    P1_REG1_REG_0_ <= n600;
    P1_REG1_REG_1_ <= n605;
    P1_REG1_REG_2_ <= n610;
    P1_REG1_REG_3_ <= n615;
    P1_REG1_REG_4_ <= n620;
    P1_REG1_REG_5_ <= n625;
    P1_REG1_REG_6_ <= n630;
    P1_REG1_REG_7_ <= n635;
    P1_REG1_REG_8_ <= n640;
    P1_REG1_REG_9_ <= n645;
    P1_REG1_REG_10_ <= n650;
    P1_REG1_REG_11_ <= n655;
    P1_REG1_REG_12_ <= n660;
    P1_REG1_REG_13_ <= n665;
    P1_REG1_REG_14_ <= n670;
    P1_REG1_REG_15_ <= n675;
    P1_REG1_REG_16_ <= n680;
    P1_REG1_REG_17_ <= n685;
    P1_REG1_REG_18_ <= n690;
    P1_REG1_REG_19_ <= n695;
    P1_REG1_REG_20_ <= n700;
    P1_REG1_REG_21_ <= n705;
    P1_REG1_REG_22_ <= n710;
    P1_REG1_REG_23_ <= n715;
    P1_REG1_REG_24_ <= n720;
    P1_REG1_REG_25_ <= n725;
    P1_REG1_REG_26_ <= n730;
    P1_REG1_REG_27_ <= n735;
    P1_REG1_REG_28_ <= n740;
    P1_REG1_REG_29_ <= n745;
    P1_REG1_REG_30_ <= n750;
    P1_REG1_REG_31_ <= n755;
    P1_REG2_REG_0_ <= n760;
    P1_REG2_REG_1_ <= n765;
    P1_REG2_REG_2_ <= n770;
    P1_REG2_REG_3_ <= n775;
    P1_REG2_REG_4_ <= n780;
    P1_REG2_REG_5_ <= n785;
    P1_REG2_REG_6_ <= n790;
    P1_REG2_REG_7_ <= n795;
    P1_REG2_REG_8_ <= n800;
    P1_REG2_REG_9_ <= n805;
    P1_REG2_REG_10_ <= n810;
    P1_REG2_REG_11_ <= n815;
    P1_REG2_REG_12_ <= n820;
    P1_REG2_REG_13_ <= n825;
    P1_REG2_REG_14_ <= n830;
    P1_REG2_REG_15_ <= n835;
    P1_REG2_REG_16_ <= n840;
    P1_REG2_REG_17_ <= n845;
    P1_REG2_REG_18_ <= n850;
    P1_REG2_REG_19_ <= n855;
    P1_REG2_REG_20_ <= n860;
    P1_REG2_REG_21_ <= n865;
    P1_REG2_REG_22_ <= n870;
    P1_REG2_REG_23_ <= n875;
    P1_REG2_REG_24_ <= n880;
    P1_REG2_REG_25_ <= n885;
    P1_REG2_REG_26_ <= n890;
    P1_REG2_REG_27_ <= n895;
    P1_REG2_REG_28_ <= n900;
    P1_REG2_REG_29_ <= n905;
    P1_REG2_REG_30_ <= n910;
    P1_REG2_REG_31_ <= n915;
    P1_ADDR_REG_19_ <= n920;
    P1_ADDR_REG_18_ <= n925;
    P1_ADDR_REG_17_ <= n930;
    P1_ADDR_REG_16_ <= n935;
    P1_ADDR_REG_15_ <= n940;
    P1_ADDR_REG_14_ <= n945;
    P1_ADDR_REG_13_ <= n950;
    P1_ADDR_REG_12_ <= n955;
    P1_ADDR_REG_11_ <= n960;
    P1_ADDR_REG_10_ <= n965;
    P1_ADDR_REG_9_ <= n970;
    P1_ADDR_REG_8_ <= n975;
    P1_ADDR_REG_7_ <= n980;
    P1_ADDR_REG_6_ <= n985;
    P1_ADDR_REG_5_ <= n990;
    P1_ADDR_REG_4_ <= n995;
    P1_ADDR_REG_3_ <= n1000;
    P1_ADDR_REG_2_ <= n1005;
    P1_ADDR_REG_1_ <= n1010;
    P1_ADDR_REG_0_ <= n1015;
    P1_DATAO_REG_0_ <= n1020;
    P1_DATAO_REG_1_ <= n1025;
    P1_DATAO_REG_2_ <= n1030;
    P1_DATAO_REG_3_ <= n1035;
    P1_DATAO_REG_4_ <= n1040;
    P1_DATAO_REG_5_ <= n1045;
    P1_DATAO_REG_6_ <= n1050;
    P1_DATAO_REG_7_ <= n1055;
    P1_DATAO_REG_8_ <= n1060;
    P1_DATAO_REG_9_ <= n1065;
    P1_DATAO_REG_10_ <= n1070;
    P1_DATAO_REG_11_ <= n1075;
    P1_DATAO_REG_12_ <= n1080;
    P1_DATAO_REG_13_ <= n1085;
    P1_DATAO_REG_14_ <= n1090;
    P1_DATAO_REG_15_ <= n1095;
    P1_DATAO_REG_16_ <= n1100;
    P1_DATAO_REG_17_ <= n1105;
    P1_DATAO_REG_18_ <= n1110;
    P1_DATAO_REG_19_ <= n1115;
    P1_DATAO_REG_20_ <= n1120;
    P1_DATAO_REG_21_ <= n1125;
    P1_DATAO_REG_22_ <= n1130;
    P1_DATAO_REG_23_ <= n1135;
    P1_DATAO_REG_24_ <= n1140;
    P1_DATAO_REG_25_ <= n1145;
    P1_DATAO_REG_26_ <= n1150;
    P1_DATAO_REG_27_ <= n1155;
    P1_DATAO_REG_28_ <= n1160;
    P1_DATAO_REG_29_ <= n1165;
    P1_DATAO_REG_30_ <= n1170;
    P1_DATAO_REG_31_ <= n1175;
    P1_B_REG <= n1180;
    P1_REG3_REG_15_ <= n1185;
    P1_REG3_REG_26_ <= n1190;
    P1_REG3_REG_6_ <= n1195;
    P1_REG3_REG_18_ <= n1200;
    P1_REG3_REG_2_ <= n1205;
    P1_REG3_REG_11_ <= n1210;
    P1_REG3_REG_22_ <= n1215;
    P1_REG3_REG_13_ <= n1220;
    P1_REG3_REG_20_ <= n1225;
    P1_REG3_REG_0_ <= n1230;
    P1_REG3_REG_9_ <= n1235;
    P1_REG3_REG_4_ <= n1240;
    P1_REG3_REG_24_ <= n1245;
    P1_REG3_REG_17_ <= n1250;
    P1_REG3_REG_5_ <= n1255;
    P1_REG3_REG_16_ <= n1260;
    P1_REG3_REG_25_ <= n1265;
    P1_REG3_REG_12_ <= n1270;
    P1_REG3_REG_21_ <= n1275;
    P1_REG3_REG_1_ <= n1280;
    P1_REG3_REG_8_ <= n1285;
    P1_REG3_REG_28_ <= n1290;
    P1_REG3_REG_19_ <= n1295;
    P1_REG3_REG_3_ <= n1300;
    P1_REG3_REG_10_ <= n1305;
    P1_REG3_REG_23_ <= n1310;
    P1_REG3_REG_14_ <= n1315;
    P1_REG3_REG_27_ <= n1320;
    P1_REG3_REG_7_ <= n1325;
    P1_STATE_REG <= n1330;
    P1_RD_REG <= n1335;
    P1_WR_REG <= n1340;
    P2_IR_REG_0_ <= n1345;
    P2_IR_REG_1_ <= n1350;
    P2_IR_REG_2_ <= n1355;
    P2_IR_REG_3_ <= n1360;
    P2_IR_REG_4_ <= n1365;
    P2_IR_REG_5_ <= n1370;
    P2_IR_REG_6_ <= n1375;
    P2_IR_REG_7_ <= n1380;
    P2_IR_REG_8_ <= n1385;
    P2_IR_REG_9_ <= n1390;
    P2_IR_REG_10_ <= n1395;
    P2_IR_REG_11_ <= n1400;
    P2_IR_REG_12_ <= n1405;
    P2_IR_REG_13_ <= n1410;
    P2_IR_REG_14_ <= n1415;
    P2_IR_REG_15_ <= n1420;
    P2_IR_REG_16_ <= n1425;
    P2_IR_REG_17_ <= n1430;
    P2_IR_REG_18_ <= n1435;
    P2_IR_REG_19_ <= n1440;
    P2_IR_REG_20_ <= n1445;
    P2_IR_REG_21_ <= n1450;
    P2_IR_REG_22_ <= n1455;
    P2_IR_REG_23_ <= n1460;
    P2_IR_REG_24_ <= n1465;
    P2_IR_REG_25_ <= n1470;
    P2_IR_REG_26_ <= n1475;
    P2_IR_REG_27_ <= n1480;
    P2_IR_REG_28_ <= n1485;
    P2_IR_REG_29_ <= n1490;
    P2_IR_REG_30_ <= n1495;
    P2_IR_REG_31_ <= n1500;
    P2_D_REG_0_ <= n1505;
    P2_D_REG_1_ <= n1510;
    P2_D_REG_2_ <= n1515;
    P2_D_REG_3_ <= n1520;
    P2_D_REG_4_ <= n1525;
    P2_D_REG_5_ <= n1530;
    P2_D_REG_6_ <= n1535;
    P2_D_REG_7_ <= n1540;
    P2_D_REG_8_ <= n1545;
    P2_D_REG_9_ <= n1550;
    P2_D_REG_10_ <= n1555;
    P2_D_REG_11_ <= n1560;
    P2_D_REG_12_ <= n1565;
    P2_D_REG_13_ <= n1570;
    P2_D_REG_14_ <= n1575;
    P2_D_REG_15_ <= n1580;
    P2_D_REG_16_ <= n1585;
    P2_D_REG_17_ <= n1590;
    P2_D_REG_18_ <= n1595;
    P2_D_REG_19_ <= n1600;
    P2_D_REG_20_ <= n1605;
    P2_D_REG_21_ <= n1610;
    P2_D_REG_22_ <= n1615;
    P2_D_REG_23_ <= n1620;
    P2_D_REG_24_ <= n1625;
    P2_D_REG_25_ <= n1630;
    P2_D_REG_26_ <= n1635;
    P2_D_REG_27_ <= n1640;
    P2_D_REG_28_ <= n1645;
    P2_D_REG_29_ <= n1650;
    P2_D_REG_30_ <= n1655;
    P2_D_REG_31_ <= n1660;
    P2_REG0_REG_0_ <= n1665;
    P2_REG0_REG_1_ <= n1670;
    P2_REG0_REG_2_ <= n1675;
    P2_REG0_REG_3_ <= n1680;
    P2_REG0_REG_4_ <= n1685;
    P2_REG0_REG_5_ <= n1690;
    P2_REG0_REG_6_ <= n1695;
    P2_REG0_REG_7_ <= n1700;
    P2_REG0_REG_8_ <= n1705;
    P2_REG0_REG_9_ <= n1710;
    P2_REG0_REG_10_ <= n1715;
    P2_REG0_REG_11_ <= n1720;
    P2_REG0_REG_12_ <= n1725;
    P2_REG0_REG_13_ <= n1730;
    P2_REG0_REG_14_ <= n1735;
    P2_REG0_REG_15_ <= n1740;
    P2_REG0_REG_16_ <= n1745;
    P2_REG0_REG_17_ <= n1750;
    P2_REG0_REG_18_ <= n1755;
    P2_REG0_REG_19_ <= n1760;
    P2_REG0_REG_20_ <= n1765;
    P2_REG0_REG_21_ <= n1770;
    P2_REG0_REG_22_ <= n1775;
    P2_REG0_REG_23_ <= n1780;
    P2_REG0_REG_24_ <= n1785;
    P2_REG0_REG_25_ <= n1790;
    P2_REG0_REG_26_ <= n1795;
    P2_REG0_REG_27_ <= n1800;
    P2_REG0_REG_28_ <= n1805;
    P2_REG0_REG_29_ <= n1810;
    P2_REG0_REG_30_ <= n1815;
    P2_REG0_REG_31_ <= n1820;
    P2_REG1_REG_0_ <= n1825;
    P2_REG1_REG_1_ <= n1830;
    P2_REG1_REG_2_ <= n1835;
    P2_REG1_REG_3_ <= n1840;
    P2_REG1_REG_4_ <= n1845;
    P2_REG1_REG_5_ <= n1850;
    P2_REG1_REG_6_ <= n1855;
    P2_REG1_REG_7_ <= n1860;
    P2_REG1_REG_8_ <= n1865;
    P2_REG1_REG_9_ <= n1870;
    P2_REG1_REG_10_ <= n1875;
    P2_REG1_REG_11_ <= n1880;
    P2_REG1_REG_12_ <= n1885;
    P2_REG1_REG_13_ <= n1890;
    P2_REG1_REG_14_ <= n1895;
    P2_REG1_REG_15_ <= n1900;
    P2_REG1_REG_16_ <= n1905;
    P2_REG1_REG_17_ <= n1910;
    P2_REG1_REG_18_ <= n1915;
    P2_REG1_REG_19_ <= n1920;
    P2_REG1_REG_20_ <= n1925;
    P2_REG1_REG_21_ <= n1930;
    P2_REG1_REG_22_ <= n1935;
    P2_REG1_REG_23_ <= n1940;
    P2_REG1_REG_24_ <= n1945;
    P2_REG1_REG_25_ <= n1950;
    P2_REG1_REG_26_ <= n1955;
    P2_REG1_REG_27_ <= n1960;
    P2_REG1_REG_28_ <= n1965;
    P2_REG1_REG_29_ <= n1970;
    P2_REG1_REG_30_ <= n1975;
    P2_REG1_REG_31_ <= n1980;
    P2_REG2_REG_0_ <= n1985;
    P2_REG2_REG_1_ <= n1990;
    P2_REG2_REG_2_ <= n1995;
    P2_REG2_REG_3_ <= n2000;
    P2_REG2_REG_4_ <= n2005;
    P2_REG2_REG_5_ <= n2010;
    P2_REG2_REG_6_ <= n2015;
    P2_REG2_REG_7_ <= n2020;
    P2_REG2_REG_8_ <= n2025;
    P2_REG2_REG_9_ <= n2030;
    P2_REG2_REG_10_ <= n2035;
    P2_REG2_REG_11_ <= n2040;
    P2_REG2_REG_12_ <= n2045;
    P2_REG2_REG_13_ <= n2050;
    P2_REG2_REG_14_ <= n2055;
    P2_REG2_REG_15_ <= n2060;
    P2_REG2_REG_16_ <= n2065;
    P2_REG2_REG_17_ <= n2070;
    P2_REG2_REG_18_ <= n2075;
    P2_REG2_REG_19_ <= n2080;
    P2_REG2_REG_20_ <= n2085;
    P2_REG2_REG_21_ <= n2090;
    P2_REG2_REG_22_ <= n2095;
    P2_REG2_REG_23_ <= n2100;
    P2_REG2_REG_24_ <= n2105;
    P2_REG2_REG_25_ <= n2110;
    P2_REG2_REG_26_ <= n2115;
    P2_REG2_REG_27_ <= n2120;
    P2_REG2_REG_28_ <= n2125;
    P2_REG2_REG_29_ <= n2130;
    P2_REG2_REG_30_ <= n2135;
    P2_REG2_REG_31_ <= n2140;
    P2_ADDR_REG_19_ <= n2145;
    P2_ADDR_REG_18_ <= n2150;
    P2_ADDR_REG_17_ <= n2155;
    P2_ADDR_REG_16_ <= n2160;
    P2_ADDR_REG_15_ <= n2165;
    P2_ADDR_REG_14_ <= n2170;
    P2_ADDR_REG_13_ <= n2175;
    P2_ADDR_REG_12_ <= n2180;
    P2_ADDR_REG_11_ <= n2185;
    P2_ADDR_REG_10_ <= n2190;
    P2_ADDR_REG_9_ <= n2195;
    P2_ADDR_REG_8_ <= n2200;
    P2_ADDR_REG_7_ <= n2205;
    P2_ADDR_REG_6_ <= n2210;
    P2_ADDR_REG_5_ <= n2215;
    P2_ADDR_REG_4_ <= n2220;
    P2_ADDR_REG_3_ <= n2225;
    P2_ADDR_REG_2_ <= n2230;
    P2_ADDR_REG_1_ <= n2235;
    P2_ADDR_REG_0_ <= n2240;
    P2_DATAO_REG_0_ <= n2245;
    P2_DATAO_REG_1_ <= n2250;
    P2_DATAO_REG_2_ <= n2255;
    P2_DATAO_REG_3_ <= n2260;
    P2_DATAO_REG_4_ <= n2265;
    P2_DATAO_REG_5_ <= n2270;
    P2_DATAO_REG_6_ <= n2275;
    P2_DATAO_REG_7_ <= n2280;
    P2_DATAO_REG_8_ <= n2285;
    P2_DATAO_REG_9_ <= n2290;
    P2_DATAO_REG_10_ <= n2295;
    P2_DATAO_REG_11_ <= n2300;
    P2_DATAO_REG_12_ <= n2305;
    P2_DATAO_REG_13_ <= n2310;
    P2_DATAO_REG_14_ <= n2315;
    P2_DATAO_REG_15_ <= n2320;
    P2_DATAO_REG_16_ <= n2325;
    P2_DATAO_REG_17_ <= n2330;
    P2_DATAO_REG_18_ <= n2335;
    P2_DATAO_REG_19_ <= n2340;
    P2_DATAO_REG_20_ <= n2345;
    P2_DATAO_REG_21_ <= n2350;
    P2_DATAO_REG_22_ <= n2355;
    P2_DATAO_REG_23_ <= n2360;
    P2_DATAO_REG_24_ <= n2365;
    P2_DATAO_REG_25_ <= n2370;
    P2_DATAO_REG_26_ <= n2375;
    P2_DATAO_REG_27_ <= n2380;
    P2_DATAO_REG_28_ <= n2385;
    P2_DATAO_REG_29_ <= n2390;
    P2_DATAO_REG_30_ <= n2395;
    P2_DATAO_REG_31_ <= n2400;
    P2_B_REG <= n2405;
    P2_REG3_REG_15_ <= n2410;
    P2_REG3_REG_26_ <= n2415;
    P2_REG3_REG_6_ <= n2420;
    P2_REG3_REG_18_ <= n2425;
    P2_REG3_REG_2_ <= n2430;
    P2_REG3_REG_11_ <= n2435;
    P2_REG3_REG_22_ <= n2440;
    P2_REG3_REG_13_ <= n2445;
    P2_REG3_REG_20_ <= n2450;
    P2_REG3_REG_0_ <= n2455;
    P2_REG3_REG_9_ <= n2460;
    P2_REG3_REG_4_ <= n2465;
    P2_REG3_REG_24_ <= n2470;
    P2_REG3_REG_17_ <= n2475;
    P2_REG3_REG_5_ <= n2480;
    P2_REG3_REG_16_ <= n2485;
    P2_REG3_REG_25_ <= n2490;
    P2_REG3_REG_12_ <= n2495;
    P2_REG3_REG_21_ <= n2500;
    P2_REG3_REG_1_ <= n2505;
    P2_REG3_REG_8_ <= n2510;
    P2_REG3_REG_28_ <= n2515;
    P2_REG3_REG_19_ <= n2520;
    P2_REG3_REG_3_ <= n2525;
    P2_REG3_REG_10_ <= n2530;
    P2_REG3_REG_23_ <= n2535;
    P2_REG3_REG_14_ <= n2540;
    P2_REG3_REG_27_ <= n2545;
    P2_REG3_REG_7_ <= n2550;
    P2_STATE_REG <= n2555;
    P2_RD_REG <= n2560;
    P2_WR_REG <= n2565;
    Q_0 <= n41480;
    Q_1 <= n41483;
    Q_2 <= n41486;
    Q_3 <= n41489;
  end
endmodule
