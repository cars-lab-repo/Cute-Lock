library ieee;
use ieee.std_logic_1164.all;

entity micks is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20,x21 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y39,y40,y41,y42,y43,y45 : out std_logic );
end micks;

architecture ARC of micks is

   type states_micks is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22 );
   signal current_micks : states_micks;

begin
   process (clk , rst)
   procedure proc_micks is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y45  <= '0' ;


   case current_micks is
   when s1 =>
      if ( x1 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_micks <= s2;

      elsif ( x1 and not x2 ) = '1' then
         y1 <= '1' ;
         current_micks <= s3;

      else
         current_micks <= s1;

      end if;

   when s2 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         current_micks <= s4;

   when s3 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_micks <= s5;

   when s4 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_micks <= s6;

   when s5 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_micks <= s7;

   when s6 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s8;

   when s7 =>
      if ( x15 and x21 and x20 and x4 and x6 ) = '1' then
         y18 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and x20 and x4 and not x6 ) = '1' then
         y38 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and x20 and not x4 and x5 and x6 and x9 ) = '1' then
         y9 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and not x8 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and x20 and not x4 and x5 and x6 and not x9 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and x20 and not x4 and x5 and not x6 and x8 ) = '1' then
         y9 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and x20 and not x4 and x5 and not x6 and not x8 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and x20 and not x4 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and x20 and not x4 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y40 <= '1' ;
         y42 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and x18 and x4 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_micks <= s10;

      elsif ( x15 and x21 and not x20 and x18 and x4 and x5 and not x6 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_micks <= s11;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and x6 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and x6 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and x6 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and x6 and not x11 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and not x6 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and not x6 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and not x6 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and x4 and not x5 and not x6 and not x10 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and x6 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and x6 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and x6 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and x6 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and x6 and not x13 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and not x6 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and not x6 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and not x6 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and not x6 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and x5 and not x6 and not x14 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and x18 and not x4 and not x5 and not x6 ) = '1' then
         y35 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and x21 and not x20 and not x18 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_micks <= s12;

      elsif ( x15 and not x21 and x18 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y29 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and not x21 and x18 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and not x21 and x18 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y10 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_micks <= s13;

      elsif ( x15 and not x21 and x18 and not x20 and x4 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and not x21 and x18 and not x20 and not x4 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( x15 and not x21 and not x18 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_micks <= s12;

      else
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_micks <= s14;

      end if;

   when s8 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_micks <= s1;

   when s9 =>
      if ( x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      else
         current_micks <= s1;

      end if;

   when s10 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y37 <= '1' ;
         current_micks <= s15;

   when s11 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

   when s12 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_micks <= s16;

      elsif ( not x3 and x19 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_micks <= s17;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_micks <= s10;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x5 and not x6 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_micks <= s11;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and x6 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and not x6 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x5 and not x6 ) = '1' then
         y35 <= '1' ;
         current_micks <= s9;

      elsif ( not x3 and x19 and not x20 and not x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_micks <= s18;

      end if;

   when s13 =>
      if ( x7 ) = '1' then
         y31 <= '1' ;
         y32 <= '1' ;
         current_micks <= s9;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      else
         current_micks <= s1;

      end if;

   when s14 =>
      if ( x16 ) = '1' then
         y12 <= '1' ;
         current_micks <= s3;

      elsif ( not x16 and x21 and x20 and x4 and x6 ) = '1' then
         y18 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and x21 and x20 and x4 and not x6 ) = '1' then
         y38 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and x6 and x9 ) = '1' then
         y9 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and not x8 ) = '1' then
         current_micks <= s1;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and x6 and not x9 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and not x6 and x8 ) = '1' then
         y9 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x16 and x21 and x20 and not x4 and x5 and not x6 and not x8 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x16 and x21 and x20 and not x4 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and x21 and x20 and not x4 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y40 <= '1' ;
         y42 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and x21 and not x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_micks <= s18;

      elsif ( not x16 and not x21 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_micks <= s18;

      elsif ( not x16 and not x21 and not x3 and x4 and x5 and x20 and x6 ) = '1' then
         y28 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and x4 and x5 and x20 and not x6 ) = '1' then
         y26 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and x4 and x5 and not x20 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and x4 and not x5 and x20 and x6 ) = '1' then
         y27 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and x4 and not x5 and x20 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y23 <= '1' ;
         current_micks <= s19;

      elsif ( not x16 and not x21 and not x3 and x4 and not x5 and not x20 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and not x4 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and not x4 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( not x16 and not x21 and not x3 and not x4 and x20 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y30 <= '1' ;
         y45 <= '1' ;
         current_micks <= s20;

      elsif ( not x16 and not x21 and not x3 and not x4 and x20 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y20 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_micks <= s21;

      else
         y5 <= '1' ;
         y20 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      end if;

   when s15 =>
      if ( x12 ) = '1' then
         y9 <= '1' ;
         current_micks <= s9;

      elsif ( not x12 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x12 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x12 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      else
         current_micks <= s1;

      end if;

   when s16 =>
      if ( x19 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_micks <= s17;

      elsif ( x19 and not x20 and x4 and x21 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_micks <= s10;

      elsif ( x19 and not x20 and x4 and x21 and x5 and not x6 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_micks <= s11;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and x6 and not x11 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and x21 and not x5 and not x6 and not x10 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and x6 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and x6 and not x13 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and not x6 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and x5 and not x6 and not x14 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( x19 and not x20 and not x4 and x21 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and not x4 and x21 and not x5 and not x6 ) = '1' then
         y35 <= '1' ;
         current_micks <= s9;

      elsif ( x19 and not x20 and not x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_micks <= s18;

      end if;

   when s17 =>
      if ( x7 ) = '1' then
         y31 <= '1' ;
         y32 <= '1' ;
         current_micks <= s9;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      else
         current_micks <= s1;

      end if;

   when s18 =>
      if ( x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_micks <= s9;

      elsif ( x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_micks <= s17;

      elsif ( not x20 and x4 and x21 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_micks <= s10;

      elsif ( not x20 and x4 and x21 and x5 and not x6 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_micks <= s11;

      elsif ( not x20 and x4 and x21 and not x5 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and x6 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and x6 and not x11 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and not x6 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and x4 and x21 and not x5 and not x6 and not x10 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      elsif ( not x20 and not x4 and x21 and x5 and x6 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and x6 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and x6 and not x13 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and not x6 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and not x6 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and x5 and not x6 and not x14 and not x17 ) = '1' then
         current_micks <= s1;

      elsif ( not x20 and not x4 and x21 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_micks <= s9;

      elsif ( not x20 and not x4 and x21 and not x5 and not x6 ) = '1' then
         y35 <= '1' ;
         current_micks <= s9;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_micks <= s9;

      end if;

   when s19 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_micks <= s22;

   when s20 =>
      if ( x7 ) = '1' then
         y33 <= '1' ;
         y34 <= '1' ;
         current_micks <= s9;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      else
         current_micks <= s1;

      end if;

   when s21 =>
      if ( x7 ) = '1' then
         y31 <= '1' ;
         y32 <= '1' ;
         current_micks <= s9;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_micks <= s1;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_micks <= s1;

      else
         current_micks <= s1;

      end if;

   when s22 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_micks <= s9;

   end case;
   end proc_micks;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y45  <= '0' ;

	current_micks <= s1;
      elsif (clk'event and clk ='1') then
        proc_micks;
      end if;
   end process;
end ARC;
