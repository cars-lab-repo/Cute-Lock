library ieee;
use ieee.std_logic_1164.all;

entity proc41616 is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y39,y40,y41,y42,y43,y44,y45,
	y46,y47 : out std_logic );
end proc41616;

architecture ARC of proc41616 is

   type states_proc41616 is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
	s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,
	s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57 );
   signal current_proc41616 : states_proc41616;

begin
   process (clk , rst)
   procedure proc_proc41616 is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;	y46  <= '0' ;	y47  <= '0' ;

   case current_proc41616 is
   when s1 =>
      if ( x3 and x5 and x17 and x18 ) = '1' then
         y23 <= '1' ;
         y24 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_proc41616 <= s1;

      elsif ( x3 and x5 and x17 and not x18 ) = '1' then
         y33 <= '1' ;
         y35 <= '1' ;
         current_proc41616 <= s1;

      elsif ( x3 and x5 and not x17 and x18 ) = '1' then
         y8 <= '1' ;
         y33 <= '1' ;
         current_proc41616 <= s1;

      elsif ( x3 and x5 and not x17 and not x18 ) = '1' then
         y23 <= '1' ;
         y33 <= '1' ;
         current_proc41616 <= s1;

      elsif ( x3 and not x5 and x6 ) = '1' then
         y7 <= '1' ;
         y24 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_proc41616 <= s2;

      elsif ( x3 and not x5 and not x6 ) = '1' then
         y32 <= '1' ;
         y39 <= '1' ;
         current_proc41616 <= s3;

      else
         current_proc41616 <= s1;

      end if;

   when s2 =>
         y7 <= '1' ;
         y25 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_proc41616 <= s1;

   when s3 =>
         y26 <= '1' ;
         current_proc41616 <= s4;

   when s4 =>
      if ( x12 and x14 and x13 and x16 ) = '1' then
         y30 <= '1' ;
         current_proc41616 <= s5;

      elsif ( x12 and x14 and x13 and not x16 ) = '1' then
         y29 <= '1' ;
         current_proc41616 <= s5;

      elsif ( x12 and x14 and not x13 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s6;

      elsif ( x12 and not x14 and x13 and x15 and x16 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s6;

      elsif ( x12 and not x14 and x13 and x15 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y27 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s7;

      elsif ( x12 and not x14 and x13 and not x15 and x16 and x11 ) = '1' then
         y26 <= '1' ;
         current_proc41616 <= s8;

      elsif ( x12 and not x14 and x13 and not x15 and x16 and not x11 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( x12 and not x14 and x13 and not x15 and x16 and not x11 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( x12 and not x14 and x13 and not x15 and x16 and not x11 and not x19 and not x10 ) = '1' then
         current_proc41616 <= s1;

      elsif ( x12 and not x14 and x13 and not x15 and not x16 and x10 ) = '1' then
         y26 <= '1' ;
         current_proc41616 <= s8;

      elsif ( x12 and not x14 and x13 and not x15 and not x16 and not x10 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( x12 and not x14 and x13 and not x15 and not x16 and not x10 and not x19 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( x12 and not x14 and x13 and not x15 and not x16 and not x10 and not x19 and not x11 ) = '1' then
         current_proc41616 <= s1;

      elsif ( x12 and not x14 and not x13 and x15 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s6;

      elsif ( x12 and not x14 and not x13 and not x15 and x1 ) = '1' then
         y19 <= '1' ;
         y23 <= '1' ;
         y32 <= '1' ;
         current_proc41616 <= s9;

      elsif ( x12 and not x14 and not x13 and not x15 and not x1 and x16 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s6;

      elsif ( x12 and not x14 and not x13 and not x15 and not x1 and not x16 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      elsif ( not x12 and x1 ) = '1' then
         y19 <= '1' ;
         y23 <= '1' ;
         y32 <= '1' ;
         current_proc41616 <= s9;

      elsif ( not x12 and not x1 and x13 and x15 and x16 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      elsif ( not x12 and not x1 and x13 and x15 and not x16 and x9 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      elsif ( not x12 and not x1 and x13 and x15 and not x16 and not x9 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and x15 and not x16 and not x9 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and x15 and not x16 and not x9 and not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and x15 and not x16 and not x9 and not x19 and not x10 and not x11 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and x16 and x8 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      elsif ( not x12 and not x1 and x13 and not x15 and x16 and not x8 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and x16 and not x8 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and x16 and not x8 and not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and x16 and not x8 and not x19 and not x10 and not x11 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and not x16 and x7 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      elsif ( not x12 and not x1 and x13 and not x15 and not x16 and not x7 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and not x16 and not x7 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and not x16 and not x7 and not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and not x1 and x13 and not x15 and not x16 and not x7 and not x19 and not x10 and not x11 ) = '1' then
         current_proc41616 <= s1;

      else
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      end if;

   when s5 =>
      if ( x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      else
         current_proc41616 <= s1;

      end if;

   when s6 =>
      if ( x15 and x13 ) = '1' then
         y3 <= '1' ;
         current_proc41616 <= s11;

      elsif ( x15 and not x13 ) = '1' then
         y3 <= '1' ;
         current_proc41616 <= s12;

      elsif ( not x15 and x14 and x13 ) = '1' then
         y3 <= '1' ;
         current_proc41616 <= s11;

      elsif ( not x15 and x14 and not x13 ) = '1' then
         y3 <= '1' ;
         current_proc41616 <= s12;

      else
         y3 <= '1' ;
         current_proc41616 <= s11;

      end if;

   when s7 =>
         y2 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s13;

   when s8 =>
         y26 <= '1' ;
         current_proc41616 <= s5;

   when s9 =>
         y26 <= '1' ;
         current_proc41616 <= s14;

   when s10 =>
      if ( x16 and x12 ) = '1' then
         y2 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s13;

      elsif ( x16 and not x12 ) = '1' then
         y3 <= '1' ;
         current_proc41616 <= s15;

      else
         y3 <= '1' ;
         current_proc41616 <= s15;

      end if;

   when s11 =>
         y37 <= '1' ;
         current_proc41616 <= s16;

   when s12 =>
         y37 <= '1' ;
         current_proc41616 <= s17;

   when s13 =>
         y37 <= '1' ;
         current_proc41616 <= s18;

   when s14 =>
      if ( x12 and x4 and x16 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( x12 and x4 and x16 and not x2 and x20 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( x12 and x4 and x16 and not x2 and not x20 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      elsif ( x12 and x4 and not x16 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s19;

      elsif ( x12 and not x4 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( x12 and not x4 and not x2 and x20 and x16 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( x12 and not x4 and not x2 and x20 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      elsif ( x12 and not x4 and not x2 and not x20 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      elsif ( not x12 and x13 and x15 and x16 and x4 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and x15 and x16 and not x4 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( not x12 and x13 and x15 and x16 and not x4 and not x2 and x20 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and x15 and x16 and not x4 and not x2 and not x20 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and x4 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and not x4 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and not x4 and not x2 and x20 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and not x4 and not x2 and not x20 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and not x19 and not x10 and not x11 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and x4 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and not x4 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and not x4 and not x2 and x20 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and not x4 and not x2 and not x20 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and not x19 and not x10 and not x11 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and x4 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and not x4 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and not x4 and not x2 and x20 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and not x4 and not x2 and not x20 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and x19 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and not x19 and x10 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and not x19 and not x10 and x11 ) = '1' then
         y40 <= '1' ;
         current_proc41616 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and not x19 and not x10 and not x11 ) = '1' then
         current_proc41616 <= s1;

      elsif ( not x12 and not x13 and x4 and x14 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s19;

      elsif ( not x12 and not x13 and x4 and not x14 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( not x12 and not x13 and not x4 and x2 ) = '1' then
         y38 <= '1' ;
         current_proc41616 <= s20;

      elsif ( not x12 and not x13 and not x4 and not x2 and x20 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      else
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      end if;

   when s15 =>
         y37 <= '1' ;
         current_proc41616 <= s24;

   when s16 =>
         y42 <= '1' ;
         current_proc41616 <= s25;

   when s17 =>
         y42 <= '1' ;
         current_proc41616 <= s26;

   when s18 =>
         y10 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s27;

   when s19 =>
      if ( x12 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      else
         y7 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_proc41616 <= s28;

      end if;

   when s20 =>
         y8 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y34 <= '1' ;
         current_proc41616 <= s29;

   when s21 =>
      if ( x12 and x16 ) = '1' then
         y3 <= '1' ;
         current_proc41616 <= s12;

      elsif ( x12 and not x16 ) = '1' then
         y2 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s13;

      else
         y3 <= '1' ;
         current_proc41616 <= s11;

      end if;

   when s22 =>
      if ( x12 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( not x12 and x14 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_proc41616 <= s28;

      else
         y19 <= '1' ;
         current_proc41616 <= s30;

      end if;

   when s23 =>
         y2 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s31;

   when s24 =>
         y42 <= '1' ;
         current_proc41616 <= s32;

   when s25 =>
         y37 <= '1' ;
         current_proc41616 <= s33;

   when s26 =>
         y37 <= '1' ;
         current_proc41616 <= s34;

   when s27 =>
         y37 <= '1' ;
         current_proc41616 <= s35;

   when s28 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s7;

   when s29 =>
      if ( x20 and x12 and x16 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( x20 and x12 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      elsif ( x20 and not x12 and x13 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( x20 and not x12 and not x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      else
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s23;

      end if;

   when s30 =>
         y9 <= '1' ;
         current_proc41616 <= s21;

   when s31 =>
         y37 <= '1' ;
         current_proc41616 <= s36;

   when s32 =>
         y37 <= '1' ;
         current_proc41616 <= s37;

   when s33 =>
         y43 <= '1' ;
         current_proc41616 <= s38;

   when s34 =>
         y43 <= '1' ;
         current_proc41616 <= s39;

   when s35 =>
         y1 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s40;

   when s36 =>
         y10 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s41;

   when s37 =>
         y43 <= '1' ;
         current_proc41616 <= s42;

   when s38 =>
         y37 <= '1' ;
         current_proc41616 <= s43;

   when s39 =>
         y37 <= '1' ;
         current_proc41616 <= s44;

   when s40 =>
         y37 <= '1' ;
         current_proc41616 <= s45;

   when s41 =>
         y37 <= '1' ;
         current_proc41616 <= s46;

   when s42 =>
         y37 <= '1' ;
         current_proc41616 <= s47;

   when s43 =>
         y44 <= '1' ;
         current_proc41616 <= s48;

   when s44 =>
         y44 <= '1' ;
         current_proc41616 <= s49;

   when s45 =>
         y36 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s5;

   when s46 =>
         y1 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s50;

   when s47 =>
         y44 <= '1' ;
         current_proc41616 <= s51;

   when s48 =>
      if ( x12 and x13 ) = '1' then
         y28 <= '1' ;
         y45 <= '1' ;
         current_proc41616 <= s5;

      elsif ( x12 and not x13 and x2 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y9 <= '1' ;
         current_proc41616 <= s52;

      elsif ( x12 and not x13 and not x2 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         current_proc41616 <= s10;

      else
         y14 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_proc41616 <= s28;

      end if;

   when s49 =>
      if ( x15 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_proc41616 <= s28;

      elsif ( not x15 and x14 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_proc41616 <= s28;

      else
         y24 <= '1' ;
         current_proc41616 <= s5;

      end if;

   when s50 =>
         y37 <= '1' ;
         current_proc41616 <= s53;

   when s51 =>
      if ( x12 and x16 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_proc41616 <= s5;

      elsif ( x12 and not x16 and x2 ) = '1' then
         y19 <= '1' ;
         current_proc41616 <= s54;

      elsif ( x12 and not x16 and not x2 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( not x12 and x13 ) = '1' then
         y7 <= '1' ;
         y25 <= '1' ;
         current_proc41616 <= s5;

      elsif ( not x12 and not x13 and x2 and x14 ) = '1' then
         y19 <= '1' ;
         current_proc41616 <= s54;

      elsif ( not x12 and not x13 and x2 and not x14 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         y19 <= '1' ;
         current_proc41616 <= s30;

      elsif ( not x12 and not x13 and not x2 and x14 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_proc41616 <= s28;

      else
         y19 <= '1' ;
         current_proc41616 <= s54;

      end if;

   when s52 =>
         y3 <= '1' ;
         current_proc41616 <= s15;

   when s53 =>
         y36 <= '1' ;
         y41 <= '1' ;
         current_proc41616 <= s55;

   when s54 =>
      if ( x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      elsif ( not x14 and x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      else
         y9 <= '1' ;
         current_proc41616 <= s21;

      end if;

   when s55 =>
         y47 <= '1' ;
         y46 <= '1' ;
         current_proc41616 <= s56;

   when s56 =>
         y8 <= '1' ;
         y19 <= '1' ;
         y34 <= '1' ;
         current_proc41616 <= s57;

   when s57 =>
      if ( x12 and x16 ) = '1' then
         y9 <= '1' ;
         current_proc41616 <= s21;

      elsif ( x12 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      elsif ( not x12 and x13 ) = '1' then
         y25 <= '1' ;
         current_proc41616 <= s5;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y42 <= '1' ;
         y5 <= '1' ;
         y43 <= '1' ;
         y6 <= '1' ;
         y44 <= '1' ;
         current_proc41616 <= s22;

      end if;

   end case;
   end proc_proc41616;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;	y46  <= '0' ;	y47  <= '0' ;
	current_proc41616 <= s1;
      elsif (clk'event and clk ='1') then
        proc_proc41616;
      end if;
   end process;
end ARC;
