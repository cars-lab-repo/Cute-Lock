library ieee;
use ieee.std_logic_1164.all;

entity otherm is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,
	x31,x32,x33,x34,x35,x36,x37,x38,x39,x40,x41,x42,x43,x44,x45,
	x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,
	x61,x62,x63,x64,x65,x66,x67 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y39,y40,y41,y42,y43,y44,y45,
	y46,y47,y48,y49,y50,y51,y52,y53,y54,y55,y56,y57,y58,y59,y60,
	y61,y62,y63,y64,y65,y66,y67,y68,y69,y70,y71,y72,y73,y74,y75,
	y77,y78,y79,y80,y81,y84,y86,y88,y90,y91,y92,y93,y94,y95,y96,
	y97,y98,y99,y100,y102,y110 : out std_logic );
end otherm;

architecture ARC of otherm is

   type states_otherm is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
	s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,
	s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,
	s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,
	s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,
	s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,
	s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,
	s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,
	s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,
	s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,
	s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,
	s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,
	s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,
	s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,
	s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,
	s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,
	s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,
	s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,
	s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,
	s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,
	s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,
	s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,
	s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,
	s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,
	s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,
	s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,
	s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,
	s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,s433,s434,s435,
	s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,
	s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,
	s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,s478,s479,s480,
	s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,
	s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,
	s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,s521,s522,s523,s524,s525,
	s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,
	s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,
	s556,s557,s558,s559,s560,s561,s562,s563,s564,s565,s566,s567,s568,s569,s570,
	s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,
	s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,
	s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,
	s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,
	s631,s632,s633,s634,s635,s636,s637,s638,s639,s640,s641,s642,s643,s644,s645,
	s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,
	s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,s673,s674,s675,
	s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,
	s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,
	s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,
	s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,
	s736,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,
	s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,
	s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,
	s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,s793,s794,s795,
	s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,
	s811,s812,s813,s814,s815,s816,s817,s818,s819,s820,s821,s822,s823,s824,s825,
	s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,
	s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,
	s856,s857,s858,s859,s860,s861,s862,s863,s864,s865,s866,s867,s868,s869,s870,
	s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,s881,s882,s883,s884,s885,
	s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,s898,s899,s900,
	s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,s913,s914,s915,
	s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,s926,s927,s928,s929,s930,
	s931,s932,s933,s934,s935,s936,s937,s938,s939,s940,s941,s942,s943,s944,s945,
	s946,s947,s948,s949,s950,s951,s952,s953,s954,s955,s956,s957,s958,s959,s960,
	s961,s962,s963,s964,s965,s966,s967,s968,s969,s970,s971,s972,s973,s974,s975,
	s976,s977,s978,s979,s980,s981,s982,s983,s984,s985,s986,s987,s988,s989,s990,
	s991,s992,s993,s994,s995,s996,s997,s998,s999,s1000,s1001,s1002,s1003,s1004,s1005,
	s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,
	s1021,s1022,s1023,s1024,s1025,s1026,s1027,s1028,s1029,s1030,s1031,s1032,s1033,s1034,s1035,
	s1036,s1037,s1038,s1039,s1040,s1041,s1042,s1043,s1044,s1045,s1046,s1047,s1048,s1049,s1050,
	s1051,s1052,s1053,s1054,s1055,s1056,s1057,s1058,s1059,s1060,s1061,s1062,s1063,s1064,s1065,
	s1066,s1067,s1068,s1069,s1070,s1071,s1072,s1073,s1074,s1075,s1076,s1077,s1078,s1079,s1080,
	s1081,s1082,s1083,s1084,s1085,s1086,s1087,s1088,s1089,s1090,s1091,s1092,s1093,s1094,s1095,
	s1096,s1097,s1098,s1099,s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,
	s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,s1120,s1121,s1122,s1123,s1124,s1125,
	s1126,s1127,s1128,s1129,s1130,s1131,s1132,s1133,s1134,s1135,s1136,s1137,s1138,s1139,s1140,
	s1141,s1142,s1143,s1144,s1145,s1146,s1147,s1148,s1149,s1150,s1151,s1152,s1153,s1154,s1155,
	s1156,s1157,s1158,s1159,s1160,s1161,s1162,s1163,s1164,s1165,s1166,s1167,s1168,s1169,s1170,
	s1171,s1172,s1173,s1174,s1175,s1176,s1177,s1178,s1179,s1180,s1181,s1182,s1183,s1184,s1185,
	s1186,s1187,s1188,s1189,s1190,s1191,s1192,s1193,s1194,s1195,s1196,s1197,s1198,s1199,s1200,
	s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,
	s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224,s1225,s1226,s1227,s1228,s1229,s1230,
	s1231,s1232,s1233,s1234,s1235,s1236,s1237,s1238,s1239,s1240,s1241,s1242,s1243,s1244,s1245,
	s1246,s1247,s1248,s1249,s1250,s1251,s1252,s1253,s1254,s1255,s1256,s1257,s1258,s1259,s1260,
	s1261,s1262,s1263,s1264,s1265,s1266,s1267,s1268,s1269,s1270,s1271,s1272,s1273,s1274,s1275
	 );
   signal current_otherm : states_otherm;

begin
   process (clk , rst)
   procedure proc_otherm is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;	y46  <= '0' ;	y47  <= '0' ;	y48  <= '0' ;
	y49  <= '0' ;	y50  <= '0' ;	y51  <= '0' ;	y52  <= '0' ;
	y53  <= '0' ;	y54  <= '0' ;	y55  <= '0' ;	y56  <= '0' ;
	y57  <= '0' ;	y58  <= '0' ;	y59  <= '0' ;	y60  <= '0' ;
	y61  <= '0' ;	y62  <= '0' ;	y63  <= '0' ;	y64  <= '0' ;
	y65  <= '0' ;	y66  <= '0' ;	y67  <= '0' ;	y68  <= '0' ;
	y69  <= '0' ;	y70  <= '0' ;	y71  <= '0' ;	y72  <= '0' ;
	y73  <= '0' ;	y74  <= '0' ;	y75  <= '0' ;	y77  <= '0' ;
	y78  <= '0' ;	y79  <= '0' ;	y80  <= '0' ;	y81  <= '0' ;
	y84  <= '0' ;	y86  <= '0' ;	y88  <= '0' ;	y90  <= '0' ;
	y91  <= '0' ;	y92  <= '0' ;	y93  <= '0' ;	y94  <= '0' ;
	y95  <= '0' ;	y96  <= '0' ;	y97  <= '0' ;	y98  <= '0' ;
	y99  <= '0' ;	y100 <= '0' ;	y102 <= '0' ;	y110 <= '0' ;


   case current_otherm is
   when s1 =>
      if ( x65 and x62 and x64 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s2;

      elsif ( x65 and x62 and x64 and x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and x62 and x64 and not x2 and x1 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s3;

      elsif ( x65 and x62 and x64 and not x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and x25 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s4;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and x26 and x27 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and x26 and not x27 and x2 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and x26 and not x27 and x2 and not x4 and x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and x26 and not x27 and x2 and not x4 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and x26 and not x27 and not x2 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and x26 and not x27 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and x14 and x12 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and x14 and not x12 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and not x14 and x15 and x12 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and not x14 and x15 and not x12 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and not x14 and not x15 and x16 and x12 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and not x14 and not x15 and x16 and not x12 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and x27 and not x14 and not x15 and not x16 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and not x27 and x12 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x65 and x62 and not x64 and x1 and x66 and x67 and not x25 and not x26 and not x27 and not x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and x62 and not x64 and x1 and x66 and not x67 and x2 ) = '1' then
         y1 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s15;

      elsif ( x65 and x62 and not x64 and x1 and x66 and not x67 and not x2 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x65 and x62 and not x64 and x1 and not x66 and x67 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x65 and x62 and not x64 and x1 and not x66 and not x67 and x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x65 and x62 and not x64 and x1 and not x66 and not x67 and not x2 and x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s19;

      elsif ( x65 and x62 and not x64 and x1 and not x66 and not x67 and not x2 and x3 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x65 and x62 and not x64 and x1 and not x66 and not x67 and not x2 and x3 and not x6 and not x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s19;

      elsif ( x65 and x62 and not x64 and x1 and not x66 and not x67 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x65 and x62 and not x64 and not x1 and x67 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and x62 and not x64 and not x1 and not x67 and x66 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and x62 and not x64 and not x1 and not x67 and not x66 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( x65 and not x62 and x63 and x66 and x67 and x64 and x13 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s22;

      elsif ( x65 and not x62 and x63 and x66 and x67 and x64 and x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and x66 and x67 and x64 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s23;

      elsif ( x65 and not x62 and x63 and x66 and x67 and x64 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and x66 and x67 and not x64 and x1 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x65 and not x62 and x63 and x66 and x67 and not x64 and not x1 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x65 and not x62 and x63 and x66 and not x67 and x64 and x9 and x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and x66 and not x67 and x64 and x9 and not x8 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s25;

      elsif ( x65 and not x62 and x63 and x66 and not x67 and x64 and not x9 and x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and x66 and not x67 and x64 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s26;

      elsif ( x65 and not x62 and x63 and x66 and not x67 and not x64 and x6 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x65 and not x62 and x63 and x66 and not x67 and not x64 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and x15 and x16 and x5 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and x15 and x16 and not x5 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and x15 and x16 and not x5 and not x6 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and x15 and not x16 and x1 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and x15 and not x16 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and not x15 and x1 and x16 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and not x15 and x1 and not x16 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and x67 and not x15 and not x1 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and x18 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and x15 and x10 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and x15 and not x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and x2 and x4 and x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and x2 and x4 and x5 and not x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and x2 and x4 and not x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and x2 and x4 and not x5 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and x2 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and x2 and not x4 and not x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and x1 and not x18 and not x15 and not x2 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and not x1 and x18 and x2 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and not x1 and x18 and not x2 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and not x1 and not x18 and x15 and x6 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and not x1 and not x18 and x15 and not x6 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and x17 and not x1 and not x18 and not x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and x15 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and x15 and not x1 and x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and x15 and not x1 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and x2 and x4 and x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and x2 and x4 and x5 and not x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and x2 and x4 and not x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and x2 and x4 and not x5 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and x2 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and x2 and not x4 and not x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and x1 and not x2 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and x18 and not x15 and not x1 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x65 and not x62 and x63 and not x66 and x64 and not x67 and not x17 and not x18 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( x65 and not x62 and x63 and not x66 and not x64 and x67 and x15 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x65 and not x62 and x63 and not x66 and not x64 and x67 and x15 and not x1 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x65 and not x62 and x63 and not x66 and not x64 and x67 and not x15 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x65 and not x62 and x63 and not x66 and not x64 and not x67 and x2 and x1 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( x65 and not x62 and x63 and not x66 and not x64 and not x67 and x2 and not x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x65 and not x62 and x63 and not x66 and not x64 and not x67 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and x66 and x67 and x1 ) = '1' then
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s40;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and x66 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and x66 and not x67 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s41;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and not x66 and x67 and x1 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s42;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and not x66 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and not x66 and not x67 and x1 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x65 and not x62 and not x63 and x2 and x64 and not x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and x66 and x67 and x1 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s44;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and x66 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and x66 and not x67 and x1 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s45;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and not x66 and x67 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s46;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and not x66 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and not x66 and not x67 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s47;

      elsif ( x65 and not x62 and not x63 and x2 and not x64 and not x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and not x2 and x1 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x65 and not x62 and not x63 and not x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and x66 and x64 and x67 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x65 and x62 and x66 and x64 and x67 and x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and x66 and x64 and x67 and not x2 and x32 and x33 and x1 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( not x65 and x62 and x66 and x64 and x67 and not x2 and x32 and x33 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and x66 and x64 and x67 and not x2 and x32 and not x33 and x1 ) = '1' then
         y3 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s49;

      elsif ( not x65 and x62 and x66 and x64 and x67 and not x2 and x32 and not x33 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and x66 and x64 and x67 and not x2 and not x32 and x1 ) = '1' then
         y3 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s49;

      elsif ( not x65 and x62 and x66 and x64 and x67 and not x2 and not x32 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and x11 and x13 and x1 and x3 and x6 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s50;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and x11 and x13 and x1 and x3 and not x6 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and x11 and x13 and x1 and not x3 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and x11 and x13 and not x1 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and x11 and not x13 and x5 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s52;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and x11 and not x13 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and not x11 and x8 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and not x11 and not x8 and x5 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and x12 and not x11 and not x8 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and x11 and x13 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and x11 and not x13 and x14 and x7 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and x11 and not x13 and x14 and not x7 and x1 and x5 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and x11 and not x13 and x14 and not x7 and x1 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and x11 and not x13 and x14 and not x7 and not x1 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and x11 and not x13 and not x14 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and x14 and x1 and x5 and x13 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and x14 and x1 and x5 and not x13 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and x14 and x1 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and x14 and not x1 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and not x14 and x13 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and not x14 and not x13 and x1 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and x10 and not x12 and not x11 and not x14 and not x13 and not x1 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( not x65 and x62 and x66 and x64 and not x67 and not x10 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( not x65 and x62 and x66 and not x64 and x67 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x65 and x62 and x66 and not x64 and not x67 and x6 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s60;

      elsif ( not x65 and x62 and x66 and not x64 and not x67 and not x6 and x7 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and x66 and not x64 and not x67 and not x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s61;

      elsif ( not x65 and x62 and not x66 and x64 and x67 and x2 and x1 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s62;

      elsif ( not x65 and x62 and not x66 and x64 and x67 and x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and x64 and x67 and not x2 and x1 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s63;

      elsif ( not x65 and x62 and not x66 and x64 and x67 and not x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and x10 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and x10 and not x1 and x2 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and x10 and not x1 and not x2 and x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and x10 and not x1 and not x2 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and x1 and x2 and x3 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and x1 and x2 and x3 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and x1 and x2 and not x3 and x4 and x5 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and x1 and x2 and not x3 and x4 and not x5 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and x1 and x2 and not x3 and not x4 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and x1 and not x2 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and x13 and not x10 and not x1 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and not x13 and not x12 and x10 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and not x13 and not x12 and x10 and not x1 and x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and not x13 and not x12 and x10 and not x1 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x65 and x62 and not x66 and x64 and not x67 and not x13 and not x12 and not x10 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( not x65 and x62 and not x66 and not x64 and x67 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( not x65 and x62 and not x66 and not x64 and x67 and x2 and not x1 ) = '1' then
         current_otherm <= s65;

      elsif ( not x65 and x62 and not x66 and not x64 and x67 and not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s66;

      elsif ( not x65 and x62 and not x66 and not x64 and x67 and not x2 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and x17 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and x17 and not x1 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and x17 and not x1 and not x2 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and x19 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and x19 and not x1 and x4 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and x19 and not x1 and not x4 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and x2 and x4 and x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and x2 and x4 and x5 and not x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and x2 and x4 and not x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and x2 and x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and x2 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and x2 and not x4 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and x1 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and x18 and not x17 and not x19 and not x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and x19 and x1 and x10 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and x19 and x1 and not x10 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and x19 and not x1 and x6 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and x19 and not x1 and not x6 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and x2 and x4 and x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and x2 and x4 and x5 and not x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and x2 and x4 and not x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and x2 and x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and x2 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and x2 and not x4 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and x1 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and x17 and not x19 and not x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x66 and not x64 and not x67 and not x18 and not x17 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and x2 and x67 and x1 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and x2 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and x2 and not x67 and x1 ) = '1' then
         y2 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s69;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and x2 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and not x2 and x67 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and not x2 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and not x2 and not x67 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( not x65 and not x62 and x63 and x66 and x64 and not x2 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and x1 and not x2 and x67 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and x1 and not x2 and not x67 and x5 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and x1 and not x2 and not x67 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and x1 and not x2 and not x67 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and not x1 and x67 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x66 and not x64 and not x1 and not x67 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and x11 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and x11 and not x14 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and x10 and x1 and x14 and x3 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and x10 and x1 and x14 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and x10 and x1 and x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and x10 and x1 and not x14 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and x10 and x1 and not x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and x10 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and not x10 and x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and not x10 and not x14 and x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and x67 and not x11 and not x10 and not x14 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and x10 and x1 and x14 and x3 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and x10 and x1 and x14 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and x10 and x1 and x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and x10 and x1 and not x14 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and x10 and x1 and not x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and x10 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and not x10 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and x15 and not x10 and not x14 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and x11 and x14 and x8 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and x11 and x14 and not x8 and x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and x11 and x14 and not x8 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and x11 and not x14 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s78;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and x11 and not x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and x14 and x10 and x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and x14 and x10 and not x7 and x1 and x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and x14 and x10 and not x7 and x1 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and x14 and x10 and not x7 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and x14 and not x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and not x14 and x1 and x10 and x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and not x14 and x1 and x10 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and not x14 and x1 and not x10 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and x13 and not x67 and not x15 and not x11 and not x14 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x65 and not x62 and x63 and not x66 and x64 and not x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and x67 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and x67 and x15 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and x67 and not x15 and x14 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and x67 and not x15 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and not x67 and x18 and x14 and x23 and x22 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and not x67 and x18 and x14 and x23 and not x22 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s81;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and not x67 and x18 and x14 and not x23 and x22 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s81;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and not x67 and x18 and x14 and not x23 and not x22 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and not x67 and x18 and not x14 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x65 and not x62 and x63 and not x66 and not x64 and not x67 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and x66 and x67 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and x66 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and x66 and not x67 and x1 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and not x66 and x67 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s83;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and not x66 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and not x66 and not x67 and x1 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s84;

      elsif ( not x65 and not x62 and not x63 and x2 and x64 and not x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and not x64 and x67 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      elsif ( not x65 and not x62 and not x63 and x2 and not x64 and x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and not x64 and not x67 and x66 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      elsif ( not x65 and not x62 and not x63 and x2 and not x64 and not x67 and x66 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x2 and not x64 and not x67 and not x66 and x1 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s45;

      elsif ( not x65 and not x62 and not x63 and x2 and not x64 and not x67 and not x66 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and not x2 and x66 and x67 and x64 and x1 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s85;

      elsif ( not x65 and not x62 and not x63 and not x2 and x66 and x67 and x64 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and not x2 and x66 and x67 and not x64 and x1 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x65 and not x62 and not x63 and not x2 and x66 and x67 and not x64 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and not x2 and x66 and not x67 and x1 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x65 and not x62 and not x63 and not x2 and x66 and not x67 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and not x2 and not x66 and x1 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      else
         current_otherm <= s1;

      end if;

   when s2 =>
      if ( x64 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s86;

      elsif ( not x64 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( not x64 and not x3 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( not x64 and not x3 and x1 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s66;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      end if;

   when s3 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s87;

      elsif ( not x62 and x64 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s88;

      elsif ( not x62 and not x64 and x65 and x66 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x62 and not x64 and x65 and not x66 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      else
         y3 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s91;

      end if;

   when s4 =>
         y12 <= '1' ;
         current_otherm <= s11;

   when s5 =>
      if ( x62 and x64 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( x62 and not x64 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x62 and not x64 and not x7 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( not x62 and x63 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s93;

      elsif ( not x62 and not x63 and x21 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      else
         y14 <= '1' ;
         current_otherm <= s95;

      end if;

   when s6 =>
      if ( x62 and x66 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x66 and x3 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( x62 and not x66 and x3 and not x2 ) = '1' then
         current_otherm <= s6;

      elsif ( x62 and not x66 and not x3 and x4 and x2 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( x62 and not x66 and not x3 and x4 and not x2 ) = '1' then
         current_otherm <= s6;

      elsif ( x62 and not x66 and not x3 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x66 and not x3 and not x4 and not x2 ) = '1' then
         current_otherm <= s6;

      elsif ( not x62 and x64 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s98;

      elsif ( not x62 and not x64 and x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and not x15 and x3 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and not x64 and not x15 and x3 and not x2 ) = '1' then
         current_otherm <= s6;

      elsif ( not x62 and not x64 and not x15 and not x3 and x4 and x2 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( not x62 and not x64 and not x15 and not x3 and x4 and not x2 ) = '1' then
         current_otherm <= s6;

      elsif ( not x62 and not x64 and not x15 and not x3 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      else
         current_otherm <= s6;

      end if;

   when s7 =>
      if ( x62 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s99;

      else
         y6 <= '1' ;
         current_otherm <= s100;

      end if;

   when s8 =>
      if ( x25 and x9 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x25 and not x9 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      end if;

   when s9 =>
      if ( x65 and x62 and x66 and x2 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x65 and x62 and x66 and x2 and not x4 and x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( x65 and x62 and x66 and x2 and not x4 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x65 and x62 and x66 and not x2 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x65 and x62 and x66 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x65 and x62 and not x66 and x5 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( x65 and x62 and not x66 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x65 and not x62 and x63 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x65 and not x62 and x63 and not x15 and x5 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( x65 and not x62 and x63 and not x15 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x65 and not x62 and not x63 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( not x65 and x62 and x18 and x17 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and x18 and x17 and not x1 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x62 and x18 and x17 and not x1 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and x18 and not x17 and x19 and x5 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x18 and not x17 and x19 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and x18 and not x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and not x18 and x17 and x7 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s104;

      elsif ( not x65 and x62 and not x18 and x17 and not x7 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s105;

      elsif ( not x65 and x62 and not x18 and not x17 and x19 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and not x18 and not x17 and not x19 and x5 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and not x18 and not x17 and not x19 and x5 and not x3 and x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x65 and x62 and not x18 and not x17 and not x19 and x5 and not x3 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and not x18 and not x17 and not x19 and not x5 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and not x62 and x63 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s99;

      elsif ( not x65 and not x62 and x63 and not x13 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s100;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and x5 and x12 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s108;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and x5 and not x12 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s109;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and x12 and x11 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and x12 and not x11 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and x12 and not x11 and x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and x12 and not x11 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and not x12 and x10 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and not x12 and not x10 and x9 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and not x12 and not x10 and x9 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and x6 and not x12 and not x10 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and not x6 and x12 ) = '1' then
         y58 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and x18 and x19 and not x3 and not x4 and not x5 and not x6 and not x12 ) = '1' then
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and x17 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s113;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and x12 and x5 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and x12 and not x5 and x14 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and x12 and not x5 and not x14 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and x12 and not x5 and not x14 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and x12 and not x5 and not x14 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and x12 and not x5 and not x14 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and not x12 and x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and not x12 and not x5 and x13 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and not x12 and not x5 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and not x12 and not x5 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and not x12 and not x5 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and x6 and not x12 and not x5 and not x13 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and x12 and x16 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and x12 and not x16 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and x12 and not x16 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and x12 and not x16 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and x12 and not x16 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and not x12 and x15 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and not x12 and not x15 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and not x12 and not x15 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and not x12 and not x15 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and x5 and not x12 and not x15 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x18 and not x19 and not x17 and not x3 and not x4 and not x6 and not x5 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and x19 and x12 and x6 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and x19 and x12 and not x6 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and x19 and not x12 and x6 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s99;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and x19 and not x12 and not x6 and x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and x19 and not x12 and not x6 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and x19 and not x12 and not x6 and not x3 and not x4 ) = '1' then
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and not x19 and x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and not x19 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and not x19 and not x3 and not x4 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x65 and not x62 and not x63 and not x18 and x5 and not x19 and not x3 and not x4 and not x6 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( not x65 and not x62 and not x63 and not x18 and not x5 and x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x65 and not x62 and not x63 and not x18 and not x5 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x62 and not x63 and not x18 and not x5 and not x3 and not x4 and x19 and x12 and x6 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x65 and not x62 and not x63 and not x18 and not x5 and not x3 and not x4 and x19 and x12 and not x6 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x65 and not x62 and not x63 and not x18 and not x5 and not x3 and not x4 and x19 and not x12 and x6 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x65 and not x62 and not x63 and not x18 and not x5 and not x3 and not x4 and x19 and not x12 and not x6 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      else
         y16 <= '1' ;
         current_otherm <= s123;

      end if;

   when s10 =>
      if ( x65 and x66 and x2 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x65 and x66 and x2 and not x4 and x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( x65 and x66 and x2 and not x4 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x65 and x66 and not x2 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x65 and x66 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x65 and not x66 and x6 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x65 and not x66 and x6 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x65 and not x66 and x6 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x65 and not x66 and x6 and not x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s125;

      elsif ( x65 and not x66 and not x6 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x66 and x4 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x65 and x66 and x4 and not x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x65 and x66 and not x4 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and not x66 and x18 and x17 and x4 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s126;

      elsif ( not x65 and not x66 and x18 and x17 and not x4 and x1 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x65 and not x66 and x18 and x17 and not x4 and x1 and not x3 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x65 and not x66 and x18 and x17 and not x4 and not x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and not x66 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and not x66 and not x18 and x17 and x11 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and not x66 and not x18 and x17 and not x11 and x16 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and not x66 and not x18 and x17 and not x11 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x66 and not x18 and not x17 and x19 and x1 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and not x66 and not x18 and not x17 and x19 and x1 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and not x66 and not x18 and not x17 and x19 and x1 and not x2 and not x3 ) = '1' then
         current_otherm <= s10;

      elsif ( not x65 and not x66 and not x18 and not x17 and x19 and not x1 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and not x66 and not x18 and not x17 and not x19 and x2 and x1 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and not x66 and not x18 and not x17 and not x19 and x2 and x1 and not x3 and x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x65 and not x66 and not x18 and not x17 and not x19 and x2 and x1 and not x3 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and not x66 and not x18 and not x17 and not x19 and x2 and not x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and not x66 and not x18 and not x17 and not x19 and not x2 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      else
         y4 <= '1' ;
         current_otherm <= s67;

      end if;

   when s11 =>
      if ( x62 and x25 and x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x62 and x25 and not x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x62 and not x25 and x26 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x62 and not x25 and x26 and not x7 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x62 and not x25 and not x26 and x12 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x62 and not x25 and not x26 and not x12 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( not x62 and x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 ) = '1' then
         y3 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s128;

      elsif ( not x62 and not x63 and not x64 and x65 and x66 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x65 and x66 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x65 and x66 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x66 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x66 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and not x64 and x65 and not x66 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and not x64 and x65 and not x66 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x66 and not x15 ) = '1' then
         current_otherm <= s1;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s12 =>
      if ( x64 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s130;

      elsif ( x64 and not x7 and x33 and x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s130;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and x13 and x5 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and x13 and not x5 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s132;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and not x13 and x8 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and not x13 and x8 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and not x13 and not x8 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and not x13 and not x8 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and not x13 and not x8 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and x14 and not x13 and not x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and x13 and x31 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and x13 and x31 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and x13 and not x31 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and x13 and not x31 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and x13 and not x31 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and x13 and not x31 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and not x13 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and x15 and not x14 and not x13 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and x14 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s136;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and x14 and not x5 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and not x14 and x16 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and not x14 and x16 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and not x14 and not x16 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and not x14 and not x16 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and not x14 and not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and x13 and not x14 and not x16 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and x14 and x30 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and x14 and x30 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and x14 and not x30 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and x14 and not x30 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and x14 and not x30 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and x14 and not x30 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and x33 and not x32 and x9 and not x15 and not x13 and not x14 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s138;

      elsif ( x64 and not x7 and x33 and not x32 and not x9 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s139;

      elsif ( x64 and not x7 and not x33 and x9 and x13 and x32 and x15 and x14 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( x64 and not x7 and not x33 and x9 and x13 and x32 and x15 and not x14 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s140;

      elsif ( x64 and not x7 and not x33 and x9 and x13 and x32 and x15 and not x14 and not x16 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s141;

      elsif ( x64 and not x7 and not x33 and x9 and x13 and x32 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s142;

      elsif ( x64 and not x7 and not x33 and x9 and x13 and x32 and not x15 and not x14 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s143;

      elsif ( x64 and not x7 and not x33 and x9 and x13 and not x32 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s144;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and x32 and x15 and x14 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s145;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and x32 and x15 and not x14 and x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and x32 and x15 and not x14 and not x17 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s146;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and x32 and not x15 and x14 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s147;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and x32 and not x15 and not x14 and x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and x32 and not x15 and not x14 and not x18 ) = '1' then
         current_otherm <= s12;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and not x32 and x4 and x6 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s148;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and not x32 and x4 and not x6 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( x64 and not x7 and not x33 and x9 and not x13 and not x32 and not x4 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s149;

      elsif ( x64 and not x7 and not x33 and not x9 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s139;

      else
         current_otherm <= s1;

      end if;

   when s13 =>
      if ( x62 and x64 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x64 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x64 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x18 and x17 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( x62 and not x64 and x18 and x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x64 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x64 and not x18 and x17 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x64 and not x18 and not x17 and x19 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x64 and not x18 and not x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x63 and x65 and x66 and x31 and x5 ) = '1' then
         y23 <= '1' ;
         y51 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s152;

      elsif ( not x62 and x63 and x65 and x66 and x31 and not x5 and x22 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s153;

      elsif ( not x62 and x63 and x65 and x66 and x31 and not x5 and not x22 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      elsif ( not x62 and x63 and x65 and x66 and not x31 and x5 ) = '1' then
         y65 <= '1' ;
         current_otherm <= s155;

      elsif ( not x62 and x63 and x65 and x66 and not x31 and not x5 ) = '1' then
         y71 <= '1' ;
         current_otherm <= s156;

      elsif ( not x62 and x63 and x65 and not x66 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y55 <= '1' ;
         y58 <= '1' ;
         y69 <= '1' ;
         current_otherm <= s157;

      elsif ( not x62 and x63 and not x65 ) = '1' then
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s158;

      else
         y2 <= '1' ;
         y15 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s159;

      end if;

   when s14 =>
      if ( x62 and x66 and x25 and x8 ) = '1' then
         y2 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s160;

      elsif ( x62 and x66 and x25 and not x8 ) = '1' then
         y1 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s160;

      elsif ( x62 and x66 and not x25 and x13 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( x62 and x66 and not x25 and not x13 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x62 and not x66 and x13 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x66 and x13 and not x11 and x6 and x4 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( x62 and not x66 and x13 and not x11 and x6 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x66 and x13 and not x11 and not x6 and x5 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( x62 and not x66 and x13 and not x11 and not x6 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( x62 and not x66 and not x13 and x14 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( x62 and not x66 and not x13 and not x14 and x9 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( x62 and not x66 and not x13 and not x14 and not x9 and x6 and x2 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( x62 and not x66 and not x13 and not x14 and not x9 and x6 and not x2 ) = '1' then
         current_otherm <= s14;

      elsif ( x62 and not x66 and not x13 and not x14 and not x9 and not x6 and x8 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( x62 and not x66 and not x13 and not x14 and not x9 and not x6 and not x8 ) = '1' then
         current_otherm <= s14;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and x67 and x11 and not x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and x64 and x67 and not x11 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and x64 and not x67 and x10 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and x64 and not x67 and not x10 and x15 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and not x10 and x15 and not x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and x64 and not x67 and not x10 and not x15 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and not x64 and x65 and x66 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and not x64 and x65 and x66 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and x13 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and x13 and not x11 and x6 and x4 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and x13 and not x11 and x6 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and x13 and not x11 and not x6 and x5 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and x13 and not x11 and not x6 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and not x13 and x14 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and not x13 and not x14 and x9 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and not x13 and not x14 and not x9 and x6 and x2 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and not x13 and not x14 and not x9 and x6 and not x2 ) = '1' then
         current_otherm <= s14;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and not x13 and not x14 and not x9 and not x6 and x8 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and x63 and not x64 and x65 and not x66 and not x15 and not x13 and not x14 and not x9 and not x6 and not x8 ) = '1' then
         current_otherm <= s14;

      elsif ( not x62 and x63 and not x64 and not x65 and x66 and x11 ) = '1' then
         y14 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s163;

      elsif ( not x62 and x63 and not x64 and not x65 and x66 and not x11 ) = '1' then
         y10 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s164;

      elsif ( not x62 and x63 and not x64 and not x65 and not x66 and x12 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( not x62 and x63 and not x64 and not x65 and not x66 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x62 and x63 and not x64 and not x65 and not x66 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x62 and x63 and not x64 and not x65 and not x66 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x64 and not x65 and not x66 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x63 and x64 and x6 and not x7 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x63 and x64 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and x23 and x24 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and x23 and x24 and x10 and not x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and x23 and x24 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and x23 and x24 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and x23 and not x24 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s167;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and x10 and x24 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and x10 and x24 and not x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and x10 and not x24 and x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and x10 and not x24 and not x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and x13 and x14 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and x13 and not x14 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and x13 and not x14 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and x13 and not x14 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and x13 and not x14 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and not x13 and x15 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and not x13 and not x15 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and not x13 and not x15 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and not x13 and not x15 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and x24 and not x13 and not x15 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and not x24 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and x9 and not x10 and not x24 and not x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and x17 and x18 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and x17 and not x18 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and x17 and not x18 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and x17 and not x18 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and x17 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and not x17 and x19 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and not x17 and not x19 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and not x17 and not x19 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and not x17 and not x19 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and x16 and not x17 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and x24 and not x16 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and not x24 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and not x24 and x8 and not x10 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 and not x23 and not x9 and not x24 and not x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( not x62 and not x63 and not x64 and x66 and not x67 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x66 and not x67 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x66 and not x67 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and not x67 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s15 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s174;

   when s16 =>
      if ( x62 and x64 and x65 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x64 and x65 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x64 and x65 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x65 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and not x65 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x64 and not x65 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x64 and not x65 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and not x65 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x66 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( x62 and not x64 and not x66 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( x62 and not x64 and not x66 and not x8 and x9 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( x62 and not x64 and not x66 and not x8 and not x9 and x10 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x62 and not x64 and not x66 and not x8 and not x9 and x10 and not x6 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x62 and not x64 and not x66 and not x8 and not x9 and not x10 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x64 and not x66 and not x8 and not x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s16;

      elsif ( not x62 and x64 and x63 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s177;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and x9 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and x3 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and x3 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and x3 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and x3 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and x6 and not x7 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and x6 and not x7 and x12 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and x6 and not x7 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and not x6 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and not x6 and not x8 and x12 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and not x6 and not x8 and x12 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and x5 and not x3 and not x6 and not x8 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and not x5 and x6 and x3 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and not x5 and x6 and not x3 ) = '1' then
         y21 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s180;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and not x5 and not x6 and x3 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and x20 and not x9 and not x5 and not x6 and not x3 ) = '1' then
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s180;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and not x20 and x4 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and not x20 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and not x20 and not x4 and not x5 and x15 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x21 and not x20 and not x4 and not x5 and not x15 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s183;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and x4 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and x9 and x8 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and x9 and x8 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and x9 and x8 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and x9 and x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and x9 and not x8 and x10 ) = '1' then
         y21 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s180;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and x9 and not x8 and not x10 ) = '1' then
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s180;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and x8 and x10 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s184;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and x8 and not x10 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s184;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and x10 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and x10 and not x11 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and x10 and not x11 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and x10 and not x11 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and x10 and not x11 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and not x10 and x12 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and not x10 and not x12 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and not x10 and not x12 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and not x10 and not x12 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and x20 and not x9 and not x8 and not x10 and not x12 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and not x20 and x6 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x21 and not x4 and not x20 and not x6 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s185;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x66 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and not x15 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and not x15 and not x8 and x9 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and not x15 and not x8 and not x9 and x10 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and not x15 and not x8 and not x9 and x10 and not x6 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and not x15 and not x8 and not x9 and not x10 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x63 and not x66 and x65 and not x15 and not x8 and not x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s16;

      elsif ( not x62 and not x64 and x63 and not x66 and not x65 and x23 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s187;

      elsif ( not x62 and not x64 and x63 and not x66 and not x65 and x23 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s188;

      elsif ( not x62 and not x64 and x63 and not x66 and not x65 and not x23 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s188;

      elsif ( not x62 and not x64 and x63 and not x66 and not x65 and not x23 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s187;

      elsif ( not x62 and not x64 and not x63 and x67 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s189;

      else
         current_otherm <= s1;

      end if;

   when s17 =>
      if ( x62 and x66 and x18 and x17 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( x62 and x66 and x18 and x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and x66 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and x66 and not x18 and x17 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and x66 and not x18 and not x17 and x19 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and x66 and not x18 and not x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x66 and x3 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( x62 and not x66 and x3 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( x62 and not x66 and not x3 and x4 and x2 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( x62 and not x66 and not x3 and x4 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( x62 and not x66 and not x3 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x66 and not x3 and not x4 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( not x62 and x65 and x63 and x66 and x67 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x62 and x65 and x63 and x66 and not x67 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x65 and x63 and not x66 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s6;

      elsif ( not x62 and x65 and x63 and not x66 and not x15 and x3 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x65 and x63 and not x66 and not x15 and x3 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( not x62 and x65 and x63 and not x66 and not x15 and not x3 and x4 and x2 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( not x62 and x65 and x63 and not x66 and not x15 and not x3 and x4 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( not x62 and x65 and x63 and not x66 and not x15 and not x3 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and x65 and x63 and not x66 and not x15 and not x3 and not x4 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( not x62 and x65 and not x63 and x66 and x64 and x67 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and x65 and not x63 and x66 and x64 and not x67 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x65 and not x63 and x66 and not x64 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x65 and not x63 and not x66 and x64 and x67 and x21 and x20 ) = '1' then
         y60 <= '1' ;
         current_otherm <= s190;

      elsif ( not x62 and x65 and not x63 and not x66 and x64 and x67 and x21 and not x20 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x65 and not x63 and not x66 and x64 and x67 and not x21 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x65 and not x63 and not x66 and x64 and not x67 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s191;

      elsif ( not x62 and x65 and not x63 and not x66 and not x64 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      elsif ( not x62 and not x65 and x63 and x66 and x67 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and x3 and x5 and x7 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s192;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and x3 and x5 and not x7 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and x3 and x5 and not x7 and x1 and not x2 ) = '1' then
         current_otherm <= s17;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and x3 and x5 and not x7 and not x1 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and x3 and not x5 and x6 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s193;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and x3 and not x5 and not x6 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s192;

      elsif ( not x62 and not x65 and x63 and x66 and not x67 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and not x65 and x63 and not x66 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      elsif ( not x62 and not x65 and not x63 and x64 and x66 and x67 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      elsif ( not x62 and not x65 and not x63 and x64 and x66 and not x67 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and not x65 and not x63 and x64 and not x66 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s18 =>
      if ( x62 and x65 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and x65 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x62 and x65 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and x65 and not x4 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s194;

      elsif ( x62 and not x65 and x3 and x1 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s195;

      elsif ( x62 and not x65 and x3 and not x1 and x4 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s195;

      elsif ( x62 and not x65 and x3 and not x1 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and not x65 and not x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      else
         y8 <= '1' ;
         current_otherm <= s127;

      end if;

   when s19 =>
      if ( x65 and x6 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x65 and x6 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x65 and x6 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x65 and x6 and not x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s125;

      elsif ( x65 and not x6 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s2;

      elsif ( not x65 and not x5 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s196;

      elsif ( not x65 and not x5 and x2 and not x1 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s197;

      elsif ( not x65 and not x5 and not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s198;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s2;

      end if;

   when s20 =>
      if ( x65 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x65 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x65 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x65 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x17 and x18 and not x1 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x17 and x18 and not x1 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x17 and not x18 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and not x17 and x18 and x2 and x19 and x4 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x65 and not x17 and x18 and x2 and x19 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and not x17 and x18 and x2 and not x19 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x17 and x18 and not x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x17 and not x18 and x19 and x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and not x17 and not x18 and x19 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x17 and not x18 and not x19 and x1 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and not x17 and not x18 and not x19 and x1 and not x3 and x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x65 and not x17 and not x18 and not x19 and x1 and not x3 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      else
         y5 <= '1' ;
         current_otherm <= s68;

      end if;

   when s21 =>
      if ( x62 and x64 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s199;

      elsif ( x62 and not x64 and x65 and x3 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and not x64 and x65 and not x3 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and not x64 and x65 and not x3 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x62 and not x64 and x65 and not x3 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x64 and x65 and not x3 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x64 and not x65 and x66 and x4 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( x62 and not x64 and not x65 and x66 and x4 and not x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x64 and not x65 and x66 and not x4 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and not x64 and not x65 and not x66 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and not x64 and not x65 and not x66 and not x3 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( x62 and not x64 and not x65 and not x66 and not x3 and x1 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s66;

      elsif ( x62 and not x64 and not x65 and not x66 and not x3 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x62 and x65 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s200;

      else
         y14 <= '1' ;
         current_otherm <= s201;

      end if;

   when s22 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s202;

   when s23 =>
      if ( x63 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      elsif ( not x63 and x64 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      elsif ( not x63 and not x64 and x67 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      else
         y24 <= '1' ;
         current_otherm <= s203;

      end if;

   when s24 =>
      if ( x62 and x17 and x18 and x65 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( x62 and x17 and x18 and x65 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and x17 and x18 and not x65 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x62 and x17 and not x18 and x65 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and x17 and not x18 and not x65 and x14 and x5 ) = '1' then
         current_otherm <= s24;

      elsif ( x62 and x17 and not x18 and not x65 and x14 and not x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and x17 and not x18 and not x65 and not x14 and x5 ) = '1' then
         current_otherm <= s24;

      elsif ( x62 and x17 and not x18 and not x65 and not x14 and not x5 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( x62 and not x17 and x18 and x65 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x17 and x18 and not x65 and x19 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x62 and not x17 and x18 and not x65 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x17 and not x18 and x19 and x65 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x17 and not x18 and x19 and not x65 and x4 and x1 ) = '1' then
         current_otherm <= s24;

      elsif ( x62 and not x17 and not x18 and x19 and not x65 and x4 and not x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x17 and not x18 and x19 and not x65 and not x4 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x62 and not x17 and not x18 and not x19 and x65 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x17 and not x18 and not x19 and not x65 ) = '1' then
         current_otherm <= s24;

      elsif ( not x62 and x64 and x63 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s205;

      elsif ( not x62 and x64 and not x63 and x66 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s206;

      elsif ( not x62 and x64 and not x63 and not x66 and x21 and x20 ) = '1' then
         y4 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s207;

      elsif ( not x62 and x64 and not x63 and not x66 and x21 and not x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x62 and x64 and not x63 and not x66 and not x21 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x62 and not x64 and x63 and x65 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x62 and not x64 and x63 and not x65 and x4 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s208;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and x5 and x7 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s192;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and x5 and not x7 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and x5 and not x7 and x1 and not x2 and x3 ) = '1' then
         current_otherm <= s24;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and x5 and not x7 and x1 and not x2 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and x5 and not x7 and not x1 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and not x5 and x6 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s193;

      elsif ( not x62 and not x64 and x63 and not x65 and not x4 and not x5 and not x6 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s192;

      elsif ( not x62 and not x64 and not x63 and x67 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      else
         y3 <= '1' ;
         current_otherm <= s208;

      end if;

   when s25 =>
         y36 <= '1' ;
         current_otherm <= s209;

   when s26 =>
         y1 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s210;

   when s27 =>
      if ( x62 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( x62 and x4 and not x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      elsif ( x62 and not x4 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and x16 and x15 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and x16 and not x15 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and x16 and not x15 and x4 and not x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      elsif ( not x62 and x16 and not x15 and not x4 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and not x16 and x15 and x6 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and not x16 and x15 and not x6 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      else
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      end if;

   when s28 =>
      if ( x62 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( x62 and x4 and not x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s214;

      elsif ( x62 and not x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      elsif ( not x62 and x15 and x6 and x16 and x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x15 and x6 and x16 and not x5 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x15 and x6 and not x16 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and x15 and not x6 and x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x15 and not x6 and not x16 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and not x15 and x16 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and not x15 and x16 and x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and not x15 and x16 and not x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      end if;

   when s29 =>
      if ( x62 and x4 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      elsif ( x62 and not x4 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and x16 and x15 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and x16 and not x15 and x4 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      elsif ( not x62 and x16 and not x15 and not x4 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and not x16 and x15 and x12 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and not x16 and x15 and not x12 ) = '1' then
         current_otherm <= s29;

      elsif ( not x62 and not x16 and not x15 and x14 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      else
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      end if;

   when s30 =>
      if ( x62 and x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( x62 and x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( x62 and x4 and not x5 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( x62 and x4 and not x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( x62 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s221;

      elsif ( not x62 and x64 and x63 and x16 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and x64 and x63 and x16 and not x15 and x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x62 and x64 and x63 and x16 and not x15 and x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and x64 and x63 and x16 and not x15 and x4 and not x5 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and x64 and x63 and x16 and not x15 and x4 and not x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and x64 and x63 and x16 and not x15 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and x64 and x63 and not x16 and x15 and x3 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x64 and x63 and not x16 and x15 and x3 and not x2 ) = '1' then
         current_otherm <= s30;

      elsif ( not x62 and x64 and x63 and not x16 and x15 and not x3 and x4 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and x64 and x63 and not x16 and x15 and not x3 and x4 and not x2 ) = '1' then
         current_otherm <= s30;

      elsif ( not x62 and x64 and x63 and not x16 and x15 and not x3 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and x64 and x63 and not x16 and x15 and not x3 and not x4 and not x2 ) = '1' then
         current_otherm <= s30;

      elsif ( not x62 and x64 and x63 and not x16 and not x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x67 and x21 and x20 ) = '1' then
         y60 <= '1' ;
         current_otherm <= s190;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x67 and x21 and not x20 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and x67 and not x21 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x62 and x64 and not x63 and x65 and not x66 and not x67 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s222;

      elsif ( not x62 and x64 and not x63 and not x65 and x67 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s223;

      elsif ( not x62 and x64 and not x63 and not x65 and not x67 and x18 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( not x62 and x64 and not x63 and not x65 and not x67 and not x18 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x65 and not x67 and not x18 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x65 and not x67 and not x18 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and not x67 and not x18 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x65 ) = '1' then
         y63 <= '1' ;
         current_otherm <= s224;

      elsif ( not x62 and not x64 and x63 and not x65 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( not x62 and not x64 and x63 and not x65 and not x7 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x62 and not x64 and not x63 and x65 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and not x63 and x65 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and not x63 and x65 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x65 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s31 =>
      if ( x15 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( x15 and not x16 and x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( x15 and not x16 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x15 and x16 and x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x15 and x16 and x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x15 and x16 and x4 and not x5 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x15 and x16 and x4 and not x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x15 and x16 and not x4 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x15 and x16 and not x4 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      else
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      end if;

   when s32 =>
      if ( x62 and x13 and x10 and x9 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x62 and x13 and x10 and not x9 and x17 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and x13 and x10 and not x9 and not x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and x13 and not x10 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and not x13 and x12 and x1 and x2 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and not x13 and x12 and x1 and not x2 and x3 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and not x13 and x12 and x1 and not x2 and not x3 ) = '1' then
         current_otherm <= s32;

      elsif ( x62 and not x13 and x12 and not x1 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x62 and not x13 and not x12 and x1 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( x62 and not x13 and not x12 and x1 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and not x13 and not x12 and x1 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x12 and x1 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and not x13 and not x12 and not x1 and x2 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and not x13 and not x12 and not x1 and not x2 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and x18 and x4 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      elsif ( not x62 and x17 and x18 and not x4 and x1 and x3 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and x17 and x18 and not x4 and x1 and not x3 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( not x62 and x17 and x18 and not x4 and not x1 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and x17 and not x18 and x11 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( not x62 and x17 and not x18 and not x11 and x16 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and x17 and not x18 and not x11 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and x18 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and not x17 and not x18 and x15 and x1 and x2 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and not x17 and not x18 and x15 and x1 and not x2 and x3 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and not x17 and not x18 and x15 and x1 and not x2 and not x3 ) = '1' then
         current_otherm <= s32;

      elsif ( not x62 and not x17 and not x18 and x15 and not x1 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x18 and not x15 and x2 and x1 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x18 and not x15 and x2 and x1 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and not x17 and not x18 and not x15 and x2 and x1 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and not x17 and not x18 and not x15 and x2 and not x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and not x17 and not x18 and not x15 and not x2 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      else
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      end if;

   when s33 =>
      if ( x62 and x13 and x10 and x17 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and x13 and x10 and not x17 and x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and x13 and x10 and not x17 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and x13 and not x10 and x3 and x15 ) = '1' then
         current_otherm <= s33;

      elsif ( x62 and x13 and not x10 and x3 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and x13 and not x10 and not x3 and x4 and x5 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and x13 and not x10 and not x3 and x4 and not x5 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x62 and x13 and not x10 and not x3 and not x4 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and not x13 and x12 and x4 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and not x13 and x12 and not x4 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and not x12 and x10 and x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and not x12 and x10 and not x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s232;

      elsif ( x62 and not x13 and not x12 and not x10 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 and x6 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( not x62 and x17 and x18 and not x6 and x8 and x4 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      elsif ( not x62 and x17 and x18 and not x6 and x8 and not x4 and x1 and x3 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and x17 and x18 and not x6 and x8 and not x4 and x1 and not x3 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( not x62 and x17 and x18 and not x6 and x8 and not x4 and not x1 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and x17 and x18 and not x6 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x17 and not x18 and x12 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( not x62 and x17 and not x18 and not x12 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and not x17 and x15 and x18 and x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and x15 and x18 and not x9 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s232;

      elsif ( not x62 and not x17 and x15 and not x18 and x2 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and x15 and not x18 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and not x15 and x18 and x4 and x5 and x3 ) = '1' then
         current_otherm <= s33;

      elsif ( not x62 and not x17 and not x15 and x18 and x4 and x5 and not x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and not x15 and x18 and x4 and not x5 and x3 ) = '1' then
         current_otherm <= s33;

      elsif ( not x62 and not x17 and not x15 and x18 and x4 and not x5 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x15 and x18 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and not x17 and not x15 and x18 and not x4 and not x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      end if;

   when s34 =>
      if ( x62 and x13 and x10 and x9 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x62 and x13 and x10 and not x9 and x17 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and x13 and x10 and not x9 and not x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and x13 and not x10 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and not x13 and x12 and x4 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and not x13 and x12 and not x4 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and not x12 and x10 and x2 and x16 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( x62 and not x13 and not x12 and x10 and x2 and not x16 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x12 and x10 and not x2 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and not x13 and not x12 and not x10 and x18 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( x62 and not x13 and not x12 and not x10 and x18 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and not x13 and not x12 and not x10 and x18 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x12 and not x10 and not x18 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x18 and not x1 and x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 and not x1 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x17 and not x18 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and not x17 and x15 and x18 and x2 and x4 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( not x62 and not x17 and x15 and x18 and x2 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and not x17 and x15 and x18 and not x2 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and x15 and not x18 and x2 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and x15 and not x18 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and not x15 and x1 and x18 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and not x15 and x1 and not x18 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x15 and x1 and not x18 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and not x17 and not x15 and x1 and not x18 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      end if;

   when s35 =>
      if ( x62 and x13 and x10 and x6 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and x13 and x10 and not x6 and x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and x13 and x10 and not x6 and not x4 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x13 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x12 and x10 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s233;

      elsif ( x62 and not x13 and not x12 and not x10 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and x17 and x18 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s234;

      elsif ( not x62 and x17 and x18 and not x7 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      elsif ( not x62 and x17 and not x18 ) = '1' then
         current_otherm <= s35;

      elsif ( not x62 and not x17 and x18 and x15 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s233;

      elsif ( not x62 and not x17 and x18 and not x15 ) = '1' then
         current_otherm <= s1;

      else
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      end if;

   when s36 =>
      if ( x62 and x13 and x10 and x7 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and x13 and x10 and not x7 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and x13 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and x12 and x15 and x9 ) = '1' then
         current_otherm <= s36;

      elsif ( x62 and not x13 and x12 and x15 and not x9 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and x12 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and not x13 and not x12 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s232;

      elsif ( not x62 and x17 and not x18 and x14 and x5 ) = '1' then
         current_otherm <= s36;

      elsif ( not x62 and x17 and not x18 and x14 and not x5 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and x17 and not x18 and not x14 and x5 ) = '1' then
         current_otherm <= s36;

      elsif ( not x62 and x17 and not x18 and not x14 and not x5 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( not x62 and not x17 and x15 and x18 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and x15 and not x18 and x4 and x1 ) = '1' then
         current_otherm <= s36;

      elsif ( not x62 and not x17 and x15 and not x18 and x4 and not x1 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and not x17 and x15 and not x18 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and not x17 and not x15 and x18 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s36;

      end if;

   when s37 =>
      if ( x62 and x13 and x10 and x3 and x5 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( x62 and x13 and x10 and x3 and not x5 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and x13 and x10 and not x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and x13 and not x10 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x62 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and not x13 and not x12 and x10 and x5 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and not x13 and not x12 and x10 and not x5 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x12 and not x10 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( x62 and not x13 and not x12 and not x10 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and not x13 and not x12 and not x10 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x12 and not x10 and not x5 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x18 and not x1 and x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 and not x1 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x17 and not x18 and x7 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s233;

      elsif ( not x62 and x17 and not x18 and not x7 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      elsif ( not x62 and not x17 and x15 and x18 and x5 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and not x17 and x15 and x18 and not x5 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and not x17 and x15 and not x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and not x17 and not x15 and x5 and x18 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x15 and x5 and not x18 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x15 and x5 and not x18 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and not x17 and not x15 and x5 and not x18 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      else
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      end if;

   when s38 =>
      if ( x63 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s236;

      elsif ( not x63 and x64 and x65 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x64 and x65 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x64 and x65 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x67 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x67 and x28 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and not x67 and x28 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and not x67 and x28 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x67 and x28 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y8 <= '1' ;
         current_otherm <= s237;

      end if;

   when s39 =>
      if ( x65 and x62 and x64 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x65 and x62 and not x64 and x66 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x65 and x62 and not x64 and x66 and not x6 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x65 and x62 and not x64 and not x66 and x67 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and x62 and not x64 and not x66 and not x67 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x65 and x62 and not x64 and not x66 and not x67 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x65 and x62 and not x64 and not x66 and not x67 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x65 and x62 and not x64 and not x66 and not x67 and not x4 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s194;

      elsif ( x65 and not x62 and x63 and x66 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x65 and not x62 and x63 and x66 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x65 and not x62 and x63 and not x66 and x67 and x15 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( x65 and not x62 and x63 and not x66 and x67 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and not x66 and not x67 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x65 and not x62 and not x63 and x64 and x67 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and x10 and x14 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and x10 and not x14 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and x14 and x8 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and x14 and not x8 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and x14 and not x8 and x6 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and x14 and not x8 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and not x14 and x7 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and not x14 and not x7 and x6 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and not x14 and not x7 and x6 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and x11 and not x14 and not x7 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and not x11 and x14 ) = '1' then
         y60 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y67 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s240;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and x21 and not x10 and not x11 and not x14 ) = '1' then
         y58 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s240;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and not x21 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and not x21 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and not x21 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and x22 and not x21 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and not x22 and x12 and x21 and x11 ) = '1' then
         y7 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s240;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and not x22 and x12 and x21 and not x11 ) = '1' then
         y7 <= '1' ;
         y62 <= '1' ;
         y74 <= '1' ;
         y110 <= '1' ;
         current_otherm <= s241;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and not x22 and x12 and not x21 and x10 ) = '1' then
         y7 <= '1' ;
         y62 <= '1' ;
         y90 <= '1' ;
         y92 <= '1' ;
         current_otherm <= s240;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and not x22 and x12 and not x21 and not x10 ) = '1' then
         y7 <= '1' ;
         y62 <= '1' ;
         y92 <= '1' ;
         y93 <= '1' ;
         y97 <= '1' ;
         current_otherm <= s240;

      elsif ( x65 and not x62 and not x63 and x64 and not x67 and not x22 and not x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s242;

      elsif ( x65 and not x62 and not x63 and not x64 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and x64 and x12 and x9 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x64 and x12 and not x9 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x65 and x62 and x64 and x12 and not x9 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and x12 and not x9 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( not x65 and x62 and x64 and x12 and not x9 and not x3 and not x1 and not x7 ) = '1' then
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and x11 and x4 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and x11 and not x4 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and not x11 and x14 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and not x11 and not x14 and x9 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and not x11 and not x14 and not x9 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and not x11 and not x14 and not x9 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and not x11 and not x14 and not x9 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and x13 and not x11 and not x14 and not x9 and not x3 and not x1 and not x7 ) = '1' then
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and not x13 and x9 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and not x13 and not x9 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and not x13 and not x9 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and not x13 and not x9 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( not x65 and x62 and x64 and not x12 and x10 and not x13 and not x9 and not x3 and not x1 and not x7 ) = '1' then
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and not x12 and not x10 and x9 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x64 and not x12 and not x10 and not x9 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x65 and x62 and x64 and not x12 and not x10 and not x9 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x65 and x62 and x64 and not x12 and not x10 and not x9 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( not x65 and x62 and x64 and not x12 and not x10 and not x9 and not x3 and not x1 and not x7 ) = '1' then
         current_otherm <= s39;

      elsif ( not x65 and x62 and not x64 and x66 and x1 and x2 and x3 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and x62 and not x64 and x66 and x1 and x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s245;

      elsif ( not x65 and x62 and not x64 and x66 and x1 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x65 and x62 and not x64 and x66 and not x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x64 and not x66 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x62 and not x64 and not x66 and x17 and x18 and not x1 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x62 and not x64 and not x66 and x17 and x18 and not x1 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and not x64 and not x66 and x17 and not x18 and x7 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x65 and x62 and not x64 and not x66 and x17 and not x18 and not x7 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x62 and not x64 and not x66 and not x17 and x18 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and not x64 and not x66 and not x17 and x18 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s246;

      elsif ( not x65 and x62 and not x64 and not x66 and not x17 and not x18 and x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x64 and not x66 and not x17 and not x18 and not x19 and x1 and x2 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x65 and x62 and not x64 and not x66 and not x17 and not x18 and not x19 and x1 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x64 and not x66 and not x17 and not x18 and not x19 and not x1 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x65 and not x62 and x63 and x66 and x8 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x65 and not x62 and x63 and x66 and not x8 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s60;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and x16 and x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s247;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and x16 and not x23 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and x16 and not x23 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and x16 and not x23 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and x16 and not x23 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and x16 and not x23 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and not x16 and x23 ) = '1' then
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s248;

      elsif ( not x65 and not x62 and x63 and not x66 and x22 and not x16 and not x23 ) = '1' then
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s249;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and x9 and x8 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and x9 and x8 and not x10 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and x9 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and x8 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and x8 and not x13 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and x8 and not x13 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and x8 and not x13 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and x8 and not x13 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and x8 and not x13 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and not x8 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and not x8 and not x3 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and not x8 and not x3 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and not x8 and not x3 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and not x8 and not x3 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and x10 and not x8 and not x3 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and x8 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and x8 and not x1 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and x8 and not x1 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and x8 and not x1 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and x8 and not x1 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and x8 and not x1 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and not x8 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and not x8 and not x15 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and not x8 and not x15 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and not x8 and not x15 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and not x8 and not x15 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and x7 and not x9 and not x10 and not x8 and not x15 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and x23 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s251;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and x16 and not x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s247;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and not x16 and x23 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s252;

      elsif ( not x65 and not x62 and x63 and not x66 and not x22 and not x16 and not x23 ) = '1' then
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s248;

      elsif ( not x65 and not x62 and not x63 and x64 and x4 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and x19 and x12 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and x19 and not x12 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s254;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and x12 and x6 ) = '1' then
         y16 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s255;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and x12 and not x6 and x16 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and not x12 and x6 ) = '1' then
         y12 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s257;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and not x12 and not x6 and x15 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and not x18 and x19 ) = '1' then
         y27 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and not x18 and not x19 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and x5 and not x18 and not x19 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and x12 and x11 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and x12 and not x11 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and not x12 and x10 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and x6 and not x12 and not x10 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and not x6 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and x19 and not x6 and not x12 ) = '1' then
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and x12 and x14 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and not x12 and x13 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and x18 and not x19 and not x6 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and not x18 and x19 and x12 and x6 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s260;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and not x18 and x19 and x12 and not x6 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s261;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and not x18 and x19 and not x12 and x6 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and not x18 and x19 and not x12 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and x8 and not x5 and not x18 and not x19 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x65 and not x62 and not x63 and x64 and not x4 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x65 and not x62 and not x63 and not x64 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x65 and not x62 and not x63 and not x64 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x65 and not x62 and not x63 and not x64 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and not x64 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s40 =>
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s264;

   when s41 =>
      if ( x62 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s265;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s266;

      end if;

   when s42 =>
      if ( x21 and x20 ) = '1' then
         y15 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s267;

      elsif ( x21 and not x20 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( not x21 and x20 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      else
         y5 <= '1' ;
         current_otherm <= s74;

      end if;

   when s43 =>
      if ( x62 and x64 and x9 and x32 and x33 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s139;

      elsif ( x62 and x64 and x9 and x32 and not x33 and x14 and x15 and x13 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( x62 and x64 and x9 and x32 and not x33 and x14 and x15 and not x13 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s145;

      elsif ( x62 and x64 and x9 and x32 and not x33 and x14 and not x15 and x13 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s142;

      elsif ( x62 and x64 and x9 and x32 and not x33 and x14 and not x15 and not x13 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s147;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and x15 and x13 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s140;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and x15 and x13 and not x16 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s141;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and x15 and not x13 and x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and x15 and not x13 and not x17 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s146;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and not x15 and x13 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s143;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and not x15 and not x13 and x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and x32 and not x33 and not x14 and not x15 and not x13 and not x18 ) = '1' then
         current_otherm <= s43;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and x14 and x5 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and x14 and not x5 and x7 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and x14 and not x5 and not x7 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s132;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and not x14 and x31 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and not x14 and x31 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and not x14 and not x31 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and not x14 and not x31 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and not x14 and not x31 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and x15 and not x14 and not x31 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and x14 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s136;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and x14 and not x5 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and not x14 and x16 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and not x14 and x16 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and not x14 and not x16 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and not x14 and not x16 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and not x14 and not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and x13 and x33 and not x15 and not x14 and not x16 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and x13 and not x33 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s144;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and x15 and x8 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and x15 and x8 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and x15 and not x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and not x15 and x30 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and not x15 and x30 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and not x14 and x15 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and not x14 and x15 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and x33 and not x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s138;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and not x33 and x4 and x6 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s148;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and not x33 and x4 and not x6 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( x62 and x64 and x9 and not x32 and not x13 and not x33 and not x4 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s149;

      elsif ( x62 and x64 and not x9 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s139;

      elsif ( x62 and not x64 and x66 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x66 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( x62 and not x64 and not x66 and not x7 and x9 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( x62 and not x64 and not x66 and not x7 and not x9 and x10 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x62 and not x64 and not x66 and not x7 and not x9 and x10 and not x6 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x62 and not x64 and not x66 and not x7 and not x9 and not x10 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x64 and not x66 and not x7 and not x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and x64 and x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x64 and x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x64 and x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and not x64 and x65 and x66 and x63 and x30 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and not x64 and x65 and x66 and x63 and not x30 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and x65 and x66 and not x63 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and x11 and x2 ) = '1' then
         y13 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s270;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and x11 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and not x11 and x4 and x12 and x13 and x2 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s271;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and not x11 and x4 and x12 and x13 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and not x11 and x4 and x12 and not x13 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and not x11 and x4 and not x12 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and x3 and not x11 and not x4 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and x11 and x2 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s272;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and x11 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and x12 and x13 and x14 and x2 ) = '1' then
         y3 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s273;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and x12 and x13 and x14 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and x12 and x13 and not x14 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and x12 and x13 and not x14 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and x12 and not x13 and x2 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and x12 and not x13 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and not x12 and x2 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and x4 and not x11 and not x12 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and x6 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and x6 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and x7 and x8 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and x7 and x8 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and x7 and not x8 and x2 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and x7 and not x8 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and not x7 and x8 and x2 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and not x7 and x8 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and not x7 and not x8 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and x5 and not x6 and not x7 and not x8 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and x7 and x9 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and x7 and x9 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and x7 and not x9 and x2 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and x7 and not x9 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and not x7 and x9 and x2 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and not x7 and x9 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and not x7 and not x9 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and x6 and not x7 and not x9 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and x7 and x10 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and x7 and x10 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and x7 and not x10 and x2 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and x7 and not x10 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and not x7 and x10 and x2 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and not x7 and x10 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and not x7 and not x10 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and x15 and not x3 and not x4 and not x5 and not x6 and not x7 and not x10 and not x2 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and not x15 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and not x15 and not x7 and x9 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and not x15 and not x7 and not x9 and x10 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and not x15 and not x7 and not x9 and x10 and not x6 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and not x15 and not x7 and not x9 and not x10 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x64 and x65 and not x66 and x63 and not x15 and not x7 and not x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s43;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and x7 and x9 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and x7 and not x9 ) = '1' then
         y75 <= '1' ;
         current_otherm <= s275;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and x9 and x12 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and x9 and not x12 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and x9 and not x12 and x20 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and x9 and not x12 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and not x9 and x13 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and not x9 and not x13 and x20 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and not x9 and not x13 and x20 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and x8 and not x9 and not x13 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s275;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and x5 and not x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s276;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and x6 and not x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s277;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and x8 and x9 and x5 and x7 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and x8 and x9 and x5 and not x7 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and x8 and x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s275;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and x8 and not x9 and x5 and x7 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and x8 and not x9 and x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and x8 and not x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s275;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and not x8 and x5 and x7 and x9 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and not x8 and x5 and x7 and not x9 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and not x8 and x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s275;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and x11 and not x8 and not x5 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s275;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and x3 and not x6 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s277;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and x67 and not x3 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s283;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and not x67 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and not x67 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and not x67 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x65 and not x66 and not x63 and not x67 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and x66 and x16 and x63 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and not x65 and x66 and x16 and x63 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and not x65 and x66 and x16 and x63 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and x66 and x16 and not x63 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s284;

      elsif ( not x62 and not x64 and not x65 and x66 and not x16 and x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and x66 and not x16 and not x63 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x65 and x66 and not x16 and not x63 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x65 and x66 and not x16 and not x63 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and x66 and not x16 and not x63 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and not x66 and x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x62 and not x64 and not x65 and not x66 and x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x62 and not x64 and not x65 and not x66 and x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and not x66 and x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and x67 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and x67 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and x67 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and x67 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and not x67 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and not x67 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and not x65 and not x66 and not x63 and not x67 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s44 =>
      if ( x62 and x32 and x33 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s285;

      elsif ( x62 and x32 and not x33 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s285;

      elsif ( x62 and x32 and not x33 and not x8 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x62 and not x32 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s285;

      elsif ( x62 and not x32 and not x8 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      else
         y9 <= '1' ;
         current_otherm <= s43;

      end if;

   when s45 =>
      if ( x64 and x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s287;

      elsif ( x64 and not x65 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( not x64 and x65 and x31 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( not x64 and x65 and x31 and not x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s289;

      elsif ( not x64 and x65 and not x31 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s199;

      elsif ( not x64 and x65 and not x31 and not x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      end if;

   when s46 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s291;

   when s47 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s292;

   when s48 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s293;

      elsif ( not x62 and x21 and x20 ) = '1' then
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s294;

      elsif ( not x62 and x21 and not x20 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s295;

      elsif ( not x62 and not x21 and x20 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s296;

      else
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s294;

      end if;

   when s49 =>
      if ( x33 and x32 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s297;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s297;

      end if;

   when s50 =>
      if ( x13 and x10 and x11 and x12 and x4 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( x13 and x10 and x11 and x12 and not x4 ) = '1' then
         current_otherm <= s50;

      elsif ( x13 and x10 and x11 and not x12 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and x10 and x11 and not x12 and not x3 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x13 and x10 and x11 and not x12 and not x3 and not x2 ) = '1' then
         current_otherm <= s50;

      elsif ( x13 and x10 and not x11 and x12 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and x10 and not x11 and x12 and not x3 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x13 and x10 and not x11 and x12 and not x3 and not x2 ) = '1' then
         current_otherm <= s50;

      elsif ( x13 and x10 and not x11 and not x12 and x14 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and x10 and not x11 and not x12 and x14 and not x3 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x13 and x10 and not x11 and not x12 and x14 and not x3 and not x2 ) = '1' then
         current_otherm <= s50;

      elsif ( x13 and x10 and not x11 and not x12 and not x14 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x13 and not x10 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and not x10 and not x3 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x13 and not x10 and not x3 and not x2 ) = '1' then
         current_otherm <= s50;

      elsif ( not x13 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x13 and not x3 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      else
         current_otherm <= s50;

      end if;

   when s51 =>
      if ( x10 and x12 and x4 and x11 and x3 and x13 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x10 and x12 and x4 and x11 and x3 and not x13 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s299;

      elsif ( x10 and x12 and x4 and x11 and not x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and x12 and x4 and not x11 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and x12 and not x4 ) = '1' then
         current_otherm <= s51;

      elsif ( x10 and not x12 and x13 and x11 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s50;

      elsif ( x10 and not x12 and x13 and not x11 and x14 and x4 and x3 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x10 and not x12 and x13 and not x11 and x14 and x4 and not x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and not x12 and x13 and not x11 and x14 and not x4 ) = '1' then
         current_otherm <= s51;

      elsif ( x10 and not x12 and x13 and not x11 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x12 and not x13 and x14 and x4 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and not x12 and not x13 and x14 and not x4 ) = '1' then
         current_otherm <= s51;

      elsif ( x10 and not x12 and not x13 and not x14 ) = '1' then
         current_otherm <= s1;

      else
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s50;

      end if;

   when s52 =>
      if ( x11 and x12 and x2 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( x11 and x12 and not x2 ) = '1' then
         current_otherm <= s52;

      elsif ( x11 and not x12 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and not x12 and not x3 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x11 and x3 ) = '1' then
         current_otherm <= s1;

      else
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      end if;

   when s53 =>
      if ( x12 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( not x12 and x11 and x13 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and x11 and x13 and not x7 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( not x12 and x11 and not x13 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( not x12 and not x11 and x14 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( not x12 and not x11 and not x14 and x7 ) = '1' then
         current_otherm <= s1;

      else
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      end if;

   when s54 =>
      if ( x12 and x11 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x12 and x11 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x12 and x11 and not x3 and not x2 ) = '1' then
         current_otherm <= s54;

      elsif ( x12 and not x11 and x10 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( x12 and not x11 and not x10 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x12 and not x11 and not x10 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x12 and not x11 and not x10 and not x3 and not x2 ) = '1' then
         current_otherm <= s54;

      elsif ( not x12 and x13 and x11 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and x13 and x11 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and x13 and x11 and not x3 and not x2 ) = '1' then
         current_otherm <= s54;

      elsif ( not x12 and x13 and not x11 and x14 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and x13 and not x11 and x14 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and x13 and not x11 and x14 and not x3 and not x2 ) = '1' then
         current_otherm <= s54;

      elsif ( not x12 and x13 and not x11 and not x14 and x10 and x5 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( not x12 and x13 and not x11 and not x14 and x10 and not x5 and x1 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and x13 and not x11 and not x14 and x10 and not x5 and not x1 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and x13 and not x11 and not x14 and not x10 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and x13 and not x11 and not x14 and not x10 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and x13 and not x11 and not x14 and not x10 and not x3 and not x2 ) = '1' then
         current_otherm <= s54;

      elsif ( not x12 and not x13 and x14 and x10 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( not x12 and not x13 and x14 and not x10 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and not x13 and x14 and not x10 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and not x13 and x14 and not x10 and not x3 and not x2 ) = '1' then
         current_otherm <= s54;

      elsif ( not x12 and not x13 and not x14 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and not x13 and not x14 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s54;

      end if;

   when s55 =>
      if ( x12 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( not x12 and x10 and x13 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x12 and x10 and x13 and not x11 and x14 and x6 and x2 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and x10 and x13 and not x11 and x14 and x6 and not x2 ) = '1' then
         current_otherm <= s55;

      elsif ( not x12 and x10 and x13 and not x11 and x14 and not x6 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x12 and x10 and x13 and not x11 and x14 and not x6 and not x2 ) = '1' then
         current_otherm <= s55;

      elsif ( not x12 and x10 and x13 and not x11 and not x14 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( not x12 and x10 and not x13 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      else
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      end if;

   when s56 =>
      if ( x10 and x12 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x10 and not x12 and x11 and x13 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x10 and not x12 and x11 and not x13 and x14 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x10 and not x12 and x11 and not x13 and not x14 and x1 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( x10 and not x12 and x11 and not x13 and not x14 and not x1 and x2 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and not x12 and x11 and not x13 and not x14 and not x1 and not x2 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( x10 and not x12 and not x11 and x13 and x14 and x6 and x2 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x10 and not x12 and not x11 and x13 and x14 and x6 and not x2 ) = '1' then
         current_otherm <= s56;

      elsif ( x10 and not x12 and not x11 and x13 and x14 and not x6 and x2 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x10 and not x12 and not x11 and x13 and x14 and not x6 and not x2 ) = '1' then
         current_otherm <= s56;

      elsif ( x10 and not x12 and not x11 and x13 and not x14 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x10 and not x12 and not x11 and not x13 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      else
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      end if;

   when s57 =>
      if ( x62 and x10 and x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x10 and not x12 and x13 and x11 and x4 and x2 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( x62 and x10 and not x12 and x13 and x11 and x4 and not x2 ) = '1' then
         current_otherm <= s57;

      elsif ( x62 and x10 and not x12 and x13 and x11 and not x4 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x62 and x10 and not x12 and x13 and x11 and not x4 and not x2 ) = '1' then
         current_otherm <= s57;

      elsif ( x62 and x10 and not x12 and x13 and not x11 and x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x10 and not x12 and x13 and not x11 and not x14 and x1 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s50;

      elsif ( x62 and x10 and not x12 and x13 and not x11 and not x14 and not x1 ) = '1' then
         y16 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s298;

      elsif ( x62 and x10 and not x12 and not x13 and x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x10 and not x12 and not x13 and not x14 and x4 and x2 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( x62 and x10 and not x12 and not x13 and not x14 and x4 and not x2 ) = '1' then
         current_otherm <= s57;

      elsif ( x62 and x10 and not x12 and not x13 and not x14 and not x4 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x62 and x10 and not x12 and not x13 and not x14 and not x4 and not x2 ) = '1' then
         current_otherm <= s57;

      elsif ( x62 and not x10 and x4 and x2 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s59;

      elsif ( x62 and not x10 and x4 and not x2 ) = '1' then
         current_otherm <= s57;

      elsif ( x62 and not x10 and not x4 and x2 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s56;

      elsif ( x62 and not x10 and not x4 and not x2 ) = '1' then
         current_otherm <= s57;

      elsif ( not x62 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s58 =>
      if ( x10 and x12 and x11 and x13 and x3 and x6 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s50;

      elsif ( x10 and x12 and x11 and x13 and x3 and not x6 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and x12 and x11 and x13 and not x3 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and x12 and x11 and not x13 and x5 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s52;

      elsif ( x10 and x12 and x11 and not x13 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and x12 and not x11 and x5 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( x10 and x12 and not x11 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and not x12 and x13 and x11 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( x10 and not x12 and x13 and not x11 and x14 and x5 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( x10 and not x12 and x13 and not x11 and x14 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and not x12 and x13 and not x11 and not x14 and x8 and x1 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( x10 and not x12 and x13 and not x11 and not x14 and x8 and not x1 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and not x12 and x13 and not x11 and not x14 and not x8 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( x10 and not x12 and not x13 and x14 and x5 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( x10 and not x12 and not x13 and x14 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and not x12 and not x13 and not x14 and x1 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s52;

      elsif ( x10 and not x12 and not x13 and not x14 and not x1 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x12 and not x13 and not x14 and not x1 and not x3 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      else
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      end if;

   when s59 =>
      if ( x12 and x11 and x10 and x13 and x2 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( x12 and x11 and x10 and x13 and not x2 ) = '1' then
         current_otherm <= s59;

      elsif ( x12 and x11 and x10 and not x13 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( x12 and x11 and not x10 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( x12 and not x11 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and x14 and x11 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and x14 and not x11 and x10 and x13 and x2 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and x14 and not x11 and x10 and x13 and not x2 ) = '1' then
         current_otherm <= s59;

      elsif ( not x12 and x14 and not x11 and x10 and not x13 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and x14 and not x11 and not x10 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and not x14 and x13 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( not x12 and not x14 and not x13 and x10 and x2 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x12 and not x14 and not x13 and x10 and not x2 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      end if;

   when s60 =>
      if ( x62 and x4 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( x62 and x4 and not x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x4 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and x63 and x9 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x9 ) = '1' then
         current_otherm <= s60;

      elsif ( not x62 and not x63 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s61 =>
      if ( x1 and x2 and x3 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x1 and x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s245;

      elsif ( x1 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      else
         y4 <= '1' ;
         current_otherm <= s67;

      end if;

   when s62 =>
         y1 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s301;

   when s63 =>
      if ( x62 and x65 and x20 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y20 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s302;

      elsif ( x62 and x65 and not x20 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s303;

      elsif ( x62 and not x65 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s304;

      elsif ( not x62 and x21 and x20 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s306;

      elsif ( not x62 and x21 and not x20 ) = '1' then
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s305;

      else
         y28 <= '1' ;
         current_otherm <= s306;

      end if;

   when s64 =>
      if ( x2 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( x2 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s19;

      elsif ( not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s66;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s70;

      end if;

   when s65 =>
      if ( x62 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x7 and x9 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x7 and not x9 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x7 and not x9 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s66 =>
      if ( x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s307;

      elsif ( not x3 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( not x3 and x2 and not x1 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s197;

      elsif ( not x3 and not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s66;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      end if;

   when s67 =>
      if ( x62 and x64 and x12 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x62 and x64 and not x12 and x10 and x13 and x11 and x5 and x6 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( x62 and x64 and not x12 and x10 and x13 and x11 and x5 and not x6 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and not x12 and x10 and x13 and x11 and x5 and not x6 and not x7 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( x62 and x64 and not x12 and x10 and x13 and x11 and not x5 and x4 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( x62 and x64 and not x12 and x10 and x13 and x11 and not x5 and not x4 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and x64 and not x12 and x10 and x13 and not x11 and x14 and x4 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( x62 and x64 and not x12 and x10 and x13 and not x11 and x14 and not x4 ) = '1' then
         current_otherm <= s67;

      elsif ( x62 and x64 and not x12 and x10 and x13 and not x11 and not x14 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x62 and x64 and not x12 and x10 and not x13 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x62 and x64 and not x12 and not x10 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x62 and not x64 and x65 and x6 and x3 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and not x64 and x65 and x6 and not x3 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and not x64 and x65 and x6 and not x3 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x62 and not x64 and x65 and not x6 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x62 and not x64 and not x65 and x66 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x65 and x66 and not x5 and x1 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s60;

      elsif ( x62 and not x64 and not x65 and x66 and not x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and x17 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s246;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and x17 and not x6 and x8 and x4 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s126;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and x17 and not x6 and x8 and not x4 and x1 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and x17 and not x6 and x8 and not x4 and x1 and not x3 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and x17 and not x6 and x8 and not x4 and not x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and x17 and not x6 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and x19 and x9 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and x19 and not x9 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and not x19 and x4 and x5 and x3 ) = '1' then
         current_otherm <= s67;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and not x19 and x4 and x5 and not x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and not x19 and x4 and not x5 and x3 ) = '1' then
         current_otherm <= s67;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and not x19 and x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and not x19 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x62 and not x64 and not x65 and not x66 and x18 and not x17 and not x19 and not x4 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x64 and not x65 and not x66 and not x18 and x17 and x12 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x62 and not x64 and not x65 and not x66 and not x18 and x17 and not x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x64 and not x65 and not x66 and not x18 and not x17 and x19 and x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x62 and not x64 and not x65 and not x66 and not x18 and not x17 and x19 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x65 and not x66 and not x18 and not x17 and not x19 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x66 and x12 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s308;

      elsif ( not x62 and x66 and x12 and not x4 and x5 ) = '1' then
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s309;

      elsif ( not x62 and x66 and x12 and not x4 and not x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s95;

      elsif ( not x62 and x66 and not x12 and x4 and x5 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x66 and not x12 and x4 and not x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x66 and not x12 and not x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s310;

      elsif ( not x62 and not x66 and x20 and x21 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x66 and x20 and x21 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x66 and x20 and x21 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x66 and x20 and x21 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x66 and x20 and not x21 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x66 and x20 and not x21 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x66 and x20 and not x21 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x66 and x20 and not x21 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x66 and not x20 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x66 and not x20 and x6 and not x7 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x66 and not x20 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s68 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s311;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and x30 and x36 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and x30 and not x36 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and x33 and x34 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and x33 and not x34 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and x33 and not x34 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and x33 and not x34 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and x33 and not x34 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and not x33 and x35 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and not x33 and not x35 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and not x33 and not x35 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and not x33 and not x35 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and x31 and not x33 and not x35 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and not x31 and x32 ) = '1' then
         y1 <= '1' ;
         y22 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s312;

      elsif ( x62 and not x64 and x65 and x4 and x5 and x6 and not x30 and not x31 and not x32 ) = '1' then
         y1 <= '1' ;
         y20 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s313;

      elsif ( x62 and not x64 and x65 and x4 and x5 and not x6 and x7 and x23 and x24 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s314;

      elsif ( x62 and not x64 and x65 and x4 and x5 and not x6 and x7 and x23 and not x24 ) = '1' then
         y1 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      elsif ( x62 and not x64 and x65 and x4 and x5 and not x6 and x7 and not x23 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      elsif ( x62 and not x64 and x65 and x4 and x5 and not x6 and not x7 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s316;

      elsif ( x62 and not x64 and x65 and x4 and not x5 and x8 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s316;

      elsif ( x62 and not x64 and x65 and x4 and not x5 and not x8 and x9 and x25 and x26 ) = '1' then
         y14 <= '1' ;
         y19 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      elsif ( x62 and not x64 and x65 and x4 and not x5 and not x8 and x9 and x25 and not x26 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      elsif ( x62 and not x64 and x65 and x4 and not x5 and not x8 and x9 and not x25 ) = '1' then
         y14 <= '1' ;
         y17 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      elsif ( x62 and not x64 and x65 and x4 and not x5 and not x8 and not x9 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s316;

      elsif ( x62 and not x64 and x65 and not x4 ) = '1' then
         y1 <= '1' ;
         y33 <= '1' ;
         y37 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s317;

      elsif ( x62 and not x64 and not x65 and x17 and x18 and x7 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s318;

      elsif ( x62 and not x64 and not x65 and x17 and x18 and not x7 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s105;

      elsif ( x62 and not x64 and not x65 and x17 and not x18 ) = '1' then
         current_otherm <= s68;

      elsif ( x62 and not x64 and not x65 and not x17 and x18 and x19 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s104;

      elsif ( x62 and not x64 and not x65 and not x17 and x18 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x65 and not x17 and not x18 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x13 and x14 and x5 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x13 and x14 and not x5 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x13 and x14 and not x5 and not x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x13 and not x14 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x13 and not x14 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and x67 and x11 and x13 and not x14 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and x67 and x11 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and x67 and x11 and not x13 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and x67 and x11 and not x13 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and x67 and not x11 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and x67 and not x11 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and x67 and not x11 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and x10 and x15 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and x10 and x15 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and x10 and x15 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and x10 and not x15 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and x15 and x5 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and x15 and not x5 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and x15 and not x5 and not x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and not x15 and x11 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and not x15 and not x11 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and not x15 and not x11 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and x13 and not x10 and not x15 and not x11 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and not x13 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and x14 and not x13 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and x9 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and x9 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and x9 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and not x9 and x15 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and not x9 and x15 and not x3 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and not x9 and x15 and not x3 and not x2 ) = '1' then
         current_otherm <= s68;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and not x9 and not x15 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x67 and not x14 and not x9 and not x15 and not x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x62 and x63 and not x64 and x66 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and not x64 and x66 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x64 and not x66 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and not x63 and x64 and x65 and x66 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and x67 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and not x67 and x21 and x15 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and not x67 and x21 and not x15 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and not x67 and x21 and not x15 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and not x67 and x21 and not x15 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and not x67 and x21 and not x15 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and not x66 and not x67 and not x21 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s319;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and x19 and x12 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and x19 and not x12 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s254;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and x6 ) = '1' then
         y16 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s255;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and x16 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and x6 ) = '1' then
         y12 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s257;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and x15 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and not x18 and x19 ) = '1' then
         y27 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and not x18 and not x19 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and not x18 and not x19 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and x11 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and not x11 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and x10 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and not x10 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and not x6 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and not x6 and not x12 ) = '1' then
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and x14 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and x13 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and not x6 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and x12 and x6 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s260;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and x12 and not x6 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s261;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and not x12 and x6 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and not x12 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and not x19 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and x24 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and x9 and x10 and x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and x9 and x10 and not x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and x9 and not x10 and x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and x9 and not x10 and not x8 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and not x9 and x10 and x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and not x9 and x10 and not x8 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s23;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and not x9 and not x10 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and x23 and not x9 and not x10 and not x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s320;

      elsif ( not x62 and not x63 and not x64 and x67 and x4 and not x24 and not x23 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and x5 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and x5 and x10 and not x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and x5 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and x5 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and x7 and x8 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and x7 and not x8 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and x7 and not x8 and x10 and not x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and x7 and not x8 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and x7 and not x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and not x7 and x9 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and not x7 and not x9 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and not x7 and not x9 and x10 and not x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and not x7 and not x9 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and x6 and not x5 and not x7 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and not x6 and x7 and x5 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and not x6 and x7 and not x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and not x6 and not x7 and x5 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and x24 and not x6 and not x7 and not x5 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and x23 and not x24 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and x24 and x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and x24 and not x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and x9 and x10 and x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and x9 and x10 and not x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and x9 and not x10 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and x9 and not x10 and not x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and not x9 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and not x9 and x8 and not x10 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and x67 and not x4 and not x23 and not x24 and not x9 and not x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and not x63 and not x64 and not x67 and x30 and x31 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s321;

      elsif ( not x62 and not x63 and not x64 and not x67 and x30 and not x31 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s322;

      else
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s146;

      end if;

   when s69 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y14 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s323;

   when s70 =>
      if ( x62 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and not x3 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( x62 and not x3 and x1 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s66;

      elsif ( x62 and not x3 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x62 and x63 and x66 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y15 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s324;

      elsif ( not x62 and x63 and not x66 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s325;

      elsif ( not x62 and not x63 and x64 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s326;

      elsif ( not x62 and not x63 and not x64 and x66 and x67 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s327;

      elsif ( not x62 and not x63 and not x64 and x66 and not x67 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s328;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s325;

      end if;

   when s71 =>
      if ( x62 and x6 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( x62 and not x6 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( not x62 and x64 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s329;

      elsif ( not x62 and not x64 and x65 and x15 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x64 and x65 and not x15 and x6 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x64 and x65 and not x15 and not x6 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( not x62 and not x64 and not x65 and x10 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x64 and not x65 and not x10 and x11 ) = '1' then
         y14 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s163;

      else
         y10 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s164;

      end if;

   when s72 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s330;

      elsif ( x62 and not x64 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      elsif ( not x62 and x63 and x67 and x11 and x14 and x13 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x62 and x63 and x67 and x11 and x14 and x13 and not x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x62 and x63 and x67 and x11 and x14 and not x13 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and x67 and x11 and x14 and not x13 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and x11 and x14 and not x13 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and x11 and x14 and not x13 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and x11 and not x14 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and x67 and x11 and not x14 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and x11 and not x14 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and x11 and not x14 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and not x11 and x10 and x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x67 and not x11 and x10 and not x13 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and x67 and not x11 and x10 and not x13 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and not x11 and x10 and not x13 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and not x11 and x10 and not x13 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and not x11 and not x10 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and x67 and not x11 and not x10 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and x67 and not x11 and not x10 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and not x11 and not x10 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and not x67 and x13 and x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and x15 and x14 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and x15 and x14 and not x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and x15 and not x14 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and x15 and not x14 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and x15 and not x14 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and x15 and not x14 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and not x15 and x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and not x15 and not x11 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and not x15 and not x11 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and not x15 and not x11 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and not x67 and x13 and not x10 and not x15 and not x11 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and not x67 and not x13 and x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x62 and x63 and not x67 and not x13 and x4 and not x2 ) = '1' then
         current_otherm <= s72;

      elsif ( not x62 and x63 and not x67 and not x13 and not x4 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and not x67 and not x13 and not x4 and not x2 ) = '1' then
         current_otherm <= s72;

      else
         y12 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s332;

      end if;

   when s73 =>
      if ( x13 and x67 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and x67 and not x14 and x11 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x13 and x67 and not x14 and not x11 and x10 and x6 and x2 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( x13 and x67 and not x14 and not x11 and x10 and x6 and not x2 ) = '1' then
         current_otherm <= s73;

      elsif ( x13 and x67 and not x14 and not x11 and x10 and not x6 and x2 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x13 and x67 and not x14 and not x11 and x10 and not x6 and not x2 ) = '1' then
         current_otherm <= s73;

      elsif ( x13 and x67 and not x14 and not x11 and not x10 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and not x67 and x15 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and not x67 and x15 and not x14 and x10 and x6 and x2 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( x13 and not x67 and x15 and not x14 and x10 and x6 and not x2 ) = '1' then
         current_otherm <= s73;

      elsif ( x13 and not x67 and x15 and not x14 and x10 and not x6 and x2 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x13 and not x67 and x15 and not x14 and x10 and not x6 and not x2 ) = '1' then
         current_otherm <= s73;

      elsif ( x13 and not x67 and x15 and not x14 and not x10 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x13 and not x67 and not x15 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      else
         y5 <= '1' ;
         current_otherm <= s68;

      end if;

   when s74 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s334;

      elsif ( x62 and not x64 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s335;

      elsif ( not x62 and x63 and x67 and x14 and x13 and x11 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and x10 and x4 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and x10 and not x4 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and not x10 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and not x10 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and not x10 and not x3 and not x2 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and x67 and x14 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and x14 and not x13 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and x14 and not x13 and not x3 and not x2 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and x67 and not x14 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and not x14 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and x67 and not x14 and not x3 and not x2 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and x14 and x10 and x4 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and x14 and x10 and not x4 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and x14 and not x10 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and not x14 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and not x14 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and not x14 and not x3 and not x2 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and not x67 and x15 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and x15 and not x13 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and not x67 and x15 and not x13 and not x3 and not x2 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and x63 and not x67 and not x15 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and not x15 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( not x62 and x63 and not x67 and not x15 and not x3 and not x2 ) = '1' then
         current_otherm <= s74;

      elsif ( not x62 and not x63 and x64 and x21 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s336;

      elsif ( not x62 and not x63 and x64 and not x21 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s337;

      else
         y33 <= '1' ;
         current_otherm <= s321;

      end if;

   when s75 =>
      if ( x13 and x67 and x11 and x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x67 and x11 and not x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( x13 and x67 and not x11 and x10 and x4 and x3 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( x13 and x67 and not x11 and x10 and x4 and x3 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( x13 and x67 and not x11 and x10 and x4 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x13 and x67 and not x11 and x10 and not x4 ) = '1' then
         current_otherm <= s75;

      elsif ( x13 and x67 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x67 and x15 and x10 and x4 and x3 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( x13 and not x67 and x15 and x10 and x4 and x3 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s76;

      elsif ( x13 and not x67 and x15 and x10 and x4 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x13 and not x67 and x15 and x10 and not x4 ) = '1' then
         current_otherm <= s75;

      elsif ( x13 and not x67 and x15 and not x10 and x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x67 and x15 and not x10 and not x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( x13 and not x67 and not x15 and x11 and x4 and x14 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x13 and not x67 and not x15 and x11 and x4 and not x14 and x3 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s338;

      elsif ( x13 and not x67 and not x15 and x11 and x4 and not x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x13 and not x67 and not x15 and x11 and not x4 ) = '1' then
         current_otherm <= s75;

      elsif ( x13 and not x67 and not x15 and not x11 and x10 and x4 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x13 and not x67 and not x15 and not x11 and x10 and not x4 ) = '1' then
         current_otherm <= s75;

      elsif ( x13 and not x67 and not x15 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         current_otherm <= s74;

      end if;

   when s76 =>
      if ( x67 and x11 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( x67 and not x11 and x13 and x14 and x10 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( x67 and not x11 and x13 and x14 and not x10 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( x67 and not x11 and x13 and x14 and not x10 and not x1 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x67 and not x11 and x13 and x14 and not x10 and not x1 and not x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x67 and not x11 and x13 and not x14 and x10 and x6 and x2 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( x67 and not x11 and x13 and not x14 and x10 and x6 and not x2 ) = '1' then
         current_otherm <= s76;

      elsif ( x67 and not x11 and x13 and not x14 and x10 and not x6 and x2 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( x67 and not x11 and x13 and not x14 and x10 and not x6 and not x2 ) = '1' then
         current_otherm <= s76;

      elsif ( x67 and not x11 and x13 and not x14 and not x10 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( x67 and not x11 and not x13 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x67 and x10 and x13 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x67 and x10 and x13 and not x14 and x15 and x6 and x2 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( not x67 and x10 and x13 and not x14 and x15 and x6 and not x2 ) = '1' then
         current_otherm <= s76;

      elsif ( not x67 and x10 and x13 and not x14 and x15 and not x6 and x2 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( not x67 and x10 and x13 and not x14 and x15 and not x6 and not x2 ) = '1' then
         current_otherm <= s76;

      elsif ( not x67 and x10 and x13 and not x14 and not x15 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x67 and x10 and not x13 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x67 and not x10 and x11 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x67 and not x10 and not x11 and x13 and x14 and x15 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x67 and not x10 and not x11 and x13 and x14 and not x15 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x67 and not x10 and not x11 and x13 and x14 and not x15 and not x1 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x67 and not x10 and not x11 and x13 and x14 and not x15 and not x1 and not x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( not x67 and not x10 and not x11 and x13 and not x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      else
         y5 <= '1' ;
         current_otherm <= s331;

      end if;

   when s77 =>
      if ( x13 and x67 and x11 and x14 and x8 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and x67 and x11 and x14 and x8 and not x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and x67 and x11 and x14 and not x8 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and x67 and x11 and not x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( x13 and x67 and not x11 and x10 and x14 and x3 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( x13 and x67 and not x11 and x10 and x14 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and x67 and not x11 and x10 and x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and x67 and not x11 and x10 and not x14 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( x13 and x67 and not x11 and x10 and not x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and x67 and not x11 and not x10 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s78;

      elsif ( x13 and x67 and not x11 and not x10 and not x1 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x67 and not x11 and not x10 and not x1 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and x15 and x10 and x14 and x3 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( x13 and not x67 and x15 and x10 and x14 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and x15 and x10 and x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and x15 and x10 and not x14 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( x13 and not x67 and x15 and x10 and not x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and x15 and not x10 and x14 and x8 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and not x67 and x15 and not x10 and x14 and x8 and not x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and x15 and not x10 and x14 and not x8 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and not x67 and x15 and not x10 and not x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( x13 and not x67 and not x15 and x11 and x5 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and not x67 and not x15 and x11 and x5 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s78;

      elsif ( x13 and not x67 and not x15 and x11 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and not x15 and not x11 and x10 and x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x13 and not x67 and not x15 and not x11 and x10 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( x13 and not x67 and not x15 and not x11 and not x10 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s78;

      elsif ( x13 and not x67 and not x15 and not x11 and not x10 and not x1 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x67 and not x15 and not x11 and not x10 and not x1 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      else
         y5 <= '1' ;
         current_otherm <= s72;

      end if;

   when s78 =>
      if ( x67 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x67 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x67 and x11 and x14 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x67 and x11 and x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x67 and x11 and not x14 and x2 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x67 and x11 and not x14 and not x2 ) = '1' then
         current_otherm <= s78;

      elsif ( not x67 and not x11 and x3 ) = '1' then
         current_otherm <= s1;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      end if;

   when s79 =>
      if ( x64 and x65 and x4 and x5 and x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and x65 and x4 and x5 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x64 and x65 and x4 and x5 and not x3 and not x6 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x64 and x65 and x4 and x5 and not x3 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s340;

      elsif ( x64 and x65 and x4 and not x5 and x3 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x64 and x65 and x4 and not x5 and not x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x64 and x65 and x4 and not x5 and not x3 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x64 and x65 and x4 and not x5 and not x3 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x65 and not x4 and x5 and x3 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x64 and x65 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x65 and not x4 and not x5 and x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x65 and not x4 and not x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and not x65 and x13 and x10 and x67 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and x13 and x10 and not x67 and x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and x13 and x10 and not x67 and not x2 and x15 ) = '1' then
         current_otherm <= s79;

      elsif ( x64 and not x65 and x13 and x10 and not x67 and not x2 and not x15 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and x13 and not x10 and x11 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and x13 and not x10 and not x11 and x67 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x64 and not x65 and x13 and not x10 and not x11 and x67 and not x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and x13 and not x10 and not x11 and not x67 and x15 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and x13 and not x10 and not x11 and not x67 and not x15 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( x64 and not x65 and x13 and not x10 and not x11 and not x67 and not x15 and not x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x65 and not x13 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      else
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s343;

      end if;

   when s80 =>
      if ( x22 and x23 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x22 and not x23 and x16 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x22 and not x23 and x16 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x22 and not x23 and x16 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x22 and not x23 and x16 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x22 and not x23 and x16 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x22 and not x23 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s344;

      elsif ( not x22 and x23 and x16 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( not x22 and x23 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s344;

      else
         y6 <= '1' ;
         current_otherm <= s39;

      end if;

   when s81 =>
      if ( x22 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s345;

      else
         y6 <= '1' ;
         current_otherm <= s346;

      end if;

   when s82 =>
      if ( x62 and x5 and x4 and x2 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x62 and x5 and x4 and not x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s221;

      elsif ( x62 and x5 and not x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s214;

      elsif ( x62 and not x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s214;

      elsif ( not x62 and x63 and x15 and x16 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and x15 and x16 and not x1 and x5 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( not x62 and x63 and x15 and x16 and not x1 and not x5 and x6 and x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and x15 and x16 and not x1 and not x5 and x6 and x2 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x15 and x16 and not x1 and not x5 and x6 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x15 and x16 and not x1 and not x5 and not x6 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x62 and x63 and x15 and not x16 and x7 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x62 and x63 and x15 and not x16 and not x7 and x9 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x62 and x63 and x15 and not x16 and not x7 and not x9 and x10 and x6 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and x63 and x15 and not x16 and not x7 and not x9 and x10 and not x6 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and x63 and x15 and not x16 and not x7 and not x9 and not x10 and x11 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and x15 and not x16 and not x7 and not x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and x16 and x5 and x4 and x2 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x63 and not x15 and x16 and x5 and x4 and not x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and x63 and not x15 and x16 and x5 and not x4 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and x16 and not x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and x11 and x2 ) = '1' then
         y13 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s270;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and x11 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and not x11 and x4 and x12 and x13 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and not x11 and x4 and x12 and x13 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and not x11 and x4 and x12 and not x13 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and not x11 and x4 and not x12 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and x3 and not x11 and not x4 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and x11 and x2 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s272;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and x11 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and x12 and x13 and x14 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s349;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and x12 and x13 and x14 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and x12 and x13 and not x14 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and x12 and x13 and not x14 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and x12 and not x13 and x2 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and x12 and not x13 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and not x12 and x2 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and x4 and not x11 and not x12 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and x6 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and x6 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and x7 and x8 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and x7 and x8 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and x7 and not x8 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and x7 and not x8 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and not x7 and x8 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and not x7 and x8 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and not x7 and not x8 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and x5 and not x6 and not x7 and not x8 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and x7 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and x7 and x9 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and x7 and not x9 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and x7 and not x9 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and not x7 and x9 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and not x7 and x9 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and not x7 and not x9 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and x6 and not x7 and not x9 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and x7 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and x7 and x10 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and x7 and not x10 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and x7 and not x10 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and not x7 and x10 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and not x7 and x10 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and not x7 and not x10 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x63 and not x15 and not x16 and not x3 and not x4 and not x5 and not x6 and not x7 and not x10 and not x2 ) = '1' then
         current_otherm <= s82;

      elsif ( not x62 and not x63 and x18 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      else
         y11 <= '1' ;
         current_otherm <= s350;

      end if;

   when s83 =>
         y2 <= '1' ;
         current_otherm <= s351;

   when s84 =>
         y19 <= '1' ;
         current_otherm <= s13;

   when s85 =>
         y1 <= '1' ;
         current_otherm <= s17;

   when s86 =>
         y5 <= '1' ;
         current_otherm <= s352;

   when s87 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s353;

   when s88 =>
      if ( x63 and x13 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( x63 and not x13 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and not x13 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and not x13 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x13 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s89 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s87;

      elsif ( not x62 and x63 and x31 and x30 and x8 ) = '1' then
         y42 <= '1' ;
         current_otherm <= s354;

      elsif ( not x62 and x63 and x31 and x30 and not x8 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s355;

      elsif ( not x62 and x63 and x31 and not x30 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and x31 and not x30 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x31 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and not x31 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x28 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x65 and x28 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x65 and x28 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x28 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x28 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s356;

      elsif ( not x62 and not x63 and not x64 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x63 and not x64 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x63 and not x64 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s90 =>
      if ( x65 and x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x65 and x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x65 and x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and x63 and x66 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x65 and not x62 and x63 and x66 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x65 and not x62 and x63 and not x66 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s343;

      elsif ( x65 and not x62 and not x63 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x65 and not x62 and not x63 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x65 and not x62 and not x63 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x62 and not x63 and not x66 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s356;

      elsif ( not x65 and x62 and x17 and x18 and x5 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x65 and x62 and x17 and x18 and not x5 and x6 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and x17 and x18 and not x5 and not x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x62 and x17 and not x18 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x65 and x62 and x17 and not x18 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x62 and not x17 and x18 and x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x62 and not x17 and x18 and not x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x65 and x62 and not x17 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and x63 and x9 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s357;

      elsif ( not x65 and not x62 and x63 and not x9 ) = '1' then
         current_otherm <= s90;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and x19 and x12 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and x19 and not x12 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s254;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and x12 and x6 ) = '1' then
         y16 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s255;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and x12 and not x6 and x16 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and x12 and not x6 and not x16 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and not x12 and x6 ) = '1' then
         y12 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s257;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and not x12 and not x6 and x15 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and not x18 and x19 ) = '1' then
         y27 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and not x18 and not x19 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and x5 and not x18 and not x19 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and x12 and x11 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and x12 and not x11 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and not x12 and x10 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and x6 and not x12 and not x10 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and not x6 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and x19 and not x6 and not x12 ) = '1' then
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s112;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and x12 and x14 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and x12 and not x14 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and not x12 and x13 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and x18 and not x19 and not x6 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and not x18 and x19 and x12 and x6 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s260;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and not x18 and x19 and x12 and not x6 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s261;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and not x18 and x19 and not x12 and x6 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and not x18 and x19 and not x12 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x65 and not x62 and not x63 and x66 and x8 and not x5 and not x18 and not x19 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x65 and not x62 and not x63 and x66 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      else
         y7 <= '1' ;
         current_otherm <= s45;

      end if;

   when s91 =>
      if ( x63 and x12 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( x63 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s358;

      end if;

   when s92 =>
      if ( x62 and x20 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x20 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x20 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x20 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x20 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s359;

      elsif ( not x62 and x63 and x65 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x65 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x65 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x65 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x67 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s361;

      elsif ( not x62 and x63 and not x65 and not x67 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x63 and not x65 and not x67 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x63 and not x65 and not x67 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and not x67 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and not x63 and x64 and not x66 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and not x63 and x64 and not x66 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x63 and not x64 and x66 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x63 and not x64 and x66 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x63 and not x64 and x66 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x66 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x66 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x66 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s93 =>
      if ( x21 and x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s362;

      elsif ( x21 and not x20 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s296;

      elsif ( not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s94 =>
      if ( x62 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s63;

      elsif ( not x62 and x63 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and x64 and x21 and x20 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s363;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and x17 and x16 and x19 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and x17 and x16 and x19 and not x11 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and x17 and x16 and not x19 and x18 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and x17 and x16 and not x19 and not x18 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and x17 and not x16 and x11 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and x17 and not x16 and not x11 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s365;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and not x17 and x16 and x19 and x14 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and not x17 and x16 and x19 and not x14 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and not x17 and x16 and not x19 and x13 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and not x17 and x16 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 and not x12 and not x17 and not x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and x64 and not x21 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      elsif ( not x62 and not x63 and not x64 and x24 and x23 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x24 and x23 and x10 and not x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x24 and x23 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and x23 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and x6 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and x10 and not x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and x13 and x14 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and x13 and not x14 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and x13 and not x14 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and x13 and not x14 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and x13 and not x14 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and not x13 and x15 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and not x13 and not x15 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and not x13 and not x15 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and not x13 and not x15 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and x9 and not x10 and not x13 and not x15 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and x17 and x18 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and x17 and not x18 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and x17 and not x18 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and x17 and not x18 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and x17 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and not x17 and x19 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and not x17 and not x19 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and not x17 and not x19 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and not x17 and not x19 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and x16 and not x17 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and x7 and not x9 and not x16 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x62 and not x63 and not x64 and x24 and not x23 and not x6 and not x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and not x64 and not x24 and x6 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s167;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and x9 and x10 and x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and x9 and x10 and not x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and x9 and not x10 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and x9 and not x10 and not x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and not x9 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and not x9 and x8 and not x10 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and not x24 and not x6 and x7 and not x23 and not x9 and not x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      else
         y16 <= '1' ;
         current_otherm <= s14;

      end if;

   when s95 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s366;

      elsif ( not x62 and x63 and x31 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and x31 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x31 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and not x31 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and x64 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x21 and x9 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and not x63 and x64 and not x66 and x21 and not x9 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x63 and x64 and not x66 and x21 and not x9 and x6 and not x7 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and not x63 and x64 and not x66 and x21 and not x9 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x21 and not x9 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x21 and x5 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s185;

      elsif ( not x62 and not x63 and x64 and not x66 and not x21 and not x5 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s363;

      elsif ( not x62 and not x63 and not x64 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s96 =>
      if ( x62 and x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      elsif ( x62 and not x12 ) = '1' then
         current_otherm <= s96;

      elsif ( not x62 and x15 and x13 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and x15 and not x13 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      elsif ( not x62 and not x15 and x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      else
         current_otherm <= s96;

      end if;

   when s97 =>
      if ( x62 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x62 and not x6 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x15 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s102;

      elsif ( not x62 and not x15 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      else
         y10 <= '1' ;
         current_otherm <= s16;

      end if;

   when s98 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s367;

   when s99 =>
      if ( x63 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x63 and x1 and not x2 and x5 and x3 ) = '1' then
         current_otherm <= s99;

      elsif ( x63 and x1 and not x2 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x63 and x1 and not x2 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( x63 and not x1 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x63 and x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x31 and x14 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x64 and x31 and not x14 ) = '1' then
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y69 <= '1' ;
         current_otherm <= s368;

      elsif ( not x63 and not x64 and not x31 and x14 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s287;

      else
         y37 <= '1' ;
         current_otherm <= s181;

      end if;

   when s100 =>
      if ( x63 and x11 ) = '1' then
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s369;

      elsif ( x63 and not x11 ) = '1' then
         y10 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s370;

      elsif ( not x63 and x64 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s371;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s372;

      end if;

   when s101 =>
      if ( x62 and x64 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s373;

      elsif ( x62 and x64 and not x17 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s374;

      elsif ( x62 and not x64 and x25 and x9 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      elsif ( x62 and not x64 and x25 and not x9 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( x62 and not x64 and not x25 and x13 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( x62 and not x64 and not x25 and not x13 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

      else
         y13 <= '1' ;
         current_otherm <= s375;

      end if;

   when s102 =>
      if ( x62 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x62 and not x6 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x15 and x6 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      else
         y10 <= '1' ;
         current_otherm <= s16;

      end if;

   when s103 =>
      if ( x62 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and x65 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x64 and x63 and x65 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x64 and x63 and x65 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and x65 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and not x65 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x64 and x63 and not x65 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x64 and x63 and not x65 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and not x65 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and x7 and x9 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and x7 and not x9 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and x9 and x11 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and x9 and not x11 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and x9 and not x11 and x14 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and x9 and not x11 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and not x9 and not x10 and x14 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and not x9 and not x10 and x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and x8 and not x9 and not x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and not x8 and x9 ) = '1' then
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s158;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and x3 and not x7 and not x8 and not x9 ) = '1' then
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s380;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and x15 and x16 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and x15 and x16 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and x15 and x16 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and x15 and x16 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and x15 and not x16 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and not x15 and x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and x9 and not x15 and not x7 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s381;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and x15 and x17 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and x15 and not x17 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and x15 and not x17 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and x15 and not x17 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and x15 and not x17 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and not x15 and x7 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and x8 and not x9 and not x15 and not x7 ) = '1' then
         y22 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s382;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and x15 and x18 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and x15 and not x18 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and x15 and not x18 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and x15 and not x18 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and x15 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and not x15 and x7 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and x9 and not x15 and not x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and x15 and x18 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and x15 and x18 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and x15 and x18 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and x15 and x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and x15 and not x18 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and not x15 and x7 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( not x62 and x64 and not x63 and x65 and x6 and not x3 and not x8 and not x9 and not x15 and not x7 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and x3 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and not x3 and x12 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s308;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and not x3 and x12 and not x4 and x5 ) = '1' then
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s309;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and not x3 and x12 and not x4 and not x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s95;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and not x3 and not x12 and x4 and x5 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and not x3 and not x12 and x4 and not x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x64 and not x63 and x65 and not x6 and not x3 and not x12 and not x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s310;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and x63 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and x63 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x65 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s383;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s104 =>
      if ( x17 and x18 and x5 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x17 and x18 and not x5 and x6 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x17 and x18 and not x5 and not x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x17 and not x18 and x14 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x17 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x17 and x6 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s126;

      else
         y7 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s105;

      end if;

   when s105 =>
      if ( x17 and x18 and x6 and x9 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s246;

      elsif ( x17 and x18 and x6 and not x9 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x17 and x18 and not x6 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s104;

      elsif ( x17 and not x18 and x10 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x17 and not x18 and not x10 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( not x17 and x8 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      else
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s126;

      end if;

   when s106 =>
      if ( x62 and x66 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s384;

      elsif ( x62 and x66 and not x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x66 and x17 and x18 and x5 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x62 and not x66 and x17 and x18 and not x5 and x6 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and not x66 and x17 and x18 and not x5 and not x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x62 and not x66 and x17 and not x18 and x9 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x66 and x17 and not x18 and x9 and not x10 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and not x66 and x17 and not x18 and not x9 and x6 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x62 and not x66 and x17 and not x18 and not x9 and not x6 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x66 and not x17 and x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and x7 and x2 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and x7 and x2 and not x3 and x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and x7 and x2 and not x3 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and x7 and not x2 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and not x7 and x8 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and not x7 and not x8 and x2 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and not x7 and not x8 and x2 and not x3 and x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and not x7 and not x8 and x2 and not x3 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x66 and not x17 and not x18 and x6 and not x7 and not x8 and not x2 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x62 and not x66 and not x17 and not x18 and not x6 and x2 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( x62 and not x66 and not x17 and not x18 and not x6 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x67 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( not x62 and x63 and not x67 and x29 and x5 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x63 and not x67 and x29 and x5 and not x4 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x62 and x63 and not x67 and x29 and not x5 and x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x63 and not x67 and x29 and not x5 and not x4 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s287;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and x31 and x15 and x5 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and x31 and x15 and not x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and x31 and not x15 and x16 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and x31 and not x15 and not x16 and x5 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and x31 and not x15 and not x16 and not x5 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and not x31 and x5 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and x4 and not x31 and not x5 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and not x4 and x5 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s385;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and not x4 and not x5 and x31 and x15 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and not x4 and not x5 and x31 and not x15 and x16 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and not x4 and not x5 and x31 and not x15 and not x16 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s386;

      elsif ( not x62 and x63 and not x67 and not x29 and x30 and not x4 and not x5 and not x31 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and x5 and x31 and x4 and x13 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and x5 and x31 and x4 and not x13 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and x5 and x31 and not x4 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and x5 and not x31 and x4 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and x5 and not x31 and x4 and not x8 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and x5 and not x31 and not x4 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s95;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and x31 and x4 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and x31 and x4 and not x8 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and x31 and not x4 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s95;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and not x31 and x4 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and not x31 and not x4 and x9 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and not x31 and not x4 and not x9 and x7 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( not x62 and x63 and not x67 and not x29 and not x30 and not x5 and not x31 and not x4 and not x9 and not x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and x64 and x65 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and x19 and x12 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s387;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and x19 and not x12 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s388;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and x12 and x6 ) = '1' then
         y50 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s389;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and x12 and not x6 and x16 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and x12 and not x6 and not x16 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and not x12 and x6 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s337;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and not x12 and not x6 and x15 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and not x18 and x19 ) = '1' then
         y27 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and not x18 and not x19 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and x5 and not x18 and not x19 and not x6 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and x12 and x11 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s390;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and x12 and not x11 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and not x12 and x10 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s390;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and x6 and not x12 and not x10 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and not x6 and x12 ) = '1' then
         y59 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and x19 and not x6 and not x12 ) = '1' then
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and x12 and x14 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and x12 and not x14 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and not x12 and x13 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and x18 and not x19 and not x6 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and not x18 and x19 and x12 and x6 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and not x18 and x19 and x12 and not x6 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and not x18 and x19 and not x12 and x6 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and not x18 and x19 and not x12 and not x6 ) = '1' then
         y42 <= '1' ;
         current_otherm <= s354;

      elsif ( not x62 and not x63 and x64 and not x65 and x7 and not x5 and not x18 and not x19 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and x64 and not x65 and not x7 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and x23 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and x23 and not x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and not x23 and x5 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and not x23 and x5 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and not x23 and x5 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and not x23 and x5 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x3 and x24 and not x23 and not x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and x5 and x11 and x12 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and x5 and x11 and x12 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and x5 and x11 and not x12 and x13 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and x5 and x11 and not x12 and x13 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and x5 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and x5 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x3 and not x24 and not x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      else
         y5 <= '1' ;
         current_otherm <= s68;

      end if;

   when s107 =>
      if ( x62 and x24 and x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x62 and x24 and x2 and not x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x62 and x24 and not x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x62 and not x24 and x2 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x62 and not x24 and not x2 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x62 and not x24 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x62 and x63 and x64 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x63 and x64 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x63 and x64 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x64 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      end if;

   when s108 =>
      if ( x63 and x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x21 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x21 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( not x63 and x65 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s393;

      elsif ( not x63 and not x65 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x65 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x65 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         y53 <= '1' ;
         current_otherm <= s394;

      end if;

   when s109 =>
      if ( x63 and x16 ) = '1' then
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s395;

      elsif ( x63 and not x16 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and not x16 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x16 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s110 =>
      if ( x65 ) = '1' then
         y4 <= '1' ;
         y20 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s396;

      elsif ( not x65 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x65 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s111 =>
      if ( x64 and x63 and x21 and x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s397;

      elsif ( x64 and x63 and x21 and not x20 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s63;

      elsif ( x64 and x63 and not x21 and x20 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( x64 and x63 and not x21 and not x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s397;

      elsif ( x64 and not x63 and x65 and x67 and x21 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s398;

      elsif ( x64 and not x63 and x65 and x67 and not x21 and x20 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s398;

      elsif ( x64 and not x63 and x65 and x67 and not x21 and not x20 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x63 and x65 and not x67 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and x66 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s399;

      elsif ( not x64 and x63 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and x23 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and x23 and x10 and not x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and x23 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and x23 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and x10 and not x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and x13 and x14 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and x13 and not x14 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and x13 and not x14 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and x13 and not x14 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and x13 and not x14 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and not x13 and x15 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and not x13 and not x15 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and not x13 and not x15 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and not x13 and not x15 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and x9 and not x10 and not x13 and not x15 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and x17 and x18 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and x17 and not x18 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and x17 and not x18 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and x17 and not x18 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and x17 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and not x17 and x19 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and not x17 and not x19 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and not x17 and not x19 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and not x17 and not x19 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and x16 and not x17 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and x7 and not x9 and not x16 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x64 and not x63 and x66 and x67 and x24 and not x23 and not x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s167;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and x9 and x10 and x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and x9 and x10 and not x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and x9 and not x10 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and x9 and not x10 and not x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and not x9 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and not x9 and x8 and not x10 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and x7 and not x23 and not x9 and not x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( not x64 and not x63 and x66 and x67 and not x24 and not x7 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and not x63 and x66 and not x67 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x63 and x66 and not x67 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x63 and x66 and not x67 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x66 and not x67 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and not x66 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and not x63 and not x66 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and not x63 and not x66 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s112 =>
      if ( x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s113 =>
      if ( x62 and x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s400;

      elsif ( x62 and not x33 and x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s400;

      elsif ( x62 and not x33 and not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and not x33 and not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and not x33 and not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x33 and not x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s114 =>
      if ( x62 and x14 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x62 and not x14 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and not x14 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and not x14 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x14 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x63 and x64 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x63 and x64 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x64 and x65 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x64 and x65 and not x18 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( not x62 and x63 and not x64 and not x65 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x62 and x63 and not x64 and not x65 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x62 and x63 and not x64 and not x65 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x64 and not x65 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x13 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s401;

      elsif ( not x62 and not x63 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s115 =>
      if ( x63 and x64 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x63 and x64 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x63 and x64 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x64 and x67 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s402;

      elsif ( x63 and not x64 and not x67 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x64 and not x67 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x64 and not x67 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x64 and not x67 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x64 and not x67 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x66 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and not x66 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and not x66 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s116 =>
      if ( x62 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s385;

      elsif ( not x62 and x64 and not x63 and x67 ) = '1' then
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s403;

      elsif ( not x62 and x64 and not x63 and not x67 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x67 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x67 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x67 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and not x64 and x63 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and not x64 and x63 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and not x64 and x63 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and not x64 and x63 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and not x64 and x63 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x65 and x67 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and not x63 and x65 and x67 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and not x63 and x65 and x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x65 and x67 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x65 and not x67 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s406;

      elsif ( not x62 and not x64 and not x63 and not x65 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and not x63 and not x65 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x64 and not x63 and not x65 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s117 =>
      if ( x62 and x64 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x64 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x64 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x67 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and not x63 and x64 and not x66 and x67 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and not x63 and x64 and not x66 and x67 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x67 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and x12 and x11 and x6 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s407;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and x12 and x11 and not x6 and x10 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and x12 and x11 and not x6 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and x12 and not x11 and x6 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and x12 and not x11 and not x6 and x10 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s409;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and x12 and not x11 and not x6 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and x11 and x6 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s410;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and x11 and not x6 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and x11 and not x6 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and x6 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and x6 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and x6 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and x6 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and not x6 and x10 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and not x6 and not x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and not x6 and not x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and not x6 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x67 and not x12 and not x11 and not x6 and not x10 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and x23 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x67 and x23 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x67 and x23 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and x23 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x67 and x30 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s413;

      elsif ( not x62 and not x63 and not x64 and not x67 and not x30 and x4 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x67 and not x30 and x4 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x67 and not x30 and x4 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x67 and not x30 and x4 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         current_otherm <= s366;

      end if;

   when s118 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x66 and x67 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x66 and x67 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x66 and x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x66 and x67 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x66 and not x67 and x28 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x66 and not x67 and x28 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x66 and not x67 and x28 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x66 and not x67 and x28 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x66 and not x67 and not x28 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s237;

      elsif ( not x63 and not x64 and not x66 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and not x64 and not x66 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and not x64 and not x66 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s119 =>
      if ( x63 and x64 and x65 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x64 and x65 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x64 and x65 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x65 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and not x65 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and x64 and not x65 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and x64 and not x65 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and not x65 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x64 and x65 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x63 and not x64 and x65 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x63 and not x64 and not x65 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s414;

      elsif ( not x63 and x64 and not x65 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x19 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x63 and not x64 and not x19 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x19 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x19 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s120 =>
      if ( x64 and x62 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x64 and x62 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x64 and x62 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and x62 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x64 and not x62 and x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x64 and not x62 and x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and not x63 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x64 and not x62 and not x63 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x64 and not x62 and not x63 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and not x63 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x62 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x65 and x63 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x64 and not x62 and x65 and not x63 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s415;

      elsif ( not x64 and not x62 and not x65 and x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x64 and not x62 and not x65 and x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x64 and not x62 and not x65 and x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and x18 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and not x18 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and not x18 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and not x18 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s121 =>
      if ( x62 and x64 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x64 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x64 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x64 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and not x64 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x64 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x66 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x63 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and x63 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x67 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s416;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x65 and not x66 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x65 and not x66 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x65 and not x66 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s122 =>
      if ( x62 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and x63 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x65 and x64 and x63 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x65 and x64 and x63 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and x63 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and not x63 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x65 and not x64 and x63 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x62 and x65 and not x64 and not x63 and x67 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and not x67 and x4 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x65 and not x64 and not x63 and not x67 and x4 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x65 and not x64 and not x63 and not x67 and x4 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and not x67 and x4 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and not x67 and not x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s352;

      elsif ( not x62 and not x65 and x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and not x63 and x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x65 and not x63 and x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x65 and not x63 and x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and not x63 and x64 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and not x63 and not x64 and x66 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x65 and not x63 and not x64 and x66 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x65 and not x63 and not x64 and x66 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and not x63 and not x64 and x66 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x65 and not x63 and not x64 and x66 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and not x63 and not x64 and not x66 and x20 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and not x65 and not x63 and not x64 and not x66 and not x20 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x65 and not x63 and not x64 and not x66 and not x20 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x65 and not x63 and not x64 and not x66 and not x20 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s123 =>
      if ( x62 and x13 and x4 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( x62 and x13 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x13 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( x62 and not x13 and not x14 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( x62 and not x13 and not x14 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( x62 and not x13 and not x14 and not x9 and not x7 and x8 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( x62 and not x13 and not x14 and not x9 and not x7 and not x8 ) = '1' then
         current_otherm <= s123;

      elsif ( not x62 and x63 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x15 and x13 and x4 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s97;

      elsif ( not x62 and x63 and not x15 and x13 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and x63 and not x15 and not x13 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x63 and not x15 and not x13 and not x14 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x63 and not x15 and not x13 and not x14 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x63 and not x15 and not x13 and not x14 and not x9 and not x7 and x8 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x63 and not x15 and not x13 and not x14 and not x9 and not x7 and not x8 ) = '1' then
         current_otherm <= s123;

      elsif ( not x62 and not x63 and x65 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x65 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x65 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x65 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x65 and not x66 ) = '1' then
         y4 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s417;

      elsif ( not x62 and not x63 and not x65 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x65 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and not x65 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s124 =>
      if ( x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s194;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s1;

      end if;

   when s125 =>
      if ( x64 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s418;

      elsif ( not x64 and x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s19;

      elsif ( not x64 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x64 and not x3 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( not x64 and not x3 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( not x64 and not x3 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      else
         y6 <= '1' ;
         current_otherm <= s39;

      end if;

   when s126 =>
      if ( x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( x17 and x18 and not x1 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x17 and x18 and not x1 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x17 and not x18 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s126;

      elsif ( x17 and not x18 and not x2 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s318;

      else
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      end if;

   when s127 =>
      if ( x62 and x65 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x65 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x65 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x65 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x65 and x17 and x11 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( x62 and not x65 and x17 and x11 and not x8 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x62 and not x65 and x17 and not x11 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( x62 and not x65 and not x17 and x18 and x8 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s318;

      elsif ( x62 and not x65 and not x17 and x18 and not x8 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s105;

      elsif ( x62 and not x65 and not x17 and not x18 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x63 and x2 and x3 and x11 ) = '1' then
         y13 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s270;

      elsif ( not x62 and x63 and x2 and x3 and not x11 ) = '1' then
         y13 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s419;

      elsif ( not x62 and x63 and x2 and not x3 and x4 and x11 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s272;

      elsif ( not x62 and x63 and x2 and not x3 and x4 and not x11 and x12 and x13 and x14 ) = '1' then
         y3 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s420;

      elsif ( not x62 and x63 and x2 and not x3 and x4 and not x11 and x12 and x13 and not x14 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s421;

      elsif ( not x62 and x63 and x2 and not x3 and x4 and not x11 and x12 and not x13 ) = '1' then
         y3 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s422;

      elsif ( not x62 and x63 and x2 and not x3 and x4 and not x11 and not x12 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s423;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and x6 and x5 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and x6 and not x5 and x9 and x7 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and x6 and not x5 and x9 and not x7 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and x6 and not x5 and not x9 and x7 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and x6 and not x5 and not x9 and not x7 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and x7 and x5 and x8 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and x7 and x5 and not x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and x7 and not x5 and x10 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and x7 and not x5 and not x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and not x7 and x5 and x8 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and not x7 and x5 and not x8 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and not x7 and not x5 and x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and x63 and x2 and not x3 and not x4 and not x6 and not x7 and not x5 and not x10 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s424;

      elsif ( not x62 and x63 and not x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x62 and not x63 and x64 and x65 and x20 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( not x62 and not x63 and x64 and x65 and x20 and not x3 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s425;

      elsif ( not x62 and not x63 and x64 and x65 and not x20 and x21 and x3 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x62 and not x63 and x64 and x65 and not x20 and x21 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s415;

      elsif ( not x62 and not x63 and x64 and x65 and not x20 and not x21 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( not x62 and not x63 and x64 and x65 and not x20 and not x21 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s427;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and x19 and x12 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and x19 and not x12 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s254;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and x6 ) = '1' then
         y16 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s255;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and x16 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and x12 and not x6 and not x16 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and x6 ) = '1' then
         y12 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s257;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and x15 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and x18 and not x19 and not x12 and not x6 and not x15 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and not x18 and x19 ) = '1' then
         y27 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and not x18 and not x19 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x62 and not x63 and x64 and not x65 and x5 and not x18 and not x19 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and x11 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and not x11 and x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and x12 and not x11 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and x10 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and not x10 and x9 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and x6 and not x12 and not x10 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and not x6 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and x19 and not x6 and not x12 ) = '1' then
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and x14 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and x12 and not x14 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and x13 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and x6 and not x12 and not x13 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and x18 and not x19 and not x6 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and x12 and x6 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s260;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and x12 and not x6 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s261;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and not x12 and x6 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and x19 and not x12 and not x6 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x62 and not x63 and x64 and not x65 and not x5 and not x18 and not x19 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      else
         y37 <= '1' ;
         current_otherm <= s428;

      end if;

   when s128 =>
      if ( x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         y9 <= '1' ;
         current_otherm <= s46;

      end if;

   when s129 =>
      if ( x64 and x63 and x4 and x5 and x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and x63 and x4 and x5 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x64 and x63 and x4 and x5 and not x3 and not x6 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x64 and x63 and x4 and x5 and not x3 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s340;

      elsif ( x64 and x63 and x4 and not x5 and x3 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x64 and x63 and x4 and not x5 and not x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x64 and x63 and x4 and not x5 and not x3 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x64 and x63 and x4 and not x5 and not x3 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and not x4 and x5 and x3 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x64 and x63 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and not x4 and not x5 and x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and not x4 and not x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and not x63 and x66 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s429;

      elsif ( x64 and not x63 and not x66 and x67 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s399;

      elsif ( x64 and not x63 and not x66 and not x67 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s430;

      elsif ( not x64 and x63 and x66 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s431;

      elsif ( not x64 and x63 and not x66 and x67 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s431;

      elsif ( not x64 and x63 and not x66 and not x67 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s432;

      elsif ( not x64 and not x63 and x65 and x67 ) = '1' then
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s433;

      elsif ( not x64 and not x63 and x65 and not x67 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s434;

      elsif ( not x64 and not x63 and not x65 and x66 and x67 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s435;

      elsif ( not x64 and not x63 and not x65 and x66 and not x67 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s432;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s434;

      end if;

   when s130 =>
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s436;

   when s131 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s142;

      end if;

   when s132 =>
         y8 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s437;

   when s133 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s438;

   when s134 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s439;

      end if;

   when s135 =>
      if ( x62 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and x63 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x65 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x65 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s440;

      end if;

   when s136 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s441;

   when s137 =>
      if ( x62 and x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x32 and x33 ) = '1' then
         y8 <= '1' ;
         y36 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s442;

      elsif ( x62 and not x32 and not x33 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and not x32 and not x33 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and not x32 and not x33 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x32 and not x33 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s138 =>
      if ( x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s139 =>
      if ( x33 and x32 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s443;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s443;

      end if;

   when s140 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s141;

      end if;

   when s141 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y12 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s444;

      else
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s144;

      end if;

   when s142 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s140;

      elsif ( not x32 and not x33 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x33 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x33 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s143 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s445;

   when s144 =>
      if ( x33 and x32 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s446;

      elsif ( x33 and not x32 and x30 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s446;

      elsif ( x33 and not x32 and not x30 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x33 and not x32 and not x30 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x33 and not x32 and not x30 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 and not x30 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s446;

      end if;

   when s145 =>
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s447;

   when s146 =>
         y30 <= '1' ;
         current_otherm <= s185;

   when s147 =>
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s448;

   when s148 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s449;

      end if;

   when s149 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s450;

      elsif ( not x62 and x20 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s451;

      elsif ( not x62 and not x20 and x21 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s452;

      else
         y28 <= '1' ;
         current_otherm <= s377;

      end if;

   when s150 =>
      if ( x62 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y48 <= '1' ;
         y57 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s453;

      end if;

   when s151 =>
      if ( x62 and x20 and x18 and x17 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( x62 and x20 and x18 and x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and x20 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and x20 and not x18 and x17 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and x20 and not x18 and not x17 and x19 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and x20 and not x18 and not x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and x22 and x18 and x17 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( x62 and not x20 and x22 and x18 and x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and x22 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and x22 and not x18 and x17 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x20 and x22 and not x18 and not x17 and x19 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x20 and x22 and not x18 and not x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and not x22 and x21 and x18 and x17 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( x62 and not x20 and not x22 and x21 and x18 and x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and not x22 and x21 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and not x22 and x21 and not x18 and x17 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x20 and not x22 and x21 and not x18 and not x17 and x19 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( x62 and not x20 and not x22 and x21 and not x18 and not x17 and not x19 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( x62 and not x20 and not x22 and not x21 and x24 and x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x62 and not x20 and not x22 and not x21 and x24 and x2 and not x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x62 and not x20 and not x22 and not x21 and x24 and not x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x62 and not x20 and not x22 and not x21 and not x24 and x2 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x62 and not x20 and not x22 and not x21 and not x24 and not x2 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x62 and not x20 and not x22 and not x21 and not x24 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s454;

      end if;

   when s152 =>
      if ( x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      else
         y60 <= '1' ;
         current_otherm <= s190;

      end if;

   when s153 =>
      if ( x63 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s455;

      elsif ( not x63 and x65 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s456;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s456;

      end if;

   when s154 =>
      if ( x63 and x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( x63 and not x19 and x4 and x22 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s153;

      elsif ( x63 and not x19 and x4 and not x22 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      elsif ( x63 and not x19 and not x4 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x63 and not x19 and not x4 and not x18 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      elsif ( not x63 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s155 =>
      if ( x63 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s156 =>
      if ( x63 ) = '1' then
         y23 <= '1' ;
         y65 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s457;

      elsif ( not x63 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s157 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s458;

   when s158 =>
      if ( x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and x65 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x14 and x65 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x14 and x65 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and not x65 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and x14 and not x65 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and x14 and not x65 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s159 =>
         y24 <= '1' ;
         current_otherm <= s406;

   when s160 =>
         y21 <= '1' ;
         current_otherm <= s459;

   when s161 =>
      if ( x67 and x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x67 and not x11 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( x67 and not x11 and not x4 ) = '1' then
         current_otherm <= s161;

      elsif ( not x67 and x10 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( not x67 and x10 and not x4 ) = '1' then
         current_otherm <= s161;

      elsif ( not x67 and not x10 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x67 and not x10 and not x15 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      else
         current_otherm <= s161;

      end if;

   when s162 =>
      if ( x63 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x65 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x63 and not x65 and x66 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s460;

      else
         y9 <= '1' ;
         current_otherm <= s43;

      end if;

   when s163 =>
      if ( x12 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x12 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      else
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s164;

      end if;

   when s164 =>
      if ( x10 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x10 and x11 ) = '1' then
         y14 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s163;

      else
         y10 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s164;

      end if;

   when s165 =>
      if ( x62 and x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x62 and not x12 ) = '1' then
         current_otherm <= s165;

      elsif ( not x62 and x63 and x15 ) = '1' then
         y11 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s461;

      elsif ( not x62 and x63 and not x15 and x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x63 and not x15 and not x12 ) = '1' then
         current_otherm <= s165;

      elsif ( not x62 and not x63 and x64 and x20 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and x64 and x20 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and x64 and x20 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x20 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x20 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         current_otherm <= s208;

      end if;

   when s166 =>
      if ( x62 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x65 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and x9 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and x9 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and x9 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and x9 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and x9 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and not x9 and x10 ) = '1' then
         y33 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and x8 and not x9 and not x10 ) = '1' then
         y37 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and x5 and x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and x5 and not x10 and x4 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and x5 and not x10 and not x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and not x5 and x4 and x10 and x6 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and not x5 and x4 and x10 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and not x5 and x4 and not x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and x9 and not x5 and not x4 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y51 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s250;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and x19 and not x8 and not x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y52 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s250;

      elsif ( not x62 and x63 and not x65 and x23 and x22 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s462;

      elsif ( not x62 and x63 and not x65 and x23 and not x22 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and not x22 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and not x22 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x23 and not x22 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and not x65 and x23 and not x22 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and not x23 and x19 and x20 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s251;

      elsif ( not x62 and x63 and not x65 and not x23 and x19 and not x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x62 and x63 and not x65 and not x23 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s462;

      elsif ( not x62 and not x63 and x64 and x65 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and x64 and x65 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and x64 and x65 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x18 ) = '1' then
         y59 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s112;

      elsif ( not x62 and not x63 and x64 and not x65 and not x18 and x19 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and not x63 and x64 and not x65 and not x18 and not x19 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and x67 and x24 and x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and x24 and not x23 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and x67 and not x24 and x11 and x12 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x67 and not x24 and x11 and x12 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and not x64 and x67 and not x24 and x11 and not x12 and x13 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and not x64 and x67 and not x24 and x11 and not x12 and x13 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and not x64 and x67 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x67 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x67 and x29 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x67 and x29 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x67 and x29 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x67 and x29 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y8 <= '1' ;
         current_otherm <= s464;

      end if;

   when s167 =>
      if ( x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x64 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x64 and not x8 and x10 and x9 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s465;

      elsif ( not x64 and not x8 and x10 and not x9 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s23;

      elsif ( not x64 and not x8 and not x10 and x9 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      else
         y23 <= '1' ;
         current_otherm <= s320;

      end if;

   when s168 =>
      if ( x62 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x23 and x22 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and x23 and x22 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and x23 and x22 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x23 and x22 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and x63 and x23 and x22 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x23 and not x22 and x19 and x20 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s251;

      elsif ( not x62 and x63 and x23 and not x22 and x19 and not x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x62 and x63 and x23 and not x22 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s462;

      elsif ( not x62 and x63 and not x23 ) = '1' then
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s158;

      elsif ( not x62 and not x63 and x64 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and x24 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and not x24 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and not x24 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x67 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x67 and x29 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x65 and not x67 and x29 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x65 and not x67 and x29 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x67 and x29 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and not x67 and not x29 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s466;

      elsif ( not x62 and not x63 and not x64 and not x65 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x65 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x65 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s169 =>
      if ( x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and x63 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x65 and x64 and x63 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x65 and x64 and x63 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and x63 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and not x63 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x65 and x64 and not x63 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x65 and x64 and not x63 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and x64 and not x63 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and x63 and x66 and x30 and x8 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x62 and x65 and not x64 and x63 and x66 and x30 and not x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and x65 and not x64 and x63 and x66 and not x30 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s3;

      elsif ( not x62 and x65 and not x64 and x63 and not x66 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and x23 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and x23 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and x23 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and x23 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and not x23 and x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and not x23 and not x24 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and not x23 and not x24 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and not x23 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and x66 and not x23 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and not x66 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and x65 and not x64 and not x63 and not x66 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and x65 and not x64 and not x63 and not x66 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x64 and not x63 and not x66 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and not x65 and x64 and x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and not x65 and x64 and x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and not x63 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x65 and x64 and not x63 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x65 and x64 and not x63 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and not x63 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and x67 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and x67 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and x67 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and x67 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and not x67 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and not x67 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and not x67 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and x64 and not x63 and not x66 and not x67 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x65 and not x64 and x63 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      else
         current_otherm <= s1;

      end if;

   when s170 =>
      if ( x63 and x20 and x21 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s467;

      elsif ( x63 and x20 and not x21 ) = '1' then
         y6 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s468;

      elsif ( x63 and not x20 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s469;

      elsif ( not x63 and x67 and x23 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s470;

      elsif ( not x63 and x67 and not x23 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and x67 and not x23 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and x67 and not x23 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x67 and not x23 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x67 and x29 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x67 and x29 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x67 and x29 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x67 and x29 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y8 <= '1' ;
         current_otherm <= s464;

      end if;

   when s171 =>
      if ( x62 and x20 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x20 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x20 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x20 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x20 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x63 and x65 and x64 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x65 and x64 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x65 and x64 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x65 and x64 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x65 and not x64 and x66 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x63 and x65 and not x64 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and x65 and not x64 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and x65 and not x64 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and x63 and x65 and not x64 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and x65 and not x64 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and x65 and not x64 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x64 and x17 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x62 and x63 and not x65 and x64 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x63 and not x65 and x64 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x63 and not x65 and x64 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and x64 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x65 and not x64 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x62 and x63 and not x65 and not x64 and not x2 and x5 and x3 and x1 ) = '1' then
         current_otherm <= s171;

      elsif ( not x62 and x63 and not x65 and not x64 and not x2 and x5 and x3 and not x1 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and x63 and not x65 and not x64 and not x2 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x62 and x63 and not x65 and not x64 and not x2 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( not x62 and not x63 and x66 and x65 and x23 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and x66 and x65 and x23 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x63 and x66 and x65 and x23 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x66 and x65 and x23 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and x24 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and x24 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and x24 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and x24 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and not x24 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and not x24 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x66 and x65 and not x23 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x66 and not x65 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      else
         current_otherm <= s1;

      end if;

   when s172 =>
      if ( x63 and x64 ) = '1' then
         y2 <= '1' ;
         y17 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s472;

      elsif ( x63 and not x64 ) = '1' then
         y66 <= '1' ;
         current_otherm <= s473;

      elsif ( not x63 and x23 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and x23 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and x23 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x23 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x23 and x24 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x23 and x24 and not x12 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x23 and x24 and not x12 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x23 and x24 and not x12 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x23 and x24 and not x12 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x23 and not x24 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x23 and not x24 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x23 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s173 =>
      if ( x64 and x63 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s474;

      elsif ( x64 and not x63 and x65 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and not x63 and x65 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and not x63 and x65 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and x65 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and x65 and not x66 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and x66 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and x10 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and x12 and x13 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s475;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and x12 and not x13 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and x12 and not x13 and x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and x12 and not x13 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and not x12 and x14 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s476;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and not x12 and not x14 and x18 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and not x12 and not x14 and x18 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and x11 and not x10 and not x12 and not x14 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and not x11 and x12 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and not x11 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s408;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and not x11 and not x12 and x10 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and x6 and not x11 and not x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y38 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s408;

      elsif ( x64 and not x63 and not x65 and not x66 and x8 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s477;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s477;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and x11 and x12 and x10 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and x11 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s479;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and x11 and not x12 and x10 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and x11 and not x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s408;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and not x11 and x12 and x10 ) = '1' then
         y42 <= '1' ;
         current_otherm <= s354;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and not x11 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and not x11 and not x12 and x10 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and x6 and not x11 and not x12 and not x10 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( x64 and not x63 and not x65 and not x66 and not x8 and not x7 and not x6 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s480;

      elsif ( not x64 and x63 and x11 and x4 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s172;

      elsif ( not x64 and x63 and x11 and not x4 ) = '1' then
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s481;

      elsif ( not x64 and x63 and not x11 and x4 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x64 and x63 and not x11 and not x4 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x64 and x63 and not x11 and not x4 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x63 and x67 and x23 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( not x64 and not x63 and x67 and not x23 and x24 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x67 and not x23 and x24 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x64 and not x63 and x67 and not x23 and x24 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x67 and not x23 and x24 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x67 and not x23 and not x24 and x11 and x12 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x64 and not x63 and x67 and not x23 and not x24 and x11 and not x12 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x64 and not x63 and x67 and not x23 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x67 and not x23 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and not x67 and x29 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x63 and not x67 and x29 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x63 and not x67 and x29 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and not x67 and x29 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y8 <= '1' ;
         current_otherm <= s466;

      end if;

   when s174 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y40 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s482;

   when s175 =>
      if ( x62 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x20 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and x63 and not x20 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x20 and not x18 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      elsif ( not x62 and not x63 and x64 and x65 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and not x63 and x64 and x65 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and not x63 and x64 and x65 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         y38 <= '1' ;
         current_otherm <= s483;

      end if;

   when s176 =>
      if ( x62 and x66 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s484;

      elsif ( x62 and not x66 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x62 and not x66 and not x11 and x10 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s271;

      elsif ( x62 and not x66 and not x11 and not x10 ) = '1' then
         current_otherm <= s176;

      elsif ( not x62 and x63 and x66 and x31 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and x66 and x31 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and x66 and not x31 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and x66 and not x31 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x66 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x66 and not x15 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and x63 and not x66 and not x15 and not x11 and x10 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s271;

      elsif ( not x62 and x63 and not x66 and not x15 and not x11 and not x10 ) = '1' then
         current_otherm <= s176;

      elsif ( not x62 and not x63 and x64 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x62 and not x63 and not x64 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s177 =>
         y14 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s485;

   when s178 =>
      if ( x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x64 and x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x64 and x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and x67 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x67 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x64 and not x63 and x65 and not x67 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x64 and not x63 and x65 and not x67 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 and not x67 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x65 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x65 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and not x64 and x63 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and not x63 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x64 and not x63 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x62 and not x64 and not x63 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s179 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x64 and x66 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x64 and x66 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x66 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and not x66 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and not x66 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x66 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and x24 and x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and x24 and not x23 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x67 and x24 and not x23 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x67 and x24 and not x23 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and x24 and not x23 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and not x24 and x11 and x12 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and not x64 and x67 and not x24 and x11 and x12 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x67 and not x24 and x11 and not x12 and x13 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and not x64 and x67 and not x24 and x11 and not x12 and x13 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x67 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x67 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x67 and x28 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and not x67 and x28 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and not x67 and x28 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x67 and x28 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y8 <= '1' ;
         current_otherm <= s356;

      end if;

   when s180 =>
      if ( x21 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x21 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x21 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x21 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x21 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s181 =>
      if ( x63 and x66 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x66 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x66 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x66 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x66 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and x66 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x65 and x66 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x65 and x66 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and x66 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x66 and x6 and x7 and x67 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x63 and x64 and x65 and not x66 and x6 and x7 and not x67 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x65 and not x66 and x6 and not x7 and x8 and x67 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x63 and x64 and x65 and not x66 and x6 and not x7 and x8 and not x67 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x65 and not x66 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x66 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and x67 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x64 and not x65 and x67 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x64 and not x65 and x67 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and x67 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and x67 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and not x67 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and not x67 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and not x67 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and not x67 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x31 and x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x63 and not x64 and x31 and not x30 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s486;

      elsif ( not x63 and not x64 and not x31 and x30 ) = '1' then
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s487;

      else
         y25 <= '1' ;
         current_otherm <= s363;

      end if;

   when s182 =>
      if ( x63 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s488;

      elsif ( not x63 and x65 and x21 and x17 and x16 and x19 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x65 and x21 and x17 and x16 and x19 and not x11 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x21 and x17 and x16 and not x19 and x18 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x65 and x21 and x17 and x16 and not x19 and not x18 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x21 and x17 and not x16 and x11 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( not x63 and x65 and x21 and x17 and not x16 and not x11 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s365;

      elsif ( not x63 and x65 and x21 and not x17 and x16 and x19 and x14 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x65 and x21 and not x17 and x16 and x19 and not x14 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x21 and not x17 and x16 and not x19 and x13 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x65 and x21 and not x17 and x16 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x21 and not x17 and not x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and not x21 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s185;

      else
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s489;

      end if;

   when s183 =>
      if ( x64 and x17 and x16 and x19 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and x17 and x16 and x19 and not x11 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and x17 and x16 and not x19 and x18 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and x17 and x16 and not x19 and not x18 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and x17 and not x16 and x11 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( x64 and x17 and not x16 and not x11 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s365;

      elsif ( x64 and not x17 and x16 and x19 and x14 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and not x17 and x16 and x19 and not x14 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and not x17 and x16 and not x19 and x13 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and not x17 and x16 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and not x17 and not x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( not x64 and not x30 and x4 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      else
         y5 <= '1' ;
         current_otherm <= s359;

      end if;

   when s184 =>
      if ( x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s185 =>
      if ( x62 ) = '1' then
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s490;

      elsif ( not x62 and x64 ) = '1' then
         current_otherm <= s65;

      else
         y35 <= '1' ;
         current_otherm <= s269;

      end if;

   when s186 =>
      if ( x63 ) = '1' then
         y60 <= '1' ;
         current_otherm <= s190;

      else
         current_otherm <= s1;

      end if;

   when s187 =>
      if ( x23 and x17 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s491;

      elsif ( x23 and x17 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s492;

      elsif ( x23 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s493;

      elsif ( not x23 and x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s492;

      elsif ( not x23 and x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s493;

      elsif ( not x23 and not x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s491;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s494;

      end if;

   when s188 =>
      if ( x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s491;

      elsif ( x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s495;

      elsif ( not x22 and x23 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s491;

      elsif ( not x22 and x23 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s496;

      elsif ( not x22 and not x23 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s497;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s493;

      end if;

   when s189 =>
      if ( x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x24 and x23 and x10 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s23;

      elsif ( not x24 and x23 and not x10 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s320;

      else
         current_otherm <= s1;

      end if;

   when s190 =>
      if ( x63 and x65 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x63 and not x65 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x65 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         y61 <= '1' ;
         current_otherm <= s498;

      end if;

   when s191 =>
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s499;

   when s192 =>
      if ( x64 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s500;

      elsif ( not x64 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x64 and x1 and not x2 and x5 and x3 ) = '1' then
         current_otherm <= s192;

      elsif ( not x64 and x1 and not x2 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      elsif ( not x64 and x1 and not x2 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      else
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      end if;

   when s193 =>
         y6 <= '1' ;
         current_otherm <= s39;

   when s194 =>
      if ( x2 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s352;

      elsif ( not x2 and x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s318;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s1;

      end if;

   when s195 =>
      if ( x3 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( x3 and x1 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s307;

      elsif ( x3 and not x1 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s1;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      end if;

   when s196 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

   when s197 =>
      if ( x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s2;

      elsif ( not x5 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s196;

      elsif ( not x5 and x2 and not x1 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s197;

      elsif ( not x5 and not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s198;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s2;

      end if;

   when s198 =>
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s66;

   when s199 =>
      if ( x62 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s41;

      elsif ( not x62 and x30 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s321;

      elsif ( not x62 and not x30 and x31 ) = '1' then
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s501;

      else
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      end if;

   when s200 =>
      if ( x19 and x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s502;

      elsif ( x19 and not x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s503;

      else
         y2 <= '1' ;
         current_otherm <= s504;

      end if;

   when s201 =>
      if ( x62 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and x63 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s505;

      elsif ( not x62 and not x63 and x64 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s123;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s506;

      end if;

   when s202 =>
         y2 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s507;

   when s203 =>
      if ( x63 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x63 and x64 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x63 and not x64 and x30 and x14 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s509;

      elsif ( not x63 and not x64 and x30 and not x14 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s510;

      elsif ( not x63 and not x64 and not x30 and x31 and x14 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x63 and not x64 and not x30 and x31 and not x14 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s511;

      elsif ( not x63 and not x64 and not x30 and not x31 and x14 ) = '1' then
         y45 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         y49 <= '1' ;
         y55 <= '1' ;
         y58 <= '1' ;
         y63 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s512;

      else
         y37 <= '1' ;
         current_otherm <= s181;

      end if;

   when s204 =>
      if ( x64 and x62 and x17 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s513;

      elsif ( x64 and x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s330;

      elsif ( x64 and not x62 and x66 and x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and not x62 and x66 and x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and not x62 and x66 and x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x66 and x21 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x66 and not x21 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x64 and not x62 and not x66 and x67 and x11 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x62 and not x66 and x67 and x11 and not x4 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( x64 and not x62 and not x66 and x67 and not x11 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and not x62 and not x66 and not x67 and x10 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and not x62 and not x66 and not x67 and not x10 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x64 and not x62 and not x66 and not x67 and not x10 and not x4 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( not x64 and x62 and x17 and x18 and x5 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x64 and x62 and x17 and x18 and not x5 and x6 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x64 and x62 and x17 and x18 and not x5 and not x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x64 and x62 and x17 and not x18 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x62 and x17 and not x18 and not x2 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s104;

      elsif ( not x64 and x62 and not x17 and x9 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x64 and x62 and not x17 and not x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and x12 and x10 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and x12 and not x10 and x11 and x13 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and x12 and not x10 and x11 and not x13 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and x12 and not x10 and x11 and not x13 and x19 and not x14 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and x12 and not x10 and x11 and not x13 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and x12 and not x10 and not x11 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y32 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s453;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and not x12 and x10 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s413;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and not x12 and not x10 and x11 and x14 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and not x12 and not x10 and x11 and not x14 and x19 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and not x12 and not x10 and x11 and not x14 and x19 and not x13 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and not x12 and not x10 and x11 and not x14 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and x6 and not x12 and not x10 and not x11 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s514;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and not x6 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s515;

      elsif ( not x64 and not x62 and x3 and x4 and x7 and not x6 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s516;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and x9 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s515;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and x11 and x12 and x6 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and x11 and x12 and not x6 ) = '1' then
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and x11 and not x12 and x6 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and x11 and not x12 and not x6 ) = '1' then
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and not x11 and x6 and x12 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and not x11 and x6 and not x12 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and x10 and not x11 and not x6 ) = '1' then
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and x11 and x12 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s517;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and x11 and x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s518;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and x11 and not x12 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y31 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and x11 and not x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y63 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s519;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and not x11 and x12 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and not x11 and x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s520;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and not x11 and not x12 and x6 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s521;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and x5 and not x9 and not x10 and not x11 and not x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s332;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and not x5 and x8 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and not x5 and x8 and not x6 and x11 and x12 ) = '1' then
         y4 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and not x5 and x8 and not x6 and x11 and not x12 ) = '1' then
         y4 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and not x5 and x8 and not x6 and not x11 ) = '1' then
         y4 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x3 and x4 and not x7 and not x5 and not x8 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s516;

      elsif ( not x64 and not x62 and x3 and not x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s522;

      else
         y5 <= '1' ;
         current_otherm <= s68;

      end if;

   when s205 =>
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1;

   when s206 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s523;

   when s207 =>
      if ( x10 ) = '1' then
         y62 <= '1' ;
         current_otherm <= s524;

      elsif ( not x10 and x11 and x4 and x5 and x3 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x10 and x11 and x4 and x5 and x3 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x10 and x11 and x4 and x5 and x3 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x4 and x5 and x3 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and x6 and not x7 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and x6 and not x7 and x12 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and x6 and not x7 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and not x6 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and not x6 and not x8 and x12 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and not x6 and not x8 and x12 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x4 and x5 and not x3 and not x6 and not x8 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x4 and not x5 and x6 and x3 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x10 and x11 and x4 and not x5 and x6 and not x3 ) = '1' then
         y21 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s180;

      elsif ( not x10 and x11 and x4 and not x5 and not x6 and x3 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x10 and x11 and x4 and not x5 and not x6 and not x3 ) = '1' then
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s180;

      elsif ( not x10 and x11 and not x4 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      else
         y62 <= '1' ;
         current_otherm <= s525;

      end if;

   when s208 =>
      if ( x63 and x64 ) = '1' then
         y21 <= '1' ;
         y27 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s526;

      elsif ( x63 and not x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      else
         y47 <= '1' ;
         y51 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s527;

      end if;

   when s209 =>
      if ( x63 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s528;

      elsif ( not x63 and x31 and x30 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x63 and x31 and not x30 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s386;

      else
         y35 <= '1' ;
         current_otherm <= s386;

      end if;

   when s210 =>
      if ( x19 and x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s351;

      elsif ( x19 and not x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s529;

      else
         y2 <= '1' ;
         current_otherm <= s502;

      end if;

   when s211 =>
      if ( x62 and x5 and x2 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( x62 and x5 and not x2 and x4 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( x62 and x5 and not x2 and x4 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( x62 and x5 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( x62 and not x5 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( not x62 and x16 and x15 and x5 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x16 and x15 and not x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      elsif ( not x62 and x16 and not x15 and x2 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( not x62 and x16 and not x15 and not x2 and x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and x16 and not x15 and not x2 and x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x16 and not x15 and not x2 and x4 and not x5 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( not x62 and x16 and not x15 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      elsif ( not x62 and not x16 and x15 and x13 and x11 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and not x16 and x15 and x13 and not x11 and x6 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and not x16 and x15 and x13 and not x11 and x6 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and not x16 and x15 and x13 and not x11 and not x6 and x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and not x16 and x15 and x13 and not x11 and not x6 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x62 and not x16 and x15 and not x13 and x14 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and not x16 and x15 and not x13 and not x14 and x9 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and not x16 and x15 and not x13 and not x14 and not x9 and x6 and x2 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and not x16 and x15 and not x13 and not x14 and not x9 and x6 and not x2 ) = '1' then
         current_otherm <= s211;

      elsif ( not x62 and not x16 and x15 and not x13 and not x14 and not x9 and not x6 and x8 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and not x16 and x15 and not x13 and not x14 and not x9 and not x6 and not x8 ) = '1' then
         current_otherm <= s211;

      else
         current_otherm <= s1;

      end if;

   when s212 =>
      if ( x62 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( x62 and not x2 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( x62 and not x2 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and x16 and x15 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s530;

      elsif ( not x62 and x16 and not x15 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x62 and x16 and not x15 and not x2 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and x16 and not x15 and not x2 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      else
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s530;

      end if;

   when s213 =>
      if ( x62 and x4 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( x62 and not x4 and not x2 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( x62 and not x4 and not x2 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and x16 and x15 and x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and x16 and x15 and not x5 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and x16 and not x15 and x4 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x16 and not x15 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x16 and not x15 and not x4 and not x2 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and x16 and not x15 and not x4 and not x2 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and not x16 and x15 and x12 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and not x16 and x15 and not x12 ) = '1' then
         current_otherm <= s213;

      else
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      end if;

   when s214 =>
      if ( x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( x4 and not x5 and x2 and x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      elsif ( x4 and not x5 and x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( x4 and not x5 and not x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x4 and x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x4 and x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      else
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      end if;

   when s215 =>
      if ( x62 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s349;

      elsif ( x62 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s221;

      elsif ( not x62 and x15 and x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and not x16 and x13 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and x15 and not x16 and x13 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and x15 and not x16 and not x13 and x14 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x15 and not x16 and not x13 and not x14 and x9 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x15 and not x16 and not x13 and not x14 and not x9 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x15 and not x16 and not x13 and not x14 and not x9 and not x7 and x8 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x15 and not x16 and not x13 and not x14 and not x9 and not x7 and not x8 ) = '1' then
         current_otherm <= s215;

      elsif ( not x62 and not x15 and x16 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s349;

      elsif ( not x62 and not x15 and x16 and not x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      else
         current_otherm <= s1;

      end if;

   when s216 =>
      if ( x62 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( not x62 and x15 and x16 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x15 and x16 and x5 and not x1 and x2 and x3 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and x15 and x16 and x5 and not x1 and x2 and x3 and not x4 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and x16 and x5 and not x1 and x2 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and x16 and x5 and not x1 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and x16 and not x5 and x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and x16 and not x5 and not x6 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and x15 and x16 and not x5 and not x6 and not x1 and x2 and x3 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and x15 and x16 and not x5 and not x6 and not x1 and x2 and x3 and not x4 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and x15 and x16 and not x5 and not x6 and not x1 and x2 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and x16 and not x5 and not x6 and not x1 and not x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x15 and not x16 and x6 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and x15 and not x16 and not x6 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and not x15 and x16 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      else
         current_otherm <= s1;

      end if;

   when s217 =>
      if ( x62 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and x16 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and not x16 and x15 and x8 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x62 and not x16 and x15 and not x8 and x9 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x62 and not x16 and x15 and not x8 and not x9 and x10 and x6 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      elsif ( not x62 and not x16 and x15 and not x8 and not x9 and x10 and not x6 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and not x16 and x15 and not x8 and not x9 and not x10 and x11 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and not x16 and x15 and not x8 and not x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s217;

      else
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s82;

      end if;

   when s218 =>
      if ( x15 and x16 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and x16 and x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x15 and x16 and x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x15 and x16 and x4 and not x5 and x2 and x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      elsif ( not x15 and x16 and x4 and not x5 and x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x15 and x16 and x4 and not x5 and not x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( not x15 and x16 and not x4 and x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x15 and x16 and not x4 and x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s216;

      elsif ( not x15 and x16 and not x4 and not x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      end if;

   when s219 =>
      if ( x62 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and x16 and x15 and x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x62 and x16 and x15 and not x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      elsif ( not x62 and x16 and not x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and not x16 and x15 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      elsif ( not x62 and not x16 and x15 and not x12 ) = '1' then
         current_otherm <= s219;

      elsif ( not x62 and not x16 and not x15 and x13 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      else
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s215;

      end if;

   when s220 =>
      if ( x62 and x1 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( x62 and not x1 and x4 and x5 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( x62 and not x1 and x4 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( x62 and not x1 and not x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x62 and x15 and x16 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and x15 and not x16 and x3 and x2 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and x15 and not x16 and x3 and not x2 ) = '1' then
         current_otherm <= s220;

      elsif ( not x62 and x15 and not x16 and not x3 and x4 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and x15 and not x16 and not x3 and x4 and not x2 ) = '1' then
         current_otherm <= s220;

      elsif ( not x62 and x15 and not x16 and not x3 and not x4 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      elsif ( not x62 and x15 and not x16 and not x3 and not x4 and not x2 ) = '1' then
         current_otherm <= s220;

      elsif ( not x62 and not x15 and x1 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and not x15 and not x1 and x16 and x4 and x5 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      elsif ( not x62 and not x15 and not x1 and x16 and x4 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and not x15 and not x1 and x16 and not x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      else
         y4 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s217;

      end if;

   when s221 =>
      if ( x4 and x5 and x1 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s220;

      elsif ( x4 and x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( x4 and not x5 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( x4 and not x5 and not x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x4 and x1 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      else
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      end if;

   when s222 =>
         y6 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1;

   when s223 =>
      if ( x17 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s531;

      else
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s223;

      end if;

   when s224 =>
      if ( x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and x10 ) = '1' then
         y62 <= '1' ;
         current_otherm <= s524;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and x3 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and x3 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and x3 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and x3 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and x6 and not x7 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and x6 and not x7 and x12 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and x6 and not x7 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and not x6 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and not x6 and not x8 and x12 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and not x6 and not x8 and x12 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and x5 and not x3 and not x6 and not x8 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and not x5 and x6 and x3 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and not x5 and x6 and not x3 ) = '1' then
         y21 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s180;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and not x5 and not x6 and x3 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x63 and x64 and x11 and not x10 and x4 and not x5 and not x6 and not x3 ) = '1' then
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s180;

      elsif ( not x63 and x64 and x11 and not x10 and not x4 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x64 and not x11 ) = '1' then
         y62 <= '1' ;
         current_otherm <= s525;

      elsif ( not x63 and not x64 and x16 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and not x16 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x16 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x16 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s225 =>
      if ( x62 and x17 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s532;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s533;

      elsif ( not x62 and x64 and x63 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x64 and x63 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x64 and x63 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x13 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s534;

      elsif ( not x62 and x64 and not x63 and not x13 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and not x13 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and x64 and not x63 and not x13 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x13 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x65 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and not x64 and x63 and x65 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and not x64 and x63 and x65 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and not x64 and x63 and x65 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and not x64 and x63 and x65 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and not x64 and x63 and x65 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and not x65 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and not x63 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and not x63 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s226 =>
      if ( x63 and x7 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      elsif ( x63 and not x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      else
         current_otherm <= s1;

      end if;

   when s227 =>
      if ( x62 and x10 and x7 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and x10 and not x7 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( x62 and not x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x13 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and not x13 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and x7 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      else
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      end if;

   when s228 =>
      if ( x62 and x13 and x8 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and x13 and x8 and not x1 and x14 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( x62 and x13 and x8 and not x1 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and x13 and not x8 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( x62 and not x13 and x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and not x10 and x6 and x7 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( x62 and not x13 and not x10 and x6 and x7 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and not x13 and not x10 and x6 and x7 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x10 and x6 and x7 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and not x13 and not x10 and x6 and not x7 and x8 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( x62 and not x13 and not x10 and x6 and not x7 and not x8 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( x62 and not x13 and not x10 and x6 and not x7 and not x8 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( x62 and not x13 and not x10 and x6 and not x7 and not x8 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( x62 and not x13 and not x10 and x6 and not x7 and not x8 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and not x13 and not x10 and not x6 and x16 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( x62 and not x13 and not x10 and not x6 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x17 and x18 and x5 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and x17 and x18 and not x5 and x6 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and x18 and not x5 and not x6 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and not x18 and x9 and x10 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and x17 and not x18 and x9 and not x10 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and not x18 and not x9 and x6 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and x17 and not x18 and not x9 and not x6 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and not x17 and x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and not x18 and x6 and x7 and x2 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x18 and x6 and x7 and x2 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and not x17 and not x18 and x6 and x7 and x2 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and not x17 and not x18 and x6 and x7 and not x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and not x17 and not x18 and x6 and not x7 and x8 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and not x17 and not x18 and x6 and not x7 and not x8 and x2 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and not x18 and x6 and not x7 and not x8 and x2 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and not x17 and not x18 and x6 and not x7 and not x8 and x2 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and not x17 and not x18 and x6 and not x7 and not x8 and not x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and not x17 and not x18 and not x6 and x2 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      else
         current_otherm <= s1;

      end if;

   when s229 =>
      if ( x62 and x13 and x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x13 and not x20 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( x62 and not x13 and x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and not x12 and x10 and x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( x62 and not x13 and not x12 and x10 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( x62 and not x13 and not x12 and not x10 and x19 and x16 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( x62 and not x13 and not x12 and not x10 and x19 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x13 and not x12 and not x10 and not x19 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( not x62 and x18 and x17 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x18 and x17 and not x1 and x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x18 and x17 and not x1 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x18 and not x17 and x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and x18 and not x17 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( not x62 and not x18 and x17 and x7 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      elsif ( not x62 and not x18 and x17 and not x7 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x18 and not x17 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x18 and not x17 and not x15 and x1 and x2 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and not x18 and not x17 and not x15 and x1 and not x2 ) = '1' then
         current_otherm <= s1;

      else
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s231;

      end if;

   when s230 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x18 and not x1 and x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 and not x1 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x17 and not x18 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      elsif ( not x62 and x17 and not x18 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s234;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      end if;

   when s231 =>
      if ( x62 and x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( x62 and not x13 and x10 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s234;

      elsif ( x62 and not x13 and x10 and not x5 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      elsif ( x62 and not x13 and not x10 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      elsif ( not x62 and x17 and x11 and x8 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and x17 and x11 and not x8 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and not x17 and x18 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s234;

      elsif ( not x62 and not x17 and x18 and not x8 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      else
         y11 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s229;

      end if;

   when s232 =>
      if ( x62 and x9 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and not x9 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      elsif ( not x62 and x17 and x18 and x5 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and x17 and x18 and not x5 and x6 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and x18 and not x5 and not x6 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and not x18 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x17 and not x18 and not x2 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s233;

      elsif ( not x62 and not x17 and x9 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      else
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s228;

      end if;

   when s233 =>
      if ( x62 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      elsif ( x62 and not x6 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      elsif ( not x62 and x17 and x18 and x5 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and x17 and x18 and not x5 and x6 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and x18 and not x5 and not x6 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and not x18 and x14 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s32;

      elsif ( not x62 and x17 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      end if;

   when s234 =>
      if ( x62 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x18 and not x1 and x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and x18 and not x1 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and x17 and not x18 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      elsif ( not x62 and x17 and not x18 and not x6 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s235;

      else
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      end if;

   when s235 =>
      if ( x62 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( x62 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      elsif ( not x62 and x17 and x18 and x6 and x9 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s227;

      elsif ( not x62 and x17 and x18 and x6 and not x9 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      elsif ( not x62 and x17 and x18 and not x6 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s233;

      elsif ( not x62 and x17 and not x18 and x10 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and not x18 and not x10 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s232;

      elsif ( not x62 and not x17 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s34;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s230;

      end if;

   when s236 =>
         y2 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s84;

   when s237 =>
      if ( x64 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( x64 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s537;

      else
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s538;

      end if;

   when s238 =>
      if ( x62 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s539;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s540;

      elsif ( not x62 and x63 and x64 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x64 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x64 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x64 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x64 and x66 and x7 and x31 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x62 and x63 and not x64 and x66 and x7 and not x31 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and not x64 and x66 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and not x64 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and not x64 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and x63 and not x64 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and x63 and not x64 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and not x64 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and x63 and not x64 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s239 =>
      if ( x63 and x22 and x16 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x22 and x16 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x22 and x16 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x22 and x16 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x22 and x16 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x22 and not x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s541;

      elsif ( x63 and not x22 and x16 and x23 ) = '1' then
         y3 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x22 and x16 and not x23 and x7 and x9 and x10 and x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x22 and x16 and not x23 and x7 and x9 and x10 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x22 and x16 and not x23 and x7 and x9 and not x10 and x8 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( x63 and not x22 and x16 and not x23 and x7 and x9 and not x10 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x22 and x16 and not x23 and x7 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s542;

      elsif ( x63 and not x22 and x16 and not x23 and x7 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x22 and x16 and not x23 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s251;

      elsif ( x63 and not x22 and not x16 and x23 ) = '1' then
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s249;

      elsif ( x63 and not x22 and not x16 and not x23 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s252;

      elsif ( not x63 and x67 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s475;

      elsif ( not x63 and not x67 and x21 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x67 and x21 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x67 and x21 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x67 and x21 and not x6 ) = '1' then
         current_otherm <= s1;

      else
         y7 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s242;

      end if;

   when s240 =>
      if ( x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s241 =>
      if ( x15 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s240;

      elsif ( not x15 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s242 =>
      if ( x9 and x21 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s543;

      elsif ( x9 and not x21 and x22 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s544;

      elsif ( x9 and not x21 and not x22 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s545;

      elsif ( not x9 and x13 and x21 and x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s546;

      elsif ( not x9 and x13 and x21 and not x10 and x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s544;

      elsif ( not x9 and x13 and x21 and not x10 and x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s547;

      elsif ( not x9 and x13 and x21 and not x10 and not x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( not x9 and x13 and x21 and not x10 and not x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s549;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and x11 and x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and x11 and not x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s545;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and x14 and x19 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and not x14 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and x10 and not x22 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s550;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and x14 and x11 and x17 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and x14 and not x11 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x13 and not x21 and not x10 and x22 and not x14 and not x11 ) = '1' then
         y102 <= '1' ;
         current_otherm <= s240;

      elsif ( not x9 and x13 and not x21 and not x10 and not x22 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s551;

      else
         y9 <= '1' ;
         y65 <= '1' ;
         y84 <= '1' ;
         y86 <= '1' ;
         y91 <= '1' ;
         current_otherm <= s552;

      end if;

   when s243 =>
      if ( x12 and x11 and x10 and x13 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x12 and x11 and x10 and x13 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x12 and x11 and x10 and x13 and not x8 and not x1 ) = '1' then
         current_otherm <= s243;

      elsif ( x12 and x11 and x10 and not x13 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( x12 and x11 and not x10 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x12 and x11 and not x10 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x12 and x11 and not x10 and not x8 and not x1 ) = '1' then
         current_otherm <= s243;

      elsif ( x12 and not x11 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x12 and not x11 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x12 and not x11 and not x8 and not x1 ) = '1' then
         current_otherm <= s243;

      elsif ( not x12 and x11 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and x11 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and x11 and not x8 and not x1 ) = '1' then
         current_otherm <= s243;

      elsif ( not x12 and not x11 and x14 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and not x11 and x14 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and not x11 and x14 and not x8 and not x1 ) = '1' then
         current_otherm <= s243;

      elsif ( not x12 and not x11 and not x14 and x13 and x10 and x9 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( not x12 and not x11 and not x14 and x13 and x10 and not x9 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and not x11 and not x14 and x13 and x10 and not x9 and not x7 ) = '1' then
         y15 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s300;

      elsif ( not x12 and not x11 and not x14 and x13 and not x10 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and not x11 and not x14 and x13 and not x10 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and not x11 and not x14 and x13 and not x10 and not x8 and not x1 ) = '1' then
         current_otherm <= s243;

      elsif ( not x12 and not x11 and not x14 and not x13 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x12 and not x11 and not x14 and not x13 and not x8 and x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      else
         current_otherm <= s243;

      end if;

   when s244 =>
      if ( x10 and x13 and x11 and x12 and x3 and x6 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s50;

      elsif ( x10 and x13 and x11 and x12 and x3 and not x6 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and x13 and x11 and x12 and not x3 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and x13 and x11 and not x12 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x10 and x13 and not x11 and x12 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and x13 and not x11 and x12 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x10 and x13 and not x11 and x12 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( x10 and x13 and not x11 and x12 and not x3 and not x1 and not x7 ) = '1' then
         current_otherm <= s244;

      elsif ( x10 and x13 and not x11 and not x12 and x14 and x5 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( x10 and x13 and not x11 and not x12 and x14 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and x13 and not x11 and not x12 and not x14 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( x10 and not x13 and x12 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x10 and not x13 and x12 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x10 and not x13 and x12 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      elsif ( x10 and not x13 and x12 and not x3 and not x1 and not x7 ) = '1' then
         current_otherm <= s244;

      elsif ( x10 and not x13 and not x12 and x14 and x5 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s54;

      elsif ( x10 and not x13 and not x12 and x14 and not x5 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( x10 and not x13 and not x12 and not x14 and x1 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s52;

      elsif ( x10 and not x13 and not x12 and not x14 and not x1 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x13 and not x12 and not x14 and not x1 and not x3 ) = '1' then
         y14 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s51;

      elsif ( not x10 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x10 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x10 and not x3 and not x1 and x7 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      else
         current_otherm <= s244;

      end if;

   when s245 =>
      if ( x62 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      elsif ( not x62 and x5 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s464;

      elsif ( not x62 and not x5 and x21 and x22 and x10 and x14 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x62 and not x5 and x21 and x22 and x10 and not x14 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and x14 and x8 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and x14 and not x8 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and x14 and not x8 and x6 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and x14 and not x8 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and not x14 and x7 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and not x14 and not x7 and x6 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and not x14 and not x7 and x6 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and x11 and not x14 and not x7 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and not x11 and x14 ) = '1' then
         y60 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y67 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and x21 and x22 and not x10 and not x11 and not x14 ) = '1' then
         y58 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and x21 and not x22 and x9 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s551;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and x11 and x14 and x10 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and x11 and x14 and not x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y90 <= '1' ;
         y95 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and x11 and not x14 and x10 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and x11 and not x14 and not x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y93 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and not x11 and x14 and x10 ) = '1' then
         y100 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and not x11 and x14 and not x10 ) = '1' then
         y46 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y73 <= '1' ;
         y95 <= '1' ;
         current_otherm <= s553;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and not x11 and not x14 and x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and x21 and not x22 and not x9 and not x11 and not x14 and not x10 ) = '1' then
         y74 <= '1' ;
         current_otherm <= s554;

      elsif ( not x62 and not x5 and not x21 and x22 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s551;

      elsif ( not x62 and not x5 and not x21 and not x22 and x10 and x11 and x9 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s555;

      elsif ( not x62 and not x5 and not x21 and not x22 and x10 and x11 and not x9 ) = '1' then
         y65 <= '1' ;
         y90 <= '1' ;
         y92 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and not x21 and not x22 and x10 and not x11 and x9 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s551;

      elsif ( not x62 and not x5 and not x21 and not x22 and x10 and not x11 and not x9 ) = '1' then
         y65 <= '1' ;
         y92 <= '1' ;
         y94 <= '1' ;
         y95 <= '1' ;
         current_otherm <= s240;

      elsif ( not x62 and not x5 and not x21 and not x22 and not x10 and x9 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s550;

      else
         y65 <= '1' ;
         y90 <= '1' ;
         y91 <= '1' ;
         y92 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s240;

      end if;

   when s246 =>
      if ( x17 and x13 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x17 and not x13 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x17 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s106;

      else
         y7 <= '1' ;
         current_otherm <= s90;

      end if;

   when s247 =>
      if ( x23 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      else
         y19 <= '1' ;
         current_otherm <= s168;

      end if;

   when s248 =>
         y10 <= '1' ;
         current_otherm <= s16;

   when s249 =>
         y10 <= '1' ;
         current_otherm <= s556;

   when s250 =>
      if ( x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      else
         current_otherm <= s1;

      end if;

   when s251 =>
      if ( x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s557;

      elsif ( not x22 and x8 and x9 and x23 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( not x22 and x8 and x9 and x23 and not x10 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x22 and x8 and x9 and not x23 and x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x8 and x9 and not x23 and not x10 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x22 and x8 and not x9 and x23 and x10 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x8 and not x9 and x23 and x10 and not x13 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x8 and not x9 and x23 and x10 and not x13 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x8 and not x9 and x23 and x10 and not x13 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x8 and not x9 and x23 and x10 and not x13 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x8 and not x9 and x23 and x10 and not x13 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x8 and not x9 and x23 and not x10 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x8 and not x9 and x23 and not x10 and not x1 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x8 and not x9 and x23 and not x10 and not x1 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x8 and not x9 and x23 and not x10 and not x1 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x8 and not x9 and x23 and not x10 and not x1 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x8 and not x9 and x23 and not x10 and not x1 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x8 and not x9 and not x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s542;

      elsif ( not x22 and not x8 and x9 and x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and not x8 and x9 and not x23 and x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and not x8 and x9 and not x23 and not x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and not x8 and not x9 and x23 and x10 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and not x8 and not x9 and x23 and x10 and not x3 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and not x8 and not x9 and x23 and x10 and not x3 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and not x8 and not x9 and x23 and x10 and not x3 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and not x8 and not x9 and x23 and x10 and not x3 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and not x8 and not x9 and x23 and x10 and not x3 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and not x8 and not x9 and x23 and not x10 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and not x8 and not x9 and x23 and not x10 and not x15 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and not x8 and not x9 and x23 and not x10 and not x15 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      end if;

   when s252 =>
      if ( x22 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s558;

      elsif ( not x22 and x23 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s559;

      else
         y10 <= '1' ;
         current_otherm <= s556;

      end if;

   when s253 =>
      if ( x63 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s395;

      elsif ( not x63 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         y52 <= '1' ;
         current_otherm <= s360;

      end if;

   when s254 =>
      if ( x63 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s255 =>
      if ( x13 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s256 =>
      if ( x63 and x65 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s387;

      elsif ( x63 and not x65 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x65 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x67 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x63 and x64 and not x67 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x67 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x67 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x67 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s257 =>
         y46 <= '1' ;
         current_otherm <= s259;

   when s258 =>
      if ( x63 and x9 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x63 and not x9 and x67 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x9 and x67 and not x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( x63 and not x9 and not x67 ) = '1' then
         current_otherm <= s258;

      elsif ( not x63 and x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and x10 and x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and x10 and not x11 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and x13 and x14 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and x13 and not x14 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and x13 and not x14 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and x13 and not x14 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and x13 and not x14 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and not x13 and x15 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and not x13 and not x15 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and not x13 and not x15 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and not x13 and not x15 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and x9 and not x10 and not x13 and not x15 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and x17 and x18 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and x17 and not x18 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and x17 and not x18 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and x17 and not x18 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and x17 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and not x17 and x19 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and not x17 and not x19 and x20 and x21 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and not x17 and not x19 and x20 and not x21 and x22 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and not x17 and not x19 and x20 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and x16 and not x17 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and x24 and not x23 and not x9 and not x16 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x63 and not x64 and x65 and x66 and not x24 and x11 and x12 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and not x64 and x65 and x66 and not x24 and x11 and x12 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x65 and x66 and not x24 and x11 and not x12 and x13 and x23 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and not x64 and x65 and x66 and not x24 and x11 and not x12 and x13 and not x23 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x63 and not x64 and x65 and x66 and not x24 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x66 and not x24 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and not x66 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and not x64 and x65 and not x66 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and not x64 and x65 and not x66 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and not x66 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x65 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x65 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x65 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s259 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s260 =>
      if ( x63 and x18 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x63 and x18 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x63 and x18 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x63 and not x18 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x63 and not x18 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x63 and not x18 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x18 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x65 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x65 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and not x65 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and not x64 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and not x64 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s261 =>
      if ( x64 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x64 and x31 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      else
         y25 <= '1' ;
         current_otherm <= s363;

      end if;

   when s262 =>
      if ( x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x65 and x4 and x5 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and x63 and x65 and x4 and not x5 ) = '1' then
         y69 <= '1' ;
         y73 <= '1' ;
         current_otherm <= s563;

      elsif ( not x62 and x63 and x65 and not x4 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x62 and x63 and not x65 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and x63 and not x65 and not x13 ) = '1' then
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s164;

      elsif ( not x62 and not x63 and x64 and x65 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and x65 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x62 and not x63 and x64 and x65 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x65 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x65 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x66 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x66 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x66 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x66 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s263 =>
      if ( x63 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and x65 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x65 and not x15 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s264 =>
         y3 <= '1' ;
         y28 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s1;

   when s265 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s564;

   when s266 =>
         y2 <= '1' ;
         y6 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s565;

   when s267 =>
         y14 <= '1' ;
         current_otherm <= s94;

   when s268 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s566;

      elsif ( x62 and not x64 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s567;

      elsif ( not x62 and x63 and x13 and x67 and x11 and x14 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x63 and x13 and x67 and x11 and not x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and x10 and x14 and x3 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and x10 and x14 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and x10 and x14 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and x10 and not x14 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and x10 and not x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and not x10 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s78;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and not x10 and not x1 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x13 and x67 and not x11 and not x10 and not x1 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and x14 and x10 and x3 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and x14 and x10 and x3 and not x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and x14 and x10 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and x14 and not x10 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and not x14 and x10 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and not x14 and x10 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and x15 and not x14 and not x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and x11 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and x11 and not x3 and x5 and x7 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and x11 and not x3 and x5 and not x7 ) = '1' then
         current_otherm <= s268;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and x11 and not x3 and not x5 and x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and x11 and not x3 and not x5 and not x12 ) = '1' then
         current_otherm <= s268;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and not x11 and x10 and x5 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and not x11 and x10 and not x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and not x11 and not x10 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s78;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and not x11 and not x10 and not x1 and x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x13 and not x67 and not x15 and not x11 and not x10 and not x1 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x13 and not x3 and x5 and x7 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and not x13 and not x3 and x5 and not x7 ) = '1' then
         current_otherm <= s268;

      elsif ( not x62 and x63 and not x13 and not x3 and not x5 and x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s75;

      elsif ( not x62 and x63 and not x13 and not x3 and not x5 and not x12 ) = '1' then
         current_otherm <= s268;

      elsif ( not x62 and not x63 and x64 and x21 and x20 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s346;

      elsif ( not x62 and not x63 and x64 and x21 and not x20 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s345;

      elsif ( not x62 and not x63 and x64 and not x21 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s346;

      else
         y47 <= '1' ;
         y51 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s527;

      end if;

   when s269 =>
      if ( x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and x8 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and x8 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and x8 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and x8 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and x10 and x25 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and x10 and not x25 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and x10 and not x25 and x23 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and x10 and not x25 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and not x10 and x24 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and not x10 and not x24 and x23 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and not x10 and not x24 and x23 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and x9 and not x8 and not x10 and not x24 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and not x9 and x10 and x8 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and not x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s356;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and not x9 and not x10 and x8 ) = '1' then
         y10 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and x31 and not x11 and not x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s287;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and x12 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and x9 and x10 and x8 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s568;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and x9 and not x10 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s569;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and not x9 and x10 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and not x9 and x10 and not x8 and x27 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and not x9 and x10 and not x8 and not x27 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and not x9 and not x10 and x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s570;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and not x9 and not x10 and not x8 and x26 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and x22 and not x9 and not x10 and not x8 and not x26 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x63 and not x64 and x65 and x4 and x30 and not x31 and not x12 and not x22 ) = '1' then
         y45 <= '1' ;
         y47 <= '1' ;
         y50 <= '1' ;
         y60 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s571;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and x12 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and x10 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and x10 and not x8 and x21 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and x10 and not x8 and not x21 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and x10 and not x8 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and not x10 and x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and not x10 and not x8 and x18 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and not x10 and not x8 and not x18 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and x9 and not x10 and not x8 and not x18 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and x10 and x19 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and x10 and not x19 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and x10 and not x19 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and not x10 and x20 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and not x10 and not x20 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and x8 and not x10 and not x20 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and x31 and not x9 and not x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and x22 and not x31 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( not x63 and not x64 and x65 and x4 and not x30 and not x12 and not x22 ) = '1' then
         y45 <= '1' ;
         y47 <= '1' ;
         y50 <= '1' ;
         y60 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s571;

      elsif ( not x63 and not x64 and x65 and not x4 and x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s359;

      elsif ( not x63 and not x64 and x65 and not x4 and not x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x63 and not x64 and not x65 and x66 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and not x64 and not x65 and x66 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and not x64 and not x65 and x66 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x65 and x66 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x65 and not x66 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x65 and not x66 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and not x65 and not x66 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s270 =>
         y9 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s272;

   when s271 =>
      if ( x62 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      elsif ( not x62 and x12 and x15 and x13 and x3 ) = '1' then
         y3 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s273;

      elsif ( not x62 and x12 and x15 and x13 and not x3 and x14 ) = '1' then
         y3 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s273;

      elsif ( not x62 and x12 and x15 and x13 and not x3 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x12 and x15 and not x13 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( not x62 and x12 and not x15 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      else
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      end if;

   when s272 =>
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

   when s273 =>
         y11 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s461;

   when s274 =>
      if ( x62 and x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x62 and not x12 ) = '1' then
         current_otherm <= s274;

      elsif ( not x62 and x63 and x15 and x14 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( not x62 and x63 and x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s96;

      elsif ( not x62 and x63 and not x15 and x12 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x63 and not x15 and not x12 ) = '1' then
         current_otherm <= s274;

      elsif ( not x62 and not x63 and x30 and x31 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s321;

      elsif ( not x62 and not x63 and x30 and not x31 ) = '1' then
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s573;

      else
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s146;

      end if;

   when s275 =>
      if ( x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s276 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s277 =>
      if ( x10 ) = '1' then
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s574;

      elsif ( not x10 and x14 and x6 and x8 and x7 ) = '1' then
         y63 <= '1' ;
         current_otherm <= s224;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and x9 and not x18 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and x9 and not x18 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and x9 and not x18 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and x9 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and not x9 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and not x9 and not x19 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and not x9 and not x19 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and not x9 and not x19 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and x8 and not x7 and not x9 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and not x8 and x9 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s575;

      elsif ( not x10 and x14 and x6 and not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( not x10 and x14 and x6 and not x8 and not x9 and x7 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( not x10 and x14 and x6 and not x8 and not x9 and x7 and not x17 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x10 and x14 and x6 and not x8 and not x9 and x7 and not x17 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x10 and x14 and x6 and not x8 and not x9 and x7 and not x17 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and not x8 and not x9 and x7 and not x17 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and not x8 and not x9 and not x7 ) = '1' then
         y65 <= '1' ;
         current_otherm <= s155;

      elsif ( not x10 and x14 and not x6 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s576;

      end if;

   when s278 =>
      if ( x64 and x63 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x64 and x63 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x64 and x63 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and x63 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s577;

      elsif ( not x64 and x20 and x63 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x20 and not x63 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x20 and not x63 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x20 and not x63 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x20 and x63 and x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x64 and not x20 and x63 and not x19 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      else
         current_otherm <= s1;

      end if;

   when s279 =>
      if ( x63 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x64 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and x64 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and x64 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s578;

      end if;

   when s280 =>
      if ( x63 and x20 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x63 and not x20 and x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( x63 and not x20 and not x19 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      elsif ( not x63 and x64 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and x64 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and x64 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s281 =>
      if ( x64 and x6 and x8 and x27 and x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and x6 and x8 and x27 and not x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and x6 and x8 and not x27 and x7 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x64 and x6 and x8 and not x27 and not x7 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( x64 and x6 and not x8 and x27 and x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and x6 and not x8 and x27 and not x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and x6 and not x8 and not x27 and x7 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( x64 and x6 and not x8 and not x27 and not x7 ) = '1' then
         y18 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s580;

      elsif ( x64 and not x6 and x7 and x27 and x8 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and not x6 and x7 and x27 and not x8 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and not x6 and x7 and not x27 and x13 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x64 and not x6 and x7 and not x27 and x13 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x64 and not x6 and x7 and not x27 and x13 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x6 and x7 and not x27 and x13 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x6 and x7 and not x27 and x13 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x6 and x7 and not x27 and not x13 and x3 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x64 and not x6 and x7 and not x27 and not x13 and x3 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x64 and not x6 and x7 and not x27 and not x13 and x3 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x6 and x7 and not x27 and not x13 and x3 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x6 and x7 and not x27 and not x13 and x3 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x6 and x7 and not x27 and not x13 and not x3 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s581;

      elsif ( x64 and not x6 and not x7 and x27 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and not x6 and not x7 and not x27 and x8 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         y32 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s579;

      elsif ( x64 and not x6 and not x7 and not x27 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s579;

      else
         y57 <= '1' ;
         current_otherm <= s582;

      end if;

   when s282 =>
      if ( x63 and x65 and x11 ) = '1' then
         y55 <= '1' ;
         current_otherm <= s254;

      elsif ( x63 and x65 and not x11 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s387;

      elsif ( x63 and not x65 and x2 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( x63 and not x65 and not x2 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and not x2 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and not x2 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x65 and not x2 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and not x2 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x65 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x63 and x64 and x65 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x65 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s583;

      elsif ( not x63 and not x64 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x64 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s283 =>
      if ( x65 and x4 ) = '1' then
         y67 <= '1' ;
         current_otherm <= s584;

      elsif ( x65 and not x4 and x6 and x5 and x7 and x9 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      elsif ( x65 and not x4 and x6 and x5 and x7 and not x9 ) = '1' then
         y75 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and x9 and x12 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and x9 and not x12 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and x9 and not x12 and x20 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and x9 and not x12 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and not x9 and x13 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and not x9 and not x13 and x20 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and not x9 and not x13 and x20 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and x8 and not x9 and not x13 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and x6 and x5 and not x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s276;

      elsif ( x65 and not x4 and x6 and not x5 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s277;

      elsif ( x65 and not x4 and x6 and not x5 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s576;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and x8 and x9 and x5 and x7 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and x8 and x9 and x5 and not x7 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and x8 and x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and x8 and not x9 and x5 and x7 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and x8 and not x9 and x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and x8 and not x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and not x8 and x5 and x7 and x9 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and not x8 and x5 and x7 and not x9 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and not x8 and x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and x3 and x11 and not x8 and not x5 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s277;

      elsif ( x65 and not x4 and not x6 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s576;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and x8 and x9 and x5 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and x8 and x9 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and x8 and not x9 and x5 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and x8 and not x9 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and not x8 and x9 and x5 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and not x8 and x9 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and not x8 and not x9 and x5 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and x7 and not x8 and not x9 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and x8 and x9 and x5 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s153;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and x8 and x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and x8 and not x9 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and x8 and not x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and not x8 and x5 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and not x8 and x5 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s275;

      elsif ( x65 and not x4 and not x6 and not x3 and not x10 and not x7 and not x8 and not x5 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s275;

      elsif ( not x65 and x16 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( not x65 and not x16 and x21 and x20 and x4 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x65 and not x16 and x21 and x20 and x4 and not x6 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and x6 and x9 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and x6 and not x9 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and not x6 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and x5 and not x6 and not x8 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s585;

      elsif ( not x65 and not x16 and x21 and x20 and not x4 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y40 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s585;

      elsif ( not x65 and not x16 and x21 and not x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s586;

      elsif ( not x65 and not x16 and not x21 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s586;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and x5 and x6 and x4 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and x5 and x6 and not x4 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s585;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and x5 and not x6 and x4 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and x5 and not x6 and not x4 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and not x5 and x6 and x4 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s385;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and not x5 and x6 and not x4 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y30 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s587;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and not x5 and not x6 and x4 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s588;

      elsif ( not x65 and not x16 and not x21 and not x3 and x20 and not x5 and not x6 and not x4 ) = '1' then
         y3 <= '1' ;
         y20 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s589;

      elsif ( not x65 and not x16 and not x21 and not x3 and not x20 and x4 and x5 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x65 and not x16 and not x21 and not x3 and not x20 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      else
         y5 <= '1' ;
         y20 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      end if;

   when s284 =>
      if ( x64 and x65 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s346;

      elsif ( x64 and not x65 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s590;

      elsif ( not x64 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x64 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x64 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s285 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s591;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s592;

      end if;

   when s286 =>
      if ( x33 and x32 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s593;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s593;

      end if;

   when s287 =>
      if ( x62 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x62 and x63 and x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x62 and x63 and not x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and x64 and x20 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s594;

      elsif ( not x62 and not x63 and x64 and x20 and not x3 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s284;

      elsif ( not x62 and not x63 and x64 and not x20 and x21 and x3 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s416;

      elsif ( not x62 and not x63 and x64 and not x20 and x21 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s486;

      elsif ( not x62 and not x63 and x64 and not x20 and not x21 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( not x62 and not x63 and x64 and not x20 and not x21 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s595;

      elsif ( not x62 and not x63 and not x64 and x31 ) = '1' then
         y47 <= '1' ;
         y54 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s596;

      else
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s597;

      end if;

   when s288 =>
      if ( x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x62 and x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s289 =>
      if ( x64 ) = '1' then
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s598;

      else
         y33 <= '1' ;
         current_otherm <= s321;

      end if;

   when s290 =>
      if ( x64 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x30 ) = '1' then
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      elsif ( not x64 and not x30 and x31 ) = '1' then
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s600;

      else
         y33 <= '1' ;
         current_otherm <= s321;

      end if;

   when s291 =>
      if ( x65 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y69 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s601;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s602;

      end if;

   when s292 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s603;

   when s293 =>
         y7 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s604;

   when s294 =>
      if ( x21 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x21 and not x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s605;

      elsif ( not x21 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s606;

      else
         y15 <= '1' ;
         current_otherm <= s111;

      end if;

   when s295 =>
         y15 <= '1' ;
         current_otherm <= s111;

   when s296 =>
      if ( x62 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x62 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x20 and x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s607;

      else
         y14 <= '1' ;
         current_otherm <= s594;

      end if;

   when s297 =>
         y3 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s608;

   when s298 =>
      if ( x13 and x10 and x12 and x11 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s53;

      elsif ( x13 and x10 and x12 and not x11 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and x10 and x12 and not x11 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( x13 and x10 and x12 and not x11 and not x3 and not x6 ) = '1' then
         current_otherm <= s298;

      elsif ( x13 and x10 and not x12 and x11 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and x10 and not x12 and x11 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( x13 and x10 and not x12 and x11 and not x3 and not x6 ) = '1' then
         current_otherm <= s298;

      elsif ( x13 and x10 and not x12 and not x11 and x14 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and x10 and not x12 and not x11 and x14 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( x13 and x10 and not x12 and not x11 and x14 and not x3 and not x6 ) = '1' then
         current_otherm <= s298;

      elsif ( x13 and x10 and not x12 and not x11 and not x14 and x1 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s244;

      elsif ( x13 and x10 and not x12 and not x11 and not x14 and not x1 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and not x10 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( x13 and not x10 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      elsif ( x13 and not x10 and not x3 and not x6 ) = '1' then
         current_otherm <= s298;

      elsif ( not x13 and x3 ) = '1' then
         y22 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s58;

      elsif ( not x13 and not x3 and x6 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s55;

      else
         current_otherm <= s298;

      end if;

   when s299 =>
      if ( x2 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s243;

      else
         current_otherm <= s299;

      end if;

   when s300 =>
      if ( x11 and x12 and x4 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( x11 and x12 and not x4 ) = '1' then
         current_otherm <= s300;

      elsif ( x11 and not x12 and x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and not x12 and not x13 and x4 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( x11 and not x12 and not x13 and not x4 ) = '1' then
         current_otherm <= s300;

      elsif ( not x11 and x14 and x4 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( not x11 and x14 and not x4 ) = '1' then
         current_otherm <= s300;

      elsif ( not x11 and not x14 and x12 and x4 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( not x11 and not x14 and x12 and not x4 ) = '1' then
         current_otherm <= s300;

      elsif ( not x11 and not x14 and not x12 and x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and not x14 and not x12 and not x13 and x4 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      else
         current_otherm <= s300;

      end if;

   when s301 =>
         y9 <= '1' ;
         y21 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s609;

   when s302 =>
      if ( x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s303 =>
         y5 <= '1' ;
         current_otherm <= s331;

   when s304 =>
         y4 <= '1' ;
         y13 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s610;

   when s305 =>
      if ( x17 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s306 =>
      if ( x9 and x21 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s611;

      elsif ( x9 and x21 and not x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s612;

      elsif ( x9 and not x21 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s607;

      elsif ( x9 and not x21 and not x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s149;

      else
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s294;

      end if;

   when s307 =>
      if ( x3 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s64;

      elsif ( x3 and x2 and not x1 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s197;

      elsif ( x3 and not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s307;

      elsif ( x3 and not x2 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      end if;

   when s308 =>
      if ( x64 and x62 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s613;

      elsif ( x64 and not x62 and x66 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( x64 and not x62 and not x66 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s614;

      elsif ( not x64 and x62 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s615;

      elsif ( not x64 and not x62 and x30 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s321;

      elsif ( not x64 and not x62 and not x30 and x31 ) = '1' then
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s501;

      else
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      end if;

   when s309 =>
         y14 <= '1' ;
         current_otherm <= s95;

   when s310 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s533;

      elsif ( x62 and not x64 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s616;

      elsif ( not x62 and x64 and x5 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s60;

      elsif ( not x62 and x64 and not x5 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x64 and x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      else
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      end if;

   when s311 =>
         y13 <= '1' ;
         current_otherm <= s617;

   when s312 =>
         y23 <= '1' ;
         current_otherm <= s169;

   when s313 =>
         y21 <= '1' ;
         current_otherm <= s262;

   when s314 =>
         y1 <= '1' ;
         y15 <= '1' ;
         y37 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s618;

   when s315 =>
      if ( x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s316 =>
      if ( x36 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s619;

      elsif ( not x36 and x38 and x39 and x41 and x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s620;

      elsif ( not x36 and x38 and x39 and x41 and not x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s315;

      elsif ( not x36 and x38 and x39 and not x41 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s539;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and x56 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and not x56 and x58 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and not x56 and not x58 and x59 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x36 and x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and x57 and x28 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and not x57 and x29 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and not x54 and x53 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x36 and x38 and not x39 and x40 and not x55 and not x54 and not x53 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x36 and x38 and not x39 and not x40 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s621;

      else
         y2 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s622;

      end if;

   when s317 =>
      if ( x10 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s623;

      elsif ( not x10 and x11 and x14 and x30 and x36 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x10 and x11 and x14 and x30 and not x36 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and x33 and x34 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s90;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and x33 and not x34 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and x33 and not x34 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and x33 and not x34 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and x33 and not x34 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and not x33 and x35 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and not x33 and not x35 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and not x33 and not x35 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and not x33 and not x35 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x14 and not x30 and x31 and not x33 and not x35 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x11 and x14 and not x30 and not x31 and x32 ) = '1' then
         y1 <= '1' ;
         y22 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s312;

      elsif ( not x10 and x11 and x14 and not x30 and not x31 and not x32 ) = '1' then
         y1 <= '1' ;
         y20 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s313;

      elsif ( not x10 and x11 and not x14 and x15 and x16 and x20 and x22 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x10 and x11 and not x14 and x15 and x16 and x20 and not x22 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s521;

      elsif ( not x10 and x11 and not x14 and x15 and x16 and not x20 and x21 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x10 and x11 and not x14 and x15 and x16 and not x20 and not x21 ) = '1' then
         y37 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s315;

      elsif ( not x10 and x11 and not x14 and x15 and not x16 and x17 and x19 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s624;

      elsif ( not x10 and x11 and not x14 and x15 and not x16 and x17 and not x19 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y44 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s315;

      elsif ( not x10 and x11 and not x14 and x15 and not x16 and not x17 and x18 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s315;

      elsif ( not x10 and x11 and not x14 and x15 and not x16 and not x17 and not x18 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x10 and x11 and not x14 and not x15 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y37 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s625;

      elsif ( not x10 and not x11 and x12 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y37 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s625;

      elsif ( not x10 and not x11 and not x12 and x13 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y37 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s625;

      elsif ( not x10 and not x11 and not x12 and not x13 and x43 and x46 and x48 ) = '1' then
         y37 <= '1' ;
         y39 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s626;

      elsif ( not x10 and not x11 and not x12 and not x13 and x43 and x46 and not x48 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s627;

      elsif ( not x10 and not x11 and not x12 and not x13 and x43 and not x46 and x47 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s628;

      elsif ( not x10 and not x11 and not x12 and not x13 and x43 and not x46 and not x47 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s629;

      elsif ( not x10 and not x11 and not x12 and not x13 and not x43 and x44 and x45 ) = '1' then
         y19 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s315;

      elsif ( not x10 and not x11 and not x12 and not x13 and not x43 and x44 and not x45 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s315;

      else
         y14 <= '1' ;
         y31 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s315;

      end if;

   when s318 =>
      if ( x65 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x17 and x18 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s20;

      elsif ( not x65 and x17 and x18 and not x1 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      elsif ( not x65 and x17 and x18 and not x1 and not x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s24;

      elsif ( not x65 and x17 and not x18 and x6 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s126;

      elsif ( not x65 and x17 and not x18 and not x6 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s105;

      else
         y2 <= '1' ;
         current_otherm <= s24;

      end if;

   when s319 =>
         y65 <= '1' ;
         y90 <= '1' ;
         y92 <= '1' ;
         y98 <= '1' ;
         y99 <= '1' ;
         current_otherm <= s240;

   when s320 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s304;

      elsif ( not x62 and x63 and x14 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s470;

      elsif ( not x62 and x63 and not x14 ) = '1' then
         y28 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s630;

      else
         y24 <= '1' ;
         current_otherm <= s117;

      end if;

   when s321 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s631;

      elsif ( not x63 and not x64 and x66 ) = '1' then
         y47 <= '1' ;
         y51 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s632;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      end if;

   when s322 =>
      if ( x64 and x66 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s633;

      elsif ( x64 and not x66 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      else
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s573;

      end if;

   when s323 =>
         y7 <= '1' ;
         y10 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1;

   when s324 =>
         y3 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s634;

   when s325 =>
      if ( x63 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x63 and x67 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s291;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s602;

      end if;

   when s326 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s635;

   when s327 =>
         y3 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s128;

   when s328 =>
         y3 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s91;

   when s329 =>
      if ( x3 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s636;

      else
         y6 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s637;

      end if;

   when s330 =>
         y13 <= '1' ;
         current_otherm <= s204;

   when s331 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s638;

      elsif ( not x62 and x63 and x67 and x14 and x13 and x11 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( not x62 and x63 and x67 and x14 and x13 and x11 and not x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and x10 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and not x10 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and not x10 and not x3 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and x67 and x14 and x13 and not x11 and not x10 and not x3 and not x6 ) = '1' then
         current_otherm <= s331;

      elsif ( not x62 and x63 and x67 and x14 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and x14 and not x13 and not x3 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and x67 and x14 and not x13 and not x3 and not x6 ) = '1' then
         current_otherm <= s331;

      elsif ( not x62 and x63 and x67 and not x14 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and x67 and not x14 and not x3 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and x67 and not x14 and not x3 and not x6 ) = '1' then
         current_otherm <= s331;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and x14 and x10 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and x14 and not x10 and x1 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and x14 and not x10 and not x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and not x14 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and not x14 and not x3 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and not x67 and x15 and x13 and not x14 and not x3 and not x6 ) = '1' then
         current_otherm <= s331;

      elsif ( not x62 and x63 and not x67 and x15 and not x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and x15 and not x13 and not x3 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and not x67 and x15 and not x13 and not x3 and not x6 ) = '1' then
         current_otherm <= s331;

      elsif ( not x62 and x63 and not x67 and not x15 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s77;

      elsif ( not x62 and x63 and not x67 and not x15 and not x3 and x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s73;

      elsif ( not x62 and x63 and not x67 and not x15 and not x3 and not x6 ) = '1' then
         current_otherm <= s331;

      elsif ( not x62 and not x63 and x64 and x21 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s639;

      elsif ( not x62 and not x63 and x64 and not x21 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s640;

      else
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      end if;

   when s332 =>
         y46 <= '1' ;
         current_otherm <= s390;

   when s333 =>
      if ( x67 and x11 and x5 and x6 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x67 and x11 and x5 and not x6 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x67 and x11 and x5 and not x6 and not x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( x67 and x11 and not x5 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      elsif ( x67 and x11 and not x5 and not x4 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      elsif ( x67 and not x11 and x4 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x67 and not x11 and not x4 ) = '1' then
         current_otherm <= s333;

      elsif ( not x67 and x10 and x4 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x67 and x10 and not x4 ) = '1' then
         current_otherm <= s333;

      elsif ( not x67 and not x10 and x5 and x6 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x67 and not x10 and x5 and not x6 and x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x67 and not x10 and x5 and not x6 and not x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s161;

      elsif ( not x67 and not x10 and not x5 and x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      else
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s333;

      end if;

   when s334 =>
         y13 <= '1' ;
         current_otherm <= s641;

   when s335 =>
      if ( x62 and x61 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( x62 and not x61 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s642;

      elsif ( not x62 and x63 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s643;

      else
         y29 <= '1' ;
         current_otherm <= s378;

      end if;

   when s336 =>
      if ( x62 and x65 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s644;

      elsif ( x62 and not x65 ) = '1' then
         y9 <= '1' ;
         y21 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s645;

      else
         y7 <= '1' ;
         current_otherm <= s646;

      end if;

   when s337 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s303;

      elsif ( not x62 and x65 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s476;

      else
         y12 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s647;

      end if;

   when s338 =>
      if ( x2 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      else
         current_otherm <= s338;

      end if;

   when s339 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

   when s340 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

   when s341 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s648;

   when s342 =>
      if ( x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s343 =>
      if ( x64 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      else
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s330;

      end if;

   when s344 =>
      if ( x22 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s650;

      else
         y10 <= '1' ;
         current_otherm <= s651;

      end if;

   when s345 =>
      if ( x63 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s247;

      elsif ( x63 and not x16 ) = '1' then
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s248;

      elsif ( not x63 and x64 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s652;

      else
         y22 <= '1' ;
         current_otherm <= s171;

      end if;

   when s346 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s359;

      elsif ( not x62 and x63 and x16 and x22 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s557;

      elsif ( not x62 and x63 and x16 and x22 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s251;

      elsif ( not x62 and x63 and x16 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s247;

      elsif ( not x62 and x63 and not x16 and x22 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s252;

      elsif ( not x62 and x63 and not x16 and not x22 ) = '1' then
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s248;

      else
         y7 <= '1' ;
         current_otherm <= s45;

      end if;

   when s347 =>
      if ( x16 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s349;

      elsif ( x16 and not x15 and x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( x16 and not x15 and not x3 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      elsif ( not x16 and x15 and x11 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x16 and x15 and not x11 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s348;

      elsif ( not x16 and x15 and not x11 and not x10 ) = '1' then
         current_otherm <= s347;

      else
         current_otherm <= s1;

      end if;

   when s348 =>
      if ( x62 and x4 and x5 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( x62 and x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s653;

      elsif ( x62 and not x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s214;

      elsif ( not x62 and x16 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x16 and not x15 and x4 and x5 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and x16 and not x15 and x4 and not x5 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x62 and x16 and not x15 and not x4 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s218;

      elsif ( not x62 and not x16 and x15 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      elsif ( not x62 and not x16 and not x15 and x12 and x13 and x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s349;

      elsif ( not x62 and not x16 and not x15 and x12 and x13 and not x3 and x14 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s349;

      elsif ( not x62 and not x16 and not x15 and x12 and x13 and not x3 and not x14 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( not x62 and not x16 and not x15 and x12 and not x13 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s29;

      else
         y4 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s27;

      end if;

   when s349 =>
      if ( x62 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s221;

      elsif ( not x62 and x15 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s28;

      elsif ( not x62 and not x15 and x16 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s31;

      else
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s212;

      end if;

   when s350 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s642;

      elsif ( not x62 and x65 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x62 and not x65 and x67 ) = '1' then
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s654;

      else
         y12 <= '1' ;
         current_otherm <= s11;

      end if;

   when s351 =>
      if ( x63 and x18 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s655;

      elsif ( x63 and not x18 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s656;

      else
         y4 <= '1' ;
         y31 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s657;

      end if;

   when s352 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s540;

      elsif ( x62 and not x64 and x66 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s658;

      elsif ( x62 and not x64 and not x66 and x6 and x3 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x62 and not x64 and not x66 and x6 and not x3 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s18;

      elsif ( x62 and not x64 and not x66 and x6 and not x3 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s124;

      elsif ( x62 and not x64 and not x66 and not x6 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( not x62 and x30 ) = '1' then
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      elsif ( not x62 and not x30 and x31 ) = '1' then
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s600;

      else
         y33 <= '1' ;
         current_otherm <= s321;

      end if;

   when s353 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s615;

   when s354 =>
      if ( x62 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x11 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x63 and x11 and not x18 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      elsif ( not x62 and x63 and not x11 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and x9 and x10 and x8 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s568;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and x9 and not x10 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s569;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and not x9 and x10 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and not x9 and x10 and not x8 and x27 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and not x9 and x10 and not x8 and not x27 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and not x9 and not x10 and x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s570;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and not x9 and not x10 and not x8 and x26 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x62 and not x63 and not x64 and x30 and x4 and not x9 and not x10 and not x8 and not x26 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x62 and not x63 and not x64 and x30 and not x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s366;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and x10 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and x10 and not x8 and x21 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and x10 and not x8 and not x21 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and x10 and not x8 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and not x10 and x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and not x10 and not x8 and x18 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and not x10 and not x8 and not x18 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and x9 and not x10 and not x8 and not x18 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and x10 and x19 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and x10 and not x19 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and x10 and not x19 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and not x10 and x20 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and not x10 and not x20 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and x8 and not x10 and not x20 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and x31 and not x9 and not x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x62 and not x63 and not x64 and not x30 and x4 and not x31 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( not x62 and not x63 and not x64 and not x30 and not x4 and x31 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s308;

      else
         y5 <= '1' ;
         current_otherm <= s359;

      end if;

   when s355 =>
      if ( x63 and x11 ) = '1' then
         y14 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s659;

      elsif ( x63 and not x11 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s660;

      elsif ( x63 and not x11 and not x15 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x63 and not x11 and not x15 and not x18 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      else
         y25 <= '1' ;
         current_otherm <= s661;

      end if;

   when s356 =>
      if ( x64 and x3 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s662;

      elsif ( x64 and not x3 and x20 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( x64 and not x3 and not x20 and x21 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and not x3 and not x20 and not x21 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s167;

      elsif ( not x64 and x31 ) = '1' then
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y69 <= '1' ;
         current_otherm <= s368;

      else
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s487;

      end if;

   when s357 =>
      if ( x66 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x66 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s663;

      elsif ( not x66 and not x22 and x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s664;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s663;

      end if;

   when s358 =>
      if ( x63 ) = '1' then
         y9 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1;

      else
         y6 <= '1' ;
         current_otherm <= s345;

      end if;

   when s359 =>
      if ( x64 and x62 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s665;

      elsif ( x64 and not x62 and x21 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s666;

      elsif ( x64 and not x62 and not x21 and x22 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s640;

      elsif ( x64 and not x62 and not x21 and not x22 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s639;

      elsif ( not x64 and x62 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s86;

      elsif ( not x64 and not x62 and x31 and x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      elsif ( not x64 and not x62 and x31 and not x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s667;

      elsif ( not x64 and not x62 and not x31 and x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s146;

      else
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s501;

      end if;

   when s360 =>
      if ( x64 and x63 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x63 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x63 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x63 and x66 and x10 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x64 and x63 and x66 and not x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      elsif ( not x64 and x63 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and x63 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and x63 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x64 and x63 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and x63 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and x63 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x65 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x63 and x65 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x63 and x65 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and x65 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and not x65 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x63 and not x65 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x63 and not x65 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x63 and not x65 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s361 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s398;

      else
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s668;

      end if;

   when s362 =>
      if ( x21 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s669;

      elsif ( not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s363 =>
      if ( x64 and x21 and x17 and x16 and x19 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and x21 and x17 and x16 and x19 and not x11 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and x21 and x17 and x16 and not x19 and x18 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and x21 and x17 and x16 and not x19 and not x18 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and x21 and x17 and not x16 and x11 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( x64 and x21 and x17 and not x16 and not x11 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s365;

      elsif ( x64 and x21 and not x17 and x16 and x19 and x14 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and x21 and not x17 and x16 and x19 and not x14 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and x21 and not x17 and x16 and not x19 and x13 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x64 and x21 and not x17 and x16 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and x21 and not x17 and not x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x64 and not x21 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s185;

      elsif ( not x64 and x30 and x31 and x14 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and x30 and x31 and not x14 ) = '1' then
         y47 <= '1' ;
         y54 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s596;

      elsif ( not x64 and x30 and not x31 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x30 and not x31 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x30 and not x31 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x30 and not x31 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x30 and not x31 and not x14 ) = '1' then
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s597;

      else
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s487;

      end if;

   when s364 =>
      if ( x64 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s606;

      elsif ( not x64 and x30 and x31 ) = '1' then
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      elsif ( not x64 and x30 and not x31 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s670;

      else
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s573;

      end if;

   when s365 =>
      if ( x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s346;

      else
         y47 <= '1' ;
         y51 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s671;

      end if;

   when s366 =>
      if ( x64 and x62 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s672;

      elsif ( x64 and not x62 and x21 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s240;

      elsif ( x64 and not x62 and not x21 and x22 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s639;

      elsif ( x64 and not x62 and not x21 and not x22 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s673;

      elsif ( not x64 and x62 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s674;

      elsif ( not x64 and not x62 and x30 ) = '1' then
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s501;

      elsif ( not x64 and not x62 and not x30 and x31 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s675;

      else
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      end if;

   when s367 =>
      if ( x6 and x3 and x7 and x9 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x6 and x3 and x7 and not x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( x6 and x3 and not x7 and x8 and x9 and x11 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( x6 and x3 and not x7 and x8 and x9 and not x11 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and x3 and not x7 and x8 and x9 and not x11 and x14 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x3 and not x7 and x8 and x9 and not x11 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x3 and not x7 and x8 and not x9 and x10 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( x6 and x3 and not x7 and x8 and not x9 and not x10 and x14 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and x3 and not x7 and x8 and not x9 and not x10 and x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x3 and not x7 and x8 and not x9 and not x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x3 and not x7 and not x8 and x9 ) = '1' then
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s676;

      elsif ( x6 and x3 and not x7 and not x8 and not x9 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s677;

      elsif ( x6 and not x3 and x8 and x9 and x15 and x16 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and x8 and x9 and x15 and x16 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and x8 and x9 and x15 and x16 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and x8 and x9 and x15 and x16 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and x8 and x9 and x15 and not x16 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s678;

      elsif ( x6 and not x3 and x8 and x9 and not x15 and x7 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x6 and not x3 and x8 and x9 and not x15 and not x7 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s677;

      elsif ( x6 and not x3 and x8 and not x9 and x15 and x17 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s678;

      elsif ( x6 and not x3 and x8 and not x9 and x15 and not x17 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and x8 and not x9 and x15 and not x17 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and x8 and not x9 and x15 and not x17 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and x8 and not x9 and x15 and not x17 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and x8 and not x9 and not x15 and x7 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x6 and not x3 and x8 and not x9 and not x15 and not x7 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s57;

      elsif ( x6 and not x3 and not x8 and x9 and x15 and x18 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s678;

      elsif ( x6 and not x3 and not x8 and x9 and x15 and not x18 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and not x8 and x9 and x15 and not x18 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and not x8 and x9 and x15 and not x18 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and not x8 and x9 and x15 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and not x8 and x9 and not x15 and x7 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( x6 and not x3 and not x8 and x9 and not x15 and not x7 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s679;

      elsif ( x6 and not x3 and not x8 and not x9 and x15 and x18 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and not x8 and not x9 and x15 and x18 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x6 and not x3 and not x8 and not x9 and x15 and x18 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and not x8 and not x9 and x15 and x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x3 and not x8 and not x9 and x15 and not x18 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s678;

      elsif ( x6 and not x3 and not x8 and not x9 and not x15 and x7 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x6 and not x3 and not x8 and not x9 and not x15 and not x7 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x6 and x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s680;

      elsif ( not x6 and not x3 and x12 and x4 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s681;

      elsif ( not x6 and not x3 and x12 and not x4 and x5 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s682;

      elsif ( not x6 and not x3 and x12 and not x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s677;

      elsif ( not x6 and not x3 and not x12 and x4 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s677;

      elsif ( not x6 and not x3 and not x12 and x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s683;

      else
         y1 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s684;

      end if;

   when s368 =>
         y43 <= '1' ;
         current_otherm <= s175;

   when s369 =>
      if ( x14 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( not x14 and x7 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s99;

      elsif ( not x14 and not x7 and x3 and x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s17;

      elsif ( not x14 and not x7 and x3 and x1 and not x2 and x5 ) = '1' then
         current_otherm <= s369;

      elsif ( not x14 and not x7 and x3 and x1 and not x2 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s7;

      elsif ( not x14 and not x7 and x3 and not x1 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s9;

      end if;

   when s370 =>
      if ( x11 ) = '1' then
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s369;

      else
         y10 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s370;

      end if;

   when s371 =>
      if ( x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s568;

      else
         y7 <= '1' ;
         current_otherm <= s288;

      end if;

   when s372 =>
      if ( x3 and x6 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x6 and not x5 and x8 and x7 and x10 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s687;

      elsif ( x3 and x6 and not x5 and x8 and x7 and x10 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( x3 and x6 and not x5 and x8 and x7 and not x10 ) = '1' then
         y72 <= '1' ;
         current_otherm <= s685;

      elsif ( x3 and x6 and not x5 and x8 and not x7 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( x3 and x6 and not x5 and x8 and not x7 and x9 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x6 and not x5 and x8 and not x7 and not x9 and x17 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( x3 and x6 and not x5 and x8 and not x7 and not x9 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x6 and not x5 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( x3 and x6 and not x5 and not x8 and not x9 and x7 and x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( x3 and x6 and not x5 and not x8 and not x9 and x7 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x6 and not x5 and not x8 and not x9 and not x7 ) = '1' then
         y71 <= '1' ;
         current_otherm <= s156;

      elsif ( x3 and not x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s687;

      elsif ( x3 and not x6 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( not x3 and x4 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s201;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s688;

      end if;

   when s373 =>
         y22 <= '1' ;
         current_otherm <= s689;

   when s374 =>
         y13 <= '1' ;
         current_otherm <= s101;

   when s375 =>
      if ( x62 and x17 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s690;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s566;

      elsif ( not x62 and x64 ) = '1' then
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s691;

      else
         y13 <= '1' ;
         current_otherm <= s692;

      end if;

   when s376 =>
      if ( x62 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and x65 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x65 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x64 and not x63 and not x65 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and x64 and not x63 and not x65 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and x64 and not x63 and not x65 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x63 and not x65 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and x63 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and not x64 and x63 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x63 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and not x63 and x65 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s623;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x64 and not x63 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s377 =>
      if ( x64 and x62 and x66 and x32 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x64 and x62 and x66 and not x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( x64 and x62 and not x66 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x64 and x62 and not x66 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x64 and x62 and not x66 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and x62 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x63 and x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( x64 and not x62 and x63 and not x9 and x20 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( x64 and not x62 and x63 and not x9 and not x20 and x21 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s63;

      elsif ( x64 and not x62 and x63 and not x9 and not x20 and not x21 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( x64 and not x62 and not x63 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and not x62 and not x63 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and not x62 and not x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and not x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x62 and x60 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s288;

      elsif ( not x64 and x62 and not x60 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x64 and x62 and not x60 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x64 and x62 and not x60 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x62 and not x60 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x65 and x63 and x66 and x30 and x4 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s660;

      elsif ( not x64 and not x62 and x65 and x63 and x66 and x30 and not x4 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x64 and not x62 and x65 and x63 and x66 and not x30 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x64 and not x62 and x65 and x63 and x66 and not x30 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x62 and x65 and x63 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and not x62 and x65 and x63 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and not x62 and x65 and x63 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x64 and not x62 and x65 and x63 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x65 and x63 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x65 and x63 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x65 and not x63 and x67 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x64 and not x62 and x65 and not x63 and x67 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x64 and not x62 and x65 and not x63 and x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x65 and not x63 and x67 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x65 and not x63 and not x67 and x17 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x64 and not x62 and x65 and not x63 and not x67 and not x17 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x62 and x65 and not x63 and not x67 and not x17 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x62 and x65 and not x63 and not x67 and not x17 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x65 and not x63 and not x67 and not x17 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and x63 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x64 and not x62 and not x65 and x63 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x64 and not x62 and not x65 and x63 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and x63 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x65 and not x63 and x66 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and not x62 and not x65 and not x63 and not x66 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s378 =>
      if ( x64 and x62 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and x62 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x64 and x62 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and x62 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x63 and x65 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s693;

      elsif ( x64 and not x62 and x63 and not x65 and x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and not x62 and x63 and not x65 and x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x64 and not x62 and x63 and not x65 and x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x63 and not x65 and x21 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and x63 and not x65 and not x21 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s375;

      elsif ( x64 and not x62 and not x63 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and not x62 and not x63 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and not x62 and not x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x62 and not x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x64 and x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x64 and x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and x63 and x66 and x14 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x64 and not x62 and x63 and x66 and x14 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x62 and x63 and x66 and not x14 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x64 and not x62 and x63 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and not x62 and x63 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x64 and not x62 and x63 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x64 and not x62 and x63 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x63 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x64 and not x62 and x63 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x63 and x65 and x67 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x64 and not x62 and not x63 and x65 and not x67 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x62 and not x63 and x65 and not x67 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and not x62 and not x63 and x65 and not x67 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x63 and x65 and not x67 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x63 and not x65 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x63 and not x65 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x64 and not x62 and not x63 and not x65 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x62 and not x63 and not x65 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s379 =>
      if ( x64 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x30 ) = '1' then
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s501;

      elsif ( not x64 and not x30 and x31 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s365;

      else
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      end if;

   when s380 =>
      if ( x14 and x65 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x14 and x65 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x14 and x65 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x65 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x14 and not x65 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x14 and not x65 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s381 =>
      if ( x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s382 =>
      if ( x63 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( not x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s383 =>
      if ( x63 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s694;

      else
         y5 <= '1' ;
         current_otherm <= s398;

      end if;

   when s384 =>
      if ( x62 and x1 and x2 and x3 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x62 and x1 and x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s245;

      elsif ( x62 and x1 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_otherm <= s10;

      elsif ( x62 and not x1 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s695;

      end if;

   when s385 =>
      if ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and x3 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and x3 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and x3 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and x3 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and x18 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and x21 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and not x4 and x5 and x3 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and not x4 and not x5 and x3 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x64 and x19 and x20 and x2 and x1 and not x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y34 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x64 and x19 and x20 and x2 and not x1 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( x63 and x64 and x19 and x20 and not x2 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s696;

      elsif ( x63 and x64 and x19 and x20 and not x2 and not x8 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( x63 and x64 and x19 and not x20 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s697;

      elsif ( x63 and x64 and not x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s698;

      elsif ( x63 and not x64 and x66 and x31 and x15 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x63 and not x64 and x66 and x31 and not x15 and x16 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x63 and not x64 and x66 and x31 and not x15 and not x16 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s386;

      elsif ( x63 and not x64 and x66 and not x31 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x63 and not x64 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x64 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x64 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and not x64 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x64 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x64 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s386 =>
      if ( x63 and x65 and x17 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( x63 and x65 and not x17 and x14 ) = '1' then
         y38 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s699;

      elsif ( x63 and x65 and not x17 and not x14 ) = '1' then
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s700;

      elsif ( x63 and not x65 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s701;

      elsif ( not x63 and x4 and x11 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x63 and x4 and not x11 and x30 and x12 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and x9 and x10 and x8 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s425;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s702;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and x9 and not x10 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s703;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and not x9 and x10 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and not x9 and x10 and not x8 and x27 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and not x9 and x10 and not x8 and not x27 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and not x9 and not x10 and x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s704;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and not x9 and not x10 and not x8 and x26 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( not x63 and x4 and not x11 and x30 and not x12 and not x9 and not x10 and not x8 and not x26 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s38;

      elsif ( not x63 and x4 and not x11 and not x30 and x31 and x15 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s95;

      elsif ( not x63 and x4 and not x11 and not x30 and x31 and not x15 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s199;

      elsif ( not x63 and x4 and not x11 and not x30 and not x31 and x8 and x9 ) = '1' then
         y47 <= '1' ;
         y55 <= '1' ;
         y63 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s512;

      elsif ( not x63 and x4 and not x11 and not x30 and not x31 and x8 and not x9 ) = '1' then
         y47 <= '1' ;
         y56 <= '1' ;
         y63 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s512;

      elsif ( not x63 and x4 and not x11 and not x30 and not x31 and not x8 and x12 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s534;

      elsif ( not x63 and x4 and not x11 and not x30 and not x31 and not x8 and not x12 ) = '1' then
         y45 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         y55 <= '1' ;
         y60 <= '1' ;
         y63 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s512;

      elsif ( not x63 and not x4 and x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s310;

      elsif ( not x63 and not x4 and not x30 and x31 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      else
         y5 <= '1' ;
         current_otherm <= s308;

      end if;

   when s387 =>
      if ( x63 and x64 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s641;

      elsif ( x63 and not x64 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s388 =>
      if ( x63 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y22 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s705;

      elsif ( not x63 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s389 =>
      if ( x13 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x13 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x13 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x13 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s390 =>
      if ( x63 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s391 =>
      if ( x63 and x66 and x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( x63 and x66 and not x19 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( x63 and not x66 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s706;

      elsif ( not x63 and x65 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s707;

      elsif ( not x63 and not x65 and x66 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x65 and x66 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x65 and x66 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x66 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x66 and x67 and x17 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( not x63 and not x65 and not x66 and x67 and not x17 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and not x65 and not x66 and x67 and not x17 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and not x65 and not x66 and x67 and not x17 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x66 and x67 and not x17 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x66 and not x67 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and not x65 and not x66 and not x67 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and not x65 and not x66 and not x67 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s392 =>
      if ( x62 and x24 and x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      elsif ( x62 and x24 and x2 and not x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x62 and x24 and not x2 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x62 and not x24 and x2 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x62 and not x24 and not x2 and x3 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x62 and not x24 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x62 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s709;

      elsif ( not x62 and x19 and not x18 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s708;

      else
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s709;

      end if;

   when s393 =>
      if ( x21 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s359;

      elsif ( x21 and not x3 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s666;

      elsif ( not x21 and x22 and x3 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y96 <= '1' ;
         current_otherm <= s710;

      elsif ( not x21 and x22 and not x3 ) = '1' then
         y60 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y79 <= '1' ;
         current_otherm <= s710;

      elsif ( not x21 and not x22 and x3 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y96 <= '1' ;
         current_otherm <= s711;

      else
         y60 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y79 <= '1' ;
         current_otherm <= s711;

      end if;

   when s394 =>
      if ( x62 and x33 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s148;

      elsif ( x62 and not x33 and x32 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s148;

      elsif ( x62 and not x33 and not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and not x33 and not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and not x33 and not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x33 and not x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s395 =>
      if ( x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s396 =>
         y6 <= '1' ;
         y25 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s712;

   when s397 =>
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s192;

   when s398 =>
      if ( x62 and x64 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s374;

      elsif ( x62 and not x64 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s713;

      elsif ( not x62 and x64 and x21 and x20 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x62 and x64 and x21 and not x20 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s432;

      elsif ( not x62 and x64 and not x21 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x62 and not x64 and x30 and x31 ) = '1' then
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      elsif ( not x62 and not x64 and x30 and not x31 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s670;

      else
         y24 <= '1' ;
         current_otherm <= s714;

      end if;

   when s399 =>
      if ( x64 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s715;

      elsif ( not x64 and x19 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s585;

      elsif ( not x64 and x19 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x64 and x19 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s716;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and x6 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and x6 and not x5 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and not x6 and x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s719;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and not x6 and not x5 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and x6 and x5 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and x6 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and not x6 and x5 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x19 and not x20 and not x4 and x21 and not x6 and not x5 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x64 and x19 and not x20 and not x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s720;

      end if;

   when s400 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x8 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s721;

      elsif ( not x32 and not x8 and x33 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s394;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s721;

      end if;

   when s401 =>
      if ( x62 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s402 =>
         y35 <= '1' ;
         current_otherm <= s386;

   when s403 =>
      if ( x17 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s406;

      else
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s403;

      end if;

   when s404 =>
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s722;

   when s405 =>
      if ( x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      else
         current_otherm <= s1;

      end if;

   when s406 =>
      if ( x64 and x66 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s723;

      elsif ( x64 and not x66 ) = '1' then
         y2 <= '1' ;
         y15 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s724;

      else
         y25 <= '1' ;
         current_otherm <= s150;

      end if;

   when s407 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s410;

   when s408 =>
      if ( x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s409 =>
      if ( x65 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      else
         y51 <= '1' ;
         current_otherm <= s279;

      end if;

   when s410 =>
         y2 <= '1' ;
         y15 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s725;

   when s411 =>
      if ( x63 and x17 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s617;

      elsif ( x63 and not x17 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x17 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x17 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and not x17 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x17 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x67 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and x64 and x67 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x63 and x64 and x67 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x67 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x67 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s108;

      else
         y38 <= '1' ;
         current_otherm <= s483;

      end if;

   when s412 =>
      if ( x63 and x66 and x23 and x25 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s582;

      elsif ( x63 and x66 and x23 and not x25 and x5 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x63 and x66 and x23 and not x25 and not x5 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s582;

      elsif ( x63 and x66 and not x23 and x5 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x63 and x66 and not x23 and x5 and not x24 ) = '1' then
         y60 <= '1' ;
         current_otherm <= s190;

      elsif ( x63 and x66 and not x23 and not x5 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s455;

      elsif ( x63 and not x66 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and not x66 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x64 and x66 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x64 and x66 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x66 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x66 ) = '1' then
         current_otherm <= s1;

      else
         y57 <= '1' ;
         current_otherm <= s582;

      end if;

   when s413 =>
      if ( x63 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y39 <= '1' ;
         current_otherm <= s726;

      end if;

   when s414 =>
      if ( x63 and x20 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s727;

      elsif ( x63 and not x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      else
         y6 <= '1' ;
         current_otherm <= s337;

      end if;

   when s415 =>
      if ( x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x64 and x4 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1;

      elsif ( not x64 and not x4 and x31 and x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s398;

      elsif ( not x64 and not x4 and x31 and not x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s310;

      elsif ( not x64 and not x4 and not x31 and x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s352;

      else
         y5 <= '1' ;
         current_otherm <= s366;

      end if;

   when s416 =>
      if ( x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x64 and x66 and x4 ) = '1' then
         y29 <= '1' ;
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y67 <= '1' ;
         current_otherm <= s728;

      elsif ( not x64 and x66 and not x4 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s268;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y69 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s729;

      end if;

   when s417 =>
      if ( x21 and x20 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x21 and x20 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x21 and x20 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and x20 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x20 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( x21 and not x20 and x6 and not x7 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( x21 and not x20 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x20 and not x6 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s418 =>
         y8 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s730;

   when s419 =>
      if ( x12 and x13 and x3 ) = '1' then
         y3 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s420;

      elsif ( x12 and x13 and not x3 and x14 ) = '1' then
         y3 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s420;

      elsif ( x12 and x13 and not x3 and not x14 ) = '1' then
         y10 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s421;

      elsif ( x12 and not x13 ) = '1' then
         y3 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s422;

      else
         y10 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s423;

      end if;

   when s420 =>
         y11 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s461;

   when s421 =>
      if ( x13 ) = '1' then
         y19 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s1;

      else
         y20 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1;

      end if;

   when s422 =>
      if ( x14 ) = '1' then
         y3 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s420;

      else
         y10 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s421;

      end if;

   when s423 =>
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

   when s424 =>
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s731;

   when s425 =>
      if ( x64 and x65 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x64 and not x65 ) = '1' then
         y5 <= '1' ;
         y13 <= '1' ;
         y30 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s732;

      elsif ( not x64 and x65 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x65 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x65 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x65 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x64 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x64 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s426 =>
      if ( x63 and x20 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s733;

      elsif ( x63 and not x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s397;

      else
         y33 <= '1' ;
         current_otherm <= s321;

      end if;

   when s427 =>
         y6 <= '1' ;
         current_otherm <= s239;

   when s428 =>
      if ( x63 ) = '1' then
         y25 <= '1' ;
         y27 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s734;

      else
         y48 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s735;

      end if;

   when s429 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s736;

   when s430 =>
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s384;

   when s431 =>
      if ( x66 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s737;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s736;

      end if;

   when s432 =>
      if ( x63 and x16 and x22 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( x63 and x16 and not x22 and x23 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( x63 and x16 and not x22 and not x23 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( x63 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s738;

      elsif ( not x63 and x64 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s739;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s740;

      end if;

   when s433 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s429;

   when s434 =>
      if ( x63 and x17 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x17 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x17 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x17 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s741;

      elsif ( not x63 and x65 and x3 and x6 and x5 and x9 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( not x63 and x65 and x3 and x6 and x5 and x9 and not x7 and x8 and x17 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x63 and x65 and x3 and x6 and x5 and x9 and not x7 and x8 and not x17 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x3 and x6 and x5 and x9 and not x7 and x8 and not x17 and x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x65 and x3 and x6 and x5 and x9 and not x7 and x8 and not x17 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x65 and x3 and x6 and x5 and x9 and not x7 and not x8 ) = '1' then
         y5 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and x7 ) = '1' then
         y68 <= '1' ;
         current_otherm <= s743;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and not x7 and x8 and x18 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and not x7 and x8 and not x18 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and not x7 and x8 and not x18 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and not x7 and x8 and not x18 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and not x7 and x8 and not x18 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x65 and x3 and x6 and x5 and not x9 and not x7 and not x8 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s744;

      elsif ( not x63 and x65 and x3 and x6 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s745;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and x8 and x7 and x9 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and x8 and x7 and not x9 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and x8 and not x7 and x11 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s746;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and x8 and not x7 and x11 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and x8 and not x7 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s747;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and not x8 and x9 and x7 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and not x8 and x9 and not x7 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and not x8 and x9 and not x7 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s747;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and not x8 and not x9 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and x65 and x3 and not x6 and x5 and not x8 and not x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s748;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and x8 and x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and x8 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s749;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and x8 and not x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and not x8 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s750;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and not x8 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y40 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s751;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and x11 and not x8 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x63 and x65 and x3 and not x6 and not x5 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s752;

      elsif ( not x63 and x65 and not x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s753;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and x4 and x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and x4 and not x6 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and x6 and x9 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and x6 and not x9 and x17 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and x6 and not x9 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and not x6 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and not x6 and not x8 and x17 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and x5 and not x6 and not x8 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s585;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and x20 and not x4 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y40 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s585;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and x6 and x4 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and x6 and not x4 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and x6 and not x4 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and x6 and not x4 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and x6 and not x4 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and x6 and not x4 and not x13 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and not x6 and x4 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s719;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and not x6 and not x4 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and not x6 and not x4 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and not x6 and not x4 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and not x6 and not x4 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and x5 and not x6 and not x4 and not x14 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and x6 and x4 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and x6 and x4 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and x6 and x4 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and x6 and x4 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and x6 and x4 and not x11 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and x6 and not x4 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and not x6 and x4 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and not x6 and x4 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and not x6 and x4 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and not x6 and x4 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and not x6 and x4 and not x10 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and x18 and not x5 and not x6 and not x4 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x63 and not x65 and x67 and x15 and x21 and not x20 and not x18 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s754;

      elsif ( not x63 and not x65 and x67 and x15 and not x21 and x18 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s585;

      elsif ( not x63 and not x65 and x67 and x15 and not x21 and x18 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s745;

      elsif ( not x63 and not x65 and x67 and x15 and not x21 and x18 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y10 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s755;

      elsif ( not x63 and not x65 and x67 and x15 and not x21 and x18 and not x20 and x4 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x63 and not x65 and x67 and x15 and not x21 and x18 and not x20 and not x4 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x63 and not x65 and x67 and x15 and not x21 and not x18 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s754;

      elsif ( not x63 and not x65 and x67 and not x15 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s283;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and x21 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and x21 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y34 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and x10 and x24 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and x10 and not x24 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and x10 and not x24 and x26 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and x10 and not x24 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and not x10 and x25 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and not x10 and not x25 and x26 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and not x10 and not x25 and x26 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and x22 and not x10 and not x25 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and not x22 and x23 and x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and not x22 and x23 and not x10 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and not x22 and not x23 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and not x22 and not x23 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and not x22 and not x23 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and x5 and not x21 and not x22 and not x23 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and x8 and x14 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and x8 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and x10 and x11 and x14 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and x10 and x11 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and x10 and not x11 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and x10 and not x11 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and x10 and not x11 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and x10 and not x11 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and not x10 and x12 and x14 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and not x10 and x12 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and x10 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s757;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and x10 and not x8 and x14 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and x10 and not x8 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and x8 and x13 and x14 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and x8 and x13 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and not x67 and x3 and x6 and not x5 and not x9 and not x10 and not x8 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and x5 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and x5 and not x7 and x8 ) = '1' then
         y5 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and x5 and not x7 and not x8 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and x5 and not x7 and not x8 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and not x5 and x8 ) = '1' then
         y5 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and not x5 and not x8 and x14 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s756;

      elsif ( not x63 and not x65 and not x67 and x3 and not x6 and not x5 and not x8 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      else
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s758;

      end if;

   when s435 =>
         y9 <= '1' ;
         current_otherm <= s759;

   when s436 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s760;

   when s437 =>
      if ( x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s143;

      elsif ( not x33 and x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s143;

      elsif ( not x33 and not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x33 and not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x33 and not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s438 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s147;

   when s439 =>
      if ( x32 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s138;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      end if;

   when s440 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s761;

   when s441 =>
         y42 <= '1' ;
         current_otherm <= s762;

   when s442 =>
      if ( x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s136;

      elsif ( not x33 and x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s136;

      elsif ( not x33 and not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x33 and not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x33 and not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s443 =>
      if ( x32 and x33 ) = '1' then
         y3 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s49;

      elsif ( x32 and not x33 and x14 and x15 and x13 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( x32 and not x33 and x14 and x15 and not x13 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s145;

      elsif ( x32 and not x33 and x14 and not x15 and x13 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s142;

      elsif ( x32 and not x33 and x14 and not x15 and not x13 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s147;

      elsif ( x32 and not x33 and not x14 and x15 and x13 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s140;

      elsif ( x32 and not x33 and not x14 and x15 and x13 and not x16 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s141;

      elsif ( x32 and not x33 and not x14 and x15 and not x13 and x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x33 and not x14 and x15 and not x13 and not x17 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s146;

      elsif ( x32 and not x33 and not x14 and not x15 and x13 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s143;

      elsif ( x32 and not x33 and not x14 and not x15 and not x13 and x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x33 and not x14 and not x15 and not x13 and not x18 ) = '1' then
         current_otherm <= s443;

      elsif ( not x32 and x13 and x33 and x15 and x14 and x5 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( not x32 and x13 and x33 and x15 and x14 and not x5 and x7 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( not x32 and x13 and x33 and x15 and x14 and not x5 and not x7 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s132;

      elsif ( not x32 and x13 and x33 and x15 and not x14 and x31 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( not x32 and x13 and x33 and x15 and not x14 and x31 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x32 and x13 and x33 and x15 and not x14 and not x31 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x13 and x33 and x15 and not x14 and not x31 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x13 and x33 and x15 and not x14 and not x31 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x13 and x33 and x15 and not x14 and not x31 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x13 and x33 and not x15 and x14 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s136;

      elsif ( not x32 and x13 and x33 and not x15 and x14 and not x5 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( not x32 and x13 and x33 and not x15 and not x14 and x16 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( not x32 and x13 and x33 and not x15 and not x14 and x16 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x32 and x13 and x33 and not x15 and not x14 and not x16 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x13 and x33 and not x15 and not x14 and not x16 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x13 and x33 and not x15 and not x14 and not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x13 and x33 and not x15 and not x14 and not x16 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and x13 and not x33 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s144;

      elsif ( not x32 and not x13 and x33 and x14 and x15 and x8 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( not x32 and not x13 and x33 and x14 and x15 and x8 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and not x13 and x33 and x14 and x15 and not x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and not x13 and x33 and x14 and not x15 and x30 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( not x32 and not x13 and x33 and x14 and not x15 and x30 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and not x13 and x33 and x14 and not x15 and not x30 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x32 and not x13 and x33 and not x14 and x15 and x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( not x32 and not x13 and x33 and not x14 and x15 and not x5 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x32 and not x13 and x33 and not x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s138;

      elsif ( not x32 and not x13 and not x33 and x4 and x6 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s148;

      elsif ( not x32 and not x13 and not x33 and x4 and not x6 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      else
         y15 <= '1' ;
         current_otherm <= s149;

      end if;

   when s444 =>
      if ( x32 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s763;

      else
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s144;

      end if;

   when s445 =>
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s764;

   when s446 =>
      if ( x32 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s132;

      elsif ( not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s447 =>
         y53 <= '1' ;
         current_otherm <= s394;

   when s448 =>
      if ( x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x32 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s765;

      end if;

   when s449 =>
      if ( x32 ) = '1' then
         y31 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s138;

      elsif ( not x32 and x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s766;

      elsif ( not x32 and not x33 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x33 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and not x33 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s450 =>
         y8 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s767;

   when s451 =>
      if ( x16 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s395;

      elsif ( not x16 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x16 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s452 =>
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s768;

   when s453 =>
         y26 <= '1' ;
         current_otherm <= s116;

   when s454 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s769;

   when s455 =>
      if ( x62 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s770;

      elsif ( not x62 and x11 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      else
         y49 <= '1' ;
         current_otherm <= s256;

      end if;

   when s456 =>
         y52 <= '1' ;
         current_otherm <= s360;

   when s457 =>
      if ( x27 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      else
         y69 <= '1' ;
         y73 <= '1' ;
         current_otherm <= s563;

      end if;

   when s458 =>
         y2 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s613;

   when s459 =>
      if ( x62 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s459;

      elsif ( x62 and x9 and not x10 and x8 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s771;

      elsif ( x62 and x9 and not x10 and not x8 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s772;

      elsif ( x62 and not x9 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s773;

      elsif ( not x62 and x65 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s460 =>
      if ( x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s461 =>
         y12 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s530;

   when s462 =>
      if ( x11 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s459;

      elsif ( not x11 and x22 and x9 and x8 and x23 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x11 and x22 and x9 and x8 and x23 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x11 and x22 and x9 and x8 and x23 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x22 and x9 and x8 and x23 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x11 and x22 and x9 and x8 and x23 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x22 and x9 and x8 and not x23 and x10 ) = '1' then
         y62 <= '1' ;
         current_otherm <= s525;

      elsif ( not x11 and x22 and x9 and x8 and not x23 and not x10 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and x10 and x5 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and x10 and not x5 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and x10 and not x5 and x6 and not x4 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and x10 and not x5 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and not x10 and x4 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and not x10 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x11 and x22 and x9 and not x8 and x23 and not x10 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x22 and x9 and not x8 and not x23 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y38 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and x22 and x9 and not x8 and not x23 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y36 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and x22 and not x9 and x10 and x23 and x8 ) = '1' then
         y33 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s1;

      elsif ( not x11 and x22 and not x9 and x10 and x23 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y51 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and x22 and not x9 and x10 and not x23 and x8 ) = '1' then
         y60 <= '1' ;
         current_otherm <= s190;

      elsif ( not x11 and x22 and not x9 and x10 and not x23 and not x8 ) = '1' then
         y58 <= '1' ;
         current_otherm <= s774;

      elsif ( not x11 and x22 and not x9 and not x10 and x23 and x8 ) = '1' then
         y37 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s1;

      elsif ( not x11 and x22 and not x9 and not x10 and x23 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y52 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and x22 and not x9 and not x10 and not x23 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s775;

      elsif ( not x11 and x22 and not x9 and not x10 and not x23 and not x8 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s577;

      elsif ( not x11 and not x22 and x23 and x21 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( not x11 and not x22 and x23 and not x21 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s776;

      elsif ( not x11 and not x22 and not x23 and x9 and x10 and x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and not x22 and not x23 and x9 and x10 and not x8 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and not x22 and not x23 and x9 and not x10 and x8 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x11 and not x22 and not x23 and x9 and not x10 and not x8 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s250;

      elsif ( not x11 and not x22 and not x23 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s542;

      else
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s250;

      end if;

   when s463 =>
      if ( x63 and x12 and x22 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s346;

      elsif ( x63 and x12 and not x22 and x23 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x63 and x12 and not x22 and not x23 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x63 and not x12 and x7 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s557;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and x9 and x23 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and x9 and x23 and not x10 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and x9 and not x23 and x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and x9 and not x23 and not x10 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and x10 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and x10 and not x13 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and x10 and not x13 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and x10 and not x13 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and x10 and not x13 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and x10 and not x13 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and not x10 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and not x10 and not x1 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and not x10 and not x1 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and not x10 and not x1 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and not x10 and not x1 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and x23 and not x10 and not x1 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and x8 and not x9 and not x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s542;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and x9 and x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and x9 and not x23 and x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and x9 and not x23 and not x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and x10 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and x10 and not x3 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and x10 and not x3 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and x10 and not x3 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and x10 and not x3 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and x10 and not x3 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and not x10 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and not x10 and not x15 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and x23 and not x10 and not x15 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x12 and x7 and not x22 and not x8 and not x9 and not x23 ) = '1' then
         y5 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( x63 and not x12 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s251;

      elsif ( not x63 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s777;

      elsif ( not x63 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s778;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      end if;

   when s464 =>
      if ( x64 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s191;

      else
         y47 <= '1' ;
         y57 <= '1' ;
         y61 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s779;

      end if;

   when s465 =>
      if ( x63 and x10 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x10 and not x2 and x3 and x4 and x5 and x1 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x10 and not x2 and x3 and x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and x3 and x4 and not x5 and x1 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x63 and x10 and not x2 and x3 and x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and x3 and not x4 and x5 and x1 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x63 and x10 and not x2 and x3 and not x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and x3 and not x4 and not x5 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and x3 and not x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and x5 and x1 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and x5 and x1 and not x6 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s340;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and not x5 and x1 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and not x5 and x1 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and not x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and not x3 and x4 and not x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and not x3 and not x4 and x1 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and not x3 and not x4 and x1 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and x10 and not x2 and not x3 and not x4 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y32 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x63 and not x10 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s780;

      elsif ( not x63 and x67 and x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and x67 and x11 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x63 and x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x67 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         y38 <= '1' ;
         current_otherm <= s261;

      end if;

   when s466 =>
      if ( x64 and x21 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s95;

      elsif ( x64 and x21 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s781;

      elsif ( x64 and not x21 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s594;

      elsif ( x64 and not x21 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s782;

      else
         y48 <= '1' ;
         y57 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s453;

      end if;

   when s467 =>
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s676;

   when s468 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s783;

   when s469 =>
         y15 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s784;

   when s470 =>
      if ( x63 and x64 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s785;

      elsif ( x63 and not x64 and x9 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s320;

      elsif ( x63 and not x64 and not x9 ) = '1' then
         current_otherm <= s470;

      else
         y27 <= '1' ;
         current_otherm <= s335;

      end if;

   when s471 =>
      if ( x20 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s786;

      elsif ( not x20 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s472 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s787;

   when s473 =>
      if ( x11 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s788;

      else
         y67 <= '1' ;
         current_otherm <= s584;

      end if;

   when s474 =>
         y14 <= '1' ;
         current_otherm <= s201;

   when s475 =>
      if ( x62 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s287;

      elsif ( not x62 and x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      else
         y7 <= '1' ;
         current_otherm <= s90;

      end if;

   when s476 =>
      if ( x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s466;

      else
         y7 <= '1' ;
         current_otherm <= s789;

      end if;

   when s477 =>
      if ( x6 and x12 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s790;

      elsif ( x6 and not x12 and x11 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s410;

      elsif ( x6 and not x12 and not x11 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x6 and not x12 and not x11 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x6 and not x12 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x12 and not x11 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and x11 and x12 and x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and x11 and x12 and x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and x11 and x12 and x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and x11 and x12 and x10 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and x11 and x12 and not x10 and x16 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and x11 and x12 and not x10 and not x16 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and x11 and not x12 and x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s791;

      elsif ( not x6 and x8 and x11 and not x12 and not x10 and x17 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and x11 and not x12 and not x10 and not x17 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and not x11 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s792;

      elsif ( not x6 and x8 and not x11 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x6 and x8 and not x11 and not x12 and x10 and x15 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and not x11 and not x12 and x10 and not x15 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x8 and not x11 and not x12 and not x10 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s790;

      end if;

   when s478 =>
      if ( x62 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x62 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x63 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x62 and x63 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and not x63 and x64 and x66 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x62 and not x63 and x64 and x66 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x66 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x62 and not x63 and x64 and not x66 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x66 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 ) = '1' then
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s793;

      elsif ( not x62 and not x63 and not x64 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x63 and not x64 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x62 and not x63 and not x64 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s479 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s794;

   when s480 =>
      if ( x11 and x12 and x10 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( x11 and x12 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( x11 and not x12 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( x11 and not x12 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x11 and x12 and x10 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s409;

      elsif ( not x11 and x12 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x11 and not x12 and x10 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x11 and not x12 and not x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x11 and not x12 and not x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x11 and not x12 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s481 =>
      if ( x7 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      else
         y10 <= '1' ;
         current_otherm <= s16;

      end if;

   when s482 =>
         y5 <= '1' ;
         current_otherm <= s359;

   when s483 =>
      if ( x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x67 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x67 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x62 and x63 and x67 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and x67 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x67 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x63 and not x67 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x63 and not x67 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x63 and not x67 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x62 and not x63 and x64 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and x64 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and x65 and x31 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s99;

      elsif ( not x62 and not x63 and not x64 and x65 and not x31 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s355;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and x6 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and x6 and not x5 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and x8 and x9 and x5 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s153;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and x8 and x9 and not x5 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y62 <= '1' ;
         y63 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and x8 and x9 and not x5 and not x7 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y57 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and x8 and not x9 and x5 ) = '1' then
         y3 <= '1' ;
         y19 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and x8 and not x9 and not x5 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y67 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and x8 and not x9 and not x5 and not x7 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y55 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and not x8 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and not x8 and not x5 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y62 <= '1' ;
         y63 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and not x8 and not x5 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and x19 and not x6 and not x8 and not x5 and not x7 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y41 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s795;

      elsif ( not x62 and not x63 and not x64 and not x65 and x66 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s796;

      elsif ( not x62 and not x63 and not x64 and not x65 and not x66 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x65 and not x66 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x62 and not x63 and not x64 and not x65 and not x66 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s484 =>
         y5 <= '1' ;
         current_otherm <= s366;

   when s485 =>
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s797;

   when s486 =>
      if ( x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s346;

      elsif ( not x64 and x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      else
         y5 <= '1' ;
         current_otherm <= s398;

      end if;

   when s487 =>
      if ( x30 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s714;

      else
         y24 <= '1' ;
         current_otherm <= s203;

      end if;

   when s488 =>
      if ( x63 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s798;

      elsif ( not x63 and x64 and x21 and x10 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s74;

      elsif ( not x63 and x64 and x21 and not x10 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s363;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and x17 and x16 and x19 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and x17 and x16 and x19 and not x11 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and x17 and x16 and not x19 and x18 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and x17 and x16 and not x19 and not x18 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and x17 and not x16 and x11 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and x17 and not x16 and not x11 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s365;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and not x17 and x16 and x19 and x14 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and not x17 and x16 and x19 and not x14 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and not x17 and x16 and not x19 and x13 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and not x17 and x16 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x64 and x21 and not x10 and not x12 and not x17 and not x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x64 and not x21 and x6 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s398;

      elsif ( not x63 and x64 and not x21 and not x6 and x5 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s185;

      elsif ( not x63 and x64 and not x21 and not x6 and not x5 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s363;

      else
         y42 <= '1' ;
         current_otherm <= s762;

      end if;

   when s489 =>
      if ( x17 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s799;

      else
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s489;

      end if;

   when s490 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y12 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s444;

   when s491 =>
      if ( x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s247;

      else
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s248;

      end if;

   when s492 =>
      if ( x16 and x22 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x16 and x22 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x16 and x22 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x16 and x22 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x16 and x22 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x16 and not x22 ) = '1' then
         y3 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      else
         y3 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s249;

      end if;

   when s493 =>
      if ( x22 ) = '1' then
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s187;

      elsif ( not x22 and x23 ) = '1' then
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s187;

      else
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s800;

      end if;

   when s494 =>
      if ( x22 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s800;

      elsif ( not x22 and x23 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s800;

      else
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s187;

      end if;

   when s495 =>
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s801;

   when s496 =>
      if ( x22 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s802;

      else
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s801;

      end if;

   when s497 =>
      if ( x22 and x16 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x22 and x16 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x22 and x16 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x22 and x16 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x22 and x16 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x22 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s344;

      elsif ( not x22 and x16 and x7 and x8 and x9 and x23 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( not x22 and x16 and x7 and x8 and x9 and x23 and not x10 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( not x22 and x16 and x7 and x8 and x9 and not x23 and x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and x8 and x9 and not x23 and not x10 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and x10 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and x10 and not x13 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and x10 and not x13 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and x10 and not x13 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and x10 and not x13 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and x10 and not x13 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and not x10 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and not x10 and not x1 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and not x10 and not x1 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and not x10 and not x1 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and not x10 and not x1 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and x23 and not x10 and not x1 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and x8 and not x9 and not x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s542;

      elsif ( not x22 and x16 and x7 and not x8 and x9 and x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and not x8 and x9 and not x23 and x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and not x8 and x9 and not x23 and not x10 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and x10 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and x10 and not x3 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and x10 and not x3 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and x10 and not x3 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and x10 and not x3 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and x10 and not x3 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and not x10 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and not x10 and not x15 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and not x10 and not x15 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and x23 and not x10 and not x15 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x22 and x16 and x7 and not x8 and not x9 and not x23 ) = '1' then
         y5 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s250;

      elsif ( not x22 and x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s251;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s252;

      end if;

   when s498 =>
      if ( x63 and x65 and x20 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x63 and x65 and not x20 ) = '1' then
         y62 <= '1' ;
         current_otherm <= s524;

      elsif ( x63 and not x65 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x65 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x65 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and x10 ) = '1' then
         y62 <= '1' ;
         current_otherm <= s524;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and x3 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and x3 and x12 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and x3 and x12 and not x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and x3 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and x6 and x7 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and x6 and not x7 and x12 and x8 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and x6 and not x7 and x12 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and x6 and not x7 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and not x6 and x8 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and not x6 and not x8 and x12 and x7 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and not x6 and not x8 and x12 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and x5 and not x3 and not x6 and not x8 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and not x5 and x6 and x3 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and not x5 and x6 and not x3 ) = '1' then
         y21 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s180;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and not x5 and not x6 and x3 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x63 and x64 and x65 and not x10 and x4 and not x5 and not x6 and not x3 ) = '1' then
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s180;

      elsif ( not x63 and x64 and x65 and not x10 and not x4 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x64 and not x65 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      elsif ( not x63 and not x64 and x65 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and not x64 and x65 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and not x64 and x65 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x65 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x65 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and not x64 and not x65 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and not x64 and not x65 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s499 =>
      if ( x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s308;

      else
         y4 <= '1' ;
         y62 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s614;

      end if;

   when s500 =>
      if ( x21 and x20 ) = '1' then
         y13 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1;

      elsif ( x21 and not x20 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x21 and not x20 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x21 and not x20 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x20 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y13 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1;

      end if;

   when s501 =>
      if ( x31 and x30 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s803;

      elsif ( x31 and not x30 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s781;

      else
         y30 <= '1' ;
         current_otherm <= s803;

      end if;

   when s502 =>
      if ( x63 and x19 and x18 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s804;

      elsif ( x63 and x19 and not x18 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s560;

      elsif ( x63 and not x19 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s655;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s805;

      end if;

   when s503 =>
         y8 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s804;

   when s504 =>
      if ( x63 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s806;

      elsif ( x63 and x19 and not x18 ) = '1' then
         y25 <= '1' ;
         y28 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s807;

      elsif ( x63 and not x19 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s804;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s808;

      end if;

   when s505 =>
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s71;

   when s506 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

   when s507 =>
         y21 <= '1' ;
         current_otherm <= s172;

   when s508 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x64 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x64 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x64 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and not x64 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and not x64 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x64 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s509 =>
      if ( x64 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s201;

      elsif ( x64 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s809;

      else
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s810;

      end if;

   when s510 =>
      if ( x63 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s560;

      elsif ( not x63 and x30 ) = '1' then
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s811;

      elsif ( not x63 and not x30 and x31 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s183;

      else
         y31 <= '1' ;
         current_otherm <= s486;

      end if;

   when s511 =>
         y25 <= '1' ;
         current_otherm <= s363;

   when s512 =>
      if ( x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s513 =>
      if ( x62 and x20 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s595;

      elsif ( x62 and not x20 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s644;

      elsif ( not x62 and x20 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s813;

      end if;

   when s514 =>
         y27 <= '1' ;
         current_otherm <= s385;

   when s515 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s814;

   when s516 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s815;

   when s517 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s816;

   when s518 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s817;

   when s519 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s818;

   when s520 =>
         y57 <= '1' ;
         current_otherm <= s135;

   when s521 =>
      if ( x62 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x62 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x64 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x62 and x64 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x64 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x64 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and not x64 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x62 and not x64 and x19 and not x14 and not x13 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x62 and not x64 and x19 and not x14 and not x13 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x62 and not x64 and x19 and not x14 and not x13 and not x11 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      else
         current_otherm <= s1;

      end if;

   when s522 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s819;

   when s523 =>
      if ( x3 and x4 and x5 and x21 and x7 and x9 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x3 and x4 and x5 and x21 and x7 and not x9 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and x9 and x12 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and x9 and not x12 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and x9 and not x12 and x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and x9 and not x12 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and not x9 and x11 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and not x9 and not x11 and x10 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and not x9 and not x11 and x10 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x5 and x21 and not x7 and x8 and not x9 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x5 and x21 and not x7 and not x8 and x9 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s820;

      elsif ( x3 and x4 and x5 and x21 and not x7 and not x8 and not x9 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y16 <= '1' ;
         y42 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s820;

      elsif ( x3 and x4 and x5 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s821;

      elsif ( x3 and x4 and not x5 and x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s822;

      elsif ( x3 and x4 and not x5 and not x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s821;

      elsif ( x3 and not x4 ) = '1' then
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s823;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s824;

      end if;

   when s524 =>
      if ( x63 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x63 and not x18 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      else
         y2 <= '1' ;
         current_otherm <= s24;

      end if;

   when s525 =>
      if ( x63 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         y63 <= '1' ;
         current_otherm <= s224;

      end if;

   when s526 =>
      if ( x18 and x19 and x14 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( x18 and x19 and not x14 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x19 and not x14 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x19 and not x14 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x19 and not x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x18 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x18 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x18 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s527 =>
         y30 <= '1' ;
         current_otherm <= s121;

   when s528 =>
         y2 <= '1' ;
         current_otherm <= s24;

   when s529 =>
         y1 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s655;

   when s530 =>
      if ( x64 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      elsif ( x64 and not x15 and x14 and x13 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

      elsif ( x64 and not x15 and x14 and not x13 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s211;

      elsif ( x64 and not x15 and not x14 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s347;

      elsif ( not x64 and x14 and x13 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x13 and x66 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x13 and not x66 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x64 and not x14 and x66 ) = '1' then
         y19 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s1;

      else
         y12 <= '1' ;
         current_otherm <= s176;

      end if;

   when s531 =>
      if ( x18 and x26 and x14 and x27 and x6 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s826;

      elsif ( x18 and x26 and x14 and x27 and x6 and not x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( x18 and x26 and x14 and x27 and not x6 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s825;

      elsif ( x18 and x26 and x14 and x27 and not x6 and not x5 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s583;

      elsif ( x18 and x26 and x14 and not x27 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s579;

      elsif ( x18 and x26 and x14 and not x27 and not x5 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s583;

      elsif ( x18 and x26 and not x14 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s826;

      elsif ( x18 and x26 and not x14 and not x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( x18 and not x26 and x27 and x14 and x5 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( x18 and not x26 and x27 and x14 and not x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s825;

      elsif ( x18 and not x26 and x27 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s826;

      elsif ( x18 and not x26 and not x27 and x7 and x6 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x18 and not x26 and not x27 and x7 and x6 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x18 and not x26 and not x27 and x7 and x6 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and x6 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and x6 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and x8 and x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s556;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and not x8 and x16 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s556;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x26 and not x27 and not x7 and x8 and x6 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x18 and not x26 and not x27 and not x7 and x8 and not x6 ) = '1' then
         y5 <= '1' ;
         y44 <= '1' ;
         y55 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s579;

      elsif ( x18 and not x26 and not x27 and not x7 and not x8 and x6 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x18 and not x26 and not x27 and not x7 and not x8 and not x6 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y53 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s579;

      else
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s827;

      end if;

   when s532 =>
      if ( x62 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s828;

      else
         y28 <= '1' ;
         current_otherm <= s780;

      end if;

   when s533 =>
         y13 <= '1' ;
         current_otherm <= s225;

   when s534 =>
      if ( x64 and x14 and x10 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and x14 and not x10 and x11 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x64 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x31 and x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      elsif ( not x64 and x31 and not x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s667;

      elsif ( not x64 and not x31 and x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s146;

      else
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s501;

      end if;

   when s535 =>
      if ( x63 and x26 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( x63 and not x26 ) = '1' then
         y66 <= '1' ;
         current_otherm <= s473;

      elsif ( not x63 and x65 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x65 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x65 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x65 and x20 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      else
         current_otherm <= s1;

      end if;

   when s536 =>
      if ( x62 and x10 and x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x10 and not x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( x62 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x17 and x18 and x5 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s536;

      elsif ( not x62 and x17 and x18 and not x5 and x6 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      elsif ( not x62 and x17 and x18 and not x5 and not x6 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s35;

      elsif ( not x62 and x17 and not x18 and x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s37;

      elsif ( not x62 and x17 and not x18 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s36;

      elsif ( not x62 and not x17 and x18 and x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and not x17 and x18 and not x1 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s33;

      else
         current_otherm <= s1;

      end if;

   when s537 =>
         y6 <= '1' ;
         current_otherm <= s336;

   when s538 =>
         y27 <= '1' ;
         current_otherm <= s488;

   when s539 =>
         y5 <= '1' ;
         current_otherm <= s310;

   when s540 =>
         y13 <= '1' ;
         current_otherm <= s238;

   when s541 =>
         y10 <= '1' ;
         current_otherm <= s559;

   when s542 =>
      if ( x63 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s829;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s742;

      end if;

   when s543 =>
      if ( x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s331;

      elsif ( not x3 and x21 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s639;

      else
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s640;

      end if;

   when s544 =>
      if ( x21 and x3 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y79 <= '1' ;
         current_otherm <= s830;

      elsif ( x21 and not x3 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y71 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s830;

      elsif ( not x21 and x22 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s366;

      elsif ( not x21 and x22 and not x3 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s639;

      elsif ( not x21 and not x22 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      else
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s319;

      end if;

   when s545 =>
      if ( x21 and x3 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y96 <= '1' ;
         current_otherm <= s710;

      elsif ( x21 and not x3 ) = '1' then
         y60 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y79 <= '1' ;
         current_otherm <= s710;

      elsif ( not x21 and x22 and x3 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s711;

      elsif ( not x21 and x22 and not x3 ) = '1' then
         y62 <= '1' ;
         y81 <= '1' ;
         current_otherm <= s711;

      elsif ( not x21 and not x22 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s359;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s639;

      end if;

   when s546 =>
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s393;

   when s547 =>
      if ( x21 and x3 ) = '1' then
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s831;

      elsif ( x21 and not x3 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y79 <= '1' ;
         y88 <= '1' ;
         y102 <= '1' ;
         current_otherm <= s831;

      elsif ( not x21 and x3 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y96 <= '1' ;
         current_otherm <= s710;

      else
         y60 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y79 <= '1' ;
         current_otherm <= s710;

      end if;

   when s548 =>
      if ( x21 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s366;

      elsif ( x21 and not x3 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y93 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x22 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s359;

      elsif ( not x21 and x22 and not x3 ) = '1' then
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s640;

      elsif ( not x21 and not x22 and x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s366;

      else
         y4 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         current_otherm <= s673;

      end if;

   when s549 =>
      if ( x3 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s68;

      else
         y4 <= '1' ;
         y62 <= '1' ;
         y73 <= '1' ;
         current_otherm <= s832;

      end if;

   when s550 =>
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s544;

   when s551 =>
      if ( x21 and x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s546;

      elsif ( x21 and not x10 and x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s544;

      elsif ( x21 and not x10 and x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s547;

      elsif ( x21 and not x10 and not x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( x21 and not x10 and not x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s549;

      elsif ( not x21 and x22 and x10 and x11 and x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( not x21 and x22 and x10 and x11 and not x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s545;

      elsif ( not x21 and x22 and x10 and not x11 and x14 and x19 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x22 and x10 and not x11 and x14 and not x19 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and x10 and not x11 and x14 and not x19 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and x10 and not x11 and x14 and not x19 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and x10 and not x11 and x14 and not x19 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and x10 and not x11 and not x14 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x22 and x10 and not x11 and not x14 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and x10 and not x11 and not x14 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and x10 and not x11 and not x14 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and x10 and not x11 and not x14 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and x14 and x11 and x17 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x22 and not x10 and x14 and x11 and not x17 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x10 and x14 and x11 and not x17 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x10 and x14 and x11 and not x17 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and x14 and x11 and not x17 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and x14 and not x11 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and x16 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and x16 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and x16 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and x16 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and x16 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and not x16 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and not x16 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and not x16 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and not x14 and x11 and not x16 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x10 and not x14 and not x11 ) = '1' then
         y102 <= '1' ;
         current_otherm <= s240;

      else
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      end if;

   when s552 =>
      if ( x21 and x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s546;

      elsif ( x21 and not x10 and x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s544;

      elsif ( x21 and not x10 and x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s547;

      elsif ( x21 and not x10 and not x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( x21 and not x10 and not x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s549;

      elsif ( not x21 and x10 and x22 and x11 and x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( not x21 and x10 and x22 and x11 and not x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s545;

      elsif ( not x21 and x10 and x22 and not x11 and x14 and x19 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x10 and x22 and not x11 and x14 and not x19 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x10 and x22 and not x11 and not x14 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x10 and x22 and not x11 and not x14 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x10 and not x22 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s550;

      elsif ( not x21 and not x10 and x22 and x14 and x11 and x17 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x10 and x22 and x14 and x11 and not x17 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x10 and x22 and x14 and not x11 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and x16 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x10 and x22 and not x14 and x11 and not x16 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x10 and x22 and not x14 and not x11 ) = '1' then
         y102 <= '1' ;
         current_otherm <= s240;

      else
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s551;

      end if;

   when s553 =>
      if ( x15 ) = '1' then
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s240;

      elsif ( not x15 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s554 =>
      if ( x63 and x28 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x63 and not x28 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x15 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      elsif ( not x63 and not x15 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x15 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x63 and not x15 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s555 =>
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s543;

   when s556 =>
      if ( x63 and x23 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s664;

      elsif ( x63 and x23 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s187;

      elsif ( x63 and not x23 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s187;

      elsif ( x63 and not x23 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s188;

      elsif ( not x63 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x63 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s557 =>
      if ( x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s833;

      elsif ( not x8 and x10 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s834;

      elsif ( not x8 and x10 and not x9 ) = '1' then
         y58 <= '1' ;
         current_otherm <= s774;

      elsif ( not x8 and not x10 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s835;

      else
         y56 <= '1' ;
         current_otherm <= s577;

      end if;

   when s558 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s836;

   when s559 =>
      if ( x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s837;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s836;

      end if;

   when s560 =>
      if ( x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s561 =>
      if ( x19 and x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s392;

      elsif ( x19 and not x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s838;

      else
         y2 <= '1' ;
         current_otherm <= s392;

      end if;

   when s562 =>
      if ( x64 and x63 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x64 and x63 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x64 and x63 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and x63 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and x65 ) = '1' then
         y4 <= '1' ;
         y20 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s396;

      elsif ( x64 and not x63 and not x65 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x64 and not x63 and not x65 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x64 and not x63 and not x65 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x63 and not x65 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x63 and x66 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x64 and x63 and x66 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x64 and x63 and x66 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x63 and x66 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x63 and not x66 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x64 and x63 and not x66 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x64 and x63 and not x66 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x63 and not x66 and not x1 ) = '1' then
         current_otherm <= s1;

      else
         y25 <= '1' ;
         current_otherm <= s363;

      end if;

   when s563 =>
      if ( x26 ) = '1' then
         y74 <= '1' ;
         current_otherm <= s554;

      elsif ( not x26 and x27 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s262;

      else
         y69 <= '1' ;
         y73 <= '1' ;
         current_otherm <= s563;

      end if;

   when s564 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s125;

   when s565 =>
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s839;

   when s566 =>
         y13 <= '1' ;
         current_otherm <= s375;

   when s567 =>
      if ( x49 and x50 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x49 and not x50 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s315;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

      end if;

   when s568 =>
      if ( x64 and x3 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s289;

      elsif ( x64 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s840;

      else
         y39 <= '1' ;
         current_otherm <= s726;

      end if;

   when s569 =>
      if ( x64 and x3 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x64 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s598;

      else
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s793;

      end if;

   when s570 =>
      if ( x64 and x3 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s594;

      elsif ( x64 and not x3 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s841;

      else
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s811;

      end if;

   when s571 =>
      if ( x30 and x9 and x10 and x8 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x30 and x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s568;

      elsif ( x30 and x9 and not x10 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x30 and x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s569;

      elsif ( x30 and not x9 and x10 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x30 and not x9 and x10 and not x8 and x27 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( x30 and not x9 and x10 and not x8 and not x27 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x30 and not x9 and not x10 and x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s570;

      elsif ( x30 and not x9 and not x10 and not x8 and x26 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( x30 and not x9 and not x10 and not x8 and not x26 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x30 and x31 and x9 and x10 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( not x30 and x31 and x9 and x10 and not x8 and x21 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x30 and x31 and x9 and x10 and not x8 and not x21 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and x9 and x10 and not x8 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and x9 and not x10 and x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( not x30 and x31 and x9 and not x10 and not x8 and x18 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x30 and x31 and x9 and not x10 and not x8 and not x18 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and x9 and not x10 and not x8 and not x18 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and not x9 and x8 and x10 and x19 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x30 and x31 and not x9 and x8 and x10 and not x19 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and not x9 and x8 and x10 and not x19 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and not x9 and x8 and not x10 and x20 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x30 and x31 and not x9 and x8 and not x10 and not x20 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x30 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and not x9 and x8 and not x10 and not x20 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x30 and x31 and not x9 and not x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      else
         y9 <= '1' ;
         current_otherm <= s572;

      end if;

   when s572 =>
      if ( x65 ) = '1' then
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s487;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s842;

      end if;

   when s573 =>
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s843;

   when s574 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y60 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s844;

   when s575 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s845;

   when s576 =>
      if ( x6 and x8 and x7 ) = '1' then
         y63 <= '1' ;
         current_otherm <= s224;

      elsif ( x6 and x8 and not x7 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x6 and x8 and not x7 and x9 and not x18 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x6 and x8 and not x7 and x9 and not x18 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x6 and x8 and not x7 and x9 and not x18 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x8 and not x7 and x9 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x8 and not x7 and not x9 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x6 and x8 and not x7 and not x9 and not x19 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x6 and x8 and not x7 and not x9 and not x19 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x6 and x8 and not x7 and not x9 and not x19 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and x8 and not x7 and not x9 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x8 and x9 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s575;

      elsif ( x6 and not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x6 and not x8 and not x9 and x7 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x6 and not x8 and not x9 and x7 and not x17 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x6 and not x8 and not x9 and x7 and not x17 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x6 and not x8 and not x9 and x7 and not x17 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x8 and not x9 and x7 and not x17 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x8 and not x9 and not x7 ) = '1' then
         y65 <= '1' ;
         current_otherm <= s155;

      else
         y57 <= '1' ;
         current_otherm <= s135;

      end if;

   when s577 =>
      if ( x63 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y38 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s250;

      else
         y55 <= '1' ;
         current_otherm <= s254;

      end if;

   when s578 =>
         y56 <= '1' ;
         current_otherm <= s412;

   when s579 =>
      if ( x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x22 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s580 =>
         y11 <= '1' ;
         current_otherm <= s425;

   when s581 =>
      if ( x8 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         y32 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s579;

      elsif ( not x8 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x8 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x8 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s582 =>
      if ( x63 and x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x63 and not x18 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      else
         y58 <= '1' ;
         current_otherm <= s774;

      end if;

   when s583 =>
      if ( x26 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x26 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x26 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x26 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x26 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x12 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x12 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x12 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x12 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x12 and not x22 ) = '1' then
         current_otherm <= s1;

      else
         y10 <= '1' ;
         current_otherm <= s16;

      end if;

   when s584 =>
      if ( x63 ) = '1' then
         y68 <= '1' ;
         current_otherm <= s743;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s585 =>
      if ( x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s586 =>
      if ( x66 and x11 and x13 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s88;

      elsif ( x66 and x11 and x13 and x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s846;

      elsif ( x66 and x11 and x13 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s847;

      elsif ( x66 and x11 and x13 and not x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s848;

      elsif ( x66 and x11 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x11 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x11 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x11 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and x15 and x13 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x66 and not x11 and x12 and x15 and x13 and not x14 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( x66 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and x15 and x13 and not x14 and not x16 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and x15 and not x13 and x14 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s460;

      elsif ( x66 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and x15 and not x13 and x14 and not x18 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and x15 and not x13 and not x14 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x66 and not x11 and x12 and not x15 and x13 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( x66 and not x11 and x12 and not x15 and x13 and not x14 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( x66 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and not x15 and not x13 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s849;

      elsif ( x66 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and x12 and not x15 and not x13 and not x14 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s850;

      elsif ( not x66 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s585;

      elsif ( not x66 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x66 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s716;

      elsif ( not x66 and not x20 and x4 and x21 and x6 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      elsif ( not x66 and not x20 and x4 and x21 and x6 and not x5 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x66 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and x4 and x21 and x6 and not x5 and not x11 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and x4 and x21 and not x6 and x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s719;

      elsif ( not x66 and not x20 and x4 and x21 and not x6 and not x5 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x66 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x66 and not x20 and not x4 and x21 and x6 and x5 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x66 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and not x4 and x21 and x6 and x5 and not x13 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and not x4 and x21 and x6 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x66 and not x20 and not x4 and x21 and not x6 and x5 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x66 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x20 and not x4 and x21 and not x6 and not x5 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      end if;

   when s587 =>
      if ( x7 ) = '1' then
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s585;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s588 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s851;

   when s589 =>
      if ( x7 ) = '1' then
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s585;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s590 =>
      if ( x17 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s852;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s590;

      end if;

   when s591 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s848;

   when s592 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s853;

   when s593 =>
      if ( x33 and x32 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s854;

      else
         y9 <= '1' ;
         current_otherm <= s854;

      end if;

   when s594 =>
      if ( x62 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s72;

      elsif ( not x62 and x63 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s855;

      else
         y15 <= '1' ;
         current_otherm <= s111;

      end if;

   when s595 =>
         y6 <= '1' ;
         current_otherm <= s346;

   when s596 =>
         y38 <= '1' ;
         current_otherm <= s261;

   when s597 =>
         y27 <= '1' ;
         current_otherm <= s465;

   when s598 =>
         y6 <= '1' ;
         current_otherm <= s856;

   when s599 =>
         y32 <= '1' ;
         current_otherm <= s120;

   when s600 =>
         y32 <= '1' ;
         current_otherm <= s857;

   when s601 =>
         y58 <= '1' ;
         current_otherm <= s858;

   when s602 =>
      if ( x66 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

      else
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1;

      end if;

   when s603 =>
         y9 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s1;

   when s604 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s859;

   when s605 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s860;

   when s606 =>
      if ( x63 and x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s397;

      elsif ( x63 and not x20 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s727;

      else
         y6 <= '1' ;
         current_otherm <= s100;

      end if;

   when s607 =>
         y28 <= '1' ;
         current_otherm <= s861;

   when s608 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s862;

   when s609 =>
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s863;

   when s610 =>
      if ( x3 and x5 and x7 and x9 and x11 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      elsif ( x3 and x5 and x7 and x9 and not x11 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( x3 and x5 and x7 and not x9 and x10 and x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( x3 and x5 and x7 and not x9 and x10 and x11 and not x12 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x3 and x5 and x7 and not x9 and x10 and x11 and not x12 and x19 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x7 and not x9 and x10 and x11 and not x12 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x7 and not x9 and x10 and not x11 and x13 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( x3 and x5 and x7 and not x9 and x10 and not x11 and not x13 and x19 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x3 and x5 and x7 and not x9 and x10 and not x11 and not x13 and x19 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x7 and not x9 and x10 and not x11 and not x13 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x7 and not x9 and not x10 and x11 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s864;

      elsif ( x3 and x5 and x7 and not x9 and not x10 and not x11 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s864;

      elsif ( x3 and x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s865;

      elsif ( x3 and not x5 and x8 and x7 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s864;

      elsif ( x3 and not x5 and x8 and not x7 and x9 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x3 and not x5 and x8 and not x7 and x9 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x3 and not x5 and x8 and not x7 and x9 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and not x5 and x8 and not x7 and x9 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and not x5 and x8 and not x7 and not x9 and x10 and x11 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s864;

      elsif ( x3 and not x5 and x8 and not x7 and not x9 and x10 and not x11 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s864;

      elsif ( x3 and not x5 and x8 and not x7 and not x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s864;

      elsif ( x3 and not x5 and not x8 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s865;

      else
         y3 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s866;

      end if;

   when s611 =>
         y28 <= '1' ;
         current_otherm <= s698;

   when s612 =>
         y28 <= '1' ;
         current_otherm <= s867;

   when s613 =>
         y13 <= '1' ;
         current_otherm <= s773;

   when s614 =>
      if ( x4 and x22 and x21 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x4 and x22 and not x21 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x4 and not x22 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s245;

      end if;

   when s615 =>
         y5 <= '1' ;
         current_otherm <= s268;

   when s616 =>
         y5 <= '1' ;
         current_otherm <= s72;

   when s617 =>
      if ( x62 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s474;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s311;

      else
         y13 <= '1' ;
         current_otherm <= s868;

      end if;

   when s618 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s869;

   when s619 =>
         y5 <= '1' ;
         current_otherm <= s398;

   when s620 =>
         y37 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s870;

   when s621 =>
         y5 <= '1' ;
         current_otherm <= s308;

   when s622 =>
      if ( x39 and x41 and x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s620;

      elsif ( x39 and x41 and not x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s315;

      elsif ( x39 and not x41 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s539;

      elsif ( not x39 and x40 and x55 and x56 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x39 and x40 and x55 and not x56 and x58 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( not x39 and x40 and x55 and not x56 and not x58 and x59 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x39 and x40 and x55 and not x56 and not x58 and not x59 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x39 and x40 and not x55 and x54 and x57 and x28 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x39 and x40 and not x55 and x54 and x57 and not x28 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x39 and x40 and not x55 and x54 and not x57 and x29 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x39 and x40 and not x55 and x54 and not x57 and not x29 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x39 and x40 and not x55 and not x54 and x53 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x39 and x40 and not x55 and not x54 and not x53 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      else
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s621;

      end if;

   when s623 =>
      if ( x62 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s176;

      elsif ( not x62 and x14 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s871;

      else
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s872;

      end if;

   when s624 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y44 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s873;

   when s625 =>
      if ( x51 and x41 and x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s620;

      elsif ( x51 and x41 and not x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s315;

      elsif ( x51 and not x41 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s539;

      elsif ( not x51 and x52 and x55 and x56 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x51 and x52 and x55 and not x56 and x58 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( not x51 and x52 and x55 and not x56 and not x58 and x59 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x51 and x52 and x55 and not x56 and not x58 and not x59 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x51 and x52 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x51 and x52 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x51 and x52 and x55 and not x56 and not x58 and not x59 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x51 and x52 and not x55 and x54 and x57 and x28 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x51 and x52 and not x55 and x54 and x57 and not x28 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x51 and x52 and not x55 and x54 and x57 and not x28 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x51 and x52 and not x55 and x54 and x57 and not x28 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x51 and x52 and not x55 and x54 and x57 and not x28 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x51 and x52 and not x55 and x54 and not x57 and x29 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x51 and x52 and not x55 and x54 and not x57 and not x29 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x51 and x52 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x51 and x52 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( not x51 and x52 and not x55 and x54 and not x57 and not x29 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( not x51 and x52 and not x55 and not x54 and x53 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( not x51 and x52 and not x55 and not x54 and not x53 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      else
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s616;

      end if;

   when s626 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s874;

   when s627 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s875;

   when s628 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s629 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s630 =>
      if ( x9 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      else
         current_otherm <= s630;

      end if;

   when s631 =>
      if ( x63 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x63 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x64 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      else
         y4 <= '1' ;
         current_otherm <= s165;

      end if;

   when s632 =>
      if ( x4 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s127;

      elsif ( not x4 and x31 and x30 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x4 and x31 and not x30 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s876;

      elsif ( not x4 and not x31 and x30 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s876;

      else
         y37 <= '1' ;
         current_otherm <= s675;

      end if;

   when s633 =>
      if ( x20 and x12 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x20 and not x12 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x20 and not x12 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x20 and not x12 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x20 and not x12 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x20 and not x12 and not x22 ) = '1' then
         current_otherm <= s1;

      else
         y26 <= '1' ;
         current_otherm <= s877;

      end if;

   when s634 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s878;

   when s635 =>
         y11 <= '1' ;
         current_otherm <= s350;

   when s636 =>
         y20 <= '1' ;
         current_otherm <= s173;

   when s637 =>
      if ( x20 and x21 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( x20 and not x21 and x4 and x6 and x14 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      elsif ( x20 and not x21 and x4 and x6 and not x14 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s879;

      elsif ( x20 and not x21 and x4 and not x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s788;

      elsif ( x20 and not x21 and not x4 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s880;

      elsif ( not x20 and x4 and x6 and x13 and x21 and x14 and x15 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x20 and x4 and x6 and x13 and x21 and x14 and not x15 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x4 and x6 and x13 and x21 and x14 and not x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and x15 and x17 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and x15 and x17 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and x15 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and x15 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and not x15 and x9 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and not x15 and x9 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and not x15 and not x9 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and x13 and x21 and not x14 and not x15 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and x13 and not x21 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s786;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and x15 and x18 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and x15 and x18 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and x15 and not x18 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and x15 and not x18 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and x15 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and x15 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and not x15 and x19 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and not x15 and x19 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and not x15 and not x19 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and not x15 and not x19 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and not x15 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and x14 and not x15 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and not x14 and x15 and x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and not x14 and x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s882;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and not x14 and not x15 and x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s883;

      elsif ( not x20 and x4 and x6 and not x13 and x21 and not x14 and not x15 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s884;

      elsif ( not x20 and x4 and x6 and not x13 and not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and not x13 and not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x4 and x6 and not x13 and not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x6 and not x13 and not x21 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and not x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s170;

      else
         y20 <= '1' ;
         current_otherm <= s788;

      end if;

   when s638 =>
         y13 <= '1' ;
         current_otherm <= s692;

   when s639 =>
      if ( x13 and x21 and x10 ) = '1' then
         y62 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y90 <= '1' ;
         current_otherm <= s546;

      elsif ( x13 and x21 and not x10 and x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s544;

      elsif ( x13 and x21 and not x10 and x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s547;

      elsif ( x13 and x21 and not x10 and not x14 and x11 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( x13 and x21 and not x10 and not x14 and not x11 ) = '1' then
         y3 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s549;

      elsif ( x13 and not x21 and x10 and x22 and x11 and x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s548;

      elsif ( x13 and not x21 and x10 and x22 and x11 and not x14 ) = '1' then
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s545;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and x14 and x19 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and x14 and not x19 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and not x14 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and x10 and x22 and not x11 and not x14 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and x10 and not x22 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s550;

      elsif ( x13 and not x21 and not x10 and x22 and x14 and x11 and x17 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and not x10 and x22 and x14 and x11 and not x17 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and not x10 and x22 and x14 and not x11 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and x18 ) = '1' then
         y12 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s240;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and x16 and not x18 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and x11 and not x16 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x21 and not x10 and x22 and not x14 and not x11 ) = '1' then
         y102 <= '1' ;
         current_otherm <= s240;

      elsif ( x13 and not x21 and not x10 and not x22 ) = '1' then
         y9 <= '1' ;
         y62 <= '1' ;
         y65 <= '1' ;
         y94 <= '1' ;
         current_otherm <= s551;

      else
         y9 <= '1' ;
         y65 <= '1' ;
         y84 <= '1' ;
         y86 <= '1' ;
         y91 <= '1' ;
         current_otherm <= s552;

      end if;

   when s640 =>
      if ( x22 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s108;

      else
         y60 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y92 <= '1' ;
         current_otherm <= s885;

      end if;

   when s641 =>
      if ( x62 and x17 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s886;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s334;

      elsif ( not x62 and x64 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s887;

      else
         y22 <= '1' ;
         current_otherm <= s888;

      end if;

   when s642 =>
         y5 <= '1' ;
         current_otherm <= s74;

   when s643 =>
      if ( x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s889;

      else
         y28 <= '1' ;
         current_otherm <= s727;

      end if;

   when s644 =>
         y14 <= '1' ;
         current_otherm <= s594;

   when s645 =>
      if ( x18 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s13;

      elsif ( not x18 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x18 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x18 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s646 =>
      if ( x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s237;

      else
         y7 <= '1' ;
         current_otherm <= s678;

      end if;

   when s647 =>
         y46 <= '1' ;
         current_otherm <= s890;

   when s648 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s891;

   when s649 =>
      if ( x64 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s465;

      elsif ( not x64 and x66 and x14 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s470;

      elsif ( not x64 and x66 and not x14 ) = '1' then
         y28 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s630;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      end if;

   when s650 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s892;

   when s651 =>
      if ( x63 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s893;

      elsif ( x63 and not x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s892;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s652 =>
      if ( x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s570;

      else
         y7 <= '1' ;
         current_otherm <= s646;

      end if;

   when s653 =>
      if ( x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s219;

      else
         y9 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s213;

      end if;

   when s654 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s894;

      else
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s654;

      end if;

   when s655 =>
      if ( x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_otherm <= s21;

      elsif ( not x5 and x6 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s895;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and x4 and x3 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y32 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s896;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and x4 and not x3 and x17 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and x4 and not x3 and not x17 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and x4 and not x3 and not x17 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and x4 and not x3 and not x17 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and x4 and not x3 and not x17 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and not x4 and x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s708;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and not x4 and not x3 and x16 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and not x4 and not x3 and not x16 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and x2 and x18 and x19 and not x4 and not x3 and not x16 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and x2 and x18 and not x19 and x3 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and x2 and x18 and not x19 and x3 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and x2 and x18 and not x19 and x3 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and x2 and x18 and not x19 and x3 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and x2 and x18 and not x19 and not x3 and x4 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x5 and not x6 and x2 and x18 and not x19 and not x3 and not x4 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( not x5 and not x6 and x2 and not x18 and x19 and x4 and x3 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( not x5 and not x6 and x2 and not x18 and x19 and x4 and not x3 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( not x5 and not x6 and x2 and not x18 and x19 and not x4 and x3 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( not x5 and not x6 and x2 and not x18 and x19 and not x4 and not x3 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s897;

      elsif ( not x5 and not x6 and x2 and not x18 and not x19 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and x19 and x3 and x15 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and x19 and x3 and not x15 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and x19 and x3 and not x15 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and x19 and x3 and not x15 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and x19 and x3 and not x15 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and x19 and not x3 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and not x19 and x3 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x5 and not x6 and not x2 and x18 and x4 and not x19 and not x3 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and x19 and x3 and x14 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and x19 and x3 and not x14 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and x19 and x3 and not x14 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and x19 and x3 and not x14 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and x19 and x3 and not x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and x19 and not x3 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and not x19 and x3 and x12 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and not x19 and x3 and not x12 and x11 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and not x19 and x3 and not x12 and x11 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and not x19 and x3 and not x12 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x6 and not x2 and x18 and not x4 and not x19 and not x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and not x18 and x19 and x4 and x3 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and not x18 and x19 and x4 and not x3 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s510;

      elsif ( not x5 and not x6 and not x2 and not x18 and x19 and not x4 and x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x5 and not x6 and not x2 and not x18 and x19 and not x4 and not x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s898;

      else
         y11 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s560;

      end if;

   when s656 =>
         y2 <= '1' ;
         current_otherm <= s502;

   when s657 =>
      if ( x3 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s899;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s900;

      end if;

   when s658 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s901;

   when s659 =>
      if ( x18 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      else
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s154;

      end if;

   when s660 =>
      if ( x63 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s460;

      end if;

   when s661 =>
      if ( x14 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s902;

      else
         y47 <= '1' ;
         y55 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s903;

      end if;

   when s662 =>
      if ( x64 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s904;

      elsif ( not x64 and x30 ) = '1' then
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      else
         y47 <= '1' ;
         y50 <= '1' ;
         y61 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s599;

      end if;

   when s663 =>
      if ( x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s905;

      elsif ( x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s906;

      elsif ( not x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s906;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s905;

      end if;

   when s664 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s905;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s906;

      end if;

   when s665 =>
         y13 <= '1' ;
         current_otherm <= s868;

   when s666 =>
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s545;

   when s667 =>
         y37 <= '1' ;
         current_otherm <= s510;

   when s668 =>
         y28 <= '1' ;
         current_otherm <= s377;

   when s669 =>
      if ( x21 and x20 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x21 and x20 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x21 and x20 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and x20 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s907;

      elsif ( not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s670 =>
      if ( x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y39 <= '1' ;
         current_otherm <= s103;

      end if;

   when s671 =>
         y48 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s908;

   when s672 =>
         y13 <= '1' ;
         current_otherm <= s909;

   when s673 =>
         y60 <= '1' ;
         y65 <= '1' ;
         y78 <= '1' ;
         y92 <= '1' ;
         current_otherm <= s546;

   when s674 =>
         y1 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s910;

   when s675 =>
      if ( x30 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s486;

      elsif ( not x30 and x31 ) = '1' then
         y47 <= '1' ;
         y51 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s671;

      else
         y5 <= '1' ;
         current_otherm <= s352;

      end if;

   when s676 =>
      if ( x63 and x67 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s911;

      elsif ( x63 and not x67 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and not x67 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and not x67 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x67 and not x14 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s912;

      end if;

   when s677 =>
      if ( x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s678 =>
      if ( x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x63 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s679 =>
      if ( x63 and x14 and x10 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and x14 and not x10 and x11 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x63 and x14 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x63 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s810;

      end if;

   when s680 =>
      if ( x12 and x4 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s681;

      elsif ( x12 and not x4 and x5 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s682;

      elsif ( x12 and not x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s677;

      elsif ( not x12 and x4 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s677;

      elsif ( not x12 and x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s683;

      else
         y1 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s684;

      end if;

   when s681 =>
         y17 <= '1' ;
         current_otherm <= s3;

   when s682 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s677;

   when s683 =>
         y3 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s677;

   when s684 =>
      if ( x5 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s677;

      else
         y9 <= '1' ;
         current_otherm <= s43;

      end if;

   when s685 =>
      if ( x15 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      else
         current_otherm <= s1;

      end if;

   when s686 =>
      if ( x10 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s913;

      elsif ( not x10 and x14 and x6 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x14 and x6 and not x5 and x7 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s890;

      elsif ( not x10 and x14 and x6 and not x5 and x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y19 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s914;

      elsif ( not x10 and x14 and x6 and not x5 and x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x10 and x14 and x6 and not x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x10 and x14 and not x6 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s890;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s915;

      end if;

   when s687 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s916;

   when s688 =>
      if ( x5 and x7 and x9 and x6 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( x5 and x7 and x9 and not x6 and x8 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x5 and x7 and x9 and not x6 and not x8 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x5 and x7 and not x9 and x6 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x5 and x7 and not x9 and not x6 and x8 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( x5 and x7 and not x9 and not x6 and not x8 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s917;

      elsif ( x5 and not x7 and x9 and x6 and x8 and x12 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x5 and not x7 and x9 and x6 and x8 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and not x7 and x9 and x6 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s918;

      elsif ( x5 and not x7 and x9 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      elsif ( x5 and not x7 and x9 and not x6 and not x10 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s919;

      elsif ( x5 and not x7 and x9 and not x6 and not x10 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y15 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s795;

      elsif ( x5 and not x7 and not x9 and x8 and x6 and x13 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x5 and not x7 and not x9 and x8 and x6 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and not x7 and not x9 and x8 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s915;

      elsif ( x5 and not x7 and not x9 and x8 and not x6 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s795;

      elsif ( x5 and not x7 and not x9 and not x8 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s708;

      elsif ( x5 and not x7 and not x9 and not x8 and not x6 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x5 and x6 and x8 and x7 and x10 and x3 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s687;

      elsif ( not x5 and x6 and x8 and x7 and x10 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( not x5 and x6 and x8 and x7 and x10 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      elsif ( not x5 and x6 and x8 and x7 and not x10 ) = '1' then
         y72 <= '1' ;
         current_otherm <= s685;

      elsif ( not x5 and x6 and x8 and not x7 and x9 and x18 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( not x5 and x6 and x8 and not x7 and x9 and x18 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      elsif ( not x5 and x6 and x8 and not x7 and x9 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and x8 and not x7 and not x9 and x17 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( not x5 and x6 and x8 and not x7 and not x9 and x17 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      elsif ( not x5 and x6 and x8 and not x7 and not x9 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and not x8 and x9 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( not x5 and x6 and not x8 and x9 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      elsif ( not x5 and x6 and not x8 and not x9 and x7 and x16 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s686;

      elsif ( not x5 and x6 and not x8 and not x9 and x7 and x16 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      elsif ( not x5 and x6 and not x8 and not x9 and x7 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and not x8 and not x9 and not x7 ) = '1' then
         y71 <= '1' ;
         current_otherm <= s156;

      elsif ( not x5 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s915;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s916;

      end if;

   when s689 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s733;

      end if;

   when s690 =>
      if ( x18 and x22 and x23 and x4 and x3 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x18 and x22 and x23 and x4 and x3 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x18 and x22 and x23 and x4 and x3 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and x4 and x3 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and x4 and not x3 and x5 and x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x18 and x22 and x23 and x4 and not x3 and x5 and not x15 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x18 and x22 and x23 and x4 and not x3 and x5 and not x15 and x21 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and x4 and not x3 and x5 and not x15 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and x4 and not x3 and not x5 and x16 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x18 and x22 and x23 and x4 and not x3 and not x5 and not x16 and x21 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x18 and x22 and x23 and x4 and not x3 and not x5 and not x16 and x21 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and x4 and not x3 and not x5 and not x16 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and not x4 and x5 and x3 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and not x4 and x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and x22 and x23 and not x4 and not x5 and x3 ) = '1' then
         y51 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s1;

      elsif ( x18 and x22 and x23 and not x4 and not x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and x22 and not x23 and x9 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and x22 and not x23 and not x9 and x3 and x5 and x4 ) = '1' then
         y42 <= '1' ;
         current_otherm <= s354;

      elsif ( x18 and x22 and not x23 and not x9 and x3 and x5 and not x4 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( x18 and x22 and not x23 and not x9 and x3 and not x5 and x4 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x22 and not x23 and not x9 and x3 and not x5 and not x4 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( x18 and x22 and not x23 and not x9 and not x3 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y11 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and x22 and not x23 and not x9 and not x3 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s920;

      elsif ( x18 and not x22 and x23 and x9 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s401;

      elsif ( x18 and not x22 and x23 and not x9 and x10 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s921;

      elsif ( x18 and not x22 and x23 and not x9 and x10 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s920;

      elsif ( x18 and not x22 and x23 and not x9 and not x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s920;

      elsif ( x18 and not x22 and not x23 and x3 and x5 and x4 ) = '1' then
         y31 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and not x22 and not x23 and x3 and x5 and not x4 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x18 and not x22 and not x23 and x3 and not x5 and x4 ) = '1' then
         y30 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and not x22 and not x23 and x3 and not x5 and not x4 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( x18 and not x22 and not x23 and not x3 and x8 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s302;

      elsif ( x18 and not x22 and not x23 and not x3 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s920;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s922;

      end if;

   when s691 =>
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s923;

   when s692 =>
      if ( x62 and x17 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s94;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s638;

      elsif ( not x62 and x63 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s693 =>
      if ( x11 and x19 and x20 and x2 and x1 and x4 and x3 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and x3 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and x3 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and x3 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and x18 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and x21 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x19 and x20 and x2 and x1 and not x4 and x5 and x3 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x11 and x19 and x20 and x2 and x1 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x19 and x20 and x2 and x1 and not x4 and not x5 and x3 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x11 and x19 and x20 and x2 and x1 and not x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y34 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x19 and x20 and x2 and not x1 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( x11 and x19 and x20 and not x2 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s696;

      elsif ( x11 and x19 and x20 and not x2 and not x8 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( x11 and x19 and not x20 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s697;

      elsif ( x11 and not x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s698;

      else
         y29 <= '1' ;
         current_otherm <= s378;

      end if;

   when s694 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s924;

   when s695 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s925;

   when s696 =>
      if ( x2 ) = '1' then
         current_otherm <= s1;

      elsif ( not x2 and x3 and x4 and x5 and x1 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x2 and x3 and x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and x3 and x4 and not x5 and x1 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x2 and x3 and x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and x3 and not x4 and x5 and x1 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x2 and x3 and not x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and x3 and not x4 and not x5 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and x3 and not x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and not x3 and x4 and x5 and x1 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( not x2 and not x3 and x4 and x5 and x1 and not x6 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( not x2 and not x3 and x4 and x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s340;

      elsif ( not x2 and not x3 and x4 and x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and not x3 and x4 and not x5 and x1 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( not x2 and not x3 and x4 and not x5 and x1 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( not x2 and not x3 and x4 and not x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and not x3 and x4 and not x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and not x3 and not x4 and x1 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( not x2 and not x3 and not x4 and x1 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      else
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y32 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      end if;

   when s697 =>
      if ( x6 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s803;

      elsif ( not x6 and x2 and x1 and x4 and x3 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x6 and x2 and x1 and x4 and x3 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x6 and x2 and x1 and x4 and x3 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x2 and x1 and x4 and x3 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and x5 and x18 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and x5 and not x18 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and not x5 and x21 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x2 and x1 and x4 and not x3 and not x5 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x2 and x1 and not x4 and x5 and x3 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x6 and x2 and x1 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and x2 and x1 and not x4 and not x5 and x3 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x2 and x1 and not x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y34 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and x2 and not x1 and x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s926;

      elsif ( not x6 and x2 and not x1 and not x3 and x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s926;

      elsif ( not x6 and x2 and not x1 and not x3 and not x4 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s926;

      elsif ( not x6 and x2 and not x1 and not x3 and not x4 and not x5 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x6 and not x2 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s927;

      elsif ( not x6 and not x2 and not x7 and x3 and x4 and x5 and x1 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x6 and not x2 and not x7 and x3 and x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and not x2 and not x7 and x3 and x4 and not x5 and x1 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( not x6 and not x2 and not x7 and x3 and x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and not x2 and not x7 and x3 and not x4 and x5 and x1 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( not x6 and not x2 and not x7 and x3 and not x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and not x2 and not x7 and x3 and not x4 and not x5 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and not x2 and not x7 and x3 and not x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s342;

      elsif ( not x6 and not x2 and not x7 and not x3 and x1 and x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      elsif ( not x6 and not x2 and not x7 and not x3 and x1 and not x5 and x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_otherm <= s79;

      elsif ( not x6 and not x2 and not x7 and not x3 and x1 and not x5 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s736;

      end if;

   when s698 =>
      if ( x65 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s928;

      elsif ( not x65 and x21 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( not x65 and x21 and not x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s929;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s929;

      end if;

   when s699 =>
      if ( x16 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x16 and not x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      else
         y35 <= '1' ;
         current_otherm <= s386;

      end if;

   when s700 =>
      if ( x15 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s631;

      else
         y35 <= '1' ;
         current_otherm <= s386;

      end if;

   when s701 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s358;

   when s702 =>
         y47 <= '1' ;
         y55 <= '1' ;
         y61 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s930;

   when s703 =>
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s931;

   when s704 =>
         y47 <= '1' ;
         y55 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s903;

   when s705 =>
         y55 <= '1' ;
         current_otherm <= s109;

   when s706 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s932;

   when s707 =>
      if ( x15 and x5 ) = '1' then
         y44 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s933;

      elsif ( x15 and not x5 and x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( x15 and not x5 and not x21 and x8 and x9 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s820;

      elsif ( x15 and not x5 and not x21 and x8 and not x9 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s820;

      elsif ( x15 and not x5 and not x21 and not x8 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s820;

      else
         y6 <= '1' ;
         y12 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s934;

      end if;

   when s708 =>
         y36 <= '1' ;
         current_otherm <= s260;

   when s709 =>
      if ( x18 and x19 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x19 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s560;

      elsif ( not x18 and x19 ) = '1' then
         y23 <= '1' ;
         y29 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s935;

      elsif ( not x18 and not x19 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s936;

      else
         y11 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s560;

      end if;

   when s710 =>
      if ( x21 ) = '1' then
         y80 <= '1' ;
         current_otherm <= s937;

      else
         y80 <= '1' ;
         current_otherm <= s938;

      end if;

   when s711 =>
         y80 <= '1' ;
         current_otherm <= s937;

   when s712 =>
      if ( x15 and x17 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x15 and not x17 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x15 and not x17 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x15 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x15 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y46 <= '1' ;
         current_otherm <= s110;

      end if;

   when s713 =>
      if ( x38 and x39 and x41 and x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s620;

      elsif ( x38 and x39 and x41 and not x42 ) = '1' then
         y1 <= '1' ;
         y37 <= '1' ;
         y40 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s315;

      elsif ( x38 and x39 and not x41 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s539;

      elsif ( x38 and not x39 and x40 and x55 and x56 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( x38 and not x39 and x40 and x55 and not x56 and x58 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( x38 and not x39 and x40 and x55 and not x56 and not x58 and x59 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x38 and not x39 and x40 and x55 and not x56 and not x58 and not x59 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and x57 and x28 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and x57 and not x28 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and not x57 and x29 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and x37 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and x3 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and x27 and not x37 and not x3 ) = '1' then
         current_otherm <= s1;

      elsif ( x38 and not x39 and x40 and not x55 and x54 and not x57 and not x29 and not x27 ) = '1' then
         current_otherm <= s1;

      elsif ( x38 and not x39 and x40 and not x55 and not x54 and x53 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s315;

      elsif ( x38 and not x39 and x40 and not x55 and not x54 and not x53 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( x38 and not x39 and not x40 ) = '1' then
         y1 <= '1' ;
         y13 <= '1' ;
         y37 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s621;

      else
         y2 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s622;

      end if;

   when s714 =>
      if ( x63 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s939;

      elsif ( not x63 and x66 and x30 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s99;

      elsif ( not x63 and x66 and not x30 ) = '1' then
         y47 <= '1' ;
         y49 <= '1' ;
         y58 <= '1' ;
         y61 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s573;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s715 =>
      if ( x3 and x4 and x6 and x8 and x9 and x12 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( x3 and x4 and x6 and x8 and x9 and not x12 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and x11 and x16 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and x11 and not x16 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and x11 and not x16 and x14 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and x11 and not x16 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and not x11 and x15 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and not x11 and not x15 and x14 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and not x11 and not x15 and x14 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x6 and x8 and not x9 and x10 and not x11 and not x15 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x6 and x8 and not x9 and not x10 and x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         y51 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and x4 and x6 and x8 and not x9 and not x10 and not x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and x4 and x6 and not x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s940;

      elsif ( x3 and x4 and not x6 and x12 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and not x6 and x12 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and not x6 and x12 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and not x6 and x12 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and x10 and x8 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and x10 and x8 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and x10 and x8 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and x10 and x8 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and x10 and not x8 and x11 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and x10 and not x8 and not x11 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and not x10 and x8 and x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and not x10 and x8 and not x11 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and not x10 and x8 and not x11 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and not x10 and x8 and not x11 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and not x10 and x8 and not x11 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and not x6 and x12 and not x9 and not x10 and not x8 ) = '1' then
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and x4 and not x6 and not x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s940;

      elsif ( x3 and not x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s941;

      else
         y14 <= '1' ;
         current_otherm <= s594;

      end if;

   when s716 =>
      if ( x7 ) = '1' then
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s585;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s717 =>
      if ( x67 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s942;

      else
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s676;

      end if;

   when s718 =>
      if ( x66 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and x67 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and x67 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and x67 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and x67 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x66 and not x67 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x67 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and not x67 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s719 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

   when s720 =>
      if ( x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s585;

      elsif ( x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s716;

      elsif ( not x20 and x4 and x21 and x6 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      elsif ( not x20 and x4 and x21 and x6 and not x5 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x21 and x6 and not x5 and not x11 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x21 and not x6 and x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s719;

      elsif ( not x20 and x4 and x21 and not x6 and not x5 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and x21 and not x6 and not x5 and not x10 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x20 and not x4 and x21 and x6 and x5 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x4 and x21 and x6 and x5 and not x13 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x4 and x21 and x6 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x20 and not x4 and x21 and not x6 and x5 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x4 and x21 and not x6 and x5 and not x14 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x4 and x21 and not x6 and not x5 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      end if;

   when s721 =>
      if ( x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s943;

      elsif ( not x33 and x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s943;

      elsif ( not x33 and not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x33 and not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x33 and not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s722 =>
         y2 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s405;

   when s723 =>
      if ( x20 and x26 and x27 and x7 and x8 and x6 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and x27 and x7 and x8 and not x6 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and x27 and x7 and not x8 and x6 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and x27 and x7 and not x8 and not x6 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and x27 and not x7 and x6 and x8 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and x27 and not x7 and x6 and not x8 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and x27 and not x7 and not x6 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( x20 and x26 and not x27 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s944;

      elsif ( x20 and not x26 ) = '1' then
         y58 <= '1' ;
         current_otherm <= s858;

      else
         y26 <= '1' ;
         current_otherm <= s116;

      end if;

   when s724 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s945;

   when s725 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s946;

   when s726 =>
      if ( x64 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s947;

      else
         y48 <= '1' ;
         y55 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s908;

      end if;

   when s727 =>
      if ( x65 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s948;

      elsif ( not x65 and x20 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      else
         y15 <= '1' ;
         current_otherm <= s414;

      end if;

   when s728 =>
      if ( x3 and x5 and x30 and x31 and x9 and x8 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x3 and x5 and x30 and x31 and x9 and x8 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x3 and x5 and x30 and x31 and x9 and x8 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and x9 and x8 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and x10 and x25 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and x10 and not x25 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and x10 and not x25 and x23 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and x10 and not x25 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and not x10 and x24 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and not x10 and not x24 and x23 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and not x10 and not x24 and x23 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and x9 and not x8 and not x10 and not x24 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and not x9 and x10 and x8 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and not x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s356;

      elsif ( x3 and x5 and x30 and x31 and not x9 and not x10 and x8 ) = '1' then
         y10 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1;

      elsif ( x3 and x5 and x30 and x31 and not x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s287;

      elsif ( x3 and x5 and x30 and not x31 and x13 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s183;

      elsif ( x3 and x5 and x30 and not x31 and not x13 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s534;

      elsif ( x3 and x5 and not x30 and x31 and x15 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x3 and x5 and not x30 and x31 and x15 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x3 and x5 and not x30 and x31 and x15 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and not x30 and x31 and x15 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x5 and not x30 and x31 and not x15 and x16 and x13 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s534;

      elsif ( x3 and x5 and not x30 and x31 and not x15 and x16 and not x13 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( x3 and x5 and not x30 and x31 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( x3 and x5 and not x30 and not x31 and x8 and x9 ) = '1' then
         y47 <= '1' ;
         y55 <= '1' ;
         y63 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s512;

      elsif ( x3 and x5 and not x30 and not x31 and x8 and not x9 ) = '1' then
         y47 <= '1' ;
         y56 <= '1' ;
         y63 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s512;

      elsif ( x3 and x5 and not x30 and not x31 and not x8 and x13 ) = '1' then
         y45 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         y55 <= '1' ;
         y59 <= '1' ;
         y63 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s512;

      elsif ( x3 and x5 and not x30 and not x31 and not x8 and not x13 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s274;

      elsif ( x3 and not x5 and x31 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s534;

      elsif ( x3 and not x5 and x31 and not x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s949;

      elsif ( x3 and not x5 and not x31 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s662;

      elsif ( x3 and not x5 and not x31 and not x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s199;

      else
         y34 <= '1' ;
         current_otherm <= s631;

      end if;

   when s729 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s950;

   when s730 =>
      if ( x3 and x4 and x33 and x32 and x13 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s854;

      elsif ( x3 and x4 and x33 and x32 and x13 and not x15 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s593;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and x15 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s951;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and x15 and not x12 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and x15 and not x12 and x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and x15 and not x12 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and not x15 and x11 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s952;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and not x15 and not x11 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and not x15 and not x11 and x10 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x33 and x32 and not x13 and x14 and not x15 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x4 and x33 and x32 and not x13 and not x14 and x15 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x3 and x4 and x33 and x32 and not x13 and not x14 and not x15 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s443;

      elsif ( x3 and x4 and x33 and not x32 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( x3 and x4 and not x33 and x6 and x32 and x14 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s765;

      elsif ( x3 and x4 and not x33 and x6 and x32 and not x14 ) = '1' then
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s953;

      elsif ( x3 and x4 and not x33 and x6 and not x32 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s148;

      elsif ( x3 and x4 and not x33 and not x6 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s48;

      elsif ( x3 and not x4 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s149;

      else
         y8 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s954;

      end if;

   when s731 =>
         y19 <= '1' ;
         current_otherm <= s166;

   when s732 =>
      if ( x17 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s955;

      else
         y5 <= '1' ;
         y13 <= '1' ;
         y30 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s732;

      end if;

   when s733 =>
      if ( x20 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y42 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s395;

      else
         y22 <= '1' ;
         current_otherm <= s92;

      end if;

   when s734 =>
         y2 <= '1' ;
         current_otherm <= s504;

   when s735 =>
         y24 <= '1' ;
         current_otherm <= s955;

   when s736 =>
      if ( x64 and x63 and x4 and x5 and x3 ) = '1' then
         y41 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and x4 and x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and x4 and not x5 and x3 ) = '1' then
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and x4 and not x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and not x4 and x3 and x5 ) = '1' then
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and not x4 and x3 and not x5 ) = '1' then
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and x63 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y32 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x64 and not x63 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( not x64 and x63 and x66 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s434;

      elsif ( not x64 and x63 and not x66 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s956;

      elsif ( not x64 and not x63 and x65 ) = '1' then
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s957;

      elsif ( not x64 and not x63 and not x65 and x67 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      else
         y6 <= '1' ;
         current_otherm <= s100;

      end if;

   when s737 =>
      if ( x18 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s736;

      else
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s737;

      end if;

   when s738 =>
      if ( x63 and x22 and x23 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s556;

      elsif ( x63 and x22 and not x23 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s357;

      elsif ( x63 and not x22 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s357;

      else
         y48 <= '1' ;
         current_otherm <= s411;

      end if;

   when s739 =>
      if ( x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s509;

      else
         y7 <= '1' ;
         current_otherm <= s652;

      end if;

   when s740 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s753;

   when s741 =>
      if ( x15 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x15 and x3 and x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      elsif ( not x15 and x3 and x6 and not x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s834;

      elsif ( not x15 and x3 and not x6 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s834;

      elsif ( not x15 and x3 and not x6 and not x5 and x10 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y32 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      elsif ( not x15 and x3 and not x6 and not x5 and not x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s834;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and x6 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and x13 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and x13 and not x8 and x12 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and x13 and not x8 and not x12 and x16 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and x13 and not x8 and not x12 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and not x13 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and not x13 and x16 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and x7 and not x6 and not x13 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x7 and x6 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( not x15 and not x3 and x4 and x1 and not x7 and not x6 and x8 ) = '1' then
         y23 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s958;

      elsif ( not x15 and not x3 and x4 and x1 and not x7 and not x6 and not x8 ) = '1' then
         y11 <= '1' ;
         y15 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s958;

      elsif ( not x15 and not x3 and x4 and not x1 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s959;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and x8 and x7 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and x8 and not x7 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and not x8 and x7 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and not x8 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      elsif ( not x15 and not x3 and not x4 and x5 and x7 and x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s960;

      elsif ( not x15 and not x3 and not x4 and x5 and x7 and not x6 and x11 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x15 and not x3 and not x4 and x5 and x7 and not x6 and not x11 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x15 and not x3 and not x4 and x5 and x7 and not x6 and not x11 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x15 and not x3 and not x4 and x5 and x7 and not x6 and not x11 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and x7 and not x6 and not x11 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and x8 and x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s961;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and x8 and not x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s962;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and not x8 and x6 and x11 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and not x8 and x6 and not x11 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and not x8 and x6 and not x11 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and not x8 and x6 and not x11 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and not x8 and x6 and not x11 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x7 and not x8 and not x6 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x15 and not x3 and not x4 and not x5 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s959;

      elsif ( not x15 and not x3 and not x4 and not x5 and not x9 and x6 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s744;

      else
         y5 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      end if;

   when s742 =>
      if ( x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s743 =>
      if ( x63 and x66 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      elsif ( x63 and not x66 and x11 and x6 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and not x66 and x11 and x6 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and x12 and x18 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and x12 and not x18 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and not x12 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x66 and x11 and not x6 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and x11 and not x6 and not x7 and not x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and not x11 and x6 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s963;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and not x12 and x10 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and not x13 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x66 and not x11 and not x6 and x7 and not x12 and not x10 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x63 and not x66 and not x11 and not x6 and not x7 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      elsif ( not x63 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s744 =>
      if ( x63 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x63 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s745 =>
      if ( x65 and x10 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s964;

      elsif ( x65 and not x10 and x18 and x8 and x7 ) = '1' then
         y5 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s965;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and x9 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and x9 and not x14 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and x9 and not x14 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and x9 and not x14 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and x9 and not x14 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and not x9 and x12 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and not x9 and not x12 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and not x9 and not x12 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and not x9 and not x12 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x10 and x18 and x8 and not x7 and not x9 and not x12 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x10 and x18 and not x8 and x9 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s966;

      elsif ( x65 and not x10 and x18 and not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( x65 and not x10 and x18 and not x8 and not x9 and x7 and x13 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x65 and not x10 and x18 and not x8 and not x9 and x7 and not x13 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x10 and x18 and not x8 and not x9 and x7 and not x13 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x10 and x18 and not x8 and not x9 and x7 and not x13 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x10 and x18 and not x8 and not x9 and x7 and not x13 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x10 and x18 and not x8 and not x9 and not x7 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      elsif ( x65 and not x10 and not x18 ) = '1' then
         y5 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s968;

      elsif ( not x65 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x65 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x65 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s746 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s969;

   when s747 =>
      if ( x10 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s970;

      elsif ( not x10 and x18 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s971;

      elsif ( not x10 and x18 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s742;

      elsif ( not x10 and x18 and not x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      else
         y5 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s972;

      end if;

   when s748 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s973;

   when s749 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y40 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s974;

   when s750 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s742;

   when s751 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s742;

   when s752 =>
      if ( x10 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s975;

      elsif ( not x10 and x18 and x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y55 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s976;

      elsif ( not x10 and x18 and x8 and x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x10 and x18 and x8 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y47 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s977;

      elsif ( not x10 and x18 and x8 and not x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x10 and x18 and not x8 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y66 <= '1' ;
         y67 <= '1' ;
         current_otherm <= s978;

      elsif ( not x10 and x18 and not x8 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s979;

      elsif ( not x10 and x18 and not x8 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      else
         y5 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s980;

      end if;

   when s753 =>
      if ( x65 and x4 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s714;

      elsif ( x65 and not x4 and x5 and x6 and x9 and x7 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x65 and not x4 and x5 and x6 and x9 and not x7 and x8 and x17 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x65 and not x4 and x5 and x6 and x9 and not x7 and x8 and not x17 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and x5 and x6 and x9 and not x7 and x8 and not x17 and x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x5 and x6 and x9 and not x7 and x8 and not x17 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x5 and x6 and x9 and not x7 and not x8 ) = '1' then
         y5 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and x7 ) = '1' then
         y68 <= '1' ;
         current_otherm <= s743;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and not x7 and x8 and x18 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and not x7 and x8 and not x18 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and not x7 and x8 and not x18 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and not x7 and x8 and not x18 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and not x7 and x8 and not x18 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and x5 and x6 and not x9 and not x7 and not x8 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s744;

      elsif ( x65 and not x4 and x5 and not x6 and x7 and x9 and x8 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( x65 and not x4 and x5 and not x6 and x7 and x9 and not x8 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s118;

      elsif ( x65 and not x4 and x5 and not x6 and x7 and not x9 and x8 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s258;

      elsif ( x65 and not x4 and x5 and not x6 and x7 and not x9 and not x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and x8 and x3 and x11 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s746;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and x8 and x3 and x11 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and x8 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s747;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and x8 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s972;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and x8 and not x3 and not x10 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y35 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s981;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and x8 and not x3 and not x10 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s982;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and not x8 and x9 and x3 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and not x8 and x9 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s747;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and not x8 and x9 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s972;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and not x8 and x9 and not x3 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s983;

      elsif ( x65 and not x4 and x5 and not x6 and not x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and not x5 and x6 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s745;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and x7 ) = '1' then
         y5 <= '1' ;
         y19 <= '1' ;
         y30 <= '1' ;
         y39 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s984;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and x9 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and x9 and not x14 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and x9 and not x14 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and x9 and not x14 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and x9 and not x14 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and not x9 and x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and not x9 and not x12 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and not x9 and not x12 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and not x9 and not x12 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and x8 and not x7 and not x9 and not x12 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s985;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s986;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and not x9 and x7 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and not x9 and x7 and not x13 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and not x9 and x7 and not x13 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and not x9 and x7 and not x13 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and not x9 and x7 and not x13 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x4 and not x5 and x6 and not x3 and not x8 and not x9 and not x7 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s748;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and x8 and x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and x8 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s749;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and x8 and not x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and not x8 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s750;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and not x8 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y40 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s751;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and x11 and not x8 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and not x5 and not x6 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s752;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s980;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s987;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and x8 and x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and x8 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s988;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and x8 and not x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and not x8 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s829;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and not x8 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s542;

      elsif ( x65 and not x4 and not x5 and not x6 and not x3 and not x10 and not x8 and not x7 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s742;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s736;

      end if;

   when s754 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s399;

      elsif ( not x3 and x19 and x20 and x5 and x6 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s585;

      elsif ( not x3 and x19 and x20 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x3 and x19 and x20 and not x5 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s716;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x6 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x6 and not x5 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and x6 and not x5 and not x11 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x6 and x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s719;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x6 and not x5 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and x21 and not x6 and not x5 and not x10 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x6 and x5 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x6 and x5 and not x13 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and x6 and not x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x6 and x5 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x6 and x5 and not x14 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x3 and x19 and not x20 and not x4 and x21 and not x6 and not x5 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x3 and x19 and not x20 and not x4 and not x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s585;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s720;

      end if;

   when s755 =>
      if ( x7 ) = '1' then
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s585;

      elsif ( not x7 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x7 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s756 =>
      if ( x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s757 =>
      if ( x14 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s756;

      elsif ( x14 and not x5 and x6 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x14 and not x5 and not x6 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s756;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s463;

      end if;

   when s758 =>
      if ( x4 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s651;

      elsif ( not x4 and x6 and x5 and x21 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s756;

      elsif ( not x4 and x6 and x5 and x21 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y34 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s756;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and x10 and x24 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and x10 and not x24 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and x10 and not x24 and x26 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and x10 and not x24 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and not x10 and x25 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s162;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and not x10 and not x25 and x26 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and not x10 and not x25 and x26 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and x5 and not x21 and x22 and not x10 and not x25 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and x5 and not x21 and not x22 and x23 and x10 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x4 and x6 and x5 and not x21 and not x22 and x23 and not x10 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( not x4 and x6 and x5 and not x21 and not x22 and not x23 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and x5 and not x21 and not x22 and not x23 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and x5 and not x21 and not x22 and not x23 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and x5 and not x21 and not x22 and not x23 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and x9 and x8 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x4 and x6 and not x5 and x9 and x8 and not x15 and x17 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x4 and x6 and not x5 and x9 and x8 and not x15 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and x11 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and x11 and not x15 and x17 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and x11 and not x15 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and not x11 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and not x11 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and not x11 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and x10 and not x11 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and x12 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and x12 and not x15 and x17 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and x12 and not x15 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and x9 and not x8 and not x10 and not x12 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and not x9 and x10 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s989;

      elsif ( not x4 and x6 and not x5 and not x9 and x10 and not x8 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x4 and x6 and not x5 and not x9 and x10 and not x8 and not x15 and x17 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x4 and x6 and not x5 and not x9 and x10 and not x8 and not x15 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and x13 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and x13 and not x15 and x17 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and x13 and not x15 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and x8 and not x13 and not x26 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x6 and not x5 and not x9 and not x10 and not x8 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x4 and not x6 and x5 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s756;

      elsif ( not x4 and not x6 and x5 and not x7 and x8 ) = '1' then
         y5 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s756;

      elsif ( not x4 and not x6 and x5 and not x7 and not x8 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x4 and not x6 and x5 and not x7 and not x8 and not x15 and x9 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s990;

      elsif ( not x4 and not x6 and x5 and not x7 and not x8 and not x15 and x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( not x4 and not x6 and x5 and not x7 and not x8 and not x15 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s756;

      elsif ( not x4 and not x6 and not x5 and x8 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s756;

      elsif ( not x4 and not x6 and not x5 and not x8 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      else
         y5 <= '1' ;
         y23 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s756;

      end if;

   when s759 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s991;

   when s760 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s44;

   when s761 =>
      if ( x15 ) = '1' then
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s992;

      else
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s440;

      end if;

   when s762 =>
      if ( x62 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s113;

      else
         y25 <= '1' ;
         current_otherm <= s993;

      end if;

   when s763 =>
      if ( x62 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x62 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y2 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s994;

      end if;

   when s764 =>
      if ( x33 and x32 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( x33 and not x32 and x30 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s446;

      elsif ( x33 and not x32 and not x30 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x33 and not x32 and not x30 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x33 and not x32 and not x30 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 and not x30 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y53 <= '1' ;
         current_otherm <= s137;

      end if;

   when s765 =>
      if ( x32 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x32 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s766 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s995;

   when s767 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s996;

   when s768 =>
      if ( x20 ) = '1' then
         y6 <= '1' ;
         y41 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s997;

      elsif ( not x20 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s689;

      else
         y22 <= '1' ;
         current_otherm <= s361;

      end if;

   when s769 =>
      if ( x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s770 =>
      if ( x62 ) = '1' then
         y18 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s998;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s999;

      end if;

   when s771 =>
      if ( x11 ) = '1' then
         y1 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s771;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      end if;

   when s772 =>
      if ( x11 ) = '1' then
         y2 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s772;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s8;

      end if;

   when s773 =>
      if ( x62 and x64 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1000;

      elsif ( x62 and x64 and not x17 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s613;

      elsif ( x62 and not x64 and x10 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s459;

      elsif ( x62 and not x64 and not x10 and x8 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s771;

      elsif ( x62 and not x64 and not x10 and not x8 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s772;

      else
         y13 <= '1' ;
         current_otherm <= s641;

      end if;

   when s774 =>
      if ( x63 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y36 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s250;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1001;

      end if;

   when s775 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y36 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s1002;

   when s776 =>
      if ( x9 and x8 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

      elsif ( x9 and x8 and not x10 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s239;

      elsif ( x9 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x9 and x10 and x8 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x9 and x10 and x8 and not x13 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and x10 and x8 and not x13 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and x10 and x8 and not x13 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x10 and x8 and not x13 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and x10 and x8 and not x13 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x10 and not x8 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x9 and x10 and not x8 and not x3 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and x10 and not x8 and not x3 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and x10 and not x8 and not x3 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x10 and not x8 and not x3 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and x10 and not x8 and not x3 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and not x10 and x8 and x1 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x9 and not x10 and x8 and not x1 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and not x10 and x8 and not x1 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and not x10 and x8 and not x1 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and not x10 and x8 and not x1 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and not x10 and x8 and not x1 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and not x10 and not x8 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s250;

      elsif ( not x9 and not x10 and not x8 and not x15 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and not x10 and not x8 and not x15 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x9 and not x10 and not x8 and not x15 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and not x10 and not x8 and not x15 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      else
         current_otherm <= s1;

      end if;

   when s777 =>
      if ( x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s778;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

      end if;

   when s778 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s717;

   when s779 =>
         y26 <= '1' ;
         current_otherm <= s877;

   when s780 =>
      if ( x65 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1003;

      elsif ( not x65 and x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s1004;

      elsif ( not x65 and not x9 and x20 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s451;

      else
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s452;

      end if;

   when s781 =>
      if ( x64 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s337;

      else
         y42 <= '1' ;
         current_otherm <= s354;

      end if;

   when s782 =>
         y6 <= '1' ;
         current_otherm <= s337;

   when s783 =>
         y6 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s395;

   when s784 =>
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1005;

   when s785 =>
      if ( x11 and x19 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1006;

      elsif ( x11 and not x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s1007;

      else
         y29 <= '1' ;
         current_otherm <= s470;

      end if;

   when s786 =>
      if ( x20 and x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x20 and x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x20 and x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x20 and x21 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x20 and not x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1008;

      elsif ( not x20 and x21 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s532;

      elsif ( not x20 and not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s787 =>
         y22 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s382;

   when s788 =>
      if ( x64 and x20 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s469;

      elsif ( x64 and not x20 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s467;

      elsif ( not x64 and x11 ) = '1' then
         y21 <= '1' ;
         current_otherm <= s459;

      else
         y68 <= '1' ;
         current_otherm <= s743;

      end if;

   when s789 =>
      if ( x65 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s569;

      else
         y7 <= '1' ;
         current_otherm <= s371;

      end if;

   when s790 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1009;

   when s791 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1010;

   when s792 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1011;

   when s793 =>
         y24 <= '1' ;
         current_otherm <= s1012;

   when s794 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s408;

   when s795 =>
      if ( x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s796 =>
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s738;

   when s797 =>
         y22 <= '1' ;
         current_otherm <= s888;

   when s798 =>
      if ( x7 and x19 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1006;

      elsif ( x7 and not x19 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s1007;

      elsif ( not x7 and x9 and x1 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( not x7 and x9 and x1 and not x3 and x4 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s343;

      elsif ( not x7 and x9 and x1 and not x3 and x4 and not x5 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( not x7 and x9 and x1 and not x3 and x4 and not x5 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( not x7 and x9 and x1 and not x3 and not x4 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s877;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and x5 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and not x5 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and x5 and x3 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1013;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and not x5 and x3 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x1 and x2 and not x4 and not x5 and not x3 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( not x7 and x9 and not x1 and not x2 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s1014;

      end if;

   when s799 =>
      if ( x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1015;

      else
         y26 <= '1' ;
         current_otherm <= s182;

      end if;

   when s800 =>
      if ( x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s1016;

      elsif ( x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s494;

      elsif ( not x22 and x23 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1017;

      elsif ( not x22 and x23 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s494;

      elsif ( not x22 and not x23 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s497;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s493;

      end if;

   when s801 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s491;

      elsif ( not x17 and x22 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s495;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s496;

      end if;

   when s802 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1017;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s496;

      end if;

   when s803 =>
      if ( x62 ) = '1' then
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1018;

      elsif ( not x62 and x63 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      else
         y42 <= '1' ;
         current_otherm <= s354;

      end if;

   when s804 =>
      if ( x7 and x19 and x18 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and x19 and x18 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and x19 and x18 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x19 and x18 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x19 and not x18 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s560;

      elsif ( x7 and not x19 and x2 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and not x19 and x2 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and not x19 and x2 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x19 and x2 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x19 and not x2 and x18 and x3 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and not x19 and not x2 and x18 and x3 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and not x19 and not x2 and x18 and x3 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x19 and not x2 and x18 and x3 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x19 and not x2 and x18 and not x3 and x4 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s560;

      elsif ( x7 and not x19 and not x2 and x18 and not x3 and not x4 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and not x19 and not x2 and x18 and not x3 and not x4 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x7 and not x19 and not x2 and x18 and not x3 and not x4 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x19 and not x2 and x18 and not x3 and not x4 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x19 and not x2 and not x18 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s560;

      else
         y5 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1019;

      end if;

   when s805 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1020;

      else
         y6 <= '1' ;
         y14 <= '1' ;
         y25 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s1021;

      end if;

   when s806 =>
         y5 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1022;

   when s807 =>
         y2 <= '1' ;
         current_otherm <= s1023;

   when s808 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s769;

      else
         y14 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1024;

      end if;

   when s809 =>
         y6 <= '1' ;
         current_otherm <= s432;

   when s810 =>
         y38 <= '1' ;
         current_otherm <= s899;

   when s811 =>
         y39 <= '1' ;
         current_otherm <= s1025;

   when s812 =>
      if ( x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x20 and x21 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s513;

      elsif ( not x20 and x21 and not x9 and x17 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x20 and x21 and not x9 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x21 and not x9 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x21 and not x9 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x21 and not x9 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s813 =>
         y22 <= '1' ;
         current_otherm <= s171;

   when s814 =>
         y68 <= '1' ;
         current_otherm <= s743;

   when s815 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s1026;

   when s816 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y32 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s405;

   when s817 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y32 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

   when s818 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y59 <= '1' ;
         y67 <= '1' ;
         current_otherm <= s405;

   when s819 =>
      if ( x5 and x7 and x6 and x12 and x10 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x5 and x7 and x6 and x12 and not x10 and x11 and x13 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( x5 and x7 and x6 and x12 and not x10 and x11 and not x13 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x5 and x7 and x6 and x12 and not x10 and x11 and not x13 and x19 and not x14 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x5 and x7 and x6 and x12 and not x10 and x11 and not x13 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and x7 and x6 and x12 and not x10 and not x11 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y32 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s453;

      elsif ( x5 and x7 and x6 and not x12 and x10 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s413;

      elsif ( x5 and x7 and x6 and not x12 and not x10 and x11 and x14 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s101;

      elsif ( x5 and x7 and x6 and not x12 and not x10 and x11 and not x14 and x19 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x5 and x7 and x6 and not x12 and not x10 and x11 and not x14 and x19 and not x13 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x5 and x7 and x6 and not x12 and not x10 and x11 and not x14 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and x7 and x6 and not x12 and not x10 and not x11 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s514;

      elsif ( x5 and x7 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s515;

      elsif ( x5 and not x7 and x9 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s515;

      elsif ( x5 and not x7 and not x9 and x10 and x11 and x12 and x6 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( x5 and not x7 and not x9 and x10 and x11 and x12 and not x6 ) = '1' then
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      elsif ( x5 and not x7 and not x9 and x10 and x11 and not x12 and x6 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( x5 and not x7 and not x9 and x10 and x11 and not x12 and not x6 ) = '1' then
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( x5 and not x7 and not x9 and x10 and not x11 and x6 and x12 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( x5 and not x7 and not x9 and x10 and not x11 and x6 and not x12 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x5 and not x7 and not x9 and x10 and not x11 and not x6 ) = '1' then
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( x5 and not x7 and not x9 and not x10 and x11 and x12 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s517;

      elsif ( x5 and not x7 and not x9 and not x10 and x11 and x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s518;

      elsif ( x5 and not x7 and not x9 and not x10 and x11 and not x12 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y31 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s405;

      elsif ( x5 and not x7 and not x9 and not x10 and x11 and not x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y63 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s519;

      elsif ( x5 and not x7 and not x9 and not x10 and not x11 and x12 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x5 and not x7 and not x9 and not x10 and not x11 and x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s520;

      elsif ( x5 and not x7 and not x9 and not x10 and not x11 and not x12 and x6 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s521;

      elsif ( x5 and not x7 and not x9 and not x10 and not x11 and not x12 and not x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s332;

      else
         y17 <= '1' ;
         current_otherm <= s3;

      end if;

   when s820 =>
      if ( x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s821 =>
      if ( x6 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s502;

      elsif ( not x6 and x14 and x21 and x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( not x6 and x14 and x21 and not x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and x7 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and x9 and x18 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and not x9 and x19 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and x7 and x9 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s1027;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and x7 and not x9 and x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x21 and x5 and not x8 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x6 and x14 and not x21 and not x5 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1028;

      end if;

   when s822 =>
         y6 <= '1' ;
         y19 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1029;

   when s823 =>
      if ( x4 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s1004;

      else
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s1030;

      end if;

   when s824 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s206;

   when s825 =>
      if ( x3 and x21 and x26 and x27 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and x26 and x27 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and x26 and x27 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and x26 and x27 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and x26 and x27 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and x26 and not x27 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1031;

      elsif ( x3 and x21 and not x26 and x7 and x8 and x6 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and x7 and x8 and x6 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and x7 and x8 and x6 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and x8 and x6 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and x8 and x6 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and x8 and not x6 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x3 and x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and x8 and not x6 and not x9 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and x6 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and x7 and not x8 and not x6 and not x10 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and not x7 and x8 and x6 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1032;

      elsif ( x3 and x21 and not x26 and not x7 and x8 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and x6 and not x11 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x21 and not x26 and not x7 and not x8 and not x6 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( x3 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1033;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1034;

      end if;

   when s826 =>
      if ( x26 and x27 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s1035;

      elsif ( x26 and not x27 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1031;

      elsif ( not x26 and x12 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x26 and not x12 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and not x12 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and not x12 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and not x12 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s827 =>
      if ( x13 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x13 and x26 and x14 and x27 and x6 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s826;

      elsif ( not x13 and x26 and x14 and x27 and x6 and not x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( not x13 and x26 and x14 and x27 and not x6 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s825;

      elsif ( not x13 and x26 and x14 and x27 and not x6 and not x5 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s583;

      elsif ( not x13 and x26 and x14 and not x27 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s579;

      elsif ( not x13 and x26 and x14 and not x27 and not x5 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s583;

      elsif ( not x13 and x26 and not x14 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s826;

      elsif ( not x13 and x26 and not x14 and not x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( not x13 and not x26 and x27 and x14 and x5 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( not x13 and not x26 and x27 and x14 and not x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s825;

      elsif ( not x13 and not x26 and x27 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s826;

      elsif ( not x13 and not x26 and not x27 and x7 and x6 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x13 and not x26 and not x27 and x7 and x6 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x13 and not x26 and not x27 and x7 and x6 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and x6 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and x6 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and x8 and x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s556;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and x8 and not x15 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and not x8 and x16 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s556;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and x7 and not x6 and not x8 and not x16 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x13 and not x26 and not x27 and not x7 and x8 and x6 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x13 and not x26 and not x27 and not x7 and x8 and not x6 ) = '1' then
         y5 <= '1' ;
         y44 <= '1' ;
         y55 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s579;

      elsif ( not x13 and not x26 and not x27 and not x7 and not x8 and x6 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y53 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s579;

      end if;

   when s828 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1036;

   when s829 =>
      if ( x63 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x63 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s742;

      end if;

   when s830 =>
         y80 <= '1' ;
         current_otherm <= s938;

   when s831 =>
         y80 <= '1' ;
         current_otherm <= s1037;

   when s832 =>
      if ( x15 ) = '1' then
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s240;

      elsif ( not x15 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s833 =>
      if ( x63 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s1038;

      elsif ( not x63 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x63 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s834 =>
      if ( x66 and x9 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1039;

      elsif ( x66 and not x9 and x19 and x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1040;

      elsif ( x66 and not x9 and x19 and not x4 and x5 and x6 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1041;

      elsif ( x66 and not x9 and x19 and not x4 and x5 and x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1042;

      elsif ( x66 and not x9 and x19 and not x4 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s958;

      elsif ( x66 and not x9 and x19 and not x4 and not x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1043;

      elsif ( x66 and not x9 and not x19 ) = '1' then
         y4 <= '1' ;
         y20 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s1044;

      else
         y6 <= '1' ;
         current_otherm <= s239;

      end if;

   when s835 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s80;

   when s836 =>
      if ( x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1017;

      elsif ( x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s496;

      elsif ( not x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s497;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1045;

      end if;

   when s837 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s1046;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1047;

      end if;

   when s838 =>
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s806;

   when s839 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1048;

      else
         y6 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s266;

      end if;

   when s840 =>
         y6 <= '1' ;
         current_otherm <= s100;

   when s841 =>
         y6 <= '1' ;
         current_otherm <= s345;

   when s842 =>
         y9 <= '1' ;
         current_otherm <= s660;

   when s843 =>
      if ( x4 and x22 and x30 and x9 and x10 and x8 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s30;

      elsif ( x4 and x22 and x30 and x9 and x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s568;

      elsif ( x4 and x22 and x30 and x9 and not x10 and x8 ) = '1' then
         y12 <= '1' ;
         current_otherm <= s11;

      elsif ( x4 and x22 and x30 and x9 and not x10 and not x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s569;

      elsif ( x4 and x22 and x30 and not x9 and x10 and x8 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x4 and x22 and x30 and not x9 and x10 and not x8 and x27 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( x4 and x22 and x30 and not x9 and x10 and not x8 and not x27 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x22 and x30 and not x9 and not x10 and x8 ) = '1' then
         y8 <= '1' ;
         current_otherm <= s570;

      elsif ( x4 and x22 and x30 and not x9 and not x10 and not x8 and x26 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( x4 and x22 and x30 and not x9 and not x10 and not x8 and not x26 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( x4 and x22 and not x30 and x31 and x9 and x10 and x8 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( x4 and x22 and not x30 and x31 and x9 and x10 and not x8 and x21 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( x4 and x22 and not x30 and x31 and x9 and x10 and not x8 and not x21 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and x9 and x10 and not x8 and not x21 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and x9 and x10 and not x8 and not x21 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and x9 and not x10 and x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      elsif ( x4 and x22 and not x30 and x31 and x9 and not x10 and not x8 and x18 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( x4 and x22 and not x30 and x31 and x9 and not x10 and not x8 and not x18 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and x9 and not x10 and not x8 and not x18 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and x9 and not x10 and not x8 and not x18 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and x10 and x19 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and x10 and not x19 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and x10 and not x19 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and x10 and not x19 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and not x10 and x20 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and not x10 and not x20 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and not x10 and not x20 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and x8 and not x10 and not x20 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x22 and not x30 and x31 and not x9 and not x8 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( x4 and x22 and not x30 and not x31 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s572;

      elsif ( x4 and not x22 ) = '1' then
         y45 <= '1' ;
         y47 <= '1' ;
         y50 <= '1' ;
         y60 <= '1' ;
         y62 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s571;

      elsif ( not x4 and x30 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s675;

      elsif ( not x4 and not x30 and x31 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      else
         y37 <= '1' ;
         current_otherm <= s510;

      end if;

   when s844 =>
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1049;

   when s845 =>
         y33 <= '1' ;
         current_otherm <= s416;

   when s846 =>
         y9 <= '1' ;
         current_otherm <= s854;

   when s847 =>
         y9 <= '1' ;
         current_otherm <= s572;

   when s848 =>
         y9 <= '1' ;
         current_otherm <= s1050;

   when s849 =>
         y9 <= '1' ;
         current_otherm <= s1051;

   when s850 =>
         y9 <= '1' ;
         current_otherm <= s1052;

   when s851 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s585;

   when s852 =>
         y24 <= '1' ;
         current_otherm <= s203;

   when s853 =>
         y9 <= '1' ;
         current_otherm <= s770;

   when s854 =>
      if ( x62 and x33 and x32 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x62 and x33 and x32 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x62 and x33 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x33 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x33 and not x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s951;

      elsif ( x62 and not x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s951;

      elsif ( not x62 and x65 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x65 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x62 and x65 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x65 and not x15 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1053;

      end if;

   when s855 =>
         y28 <= '1' ;
         current_otherm <= s917;

   when s856 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s309;

      elsif ( not x62 and x64 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s789;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s857 =>
         y31 <= '1' ;
         current_otherm <= s122;

   when s858 =>
      if ( x64 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1054;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1055;

      end if;

   when s859 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s12;

   when s860 =>
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1056;

   when s861 =>
      if ( x62 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      else
         y15 <= '1' ;
         current_otherm <= s1057;

      end if;

   when s862 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s1058;

   when s863 =>
         y19 <= '1' ;
         y24 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1;

   when s864 =>
      if ( x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s865 =>
      if ( x6 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1059;

      elsif ( not x6 and x14 and x7 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1060;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and x9 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1061;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and x11 and x16 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and not x11 and x17 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and x11 and x9 ) = '1' then
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s84;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and x11 and not x9 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and not x11 and x9 and x15 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x14 and not x7 and x5 and not x10 and not x11 and not x9 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x6 and x14 and not x7 and not x5 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1062;

      else
         y2 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1063;

      end if;

   when s866 =>
      if ( x4 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s320;

      elsif ( not x4 and x5 and x7 and x9 and x11 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s116;

      elsif ( not x4 and x5 and x7 and x9 and not x11 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s377;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and x11 and x12 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and x11 and not x12 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and x11 and not x12 and x19 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and x11 and not x12 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and not x11 and x13 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and not x11 and not x13 and x19 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and not x11 and not x13 and x19 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x5 and x7 and not x9 and x10 and not x11 and not x13 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x5 and x7 and not x9 and not x10 and x11 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and x5 and x7 and not x9 and not x10 and not x11 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and x5 and not x7 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1063;

      elsif ( not x4 and not x5 and x6 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1063;

      elsif ( not x4 and not x5 and not x6 and x9 and x10 and x11 and x7 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x4 and not x5 and not x6 and x9 and x10 and x11 and not x7 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1064;

      elsif ( not x4 and not x5 and not x6 and x9 and x10 and not x11 and x7 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x4 and not x5 and not x6 and x9 and x10 and not x11 and not x7 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s1065;

      elsif ( not x4 and not x5 and not x6 and x9 and not x10 and x11 and x7 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s1066;

      elsif ( not x4 and not x5 and not x6 and x9 and not x10 and x11 and not x7 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1067;

      elsif ( not x4 and not x5 and not x6 and x9 and not x10 and not x11 and x7 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and not x5 and not x6 and x9 and not x10 and not x11 and not x7 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         y52 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s1068;

      elsif ( not x4 and not x5 and not x6 and not x9 and x10 and x11 and x7 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1069;

      elsif ( not x4 and not x5 and not x6 and not x9 and x10 and x11 and not x7 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and not x5 and not x6 and not x9 and x10 and not x11 and x7 ) = '1' then
         y9 <= '1' ;
         y18 <= '1' ;
         y34 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and not x5 and not x6 and not x9 and x10 and not x11 and not x7 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and not x5 and not x6 and not x9 and not x10 and x7 and x11 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s864;

      elsif ( not x4 and not x5 and not x6 and not x9 and not x10 and x7 and not x11 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      else
         y11 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s864;

      end if;

   when s867 =>
         y15 <= '1' ;
         current_otherm <= s1070;

   when s868 =>
      if ( x62 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1071;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s665;

      else
         y13 <= '1' ;
         current_otherm <= s909;

      end if;

   when s869 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s870 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s1072;

   when s871 =>
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s913;

   when s872 =>
         y40 <= '1' ;
         current_otherm <= s1073;

   when s873 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s874 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s875 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s876 =>
      if ( x30 ) = '1' then
         y5 <= '1' ;
         current_otherm <= s308;

      else
         y5 <= '1' ;
         current_otherm <= s74;

      end if;

   when s877 =>
      if ( x63 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s335;

      elsif ( not x63 and x64 ) = '1' then
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1074;

      else
         y41 <= '1' ;
         current_otherm <= s1075;

      end if;

   when s878 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1031;

   when s879 =>
         y6 <= '1' ;
         y11 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1076;

   when s880 =>
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s467;

   when s881 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1077;

   when s882 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1078;

   when s883 =>
      if ( x21 and x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1077;

      elsif ( x21 and not x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1079;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1077;

      end if;

   when s884 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s362;

   when s885 =>
         y3 <= '1' ;
         y77 <= '1' ;
         current_otherm <= s547;

   when s886 =>
      if ( x62 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1080;

      else
         y28 <= '1' ;
         current_otherm <= s306;

      end if;

   when s887 =>
      if ( x65 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1081;

      else
         y13 <= '1' ;
         current_otherm <= s225;

      end if;

   when s888 =>
      if ( x62 and x20 and x23 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( x62 and x20 and not x23 ) = '1' then
         y1 <= '1' ;
         y20 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s302;

      elsif ( x62 and not x20 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s309;

      elsif ( not x62 and x64 ) = '1' then
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1082;

      else
         y23 <= '1' ;
         current_otherm <= s169;

      end if;

   when s889 =>
         y53 <= '1' ;
         current_otherm <= s763;

   when s890 =>
      if ( x64 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x64 and x9 and not x10 and x11 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x64 and x9 and not x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s738;

      end if;

   when s891 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1083;

   when s892 =>
      if ( x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s497;

      elsif ( x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1045;

      elsif ( not x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1017;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s494;

      end if;

   when s893 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s1016;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s494;

      end if;

   when s894 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1084;

   when s895 =>
      if ( x18 and x2 and x19 and x4 and x3 and x5 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x18 and x2 and x19 and x4 and x3 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x18 and x2 and x19 and x4 and x3 and not x5 and not x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y32 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s896;

      elsif ( x18 and x2 and x19 and x4 and not x3 and x17 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and x2 and x19 and x4 and not x3 and x17 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x18 and x2 and x19 and x4 and not x3 and x17 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x2 and x19 and x4 and not x3 and not x17 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x2 and x19 and not x4 and x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s708;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and x16 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and x16 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and x16 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x2 and x19 and not x4 and not x3 and not x16 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x2 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x2 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and x2 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x2 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and x3 and x19 and x4 and x15 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x2 and x3 and x19 and x4 and x15 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x18 and not x2 and x3 and x19 and x4 and x15 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and x3 and x19 and x4 and not x15 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and x14 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and x14 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and x14 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and x3 and x19 and not x4 and not x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and x3 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x2 and x3 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x18 and not x2 and x3 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and x3 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x2 and not x3 and x19 and x4 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x2 and not x3 and x19 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x18 and not x2 and not x3 and x19 and x4 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x18 and not x2 and not x3 and x19 and not x4 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( x18 and not x2 and not x3 and not x19 and x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x18 and not x2 and not x3 and not x19 and not x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s936;

      elsif ( not x18 and x19 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( not x18 and x19 and not x2 and x4 and x3 ) = '1' then
         y23 <= '1' ;
         y27 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1086;

      elsif ( not x18 and x19 and not x2 and x4 and not x3 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s428;

      elsif ( not x18 and x19 and not x2 and not x4 and x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s83;

      elsif ( not x18 and x19 and not x2 and not x4 and not x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1087;

      else
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      end if;

   when s896 =>
      if ( x14 ) = '1' then
         y1 <= '1' ;
         current_otherm <= s107;

      elsif ( not x14 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x14 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x14 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s897 =>
         y11 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1088;

   when s898 =>
         y36 <= '1' ;
         current_otherm <= s521;

   when s899 =>
      if ( x64 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1089;

      else
         y40 <= '1' ;
         current_otherm <= s1090;

      end if;

   when s900 =>
         y4 <= '1' ;
         y31 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s657;

   when s901 =>
         y7 <= '1' ;
         current_otherm <= s475;

   when s902 =>
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s872;

   when s903 =>
         y38 <= '1' ;
         current_otherm <= s483;

   when s904 =>
      if ( x4 and x20 and x9 and x8 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x20 and x9 and x8 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x20 and x9 and x8 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x20 and x9 and x8 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x20 and x9 and not x8 and x10 ) = '1' then
         y21 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s180;

      elsif ( x4 and x20 and x9 and not x8 and not x10 ) = '1' then
         y22 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s180;

      elsif ( x4 and x20 and not x9 and x8 and x10 ) = '1' then
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s184;

      elsif ( x4 and x20 and not x9 and x8 and not x10 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s184;

      elsif ( x4 and x20 and not x9 and not x8 and x10 and x11 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s67;

      elsif ( x4 and x20 and not x9 and not x8 and x10 and not x11 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x20 and not x9 and not x8 and x10 and not x11 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x20 and not x9 and not x8 and x10 and not x11 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x20 and not x9 and not x8 and x10 and not x11 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x20 and not x9 and not x8 and not x10 and x12 ) = '1' then
         y4 <= '1' ;
         current_otherm <= s165;

      elsif ( x4 and x20 and not x9 and not x8 and not x10 and not x12 and x7 and x6 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x20 and not x9 and not x8 and not x10 and not x12 and x7 and not x6 and x5 ) = '1' then
         y20 <= '1' ;
         current_otherm <= s173;

      elsif ( x4 and x20 and not x9 and not x8 and not x10 and not x12 and x7 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and x20 and not x9 and not x8 and not x10 and not x12 and not x7 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and not x20 and x21 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x4 and not x20 and x21 and not x5 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s488;

      elsif ( x4 and not x20 and not x21 and x10 ) = '1' then
         current_otherm <= s65;

      elsif ( x4 and not x20 and not x21 and not x10 ) = '1' then
         y27 <= '1' ;
         current_otherm <= s488;

      else
         y10 <= '1' ;
         current_otherm <= s16;

      end if;

   when s905 =>
      if ( x16 and x22 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      elsif ( x16 and not x22 and x23 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s168;

      elsif ( x16 and not x22 and not x23 ) = '1' then
         y19 <= '1' ;
         current_otherm <= s166;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s738;

      end if;

   when s906 =>
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1091;

   when s907 =>
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

   when s908 =>
         y24 <= '1' ;
         current_otherm <= s117;

   when s909 =>
      if ( x62 and x17 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s888;

      elsif ( x62 and not x17 ) = '1' then
         y1 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s672;

      else
         y13 <= '1' ;
         current_otherm <= s225;

      end if;

   when s910 =>
         y5 <= '1' ;
         current_otherm <= s68;

   when s911 =>
      if ( x5 ) = '1' then
         y52 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s474;

      elsif ( not x5 and x21 and x14 and x15 and x20 and x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1077;

      elsif ( not x5 and x21 and x14 and x15 and x20 and not x13 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s108;

      elsif ( not x5 and x21 and x14 and x15 and not x20 and x13 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x5 and x21 and x14 and x15 and not x20 and not x13 and x18 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x5 and x21 and x14 and x15 and not x20 and not x13 and not x18 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and x14 and x15 and not x20 and not x13 and not x18 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and x14 and x15 and not x20 and not x13 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and x14 and x15 and not x20 and not x13 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and x14 and not x15 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s513;

      elsif ( not x5 and x21 and x14 and not x15 and x20 and not x13 ) = '1' then
         y29 <= '1' ;
         current_otherm <= s378;

      elsif ( not x5 and x21 and x14 and not x15 and not x20 and x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x5 and x21 and x14 and not x15 and not x20 and not x13 and x19 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x5 and x21 and x14 and not x15 and not x20 and not x13 and not x19 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and x14 and not x15 and not x20 and not x13 and not x19 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and x14 and not x15 and not x20 and not x13 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and x14 and not x15 and not x20 and not x13 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and x15 and x11 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and x15 and not x11 and x10 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and x15 and not x11 and x10 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and x15 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and not x15 and x12 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s204;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and not x15 and not x12 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and not x15 and not x12 and x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and x20 and x13 and not x15 and not x12 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and x20 and not x13 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and x20 and not x13 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and x20 and not x13 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and x20 and not x13 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and not x20 and x15 and x13 and x17 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x5 and x21 and not x14 and not x20 and x15 and x13 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and not x20 and x15 and x13 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and not x20 and x15 and x13 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and not x20 and x15 and x13 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and not x20 and x15 and not x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s882;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and x13 and x9 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and x13 and not x9 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and x13 and not x9 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and x13 and not x9 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and x13 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and not x13 and x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s883;

      elsif ( not x5 and x21 and not x14 and not x20 and not x15 and not x13 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s884;

      elsif ( not x5 and not x21 and x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s883;

      elsif ( not x5 and not x21 and not x7 and x20 and x14 and x15 and x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s362;

      elsif ( not x5 and not x21 and not x7 and x20 and x14 and x15 and not x13 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s768;

      elsif ( not x5 and not x21 and not x7 and x20 and x14 and not x15 and x13 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s93;

      elsif ( not x5 and not x21 and not x7 and x20 and x14 and not x15 and not x13 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s387;

      elsif ( not x5 and not x21 and not x7 and x20 and not x14 and x15 and x13 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s669;

      elsif ( not x5 and not x21 and not x7 and x20 and not x14 and x15 and not x13 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1092;

      elsif ( not x5 and not x21 and not x7 and x20 and not x14 and not x15 and x13 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

      elsif ( not x5 and not x21 and not x7 and x20 and not x14 and not x15 and not x13 ) = '1' then
         y7 <= '1' ;
         y39 <= '1' ;
         y44 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1093;

      elsif ( not x5 and not x21 and not x7 and not x20 and x13 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s93;

      elsif ( not x5 and not x21 and not x7 and not x20 and not x13 and x14 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s362;

      else
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s669;

      end if;

   when s912 =>
      if ( x5 and x9 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1094;

      elsif ( x5 and x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1095;

      elsif ( x5 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s756;

      elsif ( not x5 and x6 and x17 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x5 and x6 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      else
         y5 <= '1' ;
         y26 <= '1' ;
         y29 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s756;

      end if;

   when s913 =>
         y38 <= '1' ;
         current_otherm <= s1096;

   when s914 =>
         y3 <= '1' ;
         y19 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1097;

   when s915 =>
      if ( x6 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x5 and x7 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s890;

      elsif ( x6 and not x5 and x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y19 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s914;

      elsif ( x6 and not x5 and x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x6 and not x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      else
         y46 <= '1' ;
         current_otherm <= s890;

      end if;

   when s916 =>
      if ( x6 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x6 and not x5 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      elsif ( not x6 and x8 and x9 and x5 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s153;

      elsif ( not x6 and x8 and x9 and not x5 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y62 <= '1' ;
         y63 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and x8 and x9 and not x5 and not x7 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y57 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and x8 and not x9 and x5 ) = '1' then
         y3 <= '1' ;
         y19 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and x8 and not x9 and not x5 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y67 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and x8 and not x9 and not x5 and not x7 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y55 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and not x8 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and not x8 and not x5 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y62 <= '1' ;
         y63 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s795;

      elsif ( not x6 and not x8 and not x5 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s795;

      else
         y5 <= '1' ;
         y27 <= '1' ;
         y41 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s795;

      end if;

   when s917 =>
      if ( x63 and x20 and x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s414;

      elsif ( x63 and x20 and not x9 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s733;

      elsif ( x63 and not x20 and x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s606;

      elsif ( x63 and not x20 and not x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x63 and x21 and x22 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and x21 and not x22 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      elsif ( not x63 and x21 and not x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and not x21 and x23 ) = '1' then
         y70 <= '1' ;
         current_otherm <= s263;

      else
         current_otherm <= s1;

      end if;

   when s918 =>
         y34 <= '1' ;
         current_otherm <= s178;

   when s919 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1098;

   when s920 =>
      if ( x7 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s642;

      elsif ( not x7 and x19 and x23 and x4 and x5 and x3 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and x4 and x5 and x3 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and x4 and x5 and x3 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and x4 and x5 and x3 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and x4 and x5 and not x3 and x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( not x7 and x19 and x23 and x4 and x5 and not x3 and not x12 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and x4 and x5 and not x3 and not x12 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and x4 and x5 and not x3 and not x12 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and x4 and x5 and not x3 and not x12 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and x4 and not x5 and x3 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s856;

      elsif ( not x7 and x19 and x23 and x4 and not x5 and not x3 and x11 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( not x7 and x19 and x23 and x4 and not x5 and not x3 and not x11 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and x4 and not x5 and not x3 and not x11 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and x4 and not x5 and not x3 and not x11 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and x4 and not x5 and not x3 and not x11 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and not x4 and x3 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s621;

      elsif ( not x7 and x19 and x23 and not x4 and x3 and not x5 and x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( not x7 and x19 and x23 and not x4 and x3 and not x5 and not x13 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and not x4 and x3 and not x5 and not x13 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x7 and x19 and x23 and not x4 and x3 and not x5 and not x13 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and not x4 and x3 and not x5 and not x13 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x19 and x23 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( not x7 and x19 and not x23 and x22 and x4 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1099;

      elsif ( not x7 and x19 and not x23 and x22 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x7 and x19 and not x23 and x22 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s337;

      elsif ( not x7 and x19 and not x23 and not x22 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s856;

      else
         y1 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s1100;

      end if;

   when s921 =>
         y45 <= '1' ;
         current_otherm <= s114;

   when s922 =>
      if ( x6 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x6 and x22 and x23 and x4 and x3 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x6 and x22 and x23 and x4 and x3 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x6 and x22 and x23 and x4 and x3 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and x4 and x3 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and x5 and x15 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and x5 and not x15 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and x5 and not x15 and x21 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and x5 and not x15 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and not x5 and x16 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and not x5 and not x16 and x21 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and not x5 and not x16 and x21 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and x4 and not x3 and not x5 and not x16 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and not x4 and x5 and x3 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and not x4 and x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and x22 and x23 and not x4 and not x5 and x3 ) = '1' then
         y51 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s1;

      elsif ( not x6 and x22 and x23 and not x4 and not x5 and not x3 ) = '1' then
         y1 <= '1' ;
         y19 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and x22 and not x23 and x9 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and x22 and not x23 and not x9 and x3 and x5 and x4 ) = '1' then
         y42 <= '1' ;
         current_otherm <= s354;

      elsif ( not x6 and x22 and not x23 and not x9 and x3 and x5 and not x4 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( not x6 and x22 and not x23 and not x9 and x3 and not x5 and x4 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x22 and not x23 and not x9 and x3 and not x5 and not x4 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( not x6 and x22 and not x23 and not x9 and not x3 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1100;

      elsif ( not x6 and x22 and not x23 and not x9 and not x3 and not x7 and x4 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1101;

      elsif ( not x6 and x22 and not x23 and not x9 and not x3 and not x7 and x4 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and x22 and not x23 and not x9 and not x3 and not x7 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y27 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and not x22 and x23 and x9 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s401;

      elsif ( not x6 and not x22 and x23 and not x9 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1100;

      elsif ( not x6 and not x22 and not x23 and x3 and x5 and x4 ) = '1' then
         y31 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and not x22 and not x23 and x3 and x5 and not x4 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x6 and not x22 and not x23 and x3 and not x5 and x4 ) = '1' then
         y30 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s302;

      elsif ( not x6 and not x22 and not x23 and x3 and not x5 and not x4 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s121;

      elsif ( not x6 and not x22 and not x23 and not x3 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y8 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1100;

      else
         y1 <= '1' ;
         y27 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s302;

      end if;

   when s923 =>
         y6 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1102;

   when s924 =>
      if ( x10 and x2 and x3 and x4 and x9 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and x2 and x3 and x4 and x9 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and x2 and x3 and x4 and x9 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x2 and x3 and x4 and x9 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x2 and x3 and x4 and not x9 and x8 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( x10 and x2 and x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and x2 and x3 and not x4 and x9 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s681;

      elsif ( x10 and x2 and x3 and not x4 and x9 and not x6 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x10 and x2 and x3 and not x4 and not x9 and x8 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x10 and x2 and x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and x2 and not x3 and x4 and x9 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s894;

      elsif ( x10 and x2 and not x3 and x4 and not x9 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( x10 and x2 and not x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and x2 and not x3 and not x4 and x9 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x10 and x2 and not x3 and not x4 and x9 and not x13 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x2 and not x3 and not x4 and x9 and not x13 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x2 and not x3 and not x4 and not x9 and x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and x2 and not x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and not x2 and x4 and x3 and x9 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x10 and not x2 and x4 and x3 and x9 and not x14 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x2 and x4 and x3 and x9 and not x14 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x2 and x4 and x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1104;

      elsif ( x10 and not x2 and x4 and x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and not x2 and x4 and not x3 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x10 and not x2 and x4 and not x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and not x2 and x4 and not x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and not x2 and not x4 and x9 and x3 and x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x10 and not x2 and not x4 and x9 and x3 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x10 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x2 and not x4 and x9 and x3 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x2 and not x4 and x9 and not x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( x10 and not x2 and not x4 and not x9 and x8 and x3 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and not x2 and not x4 and not x9 and x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x10 and not x2 and not x4 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y36 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1105;

      end if;

   when s925 =>
      if ( x3 and x4 and x6 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s726;

      elsif ( x3 and x4 and not x6 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s1025;

      elsif ( x3 and not x4 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1106;

      elsif ( not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s506;

      else
         y20 <= '1' ;
         current_otherm <= s173;

      end if;

   when s926 =>
      if ( x4 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s877;

      elsif ( x4 and not x3 and x5 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( x4 and not x3 and x5 and not x15 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x4 and not x3 and x5 and not x15 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x4 and not x3 and x5 and not x15 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and not x3 and x5 and not x15 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and not x3 and not x5 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( x4 and not x3 and not x5 and not x17 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x4 and not x3 and not x5 and not x17 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x4 and not x3 and not x5 and not x17 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x4 and not x3 and not x5 and not x17 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x5 and x3 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1013;

      elsif ( not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x4 and not x5 and x3 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x4 and not x5 and x3 and not x16 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x4 and not x5 and x3 and not x16 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x4 and not x5 and x3 and not x16 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and not x5 and x3 and not x16 and not x22 ) = '1' then
         current_otherm <= s1;

      else
         y38 <= '1' ;
         current_otherm <= s483;

      end if;

   when s927 =>
      if ( x1 and x4 and x5 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( x1 and x4 and not x5 and x3 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x1 and x4 and not x5 and not x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x1 and x4 and not x5 and not x3 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x1 and x4 and not x5 and not x3 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x1 and not x4 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      else
         y26 <= '1' ;
         current_otherm <= s649;

      end if;

   when s928 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1107;

   when s929 =>
         y6 <= '1' ;
         y9 <= '1' ;
         y25 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1108;

   when s930 =>
         y40 <= '1' ;
         current_otherm <= s1109;

   when s931 =>
         y40 <= '1' ;
         current_otherm <= s1110;

   when s932 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s1111;

   when s933 =>
         y4 <= '1' ;
         y20 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1112;

   when s934 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s707;

   when s935 =>
         y11 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s560;

   when s936 =>
         y21 <= '1' ;
         y29 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1113;

   when s937 =>
      if ( x21 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x21 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x21 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s409;

      elsif ( not x21 and not x22 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x22 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x22 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s938 =>
      if ( x21 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x21 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( x21 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and x20 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x21 and x22 and not x20 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x20 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and x22 and not x20 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x22 and not x20 and not x6 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and not x22 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x22 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x21 and not x22 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s939 =>
      if ( x63 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s983;

      else
         y37 <= '1' ;
         current_otherm <= s428;

      end if;

   when s940 =>
      if ( x7 and x13 and x8 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and x8 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and x8 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and x8 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and x8 and not x9 and x11 and x10 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and x8 and not x9 and x11 and x10 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and x8 and not x9 and x11 and x10 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and x8 and not x9 and x11 and x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and x8 and not x9 and x11 and not x10 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s504;

      elsif ( x7 and x13 and x8 and not x9 and not x11 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1114;

      elsif ( x7 and x13 and x8 and not x9 and not x11 and not x10 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and x8 and not x9 and not x11 and not x10 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and x8 and not x9 and not x11 and not x10 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and x8 and not x9 and not x11 and not x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and not x9 and x18 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and x10 and not x11 and x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( x7 and x13 and not x8 and x6 and x10 and not x11 and not x9 and x17 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x7 and x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and x11 and x9 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1115;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and x11 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and not x11 and x9 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x13 and not x8 and x6 and not x10 and not x11 and not x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x7 and x13 and not x8 and not x6 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s1023;

      elsif ( x7 and not x13 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1116;

      else
         y2 <= '1' ;
         current_otherm <= s1117;

      end if;

   when s941 =>
      if ( x5 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s692;

      elsif ( not x5 and x6 and x8 and x9 and x12 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x5 and x6 and x8 and x9 and not x12 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and x11 and x16 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and x11 and not x16 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and x11 and not x16 and x14 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and x11 and not x16 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and not x11 and x15 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and not x11 and not x15 and x14 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and not x11 and not x15 and x14 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and x8 and not x9 and x10 and not x11 and not x15 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x6 and x8 and not x9 and not x10 and x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         y51 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and x6 and x8 and not x9 and not x10 and not x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and x6 and not x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1116;

      elsif ( not x5 and not x6 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1116;

      elsif ( not x5 and not x6 and not x7 and x9 and x10 and x11 and x8 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s993;

      elsif ( not x5 and not x6 and not x7 and x9 and x10 and x11 and not x8 ) = '1' then
         y32 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and not x6 and not x7 and x9 and x10 and not x11 and x8 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( not x5 and not x6 and not x7 and x9 and x10 and not x11 and not x8 ) = '1' then
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and not x6 and not x7 and x9 and not x10 and x11 and x8 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( not x5 and not x6 and not x7 and x9 and not x10 and x11 and not x8 ) = '1' then
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s158;

      elsif ( not x5 and not x6 and not x7 and x9 and not x10 and not x11 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( not x5 and not x6 and not x7 and x9 and not x10 and not x11 and not x8 ) = '1' then
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s380;

      elsif ( not x5 and not x6 and not x7 and not x9 and x10 and x11 and x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s151;

      elsif ( not x5 and not x6 and not x7 and not x9 and x10 and x11 and not x8 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and not x6 and not x7 and not x9 and x10 and not x11 and x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and not x6 and not x7 and not x9 and x10 and not x11 and not x8 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and not x6 and not x7 and not x9 and not x10 and x8 and x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s769;

      elsif ( not x5 and not x6 and not x7 and not x9 and not x10 and x8 and not x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s769;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s769;

      end if;

   when s942 =>
      if ( x12 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x12 and x17 and x8 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x12 and x17 and not x8 and x9 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x12 and x17 and not x8 and not x9 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s943 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s145;

   when s944 =>
      if ( x6 and x8 and x27 and x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s579;

      elsif ( x6 and x8 and x27 and not x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s579;

      elsif ( x6 and x8 and not x27 and x7 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x6 and x8 and not x27 and not x7 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( x6 and not x8 and x27 and x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s579;

      elsif ( x6 and not x8 and x27 and not x7 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s579;

      elsif ( x6 and not x8 and not x27 and x7 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      elsif ( x6 and not x8 and not x27 and not x7 ) = '1' then
         y18 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s580;

      elsif ( not x6 and x7 and x27 and x8 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( not x6 and x7 and x27 and not x8 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( not x6 and x7 and not x27 and x13 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x6 and x7 and not x27 and x13 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x6 and x7 and not x27 and x13 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x7 and not x27 and x13 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x7 and not x27 and x13 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x7 and not x27 and not x13 and x3 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x6 and x7 and not x27 and not x13 and x3 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x6 and x7 and not x27 and not x13 and x3 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x7 and not x27 and not x13 and x3 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x7 and not x27 and not x13 and x3 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x7 and not x27 and not x13 and not x3 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s581;

      elsif ( not x6 and not x7 and x27 ) = '1' then
         y5 <= '1' ;
         y32 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s579;

      elsif ( not x6 and not x7 and not x27 and x8 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         y32 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s579;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s579;

      end if;

   when s945 =>
         y7 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1;

   when s946 =>
         y2 <= '1' ;
         y15 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s1118;

   when s947 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

   when s948 =>
      if ( x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s889;

      elsif ( not x10 and x11 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s727;

      else
         y29 <= '1' ;
         current_otherm <= s887;

      end if;

   when s949 =>
      if ( x63 ) = '1' then
         y21 <= '1' ;
         y28 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1119;

      else
         y47 <= '1' ;
         y52 <= '1' ;
         y61 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s25;

      end if;

   when s950 =>
         y33 <= '1' ;
         current_otherm <= s321;

   when s951 =>
      if ( x33 and x32 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s952;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s952;

      end if;

   when s952 =>
      if ( x33 and x32 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x33 and x32 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and x32 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x33 and not x32 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      else
         y9 <= '1' ;
         current_otherm <= s43;

      end if;

   when s953 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1120;

   when s954 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s418;

   when s955 =>
      if ( x64 and x66 ) = '1' then
         y18 <= '1' ;
         y27 <= '1' ;
         y29 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s1121;

      elsif ( x64 and not x66 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s1122;

      elsif ( not x64 and x14 and x31 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s364;

      elsif ( not x64 and x14 and x31 and not x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s662;

      elsif ( not x64 and x14 and not x31 and x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s290;

      elsif ( not x64 and x14 and not x31 and not x30 ) = '1' then
         y3 <= '1' ;
         current_otherm <= s379;

      else
         y25 <= '1' ;
         current_otherm <= s939;

      end if;

   when s956 =>
      if ( x7 and x9 and x8 and x3 and x2 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x7 and x9 and x8 and x3 and x2 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x7 and x9 and x8 and x3 and x2 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x9 and x8 and x3 and x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x9 and x8 and x3 and not x2 and x4 and x17 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( x7 and x9 and x8 and x3 and not x2 and x4 and not x17 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x7 and x9 and x8 and x3 and not x2 and x4 and not x17 and x1 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x9 and x8 and x3 and not x2 and x4 and not x17 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x9 and x8 and x3 and not x2 and not x4 and x16 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( x7 and x9 and x8 and x3 and not x2 and not x4 and not x16 and x1 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x7 and x9 and x8 and x3 and not x2 and not x4 and not x16 and x1 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x9 and x8 and x3 and not x2 and not x4 and not x16 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and x9 and x8 and not x3 and x4 and x2 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( x7 and x9 and x8 and not x3 and x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s276;

      elsif ( x7 and x9 and x8 and not x3 and not x4 and x2 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s321;

      elsif ( x7 and x9 and x8 and not x3 and not x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and x9 and not x8 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s1123;

      elsif ( x7 and not x9 and x11 and x2 and x4 and x8 and x3 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( x7 and not x9 and x11 and x2 and x4 and x8 and not x3 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( x7 and not x9 and x11 and x2 and x4 and not x8 and x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and x2 and x4 and not x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and x2 and not x4 and x8 and x3 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x7 and not x9 and x11 and x2 and not x4 and x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and x2 and not x4 and not x8 and x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and x2 and not x4 and not x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and not x2 and x8 and x3 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x7 and not x9 and x11 and not x2 and x8 and x3 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x7 and not x9 and x11 and not x2 and x8 and x3 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x9 and x11 and not x2 and x8 and x3 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x7 and not x9 and x11 and not x2 and x8 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and not x2 and x8 and not x3 and not x4 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and not x2 and not x8 and x4 and x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and not x2 and not x8 and x4 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and x11 and not x2 and not x8 and not x4 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y50 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s1103;

      elsif ( x7 and not x9 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s1123;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s1124;

      end if;

   when s957 =>
         y9 <= '1' ;
         current_otherm <= s43;

   when s958 =>
      if ( x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s959 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1043;

   when s960 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1041;

   when s961 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1042;

   when s962 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s958;

   when s963 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y55 <= '1' ;
         y58 <= '1' ;
         y69 <= '1' ;
         current_otherm <= s1125;

   when s964 =>
      if ( x18 and x8 and x7 ) = '1' then
         y5 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s965;

      elsif ( x18 and x8 and not x7 and x9 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x18 and x8 and not x7 and x9 and not x14 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x18 and x8 and not x7 and x9 and not x14 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x18 and x8 and not x7 and x9 and not x14 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x8 and not x7 and x9 and not x14 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x8 and not x7 and not x9 and x12 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x18 and x8 and not x7 and not x9 and not x12 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x18 and x8 and not x7 and not x9 and not x12 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x18 and x8 and not x7 and not x9 and not x12 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and x8 and not x7 and not x9 and not x12 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x8 and x9 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s966;

      elsif ( x18 and not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( x18 and not x8 and not x9 and x7 and x13 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x18 and not x8 and not x9 and x7 and not x13 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x18 and not x8 and not x9 and x7 and not x13 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x18 and not x8 and not x9 and x7 and not x13 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x8 and not x9 and x7 and not x13 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x18 and not x8 and not x9 and not x7 ) = '1' then
         y69 <= '1' ;
         current_otherm <= s535;

      else
         y5 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s968;

      end if;

   when s965 =>
         y5 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1126;

   when s966 =>
         y5 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1127;

   when s967 =>
      if ( x65 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x65 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x65 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x65 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x65 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x65 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s968 =>
      if ( x8 and x7 ) = '1' then
         y5 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s965;

      elsif ( x8 and not x7 and x9 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x8 and not x7 and x9 and not x14 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x8 and not x7 and x9 and not x14 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x8 and not x7 and x9 and not x14 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x7 and x9 and not x14 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x7 and not x9 and x12 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x8 and not x7 and not x9 and not x12 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x8 and not x7 and not x9 and not x12 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x8 and not x7 and not x9 and not x12 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x7 and not x9 and not x12 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x9 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s966;

      elsif ( not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

      elsif ( not x8 and not x9 and x7 and x13 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x8 and not x9 and x7 and not x13 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x8 and not x9 and x7 and not x13 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x8 and not x9 and x7 and not x13 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and not x9 and x7 and not x13 and not x15 ) = '1' then
         current_otherm <= s1;

      else
         y69 <= '1' ;
         current_otherm <= s535;

      end if;

   when s969 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s742;

   when s970 =>
      if ( x65 and x18 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s971;

      elsif ( x65 and x18 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and x18 and not x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x65 and not x18 ) = '1' then
         y5 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s972;

      else
         y9 <= '1' ;
         current_otherm <= s1128;

      end if;

   when s971 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

   when s972 =>
      if ( x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s971;

      elsif ( x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y26 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s742;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      end if;

   when s973 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y52 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s742;

   when s974 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s742;

   when s975 =>
      if ( x18 and x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y55 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s976;

      elsif ( x18 and x8 and x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x18 and x8 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y47 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s977;

      elsif ( x18 and x8 and not x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x18 and not x8 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y66 <= '1' ;
         y67 <= '1' ;
         current_otherm <= s978;

      elsif ( x18 and not x8 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s979;

      elsif ( x18 and not x8 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      else
         y5 <= '1' ;
         y19 <= '1' ;
         y23 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s980;

      end if;

   when s976 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y66 <= '1' ;
         y67 <= '1' ;
         current_otherm <= s1129;

   when s977 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s1130;

   when s978 =>
         y3 <= '1' ;
         y26 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s742;

   when s979 =>
         y3 <= '1' ;
         y26 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s742;

   when s980 =>
      if ( x8 and x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y55 <= '1' ;
         y65 <= '1' ;
         current_otherm <= s976;

      elsif ( x8 and x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( x8 and not x9 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y47 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s977;

      elsif ( x8 and not x9 and not x7 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      elsif ( not x8 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y66 <= '1' ;
         y67 <= '1' ;
         current_otherm <= s978;

      elsif ( not x8 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y56 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s979;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s742;

      end if;

   when s981 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1131;

   when s982 =>
      if ( x63 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x63 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s983 =>
      if ( x63 and x2 and x3 and x4 and x9 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x2 and x3 and x4 and x9 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x2 and x3 and x4 and x9 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x2 and x3 and x4 and x9 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x2 and x3 and x4 and not x9 and x8 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( x63 and x2 and x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and x2 and x3 and not x4 and x9 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s681;

      elsif ( x63 and x2 and x3 and not x4 and x9 and not x6 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x63 and x2 and x3 and not x4 and not x9 and x8 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x63 and x2 and x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and x2 and not x3 and x4 and x9 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s894;

      elsif ( x63 and x2 and not x3 and x4 and not x9 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( x63 and x2 and not x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and x2 and not x3 and not x4 and x9 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x63 and x2 and not x3 and not x4 and x9 and not x13 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x2 and not x3 and not x4 and x9 and not x13 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and x2 and not x3 and not x4 and not x9 and x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and x2 and not x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and not x2 and x4 and x3 and x9 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x63 and not x2 and x4 and x3 and x9 and not x14 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x2 and x4 and x3 and x9 and not x14 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x2 and x4 and x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1104;

      elsif ( x63 and not x2 and x4 and x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and not x2 and x4 and not x3 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x63 and not x2 and x4 and not x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and not x2 and x4 and not x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and not x2 and not x4 and x9 and x3 and x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x63 and not x2 and not x4 and x9 and x3 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x63 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x2 and not x4 and x9 and x3 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x63 and not x2 and not x4 and x9 and not x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( x63 and not x2 and not x4 and not x9 and x8 and x3 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and not x2 and not x4 and not x9 and x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x63 and not x2 and not x4 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x63 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x63 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s984 =>
         y5 <= '1' ;
         y19 <= '1' ;
         y30 <= '1' ;
         y39 <= '1' ;
         y60 <= '1' ;
         current_otherm <= s1132;

   when s985 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1133;

   when s986 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s967;

   when s987 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1134;

   when s988 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s1135;

   when s989 =>
      if ( x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s778;

      elsif ( not x15 and x17 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      end if;

   when s990 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1136;

   when s991 =>
      if ( x3 and x12 and x11 and x14 and x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s460;

      elsif ( x3 and x12 and x11 and x14 and x15 and not x13 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( x3 and x12 and x11 and x14 and not x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s460;

      elsif ( x3 and x12 and x11 and x14 and not x15 and not x13 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( x3 and x12 and x11 and not x14 and x13 and x15 and x9 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s425;

      elsif ( x3 and x12 and x11 and not x14 and x13 and x15 and not x9 and x8 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x3 and x12 and x11 and not x14 and x13 and x15 and not x9 and x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x12 and x11 and not x14 and x13 and x15 and not x9 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x12 and x11 and not x14 and x13 and not x15 and x10 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s425;

      elsif ( x3 and x12 and x11 and not x14 and x13 and not x15 and not x10 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x3 and x12 and x11 and not x14 and x13 and not x15 and not x10 and x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x12 and x11 and not x14 and x13 and not x15 and not x10 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x12 and x11 and not x14 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x3 and x12 and x11 and not x14 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x3 and x12 and x11 and not x14 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x12 and x11 and not x14 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x12 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1137;

      elsif ( x3 and not x12 and x6 and x11 and x13 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s460;

      elsif ( x3 and not x12 and x6 and x11 and x13 and x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s460;

      elsif ( x3 and not x12 and x6 and x11 and x13 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s460;

      elsif ( x3 and not x12 and x6 and x11 and x13 and not x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1138;

      elsif ( x3 and not x12 and x6 and x11 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x3 and not x12 and x6 and x11 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x3 and not x12 and x6 and x11 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and not x12 and x6 and x11 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and not x12 and x6 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1139;

      elsif ( x3 and not x12 and not x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1137;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1140;

      end if;

   when s992 =>
      if ( x5 and x7 and x9 and x8 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( x5 and x7 and x9 and not x8 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      elsif ( x5 and x7 and not x9 and x8 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s280;

      elsif ( x5 and x7 and not x9 and not x8 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( x5 and not x7 and x8 and x9 and x3 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x5 and not x7 and x8 and x9 and not x3 and x10 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x5 and not x7 and x8 and x9 and not x3 and not x10 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s153;

      elsif ( x5 and not x7 and x8 and not x9 and x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( x5 and not x7 and x8 and not x9 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s281;

      elsif ( x5 and not x7 and x8 and not x9 and not x3 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s275;

      elsif ( x5 and not x7 and not x8 and x3 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s275;

      elsif ( x5 and not x7 and not x8 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s275;

      elsif ( x5 and not x7 and not x8 and not x3 and x9 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s275;

      elsif ( x5 and not x7 and not x8 and not x3 and x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s275;

      elsif ( x5 and not x7 and not x8 and not x3 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s275;

      elsif ( not x5 and x8 and x9 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s275;

      elsif ( not x5 and x8 and not x9 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s275;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s275;

      end if;

   when s993 =>
      if ( x64 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x64 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x64 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y72 <= '1' ;
         current_otherm <= s538;

      end if;

   when s994 =>
         y2 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1141;

   when s995 =>
      if ( x8 ) = '1' then
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1142;

      elsif ( not x8 and x32 ) = '1' then
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1142;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      end if;

   when s996 =>
         y8 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1143;

   when s997 =>
         y29 <= '1' ;
         current_otherm <= s1144;

   when s998 =>
         y8 <= '1' ;
         y9 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s1145;

   when s999 =>
         y9 <= '1' ;
         current_otherm <= s1146;

   when s1000 =>
         y22 <= '1' ;
         current_otherm <= s361;

   when s1001 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y59 <= '1' ;
         y69 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s1147;

   when s1002 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s250;

   when s1003 =>
      if ( x10 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x2 and x3 and x4 and x5 and x1 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x10 and not x2 and x3 and x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and x3 and x4 and not x5 and x1 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x10 and not x2 and x3 and x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and x3 and not x4 and x5 and x1 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x10 and not x2 and x3 and not x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and x3 and not x4 and not x5 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and x3 and not x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and not x3 and x4 and x5 and x1 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x10 and not x2 and not x3 and x4 and x5 and x1 and not x6 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x10 and not x2 and not x3 and x4 and x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s340;

      elsif ( x10 and not x2 and not x3 and x4 and x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and not x3 and x4 and not x5 and x1 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x10 and not x2 and not x3 and x4 and not x5 and x1 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x10 and not x2 and not x3 and x4 and not x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and not x3 and x4 and not x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and not x3 and not x4 and x1 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and not x3 and not x4 and x1 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x10 and not x2 and not x3 and not x4 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y32 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( not x10 and x11 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s780;

      else
         y29 <= '1' ;
         current_otherm <= s1144;

      end if;

   when s1004 =>
      if ( x63 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s1007;

      else
         y2 <= '1' ;
         current_otherm <= s24;

      end if;

   when s1005 =>
      if ( x7 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s1148;

      elsif ( not x7 and x8 and x20 and x14 and x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s668;

      elsif ( not x7 and x8 and x20 and x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y42 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s855;

      elsif ( not x7 and x8 and x20 and not x14 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1149;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and x14 and x15 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and x14 and not x15 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and x14 and not x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and x15 and x17 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and x15 and x17 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and not x15 and x9 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and not x15 and x9 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and x13 and not x21 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and x15 and x18 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and x15 and x18 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and not x15 and x19 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and not x15 and x19 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and not x13 and x14 and not x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and x21 and x15 and x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and x21 and x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s882;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and x21 and not x15 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s884;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x8 and not x20 and not x13 and not x14 and not x21 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y6 <= '1' ;
         y9 <= '1' ;
         y25 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1150;

      end if;

   when s1006 =>
      if ( x9 and x1 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( x9 and x1 and not x3 and x4 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s343;

      elsif ( x9 and x1 and not x3 and x4 and not x5 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x9 and x1 and not x3 and x4 and not x5 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x9 and x1 and not x3 and x4 and not x5 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x9 and x1 and not x3 and not x4 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( x9 and not x1 and x2 and x4 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s877;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and x5 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and x5 and not x15 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and not x5 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x1 and x2 and x4 and not x3 and not x5 and not x17 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x1 and x2 and not x4 and x5 and x3 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1013;

      elsif ( x9 and not x1 and x2 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( x9 and not x1 and x2 and not x4 and not x5 and x3 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x1 and x2 and not x4 and not x5 and x3 and not x16 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x1 and x2 and not x4 and not x5 and not x3 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      elsif ( x9 and not x1 and not x2 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y8 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s1014;

      end if;

   when s1007 =>
      if ( x65 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1151;

      else
         y15 <= '1' ;
         current_otherm <= s149;

      end if;

   when s1008 =>
         y54 <= '1' ;
         current_otherm <= s108;

   when s1009 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1152;

   when s1010 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1153;

   when s1011 =>
         y2 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s1154;

   when s1012 =>
      if ( x64 and x12 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( x64 and not x12 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x12 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x12 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x12 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         y25 <= '1' ;
         current_otherm <= s1122;

      end if;

   when s1013 =>
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s1155;

   when s1014 =>
      if ( x1 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( x1 and not x3 and x4 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s343;

      elsif ( x1 and not x3 and x4 and not x5 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x1 and not x3 and x4 and not x5 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x1 and not x3 and x4 and not x5 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x1 and not x3 and not x4 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( not x1 and x2 and x4 and x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s877;

      elsif ( not x1 and x2 and x4 and not x3 and x5 and x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x1 and x2 and x4 and not x3 and x5 and not x15 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x1 and x2 and x4 and not x3 and x5 and not x15 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x1 and x2 and x4 and not x3 and not x5 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x1 and x2 and x4 and not x3 and not x5 and not x17 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x1 and x2 and x4 and not x3 and not x5 and not x17 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x1 and x2 and not x4 and x5 and x3 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1013;

      elsif ( not x1 and x2 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x1 and x2 and not x4 and not x5 and x3 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

      elsif ( not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x1 and x2 and not x4 and not x5 and x3 and not x16 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x1 and x2 and not x4 and not x5 and x3 and not x16 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x1 and x2 and not x4 and not x5 and not x3 ) = '1' then
         y38 <= '1' ;
         current_otherm <= s483;

      else
         y26 <= '1' ;
         current_otherm <= s649;

      end if;

   when s1015 =>
      if ( x21 and x26 and x27 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and x26 and x27 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and x26 and x27 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and x26 and x27 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and x26 and x27 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and x26 and not x27 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1031;

      elsif ( x21 and not x26 and x7 and x8 and x6 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and x7 and x8 and x6 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and x7 and x8 and x6 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and x8 and x6 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and x8 and x6 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and x8 and not x6 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and x8 and not x6 and not x9 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and x8 and not x6 and not x9 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and not x8 and x6 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( x21 and not x26 and x7 and not x8 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and not x8 and not x6 and not x10 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and x7 and not x8 and not x6 and not x10 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and not x7 and x8 and x6 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1032;

      elsif ( x21 and not x26 and not x7 and x8 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x21 and not x26 and not x7 and not x8 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and not x7 and not x8 and x6 and not x11 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and not x7 and not x8 and x6 and not x11 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x21 and not x26 and not x7 and not x8 and not x6 ) = '1' then
         y49 <= '1' ;
         current_otherm <= s256;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1033;

      end if;

   when s1016 =>
      if ( x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_otherm <= s193;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y67 <= '1' ;
         y68 <= '1' ;
         current_otherm <= s1156;

      end if;

   when s1017 =>
      if ( x16 and x22 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s557;

      elsif ( x16 and x22 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s251;

      elsif ( x16 and not x22 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( not x16 and x22 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s252;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s344;

      end if;

   when s1018 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y12 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1157;

   when s1019 =>
      if ( x6 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1158;

      elsif ( x6 and x19 and not x18 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x6 and not x19 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1158;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and x3 and x5 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and x3 and not x5 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y32 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s896;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and not x3 and x17 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and not x3 and x17 and not x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s708;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and not x3 and x16 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and not x3 and x16 and not x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and x2 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and x2 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and x2 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and x2 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and x4 and x15 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and x4 and x15 and not x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and not x4 and x14 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and not x4 and x14 and not x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and x3 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x18 and not x2 and not x3 and x19 and x4 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and not x2 and not x3 and x19 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( not x6 and x10 and x18 and not x2 and not x3 and x19 and not x4 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( not x6 and x10 and x18 and not x2 and not x3 and not x19 and x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( not x6 and x10 and x18 and not x2 and not x3 and not x19 and not x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s936;

      elsif ( not x6 and x10 and not x18 and x19 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( not x6 and x10 and not x18 and x19 and not x2 and x4 and x3 ) = '1' then
         y23 <= '1' ;
         y27 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1086;

      elsif ( not x6 and x10 and not x18 and x19 and not x2 and x4 and not x3 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s428;

      elsif ( not x6 and x10 and not x18 and x19 and not x2 and not x4 and x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s83;

      elsif ( not x6 and x10 and not x18 and x19 and not x2 and not x4 and not x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1087;

      elsif ( not x6 and x10 and not x18 and not x19 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      else
         y5 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         y30 <= '1' ;
         y35 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s895;

      end if;

   when s1020 =>
      if ( x14 and x21 and x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( x14 and x21 and not x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x14 and not x21 and x5 and x8 and x7 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and x9 and x18 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and x9 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and not x9 and x19 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x21 and x5 and x8 and not x7 and not x9 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x21 and x5 and not x8 and x7 and x9 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s1027;

      elsif ( x14 and not x21 and x5 and not x8 and x7 and not x9 and x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x21 and x5 and not x8 and x7 and not x9 and not x20 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x21 and x5 and not x8 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( x14 and not x21 and not x5 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1028;

      end if;

   when s1021 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s805;

   when s1022 =>
      if ( x10 and x18 and x2 and x19 and x4 and x3 and x5 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x10 and x18 and x2 and x19 and x4 and x3 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x10 and x18 and x2 and x19 and x4 and x3 and not x5 and not x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y32 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s896;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and x17 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and x17 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and x17 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and x2 and x19 and x4 and not x3 and not x17 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and x2 and x19 and not x4 and x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s708;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and x16 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and x16 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and x16 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and x2 and x19 and not x4 and not x3 and not x16 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and x2 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and x2 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and x2 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and x2 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and x15 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and x15 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and x15 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and x3 and x19 and x4 and not x15 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and x14 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and x14 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and x14 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and x3 and x19 and not x4 and not x14 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and x3 and not x19 and x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and not x2 and x3 and not x19 and x11 and not x12 and x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x10 and x18 and not x2 and x3 and not x19 and x11 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and x3 and not x19 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x18 and not x2 and not x3 and x19 and x4 and x5 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and not x2 and not x3 and x19 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      elsif ( x10 and x18 and not x2 and not x3 and x19 and x4 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s560;

      elsif ( x10 and x18 and not x2 and not x3 and x19 and not x4 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s115;

      elsif ( x10 and x18 and not x2 and not x3 and not x19 and x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x10 and x18 and not x2 and not x3 and not x19 and not x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s936;

      elsif ( x10 and not x18 and x19 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      elsif ( x10 and not x18 and x19 and not x2 and x4 and x3 ) = '1' then
         y23 <= '1' ;
         y27 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1086;

      elsif ( x10 and not x18 and x19 and not x2 and x4 and not x3 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s428;

      elsif ( x10 and not x18 and x19 and not x2 and not x4 and x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s83;

      elsif ( x10 and not x18 and x19 and not x2 and not x4 and not x3 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1087;

      elsif ( x10 and not x18 and not x19 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1085;

      else
         y5 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         y30 <= '1' ;
         y35 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s895;

      end if;

   when s1023 =>
      if ( x63 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1087;

      elsif ( x63 and x19 and not x18 ) = '1' then
         y25 <= '1' ;
         y29 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s560;

      elsif ( x63 and not x19 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s806;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1159;

      end if;

   when s1024 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s808;

   when s1025 =>
      if ( x64 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1160;

      else
         y48 <= '1' ;
         y55 <= '1' ;
         y61 <= '1' ;
         current_otherm <= s1035;

      end if;

   when s1026 =>
      if ( x9 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1161;

      elsif ( not x9 and x15 and x11 and x6 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x9 and x15 and x11 and x6 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and x12 and x18 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and not x12 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x15 and x11 and not x6 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and x11 and not x6 and not x7 and not x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and not x11 and x6 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s963;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and not x12 and x10 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and not x13 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x15 and not x11 and not x6 and x7 and not x12 and not x10 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x9 and x15 and not x11 and not x6 and not x7 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y33 <= '1' ;
         y40 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1162;

      end if;

   when s1027 =>
      if ( x63 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1163;

      elsif ( x63 and x19 and not x18 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1164;

      elsif ( x63 and not x19 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s561;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1165;

      end if;

   when s1028 =>
      if ( x21 and x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( x21 and not x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( not x21 and x5 and x8 and x7 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( not x21 and x5 and x8 and not x7 and x9 and x18 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x21 and x5 and x8 and not x7 and x9 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x5 and x8 and not x7 and x9 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x5 and x8 and not x7 and not x9 and x19 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x21 and x5 and x8 and not x7 and not x9 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x5 and x8 and not x7 and not x9 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x5 and not x8 and x7 and x9 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s1027;

      elsif ( not x21 and x5 and not x8 and x7 and not x9 and x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x21 and x5 and not x8 and x7 and not x9 and not x20 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x5 and not x8 and x7 and not x9 and not x20 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x21 and x5 and not x8 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      else
         y44 <= '1' ;
         current_otherm <= s391;

      end if;

   when s1029 =>
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s1166;

   when s1030 =>
      if ( x5 and x21 and x7 and x9 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x5 and x21 and x7 and not x9 ) = '1' then
         y50 <= '1' ;
         current_otherm <= s282;

      elsif ( x5 and x21 and not x7 and x8 and x9 and x12 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x5 and x21 and not x7 and x8 and x9 and not x12 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x5 and x21 and not x7 and x8 and x9 and not x12 and x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and x21 and not x7 and x8 and x9 and not x12 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and x21 and not x7 and x8 and not x9 and x11 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x5 and x21 and not x7 and x8 and not x9 and not x11 and x10 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( x5 and x21 and not x7 and x8 and not x9 and not x11 and x10 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and x21 and not x7 and x8 and not x9 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x5 and x21 and not x7 and not x8 and x9 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s820;

      elsif ( x5 and x21 and not x7 and not x8 and not x9 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y16 <= '1' ;
         y42 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s820;

      elsif ( x5 and not x21 and x16 ) = '1' then
         y34 <= '1' ;
         current_otherm <= s178;

      elsif ( x5 and not x21 and not x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1028;

      elsif ( not x5 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1028;

      elsif ( not x5 and not x6 and x8 and x9 and x21 and x7 ) = '1' then
         y36 <= '1' ;
         current_otherm <= s260;

      elsif ( not x5 and not x6 and x8 and x9 and x21 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1167;

      elsif ( not x5 and not x6 and x8 and x9 and not x21 and x7 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and x8 and x9 and not x21 and not x7 ) = '1' then
         y6 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and x8 and not x9 and x21 and x7 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( not x5 and not x6 and x8 and not x9 and x21 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y31 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and x8 and not x9 and not x21 and x7 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and x8 and not x9 and not x21 and not x7 ) = '1' then
         y6 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and not x8 and x21 and x9 and x7 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x5 and not x6 and not x8 and x21 and x9 and not x7 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and not x8 and x21 and not x9 and x7 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and not x8 and x21 and not x9 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and not x8 and not x21 and x7 and x9 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x5 and not x6 and not x8 and not x21 and x7 and not x9 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      else
         y6 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      end if;

   when s1031 =>
      if ( x63 ) = '1' then
         y9 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1;

      else
         y11 <= '1' ;
         current_otherm <= s350;

      end if;

   when s1032 =>
         y11 <= '1' ;
         current_otherm <= s284;

   when s1033 =>
      if ( x26 and x27 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x26 and x27 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x26 and x27 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x26 and x27 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x26 and x27 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x26 and not x27 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1031;

      elsif ( not x26 and x7 and x8 and x6 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x7 and x8 and x6 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x7 and x8 and x6 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and x8 and x6 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and x8 and x6 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and x8 and not x6 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x7 and x8 and not x6 and not x9 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and x8 and not x6 and not x9 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and x8 and not x6 and not x9 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and not x8 and x6 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s350;

      elsif ( not x26 and x7 and not x8 and not x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and x7 and not x8 and not x6 and not x10 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and not x8 and not x6 and not x10 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and x7 and not x8 and not x6 and not x10 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and not x7 and x8 and x6 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1032;

      elsif ( not x26 and not x7 and x8 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x26 and not x7 and not x8 and x6 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( not x26 and not x7 and not x8 and x6 and not x11 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and not x7 and not x8 and x6 and not x11 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( not x26 and not x7 and not x8 and x6 and not x11 and not x22 ) = '1' then
         current_otherm <= s1;

      else
         y49 <= '1' ;
         current_otherm <= s256;

      end if;

   when s1034 =>
         y25 <= '1' ;
         current_otherm <= s1168;

   when s1035 =>
         y25 <= '1' ;
         current_otherm <= s23;

   when s1036 =>
         y10 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1;

   when s1037 =>
         y74 <= '1' ;
         current_otherm <= s1169;

   when s1038 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1016;

   when s1039 =>
      if ( x18 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1170;

      else
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1039;

      end if;

   when s1040 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1171;

   when s1041 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s1172;

   when s1042 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s962;

   when s1043 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s1173;

   when s1044 =>
      if ( x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1040;

      elsif ( not x4 and x5 and x6 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1041;

      elsif ( not x4 and x5 and x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1042;

      elsif ( not x4 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s958;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1043;

      end if;

   when s1045 =>
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s1174;

   when s1046 =>
      if ( x16 and x6 and x4 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x16 and x6 and not x4 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x16 and x6 and not x4 and not x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x16 and not x6 and x5 ) = '1' then
         y37 <= '1' ;
         current_otherm <= s181;

      elsif ( x16 and not x6 and not x5 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y65 <= '1' ;
         y66 <= '1' ;
         current_otherm <= s541;

      end if;

   when s1047 =>
         y17 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s837;

   when s1048 =>
         y11 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1;

   when s1049 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s1175;

   when s1050 =>
      if ( x62 and x33 and x32 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and x33 and not x32 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( x62 and not x33 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1176;

      end if;

   when s1051 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s429;

   when s1052 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1177;

   when s1053 =>
         y9 <= '1' ;
         current_otherm <= s162;

   when s1054 =>
         y25 <= '1' ;
         current_otherm <= s1178;

   when s1055 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s1179;

   when s1056 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_otherm <= s1180;

   when s1057 =>
      if ( x64 and x20 ) = '1' then
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s294;

      elsif ( x64 and not x20 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s594;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_otherm <= s129;

      end if;

   when s1058 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s1181;

   when s1059 =>
      if ( x14 and x7 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1060;

      elsif ( x14 and not x7 and x5 and x10 and x9 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1061;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and x11 and x16 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and x11 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and not x11 and x17 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x7 and x5 and x10 and not x9 and not x11 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x7 and x5 and not x10 and x11 and x9 ) = '1' then
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s84;

      elsif ( x14 and not x7 and x5 and not x10 and x11 and not x9 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( x14 and not x7 and x5 and not x10 and not x11 and x9 and x15 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x7 and x5 and not x10 and not x11 and x9 and not x15 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x7 and x5 and not x10 and not x11 and not x9 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      elsif ( x14 and not x7 and not x5 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1062;

      else
         y2 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1063;

      end if;

   when s1060 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1182;

   when s1061 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1183;

   when s1062 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1184;

   when s1063 =>
      if ( x7 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1060;

      elsif ( not x7 and x5 and x10 and x9 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1061;

      elsif ( not x7 and x5 and x10 and not x9 and x11 and x16 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x7 and x5 and x10 and not x9 and x11 and not x16 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x5 and x10 and not x9 and x11 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x5 and x10 and not x9 and not x11 and x17 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x7 and x5 and x10 and not x9 and not x11 and not x17 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x5 and x10 and not x9 and not x11 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x5 and not x10 and x11 and x9 ) = '1' then
         y6 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s84;

      elsif ( not x7 and x5 and not x10 and x11 and not x9 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x7 and x5 and not x10 and not x11 and x9 and x15 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x7 and x5 and not x10 and not x11 and x9 and not x15 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x5 and not x10 and not x11 and x9 and not x15 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x5 and not x10 and not x11 and not x9 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s117;

      else
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1062;

      end if;

   when s1064 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1185;

   when s1065 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y52 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s1186;

   when s1066 =>
      if ( x62 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x62 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x62 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x62 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x62 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y47 <= '1' ;
         y57 <= '1' ;
         y61 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s779;

      end if;

   when s1067 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s864;

   when s1068 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s864;

   when s1069 =>
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1187;

   when s1070 =>
         y7 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s294;

   when s1071 =>
         y14 <= '1' ;
         current_otherm <= s5;

   when s1072 =>
         y1 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s315;

   when s1073 =>
         y41 <= '1' ;
         current_otherm <= s376;

   when s1074 =>
      if ( x17 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s322;

      else
         y5 <= '1' ;
         y13 <= '1' ;
         y17 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1074;

      end if;

   when s1075 =>
         y25 <= '1' ;
         current_otherm <= s1066;

   when s1076 =>
         y11 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s1188;

   when s1077 =>
      if ( x20 and x21 ) = '1' then
         y6 <= '1' ;
         y17 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s93;

      elsif ( x20 and not x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1189;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1190;

      end if;

   when s1078 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1191;

   when s1079 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1192;

   when s1080 =>
         y1 <= '1' ;
         y3 <= '1' ;
         y8 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1193;

   when s1081 =>
      if ( x11 and x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s889;

      elsif ( x11 and not x10 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s727;

      else
         y29 <= '1' ;
         current_otherm <= s887;

      end if;

   when s1082 =>
      if ( x21 and x20 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s63;

      elsif ( x21 and not x20 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s886;

      else
         y22 <= '1' ;
         current_otherm <= s63;

      end if;

   when s1083 =>
      if ( x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( not x5 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x5 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x5 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1084 =>
      if ( x63 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      else
         y10 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1;

      end if;

   when s1085 =>
      if ( x19 and x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s1023;

      elsif ( x19 and not x18 ) = '1' then
         y23 <= '1' ;
         y27 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1194;

      else
         y2 <= '1' ;
         current_otherm <= s1027;

      end if;

   when s1086 =>
         y2 <= '1' ;
         current_otherm <= s1195;

   when s1087 =>
         y2 <= '1' ;
         current_otherm <= s1027;

   when s1088 =>
         y12 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s560;

   when s1089 =>
         y10 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1;

   when s1090 =>
         y25 <= '1' ;
         current_otherm <= s679;

   when s1091 =>
      if ( x23 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s905;

      elsif ( x23 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s906;

      elsif ( not x23 and x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s905;

      elsif ( not x23 and x22 and not x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s906;

      elsif ( not x23 and not x22 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s906;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s905;

      end if;

   when s1092 =>
         y55 <= '1' ;
         current_otherm <= s388;

   when s1093 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1196;

   when s1094 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1197;

   when s1095 =>
      if ( x66 and x7 and x11 and x13 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s88;

      elsif ( x66 and x7 and x11 and x13 and x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s846;

      elsif ( x66 and x7 and x11 and x13 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s847;

      elsif ( x66 and x7 and x11 and x13 and not x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s848;

      elsif ( x66 and x7 and x11 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and x11 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and x11 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and x11 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and x15 and x13 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( x66 and x7 and not x11 and x12 and x15 and x13 and not x14 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( x66 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and x15 and not x13 and x14 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s460;

      elsif ( x66 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and x15 and not x13 and not x14 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and x13 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and x13 and not x14 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and not x13 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s849;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( x66 and x7 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s850;

      elsif ( x66 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1198;

      elsif ( not x66 and x26 and x25 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and x26 and not x25 and x24 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( not x66 and x26 and not x25 and not x24 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1096 =>
      if ( x65 ) = '1' then
         y42 <= '1' ;
         current_otherm <= s1034;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s1199;

      end if;

   when s1097 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

   when s1098 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s795;

   when s1099 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s537;

   when s1100 =>
      if ( x23 and x4 and x5 and x3 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and x4 and x5 and x3 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and x4 and x5 and x3 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and x4 and x5 and x3 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and x4 and x5 and not x3 and x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x23 and x4 and x5 and not x3 and not x12 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and x4 and x5 and not x3 and not x12 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and x4 and x5 and not x3 and not x12 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and x4 and x5 and not x3 and not x12 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and x4 and not x5 and x3 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s856;

      elsif ( x23 and x4 and not x5 and not x3 and x11 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x23 and x4 and not x5 and not x3 and not x11 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and x4 and not x5 and not x3 and not x11 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and x4 and not x5 and not x3 and not x11 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and x4 and not x5 and not x3 and not x11 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and not x4 and x3 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s621;

      elsif ( x23 and not x4 and x3 and not x5 and x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x23 and not x4 and x3 and not x5 and not x13 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and not x4 and x3 and not x5 and not x13 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x23 and not x4 and x3 and not x5 and not x13 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and not x4 and x3 and not x5 and not x13 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x23 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( not x23 and x22 and x4 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1099;

      elsif ( not x23 and x22 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( not x23 and x22 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s337;

      else
         y6 <= '1' ;
         current_otherm <= s856;

      end if;

   when s1101 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y27 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s1200;

   when s1102 =>
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s395;

   when s1103 =>
      if ( x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1104 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1201;

   when s1105 =>
      if ( x2 and x3 and x4 and x9 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x2 and x3 and x4 and x9 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x2 and x3 and x4 and x9 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x2 and x3 and x4 and x9 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x2 and x3 and x4 and not x9 and x8 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( x2 and x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x2 and x3 and not x4 and x9 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s681;

      elsif ( x2 and x3 and not x4 and x9 and not x6 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( x2 and x3 and not x4 and not x9 and x8 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x2 and x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x2 and not x3 and x4 and x9 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s894;

      elsif ( x2 and not x3 and x4 and not x9 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( x2 and not x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x2 and not x3 and not x4 and x9 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x2 and not x3 and not x4 and x9 and not x13 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( x2 and not x3 and not x4 and x9 and not x13 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( x2 and not x3 and not x4 and not x9 and x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( x2 and not x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x2 and x4 and x3 and x9 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x2 and x4 and x3 and x9 and not x14 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x2 and x4 and x3 and x9 and not x14 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x2 and x4 and x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1104;

      elsif ( not x2 and x4 and x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x2 and x4 and not x3 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x2 and x4 and not x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x2 and x4 and not x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x2 and not x4 and x9 and x3 and x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x2 and not x4 and x9 and x3 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x2 and not x4 and x9 and x3 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x2 and not x4 and x9 and not x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( not x2 and not x4 and not x9 and x8 and x3 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x2 and not x4 and not x9 and x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      end if;

   when s1106 =>
      if ( x7 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1202;

      elsif ( not x7 and x9 and x6 and x12 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s790;

      elsif ( not x7 and x9 and x6 and not x12 and x11 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s410;

      elsif ( not x7 and x9 and x6 and not x12 and not x11 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and x6 and not x12 and not x11 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and x6 and not x12 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and x6 and not x12 and not x11 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and x10 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and not x10 and x16 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and not x12 and x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s791;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and not x12 and not x10 and x17 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s792;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and not x12 and x10 and x15 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x7 and x9 and not x6 and x8 and not x11 and not x12 and not x10 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x7 and x9 and not x6 and not x8 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s790;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y28 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s477;

      end if;

   when s1107 =>
      if ( x19 and x20 and x2 and x1 and x4 and x3 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x19 and x20 and x2 and x1 and x4 and x3 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x19 and x20 and x2 and x1 and x4 and x3 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x20 and x2 and x1 and x4 and x3 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and x5 and x18 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and x22 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and x5 and not x18 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and x21 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and x22 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x20 and x2 and x1 and x4 and not x3 and not x5 and not x21 and not x22 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x20 and x2 and x1 and not x4 and x5 and x3 ) = '1' then
         y23 <= '1' ;
         current_otherm <= s169;

      elsif ( x19 and x20 and x2 and x1 and not x4 and x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s342;

      elsif ( x19 and x20 and x2 and x1 and not x4 and not x5 and x3 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( x19 and x20 and x2 and x1 and not x4 and not x5 and not x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y34 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s342;

      elsif ( x19 and x20 and x2 and not x1 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( x19 and x20 and not x2 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         current_otherm <= s696;

      elsif ( x19 and x20 and not x2 and not x8 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( x19 and not x20 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s697;

      elsif ( not x19 and x11 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s698;

      else
         y29 <= '1' ;
         current_otherm <= s378;

      end if;

   when s1108 =>
      if ( x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1190;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1203;

      end if;

   when s1109 =>
         y42 <= '1' ;
         current_otherm <= s1054;

   when s1110 =>
         y42 <= '1' ;
         current_otherm <= s1165;

   when s1111 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1204;

   when s1112 =>
      if ( x15 ) = '1' then
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1205;

      else
         y6 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s1206;

      end if;

   when s1113 =>
         y3 <= '1' ;
         current_otherm <= s949;

   when s1114 =>
         y4 <= '1' ;
         y31 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s1207;

   when s1115 =>
         y4 <= '1' ;
         y31 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s1208;

   when s1116 =>
      if ( x8 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x8 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x8 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x9 and x11 and x10 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x8 and not x9 and x11 and x10 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x8 and not x9 and x11 and x10 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x9 and x11 and x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x9 and x11 and not x10 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s504;

      elsif ( x8 and not x9 and not x11 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1114;

      elsif ( x8 and not x9 and not x11 and not x10 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x8 and not x9 and not x11 and not x10 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x8 and not x9 and not x11 and not x10 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x9 and not x11 and not x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and x10 and x11 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and x10 and x11 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and x10 and x11 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and x10 and x11 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and x10 and x11 and not x9 and x18 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and x10 and x11 and not x9 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and x10 and not x11 and x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( not x8 and x6 and x10 and not x11 and not x9 and x17 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and x10 and not x11 and not x9 and not x17 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and not x10 and x11 and x9 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1115;

      elsif ( not x8 and x6 and not x10 and x11 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( not x8 and x6 and not x10 and not x11 and x9 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and not x10 and not x11 and x9 and not x19 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( not x8 and x6 and not x10 and not x11 and not x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      else
         y2 <= '1' ;
         current_otherm <= s1023;

      end if;

   when s1117 =>
      if ( x63 ) = '1' then
         y23 <= '1' ;
         y29 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s560;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1209;

      end if;

   when s1118 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1210;

   when s1119 =>
         y3 <= '1' ;
         current_otherm <= s208;

   when s1120 =>
         y28 <= '1' ;
         current_otherm <= s296;

   when s1121 =>
      if ( x20 and x22 and x23 and x24 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x20 and x22 and x23 and not x24 and x25 ) = '1' then
         y59 <= '1' ;
         current_otherm <= s186;

      elsif ( x20 and x22 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( x20 and x22 and not x23 ) = '1' then
         current_otherm <= s1;

      elsif ( x20 and not x22 ) = '1' then
         current_otherm <= s1;

      else
         y11 <= '1' ;
         current_otherm <= s425;

      end if;

   when s1122 =>
      if ( x64 and x19 ) = '1' then
         y7 <= '1' ;
         current_otherm <= s739;

      elsif ( x64 and not x19 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x19 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x64 and not x19 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x64 and not x19 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y40 <= '1' ;
         current_otherm <= s478;

      end if;

   when s1123 =>
      if ( x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s1211;

      elsif ( not x6 and x10 and x2 and x3 and x4 and x9 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and x2 and x3 and x4 and x9 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and x2 and x3 and x4 and x9 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x2 and x3 and x4 and x9 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x2 and x3 and x4 and not x9 and x8 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( not x6 and x10 and x2 and x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and x2 and x3 and not x4 and x9 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x6 and x10 and x2 and x3 and not x4 and not x9 and x8 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( not x6 and x10 and x2 and x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and x2 and not x3 and x4 and x9 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s894;

      elsif ( not x6 and x10 and x2 and not x3 and x4 and not x9 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x6 and x10 and x2 and not x3 and x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and x9 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and x9 and not x13 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and x9 and not x13 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and not x9 and x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and x2 and not x3 and not x4 and not x9 and not x8 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and x9 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and x9 and not x14 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and x9 and not x14 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1104;

      elsif ( not x6 and x10 and not x2 and x4 and x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and not x2 and x4 and not x3 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x6 and x10 and not x2 and x4 and not x3 and not x9 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and not x2 and x4 and not x3 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and not x2 and not x4 and x9 and x3 and x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x6 and x10 and not x2 and not x4 and x9 and x3 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x6 and x10 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and not x2 and not x4 and x9 and x3 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x6 and x10 and not x2 and not x4 and x9 and not x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      elsif ( not x6 and x10 and not x2 and not x4 and not x9 and x8 and x3 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and not x2 and not x4 and not x9 and x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x6 and x10 and not x2 and not x4 and not x9 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y36 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1105;

      end if;

   when s1124 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1212;

   when s1125 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s1213;

   when s1126 =>
      if ( x12 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x12 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x12 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x12 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1127 =>
         y5 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1214;

   when s1128 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1215;

   when s1129 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y55 <= '1' ;
         y63 <= '1' ;
         current_otherm <= s742;

   when s1130 =>
         y3 <= '1' ;
         y26 <= '1' ;
         y55 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s742;

   when s1131 =>
      if ( x63 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s714;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y31 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s742;

      end if;

   when s1132 =>
      if ( x12 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s854;

      elsif ( not x12 and x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x12 and x15 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x12 and x15 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1133 =>
         y5 <= '1' ;
         y12 <= '1' ;
         y19 <= '1' ;
         y25 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s742;

   when s1134 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y54 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s742;

   when s1135 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y53 <= '1' ;
         y55 <= '1' ;
         current_otherm <= s742;

   when s1136 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y28 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s756;

   when s1137 =>
      if ( x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s970;

      elsif ( not x5 and x7 and x11 and x13 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s88;

      elsif ( not x5 and x7 and x11 and x13 and x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s846;

      elsif ( not x5 and x7 and x11 and x13 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s847;

      elsif ( not x5 and x7 and x11 and x13 and not x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s848;

      elsif ( not x5 and x7 and x11 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and x11 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and x11 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and x11 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and x13 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and x13 and not x14 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and x13 and not x14 and not x16 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and not x13 and x14 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s460;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and not x13 and x14 and not x18 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and x15 and not x13 and not x14 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and x13 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and x13 and not x14 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and x13 and not x14 and not x17 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and not x13 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s849;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and x12 and not x15 and not x13 and not x14 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x7 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s850;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1198;

      end if;

   when s1138 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y42 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1216;

   when s1139 =>
      if ( x14 and x13 ) = '1' then
         y5 <= '1' ;
         y29 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y53 <= '1' ;
         current_otherm <= s460;

      elsif ( x14 and not x13 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1217;

      elsif ( x14 and not x13 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s1218;

      elsif ( not x14 and x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s460;

      elsif ( not x14 and x15 and not x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s1219;

      elsif ( not x14 and not x15 and x13 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y53 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s460;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s1220;

      end if;

   when s1140 =>
      if ( x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s856;

      elsif ( not x4 and x12 and x11 and x14 and x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s460;

      elsif ( not x4 and x12 and x11 and x14 and x15 and not x13 ) = '1' then
         y35 <= '1' ;
         current_otherm <= s269;

      elsif ( not x4 and x12 and x11 and x14 and not x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s460;

      elsif ( not x4 and x12 and x11 and x14 and not x15 and not x13 ) = '1' then
         y18 <= '1' ;
         current_otherm <= s89;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and x15 and x9 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s425;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and x15 and not x9 and x8 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and x15 and not x9 and x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and x15 and not x9 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and not x15 and x10 ) = '1' then
         y11 <= '1' ;
         current_otherm <= s425;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and not x15 and not x10 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and not x15 and not x10 and x8 and not x9 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x12 and x11 and not x14 and x13 and not x15 and not x10 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x12 and x11 and not x14 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x4 and x12 and x11 and not x14 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x4 and x12 and x11 and not x14 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x12 and x11 and not x14 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x4 and x12 and not x11 and x13 and x14 and x15 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x4 and x12 and not x11 and x13 and x14 and not x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s586;

      elsif ( not x4 and x12 and not x11 and x13 and not x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s586;

      elsif ( not x4 and x12 and not x11 and not x13 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s586;

      elsif ( not x4 and not x12 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s586;

      elsif ( not x4 and not x12 and not x5 and x11 and x14 and x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s460;

      elsif ( not x4 and not x12 and not x5 and x11 and x14 and x15 and not x13 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s460;

      elsif ( not x4 and not x12 and not x5 and x11 and x14 and not x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s833;

      elsif ( not x4 and not x12 and not x5 and x11 and x14 and not x15 and not x13 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x4 and not x12 and not x5 and x11 and not x14 and x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s460;

      elsif ( not x4 and not x12 and not x5 and x11 and not x14 and x15 and not x13 ) = '1' then
         y40 <= '1' ;
         current_otherm <= s478;

      elsif ( not x4 and not x12 and not x5 and x11 and not x14 and not x15 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1221;

      elsif ( not x4 and not x12 and not x5 and x11 and not x14 and not x15 and not x13 ) = '1' then
         y39 <= '1' ;
         current_otherm <= s103;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1139;

      end if;

   when s1141 =>
         y2 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1222;

   when s1142 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s668;

   when s1143 =>
      if ( x5 ) = '1' then
         y1 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s1223;

      elsif ( not x5 and x32 and x13 and x15 and x33 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s854;

      elsif ( not x5 and x32 and x13 and x15 and not x33 and x14 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( not x5 and x32 and x13 and x15 and not x33 and not x14 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s140;

      elsif ( not x5 and x32 and x13 and x15 and not x33 and not x14 and not x16 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s141;

      elsif ( not x5 and x32 and x13 and not x15 and x33 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s593;

      elsif ( not x5 and x32 and x13 and not x15 and not x33 and x14 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s142;

      elsif ( not x5 and x32 and x13 and not x15 and not x33 and not x14 and x7 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s144;

      elsif ( not x5 and x32 and x13 and not x15 and not x33 and not x14 and not x7 ) = '1' then
         y8 <= '1' ;
         y36 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s442;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and x15 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s951;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and x15 and not x12 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and x15 and not x12 and x10 and not x11 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and x15 and not x12 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and not x15 and x11 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s952;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and not x15 and not x11 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s286;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and not x15 and not x11 and x10 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x32 and not x13 and x14 and x33 and not x15 and not x11 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x32 and not x13 and x14 and not x33 and x15 and x7 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s721;

      elsif ( not x5 and x32 and not x13 and x14 and not x33 and x15 and not x7 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s449;

      elsif ( not x5 and x32 and not x13 and x14 and not x33 and not x15 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s133;

      elsif ( not x5 and x32 and not x13 and x14 and not x33 and not x15 and not x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s439;

      elsif ( not x5 and x32 and not x13 and not x14 and x15 and x33 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x5 and x32 and not x13 and not x14 and x15 and not x33 and x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x32 and not x13 and not x14 and x15 and not x33 and not x17 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1224;

      elsif ( not x5 and x32 and not x13 and not x14 and x15 and not x33 and not x17 and not x7 ) = '1' then
         y30 <= '1' ;
         current_otherm <= s803;

      elsif ( not x5 and x32 and not x13 and not x14 and not x15 and x33 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s443;

      elsif ( not x5 and x32 and not x13 and not x14 and not x15 and not x33 and x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x32 and not x13 and not x14 and not x15 and not x33 and not x18 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s766;

      elsif ( not x5 and x32 and not x13 and not x14 and not x15 and not x33 and not x18 and not x7 ) = '1' then
         y6 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1225;

      elsif ( not x5 and not x32 and x13 and x14 and x33 and x15 and x7 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      elsif ( not x5 and not x32 and x13 and x14 and x33 and x15 and not x7 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s132;

      elsif ( not x5 and not x32 and x13 and x14 and x33 and not x15 ) = '1' then
         y53 <= '1' ;
         current_otherm <= s137;

      elsif ( not x5 and not x32 and x13 and x14 and not x33 and x7 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s132;

      elsif ( not x5 and not x32 and x13 and x14 and not x33 and not x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s143;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and x33 and x31 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and x33 and not x31 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and x33 and not x31 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and x33 and not x31 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and x33 and not x31 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and not x33 and x7 ) = '1' then
         y8 <= '1' ;
         y36 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s442;

      elsif ( not x5 and not x32 and x13 and not x14 and x15 and not x33 and not x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s136;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and x33 and x16 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and x33 and not x16 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and x33 and not x16 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and x33 and not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and x33 and not x16 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and not x33 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s400;

      elsif ( not x5 and not x32 and x13 and not x14 and not x15 and not x33 and not x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s943;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and x15 and x8 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and x15 and not x8 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and x15 and not x8 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and not x15 and x30 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and x11 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and not x11 and x12 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and not x13 and x33 and x14 and not x15 and not x30 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x32 and not x13 and x33 and not x14 and x15 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s134;

      elsif ( not x5 and not x32 and not x13 and x33 and not x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s138;

      elsif ( not x5 and not x32 and not x13 and not x33 and x7 ) = '1' then
         y6 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s131;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s140;

      end if;

   when s1144 =>
      if ( x65 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1226;

      else
         y6 <= '1' ;
         y41 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s395;

      end if;

   when s1145 =>
         y3 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1227;

   when s1146 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y57 <= '1' ;
         current_otherm <= s1228;

   when s1147 =>
      if ( x15 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s275;

      else
         y58 <= '1' ;
         current_otherm <= s774;

      end if;

   when s1148 =>
      if ( x8 and x20 and x14 and x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s668;

      elsif ( x8 and x20 and x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y42 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s855;

      elsif ( x8 and x20 and not x14 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1149;

      elsif ( x8 and not x20 and x13 and x21 and x14 and x15 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( x8 and not x20 and x13 and x21 and x14 and not x15 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( x8 and not x20 and x13 and x21 and x14 and not x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and x15 and x17 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and x15 and x17 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and x15 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and not x15 and x9 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and not x15 and x9 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and x13 and x21 and not x14 and not x15 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and x13 and not x21 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and x15 and x18 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and x15 and x18 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and x15 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and not x15 and x19 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and not x15 and x19 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and not x13 and x14 and x21 and not x15 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and not x13 and x14 and not x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( x8 and not x20 and not x13 and not x14 and x21 and x15 and x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( x8 and not x20 and not x13 and not x14 and x21 and x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s882;

      elsif ( x8 and not x20 and not x13 and not x14 and x21 and not x15 and x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s883;

      elsif ( x8 and not x20 and not x13 and not x14 and x21 and not x15 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s884;

      elsif ( x8 and not x20 and not x13 and not x14 and not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and not x13 and not x14 and not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x8 and not x20 and not x13 and not x14 and not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x8 and not x20 and not x13 and not x14 and not x21 and not x10 ) = '1' then
         current_otherm <= s1;

      else
         y6 <= '1' ;
         y9 <= '1' ;
         y25 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1150;

      end if;

   when s1149 =>
         y11 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s1229;

   when s1150 =>
      if ( x9 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s611;

      elsif ( not x9 and x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1203;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y15 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1189;

      end if;

   when s1151 =>
      if ( x19 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1006;

      elsif ( not x19 and x11 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s1007;

      else
         y29 <= '1' ;
         current_otherm <= s470;

      end if;

   when s1152 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1230;

   when s1153 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1231;

   when s1154 =>
         y24 <= '1' ;
         current_otherm <= s322;

   when s1155 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s342;

   when s1156 =>
         y10 <= '1' ;
         current_otherm <= s651;

   when s1157 =>
         y8 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s138;

   when s1158 =>
      if ( x19 and x18 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s504;

      elsif ( x19 and not x18 ) = '1' then
         y23 <= '1' ;
         y28 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1232;

      else
         y2 <= '1' ;
         current_otherm <= s1023;

      end if;

   when s1159 =>
      if ( x3 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and not x9 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         y26 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and not x9 and x10 and not x11 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         y26 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s769;

      elsif ( x3 and not x9 and not x10 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s769;

      else
         y14 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1233;

      end if;

   when s1160 =>
      if ( x12 and x11 and x6 ) = '1' then
         y5 <= '1' ;
         y27 <= '1' ;
         y49 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s407;

      elsif ( x12 and x11 and not x6 and x10 ) = '1' then
         y47 <= '1' ;
         current_otherm <= s278;

      elsif ( x12 and x11 and not x6 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( x12 and not x11 and x6 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( x12 and not x11 and not x6 and x10 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s409;

      elsif ( x12 and not x11 and not x6 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x12 and x11 and x6 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s410;

      elsif ( not x12 and x11 and not x6 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( not x12 and x11 and not x6 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_otherm <= s408;

      elsif ( not x12 and not x11 and x6 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x12 and not x11 and x6 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x12 and not x11 and x6 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and not x11 and x6 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( not x12 and not x11 and not x6 and x10 ) = '1' then
         y54 <= '1' ;
         current_otherm <= s253;

      elsif ( not x12 and not x11 and not x6 and not x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x12 and not x11 and not x6 and not x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( not x12 and not x11 and not x6 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1161 =>
         y44 <= '1' ;
         current_otherm <= s391;

   when s1162 =>
      if ( x11 and x6 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x11 and x6 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x11 and not x6 and x7 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( x11 and not x6 and x7 and not x10 and x12 and x18 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x11 and not x6 and x7 and not x10 and x12 and not x18 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and not x6 and x7 and not x10 and not x12 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x11 and not x6 and x7 and not x10 and not x12 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and not x6 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( x11 and not x6 and not x7 and not x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( not x11 and x6 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x11 and not x6 and x7 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s963;

      elsif ( not x11 and not x6 and x7 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( not x11 and not x6 and x7 and not x12 and x10 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and not x13 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( not x11 and not x6 and x7 and not x12 and x10 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and not x6 and x7 and not x12 and not x10 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      else
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      end if;

   when s1163 =>
         y9 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         y32 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s936;

   when s1164 =>
         y2 <= '1' ;
         current_otherm <= s392;

   when s1165 =>
         y25 <= '1' ;
         current_otherm <= s1234;

   when s1166 =>
      if ( x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

      elsif ( not x21 and x8 and x9 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s820;

      elsif ( not x21 and x8 and not x9 ) = '1' then
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s820;

      else
         y6 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s820;

      end if;

   when s1167 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y31 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1235;

   when s1168 =>
      if ( x64 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s182;

      elsif ( not x64 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y47 <= '1' ;
         y53 <= '1' ;
         y61 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s913;

      end if;

   when s1169 =>
      if ( x15 ) = '1' then
         y46 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s240;

      elsif ( not x15 and x6 and x7 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and x8 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s111;

      elsif ( not x15 and x6 and not x7 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1170 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1236;

   when s1171 =>
      if ( x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1171;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1237;

      end if;

   when s1172 =>
      if ( x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_otherm <= s1202;

      else
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_otherm <= s1172;

      end if;

   when s1173 =>
      if ( x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1238;

      else
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s1173;

      end if;

   when s1174 =>
      if ( x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s497;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_otherm <= s1045;

      end if;

   when s1175 =>
      if ( x14 and x6 and x8 and x7 ) = '1' then
         y63 <= '1' ;
         current_otherm <= s224;

      elsif ( x14 and x6 and x8 and not x7 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x14 and x6 and x8 and not x7 and x9 and not x18 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x14 and x6 and x8 and not x7 and x9 and not x18 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x14 and x6 and x8 and not x7 and x9 and not x18 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and x8 and not x7 and x9 and not x18 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and x8 and not x7 and not x9 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x14 and x6 and x8 and not x7 and not x9 and not x19 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x14 and x6 and x8 and not x7 and not x9 and not x19 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x14 and x6 and x8 and not x7 and not x9 and not x19 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and x8 and not x7 and not x9 and not x19 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and not x8 and x9 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_otherm <= s575;

      elsif ( x14 and x6 and not x8 and x9 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x14 and x6 and not x8 and not x9 and x7 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_otherm <= s275;

      elsif ( x14 and x6 and not x8 and not x9 and x7 and not x17 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x14 and x6 and not x8 and not x9 and x7 and not x17 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s171;

      elsif ( x14 and x6 and not x8 and not x9 and x7 and not x17 and x20 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and not x8 and not x9 and x7 and not x17 and not x20 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and not x8 and not x9 and not x7 ) = '1' then
         y65 <= '1' ;
         current_otherm <= s155;

      elsif ( x14 and not x6 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s576;

      end if;

   when s1176 =>
         y9 <= '1' ;
         current_otherm <= s285;

   when s1177 =>
         y9 <= '1' ;
         current_otherm <= s1239;

   when s1178 =>
      if ( x64 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s877;

      elsif ( not x64 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y47 <= '1' ;
         y55 <= '1' ;
         y61 <= '1' ;
         y71 <= '1' ;
         current_otherm <= s930;

      end if;

   when s1179 =>
         y23 <= '1' ;
         y72 <= '1' ;
         y73 <= '1' ;
         current_otherm <= s1;

   when s1180 =>
         y13 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1;

   when s1181 =>
         y53 <= '1' ;
         current_otherm <= s455;

   when s1182 =>
         y1 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1240;

   when s1183 =>
         y1 <= '1' ;
         y4 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s1241;

   when s1184 =>
         y1 <= '1' ;
         y4 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1242;

   when s1185 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s864;

   when s1186 =>
         y9 <= '1' ;
         y18 <= '1' ;
         y48 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s864;

   when s1187 =>
         y5 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s864;

   when s1188 =>
      if ( x16 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s395;

      elsif ( not x16 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x16 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1189 =>
      if ( x20 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1243;

      else
         y6 <= '1' ;
         y9 <= '1' ;
         y25 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1108;

      end if;

   when s1190 =>
      if ( x20 and x14 and x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s668;

      elsif ( x20 and x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y42 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s855;

      elsif ( x20 and not x14 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1149;

      elsif ( not x20 and x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1244;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1243;

      end if;

   when s1191 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1071;

   when s1192 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s1243;

   when s1193 =>
      if ( x19 and x23 and x4 and x5 and x3 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and x4 and x5 and x3 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and x4 and x5 and x3 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and x4 and x5 and x3 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and x4 and x5 and not x3 and x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x19 and x23 and x4 and x5 and not x3 and not x12 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and x4 and x5 and not x3 and not x12 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and x4 and x5 and not x3 and not x12 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and x4 and x5 and not x3 and not x12 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and x4 and not x5 and x3 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s856;

      elsif ( x19 and x23 and x4 and not x5 and not x3 and x11 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x19 and x23 and x4 and not x5 and not x3 and not x11 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and x4 and not x5 and not x3 and not x11 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and x4 and not x5 and not x3 and not x11 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and x4 and not x5 and not x3 and not x11 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and not x4 and x3 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y19 <= '1' ;
         current_otherm <= s621;

      elsif ( x19 and x23 and not x4 and x3 and not x5 and x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x19 and x23 and not x4 and x3 and not x5 and not x13 and x21 and x16 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and not x4 and x3 and not x5 and not x13 and x21 and not x16 and x15 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( x19 and x23 and not x4 and x3 and not x5 and not x13 and x21 and not x16 and not x15 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and not x4 and x3 and not x5 and not x13 and not x21 ) = '1' then
         current_otherm <= s1;

      elsif ( x19 and x23 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_otherm <= s302;

      elsif ( x19 and not x23 and x22 and x4 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1099;

      elsif ( x19 and not x23 and x22 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s39;

      elsif ( x19 and not x23 and x22 and not x4 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s337;

      elsif ( x19 and not x23 and not x22 ) = '1' then
         y6 <= '1' ;
         current_otherm <= s856;

      else
         y1 <= '1' ;
         y8 <= '1' ;
         y23 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s1100;

      end if;

   when s1194 =>
         y2 <= '1' ;
         current_otherm <= s1245;

   when s1195 =>
         y23 <= '1' ;
         y28 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s1246;

   when s1196 =>
         y7 <= '1' ;
         y39 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1247;

   when s1197 =>
         y3 <= '1' ;
         y13 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s756;

   when s1198 =>
      if ( x11 and x13 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s88;

      elsif ( x11 and x13 and x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y58 <= '1' ;
         current_otherm <= s846;

      elsif ( x11 and x13 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y59 <= '1' ;
         current_otherm <= s847;

      elsif ( x11 and x13 and not x15 and not x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s848;

      elsif ( x11 and not x13 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x11 and not x13 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( x11 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and not x13 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and x15 and x13 and x14 ) = '1' then
         y61 <= '1' ;
         current_otherm <= s498;

      elsif ( not x11 and x12 and x15 and x13 and not x14 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and x15 and x13 and not x14 and not x16 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and x15 and x13 and not x14 and not x16 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and x15 and not x13 and x14 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s460;

      elsif ( not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and x15 and not x13 and x14 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and x15 and not x13 and x14 and not x18 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and x15 and not x13 and not x14 ) = '1' then
         y9 <= '1' ;
         current_otherm <= s43;

      elsif ( not x11 and x12 and not x15 and x13 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x11 and x12 and not x15 and x13 and not x14 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_otherm <= s718;

      elsif ( not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and not x15 and x13 and not x14 and not x17 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and not x15 and x13 and not x14 and not x17 and not x8 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and not x15 and not x13 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y62 <= '1' ;
         current_otherm <= s849;

      elsif ( not x11 and x12 and not x15 and not x13 and not x14 and x8 and x9 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and x10 ) = '1' then
         y64 <= '1' ;
         current_otherm <= s226;

      elsif ( not x11 and x12 and not x15 and not x13 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x11 and x12 and not x15 and not x13 and not x14 and not x8 ) = '1' then
         current_otherm <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s850;

      end if;

   when s1199 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y26 <= '1' ;
         current_otherm <= s1248;

   when s1200 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s302;

   when s1201 =>
         y3 <= '1' ;
         y18 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s1103;

   when s1202 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1249;

   when s1203 =>
      if ( x20 ) = '1' then
         y6 <= '1' ;
         y9 <= '1' ;
         y25 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1108;

      elsif ( not x20 and x13 and x21 and x14 and x15 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s225;

      elsif ( not x20 and x13 and x21 and x14 and not x15 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x13 and x21 and x14 and not x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x13 and x21 and not x14 and x15 and x17 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x13 and x21 and not x14 and x15 and x17 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x13 and x21 and not x14 and x15 and not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x13 and x21 and not x14 and x15 and not x17 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x13 and x21 and not x14 and not x15 and x9 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and x13 and x21 and not x14 and not x15 and x9 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and x13 and x21 and not x14 and not x15 and not x9 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x13 and x21 and not x14 and not x15 and not x9 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and x13 and not x21 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

      elsif ( not x20 and not x13 and x14 and x21 and x15 and x18 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and not x13 and x14 and x21 and x15 and x18 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x13 and x14 and x21 and x15 and not x18 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x13 and x14 and x21 and x15 and not x18 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x13 and x14 and x21 and not x15 and x19 and x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s426;

      elsif ( not x20 and not x13 and x14 and x21 and not x15 and x19 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s881;

      elsif ( not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x13 and x14 and x21 and not x15 and not x19 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x13 and x14 and x21 and not x15 and not x19 and not x10 ) = '1' then
         current_otherm <= s1;

      elsif ( not x20 and not x13 and x14 and not x21 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x20 and not x13 and not x14 and x21 and x15 and x5 ) = '1' then
         y14 <= '1' ;
         current_otherm <= s5;

      elsif ( not x20 and not x13 and not x14 and x21 and x15 and not x5 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s882;

      elsif ( not x20 and not x13 and not x14 and x21 and not x15 and x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s883;

      elsif ( not x20 and not x13 and not x14 and x21 and not x15 and not x7 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s884;

      elsif ( not x20 and not x13 and not x14 and not x21 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x13 and not x14 and not x21 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x13 and not x14 and not x21 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1204 =>
      if ( x15 and x11 and x6 and x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x15 and x11 and x6 and not x12 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and x11 and not x6 and x7 and x10 ) = '1' then
         y48 <= '1' ;
         current_otherm <= s411;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and x12 and x18 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y21 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s404;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and x12 and not x18 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and not x12 and x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and x19 and not x14 and not x13 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and x11 and not x6 and x7 and not x10 and not x12 and not x17 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x15 and x11 and not x6 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and x11 and not x6 and not x7 and not x12 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and not x11 and x6 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and not x11 and not x6 and x7 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s963;

      elsif ( x15 and not x11 and not x6 and x7 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and not x11 and not x6 and x7 and not x12 and x10 and x16 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and x14 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_otherm <= s203;

      elsif ( x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and x19 and not x14 and not x13 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s405;

      elsif ( x15 and not x11 and not x6 and x7 and not x12 and x10 and not x16 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x15 and not x11 and not x6 and x7 and not x12 and not x10 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( x15 and not x11 and not x6 and not x7 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y34 <= '1' ;
         y38 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s405;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y33 <= '1' ;
         y40 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s1162;

      end if;

   when s1205 =>
      if ( x17 ) = '1' then
         y43 <= '1' ;
         current_otherm <= s175;

      elsif ( not x17 and x10 and x11 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x17 and x10 and not x11 and x12 ) = '1' then
         y41 <= '1' ;
         current_otherm <= s376;

      elsif ( not x17 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1206 =>
         y44 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s933;

   when s1207 =>
      if ( x3 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x3 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x3 and not x14 ) = '1' then
         current_otherm <= s1;

      else
         y14 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1114;

      end if;

   when s1208 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s769;

      else
         y14 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1115;

      end if;

   when s1209 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y7 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s1250;

      else
         y14 <= '1' ;
         y37 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s1251;

      end if;

   when s1210 =>
         y2 <= '1' ;
         y15 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s1252;

   when s1211 =>
         y35 <= '1' ;
         current_otherm <= s383;

   when s1212 =>
      if ( x5 ) = '1' then
         y15 <= '1' ;
         current_otherm <= s1057;

      elsif ( not x5 and x8 and x9 and x3 and x2 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and x8 and x9 and x3 and x2 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and x8 and x9 and x3 and x2 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x8 and x9 and x3 and x2 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and x4 and x17 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and x4 and not x17 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and x4 and not x17 and x1 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and x4 and not x17 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and not x4 and x16 ) = '1' then
         y17 <= '1' ;
         current_otherm <= s179;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and not x4 and not x16 and x1 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and not x4 and not x16 and x1 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x8 and x9 and x3 and not x2 and not x4 and not x16 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and x8 and x9 and not x3 and x4 and x2 ) = '1' then
         y32 <= '1' ;
         current_otherm <= s120;

      elsif ( not x5 and x8 and x9 and not x3 and x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s276;

      elsif ( not x5 and x8 and x9 and not x3 and not x4 and x2 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s321;

      elsif ( not x5 and x8 and x9 and not x3 and not x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and x8 and not x9 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1131;

      elsif ( not x5 and x8 and not x9 and not x6 and x3 and x4 and x2 ) = '1' then
         y45 <= '1' ;
         current_otherm <= s114;

      elsif ( not x5 and x8 and not x9 and not x6 and x3 and x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1253;

      elsif ( not x5 and x8 and not x9 and not x6 and x3 and not x4 and x2 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( not x5 and x8 and not x9 and not x6 and x3 and not x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y37 <= '1' ;
         y39 <= '1' ;
         current_otherm <= s982;

      elsif ( not x5 and x8 and not x9 and not x6 and not x3 and x4 and x2 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s259;

      elsif ( not x5 and x8 and not x9 and not x6 and not x3 and x4 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and x8 and not x9 and not x6 and not x3 and not x4 and x2 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and x8 and not x9 and not x6 and not x3 and not x4 and not x2 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y23 <= '1' ;
         current_otherm <= s1131;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and x4 and x9 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and x4 and x9 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and x4 and x9 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and x4 and x9 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and x4 and not x9 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and not x4 and x9 ) = '1' then
         y16 <= '1' ;
         current_otherm <= s14;

      elsif ( not x5 and not x8 and not x6 and x2 and x3 and not x4 and not x9 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and x4 and x9 ) = '1' then
         y3 <= '1' ;
         y18 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s894;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and x4 and not x9 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and not x4 and x9 and x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and not x4 and x9 and not x13 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and not x4 and x9 and not x13 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and not x4 and x9 and not x13 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and x2 and not x3 and not x4 and not x9 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and x3 and x9 and x14 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and x3 and x9 and not x14 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and x3 and x9 and not x14 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and x3 and x9 and not x14 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and x3 and not x9 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and not x3 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x5 and not x8 and not x6 and not x2 and x4 and not x3 and not x9 ) = '1' then
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1103;

      elsif ( not x5 and not x8 and not x6 and not x2 and not x4 and x9 and x3 and x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( not x5 and not x8 and not x6 and not x2 and not x4 and x9 and x3 and not x12 and x1 and x16 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and x17 ) = '1' then
         y33 <= '1' ;
         current_otherm <= s119;

      elsif ( not x5 and not x8 and not x6 and not x2 and not x4 and x9 and x3 and not x12 and x1 and not x16 and not x17 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and not x2 and not x4 and x9 and x3 and not x12 and not x1 ) = '1' then
         current_otherm <= s1;

      elsif ( not x5 and not x8 and not x6 and not x2 and not x4 and x9 and not x3 ) = '1' then
         y26 <= '1' ;
         current_otherm <= s649;

      else
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s1103;

      end if;

   when s1213 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s405;

   when s1214 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         current_otherm <= s742;

   when s1215 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y13 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1095;

   when s1216 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s460;

   when s1217 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s460;

   when s1218 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         current_otherm <= s460;

   when s1219 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s1254;

   when s1220 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1255;

   when s1221 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s1256;

   when s1222 =>
         y2 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1257;

   when s1223 =>
         y3 <= '1' ;
         current_otherm <= s199;

   when s1224 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_otherm <= s1258;

   when s1225 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s607;

   when s1226 =>
      if ( x11 and x10 and x2 ) = '1' then
         current_otherm <= s1;

      elsif ( x11 and x10 and not x2 and x3 and x4 and x5 and x1 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x11 and x10 and not x2 and x3 and x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y45 <= '1' ;
         y46 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and x3 and x4 and not x5 and x1 ) = '1' then
         y13 <= '1' ;
         current_otherm <= s238;

      elsif ( x11 and x10 and not x2 and x3 and x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and x3 and not x4 and x5 and x1 ) = '1' then
         y51 <= '1' ;
         current_otherm <= s279;

      elsif ( x11 and x10 and not x2 and x3 and not x4 and x5 and not x1 ) = '1' then
         y41 <= '1' ;
         y42 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and x3 and not x4 and not x5 and x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and x3 and not x4 and not x5 and not x1 ) = '1' then
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and x5 and x1 and x6 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and x5 and x1 and not x6 and x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_otherm <= s339;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s340;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y47 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and not x5 and x1 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and not x5 and x1 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s341;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and not x5 and x1 and not x6 and not x7 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and not x3 and x4 and not x5 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and not x3 and not x4 and x1 and x5 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and not x3 and not x4 and x1 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and x10 and not x2 and not x3 and not x4 and not x1 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         y32 <= '1' ;
         y48 <= '1' ;
         current_otherm <= s342;

      elsif ( x11 and not x10 ) = '1' then
         y28 <= '1' ;
         current_otherm <= s780;

      else
         y29 <= '1' ;
         current_otherm <= s1144;

      end if;

   when s1227 =>
         y8 <= '1' ;
         y54 <= '1' ;
         current_otherm <= s1259;

   when s1228 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s460;

   when s1229 =>
         y28 <= '1' ;
         current_otherm <= s780;

   when s1230 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1260;

   when s1231 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1261;

   when s1232 =>
         y2 <= '1' ;
         current_otherm <= s1262;

   when s1233 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1159;

   when s1234 =>
      if ( x64 and x3 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s820;

      elsif ( x64 and not x3 ) = '1' then
         y3 <= '1' ;
         y6 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_otherm <= s1263;

      elsif ( not x64 and x14 and x23 and x24 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and x25 ) = '1' then
         y10 <= '1' ;
         current_otherm <= s16;

      elsif ( not x64 and x14 and x23 and not x24 and not x25 ) = '1' then
         current_otherm <= s1;

      elsif ( not x64 and x14 and not x23 ) = '1' then
         current_otherm <= s1;

      else
         y47 <= '1' ;
         y56 <= '1' ;
         y61 <= '1' ;
         y70 <= '1' ;
         current_otherm <= s931;

      end if;

   when s1235 =>
         y4 <= '1' ;
         y6 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_otherm <= s820;

   when s1236 =>
      if ( x19 and x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1040;

      elsif ( x19 and not x4 and x5 and x6 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1041;

      elsif ( x19 and not x4 and x5 and x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1042;

      elsif ( x19 and not x4 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s958;

      elsif ( x19 and not x4 and not x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s1043;

      else
         y4 <= '1' ;
         y20 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s1044;

      end if;

   when s1237 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

   when s1238 =>
      if ( x5 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      else
         y5 <= '1' ;
         y23 <= '1' ;
         y32 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s958;

      end if;

   when s1239 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s1139;

   when s1240 =>
      if ( x9 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x9 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x9 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x9 and x11 and x10 ) = '1' then
         y9 <= '1' ;
         y21 <= '1' ;
         y30 <= '1' ;
         current_otherm <= s1264;

      elsif ( not x9 and x11 and not x10 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

      elsif ( not x9 and not x11 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1265;

      elsif ( not x9 and not x11 and not x10 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x9 and not x11 and not x10 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x9 and not x11 and not x10 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1241 =>
         y9 <= '1' ;
         y21 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s537;

   when s1242 =>
      if ( x10 and x9 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x10 and x9 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x10 and x9 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and x9 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x9 and x11 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x10 and not x9 and x11 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( x10 and not x9 and x11 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x9 and x11 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( x10 and not x9 and not x11 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         y31 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s864;

      elsif ( not x10 and x9 and x11 and x19 and x13 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x10 and x9 and x11 and x19 and not x13 and x12 ) = '1' then
         y25 <= '1' ;
         current_otherm <= s150;

      elsif ( not x10 and x9 and x11 and x19 and not x13 and not x12 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x9 and x11 and not x19 ) = '1' then
         current_otherm <= s1;

      elsif ( not x10 and x9 and not x11 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s864;

      else
         y5 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s864;

      end if;

   when s1243 =>
      if ( x20 and x14 and x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s668;

      elsif ( x20 and x14 and not x15 ) = '1' then
         y6 <= '1' ;
         y11 <= '1' ;
         y42 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s855;

      elsif ( x20 and not x14 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y44 <= '1' ;
         y45 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1149;

      elsif ( not x20 and x21 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s786;

      elsif ( not x20 and not x21 and x13 ) = '1' then
         y6 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_otherm <= s812;

      elsif ( not x20 and not x21 and not x13 and x14 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s471;

      elsif ( not x20 and not x21 and not x13 and not x14 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x21 and not x13 and not x14 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x20 and not x21 and not x13 and not x14 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1244 =>
         y15 <= '1' ;
         current_otherm <= s426;

   when s1245 =>
         y9 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s1158;

   when s1246 =>
         y2 <= '1' ;
         current_otherm <= s1117;

   when s1247 =>
      if ( x16 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         y42 <= '1' ;
         y50 <= '1' ;
         current_otherm <= s395;

      elsif ( not x16 and x10 and x11 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x16 and x10 and not x11 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( not x16 and x10 and not x11 and not x12 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1248 =>
      if ( x14 and x6 and x5 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and x6 and not x5 and x7 and x8 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s890;

      elsif ( x14 and x6 and not x5 and x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y19 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_otherm <= s914;

      elsif ( x14 and x6 and not x5 and x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x14 and x6 and not x5 and not x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_otherm <= s508;

      elsif ( x14 and not x6 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s890;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y40 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s915;

      end if;

   when s1249 =>
      if ( x63 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1266;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s1267;

      end if;

   when s1250 =>
      if ( x13 and x8 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and x8 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and x8 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x8 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x8 and not x9 and x11 and x10 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and x8 and not x9 and x11 and x10 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and x8 and not x9 and x11 and x10 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x8 and not x9 and x11 and x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x8 and not x9 and x11 and not x10 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s504;

      elsif ( x13 and x8 and not x9 and not x11 and x10 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1114;

      elsif ( x13 and x8 and not x9 and not x11 and not x10 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and x8 and not x9 and not x11 and not x10 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and x8 and not x9 and not x11 and not x10 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and x8 and not x9 and not x11 and not x10 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and x10 and x11 and x9 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and x10 and x11 and x9 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and x10 and x11 and x9 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and x10 and x11 and x9 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and x10 and x11 and not x9 and x18 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and x10 and x11 and not x9 and not x18 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and x10 and not x11 and x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s391;

      elsif ( x13 and not x8 and x6 and x10 and not x11 and not x9 and x17 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and x10 and not x11 and not x9 and not x17 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and not x10 and x11 and x9 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1115;

      elsif ( x13 and not x8 and x6 and not x10 and x11 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x13 and not x8 and x6 and not x10 and not x11 and x9 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y40 <= '1' ;
         current_otherm <= s769;

      elsif ( x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and x15 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and not x15 and x16 ) = '1' then
         y46 <= '1' ;
         current_otherm <= s110;

      elsif ( x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and x14 and not x15 and not x16 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and not x10 and not x11 and x9 and not x19 and not x14 ) = '1' then
         current_otherm <= s1;

      elsif ( x13 and not x8 and x6 and not x10 and not x11 and not x9 ) = '1' then
         y44 <= '1' ;
         current_otherm <= s562;

      elsif ( x13 and not x8 and not x6 ) = '1' then
         y2 <= '1' ;
         current_otherm <= s1023;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1116;

      end if;

   when s1251 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1209;

   when s1252 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1268;

   when s1253 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s1269;

   when s1254 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y50 <= '1' ;
         y52 <= '1' ;
         current_otherm <= s460;

   when s1255 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y47 <= '1' ;
         y51 <= '1' ;
         current_otherm <= s460;

   when s1256 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y32 <= '1' ;
         y38 <= '1' ;
         current_otherm <= s460;

   when s1257 =>
      if ( x14 ) = '1' then
         y22 <= '1' ;
         current_otherm <= s92;

      elsif ( not x14 and x22 and x21 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x14 and x22 and not x21 and x18 ) = '1' then
         y52 <= '1' ;
         current_otherm <= s360;

      elsif ( not x14 and x22 and not x21 and not x18 ) = '1' then
         current_otherm <= s1;

      else
         current_otherm <= s1;

      end if;

   when s1258 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_otherm <= s146;

   when s1259 =>
         y13 <= '1' ;
         y55 <= '1' ;
         y56 <= '1' ;
         current_otherm <= s1;

   when s1260 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1270;

   when s1261 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_otherm <= s1271;

   when s1262 =>
         y9 <= '1' ;
         y14 <= '1' ;
         y17 <= '1' ;
         y26 <= '1' ;
         y49 <= '1' ;
         current_otherm <= s709;

   when s1263 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y20 <= '1' ;
         current_otherm <= s1165;

   when s1264 =>
         y2 <= '1' ;
         y9 <= '1' ;
         y21 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1272;

   when s1265 =>
         y9 <= '1' ;
         y21 <= '1' ;
         y41 <= '1' ;
         y45 <= '1' ;
         current_otherm <= s1273;

   when s1266 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y29 <= '1' ;
         current_otherm <= s1274;

   when s1267 =>
         y2 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         current_otherm <= s1275;

   when s1268 =>
         y2 <= '1' ;
         y15 <= '1' ;
         y31 <= '1' ;
         current_otherm <= s793;

   when s1269 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y39 <= '1' ;
         y41 <= '1' ;
         current_otherm <= s1103;

   when s1270 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s908;

   when s1271 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s735;

   when s1272 =>
         y5 <= '1' ;
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_otherm <= s864;

   when s1273 =>
         y9 <= '1' ;
         y21 <= '1' ;
         y44 <= '1' ;
         current_otherm <= s864;

   when s1274 =>
      if ( x14 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x14 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_otherm <= s122;

      elsif ( x14 and x16 and not x12 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x14 and not x16 ) = '1' then
         current_otherm <= s1;

      else
         y9 <= '1' ;
         current_otherm <= s43;

      end if;

   when s1275 =>
      if ( x9 and x6 and x12 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s790;

      elsif ( x9 and x6 and not x12 and x11 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y14 <= '1' ;
         y35 <= '1' ;
         current_otherm <= s410;

      elsif ( x9 and x6 and not x12 and not x11 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and x6 and not x12 and not x11 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and x6 and not x12 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and x6 and not x12 and not x11 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and x11 and x12 and x10 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and x11 and x12 and x10 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and x11 and x12 and x10 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and x11 and x12 and x10 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and x11 and x12 and not x10 and x16 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and x11 and x12 and not x10 and not x16 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and x11 and not x12 and x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s791;

      elsif ( x9 and not x6 and x8 and x11 and not x12 and not x10 and x17 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and x11 and not x12 and not x10 and not x17 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and not x11 and x12 and x10 ) = '1' then
         y2 <= '1' ;
         y31 <= '1' ;
         y34 <= '1' ;
         current_otherm <= s792;

      elsif ( x9 and not x6 and x8 and not x11 and x12 and not x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( x9 and not x6 and x8 and not x11 and not x12 and x10 and x15 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y16 <= '1' ;
         current_otherm <= s408;

      elsif ( x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and x14 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and not x14 and x13 ) = '1' then
         y56 <= '1' ;
         current_otherm <= s412;

      elsif ( x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and x18 and not x14 and not x13 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and not x11 and not x12 and x10 and not x15 and not x18 ) = '1' then
         current_otherm <= s1;

      elsif ( x9 and not x6 and x8 and not x11 and not x12 and not x10 ) = '1' then
         y57 <= '1' ;
         current_otherm <= s135;

      elsif ( x9 and not x6 and not x8 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_otherm <= s790;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y28 <= '1' ;
         y33 <= '1' ;
         current_otherm <= s477;

      end if;

   end case;
   end proc_otherm;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;	y46  <= '0' ;	y47  <= '0' ;	y48  <= '0' ;
	y49  <= '0' ;	y50  <= '0' ;	y51  <= '0' ;	y52  <= '0' ;
	y53  <= '0' ;	y54  <= '0' ;	y55  <= '0' ;	y56  <= '0' ;
	y57  <= '0' ;	y58  <= '0' ;	y59  <= '0' ;	y60  <= '0' ;
	y61  <= '0' ;	y62  <= '0' ;	y63  <= '0' ;	y64  <= '0' ;
	y65  <= '0' ;	y66  <= '0' ;	y67  <= '0' ;	y68  <= '0' ;
	y69  <= '0' ;	y70  <= '0' ;	y71  <= '0' ;	y72  <= '0' ;
	y73  <= '0' ;	y74  <= '0' ;	y75  <= '0' ;	y77  <= '0' ;
	y78  <= '0' ;	y79  <= '0' ;	y80  <= '0' ;	y81  <= '0' ;
	y84  <= '0' ;	y86  <= '0' ;	y88  <= '0' ;	y90  <= '0' ;
	y91  <= '0' ;	y92  <= '0' ;	y93  <= '0' ;	y94  <= '0' ;
	y95  <= '0' ;	y96  <= '0' ;	y97  <= '0' ;	y98  <= '0' ;
	y99  <= '0' ;	y100 <= '0' ;	y102 <= '0' ;	y110 <= '0' ;

	current_otherm <= s1;
      elsif (clk'event and clk ='1') then
        proc_otherm;
      end if;
   end process;
end ARC;
