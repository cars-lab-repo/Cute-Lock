library ieee;
use ieee.std_logic_1164.all;

entity e4 is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,
	x31 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24 : out std_logic );
end e4;

architecture ARC of e4 is

   type states_e4 is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24 );
   signal current_e4 : states_e4;

begin
   process (clk , rst)
   procedure proc_e4 is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;


   case current_e4 is
   when s1 =>
      if ( x10 and x12 and x23 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_e4 <= s2;

      elsif ( x10 and x12 and not x23 and x4 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s3;

      elsif ( x10 and x12 and not x23 and not x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      elsif ( x10 and not x12 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s6;

      elsif ( not x10 and x1 and x22 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y12 <= '1' ;
         current_e4 <= s7;

      elsif ( not x10 and x1 and not x22 and x2 and x3 and x11 ) = '1' then
         current_e4 <= s1;

      elsif ( not x10 and x1 and not x22 and x2 and x3 and not x11 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( not x10 and x1 and not x22 and x2 and not x3 and x11 and x5 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( not x10 and x1 and not x22 and x2 and not x3 and x11 and not x5 ) = '1' then
         y1 <= '1' ;
         current_e4 <= s10;

      elsif ( not x10 and x1 and not x22 and x2 and not x3 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s3;

      elsif ( not x10 and x1 and not x22 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_e4 <= s5;

      elsif ( not x10 and not x1 and x11 and x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      elsif ( not x10 and not x1 and x11 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      else
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      end if;

   when s2 =>
      if ( x19 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s11;

      elsif ( not x19 and x26 and x5 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      elsif ( not x19 and x26 and not x5 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_e4 <= s13;

      else
         y7 <= '1' ;
         y11 <= '1' ;
         current_e4 <= s14;

      end if;

   when s3 =>
      if ( x19 and x28 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s14;

      elsif ( x19 and x28 and not x1 and x15 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x19 and x28 and not x1 and not x15 ) = '1' then
         y1 <= '1' ;
         current_e4 <= s10;

      elsif ( x19 and not x28 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      else
         y1 <= '1' ;
         current_e4 <= s10;

      end if;

   when s4 =>
      if ( x30 and x16 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s15;

      elsif ( x30 and x16 and not x6 and x8 and x19 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s11;

      elsif ( x30 and x16 and not x6 and x8 and not x19 and x26 and x5 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      elsif ( x30 and x16 and not x6 and x8 and not x19 and x26 and not x5 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_e4 <= s13;

      elsif ( x30 and x16 and not x6 and x8 and not x19 and not x26 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_e4 <= s14;

      elsif ( x30 and x16 and not x6 and not x8 ) = '1' then
         current_e4 <= s1;

      elsif ( x30 and not x16 and x10 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x30 and not x16 and not x10 ) = '1' then
         current_e4 <= s1;

      elsif ( not x30 and x5 and x9 ) = '1' then
         current_e4 <= s1;

      elsif ( not x30 and x5 and not x9 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_e4 <= s16;

      elsif ( not x30 and not x5 and x3 and x11 ) = '1' then
         current_e4 <= s4;

      elsif ( not x30 and not x5 and x3 and not x11 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( not x30 and not x5 and not x3 and x11 ) = '1' then
         y1 <= '1' ;
         current_e4 <= s10;

      else
         y9 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s3;

      end if;

   when s5 =>
      if ( x11 and x25 and x3 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s3;

      elsif ( x11 and x25 and not x3 and x5 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      elsif ( x11 and x25 and not x3 and not x5 ) = '1' then
         current_e4 <= s5;

      elsif ( x11 and not x25 ) = '1' then
         y1 <= '1' ;
         current_e4 <= s10;

      else
         y9 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s3;

      end if;

   when s6 =>
      if ( x12 and x27 and x20 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( x12 and x27 and not x20 and x13 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      elsif ( x12 and x27 and not x20 and not x13 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x12 and not x27 and x29 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_e4 <= s18;

      elsif ( x12 and not x27 and x29 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( x12 and not x27 and not x29 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s11;

      elsif ( x12 and not x27 and not x29 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s20;

      elsif ( not x12 and x29 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s11;

      else
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s21;

      end if;

   when s7 =>
      if ( x2 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      else
         y11 <= '1' ;
         y23 <= '1' ;
         current_e4 <= s19;

      end if;

   when s8 =>
      if ( x14 and x8 and x10 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x14 and x8 and not x10 ) = '1' then
         current_e4 <= s1;

      elsif ( x14 and not x8 and x30 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_e4 <= s18;

      elsif ( x14 and not x8 and x30 and not x1 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      elsif ( x14 and not x8 and x30 and not x1 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_e4 <= s19;

      elsif ( x14 and not x8 and not x30 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( not x14 and x3 and x21 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_e4 <= s13;

      elsif ( not x14 and x3 and not x21 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      end if;

   when s9 =>
      if ( x24 and x26 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s20;

      elsif ( x24 and x26 and not x7 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s22;

      elsif ( x24 and not x26 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_e4 <= s19;

      elsif ( not x24 and x28 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s6;

      else
         current_e4 <= s1;

      end if;

   when s10 =>
      if ( x19 and x13 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_e4 <= s16;

      elsif ( x19 and not x13 and x21 and x18 and x12 ) = '1' then
         current_e4 <= s10;

      elsif ( x19 and not x13 and x21 and x18 and not x12 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_e4 <= s19;

      elsif ( x19 and not x13 and x21 and not x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( x19 and not x13 and not x21 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      else
         current_e4 <= s1;

      end if;

   when s11 =>
      if ( x2 and x8 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s14;

      elsif ( x2 and x8 and not x1 and x15 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x2 and x8 and not x1 and not x15 ) = '1' then
         y1 <= '1' ;
         current_e4 <= s10;

      elsif ( x2 and not x8 and x21 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_e4 <= s18;

      elsif ( x2 and not x8 and x21 and not x1 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      elsif ( x2 and not x8 and x21 and not x1 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_e4 <= s19;

      elsif ( x2 and not x8 and not x21 ) = '1' then
         y1 <= '1' ;
         current_e4 <= s10;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      end if;

   when s12 =>
      if ( x16 and x19 and x20 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( x16 and x19 and not x20 and x13 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      elsif ( x16 and x19 and not x20 and not x13 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x16 and not x19 and x30 and x26 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_e4 <= s18;

      elsif ( x16 and not x19 and x30 and x26 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( x16 and not x19 and x30 and not x26 and x3 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( x16 and not x19 and x30 and not x26 and not x3 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_e4 <= s18;

      elsif ( x16 and not x19 and x30 and not x26 and not x3 and not x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( x16 and not x19 and not x30 and x8 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( x16 and not x19 and not x30 and not x8 ) = '1' then
         current_e4 <= s1;

      else
         current_e4 <= s1;

      end if;

   when s13 =>
      if ( x10 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_e4 <= s19;

      elsif ( not x10 and x25 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s20;

      else
         y12 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s21;

      end if;

   when s14 =>
      if ( x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s14;

      elsif ( not x1 and x15 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      else
         y1 <= '1' ;
         current_e4 <= s10;

      end if;

   when s15 =>
      if ( x16 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s15;

      elsif ( x16 and not x6 and x8 and x19 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s11;

      elsif ( x16 and not x6 and x8 and not x19 and x26 and x5 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      elsif ( x16 and not x6 and x8 and not x19 and x26 and not x5 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_e4 <= s13;

      elsif ( x16 and not x6 and x8 and not x19 and not x26 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_e4 <= s14;

      elsif ( x16 and not x6 and not x8 ) = '1' then
         current_e4 <= s1;

      elsif ( not x16 and x10 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      else
         current_e4 <= s1;

      end if;

   when s16 =>
      if ( x9 ) = '1' then
         y13 <= '1' ;
         current_e4 <= s23;

      elsif ( not x9 and x3 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      else
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      end if;

   when s17 =>
      if ( x22 and x2 and x20 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( x22 and x2 and not x20 and x13 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      elsif ( x22 and x2 and not x20 and not x13 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x22 and not x2 ) = '1' then
         current_e4 <= s1;

      elsif ( not x22 and x31 ) = '1' then
         current_e4 <= s1;

      else
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      end if;

   when s18 =>
      if ( x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      elsif ( not x5 and x17 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s12;

      else
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      end if;

   when s19 =>
      if ( x25 and x22 ) = '1' then
         current_e4 <= s1;

      elsif ( x25 and not x22 and x6 and x8 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( x25 and not x22 and x6 and not x8 ) = '1' then
         current_e4 <= s1;

      elsif ( x25 and not x22 and not x6 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_e4 <= s13;

      elsif ( not x25 and x29 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y12 <= '1' ;
         current_e4 <= s7;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_e4 <= s18;

      end if;

   when s20 =>
      if ( x7 and x15 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s14;

      elsif ( x7 and x15 and not x1 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      elsif ( x7 and not x15 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      else
         y7 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s24;

      end if;

   when s21 =>
      if ( x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_e4 <= s8;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s11;

      end if;

   when s22 =>
      if ( x16 and x9 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_e4 <= s15;

      elsif ( x16 and not x9 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_e4 <= s14;

      else
         y17 <= '1' ;
         y20 <= '1' ;
         current_e4 <= s6;

      end if;

   when s23 =>
      if ( x20 ) = '1' then
         y14 <= '1' ;
         y22 <= '1' ;
         current_e4 <= s17;

      elsif ( not x20 and x13 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_e4 <= s4;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

      end if;

   when s24 =>
         y11 <= '1' ;
         y18 <= '1' ;
         current_e4 <= s9;

   end case;
   end proc_e4;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;

	current_e4 <= s1;
      elsif (clk'event and clk ='1') then
        proc_e4;
      end if;
   end process;
end ARC;
