// Benchmark "./test_runs/structural2_nkeys_nbits--s-120240927_165956/ITC99/b22_encrypted" written by ABC on Fri Sep 27 18:34:51 2024

module b22_encrypted  ( clock, 
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, keyinput0, keyinput1, keyinput2,
    keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
    keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
    keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20,
    keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26,
    keyinput27, keyinput28, keyinput29, keyinput30, keyinput31,
    SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28  );
  input  clock;
  input  SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_,
    SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_,
    SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_,
    SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, keyinput0, keyinput1,
    keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
    keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
    keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
    keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25,
    keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28;
  reg P1_IR_REG_0_, P1_IR_REG_1_, P1_IR_REG_2_, P1_IR_REG_3_, P1_IR_REG_4_,
    P1_IR_REG_5_, P1_IR_REG_6_, P1_IR_REG_7_, P1_IR_REG_8_, P1_IR_REG_9_,
    P1_IR_REG_10_, P1_IR_REG_11_, P1_IR_REG_12_, P1_IR_REG_13_,
    P1_IR_REG_14_, P1_IR_REG_15_, P1_IR_REG_16_, P1_IR_REG_17_,
    P1_IR_REG_18_, P1_IR_REG_19_, P1_IR_REG_20_, P1_IR_REG_21_,
    P1_IR_REG_22_, P1_IR_REG_23_, P1_IR_REG_24_, P1_IR_REG_25_,
    P1_IR_REG_26_, P1_IR_REG_27_, P1_IR_REG_28_, P1_IR_REG_29_,
    P1_IR_REG_30_, P1_IR_REG_31_, P1_D_REG_0_, P1_D_REG_1_, P1_D_REG_2_,
    P1_D_REG_3_, P1_D_REG_4_, P1_D_REG_5_, P1_D_REG_6_, P1_D_REG_7_,
    P1_D_REG_8_, P1_D_REG_9_, P1_D_REG_10_, P1_D_REG_11_, P1_D_REG_12_,
    P1_D_REG_13_, P1_D_REG_14_, P1_D_REG_15_, P1_D_REG_16_, P1_D_REG_17_,
    P1_D_REG_18_, P1_D_REG_19_, P1_D_REG_20_, P1_D_REG_21_, P1_D_REG_22_,
    P1_D_REG_23_, P1_D_REG_24_, P1_D_REG_25_, P1_D_REG_26_, P1_D_REG_27_,
    P1_D_REG_28_, P1_D_REG_29_, P1_D_REG_30_, P1_D_REG_31_, P1_REG0_REG_0_,
    P1_REG0_REG_1_, P1_REG0_REG_2_, P1_REG0_REG_3_, P1_REG0_REG_4_,
    P1_REG0_REG_5_, P1_REG0_REG_6_, P1_REG0_REG_7_, P1_REG0_REG_8_,
    P1_REG0_REG_9_, P1_REG0_REG_10_, P1_REG0_REG_11_, P1_REG0_REG_12_,
    P1_REG0_REG_13_, P1_REG0_REG_14_, P1_REG0_REG_15_, P1_REG0_REG_16_,
    P1_REG0_REG_17_, P1_REG0_REG_18_, P1_REG0_REG_19_, P1_REG0_REG_20_,
    P1_REG0_REG_21_, P1_REG0_REG_22_, P1_REG0_REG_23_, P1_REG0_REG_24_,
    P1_REG0_REG_25_, P1_REG0_REG_26_, P1_REG0_REG_27_, P1_REG0_REG_28_,
    P1_REG0_REG_29_, P1_REG0_REG_30_, P1_REG0_REG_31_, P1_REG1_REG_0_,
    P1_REG1_REG_1_, P1_REG1_REG_2_, P1_REG1_REG_3_, P1_REG1_REG_4_,
    P1_REG1_REG_5_, P1_REG1_REG_6_, P1_REG1_REG_7_, P1_REG1_REG_8_,
    P1_REG1_REG_9_, P1_REG1_REG_10_, P1_REG1_REG_11_, P1_REG1_REG_12_,
    P1_REG1_REG_13_, P1_REG1_REG_14_, P1_REG1_REG_15_, P1_REG1_REG_16_,
    P1_REG1_REG_17_, P1_REG1_REG_18_, P1_REG1_REG_19_, P1_REG1_REG_20_,
    P1_REG1_REG_21_, P1_REG1_REG_22_, P1_REG1_REG_23_, P1_REG1_REG_24_,
    P1_REG1_REG_25_, P1_REG1_REG_26_, P1_REG1_REG_27_, P1_REG1_REG_28_,
    P1_REG1_REG_29_, P1_REG1_REG_30_, P1_REG1_REG_31_, P1_REG2_REG_0_,
    P1_REG2_REG_1_, P1_REG2_REG_2_, P1_REG2_REG_3_, P1_REG2_REG_4_,
    P1_REG2_REG_5_, P1_REG2_REG_6_, P1_REG2_REG_7_, P1_REG2_REG_8_,
    P1_REG2_REG_9_, P1_REG2_REG_10_, P1_REG2_REG_11_, P1_REG2_REG_12_,
    P1_REG2_REG_13_, P1_REG2_REG_14_, P1_REG2_REG_15_, P1_REG2_REG_16_,
    P1_REG2_REG_17_, P1_REG2_REG_18_, P1_REG2_REG_19_, P1_REG2_REG_20_,
    P1_REG2_REG_21_, P1_REG2_REG_22_, P1_REG2_REG_23_, P1_REG2_REG_24_,
    P1_REG2_REG_25_, P1_REG2_REG_26_, P1_REG2_REG_27_, P1_REG2_REG_28_,
    P1_REG2_REG_29_, P1_REG2_REG_30_, P1_REG2_REG_31_, P1_ADDR_REG_19_,
    P1_ADDR_REG_18_, P1_ADDR_REG_17_, P1_ADDR_REG_16_, P1_ADDR_REG_15_,
    P1_ADDR_REG_14_, P1_ADDR_REG_13_, P1_ADDR_REG_12_, P1_ADDR_REG_11_,
    P1_ADDR_REG_10_, P1_ADDR_REG_9_, P1_ADDR_REG_8_, P1_ADDR_REG_7_,
    P1_ADDR_REG_6_, P1_ADDR_REG_5_, P1_ADDR_REG_4_, P1_ADDR_REG_3_,
    P1_ADDR_REG_2_, P1_ADDR_REG_1_, P1_ADDR_REG_0_, P1_DATAO_REG_0_,
    P1_DATAO_REG_1_, P1_DATAO_REG_2_, P1_DATAO_REG_3_, P1_DATAO_REG_4_,
    P1_DATAO_REG_5_, P1_DATAO_REG_6_, P1_DATAO_REG_7_, P1_DATAO_REG_8_,
    P1_DATAO_REG_9_, P1_DATAO_REG_10_, P1_DATAO_REG_11_, P1_DATAO_REG_12_,
    P1_DATAO_REG_13_, P1_DATAO_REG_14_, P1_DATAO_REG_15_, P1_DATAO_REG_16_,
    P1_DATAO_REG_17_, P1_DATAO_REG_18_, P1_DATAO_REG_19_, P1_DATAO_REG_20_,
    P1_DATAO_REG_21_, P1_DATAO_REG_22_, P1_DATAO_REG_23_, P1_DATAO_REG_24_,
    P1_DATAO_REG_25_, P1_DATAO_REG_26_, P1_DATAO_REG_27_, P1_DATAO_REG_28_,
    P1_DATAO_REG_29_, P1_DATAO_REG_30_, P1_DATAO_REG_31_, P1_B_REG,
    P1_REG3_REG_15_, P1_REG3_REG_26_, P1_REG3_REG_6_, P1_REG3_REG_18_,
    P1_REG3_REG_2_, P1_REG3_REG_11_, P1_REG3_REG_22_, P1_REG3_REG_13_,
    P1_REG3_REG_20_, P1_REG3_REG_0_, P1_REG3_REG_9_, P1_REG3_REG_4_,
    P1_REG3_REG_24_, P1_REG3_REG_17_, P1_REG3_REG_5_, P1_REG3_REG_16_,
    P1_REG3_REG_25_, P1_REG3_REG_12_, P1_REG3_REG_21_, P1_REG3_REG_1_,
    P1_REG3_REG_8_, P1_REG3_REG_28_, P1_REG3_REG_19_, P1_REG3_REG_3_,
    P1_REG3_REG_10_, P1_REG3_REG_23_, P1_REG3_REG_14_, P1_REG3_REG_27_,
    P1_REG3_REG_7_, P1_STATE_REG, P1_RD_REG, P1_WR_REG, P2_IR_REG_0_,
    P2_IR_REG_1_, P2_IR_REG_2_, P2_IR_REG_3_, P2_IR_REG_4_, P2_IR_REG_5_,
    P2_IR_REG_6_, P2_IR_REG_7_, P2_IR_REG_8_, P2_IR_REG_9_, P2_IR_REG_10_,
    P2_IR_REG_11_, P2_IR_REG_12_, P2_IR_REG_13_, P2_IR_REG_14_,
    P2_IR_REG_15_, P2_IR_REG_16_, P2_IR_REG_17_, P2_IR_REG_18_,
    P2_IR_REG_19_, P2_IR_REG_20_, P2_IR_REG_21_, P2_IR_REG_22_,
    P2_IR_REG_23_, P2_IR_REG_24_, P2_IR_REG_25_, P2_IR_REG_26_,
    P2_IR_REG_27_, P2_IR_REG_28_, P2_IR_REG_29_, P2_IR_REG_30_,
    P2_IR_REG_31_, P2_D_REG_0_, P2_D_REG_1_, P2_D_REG_2_, P2_D_REG_3_,
    P2_D_REG_4_, P2_D_REG_5_, P2_D_REG_6_, P2_D_REG_7_, P2_D_REG_8_,
    P2_D_REG_9_, P2_D_REG_10_, P2_D_REG_11_, P2_D_REG_12_, P2_D_REG_13_,
    P2_D_REG_14_, P2_D_REG_15_, P2_D_REG_16_, P2_D_REG_17_, P2_D_REG_18_,
    P2_D_REG_19_, P2_D_REG_20_, P2_D_REG_21_, P2_D_REG_22_, P2_D_REG_23_,
    P2_D_REG_24_, P2_D_REG_25_, P2_D_REG_26_, P2_D_REG_27_, P2_D_REG_28_,
    P2_D_REG_29_, P2_D_REG_30_, P2_D_REG_31_, P2_REG0_REG_0_,
    P2_REG0_REG_1_, P2_REG0_REG_2_, P2_REG0_REG_3_, P2_REG0_REG_4_,
    P2_REG0_REG_5_, P2_REG0_REG_6_, P2_REG0_REG_7_, P2_REG0_REG_8_,
    P2_REG0_REG_9_, P2_REG0_REG_10_, P2_REG0_REG_11_, P2_REG0_REG_12_,
    P2_REG0_REG_13_, P2_REG0_REG_14_, P2_REG0_REG_15_, P2_REG0_REG_16_,
    P2_REG0_REG_17_, P2_REG0_REG_18_, P2_REG0_REG_19_, P2_REG0_REG_20_,
    P2_REG0_REG_21_, P2_REG0_REG_22_, P2_REG0_REG_23_, P2_REG0_REG_24_,
    P2_REG0_REG_25_, P2_REG0_REG_26_, P2_REG0_REG_27_, P2_REG0_REG_28_,
    P2_REG0_REG_29_, P2_REG0_REG_30_, P2_REG0_REG_31_, P2_REG1_REG_0_,
    P2_REG1_REG_1_, P2_REG1_REG_2_, P2_REG1_REG_3_, P2_REG1_REG_4_,
    P2_REG1_REG_5_, P2_REG1_REG_6_, P2_REG1_REG_7_, P2_REG1_REG_8_,
    P2_REG1_REG_9_, P2_REG1_REG_10_, P2_REG1_REG_11_, P2_REG1_REG_12_,
    P2_REG1_REG_13_, P2_REG1_REG_14_, P2_REG1_REG_15_, P2_REG1_REG_16_,
    P2_REG1_REG_17_, P2_REG1_REG_18_, P2_REG1_REG_19_, P2_REG1_REG_20_,
    P2_REG1_REG_21_, P2_REG1_REG_22_, P2_REG1_REG_23_, P2_REG1_REG_24_,
    P2_REG1_REG_25_, P2_REG1_REG_26_, P2_REG1_REG_27_, P2_REG1_REG_28_,
    P2_REG1_REG_29_, P2_REG1_REG_30_, P2_REG1_REG_31_, P2_REG2_REG_0_,
    P2_REG2_REG_1_, P2_REG2_REG_2_, P2_REG2_REG_3_, P2_REG2_REG_4_,
    P2_REG2_REG_5_, P2_REG2_REG_6_, P2_REG2_REG_7_, P2_REG2_REG_8_,
    P2_REG2_REG_9_, P2_REG2_REG_10_, P2_REG2_REG_11_, P2_REG2_REG_12_,
    P2_REG2_REG_13_, P2_REG2_REG_14_, P2_REG2_REG_15_, P2_REG2_REG_16_,
    P2_REG2_REG_17_, P2_REG2_REG_18_, P2_REG2_REG_19_, P2_REG2_REG_20_,
    P2_REG2_REG_21_, P2_REG2_REG_22_, P2_REG2_REG_23_, P2_REG2_REG_24_,
    P2_REG2_REG_25_, P2_REG2_REG_26_, P2_REG2_REG_27_, P2_REG2_REG_28_,
    P2_REG2_REG_29_, P2_REG2_REG_30_, P2_REG2_REG_31_, P2_ADDR_REG_19_,
    P2_ADDR_REG_18_, P2_ADDR_REG_17_, P2_ADDR_REG_16_, P2_ADDR_REG_15_,
    P2_ADDR_REG_14_, P2_ADDR_REG_13_, P2_ADDR_REG_12_, P2_ADDR_REG_11_,
    P2_ADDR_REG_10_, P2_ADDR_REG_9_, P2_ADDR_REG_8_, P2_ADDR_REG_7_,
    P2_ADDR_REG_6_, P2_ADDR_REG_5_, P2_ADDR_REG_4_, P2_ADDR_REG_3_,
    P2_ADDR_REG_2_, P2_ADDR_REG_1_, P2_ADDR_REG_0_, P2_DATAO_REG_0_,
    P2_DATAO_REG_1_, P2_DATAO_REG_2_, P2_DATAO_REG_3_, P2_DATAO_REG_4_,
    P2_DATAO_REG_5_, P2_DATAO_REG_6_, P2_DATAO_REG_7_, P2_DATAO_REG_8_,
    P2_DATAO_REG_9_, P2_DATAO_REG_10_, P2_DATAO_REG_11_, P2_DATAO_REG_12_,
    P2_DATAO_REG_13_, P2_DATAO_REG_14_, P2_DATAO_REG_15_, P2_DATAO_REG_16_,
    P2_DATAO_REG_17_, P2_DATAO_REG_18_, P2_DATAO_REG_19_, P2_DATAO_REG_20_,
    P2_DATAO_REG_21_, P2_DATAO_REG_22_, P2_DATAO_REG_23_, P2_DATAO_REG_24_,
    P2_DATAO_REG_25_, P2_DATAO_REG_26_, P2_DATAO_REG_27_, P2_DATAO_REG_28_,
    P2_DATAO_REG_29_, P2_DATAO_REG_30_, P2_DATAO_REG_31_, P2_B_REG,
    P2_REG3_REG_15_, P2_REG3_REG_26_, P2_REG3_REG_6_, P2_REG3_REG_18_,
    P2_REG3_REG_2_, P2_REG3_REG_11_, P2_REG3_REG_22_, P2_REG3_REG_13_,
    P2_REG3_REG_20_, P2_REG3_REG_0_, P2_REG3_REG_9_, P2_REG3_REG_4_,
    P2_REG3_REG_24_, P2_REG3_REG_17_, P2_REG3_REG_5_, P2_REG3_REG_16_,
    P2_REG3_REG_25_, P2_REG3_REG_12_, P2_REG3_REG_21_, P2_REG3_REG_1_,
    P2_REG3_REG_8_, P2_REG3_REG_28_, P2_REG3_REG_19_, P2_REG3_REG_3_,
    P2_REG3_REG_10_, P2_REG3_REG_23_, P2_REG3_REG_14_, P2_REG3_REG_27_,
    P2_REG3_REG_7_, P2_STATE_REG, P2_RD_REG, P2_WR_REG, P3_IR_REG_0_,
    P3_IR_REG_1_, P3_IR_REG_2_, P3_IR_REG_3_, P3_IR_REG_4_, P3_IR_REG_5_,
    P3_IR_REG_6_, P3_IR_REG_7_, P3_IR_REG_8_, P3_IR_REG_9_, P3_IR_REG_10_,
    P3_IR_REG_11_, P3_IR_REG_12_, P3_IR_REG_13_, P3_IR_REG_14_,
    P3_IR_REG_15_, P3_IR_REG_16_, P3_IR_REG_17_, P3_IR_REG_18_,
    P3_IR_REG_19_, P3_IR_REG_20_, P3_IR_REG_21_, P3_IR_REG_22_,
    P3_IR_REG_23_, P3_IR_REG_24_, P3_IR_REG_25_, P3_IR_REG_26_,
    P3_IR_REG_27_, P3_IR_REG_28_, P3_IR_REG_29_, P3_IR_REG_30_,
    P3_IR_REG_31_, P3_D_REG_0_, P3_D_REG_1_, P3_D_REG_2_, P3_D_REG_3_,
    P3_D_REG_4_, P3_D_REG_5_, P3_D_REG_6_, P3_D_REG_7_, P3_D_REG_8_,
    P3_D_REG_9_, P3_D_REG_10_, P3_D_REG_11_, P3_D_REG_12_, P3_D_REG_13_,
    P3_D_REG_14_, P3_D_REG_15_, P3_D_REG_16_, P3_D_REG_17_, P3_D_REG_18_,
    P3_D_REG_19_, P3_D_REG_20_, P3_D_REG_21_, P3_D_REG_22_, P3_D_REG_23_,
    P3_D_REG_24_, P3_D_REG_25_, P3_D_REG_26_, P3_D_REG_27_, P3_D_REG_28_,
    P3_D_REG_29_, P3_D_REG_30_, P3_D_REG_31_, P3_REG0_REG_0_,
    P3_REG0_REG_1_, P3_REG0_REG_2_, P3_REG0_REG_3_, P3_REG0_REG_4_,
    P3_REG0_REG_5_, P3_REG0_REG_6_, P3_REG0_REG_7_, P3_REG0_REG_8_,
    P3_REG0_REG_9_, P3_REG0_REG_10_, P3_REG0_REG_11_, P3_REG0_REG_12_,
    P3_REG0_REG_13_, P3_REG0_REG_14_, P3_REG0_REG_15_, P3_REG0_REG_16_,
    P3_REG0_REG_17_, P3_REG0_REG_18_, P3_REG0_REG_19_, P3_REG0_REG_20_,
    P3_REG0_REG_21_, P3_REG0_REG_22_, P3_REG0_REG_23_, P3_REG0_REG_24_,
    P3_REG0_REG_25_, P3_REG0_REG_26_, P3_REG0_REG_27_, P3_REG0_REG_28_,
    P3_REG0_REG_29_, P3_REG0_REG_30_, P3_REG0_REG_31_, P3_REG1_REG_0_,
    P3_REG1_REG_1_, P3_REG1_REG_2_, P3_REG1_REG_3_, P3_REG1_REG_4_,
    P3_REG1_REG_5_, P3_REG1_REG_6_, P3_REG1_REG_7_, P3_REG1_REG_8_,
    P3_REG1_REG_9_, P3_REG1_REG_10_, P3_REG1_REG_11_, P3_REG1_REG_12_,
    P3_REG1_REG_13_, P3_REG1_REG_14_, P3_REG1_REG_15_, P3_REG1_REG_16_,
    P3_REG1_REG_17_, P3_REG1_REG_18_, P3_REG1_REG_19_, P3_REG1_REG_20_,
    P3_REG1_REG_21_, P3_REG1_REG_22_, P3_REG1_REG_23_, P3_REG1_REG_24_,
    P3_REG1_REG_25_, P3_REG1_REG_26_, P3_REG1_REG_27_, P3_REG1_REG_28_,
    P3_REG1_REG_29_, P3_REG1_REG_30_, P3_REG1_REG_31_, P3_REG2_REG_0_,
    P3_REG2_REG_1_, P3_REG2_REG_2_, P3_REG2_REG_3_, P3_REG2_REG_4_,
    P3_REG2_REG_5_, P3_REG2_REG_6_, P3_REG2_REG_7_, P3_REG2_REG_8_,
    P3_REG2_REG_9_, P3_REG2_REG_10_, P3_REG2_REG_11_, P3_REG2_REG_12_,
    P3_REG2_REG_13_, P3_REG2_REG_14_, P3_REG2_REG_15_, P3_REG2_REG_16_,
    P3_REG2_REG_17_, P3_REG2_REG_18_, P3_REG2_REG_19_, P3_REG2_REG_20_,
    P3_REG2_REG_21_, P3_REG2_REG_22_, P3_REG2_REG_23_, P3_REG2_REG_24_,
    P3_REG2_REG_25_, P3_REG2_REG_26_, P3_REG2_REG_27_, P3_REG2_REG_28_,
    P3_REG2_REG_29_, P3_REG2_REG_30_, P3_REG2_REG_31_, P3_ADDR_REG_19_,
    P3_ADDR_REG_18_, P3_ADDR_REG_17_, P3_ADDR_REG_16_, P3_ADDR_REG_15_,
    P3_ADDR_REG_14_, P3_ADDR_REG_13_, P3_ADDR_REG_12_, P3_ADDR_REG_11_,
    P3_ADDR_REG_10_, P3_ADDR_REG_9_, P3_ADDR_REG_8_, P3_ADDR_REG_7_,
    P3_ADDR_REG_6_, P3_ADDR_REG_5_, P3_ADDR_REG_4_, P3_ADDR_REG_3_,
    P3_ADDR_REG_2_, P3_ADDR_REG_1_, P3_ADDR_REG_0_, P3_DATAO_REG_0_,
    P3_DATAO_REG_1_, P3_DATAO_REG_2_, P3_DATAO_REG_3_, P3_DATAO_REG_4_,
    P3_DATAO_REG_5_, P3_DATAO_REG_6_, P3_DATAO_REG_7_, P3_DATAO_REG_8_,
    P3_DATAO_REG_9_, P3_DATAO_REG_10_, P3_DATAO_REG_11_, P3_DATAO_REG_12_,
    P3_DATAO_REG_13_, P3_DATAO_REG_14_, P3_DATAO_REG_15_, P3_DATAO_REG_16_,
    P3_DATAO_REG_17_, P3_DATAO_REG_18_, P3_DATAO_REG_19_, P3_DATAO_REG_20_,
    P3_DATAO_REG_21_, P3_DATAO_REG_22_, P3_DATAO_REG_23_, P3_DATAO_REG_24_,
    P3_DATAO_REG_25_, P3_DATAO_REG_26_, P3_DATAO_REG_27_, P3_DATAO_REG_28_,
    P3_DATAO_REG_29_, P3_DATAO_REG_30_, P3_DATAO_REG_31_, P3_B_REG,
    P3_REG3_REG_15_, P3_REG3_REG_26_, P3_REG3_REG_6_, P3_REG3_REG_18_,
    P3_REG3_REG_2_, P3_REG3_REG_11_, P3_REG3_REG_22_, P3_REG3_REG_13_,
    P3_REG3_REG_20_, P3_REG3_REG_0_, P3_REG3_REG_9_, P3_REG3_REG_4_,
    P3_REG3_REG_24_, P3_REG3_REG_17_, P3_REG3_REG_5_, P3_REG3_REG_16_,
    P3_REG3_REG_25_, P3_REG3_REG_12_, P3_REG3_REG_21_, P3_REG3_REG_1_,
    P3_REG3_REG_8_, P3_REG3_REG_28_, P3_REG3_REG_19_, P3_REG3_REG_3_,
    P3_REG3_REG_10_, P3_REG3_REG_23_, P3_REG3_REG_14_, P3_REG3_REG_27_,
    P3_REG3_REG_7_, P3_STATE_REG, P3_RD_REG, P3_WR_REG, Q_0, Q_1, Q_2, Q_3,
    Q_4;
  wire new_P3_R1161_U504, new_P3_R1161_U503, new_P3_R1161_U502, new_U30,
    new_U31, new_U32, new_U33, new_U34, new_U35, new_U36, new_U37, new_U38,
    new_U39, new_U40, new_U41, new_U42, new_U43, new_U44, new_U45, new_U46,
    new_U47, new_U48, new_U49, new_U50, new_U51, new_U52, new_U53, new_U54,
    new_U55, new_U56, new_U57, new_U58, new_U59, new_U60, new_U61, new_U62,
    new_U63, new_U64, new_U65, new_U66, new_U67, new_U68, new_U69, new_U70,
    new_U71, new_U72, new_U73, new_U74, new_U75, new_U76, new_U77, new_U78,
    new_U79, new_U80, new_U81, new_U82, new_U83, new_U84, new_U85, new_U86,
    new_U87, new_U88, new_U89, new_U90, new_U91, new_U92, new_U93, new_U94,
    new_U95, new_U96, new_U97, new_U98, new_U99, new_U100, new_U101,
    new_U102, new_U103, new_U104, new_U105, new_U106, new_U107, new_U108,
    new_U109, new_U110, new_U111, new_U112, new_U113, new_U114, new_U115,
    new_U116, new_U117, new_U118, new_U119, new_U120, new_U121, new_U122,
    new_U123, new_U124, new_U125, new_U126, new_U127, new_U128, new_U129,
    new_U130, new_U131, new_U132, new_U133, new_U134, new_U135, new_U136,
    new_U137, new_U138, new_U139, new_U140, new_U141, new_U142, new_U143,
    new_U144, new_U145, new_U146, new_U147, new_U148, new_U149, new_U150,
    new_U151, new_U152, new_U153, new_U154, new_U155, new_U156, new_U157,
    new_U158, new_U159, new_U160, new_U161, new_U162, new_U163, new_U164,
    new_U165, new_U166, new_U167, new_U168, new_U169, new_U170, new_U171,
    new_U172, new_U173, new_U174, new_U175, new_U176, new_U177, new_U178,
    new_U179, new_U180, new_U181, new_U182, new_U183, new_U184, new_U185,
    new_U186, new_U187, new_U188, new_U189, new_U190, new_U191, new_U192,
    new_U193, new_U194, new_U195, new_U196, new_U197, new_U198, new_U199,
    new_U200, new_U201, new_U202, new_U203, new_U204, new_U205, new_U206,
    new_U207, new_U208, new_U209, new_U210, new_U211, new_U212, new_U213,
    new_U214, new_U215, new_U216, new_U217, new_U218, new_U219, new_U220,
    new_U221, new_U222, new_U223, new_U224, new_U225, new_U226, new_U227,
    new_U228, new_U229, new_U230, new_U231, new_U232, new_U233, new_U234,
    new_U235, new_U236, new_U237, new_U238, new_U239, new_U240, new_U241,
    new_U242, new_U243, new_U244, new_U245, new_U246, new_U247, new_U248,
    new_U249, new_U250, new_U251, new_U252, new_U253, new_U254, new_U255,
    new_U256, new_U257, new_U258, new_U259, new_U260, new_U261, new_U262,
    new_U263, new_U264, new_U265, new_U266, new_U267, new_U268, new_U269,
    new_U270, new_U271, new_U272, new_U273, new_U274, new_U275, new_U276,
    new_U277, new_U278, new_U279, new_U280, new_U281, new_U282, new_U283,
    new_U284, new_U285, new_U286, new_U287, new_U288, new_U289, new_U290,
    new_U291, new_U292, new_U293, new_U294, new_U295, new_U296, new_U297,
    new_U298, new_U299, new_U300, new_U301, new_U302, new_U303, new_U304,
    new_U305, new_U306, new_U307, new_U308, new_U309, new_U310, new_U311,
    new_U312, new_U313, new_U314, new_U315, new_U316, new_U317, new_U318,
    new_U319, new_U320, new_U321, new_U322, new_U323, new_U324, new_U325,
    new_U326, new_U327, new_U328, new_U329, new_U330, new_U331, new_U332,
    new_U333, new_U334, new_U335, new_U336, new_U337, new_U338, new_U339,
    new_U340, new_U341, new_U342, new_U343, new_U344, new_U345, new_U346,
    new_U347, new_U348, new_U349, new_U350, new_U351, new_U352, new_U353,
    new_U354, new_U355, new_U356, new_U357, new_U358, new_U359, new_U360,
    new_U361, new_U362, new_U363, new_U364, new_U365, new_U366, new_U367,
    new_U368, new_U369, new_U370, new_U371, new_U372, new_U373, new_U374,
    new_U375, new_U376, new_U377, new_U378, new_U379, new_U380, new_U381,
    new_U382, new_U383, new_U384, new_U385, new_U386, new_U387, new_U388,
    new_U389, new_U390, new_U391, new_U392, new_U393, new_U394, new_U395,
    new_U396, new_U397, new_U398, new_U399, new_U400, new_U401, new_U402,
    new_U403, new_U404, new_U405, new_U406, new_U407, new_U408, new_U409,
    new_U410, new_U411, new_U412, new_U413, new_U414, new_U415, new_U416,
    new_U417, new_U418, new_U419, new_U420, new_U421, new_U422, new_U423,
    new_U424, new_U425, new_U426, new_U427, new_P3_R1161_U501,
    new_P3_R1161_U500, new_P3_R1161_U499, new_P3_R1161_U498,
    new_P3_R1161_U497, new_P3_R1161_U496, new_P3_R1161_U495,
    new_P3_R1161_U494, new_P3_R1161_U493, new_P3_R1161_U492,
    new_P3_R1161_U491, new_P3_R1161_U490, new_P1_U3014, new_P1_U3015,
    new_P1_U3016, new_P1_U3017, new_P1_U3018, new_P1_U3019, new_P1_U3020,
    new_P1_U3021, new_P1_U3022, new_P1_U3023, new_P1_U3024, new_P1_U3025,
    new_P1_U3026, new_P1_U3027, new_P1_U3028, new_P1_U3029, new_P1_U3030,
    new_P1_U3031, new_P1_U3032, new_P1_U3033, new_P1_U3034, new_P1_U3035,
    new_P1_U3036, new_P1_U3037, new_P1_U3038, new_P1_U3039, new_P1_U3040,
    new_P1_U3041, new_P1_U3042, new_P1_U3043, new_P1_U3044, new_P1_U3045,
    new_P1_U3046, new_P1_U3047, new_P1_U3048, new_P1_U3049, new_P1_U3050,
    new_P1_U3051, new_P1_U3052, new_P1_U3053, new_P1_U3054, new_P1_U3055,
    new_P1_U3056, new_P1_U3057, new_P1_U3058, new_P1_U3059, new_P1_U3060,
    new_P1_U3061, new_P1_U3062, new_P1_U3063, new_P1_U3064, new_P1_U3065,
    new_P1_U3066, new_P1_U3067, new_P1_U3068, new_P1_U3069, new_P1_U3070,
    new_P1_U3071, new_P1_U3072, new_P1_U3073, new_P1_U3074, new_P1_U3075,
    new_P1_U3076, new_P1_U3077, new_P1_U3078, new_P1_U3079, new_P1_U3080,
    new_P1_U3081, new_P1_U3082, new_P1_U3083, new_P1_U3084, new_P1_U3087,
    new_P1_U3088, new_P1_U3089, new_P1_U3090, new_P1_U3091, new_P1_U3092,
    new_P1_U3093, new_P1_U3094, new_P1_U3095, new_P1_U3096, new_P1_U3097,
    new_P1_U3098, new_P1_U3099, new_P1_U3100, new_P1_U3101, new_P1_U3102,
    new_P1_U3103, new_P1_U3104, new_P1_U3105, new_P1_U3106, new_P1_U3107,
    new_P1_U3108, new_P1_U3109, new_P1_U3110, new_P1_U3111, new_P1_U3112,
    new_P1_U3113, new_P1_U3114, new_P1_U3115, new_P1_U3116, new_P1_U3117,
    new_P1_U3118, new_P1_U3119, new_P1_U3120, new_P1_U3121, new_P1_U3122,
    new_P1_U3123, new_P1_U3124, new_P1_U3125, new_P1_U3126, new_P1_U3127,
    new_P1_U3128, new_P1_U3129, new_P1_U3130, new_P1_U3131, new_P1_U3132,
    new_P1_U3133, new_P1_U3134, new_P1_U3135, new_P1_U3136, new_P1_U3137,
    new_P1_U3138, new_P1_U3139, new_P1_U3140, new_P1_U3141, new_P1_U3142,
    new_P1_U3143, new_P1_U3144, new_P1_U3145, new_P1_U3146, new_P1_U3147,
    new_P1_U3148, new_P1_U3149, new_P1_U3150, new_P1_U3151, new_P1_U3152,
    new_P1_U3153, new_P1_U3154, new_P1_U3155, new_P1_U3156, new_P1_U3157,
    new_P1_U3158, new_P1_U3159, new_P1_U3160, new_P1_U3161, new_P1_U3162,
    new_P1_U3163, new_P1_U3164, new_P1_U3165, new_P1_U3166, new_P1_U3167,
    new_P1_U3168, new_P1_U3169, new_P1_U3170, new_P1_U3171, new_P1_U3172,
    new_P1_U3173, new_P1_U3174, new_P1_U3175, new_P1_U3176, new_P1_U3177,
    new_P1_U3178, new_P1_U3179, new_P1_U3180, new_P1_U3181, new_P1_U3182,
    new_P1_U3183, new_P1_U3184, new_P1_U3185, new_P1_U3186, new_P1_U3187,
    new_P1_U3188, new_P1_U3189, new_P1_U3190, new_P1_U3191, new_P1_U3192,
    new_P1_U3193, new_P1_U3194, new_P1_U3195, new_P1_U3196, new_P1_U3197,
    new_P1_U3198, new_P1_U3199, new_P1_U3200, new_P1_U3201, new_P1_U3202,
    new_P1_U3203, new_P1_U3204, new_P1_U3205, new_P1_U3206, new_P1_U3207,
    new_P1_U3208, new_P1_U3209, new_P1_U3210, new_P1_U3211, new_P1_U3212,
    new_P1_U3355, new_P1_U3357, new_P1_U3358, new_P1_U3359, new_P1_U3360,
    new_P1_U3361, new_P1_U3362, new_P1_U3363, new_P1_U3364, new_P1_U3365,
    new_P1_U3366, new_P1_U3367, new_P1_U3368, new_P1_U3369, new_P1_U3370,
    new_P1_U3371, new_P1_U3372, new_P1_U3373, new_P1_U3374, new_P1_U3375,
    new_P1_U3376, new_P1_U3377, new_P1_U3378, new_P1_U3379, new_P1_U3380,
    new_P1_U3381, new_P1_U3382, new_P1_U3383, new_P1_U3384, new_P1_U3385,
    new_P1_U3386, new_P1_U3387, new_P1_U3388, new_P1_U3389, new_P1_U3390,
    new_P1_U3391, new_P1_U3392, new_P1_U3393, new_P1_U3394, new_P1_U3395,
    new_P1_U3396, new_P1_U3397, new_P1_U3398, new_P1_U3399, new_P1_U3400,
    new_P1_U3401, new_P1_U3402, new_P1_U3403, new_P1_U3404, new_P1_U3405,
    new_P1_U3406, new_P1_U3407, new_P1_U3408, new_P1_U3409, new_P1_U3410,
    new_P1_U3411, new_P1_U3412, new_P1_U3413, new_P1_U3414, new_P1_U3415,
    new_P1_U3416, new_P1_U3417, new_P1_U3418, new_P1_U3419, new_P1_U3420,
    new_P1_U3421, new_P1_U3422, new_P1_U3423, new_P1_U3424, new_P1_U3425,
    new_P1_U3426, new_P1_U3427, new_P1_U3428, new_P1_U3429, new_P1_U3430,
    new_P1_U3431, new_P1_U3432, new_P1_U3433, new_P1_U3434, new_P1_U3435,
    new_P1_U3436, new_P1_U3437, new_P1_U3438, new_P1_U3439, new_P1_U3440,
    new_P1_U3441, new_P1_U3442, new_P1_U3443, new_P1_U3444, new_P1_U3447,
    new_P1_U3448, new_P1_U3449, new_P1_U3450, new_P1_U3451, new_P1_U3452,
    new_P1_U3453, new_P1_U3454, new_P1_U3455, new_P1_U3456, new_P1_U3457,
    new_P1_U3458, new_P1_U3460, new_P1_U3461, new_P1_U3463, new_P1_U3464,
    new_P1_U3466, new_P1_U3467, new_P1_U3469, new_P1_U3470, new_P1_U3472,
    new_P1_U3473, new_P1_U3475, new_P1_U3476, new_P1_U3478, new_P1_U3479,
    new_P1_U3481, new_P1_U3482, new_P1_U3484, new_P1_U3485, new_P1_U3487,
    new_P1_U3488, new_P1_U3490, new_P1_U3491, new_P1_U3493, new_P1_U3494,
    new_P1_U3496, new_P1_U3497, new_P1_U3499, new_P1_U3500, new_P1_U3502,
    new_P1_U3503, new_P1_U3505, new_P1_U3506, new_P1_U3508, new_P1_U3509,
    new_P1_U3511, new_P1_U3512, new_P1_U3514, new_P1_U3592, new_P1_U3593,
    new_P1_U3594, new_P1_U3595, new_P1_U3596, new_P1_U3597, new_P1_U3598,
    new_P1_U3599, new_P1_U3600, new_P1_U3601, new_P1_U3602, new_P1_U3603,
    new_P1_U3604, new_P1_U3605, new_P1_U3606, new_P1_U3607, new_P1_U3608,
    new_P1_U3609, new_P1_U3610, new_P1_U3611, new_P1_U3612, new_P1_U3613,
    new_P1_U3614, new_P1_U3615, new_P1_U3616, new_P1_U3617, new_P1_U3618,
    new_P1_U3619, new_P1_U3620, new_P1_U3621, new_P1_U3622, new_P1_U3623,
    new_P1_U3624, new_P1_U3625, new_P1_U3626, new_P1_U3627, new_P1_U3628,
    new_P1_U3629, new_P1_U3630, new_P1_U3631, new_P1_U3632, new_P1_U3633,
    new_P1_U3634, new_P1_U3635, new_P1_U3636, new_P1_U3637, new_P1_U3638,
    new_P1_U3639, new_P1_U3640, new_P1_U3641, new_P1_U3642, new_P1_U3643,
    new_P1_U3644, new_P1_U3645, new_P1_U3646, new_P1_U3647, new_P1_U3648,
    new_P1_U3649, new_P1_U3650, new_P1_U3651, new_P1_U3652, new_P1_U3653,
    new_P1_U3654, new_P1_U3655, new_P1_U3656, new_P1_U3657, new_P1_U3658,
    new_P1_U3659, new_P1_U3660, new_P1_U3661, new_P1_U3662, new_P1_U3663,
    new_P1_U3664, new_P1_U3665, new_P1_U3666, new_P1_U3667, new_P1_U3668,
    new_P1_U3669, new_P1_U3670, new_P1_U3671, new_P1_U3672, new_P1_U3673,
    new_P1_U3674, new_P1_U3675, new_P1_U3676, new_P1_U3677, new_P1_U3678,
    new_P1_U3679, new_P1_U3680, new_P1_U3681, new_P1_U3682, new_P1_U3683,
    new_P1_U3684, new_P1_U3685, new_P1_U3686, new_P1_U3687, new_P1_U3688,
    new_P1_U3689, new_P1_U3690, new_P1_U3691, new_P1_U3692, new_P1_U3693,
    new_P1_U3694, new_P1_U3695, new_P1_U3696, new_P1_U3697, new_P1_U3698,
    new_P1_U3699, new_P1_U3700, new_P1_U3701, new_P1_U3702, new_P1_U3703,
    new_P1_U3704, new_P1_U3705, new_P1_U3706, new_P1_U3707, new_P1_U3708,
    new_P1_U3709, new_P1_U3710, new_P1_U3711, new_P1_U3712, new_P1_U3713,
    new_P1_U3714, new_P1_U3715, new_P1_U3716, new_P1_U3717, new_P1_U3718,
    new_P1_U3719, new_P1_U3720, new_P1_U3721, new_P1_U3722, new_P1_U3723,
    new_P1_U3724, new_P1_U3725, new_P1_U3726, new_P1_U3727, new_P1_U3728,
    new_P1_U3729, new_P1_U3730, new_P1_U3731, new_P1_U3732, new_P1_U3733,
    new_P1_U3734, new_P1_U3735, new_P1_U3736, new_P1_U3737, new_P1_U3738,
    new_P1_U3739, new_P1_U3740, new_P1_U3741, new_P1_U3742, new_P1_U3743,
    new_P1_U3744, new_P1_U3745, new_P1_U3746, new_P1_U3747, new_P1_U3748,
    new_P1_U3749, new_P1_U3750, new_P1_U3751, new_P1_U3752, new_P1_U3753,
    new_P1_U3754, new_P1_U3755, new_P1_U3756, new_P1_U3757, new_P1_U3758,
    new_P1_U3759, new_P1_U3760, new_P1_U3761, new_P1_U3762, new_P1_U3763,
    new_P1_U3764, new_P1_U3765, new_P1_U3766, new_P1_U3767, new_P1_U3768,
    new_P1_U3769, new_P1_U3770, new_P1_U3771, new_P1_U3772, new_P1_U3773,
    new_P1_U3774, new_P1_U3775, new_P1_U3776, new_P1_U3777, new_P1_U3778,
    new_P1_U3779, new_P1_U3780, new_P1_U3781, new_P1_U3782, new_P1_U3783,
    new_P1_U3784, new_P1_U3785, new_P1_U3786, new_P1_U3787, new_P1_U3788,
    new_P1_U3789, new_P1_U3790, new_P1_U3791, new_P1_U3792, new_P1_U3793,
    new_P1_U3794, new_P1_U3795, new_P1_U3796, new_P1_U3797, new_P1_U3798,
    new_P1_U3799, new_P1_U3800, new_P1_U3801, new_P1_U3802, new_P1_U3803,
    new_P1_U3804, new_P1_U3805, new_P1_U3806, new_P1_U3807, new_P1_U3808,
    new_P1_U3809, new_P1_U3810, new_P1_U3811, new_P1_U3812, new_P1_U3813,
    new_P1_U3814, new_P1_U3815, new_P1_U3816, new_P1_U3817, new_P1_U3818,
    new_P1_U3819, new_P1_U3820, new_P1_U3821, new_P1_U3822, new_P1_U3823,
    new_P1_U3824, new_P1_U3825, new_P1_U3826, new_P1_U3827, new_P1_U3828,
    new_P1_U3829, new_P1_U3830, new_P1_U3831, new_P1_U3832, new_P1_U3833,
    new_P1_U3834, new_P1_U3835, new_P1_U3836, new_P1_U3837, new_P1_U3838,
    new_P1_U3839, new_P1_U3840, new_P1_U3841, new_P1_U3842, new_P1_U3843,
    new_P1_U3844, new_P1_U3845, new_P1_U3846, new_P1_U3847, new_P1_U3848,
    new_P1_U3849, new_P1_U3850, new_P1_U3851, new_P1_U3852, new_P1_U3853,
    new_P1_U3854, new_P1_U3855, new_P1_U3856, new_P1_U3857, new_P1_U3858,
    new_P1_U3859, new_P1_U3860, new_P1_U3861, new_P1_U3862, new_P1_U3863,
    new_P1_U3864, new_P1_U3865, new_P1_U3866, new_P1_U3867, new_P1_U3868,
    new_P1_U3869, new_P1_U3870, new_P1_U3871, new_P1_U3872, new_P1_U3873,
    new_P1_U3874, new_P1_U3875, new_P1_U3876, new_P1_U3877, new_P1_U3878,
    new_P1_U3879, new_P1_U3880, new_P1_U3881, new_P1_U3882, new_P1_U3883,
    new_P1_U3884, new_P1_U3885, new_P1_U3886, new_P1_U3887, new_P1_U3888,
    new_P1_U3889, new_P1_U3890, new_P1_U3891, new_P1_U3892, new_P1_U3893,
    new_P1_U3894, new_P1_U3895, new_P1_U3896, new_P1_U3897, new_P1_U3898,
    new_P1_U3899, new_P1_U3900, new_P1_U3901, new_P1_U3902, new_P1_U3903,
    new_P1_U3904, new_P1_U3905, new_P1_U3906, new_P1_U3907, new_P1_U3908,
    new_P1_U3909, new_P1_U3910, new_P1_U3911, new_P1_U3912, new_P1_U3913,
    new_P1_U3914, new_P1_U3915, new_P1_U3916, new_P1_U3917, new_P1_U3918,
    new_P1_U3919, new_P1_U3920, new_P1_U3921, new_P1_U3922, new_P1_U3923,
    new_P1_U3924, new_P1_U3925, new_P1_U3926, new_P1_U3927, new_P1_U3928,
    new_P1_U3929, new_P1_U3930, new_P1_U3931, new_P1_U3932, new_P1_U3933,
    new_P1_U3934, new_P1_U3935, new_P1_U3936, new_P1_U3937, new_P1_U3938,
    new_P1_U3939, new_P1_U3940, new_P1_U3941, new_P1_U3942, new_P1_U3943,
    new_P1_U3944, new_P1_U3945, new_P1_U3946, new_P1_U3947, new_P1_U3948,
    new_P1_U3949, new_P1_U3950, new_P1_U3951, new_P1_U3952, new_P1_U3953,
    new_P1_U3954, new_P1_U3955, new_P1_U3956, new_P1_U3957, new_P1_U3958,
    new_P1_U3959, new_P1_U3960, new_P1_U3961, new_P1_U3962, new_P1_U3963,
    new_P1_U3964, new_P1_U3965, new_P1_U3966, new_P1_U3967, new_P1_U3968,
    new_P1_U3969, new_P1_U3970, new_P1_U3971, new_P1_U3972, new_P1_U3973,
    new_P1_U3974, new_P1_U3975, new_P1_U3976, new_P1_U3977, new_P1_U3978,
    new_P1_U3979, new_P1_U3980, new_P1_U3981, new_P1_U3982, new_P1_U3983,
    new_P1_U3984, new_P1_U3985, new_P1_U3986, new_P1_U3987, new_P1_U3988,
    new_P1_U3989, new_P1_U3990, new_P1_U3991, new_P1_U3992, new_P1_U3993,
    new_P1_U3994, new_P1_U3995, new_P1_U3996, new_P1_U3997, new_P1_U3998,
    new_P1_U3999, new_P1_U4000, new_P1_U4001, new_P1_U4002, new_P1_U4003,
    new_P1_U4004, new_P1_U4005, new_P1_U4006, new_P1_U4007, new_P1_U4008,
    new_P1_U4009, new_P1_U4010, new_P1_U4011, new_P1_U4012, new_P1_U4013,
    new_P1_U4014, new_P1_U4015, new_P1_U4017, new_P1_U4018, new_P1_U4019,
    new_P1_U4020, new_P1_U4021, new_P1_U4022, new_P1_U4023, new_P1_U4024,
    new_P1_U4025, new_P1_U4026, new_P1_U4027, new_P1_U4028, new_P1_U4029,
    new_P1_U4030, new_P1_U4031, new_P1_U4032, new_P1_U4033, new_P1_U4034,
    new_P1_U4035, new_P1_U4036, new_P1_U4037, new_P1_U4038, new_P1_U4039,
    new_P1_U4040, new_P1_U4041, new_P1_U4042, new_P1_U4043, new_P1_U4044,
    new_P1_U4045, new_P1_U4046, new_P1_U4047, new_P1_U4048, new_P1_U4049,
    new_P1_U4050, new_P1_U4051, new_P1_U4052, new_P1_U4053, new_P1_U4054,
    new_P1_U4055, new_P1_U4056, new_P1_U4057, new_P1_U4058, new_P1_U4059,
    new_P1_U4060, new_P1_U4061, new_P1_U4062, new_P1_U4063, new_P1_U4064,
    new_P1_U4065, new_P1_U4066, new_P1_U4067, new_P1_U4068, new_P1_U4069,
    new_P1_U4070, new_P1_U4071, new_P1_U4072, new_P1_U4073, new_P1_U4074,
    new_P1_U4075, new_P1_U4076, new_P1_U4077, new_P1_U4078, new_P1_U4079,
    new_P1_U4080, new_P1_U4081, new_P1_U4082, new_P1_U4083, new_P1_U4084,
    new_P1_U4085, new_P1_U4086, new_P1_U4087, new_P1_U4088, new_P1_U4089,
    new_P1_U4090, new_P1_U4091, new_P1_U4092, new_P1_U4093, new_P1_U4094,
    new_P1_U4095, new_P1_U4096, new_P1_U4097, new_P1_U4098, new_P1_U4099,
    new_P1_U4100, new_P1_U4101, new_P1_U4102, new_P1_U4103, new_P1_U4104,
    new_P1_U4105, new_P1_U4106, new_P1_U4107, new_P1_U4108, new_P1_U4109,
    new_P1_U4110, new_P1_U4111, new_P1_U4112, new_P1_U4113, new_P1_U4114,
    new_P1_U4115, new_P1_U4116, new_P1_U4117, new_P1_U4118, new_P1_U4119,
    new_P1_U4120, new_P1_U4121, new_P1_U4122, new_P1_U4123, new_P1_U4124,
    new_P1_U4125, new_P1_U4126, new_P1_U4127, new_P1_U4128, new_P1_U4129,
    new_P1_U4130, new_P1_U4131, new_P1_U4132, new_P1_U4133, new_P1_U4134,
    new_P1_U4135, new_P1_U4136, new_P1_U4137, new_P1_U4138, new_P1_U4139,
    new_P1_U4140, new_P1_U4141, new_P1_U4142, new_P1_U4143, new_P1_U4144,
    new_P1_U4145, new_P1_U4146, new_P1_U4147, new_P1_U4148, new_P1_U4149,
    new_P1_U4150, new_P1_U4151, new_P1_U4152, new_P1_U4153, new_P1_U4154,
    new_P1_U4155, new_P1_U4156, new_P1_U4157, new_P1_U4158, new_P1_U4159,
    new_P1_U4160, new_P1_U4161, new_P1_U4162, new_P1_U4163, new_P1_U4164,
    new_P1_U4165, new_P1_U4166, new_P1_U4167, new_P1_U4168, new_P1_U4169,
    new_P1_U4170, new_P1_U4171, new_P1_U4172, new_P1_U4173, new_P1_U4174,
    new_P1_U4175, new_P1_U4176, new_P1_U4177, new_P1_U4178, new_P1_U4179,
    new_P1_U4180, new_P1_U4181, new_P1_U4182, new_P1_U4183, new_P1_U4184,
    new_P1_U4185, new_P1_U4186, new_P1_U4187, new_P1_U4188, new_P1_U4189,
    new_P1_U4190, new_P1_U4191, new_P1_U4192, new_P1_U4193, new_P1_U4194,
    new_P1_U4195, new_P1_U4196, new_P1_U4197, new_P1_U4198, new_P1_U4199,
    new_P1_U4200, new_P1_U4201, new_P1_U4202, new_P1_U4203, new_P1_U4204,
    new_P1_U4205, new_P1_U4206, new_P1_U4207, new_P1_U4208, new_P1_U4209,
    new_P1_U4210, new_P1_U4211, new_P1_U4212, new_P1_U4213, new_P1_U4214,
    new_P1_U4215, new_P1_U4216, new_P1_U4217, new_P1_U4218, new_P1_U4219,
    new_P1_U4220, new_P1_U4221, new_P1_U4222, new_P1_U4223, new_P1_U4224,
    new_P1_U4225, new_P1_U4226, new_P1_U4227, new_P1_U4228, new_P1_U4229,
    new_P1_U4230, new_P1_U4231, new_P1_U4232, new_P1_U4233, new_P1_U4234,
    new_P1_U4235, new_P1_U4236, new_P1_U4237, new_P1_U4238, new_P1_U4239,
    new_P1_U4240, new_P1_U4241, new_P1_U4242, new_P1_U4243, new_P1_U4244,
    new_P1_U4245, new_P1_U4246, new_P1_U4247, new_P1_U4248, new_P1_U4249,
    new_P1_U4250, new_P1_U4251, new_P1_U4252, new_P1_U4253, new_P1_U4254,
    new_P1_U4255, new_P1_U4256, new_P1_U4257, new_P1_U4258, new_P1_U4259,
    new_P1_U4260, new_P1_U4261, new_P1_U4262, new_P1_U4263, new_P1_U4264,
    new_P1_U4265, new_P1_U4266, new_P1_U4267, new_P1_U4268, new_P1_U4269,
    new_P1_U4270, new_P1_U4271, new_P1_U4272, new_P1_U4273, new_P1_U4274,
    new_P1_U4275, new_P1_U4276, new_P1_U4277, new_P1_U4278, new_P1_U4279,
    new_P1_U4280, new_P1_U4281, new_P1_U4282, new_P1_U4283, new_P1_U4284,
    new_P1_U4285, new_P1_U4286, new_P1_U4287, new_P1_U4288, new_P1_U4289,
    new_P1_U4290, new_P1_U4291, new_P1_U4292, new_P1_U4293, new_P1_U4294,
    new_P1_U4295, new_P1_U4296, new_P1_U4297, new_P1_U4298, new_P1_U4299,
    new_P1_U4300, new_P1_U4301, new_P1_U4302, new_P1_U4303, new_P1_U4304,
    new_P1_U4305, new_P1_U4306, new_P1_U4307, new_P1_U4308, new_P1_U4309,
    new_P1_U4310, new_P1_U4311, new_P1_U4312, new_P1_U4313, new_P1_U4314,
    new_P1_U4315, new_P1_U4316, new_P1_U4317, new_P1_U4318, new_P1_U4319,
    new_P1_U4320, new_P1_U4321, new_P1_U4322, new_P1_U4323, new_P1_U4324,
    new_P1_U4325, new_P1_U4326, new_P1_U4327, new_P1_U4328, new_P1_U4329,
    new_P1_U4330, new_P1_U4331, new_P1_U4332, new_P1_U4333, new_P1_U4334,
    new_P1_U4335, new_P1_U4336, new_P1_U4337, new_P1_U4338, new_P1_U4339,
    new_P1_U4340, new_P1_U4341, new_P1_U4342, new_P1_U4343, new_P1_U4344,
    new_P1_U4345, new_P1_U4346, new_P1_U4347, new_P1_U4348, new_P1_U4349,
    new_P1_U4350, new_P1_U4351, new_P1_U4352, new_P1_U4353, new_P1_U4354,
    new_P1_U4355, new_P1_U4356, new_P1_U4357, new_P1_U4358, new_P1_U4359,
    new_P1_U4360, new_P1_U4361, new_P1_U4362, new_P1_U4363, new_P1_U4364,
    new_P1_U4365, new_P1_U4366, new_P1_U4367, new_P1_U4368, new_P1_U4369,
    new_P1_U4370, new_P1_U4371, new_P1_U4372, new_P1_U4373, new_P1_U4374,
    new_P1_U4375, new_P1_U4376, new_P1_U4377, new_P1_U4378, new_P1_U4379,
    new_P1_U4380, new_P1_U4381, new_P1_U4382, new_P1_U4383, new_P1_U4384,
    new_P1_U4385, new_P1_U4386, new_P1_U4387, new_P1_U4388, new_P1_U4389,
    new_P1_U4390, new_P1_U4391, new_P1_U4392, new_P1_U4393, new_P1_U4394,
    new_P1_U4395, new_P1_U4396, new_P1_U4397, new_P1_U4398, new_P1_U4399,
    new_P1_U4400, new_P1_U4401, new_P1_U4402, new_P1_U4403, new_P1_U4404,
    new_P1_U4405, new_P1_U4406, new_P1_U4407, new_P1_U4408, new_P1_U4409,
    new_P1_U4410, new_P1_U4411, new_P1_U4412, new_P1_U4413, new_P1_U4414,
    new_P1_U4415, new_P1_U4416, new_P1_U4417, new_P1_U4418, new_P1_U4419,
    new_P1_U4420, new_P1_U4421, new_P1_U4422, new_P1_U4423, new_P1_U4424,
    new_P1_U4425, new_P1_U4426, new_P1_U4427, new_P1_U4428, new_P1_U4429,
    new_P1_U4430, new_P1_U4431, new_P1_U4432, new_P1_U4433, new_P1_U4434,
    new_P1_U4435, new_P1_U4436, new_P1_U4437, new_P1_U4438, new_P1_U4439,
    new_P1_U4440, new_P1_U4441, new_P1_U4442, new_P1_U4443, new_P1_U4444,
    new_P1_U4445, new_P1_U4446, new_P1_U4447, new_P1_U4448, new_P1_U4449,
    new_P1_U4450, new_P1_U4451, new_P1_U4452, new_P1_U4453, new_P1_U4454,
    new_P1_U4455, new_P1_U4456, new_P1_U4457, new_P1_U4458, new_P1_U4459,
    new_P1_U4460, new_P1_U4461, new_P1_U4462, new_P1_U4463, new_P1_U4464,
    new_P1_U4465, new_P1_U4466, new_P1_U4467, new_P1_U4468, new_P1_U4469,
    new_P1_U4470, new_P1_U4471, new_P1_U4472, new_P1_U4473, new_P1_U4474,
    new_P1_U4475, new_P1_U4476, new_P1_U4477, new_P1_U4478, new_P1_U4479,
    new_P1_U4480, new_P1_U4481, new_P1_U4482, new_P1_U4483, new_P1_U4484,
    new_P1_U4485, new_P1_U4486, new_P1_U4487, new_P1_U4488, new_P1_U4489,
    new_P1_U4490, new_P1_U4491, new_P1_U4492, new_P1_U4493, new_P1_U4494,
    new_P1_U4495, new_P1_U4496, new_P1_U4497, new_P1_U4498, new_P1_U4499,
    new_P1_U4500, new_P1_U4501, new_P1_U4502, new_P1_U4503, new_P1_U4504,
    new_P1_U4505, new_P1_U4506, new_P1_U4507, new_P1_U4508, new_P1_U4509,
    new_P1_U4510, new_P1_U4511, new_P1_U4512, new_P1_U4513, new_P1_U4514,
    new_P1_U4515, new_P1_U4516, new_P1_U4517, new_P1_U4518, new_P1_U4519,
    new_P1_U4520, new_P1_U4521, new_P1_U4522, new_P1_U4523, new_P1_U4524,
    new_P1_U4525, new_P1_U4526, new_P1_U4527, new_P1_U4528, new_P1_U4529,
    new_P1_U4530, new_P1_U4531, new_P1_U4532, new_P1_U4533, new_P1_U4534,
    new_P1_U4535, new_P1_U4536, new_P1_U4537, new_P1_U4538, new_P1_U4539,
    new_P1_U4540, new_P1_U4541, new_P1_U4542, new_P1_U4543, new_P1_U4544,
    new_P1_U4545, new_P1_U4546, new_P1_U4547, new_P1_U4548, new_P1_U4549,
    new_P1_U4550, new_P1_U4551, new_P1_U4552, new_P1_U4553, new_P1_U4554,
    new_P1_U4555, new_P1_U4556, new_P1_U4557, new_P1_U4558, new_P1_U4559,
    new_P1_U4560, new_P1_U4561, new_P1_U4562, new_P1_U4563, new_P1_U4564,
    new_P1_U4565, new_P1_U4566, new_P1_U4567, new_P1_U4568, new_P1_U4569,
    new_P1_U4570, new_P1_U4571, new_P1_U4572, new_P1_U4573, new_P1_U4574,
    new_P1_U4575, new_P1_U4576, new_P1_U4577, new_P1_U4578, new_P1_U4579,
    new_P1_U4580, new_P1_U4581, new_P1_U4582, new_P1_U4583, new_P1_U4584,
    new_P1_U4585, new_P1_U4586, new_P1_U4587, new_P1_U4588, new_P1_U4589,
    new_P1_U4590, new_P1_U4591, new_P1_U4592, new_P1_U4593, new_P1_U4594,
    new_P1_U4595, new_P1_U4596, new_P1_U4597, new_P1_U4598, new_P1_U4599,
    new_P1_U4600, new_P1_U4601, new_P1_U4602, new_P1_U4603, new_P1_U4604,
    new_P1_U4605, new_P1_U4606, new_P1_U4607, new_P1_U4608, new_P1_U4609,
    new_P1_U4610, new_P1_U4611, new_P1_U4612, new_P1_U4613, new_P1_U4614,
    new_P1_U4615, new_P1_U4616, new_P1_U4617, new_P1_U4618, new_P1_U4619,
    new_P1_U4620, new_P1_U4621, new_P1_U4622, new_P1_U4623, new_P1_U4624,
    new_P1_U4625, new_P1_U4626, new_P1_U4627, new_P1_U4628, new_P1_U4629,
    new_P1_U4630, new_P1_U4631, new_P1_U4632, new_P1_U4633, new_P1_U4634,
    new_P1_U4635, new_P1_U4636, new_P1_U4637, new_P1_U4638, new_P1_U4639,
    new_P1_U4640, new_P1_U4641, new_P1_U4642, new_P1_U4643, new_P1_U4644,
    new_P1_U4645, new_P1_U4646, new_P1_U4647, new_P1_U4648, new_P1_U4649,
    new_P1_U4650, new_P1_U4651, new_P1_U4652, new_P1_U4653, new_P1_U4654,
    new_P1_U4655, new_P1_U4656, new_P1_U4657, new_P1_U4658, new_P1_U4659,
    new_P1_U4660, new_P1_U4661, new_P1_U4662, new_P1_U4663, new_P1_U4664,
    new_P1_U4665, new_P1_U4666, new_P1_U4667, new_P1_U4668, new_P1_U4669,
    new_P1_U4670, new_P1_U4671, new_P1_U4672, new_P1_U4673, new_P1_U4674,
    new_P1_U4675, new_P1_U4676, new_P1_U4677, new_P1_U4678, new_P1_U4679,
    new_P1_U4680, new_P1_U4681, new_P1_U4682, new_P1_U4683, new_P1_U4684,
    new_P1_U4685, new_P1_U4686, new_P1_U4687, new_P1_U4688, new_P1_U4689,
    new_P1_U4690, new_P1_U4691, new_P1_U4692, new_P1_U4693, new_P1_U4694,
    new_P1_U4695, new_P1_U4696, new_P1_U4697, new_P1_U4698, new_P1_U4699,
    new_P1_U4700, new_P1_U4701, new_P1_U4702, new_P1_U4703, new_P1_U4704,
    new_P1_U4705, new_P1_U4706, new_P1_U4707, new_P1_U4708, new_P1_U4709,
    new_P1_U4710, new_P1_U4711, new_P1_U4712, new_P1_U4713, new_P1_U4714,
    new_P1_U4715, new_P1_U4716, new_P1_U4717, new_P1_U4718, new_P1_U4719,
    new_P1_U4720, new_P1_U4721, new_P1_U4722, new_P1_U4723, new_P1_U4724,
    new_P1_U4725, new_P1_U4726, new_P1_U4727, new_P1_U4728, new_P1_U4729,
    new_P1_U4730, new_P1_U4731, new_P1_U4732, new_P1_U4733, new_P1_U4734,
    new_P1_U4735, new_P1_U4736, new_P1_U4737, new_P1_U4738, new_P1_U4739,
    new_P1_U4740, new_P1_U4741, new_P1_U4742, new_P1_U4743, new_P1_U4744,
    new_P1_U4745, new_P1_U4746, new_P1_U4747, new_P1_U4748, new_P1_U4749,
    new_P1_U4750, new_P1_U4751, new_P1_U4752, new_P1_U4753, new_P1_U4754,
    new_P1_U4755, new_P1_U4756, new_P1_U4757, new_P1_U4758, new_P1_U4759,
    new_P1_U4760, new_P1_U4761, new_P1_U4762, new_P1_U4763, new_P1_U4764,
    new_P1_U4765, new_P1_U4766, new_P1_U4767, new_P1_U4768, new_P1_U4769,
    new_P1_U4770, new_P1_U4771, new_P1_U4772, new_P1_U4773, new_P1_U4774,
    new_P1_U4775, new_P1_U4776, new_P1_U4777, new_P1_U4778, new_P1_U4779,
    new_P1_U4780, new_P1_U4781, new_P1_U4782, new_P1_U4783, new_P1_U4784,
    new_P1_U4785, new_P1_U4786, new_P1_U4787, new_P1_U4788, new_P1_U4789,
    new_P1_U4790, new_P1_U4791, new_P1_U4792, new_P1_U4793, new_P1_U4794,
    new_P1_U4795, new_P1_U4796, new_P1_U4797, new_P1_U4798, new_P1_U4799,
    new_P1_U4800, new_P1_U4801, new_P1_U4802, new_P1_U4803, new_P1_U4804,
    new_P1_U4805, new_P1_U4806, new_P1_U4807, new_P1_U4808, new_P1_U4809,
    new_P1_U4810, new_P1_U4811, new_P1_U4812, new_P1_U4813, new_P1_U4814,
    new_P1_U4815, new_P1_U4816, new_P1_U4817, new_P1_U4818, new_P1_U4819,
    new_P1_U4820, new_P1_U4821, new_P1_U4822, new_P1_U4823, new_P1_U4824,
    new_P1_U4825, new_P1_U4826, new_P1_U4827, new_P1_U4828, new_P1_U4829,
    new_P1_U4830, new_P1_U4831, new_P1_U4832, new_P1_U4833, new_P1_U4834,
    new_P1_U4835, new_P1_U4836, new_P1_U4837, new_P1_U4838, new_P1_U4839,
    new_P1_U4840, new_P1_U4841, new_P1_U4842, new_P1_U4843, new_P1_U4844,
    new_P1_U4845, new_P1_U4846, new_P1_U4847, new_P1_U4848, new_P1_U4849,
    new_P1_U4850, new_P1_U4851, new_P1_U4852, new_P1_U4853, new_P1_U4854,
    new_P1_U4855, new_P1_U4856, new_P1_U4857, new_P1_U4858, new_P1_U4859,
    new_P1_U4860, new_P1_U4861, new_P1_U4862, new_P1_U4863, new_P1_U4864,
    new_P1_U4865, new_P1_U4866, new_P1_U4867, new_P1_U4868, new_P1_U4869,
    new_P1_U4870, new_P1_U4871, new_P1_U4872, new_P1_U4873, new_P1_U4874,
    new_P1_U4875, new_P1_U4876, new_P1_U4877, new_P1_U4878, new_P1_U4879,
    new_P1_U4880, new_P1_U4881, new_P1_U4882, new_P1_U4883, new_P1_U4884,
    new_P1_U4885, new_P1_U4886, new_P1_U4887, new_P1_U4888, new_P1_U4889,
    new_P1_U4890, new_P1_U4891, new_P1_U4892, new_P1_U4893, new_P1_U4894,
    new_P1_U4895, new_P1_U4896, new_P1_U4897, new_P1_U4898, new_P1_U4899,
    new_P1_U4900, new_P1_U4901, new_P1_U4902, new_P1_U4903, new_P1_U4904,
    new_P1_U4905, new_P1_U4906, new_P1_U4907, new_P1_U4908, new_P1_U4909,
    new_P1_U4910, new_P1_U4911, new_P1_U4912, new_P1_U4913, new_P1_U4914,
    new_P1_U4915, new_P1_U4916, new_P1_U4917, new_P1_U4918, new_P1_U4919,
    new_P1_U4920, new_P1_U4921, new_P1_U4922, new_P1_U4923, new_P1_U4924,
    new_P1_U4925, new_P1_U4926, new_P1_U4927, new_P1_U4928, new_P1_U4929,
    new_P1_U4930, new_P1_U4931, new_P1_U4932, new_P1_U4933, new_P1_U4934,
    new_P1_U4935, new_P1_U4936, new_P1_U4937, new_P1_U4938, new_P1_U4939,
    new_P1_U4940, new_P1_U4941, new_P1_U4942, new_P1_U4943, new_P1_U4944,
    new_P1_U4945, new_P1_U4946, new_P1_U4947, new_P1_U4948, new_P1_U4949,
    new_P1_U4950, new_P1_U4951, new_P1_U4952, new_P1_U4953, new_P1_U4954,
    new_P1_U4955, new_P1_U4956, new_P1_U4957, new_P1_U4958, new_P1_U4959,
    new_P1_U4960, new_P1_U4961, new_P1_U4962, new_P1_U4963, new_P1_U4964,
    new_P1_U4965, new_P1_U4966, new_P1_U4967, new_P1_U4968, new_P1_U4969,
    new_P1_U4970, new_P1_U4971, new_P1_U4972, new_P1_U4973, new_P1_U4974,
    new_P1_U4975, new_P1_U4976, new_P1_U4977, new_P1_U4978, new_P1_U4979,
    new_P1_U4980, new_P1_U4981, new_P1_U4982, new_P1_U4983, new_P1_U4984,
    new_P1_U4985, new_P1_U4986, new_P1_U4987, new_P1_U4988, new_P1_U4989,
    new_P1_U4990, new_P1_U4991, new_P1_U4992, new_P1_U4993, new_P1_U4994,
    new_P1_U4995, new_P1_U4996, new_P1_U4997, new_P1_U4998, new_P1_U4999,
    new_P1_U5000, new_P1_U5001, new_P1_U5002, new_P1_U5003, new_P1_U5004,
    new_P1_U5005, new_P1_U5006, new_P1_U5007, new_P1_U5008, new_P1_U5009,
    new_P1_U5010, new_P1_U5011, new_P1_U5012, new_P1_U5013, new_P1_U5014,
    new_P1_U5015, new_P1_U5016, new_P1_U5017, new_P1_U5018, new_P1_U5019,
    new_P1_U5020, new_P1_U5021, new_P1_U5022, new_P1_U5023, new_P1_U5024,
    new_P1_U5025, new_P1_U5026, new_P1_U5027, new_P1_U5028, new_P1_U5029,
    new_P1_U5030, new_P1_U5031, new_P1_U5032, new_P1_U5033, new_P1_U5034,
    new_P1_U5035, new_P1_U5036, new_P1_U5037, new_P1_U5038, new_P1_U5039,
    new_P1_U5040, new_P1_U5041, new_P1_U5042, new_P1_U5043, new_P1_U5044,
    new_P1_U5045, new_P1_U5046, new_P1_U5047, new_P1_U5048, new_P1_U5049,
    new_P1_U5050, new_P1_U5051, new_P1_U5052, new_P1_U5053, new_P1_U5054,
    new_P1_U5055, new_P1_U5056, new_P1_U5057, new_P1_U5058, new_P1_U5059,
    new_P1_U5060, new_P1_U5061, new_P1_U5062, new_P1_U5063, new_P1_U5064,
    new_P1_U5065, new_P1_U5066, new_P1_U5067, new_P1_U5068, new_P1_U5069,
    new_P1_U5070, new_P1_U5071, new_P1_U5072, new_P1_U5073, new_P1_U5074,
    new_P1_U5075, new_P1_U5076, new_P1_U5077, new_P1_U5078, new_P1_U5079,
    new_P1_U5080, new_P1_U5081, new_P1_U5082, new_P1_U5083, new_P1_U5084,
    new_P1_U5085, new_P1_U5086, new_P1_U5087, new_P1_U5088, new_P1_U5089,
    new_P1_U5090, new_P1_U5091, new_P1_U5092, new_P1_U5093, new_P1_U5094,
    new_P1_U5095, new_P1_U5096, new_P1_U5097, new_P1_U5098, new_P1_U5099,
    new_P1_U5100, new_P1_U5101, new_P1_U5102, new_P1_U5103, new_P1_U5104,
    new_P1_U5105, new_P1_U5106, new_P1_U5107, new_P1_U5108, new_P1_U5109,
    new_P1_U5110, new_P1_U5111, new_P1_U5112, new_P1_U5113, new_P1_U5114,
    new_P1_U5115, new_P1_U5116, new_P1_U5117, new_P1_U5118, new_P1_U5119,
    new_P1_U5120, new_P1_U5121, new_P1_U5122, new_P1_U5123, new_P1_U5124,
    new_P1_U5125, new_P1_U5126, new_P1_U5127, new_P1_U5128, new_P1_U5129,
    new_P1_U5130, new_P1_U5131, new_P1_U5132, new_P1_U5133, new_P1_U5134,
    new_P1_U5135, new_P1_U5136, new_P1_U5137, new_P1_U5138, new_P1_U5139,
    new_P1_U5140, new_P1_U5141, new_P1_U5142, new_P1_U5143, new_P1_U5144,
    new_P1_U5145, new_P1_U5146, new_P1_U5147, new_P1_U5148, new_P1_U5149,
    new_P1_U5150, new_P1_U5151, new_P1_U5152, new_P1_U5153, new_P1_U5154,
    new_P1_U5155, new_P1_U5156, new_P1_U5157, new_P1_U5158, new_P1_U5159,
    new_P1_U5160, new_P1_U5161, new_P1_U5162, new_P1_U5163, new_P1_U5164,
    new_P1_U5165, new_P1_U5166, new_P1_U5167, new_P1_U5168, new_P1_U5169,
    new_P1_U5170, new_P1_U5171, new_P1_U5172, new_P1_U5173, new_P1_U5174,
    new_P1_U5175, new_P1_U5176, new_P1_U5177, new_P1_U5178, new_P1_U5179,
    new_P1_U5180, new_P1_U5181, new_P1_U5182, new_P1_U5183, new_P1_U5184,
    new_P1_U5185, new_P1_U5186, new_P1_U5187, new_P1_U5188, new_P1_U5189,
    new_P1_U5190, new_P1_U5191, new_P1_U5192, new_P1_U5193, new_P1_U5194,
    new_P1_U5195, new_P1_U5196, new_P1_U5197, new_P1_U5198, new_P1_U5199,
    new_P1_U5200, new_P1_U5201, new_P1_U5202, new_P1_U5203, new_P1_U5204,
    new_P1_U5205, new_P1_U5206, new_P1_U5207, new_P1_U5208, new_P1_U5209,
    new_P1_U5210, new_P1_U5211, new_P1_U5212, new_P1_U5213, new_P1_U5214,
    new_P1_U5215, new_P1_U5216, new_P1_U5217, new_P1_U5218, new_P1_U5219,
    new_P1_U5220, new_P1_U5221, new_P1_U5222, new_P1_U5223, new_P1_U5224,
    new_P1_U5225, new_P1_U5226, new_P1_U5227, new_P1_U5228, new_P1_U5229,
    new_P1_U5230, new_P1_U5231, new_P1_U5232, new_P1_U5233, new_P1_U5234,
    new_P1_U5235, new_P1_U5236, new_P1_U5237, new_P1_U5238, new_P1_U5239,
    new_P1_U5240, new_P1_U5241, new_P1_U5242, new_P1_U5243, new_P1_U5244,
    new_P1_U5245, new_P1_U5246, new_P1_U5247, new_P1_U5248, new_P1_U5249,
    new_P1_U5250, new_P1_U5251, new_P1_U5252, new_P1_U5253, new_P1_U5254,
    new_P1_U5255, new_P1_U5256, new_P1_U5257, new_P1_U5258, new_P1_U5259,
    new_P1_U5260, new_P1_U5261, new_P1_U5262, new_P1_U5263, new_P1_U5264,
    new_P1_U5265, new_P1_U5266, new_P1_U5267, new_P1_U5268, new_P1_U5269,
    new_P1_U5270, new_P1_U5271, new_P1_U5272, new_P1_U5273, new_P1_U5274,
    new_P1_U5275, new_P1_U5276, new_P1_U5277, new_P1_U5278, new_P1_U5279,
    new_P1_U5280, new_P1_U5281, new_P1_U5282, new_P1_U5283, new_P1_U5284,
    new_P1_U5285, new_P1_U5286, new_P1_U5287, new_P1_U5288, new_P1_U5289,
    new_P1_U5290, new_P1_U5291, new_P1_U5292, new_P1_U5293, new_P1_U5294,
    new_P1_U5295, new_P1_U5296, new_P1_U5297, new_P1_U5298, new_P1_U5299,
    new_P1_U5300, new_P1_U5301, new_P1_U5302, new_P1_U5303, new_P1_U5304,
    new_P1_U5305, new_P1_U5306, new_P1_U5307, new_P1_U5308, new_P1_U5309,
    new_P1_U5310, new_P1_U5311, new_P1_U5312, new_P1_U5313, new_P1_U5314,
    new_P1_U5315, new_P1_U5316, new_P1_U5317, new_P1_U5318, new_P1_U5319,
    new_P1_U5320, new_P1_U5321, new_P1_U5322, new_P1_U5323, new_P1_U5324,
    new_P1_U5325, new_P1_U5326, new_P1_U5327, new_P1_U5328, new_P1_U5329,
    new_P1_U5330, new_P1_U5331, new_P1_U5332, new_P1_U5333, new_P1_U5334,
    new_P1_U5335, new_P1_U5336, new_P1_U5337, new_P1_U5338, new_P1_U5339,
    new_P1_U5340, new_P1_U5341, new_P1_U5342, new_P1_U5343, new_P1_U5344,
    new_P1_U5345, new_P1_U5346, new_P1_U5347, new_P1_U5348, new_P1_U5349,
    new_P1_U5350, new_P1_U5351, new_P1_U5352, new_P1_U5353, new_P1_U5354,
    new_P1_U5355, new_P1_U5356, new_P1_U5357, new_P1_U5358, new_P1_U5359,
    new_P1_U5360, new_P1_U5361, new_P1_U5362, new_P1_U5363, new_P1_U5364,
    new_P1_U5365, new_P1_U5366, new_P1_U5367, new_P1_U5368, new_P1_U5369,
    new_P1_U5370, new_P1_U5371, new_P1_U5372, new_P1_U5373, new_P1_U5374,
    new_P1_U5375, new_P1_U5376, new_P1_U5377, new_P1_U5378, new_P1_U5379,
    new_P1_U5380, new_P1_U5381, new_P1_U5382, new_P1_U5383, new_P1_U5384,
    new_P1_U5385, new_P1_U5386, new_P1_U5387, new_P1_U5388, new_P1_U5389,
    new_P1_U5390, new_P1_U5391, new_P1_U5392, new_P1_U5393, new_P1_U5394,
    new_P1_U5395, new_P1_U5396, new_P1_U5397, new_P1_U5398, new_P1_U5399,
    new_P1_U5400, new_P1_U5401, new_P1_U5402, new_P1_U5403, new_P1_U5404,
    new_P1_U5405, new_P1_U5406, new_P1_U5407, new_P1_U5408, new_P1_U5409,
    new_P1_U5410, new_P1_U5411, new_P1_U5412, new_P1_U5413, new_P1_U5414,
    new_P1_U5415, new_P1_U5416, new_P1_U5417, new_P1_U5418, new_P1_U5419,
    new_P1_U5420, new_P1_U5421, new_P1_U5422, new_P1_U5423, new_P1_U5424,
    new_P1_U5425, new_P1_U5426, new_P1_U5427, new_P1_U5428, new_P1_U5429,
    new_P1_U5430, new_P1_U5431, new_P1_U5432, new_P1_U5433, new_P1_U5434,
    new_P1_U5435, new_P1_U5436, new_P1_U5437, new_P1_U5438, new_P1_U5439,
    new_P1_U5440, new_P1_U5441, new_P1_U5442, new_P1_U5443, new_P1_U5444,
    new_P1_U5445, new_P1_U5446, new_P1_U5447, new_P1_U5448, new_P1_U5449,
    new_P1_U5450, new_P1_U5451, new_P1_U5452, new_P1_U5453, new_P1_U5454,
    new_P1_U5455, new_P1_U5456, new_P1_U5457, new_P1_U5458, new_P1_U5459,
    new_P1_U5460, new_P1_U5461, new_P1_U5462, new_P1_U5463, new_P1_U5464,
    new_P1_U5465, new_P1_U5466, new_P1_U5467, new_P1_U5468, new_P1_U5469,
    new_P1_U5470, new_P1_U5471, new_P1_U5472, new_P1_U5473, new_P1_U5474,
    new_P1_U5475, new_P1_U5476, new_P1_U5477, new_P1_U5478, new_P1_U5479,
    new_P1_U5480, new_P1_U5481, new_P1_U5482, new_P1_U5483, new_P1_U5484,
    new_P1_U5485, new_P1_U5486, new_P1_U5487, new_P1_U5488, new_P1_U5489,
    new_P1_U5490, new_P1_U5491, new_P1_U5492, new_P1_U5493, new_P1_U5494,
    new_P1_U5495, new_P1_U5496, new_P1_U5497, new_P1_U5498, new_P1_U5499,
    new_P1_U5500, new_P1_U5501, new_P1_U5502, new_P1_U5503, new_P1_U5504,
    new_P1_U5505, new_P1_U5506, new_P1_U5507, new_P1_U5508, new_P1_U5509,
    new_P1_U5510, new_P1_U5511, new_P1_U5512, new_P1_U5513, new_P1_U5514,
    new_P1_U5515, new_P1_U5516, new_P1_U5517, new_P1_U5518, new_P1_U5519,
    new_P1_U5520, new_P1_U5521, new_P1_U5522, new_P1_U5523, new_P1_U5524,
    new_P1_U5525, new_P1_U5526, new_P1_U5527, new_P1_U5528, new_P1_U5529,
    new_P1_U5530, new_P1_U5531, new_P1_U5532, new_P1_U5533, new_P1_U5534,
    new_P1_U5535, new_P1_U5536, new_P1_U5537, new_P1_U5538, new_P1_U5539,
    new_P1_U5540, new_P1_U5541, new_P1_U5542, new_P1_U5543, new_P1_U5544,
    new_P1_U5545, new_P1_U5546, new_P1_U5547, new_P1_U5548, new_P1_U5549,
    new_P1_U5550, new_P1_U5551, new_P1_U5552, new_P1_U5553, new_P1_U5554,
    new_P1_U5555, new_P1_U5556, new_P1_U5557, new_P1_U5558, new_P1_U5559,
    new_P1_U5560, new_P1_U5561, new_P1_U5562, new_P1_U5563, new_P1_U5564,
    new_P1_U5565, new_P1_U5566, new_P1_U5567, new_P1_U5568, new_P1_U5569,
    new_P1_U5570, new_P1_U5571, new_P1_U5572, new_P1_U5573, new_P1_U5574,
    new_P1_U5575, new_P1_U5576, new_P1_U5577, new_P1_U5578, new_P1_U5579,
    new_P1_U5580, new_P1_U5581, new_P1_U5582, new_P1_U5583, new_P1_U5584,
    new_P1_U5585, new_P1_U5586, new_P1_U5587, new_P1_U5588, new_P1_U5589,
    new_P1_U5590, new_P1_U5591, new_P1_U5592, new_P1_U5593, new_P1_U5594,
    new_P1_U5595, new_P1_U5596, new_P1_U5597, new_P1_U5598, new_P1_U5599,
    new_P1_U5600, new_P1_U5601, new_P1_U5602, new_P1_U5603, new_P1_U5604,
    new_P1_U5605, new_P1_U5606, new_P1_U5607, new_P1_U5608, new_P1_U5609,
    new_P1_U5610, new_P1_U5611, new_P1_U5612, new_P1_U5613, new_P1_U5614,
    new_P1_U5615, new_P1_U5616, new_P1_U5617, new_P1_U5618, new_P1_U5619,
    new_P1_U5620, new_P1_U5621, new_P1_U5622, new_P1_U5623, new_P1_U5624,
    new_P1_U5625, new_P1_U5626, new_P1_U5627, new_P1_U5628, new_P1_U5629,
    new_P1_U5630, new_P1_U5631, new_P1_U5632, new_P1_U5633, new_P1_U5634,
    new_P1_U5635, new_P1_U5636, new_P1_U5637, new_P1_U5638, new_P1_U5639,
    new_P1_U5640, new_P1_U5641, new_P1_U5642, new_P1_U5643, new_P1_U5644,
    new_P1_U5645, new_P1_U5646, new_P1_U5647, new_P1_U5648, new_P1_U5649,
    new_P1_U5650, new_P1_U5651, new_P1_U5652, new_P1_U5653, new_P1_U5654,
    new_P1_U5655, new_P1_U5656, new_P1_U5657, new_P1_U5658, new_P1_U5659,
    new_P1_U5660, new_P1_U5661, new_P1_U5662, new_P1_U5663, new_P1_U5664,
    new_P1_U5665, new_P1_U5666, new_P1_U5667, new_P1_U5668, new_P1_U5669,
    new_P1_U5670, new_P1_U5671, new_P1_U5672, new_P1_U5673, new_P1_U5674,
    new_P1_U5675, new_P1_U5676, new_P1_U5677, new_P1_U5678, new_P1_U5679,
    new_P1_U5680, new_P1_U5681, new_P1_U5682, new_P1_U5683, new_P1_U5684,
    new_P1_U5685, new_P1_U5686, new_P1_U5687, new_P1_U5688, new_P1_U5689,
    new_P1_U5690, new_P1_U5691, new_P1_U5692, new_P1_U5693, new_P1_U5694,
    new_P1_U5695, new_P1_U5696, new_P1_U5697, new_P1_U5698, new_P1_U5699,
    new_P1_U5700, new_P1_U5701, new_P1_U5702, new_P1_U5703, new_P1_U5704,
    new_P1_U5705, new_P1_U5706, new_P1_U5707, new_P1_U5708, new_P1_U5709,
    new_P1_U5710, new_P1_U5711, new_P1_U5712, new_P1_U5713, new_P1_U5714,
    new_P1_U5715, new_P1_U5716, new_P1_U5717, new_P1_U5718, new_P1_U5719,
    new_P1_U5720, new_P1_U5721, new_P1_U5722, new_P1_U5723, new_P1_U5724,
    new_P1_U5725, new_P1_U5726, new_P1_U5727, new_P1_U5728, new_P1_U5729,
    new_P1_U5730, new_P1_U5731, new_P1_U5732, new_P1_U5733, new_P1_U5734,
    new_P1_U5735, new_P1_U5736, new_P1_U5737, new_P1_U5738, new_P1_U5739,
    new_P1_U5740, new_P1_U5741, new_P1_U5742, new_P1_U5743, new_P1_U5744,
    new_P1_U5745, new_P1_U5746, new_P1_U5747, new_P1_U5748, new_P1_U5749,
    new_P1_U5750, new_P1_U5751, new_P1_U5752, new_P1_U5753, new_P1_U5754,
    new_P1_U5755, new_P1_U5756, new_P1_U5757, new_P1_U5758, new_P1_U5759,
    new_P1_U5760, new_P1_U5761, new_P1_U5762, new_P1_U5763, new_P1_U5764,
    new_P1_U5765, new_P1_U5766, new_P1_U5767, new_P1_U5768, new_P1_U5769,
    new_P1_U5770, new_P1_U5771, new_P1_U5772, new_P1_U5773, new_P1_U5774,
    new_P1_U5775, new_P1_U5776, new_P1_U5777, new_P1_U5778, new_P1_U5779,
    new_P1_U5780, new_P1_U5781, new_P1_U5782, new_P1_U5783, new_P1_U5784,
    new_P1_U5785, new_P1_U5786, new_P1_U5787, new_P1_U5788, new_P1_U5789,
    new_P1_U5790, new_P1_U5791, new_P1_U5792, new_P1_U5793, new_P1_U5794,
    new_P1_U5795, new_P1_U5796, new_P1_U5797, new_P1_U5798, new_P1_U5799,
    new_P1_U5800, new_P1_U5801, new_P1_U5802, new_P1_U5803, new_P1_U5804,
    new_P1_U5805, new_P1_U5806, new_P1_U5807, new_P1_U5808, new_P1_U5809,
    new_P1_U5810, new_P1_U5811, new_P1_U5812, new_P1_U5813, new_P1_U5814,
    new_P1_U5815, new_P1_U5816, new_P1_U5817, new_P1_U5818, new_P1_U5819,
    new_P1_U5820, new_P1_U5821, new_P1_U5822, new_P1_U5823, new_P1_U5824,
    new_P1_U5825, new_P1_U5826, new_P1_U5827, new_P1_U5828, new_P1_U5829,
    new_P1_U5830, new_P1_U5831, new_P1_U5832, new_P1_U5833, new_P1_U5834,
    new_P1_U5835, new_P1_U5836, new_P1_U5837, new_P1_U5838, new_P1_U5839,
    new_P1_U5840, new_P1_U5841, new_P1_U5842, new_P1_U5843, new_P1_U5844,
    new_P1_U5845, new_P1_U5846, new_P1_U5847, new_P1_U5848, new_P1_U5849,
    new_P1_U5850, new_P1_U5851, new_P1_U5852, new_P1_U5853, new_P1_U5854,
    new_P1_U5855, new_P1_U5856, new_P1_U5857, new_P1_U5858, new_P1_U5859,
    new_P1_U5860, new_P1_U5861, new_P1_U5862, new_P1_U5863, new_P1_U5864,
    new_P1_U5865, new_P1_U5866, new_P1_U5867, new_P1_U5868, new_P1_U5869,
    new_P1_U5870, new_P1_U5871, new_P1_U5872, new_P1_U5873, new_P1_U5874,
    new_P1_U5875, new_P1_U5876, new_P1_U5877, new_P1_U5878, new_P1_U5879,
    new_P1_U5880, new_P1_U5881, new_P1_U5882, new_P1_U5883, new_P1_U5884,
    new_P1_U5885, new_P1_U5886, new_P1_U5887, new_P1_U5888, new_P1_U5889,
    new_P1_U5890, new_P1_U5891, new_P1_U5892, new_P1_U5893, new_P1_U5894,
    new_P1_U5895, new_P1_U5896, new_P1_U5897, new_P1_U5898, new_P1_U5899,
    new_P1_U5900, new_P1_U5901, new_P1_U5902, new_P1_U5903, new_P1_U5904,
    new_P1_U5905, new_P1_U5906, new_P1_U5907, new_P1_U5908, new_P1_U5909,
    new_P1_U5910, new_P1_U5911, new_P1_U5912, new_P1_U5913, new_P1_U5914,
    new_P1_U5915, new_P1_U5916, new_P1_U5917, new_P1_U5918, new_P1_U5919,
    new_P1_U5920, new_P1_U5921, new_P1_U5922, new_P1_U5923, new_P1_U5924,
    new_P1_U5925, new_P1_U5926, new_P1_U5927, new_P1_U5928, new_P1_U5929,
    new_P1_U5930, new_P1_U5931, new_P1_U5932, new_P1_U5933, new_P1_U5934,
    new_P1_U5935, new_P1_U5936, new_P1_U5937, new_P1_U5938, new_P1_U5939,
    new_P1_U5940, new_P1_U5941, new_P1_U5942, new_P1_U5943, new_P1_U5944,
    new_P1_U5945, new_P1_U5946, new_P1_U5947, new_P1_U5948, new_P1_U5949,
    new_P1_U5950, new_P1_U5951, new_P1_U5952, new_P1_U5953, new_P1_U5954,
    new_P1_U5955, new_P1_U5956, new_P1_U5957, new_P1_U5958, new_P1_U5959,
    new_P1_U5960, new_P1_U5961, new_P1_U5962, new_P1_U5963, new_P1_U5964,
    new_P1_U5965, new_P1_U5966, new_P1_U5967, new_P1_U5968, new_P1_U5969,
    new_P1_U5970, new_P1_U5971, new_P1_U5972, new_P1_U5973, new_P1_U5974,
    new_P1_U5975, new_P1_U5976, new_P1_U5977, new_P1_U5978, new_P1_U5979,
    new_P1_U5980, new_P1_U5981, new_P1_U5982, new_P1_U5983, new_P1_U5984,
    new_P1_U5985, new_P1_U5986, new_P1_U5987, new_P1_U5988, new_P1_U5989,
    new_P1_U5990, new_P1_U5991, new_P1_U5992, new_P1_U5993, new_P1_U5994,
    new_P1_U5995, new_P1_U5996, new_P1_U5997, new_P1_U5998, new_P1_U5999,
    new_P1_U6000, new_P1_U6001, new_P1_U6002, new_P1_U6003, new_P1_U6004,
    new_P1_U6005, new_P1_U6006, new_P1_U6007, new_P1_U6008, new_P1_U6009,
    new_P1_U6010, new_P1_U6011, new_P1_U6012, new_P1_U6013, new_P1_U6014,
    new_P1_U6015, new_P1_U6016, new_P1_U6017, new_P1_U6018, new_P1_U6019,
    new_P1_U6020, new_P1_U6021, new_P1_U6022, new_P1_U6023, new_P1_U6024,
    new_P1_U6025, new_P1_U6026, new_P1_U6027, new_P1_U6028, new_P1_U6029,
    new_P1_U6030, new_P1_U6031, new_P1_U6032, new_P1_U6033, new_P1_U6034,
    new_P1_U6035, new_P1_U6036, new_P1_U6037, new_P1_U6038, new_P1_U6039,
    new_P1_U6040, new_P1_U6041, new_P1_U6042, new_P1_U6043, new_P1_U6044,
    new_P1_U6045, new_P1_U6046, new_P1_U6047, new_P1_U6048, new_P1_U6049,
    new_P1_U6050, new_P1_U6051, new_P1_U6052, new_P1_U6053, new_P1_U6054,
    new_P1_U6055, new_P1_U6056, new_P1_U6057, new_P1_U6058, new_P1_U6059,
    new_P1_U6060, new_P1_U6061, new_P1_U6062, new_P1_U6063, new_P1_U6064,
    new_P1_U6065, new_P1_U6066, new_P1_U6067, new_P1_U6068, new_P1_U6069,
    new_P1_U6070, new_P1_U6071, new_P1_U6072, new_P1_U6073, new_P1_U6074,
    new_P1_U6075, new_P1_U6076, new_P1_U6077, new_P1_U6078, new_P1_U6079,
    new_P1_U6080, new_P1_U6081, new_P1_U6082, new_P1_U6083, new_P1_U6084,
    new_P1_U6085, new_P1_U6086, new_P1_U6087, new_P1_U6088, new_P1_U6089,
    new_P1_U6090, new_P1_U6091, new_P1_U6092, new_P1_U6093, new_P1_U6094,
    new_P1_U6095, new_P1_U6096, new_P1_U6097, new_P1_U6098, new_P1_U6099,
    new_P1_U6100, new_P1_U6101, new_P1_U6102, new_P1_U6103, new_P1_U6104,
    new_P1_U6105, new_P1_U6106, new_P1_U6107, new_P1_U6108, new_P1_U6109,
    new_P1_U6110, new_P1_U6111, new_P1_U6112, new_P1_U6113, new_P1_U6114,
    new_P1_U6115, new_P1_U6116, new_P1_U6117, new_P1_U6118, new_P1_U6119,
    new_P1_U6120, new_P1_U6121, new_P1_U6122, new_P1_U6123, new_P1_U6124,
    new_P1_U6125, new_P1_U6126, new_P1_U6127, new_P1_U6128, new_P1_U6129,
    new_P1_U6130, new_P1_U6131, new_P1_U6132, new_P1_U6133, new_P1_U6134,
    new_P1_U6135, new_P1_U6136, new_P1_U6137, new_P1_U6138, new_P1_U6139,
    new_P1_U6140, new_P1_U6141, new_P1_U6142, new_P1_U6143, new_P1_U6144,
    new_P1_U6145, new_P1_U6146, new_P1_U6147, new_P1_U6148, new_P1_U6149,
    new_P1_U6150, new_P1_U6151, new_P1_U6152, new_P1_U6153, new_P1_U6154,
    new_P1_U6155, new_P1_U6156, new_P1_U6157, new_P1_U6158, new_P1_U6159,
    new_P1_U6160, new_P1_U6161, new_P1_U6162, new_P1_U6163, new_P1_U6164,
    new_P1_U6165, new_P1_U6166, new_P1_U6167, new_P1_U6168, new_P1_U6169,
    new_P1_U6170, new_P1_U6171, new_P1_U6172, new_P1_U6173, new_P1_U6174,
    new_P1_U6175, new_P1_U6176, new_P1_U6177, new_P1_U6178, new_P1_U6179,
    new_P1_U6180, new_P1_U6181, new_P1_U6182, new_P1_U6183, new_P1_U6184,
    new_P1_U6185, new_P1_U6186, new_P1_U6187, new_P1_U6188, new_P1_U6189,
    new_P1_U6190, new_P1_U6191, new_P1_U6192, new_P1_U6193, new_P1_U6194,
    new_P1_U6195, new_P1_U6196, new_P1_U6197, new_P1_U6198, new_P1_U6199,
    new_P1_U6200, new_P1_U6201, new_P1_U6202, new_P1_U6203, new_P1_U6204,
    new_P1_U6205, new_P1_U6206, new_P1_U6207, new_P1_U6208, new_P1_U6209,
    new_P1_U6210, new_P1_U6211, new_P1_U6212, new_P1_U6213, new_P1_U6214,
    new_P1_U6215, new_P1_U6216, new_P1_U6217, new_P1_U6218, new_P1_U6219,
    new_P1_U6220, new_P1_U6221, new_P1_U6222, new_P1_U6223, new_P1_U6224,
    new_P1_U6225, new_P1_U6226, new_P1_U6227, new_P1_U6228, new_P1_U6229,
    new_P1_U6230, new_P1_U6231, new_P1_U6232, new_P1_U6233, new_P1_U6234,
    new_P1_U6235, new_P1_U6236, new_P1_U6237, new_P1_U6238, new_P1_U6239,
    new_P1_U6240, new_P1_U6241, new_P1_U6242, new_P1_U6243, new_P1_U6244,
    new_P1_U6245, new_P1_U6246, new_P1_U6247, new_P1_U6248, new_P1_U6249,
    new_P1_U6250, new_P1_U6251, new_P1_U6252, new_P1_U6253, new_P1_U6254,
    new_P1_U6255, new_P1_U6256, new_P1_U6257, new_P1_U6258, new_P1_U6259,
    new_P1_U6260, new_P1_U6261, new_P1_U6262, new_P1_U6263, new_P1_U6264,
    new_P1_U6265, new_P1_U6266, new_P1_U6267, new_P1_U6268, new_P1_U6269,
    new_P1_U6270, new_P1_U6271, new_P1_U6272, new_P1_U6273, new_P1_U6274,
    new_P1_U6275, new_P1_U6276, new_P1_U6277, new_P1_U6278, new_P1_U6279,
    new_P1_U6280, new_P1_U6281, new_P1_U6282, new_P1_U6283, new_P1_U6284,
    new_P1_U6285, new_P3_R1161_U489, new_P3_R1161_U488, new_P3_R1161_U487,
    new_P3_R1161_U486, new_P3_R1161_U485, new_P3_R1161_U484,
    new_P3_R1161_U483, new_P3_R1161_U482, new_P3_R1161_U481,
    new_P3_R1161_U480, new_P3_R1161_U479, new_P3_R1161_U478,
    new_P3_R1161_U477, new_P3_R1161_U476, new_P3_R1161_U475,
    new_P3_R1161_U474, new_P3_R1161_U473, new_P3_R1161_U472,
    new_P3_R1161_U471, new_P3_R1161_U470, new_P3_R1161_U469, new_P2_U3014,
    new_P2_U3015, new_P2_U3016, new_P2_U3017, new_P2_U3018, new_P2_U3019,
    new_P2_U3020, new_P2_U3021, new_P2_U3022, new_P2_U3023, new_P2_U3024,
    new_P2_U3025, new_P2_U3026, new_P2_U3027, new_P2_U3028, new_P2_U3029,
    new_P2_U3030, new_P2_U3031, new_P2_U3032, new_P2_U3033, new_P2_U3034,
    new_P2_U3035, new_P2_U3036, new_P2_U3037, new_P2_U3038, new_P2_U3039,
    new_P2_U3040, new_P2_U3041, new_P2_U3042, new_P2_U3043, new_P2_U3044,
    new_P2_U3045, new_P2_U3046, new_P2_U3047, new_P2_U3048, new_P2_U3049,
    new_P2_U3050, new_P2_U3051, new_P2_U3052, new_P2_U3053, new_P2_U3054,
    new_P2_U3055, new_P2_U3056, new_P2_U3057, new_P2_U3058, new_P2_U3059,
    new_P2_U3060, new_P2_U3061, new_P2_U3062, new_P2_U3063, new_P2_U3064,
    new_P2_U3065, new_P2_U3066, new_P2_U3067, new_P2_U3068, new_P2_U3069,
    new_P2_U3070, new_P2_U3071, new_P2_U3072, new_P2_U3073, new_P2_U3074,
    new_P2_U3075, new_P2_U3076, new_P2_U3077, new_P2_U3078, new_P2_U3079,
    new_P2_U3080, new_P2_U3081, new_P2_U3082, new_P2_U3083, new_P2_U3084,
    new_P2_U3085, new_P2_U3086, new_P2_U3089, new_P2_U3090, new_P2_U3091,
    new_P2_U3092, new_P2_U3093, new_P2_U3094, new_P2_U3095, new_P2_U3096,
    new_P2_U3097, new_P2_U3098, new_P2_U3099, new_P2_U3100, new_P2_U3101,
    new_P2_U3102, new_P2_U3103, new_P2_U3104, new_P2_U3105, new_P2_U3106,
    new_P2_U3107, new_P2_U3108, new_P2_U3109, new_P2_U3110, new_P2_U3111,
    new_P2_U3112, new_P2_U3113, new_P2_U3114, new_P2_U3115, new_P2_U3116,
    new_P2_U3117, new_P2_U3118, new_P2_U3119, new_P2_U3120, new_P2_U3121,
    new_P2_U3122, new_P2_U3123, new_P2_U3124, new_P2_U3125, new_P2_U3126,
    new_P2_U3127, new_P2_U3128, new_P2_U3129, new_P2_U3130, new_P2_U3131,
    new_P2_U3132, new_P2_U3133, new_P2_U3134, new_P2_U3135, new_P2_U3136,
    new_P2_U3137, new_P2_U3138, new_P2_U3139, new_P2_U3140, new_P2_U3141,
    new_P2_U3142, new_P2_U3143, new_P2_U3144, new_P2_U3145, new_P2_U3146,
    new_P2_U3147, new_P2_U3148, new_P2_U3149, new_P2_U3150, new_P2_U3151,
    new_P2_U3152, new_P2_U3153, new_P2_U3154, new_P2_U3155, new_P2_U3156,
    new_P2_U3157, new_P2_U3158, new_P2_U3159, new_P2_U3160, new_P2_U3161,
    new_P2_U3162, new_P2_U3163, new_P2_U3164, new_P2_U3165, new_P2_U3166,
    new_P2_U3167, new_P2_U3168, new_P2_U3169, new_P2_U3170, new_P2_U3171,
    new_P2_U3172, new_P2_U3173, new_P2_U3174, new_P2_U3175, new_P2_U3176,
    new_P2_U3177, new_P2_U3178, new_P2_U3179, new_P2_U3180, new_P2_U3181,
    new_P2_U3182, new_P2_U3183, new_P2_U3184, new_P2_U3329, new_P2_U3330,
    new_P2_U3331, new_P2_U3332, new_P2_U3333, new_P2_U3334, new_P2_U3335,
    new_P2_U3336, new_P2_U3337, new_P2_U3338, new_P2_U3339, new_P2_U3340,
    new_P2_U3341, new_P2_U3342, new_P2_U3343, new_P2_U3344, new_P2_U3345,
    new_P2_U3346, new_P2_U3347, new_P2_U3348, new_P2_U3349, new_P2_U3350,
    new_P2_U3351, new_P2_U3352, new_P2_U3353, new_P2_U3354, new_P2_U3355,
    new_P2_U3356, new_P2_U3357, new_P2_U3358, new_P2_U3359, new_P2_U3360,
    new_P2_U3361, new_P2_U3362, new_P2_U3363, new_P2_U3364, new_P2_U3365,
    new_P2_U3366, new_P2_U3367, new_P2_U3368, new_P2_U3369, new_P2_U3370,
    new_P2_U3371, new_P2_U3372, new_P2_U3373, new_P2_U3374, new_P2_U3375,
    new_P2_U3376, new_P2_U3377, new_P2_U3378, new_P2_U3379, new_P2_U3380,
    new_P2_U3381, new_P2_U3382, new_P2_U3383, new_P2_U3384, new_P2_U3385,
    new_P2_U3386, new_P2_U3387, new_P2_U3388, new_P2_U3389, new_P2_U3390,
    new_P2_U3391, new_P2_U3392, new_P2_U3393, new_P2_U3394, new_P2_U3395,
    new_P2_U3396, new_P2_U3397, new_P2_U3398, new_P2_U3399, new_P2_U3400,
    new_P2_U3401, new_P2_U3402, new_P2_U3403, new_P2_U3404, new_P2_U3405,
    new_P2_U3406, new_P2_U3407, new_P2_U3408, new_P2_U3409, new_P2_U3410,
    new_P2_U3411, new_P2_U3412, new_P2_U3413, new_P2_U3414, new_P2_U3415,
    new_P2_U3418, new_P2_U3419, new_P2_U3420, new_P2_U3421, new_P2_U3422,
    new_P2_U3423, new_P2_U3424, new_P2_U3425, new_P2_U3426, new_P2_U3427,
    new_P2_U3428, new_P2_U3429, new_P2_U3431, new_P2_U3432, new_P2_U3434,
    new_P2_U3435, new_P2_U3437, new_P2_U3438, new_P2_U3440, new_P2_U3441,
    new_P2_U3443, new_P2_U3444, new_P2_U3446, new_P2_U3447, new_P2_U3449,
    new_P2_U3450, new_P2_U3452, new_P2_U3453, new_P2_U3455, new_P2_U3456,
    new_P2_U3458, new_P2_U3459, new_P2_U3461, new_P2_U3462, new_P2_U3464,
    new_P2_U3465, new_P2_U3467, new_P2_U3468, new_P2_U3470, new_P2_U3471,
    new_P2_U3473, new_P2_U3474, new_P2_U3476, new_P2_U3477, new_P2_U3479,
    new_P2_U3480, new_P2_U3482, new_P2_U3483, new_P2_U3485, new_P2_U3563,
    new_P2_U3564, new_P2_U3565, new_P2_U3566, new_P2_U3567, new_P2_U3568,
    new_P2_U3569, new_P2_U3570, new_P2_U3571, new_P2_U3572, new_P2_U3573,
    new_P2_U3574, new_P2_U3575, new_P2_U3576, new_P2_U3577, new_P2_U3578,
    new_P2_U3579, new_P2_U3580, new_P2_U3581, new_P2_U3582, new_P2_U3583,
    new_P2_U3584, new_P2_U3585, new_P2_U3586, new_P2_U3587, new_P2_U3588,
    new_P2_U3589, new_P2_U3590, new_P2_U3591, new_P2_U3592, new_P2_U3593,
    new_P2_U3594, new_P2_U3595, new_P2_U3596, new_P2_U3597, new_P2_U3598,
    new_P2_U3599, new_P2_U3600, new_P2_U3601, new_P2_U3602, new_P2_U3603,
    new_P2_U3604, new_P2_U3605, new_P2_U3606, new_P2_U3607, new_P2_U3608,
    new_P2_U3609, new_P2_U3610, new_P2_U3611, new_P2_U3612, new_P2_U3613,
    new_P2_U3614, new_P2_U3615, new_P2_U3616, new_P2_U3617, new_P2_U3618,
    new_P2_U3619, new_P2_U3620, new_P2_U3621, new_P2_U3622, new_P2_U3623,
    new_P2_U3624, new_P2_U3625, new_P2_U3626, new_P2_U3627, new_P2_U3628,
    new_P2_U3629, new_P2_U3630, new_P2_U3631, new_P2_U3632, new_P2_U3633,
    new_P2_U3634, new_P2_U3635, new_P2_U3636, new_P2_U3637, new_P2_U3638,
    new_P2_U3639, new_P2_U3640, new_P2_U3641, new_P2_U3642, new_P2_U3643,
    new_P2_U3644, new_P2_U3645, new_P2_U3646, new_P2_U3647, new_P2_U3648,
    new_P2_U3649, new_P2_U3650, new_P2_U3651, new_P2_U3652, new_P2_U3653,
    new_P2_U3654, new_P2_U3655, new_P2_U3656, new_P2_U3657, new_P2_U3658,
    new_P2_U3659, new_P2_U3660, new_P2_U3661, new_P2_U3662, new_P2_U3663,
    new_P2_U3664, new_P2_U3665, new_P2_U3666, new_P2_U3667, new_P2_U3668,
    new_P2_U3669, new_P2_U3670, new_P2_U3671, new_P2_U3672, new_P2_U3673,
    new_P2_U3674, new_P2_U3675, new_P2_U3676, new_P2_U3677, new_P2_U3678,
    new_P2_U3679, new_P2_U3680, new_P2_U3681, new_P2_U3682, new_P2_U3683,
    new_P2_U3684, new_P2_U3685, new_P2_U3686, new_P2_U3687, new_P2_U3688,
    new_P2_U3689, new_P2_U3690, new_P2_U3691, new_P2_U3692, new_P2_U3693,
    new_P2_U3694, new_P2_U3695, new_P2_U3696, new_P2_U3697, new_P2_U3698,
    new_P2_U3699, new_P2_U3700, new_P2_U3701, new_P2_U3702, new_P2_U3703,
    new_P2_U3704, new_P2_U3705, new_P2_U3706, new_P2_U3707, new_P2_U3708,
    new_P2_U3709, new_P2_U3710, new_P2_U3711, new_P2_U3712, new_P2_U3713,
    new_P2_U3714, new_P2_U3715, new_P2_U3716, new_P2_U3717, new_P2_U3718,
    new_P2_U3719, new_P2_U3720, new_P2_U3721, new_P2_U3722, new_P2_U3723,
    new_P2_U3724, new_P2_U3725, new_P2_U3726, new_P2_U3727, new_P2_U3728,
    new_P2_U3729, new_P2_U3730, new_P2_U3731, new_P2_U3732, new_P2_U3733,
    new_P2_U3734, new_P2_U3735, new_P2_U3736, new_P2_U3737, new_P2_U3738,
    new_P2_U3739, new_P2_U3740, new_P2_U3741, new_P2_U3742, new_P2_U3743,
    new_P2_U3744, new_P2_U3745, new_P2_U3746, new_P2_U3747, new_P2_U3748,
    new_P2_U3749, new_P2_U3750, new_P2_U3751, new_P2_U3752, new_P2_U3753,
    new_P2_U3754, new_P2_U3755, new_P2_U3756, new_P2_U3757, new_P2_U3758,
    new_P2_U3759, new_P2_U3760, new_P2_U3761, new_P2_U3762, new_P2_U3763,
    new_P2_U3764, new_P2_U3765, new_P2_U3766, new_P2_U3767, new_P2_U3768,
    new_P2_U3769, new_P2_U3770, new_P2_U3771, new_P2_U3772, new_P2_U3773,
    new_P2_U3774, new_P2_U3775, new_P2_U3776, new_P2_U3777, new_P2_U3778,
    new_P2_U3779, new_P2_U3780, new_P2_U3781, new_P2_U3782, new_P2_U3783,
    new_P2_U3784, new_P2_U3785, new_P2_U3786, new_P2_U3787, new_P2_U3788,
    new_P2_U3789, new_P2_U3790, new_P2_U3791, new_P2_U3792, new_P2_U3793,
    new_P2_U3794, new_P2_U3795, new_P2_U3796, new_P2_U3797, new_P2_U3798,
    new_P2_U3799, new_P2_U3800, new_P2_U3801, new_P2_U3802, new_P2_U3803,
    new_P2_U3804, new_P2_U3805, new_P2_U3806, new_P2_U3807, new_P2_U3808,
    new_P2_U3809, new_P2_U3810, new_P2_U3811, new_P2_U3812, new_P2_U3813,
    new_P2_U3814, new_P2_U3815, new_P2_U3816, new_P2_U3817, new_P2_U3818,
    new_P2_U3819, new_P2_U3820, new_P2_U3821, new_P2_U3822, new_P2_U3823,
    new_P2_U3824, new_P2_U3825, new_P2_U3826, new_P2_U3827, new_P2_U3828,
    new_P2_U3829, new_P2_U3830, new_P2_U3831, new_P2_U3832, new_P2_U3833,
    new_P2_U3834, new_P2_U3835, new_P2_U3836, new_P2_U3837, new_P2_U3838,
    new_P2_U3839, new_P2_U3840, new_P2_U3841, new_P2_U3842, new_P2_U3843,
    new_P2_U3844, new_P2_U3845, new_P2_U3846, new_P2_U3847, new_P2_U3848,
    new_P2_U3849, new_P2_U3850, new_P2_U3851, new_P2_U3852, new_P2_U3853,
    new_P2_U3854, new_P2_U3855, new_P2_U3856, new_P2_U3857, new_P2_U3858,
    new_P2_U3859, new_P2_U3860, new_P2_U3861, new_P2_U3862, new_P2_U3863,
    new_P2_U3864, new_P2_U3865, new_P2_U3866, new_P2_U3867, new_P2_U3868,
    new_P2_U3869, new_P2_U3870, new_P2_U3871, new_P2_U3872, new_P2_U3873,
    new_P2_U3874, new_P2_U3875, new_P2_U3876, new_P2_U3877, new_P2_U3878,
    new_P2_U3879, new_P2_U3880, new_P2_U3881, new_P2_U3882, new_P2_U3883,
    new_P2_U3884, new_P2_U3885, new_P2_U3886, new_P2_U3887, new_P2_U3888,
    new_P2_U3889, new_P2_U3890, new_P2_U3891, new_P2_U3892, new_P2_U3893,
    new_P2_U3894, new_P2_U3895, new_P2_U3896, new_P2_U3897, new_P2_U3898,
    new_P2_U3899, new_P2_U3900, new_P2_U3901, new_P2_U3902, new_P2_U3903,
    new_P2_U3904, new_P2_U3905, new_P2_U3906, new_P2_U3907, new_P2_U3908,
    new_P2_U3909, new_P2_U3910, new_P2_U3911, new_P2_U3912, new_P2_U3913,
    new_P2_U3914, new_P2_U3915, new_P2_U3916, new_P2_U3917, new_P2_U3918,
    new_P2_U3919, new_P2_U3920, new_P2_U3921, new_P2_U3922, new_P2_U3923,
    new_P2_U3924, new_P2_U3925, new_P2_U3926, new_P2_U3927, new_P2_U3928,
    new_P2_U3929, new_P2_U3930, new_P2_U3931, new_P2_U3932, new_P2_U3933,
    new_P2_U3934, new_P2_U3935, new_P2_U3936, new_P2_U3937, new_P2_U3938,
    new_P2_U3939, new_P2_U3940, new_P2_U3941, new_P2_U3942, new_P2_U3943,
    new_P2_U3944, new_P2_U3945, new_P2_U3946, new_P2_U3948, new_P2_U3949,
    new_P2_U3950, new_P2_U3951, new_P2_U3952, new_P2_U3953, new_P2_U3954,
    new_P2_U3955, new_P2_U3956, new_P2_U3957, new_P2_U3958, new_P2_U3959,
    new_P2_U3960, new_P2_U3961, new_P2_U3962, new_P2_U3963, new_P2_U3964,
    new_P2_U3965, new_P2_U3966, new_P2_U3967, new_P2_U3968, new_P2_U3969,
    new_P2_U3970, new_P2_U3971, new_P2_U3972, new_P2_U3973, new_P2_U3974,
    new_P2_U3975, new_P2_U3976, new_P2_U3977, new_P2_U3978, new_P2_U3979,
    new_P2_U3980, new_P2_U3981, new_P2_U3982, new_P2_U3983, new_P2_U3984,
    new_P2_U3985, new_P2_U3986, new_P2_U3987, new_P2_U3988, new_P2_U3989,
    new_P2_U3990, new_P2_U3991, new_P2_U3992, new_P2_U3993, new_P2_U3994,
    new_P2_U3995, new_P2_U3996, new_P2_U3997, new_P2_U3998, new_P2_U3999,
    new_P2_U4000, new_P2_U4001, new_P2_U4002, new_P2_U4003, new_P2_U4004,
    new_P2_U4005, new_P2_U4006, new_P2_U4007, new_P2_U4008, new_P2_U4009,
    new_P2_U4010, new_P2_U4011, new_P2_U4012, new_P2_U4013, new_P2_U4014,
    new_P2_U4015, new_P2_U4016, new_P2_U4017, new_P2_U4018, new_P2_U4019,
    new_P2_U4020, new_P2_U4021, new_P2_U4022, new_P2_U4023, new_P2_U4024,
    new_P2_U4025, new_P2_U4026, new_P2_U4027, new_P2_U4028, new_P2_U4029,
    new_P2_U4030, new_P2_U4031, new_P2_U4032, new_P2_U4033, new_P2_U4034,
    new_P2_U4035, new_P2_U4036, new_P2_U4037, new_P2_U4038, new_P2_U4039,
    new_P2_U4040, new_P2_U4041, new_P2_U4042, new_P2_U4043, new_P2_U4044,
    new_P2_U4045, new_P2_U4046, new_P2_U4047, new_P2_U4048, new_P2_U4049,
    new_P2_U4050, new_P2_U4051, new_P2_U4052, new_P2_U4053, new_P2_U4054,
    new_P2_U4055, new_P2_U4056, new_P2_U4057, new_P2_U4058, new_P2_U4059,
    new_P2_U4060, new_P2_U4061, new_P2_U4062, new_P2_U4063, new_P2_U4064,
    new_P2_U4065, new_P2_U4066, new_P2_U4067, new_P2_U4068, new_P2_U4069,
    new_P2_U4070, new_P2_U4071, new_P2_U4072, new_P2_U4073, new_P2_U4074,
    new_P2_U4075, new_P2_U4076, new_P2_U4077, new_P2_U4078, new_P2_U4079,
    new_P2_U4080, new_P2_U4081, new_P2_U4082, new_P2_U4083, new_P2_U4084,
    new_P2_U4085, new_P2_U4086, new_P2_U4087, new_P2_U4088, new_P2_U4089,
    new_P2_U4090, new_P2_U4091, new_P2_U4092, new_P2_U4093, new_P2_U4094,
    new_P2_U4095, new_P2_U4096, new_P2_U4097, new_P2_U4098, new_P2_U4099,
    new_P2_U4100, new_P2_U4101, new_P2_U4102, new_P2_U4103, new_P2_U4104,
    new_P2_U4105, new_P2_U4106, new_P2_U4107, new_P2_U4108, new_P2_U4109,
    new_P2_U4110, new_P2_U4111, new_P2_U4112, new_P2_U4113, new_P2_U4114,
    new_P2_U4115, new_P2_U4116, new_P2_U4117, new_P2_U4118, new_P2_U4119,
    new_P2_U4120, new_P2_U4121, new_P2_U4122, new_P2_U4123, new_P2_U4124,
    new_P2_U4125, new_P2_U4126, new_P2_U4127, new_P2_U4128, new_P2_U4129,
    new_P2_U4130, new_P2_U4131, new_P2_U4132, new_P2_U4133, new_P2_U4134,
    new_P2_U4135, new_P2_U4136, new_P2_U4137, new_P2_U4138, new_P2_U4139,
    new_P2_U4140, new_P2_U4141, new_P2_U4142, new_P2_U4143, new_P2_U4144,
    new_P2_U4145, new_P2_U4146, new_P2_U4147, new_P2_U4148, new_P2_U4149,
    new_P2_U4150, new_P2_U4151, new_P2_U4152, new_P2_U4153, new_P2_U4154,
    new_P2_U4155, new_P2_U4156, new_P2_U4157, new_P2_U4158, new_P2_U4159,
    new_P2_U4160, new_P2_U4161, new_P2_U4162, new_P2_U4163, new_P2_U4164,
    new_P2_U4165, new_P2_U4166, new_P2_U4167, new_P2_U4168, new_P2_U4169,
    new_P2_U4170, new_P2_U4171, new_P2_U4172, new_P2_U4173, new_P2_U4174,
    new_P2_U4175, new_P2_U4176, new_P2_U4177, new_P2_U4178, new_P2_U4179,
    new_P2_U4180, new_P2_U4181, new_P2_U4182, new_P2_U4183, new_P2_U4184,
    new_P2_U4185, new_P2_U4186, new_P2_U4187, new_P2_U4188, new_P2_U4189,
    new_P2_U4190, new_P2_U4191, new_P2_U4192, new_P2_U4193, new_P2_U4194,
    new_P2_U4195, new_P2_U4196, new_P2_U4197, new_P2_U4198, new_P2_U4199,
    new_P2_U4200, new_P2_U4201, new_P2_U4202, new_P2_U4203, new_P2_U4204,
    new_P2_U4205, new_P2_U4206, new_P2_U4207, new_P2_U4208, new_P2_U4209,
    new_P2_U4210, new_P2_U4211, new_P2_U4212, new_P2_U4213, new_P2_U4214,
    new_P2_U4215, new_P2_U4216, new_P2_U4217, new_P2_U4218, new_P2_U4219,
    new_P2_U4220, new_P2_U4221, new_P2_U4222, new_P2_U4223, new_P2_U4224,
    new_P2_U4225, new_P2_U4226, new_P2_U4227, new_P2_U4228, new_P2_U4229,
    new_P2_U4230, new_P2_U4231, new_P2_U4232, new_P2_U4233, new_P2_U4234,
    new_P2_U4235, new_P2_U4236, new_P2_U4237, new_P2_U4238, new_P2_U4239,
    new_P2_U4240, new_P2_U4241, new_P2_U4242, new_P2_U4243, new_P2_U4244,
    new_P2_U4245, new_P2_U4246, new_P2_U4247, new_P2_U4248, new_P2_U4249,
    new_P2_U4250, new_P2_U4251, new_P2_U4252, new_P2_U4253, new_P2_U4254,
    new_P2_U4255, new_P2_U4256, new_P2_U4257, new_P2_U4258, new_P2_U4259,
    new_P2_U4260, new_P2_U4261, new_P2_U4262, new_P2_U4263, new_P2_U4264,
    new_P2_U4265, new_P2_U4266, new_P2_U4267, new_P2_U4268, new_P2_U4269,
    new_P2_U4270, new_P2_U4271, new_P2_U4272, new_P2_U4273, new_P2_U4274,
    new_P2_U4275, new_P2_U4276, new_P2_U4277, new_P2_U4278, new_P2_U4279,
    new_P2_U4280, new_P2_U4281, new_P2_U4282, new_P2_U4283, new_P2_U4284,
    new_P2_U4285, new_P2_U4286, new_P2_U4287, new_P2_U4288, new_P2_U4289,
    new_P2_U4290, new_P2_U4291, new_P2_U4292, new_P2_U4293, new_P2_U4294,
    new_P2_U4295, new_P2_U4296, new_P2_U4297, new_P2_U4298, new_P2_U4299,
    new_P2_U4300, new_P2_U4301, new_P2_U4302, new_P2_U4303, new_P2_U4304,
    new_P2_U4305, new_P2_U4306, new_P2_U4307, new_P2_U4308, new_P2_U4309,
    new_P2_U4310, new_P2_U4311, new_P2_U4312, new_P2_U4313, new_P2_U4314,
    new_P2_U4315, new_P2_U4316, new_P2_U4317, new_P2_U4318, new_P2_U4319,
    new_P2_U4320, new_P2_U4321, new_P2_U4322, new_P2_U4323, new_P2_U4324,
    new_P2_U4325, new_P2_U4326, new_P2_U4327, new_P2_U4328, new_P2_U4329,
    new_P2_U4330, new_P2_U4331, new_P2_U4332, new_P2_U4333, new_P2_U4334,
    new_P2_U4335, new_P2_U4336, new_P2_U4337, new_P2_U4338, new_P2_U4339,
    new_P2_U4340, new_P2_U4341, new_P2_U4342, new_P2_U4343, new_P2_U4344,
    new_P2_U4345, new_P2_U4346, new_P2_U4347, new_P2_U4348, new_P2_U4349,
    new_P2_U4350, new_P2_U4351, new_P2_U4352, new_P2_U4353, new_P2_U4354,
    new_P2_U4355, new_P2_U4356, new_P2_U4357, new_P2_U4358, new_P2_U4359,
    new_P2_U4360, new_P2_U4361, new_P2_U4362, new_P2_U4363, new_P2_U4364,
    new_P2_U4365, new_P2_U4366, new_P2_U4367, new_P2_U4368, new_P2_U4369,
    new_P2_U4370, new_P2_U4371, new_P2_U4372, new_P2_U4373, new_P2_U4374,
    new_P2_U4375, new_P2_U4376, new_P2_U4377, new_P2_U4378, new_P2_U4379,
    new_P2_U4380, new_P2_U4381, new_P2_U4382, new_P2_U4383, new_P2_U4384,
    new_P2_U4385, new_P2_U4386, new_P2_U4387, new_P2_U4388, new_P2_U4389,
    new_P2_U4390, new_P2_U4391, new_P2_U4392, new_P2_U4393, new_P2_U4394,
    new_P2_U4395, new_P2_U4396, new_P2_U4397, new_P2_U4398, new_P2_U4399,
    new_P2_U4400, new_P2_U4401, new_P2_U4402, new_P2_U4403, new_P2_U4404,
    new_P2_U4405, new_P2_U4406, new_P2_U4407, new_P2_U4408, new_P2_U4409,
    new_P2_U4410, new_P2_U4411, new_P2_U4412, new_P2_U4413, new_P2_U4414,
    new_P2_U4415, new_P2_U4416, new_P2_U4417, new_P2_U4418, new_P2_U4419,
    new_P2_U4420, new_P2_U4421, new_P2_U4422, new_P2_U4423, new_P2_U4424,
    new_P2_U4425, new_P2_U4426, new_P2_U4427, new_P2_U4428, new_P2_U4429,
    new_P2_U4430, new_P2_U4431, new_P2_U4432, new_P2_U4433, new_P2_U4434,
    new_P2_U4435, new_P2_U4436, new_P2_U4437, new_P2_U4438, new_P2_U4439,
    new_P2_U4440, new_P2_U4441, new_P2_U4442, new_P2_U4443, new_P2_U4444,
    new_P2_U4445, new_P2_U4446, new_P2_U4447, new_P2_U4448, new_P2_U4449,
    new_P2_U4450, new_P2_U4451, new_P2_U4452, new_P2_U4453, new_P2_U4454,
    new_P2_U4455, new_P2_U4456, new_P2_U4457, new_P2_U4458, new_P2_U4459,
    new_P2_U4460, new_P2_U4461, new_P2_U4462, new_P2_U4463, new_P2_U4464,
    new_P2_U4465, new_P2_U4466, new_P2_U4467, new_P2_U4468, new_P2_U4469,
    new_P2_U4470, new_P2_U4471, new_P2_U4472, new_P2_U4473, new_P2_U4474,
    new_P2_U4475, new_P2_U4476, new_P2_U4477, new_P2_U4478, new_P2_U4479,
    new_P2_U4480, new_P2_U4481, new_P2_U4482, new_P2_U4483, new_P2_U4484,
    new_P2_U4485, new_P2_U4486, new_P2_U4487, new_P2_U4488, new_P2_U4489,
    new_P2_U4490, new_P2_U4491, new_P2_U4492, new_P2_U4493, new_P2_U4494,
    new_P2_U4495, new_P2_U4496, new_P2_U4497, new_P2_U4498, new_P2_U4499,
    new_P2_U4500, new_P2_U4501, new_P2_U4502, new_P2_U4503, new_P2_U4504,
    new_P2_U4505, new_P2_U4506, new_P2_U4507, new_P2_U4508, new_P2_U4509,
    new_P2_U4510, new_P2_U4511, new_P2_U4512, new_P2_U4513, new_P2_U4514,
    new_P2_U4515, new_P2_U4516, new_P2_U4517, new_P2_U4518, new_P2_U4519,
    new_P2_U4520, new_P2_U4521, new_P2_U4522, new_P2_U4523, new_P2_U4524,
    new_P2_U4525, new_P2_U4526, new_P2_U4527, new_P2_U4528, new_P2_U4529,
    new_P2_U4530, new_P2_U4531, new_P2_U4532, new_P2_U4533, new_P2_U4534,
    new_P2_U4535, new_P2_U4536, new_P2_U4537, new_P2_U4538, new_P2_U4539,
    new_P2_U4540, new_P2_U4541, new_P2_U4542, new_P2_U4543, new_P2_U4544,
    new_P2_U4545, new_P2_U4546, new_P2_U4547, new_P2_U4548, new_P2_U4549,
    new_P2_U4550, new_P2_U4551, new_P2_U4552, new_P2_U4553, new_P2_U4554,
    new_P2_U4555, new_P2_U4556, new_P2_U4557, new_P2_U4558, new_P2_U4559,
    new_P2_U4560, new_P2_U4561, new_P2_U4562, new_P2_U4563, new_P2_U4564,
    new_P2_U4565, new_P2_U4566, new_P2_U4567, new_P2_U4568, new_P2_U4569,
    new_P2_U4570, new_P2_U4571, new_P2_U4572, new_P2_U4573, new_P2_U4574,
    new_P2_U4575, new_P2_U4576, new_P2_U4577, new_P2_U4578, new_P2_U4579,
    new_P2_U4580, new_P2_U4581, new_P2_U4582, new_P2_U4583, new_P2_U4584,
    new_P2_U4585, new_P2_U4586, new_P2_U4587, new_P2_U4588, new_P2_U4589,
    new_P2_U4590, new_P2_U4591, new_P2_U4592, new_P2_U4593, new_P2_U4594,
    new_P2_U4595, new_P2_U4596, new_P2_U4597, new_P2_U4598, new_P2_U4599,
    new_P2_U4600, new_P2_U4601, new_P2_U4602, new_P2_U4603, new_P2_U4604,
    new_P2_U4605, new_P2_U4606, new_P2_U4607, new_P2_U4608, new_P2_U4609,
    new_P2_U4610, new_P2_U4611, new_P2_U4612, new_P2_U4613, new_P2_U4614,
    new_P2_U4615, new_P2_U4616, new_P2_U4617, new_P2_U4618, new_P2_U4619,
    new_P2_U4620, new_P2_U4621, new_P2_U4622, new_P2_U4623, new_P2_U4624,
    new_P2_U4625, new_P2_U4626, new_P2_U4627, new_P2_U4628, new_P2_U4629,
    new_P2_U4630, new_P2_U4631, new_P2_U4632, new_P2_U4633, new_P2_U4634,
    new_P2_U4635, new_P2_U4636, new_P2_U4637, new_P2_U4638, new_P2_U4639,
    new_P2_U4640, new_P2_U4641, new_P2_U4642, new_P2_U4643, new_P2_U4644,
    new_P2_U4645, new_P2_U4646, new_P2_U4647, new_P2_U4648, new_P2_U4649,
    new_P2_U4650, new_P2_U4651, new_P2_U4652, new_P2_U4653, new_P2_U4654,
    new_P2_U4655, new_P2_U4656, new_P2_U4657, new_P2_U4658, new_P2_U4659,
    new_P2_U4660, new_P2_U4661, new_P2_U4662, new_P2_U4663, new_P2_U4664,
    new_P2_U4665, new_P2_U4666, new_P2_U4667, new_P2_U4668, new_P2_U4669,
    new_P2_U4670, new_P2_U4671, new_P2_U4672, new_P2_U4673, new_P2_U4674,
    new_P2_U4675, new_P2_U4676, new_P2_U4677, new_P2_U4678, new_P2_U4679,
    new_P2_U4680, new_P2_U4681, new_P2_U4682, new_P2_U4683, new_P2_U4684,
    new_P2_U4685, new_P2_U4686, new_P2_U4687, new_P2_U4688, new_P2_U4689,
    new_P2_U4690, new_P2_U4691, new_P2_U4692, new_P2_U4693, new_P2_U4694,
    new_P2_U4695, new_P2_U4696, new_P2_U4697, new_P2_U4698, new_P2_U4699,
    new_P2_U4700, new_P2_U4701, new_P2_U4702, new_P2_U4703, new_P2_U4704,
    new_P2_U4705, new_P2_U4706, new_P2_U4707, new_P2_U4708, new_P2_U4709,
    new_P2_U4710, new_P2_U4711, new_P2_U4712, new_P2_U4713, new_P2_U4714,
    new_P2_U4715, new_P2_U4716, new_P2_U4717, new_P2_U4718, new_P2_U4719,
    new_P2_U4720, new_P2_U4721, new_P2_U4722, new_P2_U4723, new_P2_U4724,
    new_P2_U4725, new_P2_U4726, new_P2_U4727, new_P2_U4728, new_P2_U4729,
    new_P2_U4730, new_P2_U4731, new_P2_U4732, new_P2_U4733, new_P2_U4734,
    new_P2_U4735, new_P2_U4736, new_P2_U4737, new_P2_U4738, new_P2_U4739,
    new_P2_U4740, new_P2_U4741, new_P2_U4742, new_P2_U4743, new_P2_U4744,
    new_P2_U4745, new_P2_U4746, new_P2_U4747, new_P2_U4748, new_P2_U4749,
    new_P2_U4750, new_P2_U4751, new_P2_U4752, new_P2_U4753, new_P2_U4754,
    new_P2_U4755, new_P2_U4756, new_P2_U4757, new_P2_U4758, new_P2_U4759,
    new_P2_U4760, new_P2_U4761, new_P2_U4762, new_P2_U4763, new_P2_U4764,
    new_P2_U4765, new_P2_U4766, new_P2_U4767, new_P2_U4768, new_P2_U4769,
    new_P2_U4770, new_P2_U4771, new_P2_U4772, new_P2_U4773, new_P2_U4774,
    new_P2_U4775, new_P2_U4776, new_P2_U4777, new_P2_U4778, new_P2_U4779,
    new_P2_U4780, new_P2_U4781, new_P2_U4782, new_P2_U4783, new_P2_U4784,
    new_P2_U4785, new_P2_U4786, new_P2_U4787, new_P2_U4788, new_P2_U4789,
    new_P2_U4790, new_P2_U4791, new_P2_U4792, new_P2_U4793, new_P2_U4794,
    new_P2_U4795, new_P2_U4796, new_P2_U4797, new_P2_U4798, new_P2_U4799,
    new_P2_U4800, new_P2_U4801, new_P2_U4802, new_P2_U4803, new_P2_U4804,
    new_P2_U4805, new_P2_U4806, new_P2_U4807, new_P2_U4808, new_P2_U4809,
    new_P2_U4810, new_P2_U4811, new_P2_U4812, new_P2_U4813, new_P2_U4814,
    new_P2_U4815, new_P2_U4816, new_P2_U4817, new_P2_U4818, new_P2_U4819,
    new_P2_U4820, new_P2_U4821, new_P2_U4822, new_P2_U4823, new_P2_U4824,
    new_P2_U4825, new_P2_U4826, new_P2_U4827, new_P2_U4828, new_P2_U4829,
    new_P2_U4830, new_P2_U4831, new_P2_U4832, new_P2_U4833, new_P2_U4834,
    new_P2_U4835, new_P2_U4836, new_P2_U4837, new_P2_U4838, new_P2_U4839,
    new_P2_U4840, new_P2_U4841, new_P2_U4842, new_P2_U4843, new_P2_U4844,
    new_P2_U4845, new_P2_U4846, new_P2_U4847, new_P2_U4848, new_P2_U4849,
    new_P2_U4850, new_P2_U4851, new_P2_U4852, new_P2_U4853, new_P2_U4854,
    new_P2_U4855, new_P2_U4856, new_P2_U4857, new_P2_U4858, new_P2_U4859,
    new_P2_U4860, new_P2_U4861, new_P2_U4862, new_P2_U4863, new_P2_U4864,
    new_P2_U4865, new_P2_U4866, new_P2_U4867, new_P2_U4868, new_P2_U4869,
    new_P2_U4870, new_P2_U4871, new_P2_U4872, new_P2_U4873, new_P2_U4874,
    new_P2_U4875, new_P2_U4876, new_P2_U4877, new_P2_U4878, new_P2_U4879,
    new_P2_U4880, new_P2_U4881, new_P2_U4882, new_P2_U4883, new_P2_U4884,
    new_P2_U4885, new_P2_U4886, new_P2_U4887, new_P2_U4888, new_P2_U4889,
    new_P2_U4890, new_P2_U4891, new_P2_U4892, new_P2_U4893, new_P2_U4894,
    new_P2_U4895, new_P2_U4896, new_P2_U4897, new_P2_U4898, new_P2_U4899,
    new_P2_U4900, new_P2_U4901, new_P2_U4902, new_P2_U4903, new_P2_U4904,
    new_P2_U4905, new_P2_U4906, new_P2_U4907, new_P2_U4908, new_P2_U4909,
    new_P2_U4910, new_P2_U4911, new_P2_U4912, new_P2_U4913, new_P2_U4914,
    new_P2_U4915, new_P2_U4916, new_P2_U4917, new_P2_U4918, new_P2_U4919,
    new_P2_U4920, new_P2_U4921, new_P2_U4922, new_P2_U4923, new_P2_U4924,
    new_P2_U4925, new_P2_U4926, new_P2_U4927, new_P2_U4928, new_P2_U4929,
    new_P2_U4930, new_P2_U4931, new_P2_U4932, new_P2_U4933, new_P2_U4934,
    new_P2_U4935, new_P2_U4936, new_P2_U4937, new_P2_U4938, new_P2_U4939,
    new_P2_U4940, new_P2_U4941, new_P2_U4942, new_P2_U4943, new_P2_U4944,
    new_P2_U4945, new_P2_U4946, new_P2_U4947, new_P2_U4948, new_P2_U4949,
    new_P2_U4950, new_P2_U4951, new_P2_U4952, new_P2_U4953, new_P2_U4954,
    new_P2_U4955, new_P2_U4956, new_P2_U4957, new_P2_U4958, new_P2_U4959,
    new_P2_U4960, new_P2_U4961, new_P2_U4962, new_P2_U4963, new_P2_U4964,
    new_P2_U4965, new_P2_U4966, new_P2_U4967, new_P2_U4968, new_P2_U4969,
    new_P2_U4970, new_P2_U4971, new_P2_U4972, new_P2_U4973, new_P2_U4974,
    new_P2_U4975, new_P2_U4976, new_P2_U4977, new_P2_U4978, new_P2_U4979,
    new_P2_U4980, new_P2_U4981, new_P2_U4982, new_P2_U4983, new_P2_U4984,
    new_P2_U4985, new_P2_U4986, new_P2_U4987, new_P2_U4988, new_P2_U4989,
    new_P2_U4990, new_P2_U4991, new_P2_U4992, new_P2_U4993, new_P2_U4994,
    new_P2_U4995, new_P2_U4996, new_P2_U4997, new_P2_U4998, new_P2_U4999,
    new_P2_U5000, new_P2_U5001, new_P2_U5002, new_P2_U5003, new_P2_U5004,
    new_P2_U5005, new_P2_U5006, new_P2_U5007, new_P2_U5008, new_P2_U5009,
    new_P2_U5010, new_P2_U5011, new_P2_U5012, new_P2_U5013, new_P2_U5014,
    new_P2_U5015, new_P2_U5016, new_P2_U5017, new_P2_U5018, new_P2_U5019,
    new_P2_U5020, new_P2_U5021, new_P2_U5022, new_P2_U5023, new_P2_U5024,
    new_P2_U5025, new_P2_U5026, new_P2_U5027, new_P2_U5028, new_P2_U5029,
    new_P2_U5030, new_P2_U5031, new_P2_U5032, new_P2_U5033, new_P2_U5034,
    new_P2_U5035, new_P2_U5036, new_P2_U5037, new_P2_U5038, new_P2_U5039,
    new_P2_U5040, new_P2_U5041, new_P2_U5042, new_P2_U5043, new_P2_U5044,
    new_P2_U5045, new_P2_U5046, new_P2_U5047, new_P2_U5048, new_P2_U5049,
    new_P2_U5050, new_P2_U5051, new_P2_U5052, new_P2_U5053, new_P2_U5054,
    new_P2_U5055, new_P2_U5056, new_P2_U5057, new_P2_U5058, new_P2_U5059,
    new_P2_U5060, new_P2_U5061, new_P2_U5062, new_P2_U5063, new_P2_U5064,
    new_P2_U5065, new_P2_U5066, new_P2_U5067, new_P2_U5068, new_P2_U5069,
    new_P2_U5070, new_P2_U5071, new_P2_U5072, new_P2_U5073, new_P2_U5074,
    new_P2_U5075, new_P2_U5076, new_P2_U5077, new_P2_U5078, new_P2_U5079,
    new_P2_U5080, new_P2_U5081, new_P2_U5082, new_P2_U5083, new_P2_U5084,
    new_P2_U5085, new_P2_U5086, new_P2_U5087, new_P2_U5088, new_P2_U5089,
    new_P2_U5090, new_P2_U5091, new_P2_U5092, new_P2_U5093, new_P2_U5094,
    new_P2_U5095, new_P2_U5096, new_P2_U5097, new_P2_U5098, new_P2_U5099,
    new_P2_U5100, new_P2_U5101, new_P2_U5102, new_P2_U5103, new_P2_U5104,
    new_P2_U5105, new_P2_U5106, new_P2_U5107, new_P2_U5108, new_P2_U5109,
    new_P2_U5110, new_P2_U5111, new_P2_U5112, new_P2_U5113, new_P2_U5114,
    new_P2_U5115, new_P2_U5116, new_P2_U5117, new_P2_U5118, new_P2_U5119,
    new_P2_U5120, new_P2_U5121, new_P2_U5122, new_P2_U5123, new_P2_U5124,
    new_P2_U5125, new_P2_U5126, new_P2_U5127, new_P2_U5128, new_P2_U5129,
    new_P2_U5130, new_P2_U5131, new_P2_U5132, new_P2_U5133, new_P2_U5134,
    new_P2_U5135, new_P2_U5136, new_P2_U5137, new_P2_U5138, new_P2_U5139,
    new_P2_U5140, new_P2_U5141, new_P2_U5142, new_P2_U5143, new_P2_U5144,
    new_P2_U5145, new_P2_U5146, new_P2_U5147, new_P2_U5148, new_P2_U5149,
    new_P2_U5150, new_P2_U5151, new_P2_U5152, new_P2_U5153, new_P2_U5154,
    new_P2_U5155, new_P2_U5156, new_P2_U5157, new_P2_U5158, new_P2_U5159,
    new_P2_U5160, new_P2_U5161, new_P2_U5162, new_P2_U5163, new_P2_U5164,
    new_P2_U5165, new_P2_U5166, new_P2_U5167, new_P2_U5168, new_P2_U5169,
    new_P2_U5170, new_P2_U5171, new_P2_U5172, new_P2_U5173, new_P2_U5174,
    new_P2_U5175, new_P2_U5176, new_P2_U5177, new_P2_U5178, new_P2_U5179,
    new_P2_U5180, new_P2_U5181, new_P2_U5182, new_P2_U5183, new_P2_U5184,
    new_P2_U5185, new_P2_U5186, new_P2_U5187, new_P2_U5188, new_P2_U5189,
    new_P2_U5190, new_P2_U5191, new_P2_U5192, new_P2_U5193, new_P2_U5194,
    new_P2_U5195, new_P2_U5196, new_P2_U5197, new_P2_U5198, new_P2_U5199,
    new_P2_U5200, new_P2_U5201, new_P2_U5202, new_P2_U5203, new_P2_U5204,
    new_P2_U5205, new_P2_U5206, new_P2_U5207, new_P2_U5208, new_P2_U5209,
    new_P2_U5210, new_P2_U5211, new_P2_U5212, new_P2_U5213, new_P2_U5214,
    new_P2_U5215, new_P2_U5216, new_P2_U5217, new_P2_U5218, new_P2_U5219,
    new_P2_U5220, new_P2_U5221, new_P2_U5222, new_P2_U5223, new_P2_U5224,
    new_P2_U5225, new_P2_U5226, new_P2_U5227, new_P2_U5228, new_P2_U5229,
    new_P2_U5230, new_P2_U5231, new_P2_U5232, new_P2_U5233, new_P2_U5234,
    new_P2_U5235, new_P2_U5236, new_P2_U5237, new_P2_U5238, new_P2_U5239,
    new_P2_U5240, new_P2_U5241, new_P2_U5242, new_P2_U5243, new_P2_U5244,
    new_P2_U5245, new_P2_U5246, new_P2_U5247, new_P2_U5248, new_P2_U5249,
    new_P2_U5250, new_P2_U5251, new_P2_U5252, new_P2_U5253, new_P2_U5254,
    new_P2_U5255, new_P2_U5256, new_P2_U5257, new_P2_U5258, new_P2_U5259,
    new_P2_U5260, new_P2_U5261, new_P2_U5262, new_P2_U5263, new_P2_U5264,
    new_P2_U5265, new_P2_U5266, new_P2_U5267, new_P2_U5268, new_P2_U5269,
    new_P2_U5270, new_P2_U5271, new_P2_U5272, new_P2_U5273, new_P2_U5274,
    new_P2_U5275, new_P2_U5276, new_P2_U5277, new_P2_U5278, new_P2_U5279,
    new_P2_U5280, new_P2_U5281, new_P2_U5282, new_P2_U5283, new_P2_U5284,
    new_P2_U5285, new_P2_U5286, new_P2_U5287, new_P2_U5288, new_P2_U5289,
    new_P2_U5290, new_P2_U5291, new_P2_U5292, new_P2_U5293, new_P2_U5294,
    new_P2_U5295, new_P2_U5296, new_P2_U5297, new_P2_U5298, new_P2_U5299,
    new_P2_U5300, new_P2_U5301, new_P2_U5302, new_P2_U5303, new_P2_U5304,
    new_P2_U5305, new_P2_U5306, new_P2_U5307, new_P2_U5308, new_P2_U5309,
    new_P2_U5310, new_P2_U5311, new_P2_U5312, new_P2_U5313, new_P2_U5314,
    new_P2_U5315, new_P2_U5316, new_P2_U5317, new_P2_U5318, new_P2_U5319,
    new_P2_U5320, new_P2_U5321, new_P2_U5322, new_P2_U5323, new_P2_U5324,
    new_P2_U5325, new_P2_U5326, new_P2_U5327, new_P2_U5328, new_P2_U5329,
    new_P2_U5330, new_P2_U5331, new_P2_U5332, new_P2_U5333, new_P2_U5334,
    new_P2_U5335, new_P2_U5336, new_P2_U5337, new_P2_U5338, new_P2_U5339,
    new_P2_U5340, new_P2_U5341, new_P2_U5342, new_P2_U5343, new_P2_U5344,
    new_P2_U5345, new_P2_U5346, new_P2_U5347, new_P2_U5348, new_P2_U5349,
    new_P2_U5350, new_P2_U5351, new_P2_U5352, new_P2_U5353, new_P2_U5354,
    new_P2_U5355, new_P2_U5356, new_P2_U5357, new_P2_U5358, new_P2_U5359,
    new_P2_U5360, new_P2_U5361, new_P2_U5362, new_P2_U5363, new_P2_U5364,
    new_P2_U5365, new_P2_U5366, new_P2_U5367, new_P2_U5368, new_P2_U5369,
    new_P2_U5370, new_P2_U5371, new_P2_U5372, new_P2_U5373, new_P2_U5374,
    new_P2_U5375, new_P2_U5376, new_P2_U5377, new_P2_U5378, new_P2_U5379,
    new_P2_U5380, new_P2_U5381, new_P2_U5382, new_P2_U5383, new_P2_U5384,
    new_P2_U5385, new_P2_U5386, new_P2_U5387, new_P2_U5388, new_P2_U5389,
    new_P2_U5390, new_P2_U5391, new_P2_U5392, new_P2_U5393, new_P2_U5394,
    new_P2_U5395, new_P2_U5396, new_P2_U5397, new_P2_U5398, new_P2_U5399,
    new_P2_U5400, new_P2_U5401, new_P2_U5402, new_P2_U5403, new_P2_U5404,
    new_P2_U5405, new_P2_U5406, new_P2_U5407, new_P2_U5408, new_P2_U5409,
    new_P2_U5410, new_P2_U5411, new_P2_U5412, new_P2_U5413, new_P2_U5414,
    new_P2_U5415, new_P2_U5416, new_P2_U5417, new_P2_U5418, new_P2_U5419,
    new_P2_U5420, new_P2_U5421, new_P2_U5422, new_P2_U5423, new_P2_U5424,
    new_P2_U5425, new_P2_U5426, new_P2_U5427, new_P2_U5428, new_P2_U5429,
    new_P2_U5430, new_P2_U5431, new_P2_U5432, new_P2_U5433, new_P2_U5434,
    new_P2_U5435, new_P2_U5436, new_P2_U5437, new_P2_U5438, new_P2_U5439,
    new_P2_U5440, new_P2_U5441, new_P2_U5442, new_P2_U5443, new_P2_U5444,
    new_P2_U5445, new_P2_U5446, new_P2_U5447, new_P2_U5448, new_P2_U5449,
    new_P2_U5450, new_P2_U5451, new_P2_U5452, new_P2_U5453, new_P2_U5454,
    new_P2_U5455, new_P2_U5456, new_P2_U5457, new_P2_U5458, new_P2_U5459,
    new_P2_U5460, new_P2_U5461, new_P2_U5462, new_P2_U5463, new_P2_U5464,
    new_P2_U5465, new_P2_U5466, new_P2_U5467, new_P2_U5468, new_P2_U5469,
    new_P2_U5470, new_P2_U5471, new_P2_U5472, new_P2_U5473, new_P2_U5474,
    new_P2_U5475, new_P2_U5476, new_P2_U5477, new_P2_U5478, new_P2_U5479,
    new_P2_U5480, new_P2_U5481, new_P2_U5482, new_P2_U5483, new_P2_U5484,
    new_P2_U5485, new_P2_U5486, new_P2_U5487, new_P2_U5488, new_P2_U5489,
    new_P2_U5490, new_P2_U5491, new_P2_U5492, new_P2_U5493, new_P2_U5494,
    new_P2_U5495, new_P2_U5496, new_P2_U5497, new_P2_U5498, new_P2_U5499,
    new_P2_U5500, new_P2_U5501, new_P2_U5502, new_P2_U5503, new_P2_U5504,
    new_P2_U5505, new_P2_U5506, new_P2_U5507, new_P2_U5508, new_P2_U5509,
    new_P2_U5510, new_P2_U5511, new_P2_U5512, new_P2_U5513, new_P2_U5514,
    new_P2_U5515, new_P2_U5516, new_P2_U5517, new_P2_U5518, new_P2_U5519,
    new_P2_U5520, new_P2_U5521, new_P2_U5522, new_P2_U5523, new_P2_U5524,
    new_P2_U5525, new_P2_U5526, new_P2_U5527, new_P2_U5528, new_P2_U5529,
    new_P2_U5530, new_P2_U5531, new_P2_U5532, new_P2_U5533, new_P2_U5534,
    new_P2_U5535, new_P2_U5536, new_P2_U5537, new_P2_U5538, new_P2_U5539,
    new_P2_U5540, new_P2_U5541, new_P2_U5542, new_P2_U5543, new_P2_U5544,
    new_P2_U5545, new_P2_U5546, new_P2_U5547, new_P2_U5548, new_P2_U5549,
    new_P2_U5550, new_P2_U5551, new_P2_U5552, new_P2_U5553, new_P2_U5554,
    new_P2_U5555, new_P2_U5556, new_P2_U5557, new_P2_U5558, new_P2_U5559,
    new_P2_U5560, new_P2_U5561, new_P2_U5562, new_P2_U5563, new_P2_U5564,
    new_P2_U5565, new_P2_U5566, new_P2_U5567, new_P2_U5568, new_P2_U5569,
    new_P2_U5570, new_P2_U5571, new_P2_U5572, new_P2_U5573, new_P2_U5574,
    new_P2_U5575, new_P2_U5576, new_P2_U5577, new_P2_U5578, new_P2_U5579,
    new_P2_U5580, new_P2_U5581, new_P2_U5582, new_P2_U5583, new_P2_U5584,
    new_P2_U5585, new_P2_U5586, new_P2_U5587, new_P2_U5588, new_P2_U5589,
    new_P2_U5590, new_P2_U5591, new_P2_U5592, new_P2_U5593, new_P2_U5594,
    new_P2_U5595, new_P2_U5596, new_P2_U5597, new_P2_U5598, new_P2_U5599,
    new_P2_U5600, new_P2_U5601, new_P2_U5602, new_P2_U5603, new_P2_U5604,
    new_P2_U5605, new_P2_U5606, new_P2_U5607, new_P2_U5608, new_P2_U5609,
    new_P2_U5610, new_P2_U5611, new_P2_U5612, new_P2_U5613, new_P2_U5614,
    new_P2_U5615, new_P2_U5616, new_P2_U5617, new_P2_U5618, new_P2_U5619,
    new_P2_U5620, new_P2_U5621, new_P2_U5622, new_P2_U5623, new_P2_U5624,
    new_P2_U5625, new_P2_U5626, new_P2_U5627, new_P2_U5628, new_P2_U5629,
    new_P2_U5630, new_P2_U5631, new_P2_U5632, new_P2_U5633, new_P2_U5634,
    new_P2_U5635, new_P2_U5636, new_P2_U5637, new_P2_U5638, new_P2_U5639,
    new_P2_U5640, new_P2_U5641, new_P2_U5642, new_P2_U5643, new_P2_U5644,
    new_P2_U5645, new_P2_U5646, new_P2_U5647, new_P2_U5648, new_P2_U5649,
    new_P2_U5650, new_P2_U5651, new_P2_U5652, new_P2_U5653, new_P2_U5654,
    new_P2_U5655, new_P2_U5656, new_P2_U5657, new_P2_U5658, new_P2_U5659,
    new_P2_U5660, new_P2_U5661, new_P2_U5662, new_P2_U5663, new_P2_U5664,
    new_P2_U5665, new_P2_U5666, new_P2_U5667, new_P2_U5668, new_P2_U5669,
    new_P2_U5670, new_P2_U5671, new_P2_U5672, new_P2_U5673, new_P2_U5674,
    new_P2_U5675, new_P2_U5676, new_P2_U5677, new_P2_U5678, new_P2_U5679,
    new_P2_U5680, new_P2_U5681, new_P2_U5682, new_P2_U5683, new_P2_U5684,
    new_P2_U5685, new_P2_U5686, new_P2_U5687, new_P2_U5688, new_P2_U5689,
    new_P2_U5690, new_P2_U5691, new_P2_U5692, new_P2_U5693, new_P2_U5694,
    new_P2_U5695, new_P2_U5696, new_P2_U5697, new_P2_U5698, new_P2_U5699,
    new_P2_U5700, new_P2_U5701, new_P2_U5702, new_P2_U5703, new_P2_U5704,
    new_P2_U5705, new_P2_U5706, new_P2_U5707, new_P2_U5708, new_P2_U5709,
    new_P2_U5710, new_P2_U5711, new_P2_U5712, new_P2_U5713, new_P2_U5714,
    new_P2_U5715, new_P2_U5716, new_P2_U5717, new_P2_U5718, new_P2_U5719,
    new_P2_U5720, new_P2_U5721, new_P2_U5722, new_P2_U5723, new_P2_U5724,
    new_P2_U5725, new_P2_U5726, new_P2_U5727, new_P2_U5728, new_P2_U5729,
    new_P2_U5730, new_P2_U5731, new_P2_U5732, new_P2_U5733, new_P2_U5734,
    new_P2_U5735, new_P2_U5736, new_P2_U5737, new_P2_U5738, new_P2_U5739,
    new_P2_U5740, new_P2_U5741, new_P2_U5742, new_P2_U5743, new_P2_U5744,
    new_P2_U5745, new_P2_U5746, new_P2_U5747, new_P2_U5748, new_P2_U5749,
    new_P2_U5750, new_P2_U5751, new_P2_U5752, new_P2_U5753, new_P2_U5754,
    new_P2_U5755, new_P2_U5756, new_P2_U5757, new_P2_U5758, new_P2_U5759,
    new_P2_U5760, new_P2_U5761, new_P2_U5762, new_P2_U5763, new_P2_U5764,
    new_P2_U5765, new_P2_U5766, new_P2_U5767, new_P2_U5768, new_P2_U5769,
    new_P2_U5770, new_P2_U5771, new_P2_U5772, new_P2_U5773, new_P2_U5774,
    new_P2_U5775, new_P2_U5776, new_P2_U5777, new_P2_U5778, new_P2_U5779,
    new_P2_U5780, new_P2_U5781, new_P2_U5782, new_P2_U5783, new_P2_U5784,
    new_P2_U5785, new_P2_U5786, new_P2_U5787, new_P2_U5788, new_P2_U5789,
    new_P2_U5790, new_P2_U5791, new_P2_U5792, new_P2_U5793, new_P2_U5794,
    new_P2_U5795, new_P2_U5796, new_P2_U5797, new_P2_U5798, new_P2_U5799,
    new_P2_U5800, new_P2_U5801, new_P2_U5802, new_P2_U5803, new_P2_U5804,
    new_P2_U5805, new_P2_U5806, new_P2_U5807, new_P2_U5808, new_P2_U5809,
    new_P2_U5810, new_P2_U5811, new_P2_U5812, new_P2_U5813, new_P2_U5814,
    new_P2_U5815, new_P2_U5816, new_P2_U5817, new_P2_U5818, new_P2_U5819,
    new_P2_U5820, new_P2_U5821, new_P2_U5822, new_P2_U5823, new_P2_U5824,
    new_P2_U5825, new_P2_U5826, new_P2_U5827, new_P2_U5828, new_P2_U5829,
    new_P2_U5830, new_P2_U5831, new_P2_U5832, new_P2_U5833, new_P2_U5834,
    new_P2_U5835, new_P2_U5836, new_P2_U5837, new_P2_U5838, new_P2_U5839,
    new_P2_U5840, new_P2_U5841, new_P2_U5842, new_P2_U5843, new_P2_U5844,
    new_P2_U5845, new_P2_U5846, new_P2_U5847, new_P2_U5848, new_P2_U5849,
    new_P2_U5850, new_P2_U5851, new_P2_U5852, new_P2_U5853, new_P2_U5854,
    new_P2_U5855, new_P2_U5856, new_P2_U5857, new_P2_U5858, new_P2_U5859,
    new_P2_U5860, new_P2_U5861, new_P2_U5862, new_P2_U5863, new_P2_U5864,
    new_P2_U5865, new_P2_U5866, new_P2_U5867, new_P2_U5868, new_P2_U5869,
    new_P2_U5870, new_P2_U5871, new_P2_U5872, new_P2_U5873, new_P2_U5874,
    new_P2_U5875, new_P2_U5876, new_P2_U5877, new_P2_U5878, new_P2_U5879,
    new_P2_U5880, new_P2_U5881, new_P2_U5882, new_P2_U5883, new_P2_U5884,
    new_P2_U5885, new_P2_U5886, new_P2_U5887, new_P2_U5888, new_P2_U5889,
    new_P2_U5890, new_P2_U5891, new_P2_U5892, new_P2_U5893, new_P2_U5894,
    new_P2_U5895, new_P2_U5896, new_P2_U5897, new_P2_U5898, new_P2_U5899,
    new_P2_U5900, new_P2_U5901, new_P2_U5902, new_P2_U5903, new_P2_U5904,
    new_P2_U5905, new_P2_U5906, new_P2_U5907, new_P2_U5908, new_P2_U5909,
    new_P2_U5910, new_P2_U5911, new_P2_U5912, new_P2_U5913, new_P2_U5914,
    new_P2_U5915, new_P2_U5916, new_P2_U5917, new_P2_U5918, new_P2_U5919,
    new_P2_U5920, new_P2_U5921, new_P2_U5922, new_P2_U5923, new_P2_U5924,
    new_P2_U5925, new_P2_U5926, new_P2_U5927, new_P2_U5928, new_P2_U5929,
    new_P2_U5930, new_P2_U5931, new_P2_U5932, new_P2_U5933, new_P2_U5934,
    new_P2_U5935, new_P2_U5936, new_P2_U5937, new_P2_U5938, new_P2_U5939,
    new_P2_U5940, new_P2_U5941, new_P2_U5942, new_P2_U5943, new_P2_U5944,
    new_P2_U5945, new_P2_U5946, new_P2_U5947, new_P2_U5948, new_P2_U5949,
    new_P2_U5950, new_P2_U5951, new_P2_U5952, new_P2_U5953, new_P2_U5954,
    new_P2_U5955, new_P2_U5956, new_P2_U5957, new_P2_U5958, new_P2_U5959,
    new_P2_U5960, new_P2_U5961, new_P2_U5962, new_P2_U5963, new_P2_U5964,
    new_P2_U5965, new_P2_U5966, new_P2_U5967, new_P2_U5968, new_P2_U5969,
    new_P2_U5970, new_P2_U5971, new_P2_U5972, new_P2_U5973, new_P2_U5974,
    new_P2_U5975, new_P2_U5976, new_P2_U5977, new_P2_U5978, new_P2_U5979,
    new_P2_U5980, new_P2_U5981, new_P2_U5982, new_P2_U5983, new_P2_U5984,
    new_P2_U5985, new_P2_U5986, new_P2_U5987, new_P2_U5988, new_P2_U5989,
    new_P2_U5990, new_P2_U5991, new_P2_U5992, new_P2_U5993, new_P2_U5994,
    new_P2_U5995, new_P2_U5996, new_P2_U5997, new_P2_U5998, new_P2_U5999,
    new_P2_U6000, new_P2_U6001, new_P2_U6002, new_P2_U6003, new_P2_U6004,
    new_P2_U6005, new_P2_U6006, new_P2_U6007, new_P2_U6008, new_P2_U6009,
    new_P2_U6010, new_P2_U6011, new_P2_U6012, new_P2_U6013, new_P2_U6014,
    new_P2_U6015, new_P2_U6016, new_P2_U6017, new_P2_U6018, new_P2_U6019,
    new_P2_U6020, new_P2_U6021, new_P2_U6022, new_P2_U6023, new_P2_U6024,
    new_P2_U6025, new_P2_U6026, new_P2_U6027, new_P2_U6028, new_P2_U6029,
    new_P2_U6030, new_P2_U6031, new_P2_U6032, new_P2_U6033, new_P2_U6034,
    new_P2_U6035, new_P2_U6036, new_P2_U6037, new_P2_U6038, new_P2_U6039,
    new_P2_U6040, new_P2_U6041, new_P2_U6042, new_P2_U6043, new_P2_U6044,
    new_P2_U6045, new_P2_U6046, new_P2_U6047, new_P2_U6048, new_P2_U6049,
    new_P2_U6050, new_P2_U6051, new_P2_U6052, new_P2_U6053, new_P2_U6054,
    new_P2_U6055, new_P2_U6056, new_P2_U6057, new_P2_U6058, new_P2_U6059,
    new_P2_U6060, new_P2_U6061, new_P2_U6062, new_P2_U6063, new_P2_U6064,
    new_P2_U6065, new_P2_U6066, new_P2_U6067, new_P2_U6068, new_P2_U6069,
    new_P2_U6070, new_P2_U6071, new_P2_U6072, new_P2_U6073, new_P2_U6074,
    new_P2_U6075, new_P2_U6076, new_P2_U6077, new_P2_U6078, new_P2_U6079,
    new_P2_U6080, new_P2_U6081, new_P2_U6082, new_P2_U6083, new_P2_U6084,
    new_P2_U6085, new_P2_U6086, new_P2_U6087, new_P2_U6088, new_P2_U6089,
    new_P2_U6090, new_P2_U6091, new_P2_U6092, new_P2_U6093, new_P2_U6094,
    new_P2_U6095, new_P2_U6096, new_P2_U6097, new_P2_U6098, new_P2_U6099,
    new_P2_U6100, new_P2_U6101, new_P2_U6102, new_P2_U6103, new_P2_U6104,
    new_P2_U6105, new_P2_U6106, new_P2_U6107, new_P2_U6108, new_P2_U6109,
    new_P2_U6110, new_P2_U6111, new_P2_U6112, new_P2_U6113, new_P2_U6114,
    new_P2_U6115, new_P2_U6116, new_P2_U6117, new_P2_U6118, new_P2_U6119,
    new_P2_U6120, new_P2_U6121, new_P2_U6122, new_P2_U6123, new_P2_U6124,
    new_P2_U6125, new_P2_U6126, new_P2_U6127, new_P2_U6128, new_P2_U6129,
    new_P2_U6130, new_P2_U6131, new_P2_U6132, new_P2_U6133, new_P2_U6134,
    new_P2_U6135, new_P2_U6136, new_P2_U6137, new_P2_U6138, new_P2_U6139,
    new_P2_U6140, new_P2_U6141, new_P2_U6142, new_P2_U6143, new_P2_U6144,
    new_P2_U6145, new_P2_U6146, new_P2_U6147, new_P2_U6148, new_P2_U6149,
    new_P2_U6150, new_P3_R1161_U468, new_P3_R1161_U467, new_P3_R1161_U466,
    new_P3_R1161_U465, new_P3_R1161_U464, new_P3_R1161_U463,
    new_P3_R1161_U462, new_P3_R1161_U461, new_P3_R1161_U460,
    new_P3_R1161_U459, new_P3_R1161_U458, new_P3_R1161_U457,
    new_P3_R1161_U456, new_P3_R1161_U455, new_P3_R1161_U454,
    new_P3_R1161_U453, new_P3_R1161_U452, new_P3_R1161_U451,
    new_P3_R1161_U450, new_P3_R1161_U449, new_P3_U3013, new_P3_U3014,
    new_P3_U3015, new_P3_U3016, new_P3_U3017, new_P3_U3018, new_P3_U3019,
    new_P3_U3020, new_P3_U3021, new_P3_U3022, new_P3_U3023, new_P3_U3024,
    new_P3_U3025, new_P3_U3026, new_P3_U3027, new_P3_U3028, new_P3_U3029,
    new_P3_U3030, new_P3_U3031, new_P3_U3032, new_P3_U3033, new_P3_U3034,
    new_P3_U3035, new_P3_U3036, new_P3_U3037, new_P3_U3038, new_P3_U3039,
    new_P3_U3040, new_P3_U3041, new_P3_U3042, new_P3_U3043, new_P3_U3044,
    new_P3_U3045, new_P3_U3046, new_P3_U3047, new_P3_U3048, new_P3_U3049,
    new_P3_U3050, new_P3_U3051, new_P3_U3052, new_P3_U3053, new_P3_U3054,
    new_P3_U3055, new_P3_U3056, new_P3_U3057, new_P3_U3058, new_P3_U3059,
    new_P3_U3060, new_P3_U3061, new_P3_U3062, new_P3_U3063, new_P3_U3064,
    new_P3_U3065, new_P3_U3066, new_P3_U3067, new_P3_U3068, new_P3_U3069,
    new_P3_U3070, new_P3_U3071, new_P3_U3072, new_P3_U3073, new_P3_U3074,
    new_P3_U3075, new_P3_U3076, new_P3_U3077, new_P3_U3078, new_P3_U3079,
    new_P3_U3080, new_P3_U3081, new_P3_U3082, new_P3_U3083, new_P3_U3084,
    new_P3_U3085, new_P3_U3086, new_P3_U3087, new_P3_U3088, new_P3_U3089,
    new_P3_U3090, new_P3_U3091, new_P3_U3092, new_P3_U3093, new_P3_U3094,
    new_P3_U3095, new_P3_U3096, new_P3_U3097, new_P3_U3098, new_P3_U3099,
    new_P3_U3100, new_P3_U3101, new_P3_U3102, new_P3_U3103, new_P3_U3104,
    new_P3_U3105, new_P3_U3106, new_P3_U3107, new_P3_U3108, new_P3_U3109,
    new_P3_U3110, new_P3_U3111, new_P3_U3112, new_P3_U3113, new_P3_U3114,
    new_P3_U3115, new_P3_U3116, new_P3_U3117, new_P3_U3118, new_P3_U3119,
    new_P3_U3120, new_P3_U3121, new_P3_U3122, new_P3_U3123, new_P3_U3124,
    new_P3_U3125, new_P3_U3126, new_P3_U3127, new_P3_U3128, new_P3_U3129,
    new_P3_U3130, new_P3_U3131, new_P3_U3132, new_P3_U3133, new_P3_U3134,
    new_P3_U3135, new_P3_U3136, new_P3_U3137, new_P3_U3138, new_P3_U3139,
    new_P3_U3140, new_P3_U3141, new_P3_U3142, new_P3_U3143, new_P3_U3144,
    new_P3_U3145, new_P3_U3146, new_P3_U3147, new_P3_U3148, new_P3_U3149,
    new_P3_U3152, new_P3_U3297, new_P3_U3298, new_P3_U3299, new_P3_U3300,
    new_P3_U3301, new_P3_U3302, new_P3_U3303, new_P3_U3304, new_P3_U3305,
    new_P3_U3306, new_P3_U3307, new_P3_U3308, new_P3_U3309, new_P3_U3310,
    new_P3_U3311, new_P3_U3312, new_P3_U3313, new_P3_U3314, new_P3_U3315,
    new_P3_U3316, new_P3_U3317, new_P3_U3318, new_P3_U3319, new_P3_U3320,
    new_P3_U3321, new_P3_U3322, new_P3_U3323, new_P3_U3324, new_P3_U3325,
    new_P3_U3326, new_P3_U3327, new_P3_U3328, new_P3_U3329, new_P3_U3330,
    new_P3_U3331, new_P3_U3332, new_P3_U3333, new_P3_U3334, new_P3_U3335,
    new_P3_U3336, new_P3_U3337, new_P3_U3338, new_P3_U3339, new_P3_U3340,
    new_P3_U3341, new_P3_U3342, new_P3_U3343, new_P3_U3344, new_P3_U3345,
    new_P3_U3346, new_P3_U3347, new_P3_U3348, new_P3_U3349, new_P3_U3350,
    new_P3_U3351, new_P3_U3352, new_P3_U3353, new_P3_U3354, new_P3_U3355,
    new_P3_U3356, new_P3_U3357, new_P3_U3358, new_P3_U3359, new_P3_U3360,
    new_P3_U3361, new_P3_U3362, new_P3_U3363, new_P3_U3364, new_P3_U3365,
    new_P3_U3366, new_P3_U3367, new_P3_U3368, new_P3_U3369, new_P3_U3370,
    new_P3_U3371, new_P3_U3372, new_P3_U3373, new_P3_U3374, new_P3_U3375,
    new_P3_U3378, new_P3_U3379, new_P3_U3380, new_P3_U3381, new_P3_U3382,
    new_P3_U3383, new_P3_U3384, new_P3_U3385, new_P3_U3386, new_P3_U3387,
    new_P3_U3388, new_P3_U3389, new_P3_U3391, new_P3_U3392, new_P3_U3394,
    new_P3_U3395, new_P3_U3397, new_P3_U3398, new_P3_U3400, new_P3_U3401,
    new_P3_U3403, new_P3_U3404, new_P3_U3406, new_P3_U3407, new_P3_U3409,
    new_P3_U3410, new_P3_U3412, new_P3_U3413, new_P3_U3415, new_P3_U3416,
    new_P3_U3418, new_P3_U3419, new_P3_U3421, new_P3_U3422, new_P3_U3424,
    new_P3_U3425, new_P3_U3427, new_P3_U3428, new_P3_U3430, new_P3_U3431,
    new_P3_U3433, new_P3_U3434, new_P3_U3436, new_P3_U3437, new_P3_U3439,
    new_P3_U3440, new_P3_U3442, new_P3_U3443, new_P3_U3445, new_P3_U3523,
    new_P3_U3524, new_P3_U3525, new_P3_U3526, new_P3_U3527, new_P3_U3528,
    new_P3_U3529, new_P3_U3530, new_P3_U3531, new_P3_U3532, new_P3_U3533,
    new_P3_U3534, new_P3_U3535, new_P3_U3536, new_P3_U3537, new_P3_U3538,
    new_P3_U3539, new_P3_U3540, new_P3_U3541, new_P3_U3542, new_P3_U3543,
    new_P3_U3544, new_P3_U3545, new_P3_U3546, new_P3_U3547, new_P3_U3548,
    new_P3_U3549, new_P3_U3550, new_P3_U3551, new_P3_U3552, new_P3_U3553,
    new_P3_U3554, new_P3_U3555, new_P3_U3556, new_P3_U3557, new_P3_U3558,
    new_P3_U3559, new_P3_U3560, new_P3_U3561, new_P3_U3562, new_P3_U3563,
    new_P3_U3564, new_P3_U3565, new_P3_U3566, new_P3_U3567, new_P3_U3568,
    new_P3_U3569, new_P3_U3570, new_P3_U3571, new_P3_U3572, new_P3_U3573,
    new_P3_U3574, new_P3_U3575, new_P3_U3576, new_P3_U3577, new_P3_U3578,
    new_P3_U3579, new_P3_U3580, new_P3_U3581, new_P3_U3582, new_P3_U3583,
    new_P3_U3584, new_P3_U3585, new_P3_U3586, new_P3_U3587, new_P3_U3588,
    new_P3_U3589, new_P3_U3590, new_P3_U3591, new_P3_U3592, new_P3_U3593,
    new_P3_U3594, new_P3_U3595, new_P3_U3596, new_P3_U3597, new_P3_U3598,
    new_P3_U3599, new_P3_U3600, new_P3_U3601, new_P3_U3602, new_P3_U3603,
    new_P3_U3604, new_P3_U3605, new_P3_U3606, new_P3_U3607, new_P3_U3608,
    new_P3_U3609, new_P3_U3610, new_P3_U3611, new_P3_U3612, new_P3_U3613,
    new_P3_U3614, new_P3_U3615, new_P3_U3616, new_P3_U3617, new_P3_U3618,
    new_P3_U3619, new_P3_U3620, new_P3_U3621, new_P3_U3622, new_P3_U3623,
    new_P3_U3624, new_P3_U3625, new_P3_U3626, new_P3_U3627, new_P3_U3628,
    new_P3_U3629, new_P3_U3630, new_P3_U3631, new_P3_U3632, new_P3_U3633,
    new_P3_U3634, new_P3_U3635, new_P3_U3636, new_P3_U3637, new_P3_U3638,
    new_P3_U3639, new_P3_U3640, new_P3_U3641, new_P3_U3642, new_P3_U3643,
    new_P3_U3644, new_P3_U3645, new_P3_U3646, new_P3_U3647, new_P3_U3648,
    new_P3_U3649, new_P3_U3650, new_P3_U3651, new_P3_U3652, new_P3_U3653,
    new_P3_U3654, new_P3_U3655, new_P3_U3656, new_P3_U3657, new_P3_U3658,
    new_P3_U3659, new_P3_U3660, new_P3_U3661, new_P3_U3662, new_P3_U3663,
    new_P3_U3664, new_P3_U3665, new_P3_U3666, new_P3_U3667, new_P3_U3668,
    new_P3_U3669, new_P3_U3670, new_P3_U3671, new_P3_U3672, new_P3_U3673,
    new_P3_U3674, new_P3_U3675, new_P3_U3676, new_P3_U3677, new_P3_U3678,
    new_P3_U3679, new_P3_U3680, new_P3_U3681, new_P3_U3682, new_P3_U3683,
    new_P3_U3684, new_P3_U3685, new_P3_U3686, new_P3_U3687, new_P3_U3688,
    new_P3_U3689, new_P3_U3690, new_P3_U3691, new_P3_U3692, new_P3_U3693,
    new_P3_U3694, new_P3_U3695, new_P3_U3696, new_P3_U3697, new_P3_U3698,
    new_P3_U3699, new_P3_U3700, new_P3_U3701, new_P3_U3702, new_P3_U3703,
    new_P3_U3704, new_P3_U3705, new_P3_U3706, new_P3_U3707, new_P3_U3708,
    new_P3_U3709, new_P3_U3710, new_P3_U3711, new_P3_U3712, new_P3_U3713,
    new_P3_U3714, new_P3_U3715, new_P3_U3716, new_P3_U3717, new_P3_U3718,
    new_P3_U3719, new_P3_U3720, new_P3_U3721, new_P3_U3722, new_P3_U3723,
    new_P3_U3724, new_P3_U3725, new_P3_U3726, new_P3_U3727, new_P3_U3728,
    new_P3_U3729, new_P3_U3730, new_P3_U3731, new_P3_U3732, new_P3_U3733,
    new_P3_U3734, new_P3_U3735, new_P3_U3736, new_P3_U3737, new_P3_U3738,
    new_P3_U3739, new_P3_U3740, new_P3_U3741, new_P3_U3742, new_P3_U3743,
    new_P3_U3744, new_P3_U3745, new_P3_U3746, new_P3_U3747, new_P3_U3748,
    new_P3_U3749, new_P3_U3750, new_P3_U3751, new_P3_U3752, new_P3_U3753,
    new_P3_U3754, new_P3_U3755, new_P3_U3756, new_P3_U3757, new_P3_U3758,
    new_P3_U3759, new_P3_U3760, new_P3_U3761, new_P3_U3762, new_P3_U3763,
    new_P3_U3764, new_P3_U3765, new_P3_U3766, new_P3_U3767, new_P3_U3768,
    new_P3_U3769, new_P3_U3770, new_P3_U3771, new_P3_U3772, new_P3_U3773,
    new_P3_U3774, new_P3_U3775, new_P3_U3776, new_P3_U3777, new_P3_U3778,
    new_P3_U3779, new_P3_U3780, new_P3_U3781, new_P3_U3782, new_P3_U3783,
    new_P3_U3784, new_P3_U3785, new_P3_U3786, new_P3_U3787, new_P3_U3788,
    new_P3_U3789, new_P3_U3790, new_P3_U3791, new_P3_U3792, new_P3_U3793,
    new_P3_U3794, new_P3_U3795, new_P3_U3796, new_P3_U3797, new_P3_U3798,
    new_P3_U3799, new_P3_U3800, new_P3_U3801, new_P3_U3802, new_P3_U3803,
    new_P3_U3804, new_P3_U3805, new_P3_U3806, new_P3_U3807, new_P3_U3808,
    new_P3_U3809, new_P3_U3810, new_P3_U3811, new_P3_U3812, new_P3_U3813,
    new_P3_U3814, new_P3_U3815, new_P3_U3816, new_P3_U3817, new_P3_U3818,
    new_P3_U3819, new_P3_U3820, new_P3_U3821, new_P3_U3822, new_P3_U3823,
    new_P3_U3824, new_P3_U3825, new_P3_U3826, new_P3_U3827, new_P3_U3828,
    new_P3_U3829, new_P3_U3830, new_P3_U3831, new_P3_U3832, new_P3_U3833,
    new_P3_U3834, new_P3_U3835, new_P3_U3836, new_P3_U3837, new_P3_U3838,
    new_P3_U3839, new_P3_U3840, new_P3_U3841, new_P3_U3842, new_P3_U3843,
    new_P3_U3844, new_P3_U3845, new_P3_U3846, new_P3_U3847, new_P3_U3848,
    new_P3_U3849, new_P3_U3850, new_P3_U3851, new_P3_U3852, new_P3_U3853,
    new_P3_U3854, new_P3_U3855, new_P3_U3856, new_P3_U3857, new_P3_U3858,
    new_P3_U3859, new_P3_U3860, new_P3_U3861, new_P3_U3862, new_P3_U3863,
    new_P3_U3864, new_P3_U3865, new_P3_U3866, new_P3_U3867, new_P3_U3868,
    new_P3_U3869, new_P3_U3870, new_P3_U3871, new_P3_U3872, new_P3_U3873,
    new_P3_U3874, new_P3_U3875, new_P3_U3876, new_P3_U3877, new_P3_U3878,
    new_P3_U3879, new_P3_U3880, new_P3_U3881, new_P3_U3882, new_P3_U3883,
    new_P3_U3884, new_P3_U3885, new_P3_U3886, new_P3_U3887, new_P3_U3888,
    new_P3_U3889, new_P3_U3890, new_P3_U3891, new_P3_U3892, new_P3_U3893,
    new_P3_U3894, new_P3_U3895, new_P3_U3896, new_P3_U3898, new_P3_U3899,
    new_P3_U3900, new_P3_U3901, new_P3_U3902, new_P3_U3903, new_P3_U3904,
    new_P3_U3905, new_P3_U3906, new_P3_U3907, new_P3_U3908, new_P3_U3909,
    new_P3_U3910, new_P3_U3911, new_P3_U3912, new_P3_U3913, new_P3_U3914,
    new_P3_U3915, new_P3_U3916, new_P3_U3917, new_P3_U3918, new_P3_U3919,
    new_P3_U3920, new_P3_U3921, new_P3_U3922, new_P3_U3923, new_P3_U3924,
    new_P3_U3925, new_P3_U3926, new_P3_U3927, new_P3_U3928, new_P3_U3929,
    new_P3_U3930, new_P3_U3931, new_P3_U3932, new_P3_U3933, new_P3_U3934,
    new_P3_U3935, new_P3_U3936, new_P3_U3937, new_P3_U3938, new_P3_U3939,
    new_P3_U3940, new_P3_U3941, new_P3_U3942, new_P3_U3943, new_P3_U3944,
    new_P3_U3945, new_P3_U3946, new_P3_U3947, new_P3_U3948, new_P3_U3949,
    new_P3_U3950, new_P3_U3951, new_P3_U3952, new_P3_U3953, new_P3_U3954,
    new_P3_U3955, new_P3_U3956, new_P3_U3957, new_P3_U3958, new_P3_U3959,
    new_P3_U3960, new_P3_U3961, new_P3_U3962, new_P3_U3963, new_P3_U3964,
    new_P3_U3965, new_P3_U3966, new_P3_U3967, new_P3_U3968, new_P3_U3969,
    new_P3_U3970, new_P3_U3971, new_P3_U3972, new_P3_U3973, new_P3_U3974,
    new_P3_U3975, new_P3_U3976, new_P3_U3977, new_P3_U3978, new_P3_U3979,
    new_P3_U3980, new_P3_U3981, new_P3_U3982, new_P3_U3983, new_P3_U3984,
    new_P3_U3985, new_P3_U3986, new_P3_U3987, new_P3_U3988, new_P3_U3989,
    new_P3_U3990, new_P3_U3991, new_P3_U3992, new_P3_U3993, new_P3_U3994,
    new_P3_U3995, new_P3_U3996, new_P3_U3997, new_P3_U3998, new_P3_U3999,
    new_P3_U4000, new_P3_U4001, new_P3_U4002, new_P3_U4003, new_P3_U4004,
    new_P3_U4005, new_P3_U4006, new_P3_U4007, new_P3_U4008, new_P3_U4009,
    new_P3_U4010, new_P3_U4011, new_P3_U4012, new_P3_U4013, new_P3_U4014,
    new_P3_U4015, new_P3_U4016, new_P3_U4017, new_P3_U4018, new_P3_U4019,
    new_P3_U4020, new_P3_U4021, new_P3_U4022, new_P3_U4023, new_P3_U4024,
    new_P3_U4025, new_P3_U4026, new_P3_U4027, new_P3_U4028, new_P3_U4029,
    new_P3_U4030, new_P3_U4031, new_P3_U4032, new_P3_U4033, new_P3_U4034,
    new_P3_U4035, new_P3_U4036, new_P3_U4037, new_P3_U4038, new_P3_U4039,
    new_P3_U4040, new_P3_U4041, new_P3_U4042, new_P3_U4043, new_P3_U4044,
    new_P3_U4045, new_P3_U4046, new_P3_U4047, new_P3_U4048, new_P3_U4049,
    new_P3_U4050, new_P3_U4051, new_P3_U4052, new_P3_U4053, new_P3_U4054,
    new_P3_U4055, new_P3_U4056, new_P3_U4057, new_P3_U4058, new_P3_U4059,
    new_P3_U4060, new_P3_U4061, new_P3_U4062, new_P3_U4063, new_P3_U4064,
    new_P3_U4065, new_P3_U4066, new_P3_U4067, new_P3_U4068, new_P3_U4069,
    new_P3_U4070, new_P3_U4071, new_P3_U4072, new_P3_U4073, new_P3_U4074,
    new_P3_U4075, new_P3_U4076, new_P3_U4077, new_P3_U4078, new_P3_U4079,
    new_P3_U4080, new_P3_U4081, new_P3_U4082, new_P3_U4083, new_P3_U4084,
    new_P3_U4085, new_P3_U4086, new_P3_U4087, new_P3_U4088, new_P3_U4089,
    new_P3_U4090, new_P3_U4091, new_P3_U4092, new_P3_U4093, new_P3_U4094,
    new_P3_U4095, new_P3_U4096, new_P3_U4097, new_P3_U4098, new_P3_U4099,
    new_P3_U4100, new_P3_U4101, new_P3_U4102, new_P3_U4103, new_P3_U4104,
    new_P3_U4105, new_P3_U4106, new_P3_U4107, new_P3_U4108, new_P3_U4109,
    new_P3_U4110, new_P3_U4111, new_P3_U4112, new_P3_U4113, new_P3_U4114,
    new_P3_U4115, new_P3_U4116, new_P3_U4117, new_P3_U4118, new_P3_U4119,
    new_P3_U4120, new_P3_U4121, new_P3_U4122, new_P3_U4123, new_P3_U4124,
    new_P3_U4125, new_P3_U4126, new_P3_U4127, new_P3_U4128, new_P3_U4129,
    new_P3_U4130, new_P3_U4131, new_P3_U4132, new_P3_U4133, new_P3_U4134,
    new_P3_U4135, new_P3_U4136, new_P3_U4137, new_P3_U4138, new_P3_U4139,
    new_P3_U4140, new_P3_U4141, new_P3_U4142, new_P3_U4143, new_P3_U4144,
    new_P3_U4145, new_P3_U4146, new_P3_U4147, new_P3_U4148, new_P3_U4149,
    new_P3_U4150, new_P3_U4151, new_P3_U4152, new_P3_U4153, new_P3_U4154,
    new_P3_U4155, new_P3_U4156, new_P3_U4157, new_P3_U4158, new_P3_U4159,
    new_P3_U4160, new_P3_U4161, new_P3_U4162, new_P3_U4163, new_P3_U4164,
    new_P3_U4165, new_P3_U4166, new_P3_U4167, new_P3_U4168, new_P3_U4169,
    new_P3_U4170, new_P3_U4171, new_P3_U4172, new_P3_U4173, new_P3_U4174,
    new_P3_U4175, new_P3_U4176, new_P3_U4177, new_P3_U4178, new_P3_U4179,
    new_P3_U4180, new_P3_U4181, new_P3_U4182, new_P3_U4183, new_P3_U4184,
    new_P3_U4185, new_P3_U4186, new_P3_U4187, new_P3_U4188, new_P3_U4189,
    new_P3_U4190, new_P3_U4191, new_P3_U4192, new_P3_U4193, new_P3_U4194,
    new_P3_U4195, new_P3_U4196, new_P3_U4197, new_P3_U4198, new_P3_U4199,
    new_P3_U4200, new_P3_U4201, new_P3_U4202, new_P3_U4203, new_P3_U4204,
    new_P3_U4205, new_P3_U4206, new_P3_U4207, new_P3_U4208, new_P3_U4209,
    new_P3_U4210, new_P3_U4211, new_P3_U4212, new_P3_U4213, new_P3_U4214,
    new_P3_U4215, new_P3_U4216, new_P3_U4217, new_P3_U4218, new_P3_U4219,
    new_P3_U4220, new_P3_U4221, new_P3_U4222, new_P3_U4223, new_P3_U4224,
    new_P3_U4225, new_P3_U4226, new_P3_U4227, new_P3_U4228, new_P3_U4229,
    new_P3_U4230, new_P3_U4231, new_P3_U4232, new_P3_U4233, new_P3_U4234,
    new_P3_U4235, new_P3_U4236, new_P3_U4237, new_P3_U4238, new_P3_U4239,
    new_P3_U4240, new_P3_U4241, new_P3_U4242, new_P3_U4243, new_P3_U4244,
    new_P3_U4245, new_P3_U4246, new_P3_U4247, new_P3_U4248, new_P3_U4249,
    new_P3_U4250, new_P3_U4251, new_P3_U4252, new_P3_U4253, new_P3_U4254,
    new_P3_U4255, new_P3_U4256, new_P3_U4257, new_P3_U4258, new_P3_U4259,
    new_P3_U4260, new_P3_U4261, new_P3_U4262, new_P3_U4263, new_P3_U4264,
    new_P3_U4265, new_P3_U4266, new_P3_U4267, new_P3_U4268, new_P3_U4269,
    new_P3_U4270, new_P3_U4271, new_P3_U4272, new_P3_U4273, new_P3_U4274,
    new_P3_U4275, new_P3_U4276, new_P3_U4277, new_P3_U4278, new_P3_U4279,
    new_P3_U4280, new_P3_U4281, new_P3_U4282, new_P3_U4283, new_P3_U4284,
    new_P3_U4285, new_P3_U4286, new_P3_U4287, new_P3_U4288, new_P3_U4289,
    new_P3_U4290, new_P3_U4291, new_P3_U4292, new_P3_U4293, new_P3_U4294,
    new_P3_U4295, new_P3_U4296, new_P3_U4297, new_P3_U4298, new_P3_U4299,
    new_P3_U4300, new_P3_U4301, new_P3_U4302, new_P3_U4303, new_P3_U4304,
    new_P3_U4305, new_P3_U4306, new_P3_U4307, new_P3_U4308, new_P3_U4309,
    new_P3_U4310, new_P3_U4311, new_P3_U4312, new_P3_U4313, new_P3_U4314,
    new_P3_U4315, new_P3_U4316, new_P3_U4317, new_P3_U4318, new_P3_U4319,
    new_P3_U4320, new_P3_U4321, new_P3_U4322, new_P3_U4323, new_P3_U4324,
    new_P3_U4325, new_P3_U4326, new_P3_U4327, new_P3_U4328, new_P3_U4329,
    new_P3_U4330, new_P3_U4331, new_P3_U4332, new_P3_U4333, new_P3_U4334,
    new_P3_U4335, new_P3_U4336, new_P3_U4337, new_P3_U4338, new_P3_U4339,
    new_P3_U4340, new_P3_U4341, new_P3_U4342, new_P3_U4343, new_P3_U4344,
    new_P3_U4345, new_P3_U4346, new_P3_U4347, new_P3_U4348, new_P3_U4349,
    new_P3_U4350, new_P3_U4351, new_P3_U4352, new_P3_U4353, new_P3_U4354,
    new_P3_U4355, new_P3_U4356, new_P3_U4357, new_P3_U4358, new_P3_U4359,
    new_P3_U4360, new_P3_U4361, new_P3_U4362, new_P3_U4363, new_P3_U4364,
    new_P3_U4365, new_P3_U4366, new_P3_U4367, new_P3_U4368, new_P3_U4369,
    new_P3_U4370, new_P3_U4371, new_P3_U4372, new_P3_U4373, new_P3_U4374,
    new_P3_U4375, new_P3_U4376, new_P3_U4377, new_P3_U4378, new_P3_U4379,
    new_P3_U4380, new_P3_U4381, new_P3_U4382, new_P3_U4383, new_P3_U4384,
    new_P3_U4385, new_P3_U4386, new_P3_U4387, new_P3_U4388, new_P3_U4389,
    new_P3_U4390, new_P3_U4391, new_P3_U4392, new_P3_U4393, new_P3_U4394,
    new_P3_U4395, new_P3_U4396, new_P3_U4397, new_P3_U4398, new_P3_U4399,
    new_P3_U4400, new_P3_U4401, new_P3_U4402, new_P3_U4403, new_P3_U4404,
    new_P3_U4405, new_P3_U4406, new_P3_U4407, new_P3_U4408, new_P3_U4409,
    new_P3_U4410, new_P3_U4411, new_P3_U4412, new_P3_U4413, new_P3_U4414,
    new_P3_U4415, new_P3_U4416, new_P3_U4417, new_P3_U4418, new_P3_U4419,
    new_P3_U4420, new_P3_U4421, new_P3_U4422, new_P3_U4423, new_P3_U4424,
    new_P3_U4425, new_P3_U4426, new_P3_U4427, new_P3_U4428, new_P3_U4429,
    new_P3_U4430, new_P3_U4431, new_P3_U4432, new_P3_U4433, new_P3_U4434,
    new_P3_U4435, new_P3_U4436, new_P3_U4437, new_P3_U4438, new_P3_U4439,
    new_P3_U4440, new_P3_U4441, new_P3_U4442, new_P3_U4443, new_P3_U4444,
    new_P3_U4445, new_P3_U4446, new_P3_U4447, new_P3_U4448, new_P3_U4449,
    new_P3_U4450, new_P3_U4451, new_P3_U4452, new_P3_U4453, new_P3_U4454,
    new_P3_U4455, new_P3_U4456, new_P3_U4457, new_P3_U4458, new_P3_U4459,
    new_P3_U4460, new_P3_U4461, new_P3_U4462, new_P3_U4463, new_P3_U4464,
    new_P3_U4465, new_P3_U4466, new_P3_U4467, new_P3_U4468, new_P3_U4469,
    new_P3_U4470, new_P3_U4471, new_P3_U4472, new_P3_U4473, new_P3_U4474,
    new_P3_U4475, new_P3_U4476, new_P3_U4477, new_P3_U4478, new_P3_U4479,
    new_P3_U4480, new_P3_U4481, new_P3_U4482, new_P3_U4483, new_P3_U4484,
    new_P3_U4485, new_P3_U4486, new_P3_U4487, new_P3_U4488, new_P3_U4489,
    new_P3_U4490, new_P3_U4491, new_P3_U4492, new_P3_U4493, new_P3_U4494,
    new_P3_U4495, new_P3_U4496, new_P3_U4497, new_P3_U4498, new_P3_U4499,
    new_P3_U4500, new_P3_U4501, new_P3_U4502, new_P3_U4503, new_P3_U4504,
    new_P3_U4505, new_P3_U4506, new_P3_U4507, new_P3_U4508, new_P3_U4509,
    new_P3_U4510, new_P3_U4511, new_P3_U4512, new_P3_U4513, new_P3_U4514,
    new_P3_U4515, new_P3_U4516, new_P3_U4517, new_P3_U4518, new_P3_U4519,
    new_P3_U4520, new_P3_U4521, new_P3_U4522, new_P3_U4523, new_P3_U4524,
    new_P3_U4525, new_P3_U4526, new_P3_U4527, new_P3_U4528, new_P3_U4529,
    new_P3_U4530, new_P3_U4531, new_P3_U4532, new_P3_U4533, new_P3_U4534,
    new_P3_U4535, new_P3_U4536, new_P3_U4537, new_P3_U4538, new_P3_U4539,
    new_P3_U4540, new_P3_U4541, new_P3_U4542, new_P3_U4543, new_P3_U4544,
    new_P3_U4545, new_P3_U4546, new_P3_U4547, new_P3_U4548, new_P3_U4549,
    new_P3_U4550, new_P3_U4551, new_P3_U4552, new_P3_U4553, new_P3_U4554,
    new_P3_U4555, new_P3_U4556, new_P3_U4557, new_P3_U4558, new_P3_U4559,
    new_P3_U4560, new_P3_U4561, new_P3_U4562, new_P3_U4563, new_P3_U4564,
    new_P3_U4565, new_P3_U4566, new_P3_U4567, new_P3_U4568, new_P3_U4569,
    new_P3_U4570, new_P3_U4571, new_P3_U4572, new_P3_U4573, new_P3_U4574,
    new_P3_U4575, new_P3_U4576, new_P3_U4577, new_P3_U4578, new_P3_U4579,
    new_P3_U4580, new_P3_U4581, new_P3_U4582, new_P3_U4583, new_P3_U4584,
    new_P3_U4585, new_P3_U4586, new_P3_U4587, new_P3_U4588, new_P3_U4589,
    new_P3_U4590, new_P3_U4591, new_P3_U4592, new_P3_U4593, new_P3_U4594,
    new_P3_U4595, new_P3_U4596, new_P3_U4597, new_P3_U4598, new_P3_U4599,
    new_P3_U4600, new_P3_U4601, new_P3_U4602, new_P3_U4603, new_P3_U4604,
    new_P3_U4605, new_P3_U4606, new_P3_U4607, new_P3_U4608, new_P3_U4609,
    new_P3_U4610, new_P3_U4611, new_P3_U4612, new_P3_U4613, new_P3_U4614,
    new_P3_U4615, new_P3_U4616, new_P3_U4617, new_P3_U4618, new_P3_U4619,
    new_P3_U4620, new_P3_U4621, new_P3_U4622, new_P3_U4623, new_P3_U4624,
    new_P3_U4625, new_P3_U4626, new_P3_U4627, new_P3_U4628, new_P3_U4629,
    new_P3_U4630, new_P3_U4631, new_P3_U4632, new_P3_U4633, new_P3_U4634,
    new_P3_U4635, new_P3_U4636, new_P3_U4637, new_P3_U4638, new_P3_U4639,
    new_P3_U4640, new_P3_U4641, new_P3_U4642, new_P3_U4643, new_P3_U4644,
    new_P3_U4645, new_P3_U4646, new_P3_U4647, new_P3_U4648, new_P3_U4649,
    new_P3_U4650, new_P3_U4651, new_P3_U4652, new_P3_U4653, new_P3_U4654,
    new_P3_U4655, new_P3_U4656, new_P3_U4657, new_P3_U4658, new_P3_U4659,
    new_P3_U4660, new_P3_U4661, new_P3_U4662, new_P3_U4663, new_P3_U4664,
    new_P3_U4665, new_P3_U4666, new_P3_U4667, new_P3_U4668, new_P3_U4669,
    new_P3_U4670, new_P3_U4671, new_P3_U4672, new_P3_U4673, new_P3_U4674,
    new_P3_U4675, new_P3_U4676, new_P3_U4677, new_P3_U4678, new_P3_U4679,
    new_P3_U4680, new_P3_U4681, new_P3_U4682, new_P3_U4683, new_P3_U4684,
    new_P3_U4685, new_P3_U4686, new_P3_U4687, new_P3_U4688, new_P3_U4689,
    new_P3_U4690, new_P3_U4691, new_P3_U4692, new_P3_U4693, new_P3_U4694,
    new_P3_U4695, new_P3_U4696, new_P3_U4697, new_P3_U4698, new_P3_U4699,
    new_P3_U4700, new_P3_U4701, new_P3_U4702, new_P3_U4703, new_P3_U4704,
    new_P3_U4705, new_P3_U4706, new_P3_U4707, new_P3_U4708, new_P3_U4709,
    new_P3_U4710, new_P3_U4711, new_P3_U4712, new_P3_U4713, new_P3_U4714,
    new_P3_U4715, new_P3_U4716, new_P3_U4717, new_P3_U4718, new_P3_U4719,
    new_P3_U4720, new_P3_U4721, new_P3_U4722, new_P3_U4723, new_P3_U4724,
    new_P3_U4725, new_P3_U4726, new_P3_U4727, new_P3_U4728, new_P3_U4729,
    new_P3_U4730, new_P3_U4731, new_P3_U4732, new_P3_U4733, new_P3_U4734,
    new_P3_U4735, new_P3_U4736, new_P3_U4737, new_P3_U4738, new_P3_U4739,
    new_P3_U4740, new_P3_U4741, new_P3_U4742, new_P3_U4743, new_P3_U4744,
    new_P3_U4745, new_P3_U4746, new_P3_U4747, new_P3_U4748, new_P3_U4749,
    new_P3_U4750, new_P3_U4751, new_P3_U4752, new_P3_U4753, new_P3_U4754,
    new_P3_U4755, new_P3_U4756, new_P3_U4757, new_P3_U4758, new_P3_U4759,
    new_P3_U4760, new_P3_U4761, new_P3_U4762, new_P3_U4763, new_P3_U4764,
    new_P3_U4765, new_P3_U4766, new_P3_U4767, new_P3_U4768, new_P3_U4769,
    new_P3_U4770, new_P3_U4771, new_P3_U4772, new_P3_U4773, new_P3_U4774,
    new_P3_U4775, new_P3_U4776, new_P3_U4777, new_P3_U4778, new_P3_U4779,
    new_P3_U4780, new_P3_U4781, new_P3_U4782, new_P3_U4783, new_P3_U4784,
    new_P3_U4785, new_P3_U4786, new_P3_U4787, new_P3_U4788, new_P3_U4789,
    new_P3_U4790, new_P3_U4791, new_P3_U4792, new_P3_U4793, new_P3_U4794,
    new_P3_U4795, new_P3_U4796, new_P3_U4797, new_P3_U4798, new_P3_U4799,
    new_P3_U4800, new_P3_U4801, new_P3_U4802, new_P3_U4803, new_P3_U4804,
    new_P3_U4805, new_P3_U4806, new_P3_U4807, new_P3_U4808, new_P3_U4809,
    new_P3_U4810, new_P3_U4811, new_P3_U4812, new_P3_U4813, new_P3_U4814,
    new_P3_U4815, new_P3_U4816, new_P3_U4817, new_P3_U4818, new_P3_U4819,
    new_P3_U4820, new_P3_U4821, new_P3_U4822, new_P3_U4823, new_P3_U4824,
    new_P3_U4825, new_P3_U4826, new_P3_U4827, new_P3_U4828, new_P3_U4829,
    new_P3_U4830, new_P3_U4831, new_P3_U4832, new_P3_U4833, new_P3_U4834,
    new_P3_U4835, new_P3_U4836, new_P3_U4837, new_P3_U4838, new_P3_U4839,
    new_P3_U4840, new_P3_U4841, new_P3_U4842, new_P3_U4843, new_P3_U4844,
    new_P3_U4845, new_P3_U4846, new_P3_U4847, new_P3_U4848, new_P3_U4849,
    new_P3_U4850, new_P3_U4851, new_P3_U4852, new_P3_U4853, new_P3_U4854,
    new_P3_U4855, new_P3_U4856, new_P3_U4857, new_P3_U4858, new_P3_U4859,
    new_P3_U4860, new_P3_U4861, new_P3_U4862, new_P3_U4863, new_P3_U4864,
    new_P3_U4865, new_P3_U4866, new_P3_U4867, new_P3_U4868, new_P3_U4869,
    new_P3_U4870, new_P3_U4871, new_P3_U4872, new_P3_U4873, new_P3_U4874,
    new_P3_U4875, new_P3_U4876, new_P3_U4877, new_P3_U4878, new_P3_U4879,
    new_P3_U4880, new_P3_U4881, new_P3_U4882, new_P3_U4883, new_P3_U4884,
    new_P3_U4885, new_P3_U4886, new_P3_U4887, new_P3_U4888, new_P3_U4889,
    new_P3_U4890, new_P3_U4891, new_P3_U4892, new_P3_U4893, new_P3_U4894,
    new_P3_U4895, new_P3_U4896, new_P3_U4897, new_P3_U4898, new_P3_U4899,
    new_P3_U4900, new_P3_U4901, new_P3_U4902, new_P3_U4903, new_P3_U4904,
    new_P3_U4905, new_P3_U4906, new_P3_U4907, new_P3_U4908, new_P3_U4909,
    new_P3_U4910, new_P3_U4911, new_P3_U4912, new_P3_U4913, new_P3_U4914,
    new_P3_U4915, new_P3_U4916, new_P3_U4917, new_P3_U4918, new_P3_U4919,
    new_P3_U4920, new_P3_U4921, new_P3_U4922, new_P3_U4923, new_P3_U4924,
    new_P3_U4925, new_P3_U4926, new_P3_U4927, new_P3_U4928, new_P3_U4929,
    new_P3_U4930, new_P3_U4931, new_P3_U4932, new_P3_U4933, new_P3_U4934,
    new_P3_U4935, new_P3_U4936, new_P3_U4937, new_P3_U4938, new_P3_U4939,
    new_P3_U4940, new_P3_U4941, new_P3_U4942, new_P3_U4943, new_P3_U4944,
    new_P3_U4945, new_P3_U4946, new_P3_U4947, new_P3_U4948, new_P3_U4949,
    new_P3_U4950, new_P3_U4951, new_P3_U4952, new_P3_U4953, new_P3_U4954,
    new_P3_U4955, new_P3_U4956, new_P3_U4957, new_P3_U4958, new_P3_U4959,
    new_P3_U4960, new_P3_U4961, new_P3_U4962, new_P3_U4963, new_P3_U4964,
    new_P3_U4965, new_P3_U4966, new_P3_U4967, new_P3_U4968, new_P3_U4969,
    new_P3_U4970, new_P3_U4971, new_P3_U4972, new_P3_U4973, new_P3_U4974,
    new_P3_U4975, new_P3_U4976, new_P3_U4977, new_P3_U4978, new_P3_U4979,
    new_P3_U4980, new_P3_U4981, new_P3_U4982, new_P3_U4983, new_P3_U4984,
    new_P3_U4985, new_P3_U4986, new_P3_U4987, new_P3_U4988, new_P3_U4989,
    new_P3_U4990, new_P3_U4991, new_P3_U4992, new_P3_U4993, new_P3_U4994,
    new_P3_U4995, new_P3_U4996, new_P3_U4997, new_P3_U4998, new_P3_U4999,
    new_P3_U5000, new_P3_U5001, new_P3_U5002, new_P3_U5003, new_P3_U5004,
    new_P3_U5005, new_P3_U5006, new_P3_U5007, new_P3_U5008, new_P3_U5009,
    new_P3_U5010, new_P3_U5011, new_P3_U5012, new_P3_U5013, new_P3_U5014,
    new_P3_U5015, new_P3_U5016, new_P3_U5017, new_P3_U5018, new_P3_U5019,
    new_P3_U5020, new_P3_U5021, new_P3_U5022, new_P3_U5023, new_P3_U5024,
    new_P3_U5025, new_P3_U5026, new_P3_U5027, new_P3_U5028, new_P3_U5029,
    new_P3_U5030, new_P3_U5031, new_P3_U5032, new_P3_U5033, new_P3_U5034,
    new_P3_U5035, new_P3_U5036, new_P3_U5037, new_P3_U5038, new_P3_U5039,
    new_P3_U5040, new_P3_U5041, new_P3_U5042, new_P3_U5043, new_P3_U5044,
    new_P3_U5045, new_P3_U5046, new_P3_U5047, new_P3_U5048, new_P3_U5049,
    new_P3_U5050, new_P3_U5051, new_P3_U5052, new_P3_U5053, new_P3_U5054,
    new_P3_U5055, new_P3_U5056, new_P3_U5057, new_P3_U5058, new_P3_U5059,
    new_P3_U5060, new_P3_U5061, new_P3_U5062, new_P3_U5063, new_P3_U5064,
    new_P3_U5065, new_P3_U5066, new_P3_U5067, new_P3_U5068, new_P3_U5069,
    new_P3_U5070, new_P3_U5071, new_P3_U5072, new_P3_U5073, new_P3_U5074,
    new_P3_U5075, new_P3_U5076, new_P3_U5077, new_P3_U5078, new_P3_U5079,
    new_P3_U5080, new_P3_U5081, new_P3_U5082, new_P3_U5083, new_P3_U5084,
    new_P3_U5085, new_P3_U5086, new_P3_U5087, new_P3_U5088, new_P3_U5089,
    new_P3_U5090, new_P3_U5091, new_P3_U5092, new_P3_U5093, new_P3_U5094,
    new_P3_U5095, new_P3_U5096, new_P3_U5097, new_P3_U5098, new_P3_U5099,
    new_P3_U5100, new_P3_U5101, new_P3_U5102, new_P3_U5103, new_P3_U5104,
    new_P3_U5105, new_P3_U5106, new_P3_U5107, new_P3_U5108, new_P3_U5109,
    new_P3_U5110, new_P3_U5111, new_P3_U5112, new_P3_U5113, new_P3_U5114,
    new_P3_U5115, new_P3_U5116, new_P3_U5117, new_P3_U5118, new_P3_U5119,
    new_P3_U5120, new_P3_U5121, new_P3_U5122, new_P3_U5123, new_P3_U5124,
    new_P3_U5125, new_P3_U5126, new_P3_U5127, new_P3_U5128, new_P3_U5129,
    new_P3_U5130, new_P3_U5131, new_P3_U5132, new_P3_U5133, new_P3_U5134,
    new_P3_U5135, new_P3_U5136, new_P3_U5137, new_P3_U5138, new_P3_U5139,
    new_P3_U5140, new_P3_U5141, new_P3_U5142, new_P3_U5143, new_P3_U5144,
    new_P3_U5145, new_P3_U5146, new_P3_U5147, new_P3_U5148, new_P3_U5149,
    new_P3_U5150, new_P3_U5151, new_P3_U5152, new_P3_U5153, new_P3_U5154,
    new_P3_U5155, new_P3_U5156, new_P3_U5157, new_P3_U5158, new_P3_U5159,
    new_P3_U5160, new_P3_U5161, new_P3_U5162, new_P3_U5163, new_P3_U5164,
    new_P3_U5165, new_P3_U5166, new_P3_U5167, new_P3_U5168, new_P3_U5169,
    new_P3_U5170, new_P3_U5171, new_P3_U5172, new_P3_U5173, new_P3_U5174,
    new_P3_U5175, new_P3_U5176, new_P3_U5177, new_P3_U5178, new_P3_U5179,
    new_P3_U5180, new_P3_U5181, new_P3_U5182, new_P3_U5183, new_P3_U5184,
    new_P3_U5185, new_P3_U5186, new_P3_U5187, new_P3_U5188, new_P3_U5189,
    new_P3_U5190, new_P3_U5191, new_P3_U5192, new_P3_U5193, new_P3_U5194,
    new_P3_U5195, new_P3_U5196, new_P3_U5197, new_P3_U5198, new_P3_U5199,
    new_P3_U5200, new_P3_U5201, new_P3_U5202, new_P3_U5203, new_P3_U5204,
    new_P3_U5205, new_P3_U5206, new_P3_U5207, new_P3_U5208, new_P3_U5209,
    new_P3_U5210, new_P3_U5211, new_P3_U5212, new_P3_U5213, new_P3_U5214,
    new_P3_U5215, new_P3_U5216, new_P3_U5217, new_P3_U5218, new_P3_U5219,
    new_P3_U5220, new_P3_U5221, new_P3_U5222, new_P3_U5223, new_P3_U5224,
    new_P3_U5225, new_P3_U5226, new_P3_U5227, new_P3_U5228, new_P3_U5229,
    new_P3_U5230, new_P3_U5231, new_P3_U5232, new_P3_U5233, new_P3_U5234,
    new_P3_U5235, new_P3_U5236, new_P3_U5237, new_P3_U5238, new_P3_U5239,
    new_P3_U5240, new_P3_U5241, new_P3_U5242, new_P3_U5243, new_P3_U5244,
    new_P3_U5245, new_P3_U5246, new_P3_U5247, new_P3_U5248, new_P3_U5249,
    new_P3_U5250, new_P3_U5251, new_P3_U5252, new_P3_U5253, new_P3_U5254,
    new_P3_U5255, new_P3_U5256, new_P3_U5257, new_P3_U5258, new_P3_U5259,
    new_P3_U5260, new_P3_U5261, new_P3_U5262, new_P3_U5263, new_P3_U5264,
    new_P3_U5265, new_P3_U5266, new_P3_U5267, new_P3_U5268, new_P3_U5269,
    new_P3_U5270, new_P3_U5271, new_P3_U5272, new_P3_U5273, new_P3_U5274,
    new_P3_U5275, new_P3_U5276, new_P3_U5277, new_P3_U5278, new_P3_U5279,
    new_P3_U5280, new_P3_U5281, new_P3_U5282, new_P3_U5283, new_P3_U5284,
    new_P3_U5285, new_P3_U5286, new_P3_U5287, new_P3_U5288, new_P3_U5289,
    new_P3_U5290, new_P3_U5291, new_P3_U5292, new_P3_U5293, new_P3_U5294,
    new_P3_U5295, new_P3_U5296, new_P3_U5297, new_P3_U5298, new_P3_U5299,
    new_P3_U5300, new_P3_U5301, new_P3_U5302, new_P3_U5303, new_P3_U5304,
    new_P3_U5305, new_P3_U5306, new_P3_U5307, new_P3_U5308, new_P3_U5309,
    new_P3_U5310, new_P3_U5311, new_P3_U5312, new_P3_U5313, new_P3_U5314,
    new_P3_U5315, new_P3_U5316, new_P3_U5317, new_P3_U5318, new_P3_U5319,
    new_P3_U5320, new_P3_U5321, new_P3_U5322, new_P3_U5323, new_P3_U5324,
    new_P3_U5325, new_P3_U5326, new_P3_U5327, new_P3_U5328, new_P3_U5329,
    new_P3_U5330, new_P3_U5331, new_P3_U5332, new_P3_U5333, new_P3_U5334,
    new_P3_U5335, new_P3_U5336, new_P3_U5337, new_P3_U5338, new_P3_U5339,
    new_P3_U5340, new_P3_U5341, new_P3_U5342, new_P3_U5343, new_P3_U5344,
    new_P3_U5345, new_P3_U5346, new_P3_U5347, new_P3_U5348, new_P3_U5349,
    new_P3_U5350, new_P3_U5351, new_P3_U5352, new_P3_U5353, new_P3_U5354,
    new_P3_U5355, new_P3_U5356, new_P3_U5357, new_P3_U5358, new_P3_U5359,
    new_P3_U5360, new_P3_U5361, new_P3_U5362, new_P3_U5363, new_P3_U5364,
    new_P3_U5365, new_P3_U5366, new_P3_U5367, new_P3_U5368, new_P3_U5369,
    new_P3_U5370, new_P3_U5371, new_P3_U5372, new_P3_U5373, new_P3_U5374,
    new_P3_U5375, new_P3_U5376, new_P3_U5377, new_P3_U5378, new_P3_U5379,
    new_P3_U5380, new_P3_U5381, new_P3_U5382, new_P3_U5383, new_P3_U5384,
    new_P3_U5385, new_P3_U5386, new_P3_U5387, new_P3_U5388, new_P3_U5389,
    new_P3_U5390, new_P3_U5391, new_P3_U5392, new_P3_U5393, new_P3_U5394,
    new_P3_U5395, new_P3_U5396, new_P3_U5397, new_P3_U5398, new_P3_U5399,
    new_P3_U5400, new_P3_U5401, new_P3_U5402, new_P3_U5403, new_P3_U5404,
    new_P3_U5405, new_P3_U5406, new_P3_U5407, new_P3_U5408, new_P3_U5409,
    new_P3_U5410, new_P3_U5411, new_P3_U5412, new_P3_U5413, new_P3_U5414,
    new_P3_U5415, new_P3_U5416, new_P3_U5417, new_P3_U5418, new_P3_U5419,
    new_P3_U5420, new_P3_U5421, new_P3_U5422, new_P3_U5423, new_P3_U5424,
    new_P3_U5425, new_P3_U5426, new_P3_U5427, new_P3_U5428, new_P3_U5429,
    new_P3_U5430, new_P3_U5431, new_P3_U5432, new_P3_U5433, new_P3_U5434,
    new_P3_U5435, new_P3_U5436, new_P3_U5437, new_P3_U5438, new_P3_U5439,
    new_P3_U5440, new_P3_U5441, new_P3_U5442, new_P3_U5443, new_P3_U5444,
    new_P3_U5445, new_P3_U5446, new_P3_U5447, new_P3_U5448, new_P3_U5449,
    new_P3_U5450, new_P3_U5451, new_P3_U5452, new_P3_U5453, new_P3_U5454,
    new_P3_U5455, new_P3_U5456, new_P3_U5457, new_P3_U5458, new_P3_U5459,
    new_P3_U5460, new_P3_U5461, new_P3_U5462, new_P3_U5463, new_P3_U5464,
    new_P3_U5465, new_P3_U5466, new_P3_U5467, new_P3_U5468, new_P3_U5469,
    new_P3_U5470, new_P3_U5471, new_P3_U5472, new_P3_U5473, new_P3_U5474,
    new_P3_U5475, new_P3_U5476, new_P3_U5477, new_P3_U5478, new_P3_U5479,
    new_P3_U5480, new_P3_U5481, new_P3_U5482, new_P3_U5483, new_P3_U5484,
    new_P3_U5485, new_P3_U5486, new_P3_U5487, new_P3_U5488, new_P3_U5489,
    new_P3_U5490, new_P3_U5491, new_P3_U5492, new_P3_U5493, new_P3_U5494,
    new_P3_U5495, new_P3_U5496, new_P3_U5497, new_P3_U5498, new_P3_U5499,
    new_P3_U5500, new_P3_U5501, new_P3_U5502, new_P3_U5503, new_P3_U5504,
    new_P3_U5505, new_P3_U5506, new_P3_U5507, new_P3_U5508, new_P3_U5509,
    new_P3_U5510, new_P3_U5511, new_P3_U5512, new_P3_U5513, new_P3_U5514,
    new_P3_U5515, new_P3_U5516, new_P3_U5517, new_P3_U5518, new_P3_U5519,
    new_P3_U5520, new_P3_U5521, new_P3_U5522, new_P3_U5523, new_P3_U5524,
    new_P3_U5525, new_P3_U5526, new_P3_U5527, new_P3_U5528, new_P3_U5529,
    new_P3_U5530, new_P3_U5531, new_P3_U5532, new_P3_U5533, new_P3_U5534,
    new_P3_U5535, new_P3_U5536, new_P3_U5537, new_P3_U5538, new_P3_U5539,
    new_P3_U5540, new_P3_U5541, new_P3_U5542, new_P3_U5543, new_P3_U5544,
    new_P3_U5545, new_P3_U5546, new_P3_U5547, new_P3_U5548, new_P3_U5549,
    new_P3_U5550, new_P3_U5551, new_P3_U5552, new_P3_U5553, new_P3_U5554,
    new_P3_U5555, new_P3_U5556, new_P3_U5557, new_P3_U5558, new_P3_U5559,
    new_P3_U5560, new_P3_U5561, new_P3_U5562, new_P3_U5563, new_P3_U5564,
    new_P3_U5565, new_P3_U5566, new_P3_U5567, new_P3_U5568, new_P3_U5569,
    new_P3_U5570, new_P3_U5571, new_P3_U5572, new_P3_U5573, new_P3_U5574,
    new_P3_U5575, new_P3_U5576, new_P3_U5577, new_P3_U5578, new_P3_U5579,
    new_P3_U5580, new_P3_U5581, new_P3_U5582, new_P3_U5583, new_P3_U5584,
    new_P3_U5585, new_P3_U5586, new_P3_U5587, new_P3_U5588, new_P3_U5589,
    new_P3_U5590, new_P3_U5591, new_P3_U5592, new_P3_U5593, new_P3_U5594,
    new_P3_U5595, new_P3_U5596, new_P3_U5597, new_P3_U5598, new_P3_U5599,
    new_P3_U5600, new_P3_U5601, new_P3_U5602, new_P3_U5603, new_P3_U5604,
    new_P3_U5605, new_P3_U5606, new_P3_U5607, new_P3_U5608, new_P3_U5609,
    new_P3_U5610, new_P3_U5611, new_P3_U5612, new_P3_U5613, new_P3_U5614,
    new_P3_U5615, new_P3_U5616, new_P3_U5617, new_P3_U5618, new_P3_U5619,
    new_P3_U5620, new_P3_U5621, new_P3_U5622, new_P3_U5623, new_P3_U5624,
    new_P3_U5625, new_P3_U5626, new_P3_U5627, new_P3_U5628, new_P3_U5629,
    new_P3_U5630, new_P3_U5631, new_P3_U5632, new_P3_U5633, new_P3_U5634,
    new_P3_U5635, new_P3_U5636, new_P3_U5637, new_P3_U5638, new_P3_U5639,
    new_P3_U5640, new_P3_U5641, new_P3_U5642, new_P3_U5643, new_P3_U5644,
    new_P3_U5645, new_P3_U5646, new_P3_U5647, new_P3_U5648, new_P3_U5649,
    new_P3_U5650, new_P3_U5651, new_P3_U5652, new_P3_U5653, new_P3_U5654,
    new_P3_U5655, new_P3_U5656, new_P3_U5657, new_P3_U5658, new_P3_U5659,
    new_P3_U5660, new_P3_U5661, new_P3_U5662, new_P3_U5663, new_P3_U5664,
    new_P3_U5665, new_P3_U5666, new_P3_U5667, new_P3_U5668, new_P3_U5669,
    new_P3_U5670, new_P3_U5671, new_P3_U5672, new_P3_U5673, new_P3_U5674,
    new_P3_U5675, new_P3_U5676, new_P3_U5677, new_P3_U5678, new_P3_U5679,
    new_P3_U5680, new_P3_U5681, new_P3_U5682, new_P3_U5683, new_P3_U5684,
    new_P3_U5685, new_P3_U5686, new_P3_U5687, new_P3_U5688, new_P3_U5689,
    new_P3_U5690, new_P3_U5691, new_P3_U5692, new_P3_U5693, new_P3_U5694,
    new_P3_U5695, new_P3_U5696, new_P3_U5697, new_P3_U5698, new_P3_U5699,
    new_P3_U5700, new_P3_U5701, new_P3_U5702, new_P3_U5703, new_P3_U5704,
    new_P3_U5705, new_P3_U5706, new_P3_U5707, new_P3_U5708, new_P3_U5709,
    new_P3_U5710, new_P3_U5711, new_P3_U5712, new_P3_U5713, new_P3_U5714,
    new_P3_U5715, new_P3_U5716, new_P3_U5717, new_P3_U5718, new_P3_U5719,
    new_P3_U5720, new_P3_U5721, new_P3_U5722, new_P3_U5723, new_P3_U5724,
    new_P3_U5725, new_P3_U5726, new_P3_U5727, new_P3_U5728, new_P3_U5729,
    new_P3_U5730, new_P3_U5731, new_P3_U5732, new_P3_U5733, new_P3_U5734,
    new_P3_U5735, new_P3_U5736, new_P3_U5737, new_P3_U5738, new_P3_U5739,
    new_P3_U5740, new_P3_U5741, new_P3_U5742, new_P3_U5743, new_P3_U5744,
    new_P3_U5745, new_P3_U5746, new_P3_U5747, new_P3_U5748, new_P3_U5749,
    new_P3_U5750, new_P3_U5751, new_P3_U5752, new_P3_U5753, new_P3_U5754,
    new_P3_U5755, new_P3_U5756, new_P3_U5757, new_P3_U5758, new_P3_U5759,
    new_P3_U5760, new_P3_U5761, new_P3_U5762, new_P3_U5763, new_P3_U5764,
    new_P3_U5765, new_P3_U5766, new_P3_U5767, new_P3_U5768, new_P3_U5769,
    new_P3_U5770, new_P3_U5771, new_P3_U5772, new_P3_U5773, new_P3_U5774,
    new_P3_U5775, new_P3_U5776, new_P3_U5777, new_P3_U5778, new_P3_U5779,
    new_P3_U5780, new_P3_U5781, new_P3_U5782, new_P3_U5783, new_P3_U5784,
    new_P3_U5785, new_P3_U5786, new_P3_U5787, new_P3_U5788, new_P3_U5789,
    new_P3_U5790, new_P3_U5791, new_P3_U5792, new_P3_U5793, new_P3_U5794,
    new_P3_U5795, new_P3_U5796, new_P3_U5797, new_P3_U5798, new_P3_U5799,
    new_P3_U5800, new_P3_U5801, new_P3_U5802, new_P3_U5803, new_P3_U5804,
    new_P3_U5805, new_P3_U5806, new_P3_U5807, new_P3_U5808, new_P3_U5809,
    new_P3_U5810, new_P3_U5811, new_P3_U5812, new_P3_U5813, new_P3_U5814,
    new_P3_U5815, new_P3_U5816, new_P3_U5817, new_P3_U5818, new_P3_U5819,
    new_P3_U5820, new_P3_U5821, new_P3_U5822, new_P3_U5823, new_P3_U5824,
    new_P3_U5825, new_P3_U5826, new_P3_U5827, new_P3_U5828, new_P3_U5829,
    new_P3_U5830, new_P3_U5831, new_P3_U5832, new_P3_U5833, new_P3_U5834,
    new_P3_U5835, new_P3_U5836, new_P3_U5837, new_P3_U5838, new_P3_U5839,
    new_P3_U5840, new_P3_U5841, new_P3_U5842, new_P3_U5843, new_P3_U5844,
    new_P3_U5845, new_P3_U5846, new_P3_U5847, new_P3_U5848, new_P3_U5849,
    new_P3_U5850, new_P3_U5851, new_P3_U5852, new_P3_U5853, new_P3_U5854,
    new_P3_U5855, new_P3_U5856, new_P3_U5857, new_P3_U5858, new_P3_U5859,
    new_P3_U5860, new_P3_U5861, new_P3_U5862, new_P3_U5863, new_P3_U5864,
    new_P3_U5865, new_P3_U5866, new_P3_U5867, new_P3_U5868, new_P3_U5869,
    new_P3_U5870, new_P3_U5871, new_P3_U5872, new_P3_U5873, new_P3_U5874,
    new_P3_U5875, new_P3_U5876, new_P3_U5877, new_P3_U5878, new_P3_U5879,
    new_P3_U5880, new_P3_U5881, new_P3_U5882, new_P3_U5883, new_P3_U5884,
    new_P3_U5885, new_P3_U5886, new_P3_U5887, new_P3_U5888, new_P3_U5889,
    new_P3_U5890, new_P3_U5891, new_P3_U5892, new_P3_U5893, new_P3_U5894,
    new_P3_U5895, new_P3_U5896, new_P3_U5897, new_P3_U5898, new_P3_U5899,
    new_P3_U5900, new_P3_U5901, new_P3_U5902, new_P3_U5903, new_P3_U5904,
    new_P3_U5905, new_P3_U5906, new_P3_U5907, new_P3_U5908, new_P3_U5909,
    new_P3_U5910, new_P3_U5911, new_P3_U5912, new_P3_U5913, new_P3_U5914,
    new_P3_U5915, new_P3_U5916, new_P3_U5917, new_P3_U5918, new_P3_U5919,
    new_P3_U5920, new_P3_U5921, new_P3_U5922, new_P3_U5923, new_P3_U5924,
    new_P3_U5925, new_P3_U5926, new_P3_U5927, new_P3_U5928, new_P3_U5929,
    new_P3_U5930, new_P3_U5931, new_P3_U5932, new_P3_U5933, new_P3_U5934,
    new_P3_U5935, new_P3_U5936, new_P3_U5937, new_P3_U5938, new_P3_U5939,
    new_P3_U5940, new_P3_U5941, new_P3_U5942, new_P3_U5943, new_P3_U5944,
    new_P3_U5945, new_P3_U5946, new_P3_U5947, new_P3_U5948, new_P3_U5949,
    new_P3_U5950, new_P3_U5951, new_P3_U5952, new_P3_U5953, new_P3_U5954,
    new_P3_U5955, new_P3_U5956, new_P3_U5957, new_P3_U5958, new_P3_U5959,
    new_P3_U5960, new_P3_U5961, new_P3_U5962, new_P3_U5963, new_P3_U5964,
    new_P3_U5965, new_P3_U5966, new_P3_U5967, new_P3_U5968, new_P3_U5969,
    new_P3_U5970, new_P3_U5971, new_P3_U5972, new_P3_U5973, new_P3_U5974,
    new_P3_U5975, new_P3_U5976, new_P3_U5977, new_P3_U5978, new_P3_U5979,
    new_P3_U5980, new_P3_U5981, new_P3_U5982, new_P3_U5983, new_P3_U5984,
    new_P3_U5985, new_P3_U5986, new_P3_U5987, new_P3_U5988, new_P3_U5989,
    new_P3_U5990, new_P3_U5991, new_P3_U5992, new_P3_U5993, new_P3_U5994,
    new_P3_U5995, new_P3_U5996, new_P3_U5997, new_P3_U5998, new_P3_U5999,
    new_P3_U6000, new_P3_U6001, new_P3_U6002, new_P3_U6003, new_P3_U6004,
    new_P3_U6005, new_P3_U6006, new_P3_U6007, new_P3_U6008, new_P3_U6009,
    new_P3_U6010, new_P3_U6011, new_P3_U6012, new_P3_U6013, new_P3_U6014,
    new_P3_U6015, new_P3_U6016, new_P3_U6017, new_P3_U6018, new_P3_U6019,
    new_P3_U6020, new_P3_U6021, new_P3_U6022, new_P3_U6023, new_P3_U6024,
    new_P3_U6025, new_P3_U6026, new_P3_U6027, new_P3_U6028, new_P3_U6029,
    new_P3_U6030, new_P3_U6031, new_P3_U6032, new_P3_U6033, new_P3_U6034,
    new_P3_U6035, new_P3_U6036, new_P3_U6037, new_P3_U6038, new_P3_U6039,
    new_P3_U6040, new_P3_U6041, new_P3_U6042, new_P3_U6043, new_P3_U6044,
    new_P3_U6045, new_P3_U6046, new_P3_U6047, new_P3_U6048,
    new_P3_R1161_U448, new_P3_R1161_U447, new_P3_R1161_U446,
    new_P3_R1161_U445, new_P3_R1161_U444, new_P3_R1161_U443,
    new_P3_R1161_U442, new_P3_R1161_U441, new_P3_R1161_U440,
    new_P3_R1161_U439, new_P3_R1161_U438, new_P3_R1161_U437,
    new_P3_R1161_U436, new_P3_R1161_U435, new_P3_R1161_U434,
    new_P3_R1161_U433, new_P3_R1161_U432, new_P3_R1161_U431,
    new_P3_R1161_U430, new_SUB_1605_U6, new_SUB_1605_U7, new_SUB_1605_U8,
    new_SUB_1605_U9, new_SUB_1605_U10, new_SUB_1605_U11, new_SUB_1605_U12,
    new_SUB_1605_U13, new_SUB_1605_U14, new_SUB_1605_U15, new_SUB_1605_U16,
    new_SUB_1605_U17, new_SUB_1605_U18, new_SUB_1605_U19, new_SUB_1605_U20,
    new_SUB_1605_U21, new_SUB_1605_U22, new_SUB_1605_U23, new_SUB_1605_U24,
    new_SUB_1605_U25, new_SUB_1605_U26, new_SUB_1605_U27, new_SUB_1605_U28,
    new_SUB_1605_U29, new_SUB_1605_U30, new_SUB_1605_U31, new_SUB_1605_U32,
    new_SUB_1605_U33, new_SUB_1605_U34, new_SUB_1605_U35, new_SUB_1605_U36,
    new_SUB_1605_U37, new_SUB_1605_U38, new_SUB_1605_U39, new_SUB_1605_U40,
    new_SUB_1605_U41, new_SUB_1605_U42, new_SUB_1605_U43, new_SUB_1605_U44,
    new_SUB_1605_U45, new_SUB_1605_U46, new_SUB_1605_U47, new_SUB_1605_U48,
    new_SUB_1605_U49, new_SUB_1605_U50, new_SUB_1605_U51, new_SUB_1605_U52,
    new_SUB_1605_U53, new_SUB_1605_U54, new_SUB_1605_U55, new_SUB_1605_U56,
    new_SUB_1605_U57, new_SUB_1605_U58, new_SUB_1605_U59, new_SUB_1605_U60,
    new_SUB_1605_U61, new_SUB_1605_U62, new_SUB_1605_U63, new_SUB_1605_U64,
    new_SUB_1605_U65, new_SUB_1605_U66, new_SUB_1605_U67, new_SUB_1605_U68,
    new_SUB_1605_U69, new_SUB_1605_U70, new_SUB_1605_U71, new_SUB_1605_U72,
    new_SUB_1605_U73, new_SUB_1605_U74, new_SUB_1605_U75, new_SUB_1605_U76,
    new_SUB_1605_U77, new_SUB_1605_U78, new_SUB_1605_U79, new_SUB_1605_U80,
    new_SUB_1605_U81, new_SUB_1605_U82, new_SUB_1605_U83, new_SUB_1605_U84,
    new_SUB_1605_U85, new_SUB_1605_U86, new_SUB_1605_U87, new_SUB_1605_U88,
    new_SUB_1605_U89, new_SUB_1605_U90, new_SUB_1605_U91, new_SUB_1605_U92,
    new_SUB_1605_U93, new_SUB_1605_U94, new_SUB_1605_U95, new_SUB_1605_U96,
    new_SUB_1605_U97, new_SUB_1605_U98, new_SUB_1605_U99,
    new_SUB_1605_U100, new_SUB_1605_U101, new_SUB_1605_U102,
    new_SUB_1605_U103, new_SUB_1605_U104, new_SUB_1605_U105,
    new_SUB_1605_U106, new_SUB_1605_U107, new_SUB_1605_U108,
    new_SUB_1605_U109, new_SUB_1605_U110, new_SUB_1605_U111,
    new_SUB_1605_U112, new_SUB_1605_U113, new_SUB_1605_U114,
    new_SUB_1605_U115, new_SUB_1605_U116, new_SUB_1605_U117,
    new_SUB_1605_U118, new_SUB_1605_U119, new_SUB_1605_U120,
    new_SUB_1605_U121, new_SUB_1605_U122, new_SUB_1605_U123,
    new_SUB_1605_U124, new_SUB_1605_U125, new_SUB_1605_U126,
    new_SUB_1605_U127, new_SUB_1605_U128, new_SUB_1605_U129,
    new_SUB_1605_U130, new_SUB_1605_U131, new_SUB_1605_U132,
    new_SUB_1605_U133, new_SUB_1605_U134, new_SUB_1605_U135,
    new_SUB_1605_U136, new_SUB_1605_U137, new_SUB_1605_U138,
    new_SUB_1605_U139, new_SUB_1605_U140, new_SUB_1605_U141,
    new_SUB_1605_U142, new_SUB_1605_U143, new_SUB_1605_U144,
    new_SUB_1605_U145, new_SUB_1605_U146, new_SUB_1605_U147,
    new_SUB_1605_U148, new_SUB_1605_U149, new_SUB_1605_U150,
    new_SUB_1605_U151, new_SUB_1605_U152, new_SUB_1605_U153,
    new_SUB_1605_U154, new_SUB_1605_U155, new_SUB_1605_U156,
    new_SUB_1605_U157, new_SUB_1605_U158, new_SUB_1605_U159,
    new_SUB_1605_U160, new_SUB_1605_U161, new_SUB_1605_U162,
    new_SUB_1605_U163, new_SUB_1605_U164, new_SUB_1605_U165,
    new_SUB_1605_U166, new_SUB_1605_U167, new_SUB_1605_U168,
    new_SUB_1605_U169, new_SUB_1605_U170, new_SUB_1605_U171,
    new_SUB_1605_U172, new_SUB_1605_U173, new_SUB_1605_U174,
    new_SUB_1605_U175, new_SUB_1605_U176, new_SUB_1605_U177,
    new_SUB_1605_U178, new_SUB_1605_U179, new_SUB_1605_U180,
    new_SUB_1605_U181, new_SUB_1605_U182, new_SUB_1605_U183,
    new_SUB_1605_U184, new_SUB_1605_U185, new_SUB_1605_U186,
    new_SUB_1605_U187, new_SUB_1605_U188, new_SUB_1605_U189,
    new_SUB_1605_U190, new_SUB_1605_U191, new_SUB_1605_U192,
    new_SUB_1605_U193, new_SUB_1605_U194, new_SUB_1605_U195,
    new_SUB_1605_U196, new_SUB_1605_U197, new_SUB_1605_U198,
    new_SUB_1605_U199, new_SUB_1605_U200, new_SUB_1605_U201,
    new_SUB_1605_U202, new_SUB_1605_U203, new_SUB_1605_U204,
    new_SUB_1605_U205, new_SUB_1605_U206, new_SUB_1605_U207,
    new_SUB_1605_U208, new_SUB_1605_U209, new_SUB_1605_U210,
    new_SUB_1605_U211, new_SUB_1605_U212, new_SUB_1605_U213,
    new_SUB_1605_U214, new_SUB_1605_U215, new_SUB_1605_U216,
    new_SUB_1605_U217, new_SUB_1605_U218, new_SUB_1605_U219,
    new_SUB_1605_U220, new_SUB_1605_U221, new_SUB_1605_U222,
    new_SUB_1605_U223, new_SUB_1605_U224, new_SUB_1605_U225,
    new_SUB_1605_U226, new_SUB_1605_U227, new_SUB_1605_U228,
    new_SUB_1605_U229, new_SUB_1605_U230, new_SUB_1605_U231,
    new_SUB_1605_U232, new_SUB_1605_U233, new_SUB_1605_U234,
    new_SUB_1605_U235, new_SUB_1605_U236, new_SUB_1605_U237,
    new_SUB_1605_U238, new_SUB_1605_U239, new_SUB_1605_U240,
    new_SUB_1605_U241, new_SUB_1605_U242, new_SUB_1605_U243,
    new_SUB_1605_U244, new_SUB_1605_U245, new_SUB_1605_U246,
    new_SUB_1605_U247, new_SUB_1605_U248, new_SUB_1605_U249,
    new_SUB_1605_U250, new_SUB_1605_U251, new_SUB_1605_U252,
    new_SUB_1605_U253, new_SUB_1605_U254, new_SUB_1605_U255,
    new_SUB_1605_U256, new_SUB_1605_U257, new_SUB_1605_U258,
    new_SUB_1605_U259, new_SUB_1605_U260, new_SUB_1605_U261,
    new_SUB_1605_U262, new_SUB_1605_U263, new_SUB_1605_U264,
    new_SUB_1605_U265, new_SUB_1605_U266, new_SUB_1605_U267,
    new_SUB_1605_U268, new_SUB_1605_U269, new_SUB_1605_U270,
    new_SUB_1605_U271, new_SUB_1605_U272, new_SUB_1605_U273,
    new_SUB_1605_U274, new_SUB_1605_U275, new_SUB_1605_U276,
    new_SUB_1605_U277, new_SUB_1605_U278, new_SUB_1605_U279,
    new_SUB_1605_U280, new_SUB_1605_U281, new_SUB_1605_U282,
    new_SUB_1605_U283, new_SUB_1605_U284, new_SUB_1605_U285,
    new_SUB_1605_U286, new_SUB_1605_U287, new_SUB_1605_U288,
    new_SUB_1605_U289, new_SUB_1605_U290, new_SUB_1605_U291,
    new_SUB_1605_U292, new_SUB_1605_U293, new_SUB_1605_U294,
    new_SUB_1605_U295, new_SUB_1605_U296, new_SUB_1605_U297,
    new_SUB_1605_U298, new_SUB_1605_U299, new_SUB_1605_U300,
    new_SUB_1605_U301, new_SUB_1605_U302, new_SUB_1605_U303,
    new_SUB_1605_U304, new_SUB_1605_U305, new_SUB_1605_U306,
    new_SUB_1605_U307, new_SUB_1605_U308, new_SUB_1605_U309,
    new_SUB_1605_U310, new_SUB_1605_U311, new_SUB_1605_U312,
    new_SUB_1605_U313, new_SUB_1605_U314, new_SUB_1605_U315,
    new_SUB_1605_U316, new_SUB_1605_U317, new_SUB_1605_U318,
    new_SUB_1605_U319, new_SUB_1605_U320, new_SUB_1605_U321,
    new_SUB_1605_U322, new_SUB_1605_U323, new_SUB_1605_U324,
    new_SUB_1605_U325, new_SUB_1605_U326, new_SUB_1605_U327,
    new_SUB_1605_U328, new_SUB_1605_U329, new_SUB_1605_U330,
    new_SUB_1605_U331, new_SUB_1605_U332, new_SUB_1605_U333,
    new_SUB_1605_U334, new_SUB_1605_U335, new_SUB_1605_U336,
    new_SUB_1605_U337, new_SUB_1605_U338, new_SUB_1605_U339,
    new_SUB_1605_U340, new_SUB_1605_U341, new_SUB_1605_U342,
    new_SUB_1605_U343, new_SUB_1605_U344, new_SUB_1605_U345,
    new_SUB_1605_U346, new_SUB_1605_U347, new_SUB_1605_U348,
    new_SUB_1605_U349, new_SUB_1605_U350, new_SUB_1605_U351,
    new_SUB_1605_U352, new_SUB_1605_U353, new_SUB_1605_U354,
    new_SUB_1605_U355, new_SUB_1605_U356, new_SUB_1605_U357,
    new_SUB_1605_U358, new_SUB_1605_U359, new_SUB_1605_U360,
    new_SUB_1605_U361, new_SUB_1605_U362, new_SUB_1605_U363,
    new_SUB_1605_U364, new_SUB_1605_U365, new_SUB_1605_U366,
    new_SUB_1605_U367, new_SUB_1605_U368, new_SUB_1605_U369,
    new_SUB_1605_U370, new_SUB_1605_U371, new_SUB_1605_U372,
    new_SUB_1605_U373, new_SUB_1605_U374, new_SUB_1605_U375,
    new_SUB_1605_U376, new_SUB_1605_U377, new_SUB_1605_U378,
    new_SUB_1605_U379, new_SUB_1605_U380, new_SUB_1605_U381,
    new_SUB_1605_U382, new_SUB_1605_U383, new_SUB_1605_U384,
    new_SUB_1605_U385, new_SUB_1605_U386, new_SUB_1605_U387,
    new_SUB_1605_U388, new_SUB_1605_U389, new_SUB_1605_U390,
    new_SUB_1605_U391, new_SUB_1605_U392, new_SUB_1605_U393,
    new_SUB_1605_U394, new_SUB_1605_U395, new_SUB_1605_U396,
    new_SUB_1605_U397, new_SUB_1605_U398, new_SUB_1605_U399,
    new_SUB_1605_U400, new_SUB_1605_U401, new_SUB_1605_U402,
    new_SUB_1605_U403, new_SUB_1605_U404, new_SUB_1605_U405,
    new_SUB_1605_U406, new_SUB_1605_U407, new_SUB_1605_U408,
    new_SUB_1605_U409, new_SUB_1605_U410, new_SUB_1605_U411,
    new_SUB_1605_U412, new_SUB_1605_U413, new_SUB_1605_U414,
    new_SUB_1605_U415, new_SUB_1605_U416, new_SUB_1605_U417,
    new_SUB_1605_U418, new_SUB_1605_U419, new_SUB_1605_U420,
    new_SUB_1605_U421, new_SUB_1605_U422, new_SUB_1605_U423,
    new_SUB_1605_U424, new_SUB_1605_U425, new_SUB_1605_U426,
    new_SUB_1605_U427, new_SUB_1605_U428, new_SUB_1605_U429,
    new_SUB_1605_U430, new_SUB_1605_U431, new_SUB_1605_U432,
    new_SUB_1605_U433, new_SUB_1605_U434, new_SUB_1605_U435,
    new_SUB_1605_U436, new_SUB_1605_U437, new_SUB_1605_U438,
    new_SUB_1605_U439, new_SUB_1605_U440, new_SUB_1605_U441,
    new_SUB_1605_U442, new_SUB_1605_U443, new_SUB_1605_U444,
    new_SUB_1605_U445, new_SUB_1605_U446, new_SUB_1605_U447,
    new_SUB_1605_U448, new_SUB_1605_U449, new_SUB_1605_U450,
    new_SUB_1605_U451, new_SUB_1605_U452, new_SUB_1605_U453,
    new_SUB_1605_U454, new_SUB_1605_U455, new_SUB_1605_U456,
    new_SUB_1605_U457, new_SUB_1605_U458, new_SUB_1605_U459,
    new_SUB_1605_U460, new_SUB_1605_U461, new_SUB_1605_U462,
    new_SUB_1605_U463, new_SUB_1605_U464, new_SUB_1605_U465,
    new_SUB_1605_U466, new_SUB_1605_U467, new_SUB_1605_U468,
    new_SUB_1605_U469, new_SUB_1605_U470, new_SUB_1605_U471,
    new_SUB_1605_U472, new_SUB_1605_U473, new_SUB_1605_U474,
    new_SUB_1605_U475, new_SUB_1605_U476, new_SUB_1605_U477,
    new_SUB_1605_U478, new_SUB_1605_U479, new_SUB_1605_U480, new_R152_U4,
    new_R152_U5, new_R152_U6, new_R152_U7, new_R152_U8, new_R152_U9,
    new_R152_U10, new_R152_U11, new_R152_U12, new_R152_U13, new_R152_U14,
    new_R152_U15, new_R152_U16, new_R152_U17, new_R152_U18, new_R152_U19,
    new_R152_U20, new_R152_U21, new_R152_U22, new_R152_U23, new_R152_U24,
    new_R152_U25, new_R152_U26, new_R152_U27, new_R152_U28, new_R152_U29,
    new_R152_U30, new_R152_U31, new_R152_U32, new_R152_U33, new_R152_U34,
    new_R152_U35, new_R152_U36, new_R152_U37, new_R152_U38, new_R152_U39,
    new_R152_U40, new_R152_U41, new_R152_U42, new_R152_U43, new_R152_U44,
    new_R152_U45, new_R152_U46, new_R152_U47, new_R152_U48, new_R152_U49,
    new_R152_U50, new_R152_U51, new_R152_U52, new_R152_U53, new_R152_U54,
    new_R152_U55, new_R152_U56, new_R152_U57, new_R152_U58, new_R152_U59,
    new_R152_U60, new_R152_U61, new_R152_U62, new_R152_U63, new_R152_U64,
    new_R152_U65, new_R152_U66, new_R152_U67, new_R152_U68, new_R152_U69,
    new_R152_U70, new_R152_U71, new_R152_U72, new_R152_U73, new_R152_U74,
    new_R152_U75, new_R152_U76, new_R152_U77, new_R152_U78, new_R152_U79,
    new_R152_U80, new_R152_U81, new_R152_U82, new_R152_U83, new_R152_U84,
    new_R152_U85, new_R152_U86, new_R152_U87, new_R152_U88, new_R152_U89,
    new_R152_U90, new_R152_U91, new_R152_U92, new_R152_U93, new_R152_U94,
    new_R152_U95, new_R152_U96, new_R152_U97, new_R152_U98, new_R152_U99,
    new_R152_U100, new_R152_U101, new_R152_U102, new_R152_U103,
    new_R152_U104, new_R152_U105, new_R152_U106, new_R152_U107,
    new_R152_U108, new_R152_U109, new_R152_U110, new_R152_U111,
    new_R152_U112, new_R152_U113, new_R152_U114, new_R152_U115,
    new_R152_U116, new_R152_U117, new_R152_U118, new_R152_U119,
    new_R152_U120, new_R152_U121, new_R152_U122, new_R152_U123,
    new_R152_U124, new_R152_U125, new_R152_U126, new_R152_U127,
    new_R152_U128, new_R152_U129, new_R152_U130, new_R152_U131,
    new_R152_U132, new_R152_U133, new_R152_U134, new_R152_U135,
    new_R152_U136, new_R152_U137, new_R152_U138, new_R152_U139,
    new_R152_U140, new_R152_U141, new_R152_U142, new_R152_U143,
    new_R152_U144, new_R152_U145, new_R152_U146, new_R152_U147,
    new_R152_U148, new_R152_U149, new_R152_U150, new_R152_U151,
    new_R152_U152, new_R152_U153, new_R152_U154, new_R152_U155,
    new_R152_U156, new_R152_U157, new_R152_U158, new_R152_U159,
    new_R152_U160, new_R152_U161, new_R152_U162, new_R152_U163,
    new_R152_U164, new_R152_U165, new_R152_U166, new_R152_U167,
    new_R152_U168, new_R152_U169, new_R152_U170, new_R152_U171,
    new_R152_U172, new_R152_U173, new_R152_U174, new_R152_U175,
    new_R152_U176, new_R152_U177, new_R152_U178, new_R152_U179,
    new_R152_U180, new_R152_U181, new_R152_U182, new_R152_U183,
    new_R152_U184, new_R152_U185, new_R152_U186, new_R152_U187,
    new_R152_U188, new_R152_U189, new_R152_U190, new_R152_U191,
    new_R152_U192, new_R152_U193, new_R152_U194, new_R152_U195,
    new_R152_U196, new_R152_U197, new_R152_U198, new_R152_U199,
    new_R152_U200, new_R152_U201, new_R152_U202, new_R152_U203,
    new_R152_U204, new_R152_U205, new_R152_U206, new_R152_U207,
    new_R152_U208, new_R152_U209, new_R152_U210, new_R152_U211,
    new_R152_U212, new_R152_U213, new_R152_U214, new_R152_U215,
    new_R152_U216, new_R152_U217, new_R152_U218, new_R152_U219,
    new_R152_U220, new_R152_U221, new_R152_U222, new_R152_U223,
    new_R152_U224, new_R152_U225, new_R152_U226, new_R152_U227,
    new_R152_U228, new_R152_U229, new_R152_U230, new_R152_U231,
    new_R152_U232, new_R152_U233, new_R152_U234, new_R152_U235,
    new_R152_U236, new_R152_U237, new_R152_U238, new_R152_U239,
    new_R152_U240, new_R152_U241, new_R152_U242, new_R152_U243,
    new_R152_U244, new_R152_U245, new_R152_U246, new_R152_U247,
    new_R152_U248, new_R152_U249, new_R152_U250, new_R152_U251,
    new_R152_U252, new_R152_U253, new_R152_U254, new_R152_U255,
    new_R152_U256, new_R152_U257, new_R152_U258, new_R152_U259,
    new_R152_U260, new_R152_U261, new_R152_U262, new_R152_U263,
    new_R152_U264, new_R152_U265, new_R152_U266, new_R152_U267,
    new_R152_U268, new_R152_U269, new_R152_U270, new_R152_U271,
    new_R152_U272, new_R152_U273, new_R152_U274, new_R152_U275,
    new_R152_U276, new_R152_U277, new_R152_U278, new_R152_U279,
    new_R152_U280, new_R152_U281, new_R152_U282, new_R152_U283,
    new_R152_U284, new_R152_U285, new_R152_U286, new_R152_U287,
    new_R152_U288, new_R152_U289, new_R152_U290, new_R152_U291,
    new_R152_U292, new_R152_U293, new_R152_U294, new_R152_U295,
    new_R152_U296, new_R152_U297, new_R152_U298, new_R152_U299,
    new_R152_U300, new_R152_U301, new_R152_U302, new_R152_U303,
    new_R152_U304, new_R152_U305, new_R152_U306, new_R152_U307,
    new_R152_U308, new_R152_U309, new_R152_U310, new_R152_U311,
    new_R152_U312, new_R152_U313, new_R152_U314, new_R152_U315,
    new_R152_U316, new_R152_U317, new_R152_U318, new_R152_U319,
    new_R152_U320, new_R152_U321, new_R152_U322, new_R152_U323,
    new_R152_U324, new_R152_U325, new_R152_U326, new_R152_U327,
    new_R152_U328, new_R152_U329, new_R152_U330, new_R152_U331,
    new_R152_U332, new_R152_U333, new_R152_U334, new_R152_U335,
    new_R152_U336, new_R152_U337, new_R152_U338, new_R152_U339,
    new_R152_U340, new_R152_U341, new_R152_U342, new_R152_U343,
    new_R152_U344, new_R152_U345, new_R152_U346, new_R152_U347,
    new_R152_U348, new_R152_U349, new_R152_U350, new_R152_U351,
    new_R152_U352, new_R152_U353, new_R152_U354, new_R152_U355,
    new_R152_U356, new_R152_U357, new_R152_U358, new_R152_U359,
    new_R152_U360, new_R152_U361, new_R152_U362, new_R152_U363,
    new_R152_U364, new_R152_U365, new_R152_U366, new_R152_U367,
    new_R152_U368, new_R152_U369, new_R152_U370, new_R152_U371,
    new_R152_U372, new_R152_U373, new_R152_U374, new_R152_U375,
    new_R152_U376, new_R152_U377, new_R152_U378, new_R152_U379,
    new_R152_U380, new_R152_U381, new_R152_U382, new_R152_U383,
    new_R152_U384, new_R152_U385, new_R152_U386, new_R152_U387,
    new_R152_U388, new_R152_U389, new_R152_U390, new_R152_U391,
    new_R152_U392, new_R152_U393, new_R152_U394, new_R152_U395,
    new_R152_U396, new_R152_U397, new_R152_U398, new_R152_U399,
    new_R152_U400, new_R152_U401, new_R152_U402, new_R152_U403,
    new_R152_U404, new_R152_U405, new_R152_U406, new_R152_U407,
    new_R152_U408, new_R152_U409, new_R152_U410, new_R152_U411,
    new_R152_U412, new_R152_U413, new_R152_U414, new_R152_U415,
    new_R152_U416, new_R152_U417, new_R152_U418, new_R152_U419,
    new_R152_U420, new_R152_U421, new_R152_U422, new_R152_U423,
    new_R152_U424, new_R152_U425, new_R152_U426, new_R152_U427,
    new_R152_U428, new_R152_U429, new_R152_U430, new_R152_U431,
    new_R152_U432, new_R152_U433, new_R152_U434, new_R152_U435,
    new_R152_U436, new_R152_U437, new_R152_U438, new_R152_U439,
    new_R152_U440, new_R152_U441, new_R152_U442, new_R152_U443,
    new_R152_U444, new_R152_U445, new_R152_U446, new_R152_U447,
    new_R152_U448, new_R152_U449, new_R152_U450, new_R152_U451,
    new_R152_U452, new_R152_U453, new_R152_U454, new_R152_U455,
    new_R152_U456, new_R152_U457, new_R152_U458, new_R152_U459,
    new_R152_U460, new_R152_U461, new_R152_U462, new_R152_U463,
    new_R152_U464, new_R152_U465, new_R152_U466, new_R152_U467,
    new_R152_U468, new_R152_U469, new_R152_U470, new_R152_U471,
    new_R152_U472, new_R152_U473, new_R152_U474, new_R152_U475,
    new_R152_U476, new_R152_U477, new_R152_U478, new_R152_U479,
    new_R152_U480, new_R152_U481, new_R152_U482, new_R152_U483,
    new_R152_U484, new_R152_U485, new_R152_U486, new_R152_U487,
    new_R152_U488, new_R152_U489, new_R152_U490, new_R152_U491,
    new_R152_U492, new_R152_U493, new_R152_U494, new_R152_U495,
    new_R152_U496, new_R152_U497, new_R152_U498, new_R152_U499,
    new_R152_U500, new_R152_U501, new_R152_U502, new_R152_U503,
    new_R152_U504, new_R152_U505, new_R152_U506, new_R152_U507,
    new_R152_U508, new_R152_U509, new_R152_U510, new_R152_U511,
    new_R152_U512, new_R152_U513, new_R152_U514, new_R152_U515,
    new_R152_U516, new_R152_U517, new_R152_U518, new_R152_U519,
    new_R152_U520, new_R152_U521, new_R152_U522, new_R152_U523,
    new_R152_U524, new_R152_U525, new_R152_U526, new_R152_U527,
    new_R152_U528, new_R152_U529, new_R152_U530, new_R152_U531,
    new_R152_U532, new_R152_U533, new_R152_U534, new_R152_U535,
    new_R152_U536, new_R152_U537, new_R152_U538, new_R152_U539,
    new_R152_U540, new_R152_U541, new_R152_U542, new_R152_U543,
    new_R152_U544, new_R152_U545, new_R152_U546, new_R152_U547,
    new_R152_U548, new_R152_U549, new_R152_U550, new_R152_U551,
    new_R152_U552, new_R152_U553, new_R152_U554, new_LT_1602_U6,
    new_LT_1601_U6, new_SUB_1596_U6, new_SUB_1596_U7, new_SUB_1596_U8,
    new_SUB_1596_U9, new_SUB_1596_U10, new_SUB_1596_U11, new_SUB_1596_U12,
    new_SUB_1596_U13, new_SUB_1596_U14, new_SUB_1596_U15, new_SUB_1596_U16,
    new_SUB_1596_U17, new_SUB_1596_U18, new_SUB_1596_U19, new_SUB_1596_U20,
    new_SUB_1596_U21, new_SUB_1596_U22, new_SUB_1596_U23, new_SUB_1596_U24,
    new_SUB_1596_U25, new_SUB_1596_U26, new_SUB_1596_U27, new_SUB_1596_U28,
    new_SUB_1596_U29, new_SUB_1596_U30, new_SUB_1596_U31, new_SUB_1596_U32,
    new_SUB_1596_U33, new_SUB_1596_U34, new_SUB_1596_U35, new_SUB_1596_U36,
    new_SUB_1596_U37, new_SUB_1596_U38, new_SUB_1596_U39, new_SUB_1596_U40,
    new_SUB_1596_U41, new_SUB_1596_U42, new_SUB_1596_U43, new_SUB_1596_U44,
    new_SUB_1596_U45, new_SUB_1596_U46, new_SUB_1596_U47, new_SUB_1596_U48,
    new_SUB_1596_U49, new_SUB_1596_U50, new_SUB_1596_U51, new_SUB_1596_U52,
    new_SUB_1596_U71, new_SUB_1596_U72, new_SUB_1596_U73, new_SUB_1596_U74,
    new_SUB_1596_U75, new_SUB_1596_U76, new_SUB_1596_U77, new_SUB_1596_U78,
    new_SUB_1596_U79, new_SUB_1596_U80, new_SUB_1596_U81, new_SUB_1596_U82,
    new_SUB_1596_U83, new_SUB_1596_U84, new_SUB_1596_U85, new_SUB_1596_U86,
    new_SUB_1596_U87, new_SUB_1596_U88, new_SUB_1596_U89, new_SUB_1596_U90,
    new_SUB_1596_U91, new_SUB_1596_U92, new_SUB_1596_U93, new_SUB_1596_U94,
    new_SUB_1596_U95, new_SUB_1596_U96, new_SUB_1596_U97, new_SUB_1596_U98,
    new_SUB_1596_U99, new_SUB_1596_U100, new_SUB_1596_U101,
    new_SUB_1596_U102, new_SUB_1596_U103, new_SUB_1596_U104,
    new_SUB_1596_U105, new_SUB_1596_U106, new_SUB_1596_U107,
    new_SUB_1596_U108, new_SUB_1596_U109, new_SUB_1596_U110,
    new_SUB_1596_U111, new_SUB_1596_U112, new_SUB_1596_U113,
    new_SUB_1596_U114, new_SUB_1596_U115, new_SUB_1596_U116,
    new_SUB_1596_U117, new_SUB_1596_U118, new_SUB_1596_U119,
    new_SUB_1596_U120, new_SUB_1596_U121, new_SUB_1596_U122,
    new_SUB_1596_U123, new_SUB_1596_U124, new_SUB_1596_U125,
    new_SUB_1596_U126, new_SUB_1596_U127, new_SUB_1596_U128,
    new_SUB_1596_U129, new_SUB_1596_U130, new_SUB_1596_U131,
    new_SUB_1596_U132, new_SUB_1596_U133, new_SUB_1596_U134,
    new_SUB_1596_U135, new_SUB_1596_U136, new_SUB_1596_U137,
    new_SUB_1596_U138, new_SUB_1596_U139, new_SUB_1596_U140,
    new_SUB_1596_U141, new_SUB_1596_U142, new_SUB_1596_U143,
    new_SUB_1596_U144, new_SUB_1596_U145, new_SUB_1596_U146,
    new_SUB_1596_U147, new_SUB_1596_U148, new_SUB_1596_U149,
    new_SUB_1596_U150, new_SUB_1596_U151, new_SUB_1596_U152,
    new_SUB_1596_U153, new_SUB_1596_U154, new_SUB_1596_U155,
    new_SUB_1596_U156, new_SUB_1596_U157, new_SUB_1596_U158,
    new_SUB_1596_U159, new_SUB_1596_U160, new_SUB_1596_U161,
    new_SUB_1596_U162, new_SUB_1596_U163, new_SUB_1596_U164,
    new_SUB_1596_U165, new_SUB_1596_U166, new_SUB_1596_U167,
    new_SUB_1596_U168, new_SUB_1596_U169, new_SUB_1596_U170,
    new_SUB_1596_U171, new_SUB_1596_U172, new_SUB_1596_U173,
    new_SUB_1596_U174, new_SUB_1596_U175, new_SUB_1596_U176,
    new_SUB_1596_U177, new_SUB_1596_U178, new_SUB_1596_U179,
    new_SUB_1596_U180, new_SUB_1596_U181, new_SUB_1596_U182,
    new_SUB_1596_U183, new_SUB_1596_U184, new_SUB_1596_U185,
    new_SUB_1596_U186, new_SUB_1596_U187, new_SUB_1596_U188,
    new_SUB_1596_U189, new_SUB_1596_U190, new_SUB_1596_U191,
    new_SUB_1596_U192, new_SUB_1596_U193, new_SUB_1596_U194,
    new_SUB_1596_U195, new_SUB_1596_U196, new_SUB_1596_U197,
    new_SUB_1596_U198, new_SUB_1596_U199, new_SUB_1596_U200,
    new_SUB_1596_U201, new_SUB_1596_U202, new_SUB_1596_U203,
    new_SUB_1596_U204, new_SUB_1596_U205, new_SUB_1596_U206,
    new_SUB_1596_U207, new_SUB_1596_U208, new_SUB_1596_U209,
    new_SUB_1596_U210, new_SUB_1596_U211, new_SUB_1596_U212,
    new_SUB_1596_U213, new_SUB_1596_U214, new_SUB_1596_U215,
    new_SUB_1596_U216, new_SUB_1596_U217, new_SUB_1596_U218,
    new_SUB_1596_U219, new_SUB_1596_U220, new_SUB_1596_U221,
    new_SUB_1596_U222, new_SUB_1596_U223, new_SUB_1596_U224,
    new_SUB_1596_U225, new_SUB_1596_U226, new_SUB_1596_U227,
    new_SUB_1596_U228, new_SUB_1596_U229, new_SUB_1596_U230,
    new_SUB_1596_U231, new_SUB_1596_U232, new_SUB_1596_U233,
    new_SUB_1596_U234, new_SUB_1596_U235, new_SUB_1596_U236,
    new_SUB_1596_U237, new_SUB_1596_U238, new_SUB_1596_U239,
    new_SUB_1596_U240, new_SUB_1596_U241, new_SUB_1596_U242,
    new_SUB_1596_U243, new_SUB_1596_U244, new_SUB_1596_U245,
    new_SUB_1596_U246, new_SUB_1596_U247, new_SUB_1596_U248,
    new_SUB_1596_U249, new_SUB_1596_U250, new_SUB_1596_U251,
    new_SUB_1596_U252, new_SUB_1596_U253, new_SUB_1596_U254,
    new_SUB_1596_U255, new_SUB_1596_U256, new_SUB_1596_U257,
    new_SUB_1596_U258, new_SUB_1596_U259, new_SUB_1596_U260,
    new_SUB_1596_U261, new_SUB_1596_U262, new_SUB_1596_U263,
    new_SUB_1596_U264, new_SUB_1596_U265, new_SUB_1596_U266,
    new_SUB_1596_U267, new_SUB_1596_U268, new_SUB_1596_U269,
    new_SUB_1596_U270, new_SUB_1596_U271, new_SUB_1596_U272,
    new_SUB_1596_U273, new_SUB_1596_U274, new_SUB_1596_U275,
    new_SUB_1596_U276, new_SUB_1596_U277, new_SUB_1596_U278,
    new_SUB_1596_U279, new_SUB_1596_U280, new_SUB_1596_U281,
    new_SUB_1596_U282, new_SUB_1596_U283, new_SUB_1596_U284,
    new_SUB_1596_U285, new_SUB_1596_U286, new_SUB_1596_U287,
    new_SUB_1596_U288, new_SUB_1596_U289, new_SUB_1596_U290,
    new_SUB_1596_U291, new_ADD_1596_U6, new_ADD_1596_U7, new_ADD_1596_U8,
    new_ADD_1596_U9, new_ADD_1596_U10, new_ADD_1596_U11, new_ADD_1596_U12,
    new_ADD_1596_U13, new_ADD_1596_U14, new_ADD_1596_U15, new_ADD_1596_U16,
    new_ADD_1596_U17, new_ADD_1596_U18, new_ADD_1596_U19, new_ADD_1596_U20,
    new_ADD_1596_U21, new_ADD_1596_U22, new_ADD_1596_U23, new_ADD_1596_U24,
    new_ADD_1596_U25, new_ADD_1596_U26, new_ADD_1596_U27, new_ADD_1596_U28,
    new_ADD_1596_U29, new_ADD_1596_U30, new_ADD_1596_U31, new_ADD_1596_U32,
    new_ADD_1596_U33, new_ADD_1596_U34, new_ADD_1596_U35, new_ADD_1596_U36,
    new_ADD_1596_U37, new_ADD_1596_U38, new_ADD_1596_U39, new_ADD_1596_U40,
    new_ADD_1596_U41, new_ADD_1596_U42, new_ADD_1596_U43, new_ADD_1596_U44,
    new_ADD_1596_U45, new_ADD_1596_U46, new_ADD_1596_U47, new_ADD_1596_U48,
    new_ADD_1596_U49, new_ADD_1596_U50, new_ADD_1596_U51, new_ADD_1596_U52,
    new_ADD_1596_U53, new_ADD_1596_U54, new_ADD_1596_U55, new_ADD_1596_U56,
    new_ADD_1596_U57, new_ADD_1596_U58, new_ADD_1596_U59, new_ADD_1596_U60,
    new_ADD_1596_U61, new_ADD_1596_U62, new_ADD_1596_U63, new_ADD_1596_U64,
    new_ADD_1596_U65, new_ADD_1596_U66, new_ADD_1596_U67, new_ADD_1596_U68,
    new_ADD_1596_U69, new_ADD_1596_U70, new_ADD_1596_U71, new_ADD_1596_U72,
    new_ADD_1596_U73, new_ADD_1596_U74, new_ADD_1596_U75, new_ADD_1596_U76,
    new_ADD_1596_U77, new_ADD_1596_U78, new_ADD_1596_U79, new_ADD_1596_U80,
    new_ADD_1596_U81, new_ADD_1596_U82, new_ADD_1596_U83, new_ADD_1596_U84,
    new_ADD_1596_U85, new_ADD_1596_U86, new_ADD_1596_U87, new_ADD_1596_U88,
    new_ADD_1596_U89, new_ADD_1596_U90, new_ADD_1596_U91, new_ADD_1596_U92,
    new_ADD_1596_U93, new_ADD_1596_U94, new_ADD_1596_U95, new_ADD_1596_U96,
    new_ADD_1596_U97, new_ADD_1596_U98, new_ADD_1596_U99,
    new_ADD_1596_U100, new_ADD_1596_U101, new_ADD_1596_U102,
    new_ADD_1596_U103, new_ADD_1596_U104, new_ADD_1596_U105,
    new_ADD_1596_U106, new_ADD_1596_U107, new_ADD_1596_U108,
    new_ADD_1596_U109, new_ADD_1596_U110, new_ADD_1596_U111,
    new_ADD_1596_U112, new_ADD_1596_U113, new_ADD_1596_U114,
    new_ADD_1596_U115, new_ADD_1596_U116, new_ADD_1596_U117,
    new_ADD_1596_U118, new_ADD_1596_U119, new_ADD_1596_U120,
    new_ADD_1596_U121, new_ADD_1596_U122, new_ADD_1596_U123,
    new_ADD_1596_U124, new_ADD_1596_U125, new_ADD_1596_U126,
    new_ADD_1596_U127, new_ADD_1596_U128, new_ADD_1596_U129,
    new_ADD_1596_U130, new_ADD_1596_U131, new_ADD_1596_U132,
    new_ADD_1596_U133, new_ADD_1596_U134, new_ADD_1596_U135,
    new_ADD_1596_U136, new_ADD_1596_U137, new_ADD_1596_U138,
    new_ADD_1596_U139, new_ADD_1596_U140, new_ADD_1596_U141,
    new_ADD_1596_U142, new_ADD_1596_U143, new_ADD_1596_U144,
    new_ADD_1596_U145, new_ADD_1596_U146, new_ADD_1596_U147,
    new_ADD_1596_U148, new_ADD_1596_U149, new_ADD_1596_U150,
    new_ADD_1596_U151, new_ADD_1596_U152, new_ADD_1596_U153,
    new_ADD_1596_U154, new_ADD_1596_U155, new_ADD_1596_U156,
    new_ADD_1596_U157, new_ADD_1596_U158, new_ADD_1596_U159,
    new_ADD_1596_U160, new_ADD_1596_U161, new_ADD_1596_U162,
    new_ADD_1596_U163, new_ADD_1596_U164, new_ADD_1596_U165,
    new_ADD_1596_U166, new_ADD_1596_U167, new_ADD_1596_U168,
    new_ADD_1596_U169, new_ADD_1596_U170, new_ADD_1596_U171,
    new_ADD_1596_U172, new_ADD_1596_U173, new_ADD_1596_U174,
    new_ADD_1596_U175, new_ADD_1596_U176, new_ADD_1596_U177,
    new_ADD_1596_U178, new_ADD_1596_U179, new_ADD_1596_U180,
    new_ADD_1596_U181, new_ADD_1596_U182, new_ADD_1596_U183,
    new_ADD_1596_U184, new_ADD_1596_U185, new_ADD_1596_U186,
    new_ADD_1596_U187, new_ADD_1596_U188, new_ADD_1596_U189,
    new_ADD_1596_U190, new_ADD_1596_U191, new_ADD_1596_U192,
    new_ADD_1596_U193, new_ADD_1596_U194, new_ADD_1596_U195,
    new_ADD_1596_U196, new_ADD_1596_U197, new_ADD_1596_U198,
    new_ADD_1596_U199, new_ADD_1596_U200, new_ADD_1596_U201,
    new_ADD_1596_U202, new_ADD_1596_U203, new_ADD_1596_U204,
    new_ADD_1596_U205, new_ADD_1596_U206, new_ADD_1596_U207,
    new_ADD_1596_U208, new_ADD_1596_U209, new_ADD_1596_U210,
    new_ADD_1596_U211, new_ADD_1596_U212, new_ADD_1596_U213,
    new_ADD_1596_U214, new_ADD_1596_U215, new_ADD_1596_U216,
    new_ADD_1596_U217, new_ADD_1596_U218, new_ADD_1596_U219,
    new_ADD_1596_U220, new_ADD_1596_U221, new_ADD_1596_U222,
    new_ADD_1596_U223, new_ADD_1596_U224, new_ADD_1596_U225,
    new_ADD_1596_U226, new_ADD_1596_U227, new_ADD_1596_U228,
    new_ADD_1596_U229, new_ADD_1596_U230, new_ADD_1596_U231,
    new_ADD_1596_U232, new_ADD_1596_U233, new_ADD_1596_U234,
    new_ADD_1596_U235, new_ADD_1596_U236, new_ADD_1596_U237,
    new_ADD_1596_U238, new_ADD_1596_U239, new_ADD_1596_U240,
    new_ADD_1596_U241, new_ADD_1596_U242, new_ADD_1596_U243,
    new_ADD_1596_U244, new_ADD_1596_U245, new_ADD_1596_U246,
    new_ADD_1596_U247, new_ADD_1596_U248, new_ADD_1596_U249,
    new_ADD_1596_U250, new_ADD_1596_U251, new_ADD_1596_U252,
    new_ADD_1596_U253, new_ADD_1596_U254, new_ADD_1596_U255,
    new_ADD_1596_U256, new_ADD_1596_U257, new_ADD_1596_U258,
    new_ADD_1596_U259, new_ADD_1596_U260, new_ADD_1596_U261,
    new_ADD_1596_U262, new_ADD_1596_U263, new_ADD_1596_U264,
    new_ADD_1596_U265, new_ADD_1596_U266, new_ADD_1596_U267,
    new_ADD_1596_U268, new_ADD_1596_U269, new_ADD_1596_U270,
    new_ADD_1596_U271, new_ADD_1596_U272, new_ADD_1596_U273,
    new_ADD_1596_U274, new_LT_1601_21_U6, new_P1_ADD_99_U4,
    new_P1_ADD_99_U5, new_P1_ADD_99_U6, new_P1_ADD_99_U7, new_P1_ADD_99_U8,
    new_P1_ADD_99_U9, new_P1_ADD_99_U10, new_P1_ADD_99_U11,
    new_P1_ADD_99_U12, new_P1_ADD_99_U13, new_P1_ADD_99_U14,
    new_P1_ADD_99_U15, new_P1_ADD_99_U16, new_P1_ADD_99_U17,
    new_P1_ADD_99_U18, new_P1_ADD_99_U19, new_P1_ADD_99_U20,
    new_P1_ADD_99_U21, new_P1_ADD_99_U22, new_P1_ADD_99_U23,
    new_P1_ADD_99_U24, new_P1_ADD_99_U25, new_P1_ADD_99_U26,
    new_P1_ADD_99_U27, new_P1_ADD_99_U28, new_P1_ADD_99_U29,
    new_P1_ADD_99_U30, new_P1_ADD_99_U31, new_P1_ADD_99_U32,
    new_P1_ADD_99_U33, new_P1_ADD_99_U34, new_P1_ADD_99_U35,
    new_P1_ADD_99_U36, new_P1_ADD_99_U37, new_P1_ADD_99_U38,
    new_P1_ADD_99_U39, new_P1_ADD_99_U40, new_P1_ADD_99_U41,
    new_P1_ADD_99_U42, new_P1_ADD_99_U43, new_P1_ADD_99_U44,
    new_P1_ADD_99_U45, new_P1_ADD_99_U46, new_P1_ADD_99_U47,
    new_P1_ADD_99_U48, new_P1_ADD_99_U49, new_P1_ADD_99_U50,
    new_P1_ADD_99_U51, new_P1_ADD_99_U52, new_P1_ADD_99_U53,
    new_P1_ADD_99_U54, new_P1_ADD_99_U55, new_P1_ADD_99_U56,
    new_P1_ADD_99_U57, new_P1_ADD_99_U58, new_P1_ADD_99_U59,
    new_P1_ADD_99_U60, new_P1_ADD_99_U61, new_P1_ADD_99_U62,
    new_P1_ADD_99_U63, new_P1_ADD_99_U64, new_P1_ADD_99_U65,
    new_P1_ADD_99_U66, new_P1_ADD_99_U67, new_P1_ADD_99_U68,
    new_P1_ADD_99_U69, new_P1_ADD_99_U70, new_P1_ADD_99_U71,
    new_P1_ADD_99_U72, new_P1_ADD_99_U73, new_P1_ADD_99_U74,
    new_P1_ADD_99_U75, new_P1_ADD_99_U76, new_P1_ADD_99_U77,
    new_P1_ADD_99_U78, new_P1_ADD_99_U79, new_P1_ADD_99_U80,
    new_P1_ADD_99_U81, new_P1_ADD_99_U82, new_P1_ADD_99_U83,
    new_P1_ADD_99_U84, new_P1_ADD_99_U85, new_P1_ADD_99_U86,
    new_P1_ADD_99_U87, new_P1_ADD_99_U88, new_P1_ADD_99_U89,
    new_P1_ADD_99_U90, new_P1_ADD_99_U91, new_P1_ADD_99_U92,
    new_P1_ADD_99_U93, new_P1_ADD_99_U94, new_P1_ADD_99_U95,
    new_P1_ADD_99_U96, new_P1_ADD_99_U97, new_P1_ADD_99_U98,
    new_P1_ADD_99_U99, new_P1_ADD_99_U100, new_P1_ADD_99_U101,
    new_P1_ADD_99_U102, new_P1_ADD_99_U103, new_P1_ADD_99_U104,
    new_P1_ADD_99_U105, new_P1_ADD_99_U106, new_P1_ADD_99_U107,
    new_P1_ADD_99_U108, new_P1_ADD_99_U109, new_P1_ADD_99_U110,
    new_P1_ADD_99_U111, new_P1_ADD_99_U112, new_P1_ADD_99_U113,
    new_P1_ADD_99_U114, new_P1_ADD_99_U115, new_P1_ADD_99_U116,
    new_P1_ADD_99_U117, new_P1_ADD_99_U118, new_P1_ADD_99_U119,
    new_P1_ADD_99_U120, new_P1_ADD_99_U121, new_P1_ADD_99_U122,
    new_P1_ADD_99_U123, new_P1_ADD_99_U124, new_P1_ADD_99_U125,
    new_P1_ADD_99_U126, new_P1_ADD_99_U127, new_P1_ADD_99_U128,
    new_P1_ADD_99_U129, new_P1_ADD_99_U130, new_P1_ADD_99_U131,
    new_P1_ADD_99_U132, new_P1_ADD_99_U133, new_P1_ADD_99_U134,
    new_P1_ADD_99_U135, new_P1_ADD_99_U136, new_P1_ADD_99_U137,
    new_P1_ADD_99_U138, new_P1_ADD_99_U139, new_P1_ADD_99_U140,
    new_P1_ADD_99_U141, new_P1_ADD_99_U142, new_P1_ADD_99_U143,
    new_P1_ADD_99_U144, new_P1_ADD_99_U145, new_P1_ADD_99_U146,
    new_P1_ADD_99_U147, new_P1_ADD_99_U148, new_P1_ADD_99_U149,
    new_P1_ADD_99_U150, new_P1_ADD_99_U151, new_P1_ADD_99_U152,
    new_P1_ADD_99_U153, new_P1_R1105_U4, new_P1_R1105_U5, new_P1_R1105_U6,
    new_P1_R1105_U7, new_P1_R1105_U8, new_P1_R1105_U9, new_P1_R1105_U10,
    new_P1_R1105_U11, new_P1_R1105_U12, new_P1_R1105_U13, new_P1_R1105_U14,
    new_P1_R1105_U15, new_P1_R1105_U16, new_P1_R1105_U17, new_P1_R1105_U18,
    new_P1_R1105_U19, new_P1_R1105_U20, new_P1_R1105_U21, new_P1_R1105_U22,
    new_P1_R1105_U23, new_P1_R1105_U24, new_P1_R1105_U25, new_P1_R1105_U26,
    new_P1_R1105_U27, new_P1_R1105_U28, new_P1_R1105_U29, new_P1_R1105_U30,
    new_P1_R1105_U31, new_P1_R1105_U32, new_P1_R1105_U33, new_P1_R1105_U34,
    new_P1_R1105_U35, new_P1_R1105_U36, new_P1_R1105_U37, new_P1_R1105_U38,
    new_P1_R1105_U39, new_P1_R1105_U40, new_P1_R1105_U41, new_P1_R1105_U42,
    new_P1_R1105_U43, new_P1_R1105_U44, new_P1_R1105_U45, new_P1_R1105_U46,
    new_P1_R1105_U47, new_P1_R1105_U48, new_P1_R1105_U49, new_P1_R1105_U50,
    new_P1_R1105_U51, new_P1_R1105_U52, new_P1_R1105_U53, new_P1_R1105_U54,
    new_P1_R1105_U55, new_P1_R1105_U56, new_P1_R1105_U57, new_P1_R1105_U58,
    new_P1_R1105_U59, new_P1_R1105_U60, new_P1_R1105_U61, new_P1_R1105_U62,
    new_P1_R1105_U63, new_P1_R1105_U64, new_P1_R1105_U65, new_P1_R1105_U66,
    new_P1_R1105_U67, new_P1_R1105_U68, new_P1_R1105_U69, new_P1_R1105_U70,
    new_P1_R1105_U71, new_P1_R1105_U72, new_P1_R1105_U73, new_P1_R1105_U74,
    new_P1_R1105_U75, new_P1_R1105_U76, new_P1_R1105_U77, new_P1_R1105_U78,
    new_P1_R1105_U79, new_P1_R1105_U80, new_P1_R1105_U81, new_P1_R1105_U82,
    new_P1_R1105_U83, new_P1_R1105_U84, new_P1_R1105_U85, new_P1_R1105_U86,
    new_P1_R1105_U87, new_P1_R1105_U88, new_P1_R1105_U89, new_P1_R1105_U90,
    new_P1_R1105_U91, new_P1_R1105_U92, new_P1_R1105_U93, new_P1_R1105_U94,
    new_P1_R1105_U95, new_P1_R1105_U96, new_P1_R1105_U97, new_P1_R1105_U98,
    new_P1_R1105_U99, new_P1_R1105_U100, new_P1_R1105_U101,
    new_P1_R1105_U102, new_P1_R1105_U103, new_P1_R1105_U104,
    new_P1_R1105_U105, new_P1_R1105_U106, new_P1_R1105_U107,
    new_P1_R1105_U108, new_P1_R1105_U109, new_P1_R1105_U110,
    new_P1_R1105_U111, new_P1_R1105_U112, new_P1_R1105_U113,
    new_P1_R1105_U114, new_P1_R1105_U115, new_P1_R1105_U116,
    new_P1_R1105_U117, new_P1_R1105_U118, new_P1_R1105_U119,
    new_P1_R1105_U120, new_P1_R1105_U121, new_P1_R1105_U122,
    new_P1_R1105_U123, new_P1_R1105_U124, new_P1_R1105_U125,
    new_P1_R1105_U126, new_P1_R1105_U127, new_P1_R1105_U128,
    new_P1_R1105_U129, new_P1_R1105_U130, new_P1_R1105_U131,
    new_P1_R1105_U132, new_P1_R1105_U133, new_P1_R1105_U134,
    new_P1_R1105_U135, new_P1_R1105_U136, new_P1_R1105_U137,
    new_P1_R1105_U138, new_P1_R1105_U139, new_P1_R1105_U140,
    new_P1_R1105_U141, new_P1_R1105_U142, new_P1_R1105_U143,
    new_P1_R1105_U144, new_P1_R1105_U145, new_P1_R1105_U146,
    new_P1_R1105_U147, new_P1_R1105_U148, new_P1_R1105_U149,
    new_P1_R1105_U150, new_P1_R1105_U151, new_P1_R1105_U152,
    new_P1_R1105_U153, new_P1_R1105_U154, new_P1_R1105_U155,
    new_P1_R1105_U156, new_P1_R1105_U157, new_P1_R1105_U158,
    new_P1_R1105_U159, new_P1_R1105_U160, new_P1_R1105_U161,
    new_P1_R1105_U162, new_P1_R1105_U163, new_P1_R1105_U164,
    new_P1_R1105_U165, new_P1_R1105_U166, new_P1_R1105_U167,
    new_P1_R1105_U168, new_P1_R1105_U169, new_P1_R1105_U170,
    new_P1_R1105_U171, new_P1_R1105_U172, new_P1_R1105_U173,
    new_P1_R1105_U174, new_P1_R1105_U175, new_P1_R1105_U176,
    new_P1_R1105_U177, new_P1_R1105_U178, new_P1_R1105_U179,
    new_P1_R1105_U180, new_P1_R1105_U181, new_P1_R1105_U182,
    new_P1_R1105_U183, new_P1_R1105_U184, new_P1_R1105_U185,
    new_P1_R1105_U186, new_P1_R1105_U187, new_P1_R1105_U188,
    new_P1_R1105_U189, new_P1_R1105_U190, new_P1_R1105_U191,
    new_P1_R1105_U192, new_P1_R1105_U193, new_P1_R1105_U194,
    new_P1_R1105_U195, new_P1_R1105_U196, new_P1_R1105_U197,
    new_P1_R1105_U198, new_P1_R1105_U199, new_P1_R1105_U200,
    new_P1_R1105_U201, new_P1_R1105_U202, new_P1_R1105_U203,
    new_P1_R1105_U204, new_P1_R1105_U205, new_P1_R1105_U206,
    new_P1_R1105_U207, new_P1_R1105_U208, new_P1_R1105_U209,
    new_P1_R1105_U210, new_P1_R1105_U211, new_P1_R1105_U212,
    new_P1_R1105_U213, new_P1_R1105_U214, new_P1_R1105_U215,
    new_P1_R1105_U216, new_P1_R1105_U217, new_P1_R1105_U218,
    new_P1_R1105_U219, new_P1_R1105_U220, new_P1_R1105_U221,
    new_P1_R1105_U222, new_P1_R1105_U223, new_P1_R1105_U224,
    new_P1_R1105_U225, new_P1_R1105_U226, new_P1_R1105_U227,
    new_P1_R1105_U228, new_P1_R1105_U229, new_P1_R1105_U230,
    new_P1_R1105_U231, new_P1_R1105_U232, new_P1_R1105_U233,
    new_P1_R1105_U234, new_P1_R1105_U235, new_P1_R1105_U236,
    new_P1_R1105_U237, new_P1_R1105_U238, new_P1_R1105_U239,
    new_P1_R1105_U240, new_P1_R1105_U241, new_P1_R1105_U242,
    new_P1_R1105_U243, new_P1_R1105_U244, new_P1_R1105_U245,
    new_P1_R1105_U246, new_P1_R1105_U247, new_P1_R1105_U248,
    new_P1_R1105_U249, new_P1_R1105_U250, new_P1_R1105_U251,
    new_P1_R1105_U252, new_P1_R1105_U253, new_P1_R1105_U254,
    new_P1_R1105_U255, new_P1_R1105_U256, new_P1_R1105_U257,
    new_P1_R1105_U258, new_P1_R1105_U259, new_P1_R1105_U260,
    new_P1_R1105_U261, new_P1_R1105_U262, new_P1_R1105_U263,
    new_P1_R1105_U264, new_P1_R1105_U265, new_P1_R1105_U266,
    new_P1_R1105_U267, new_P1_R1105_U268, new_P1_R1105_U269,
    new_P1_R1105_U270, new_P1_R1105_U271, new_P1_R1105_U272,
    new_P1_R1105_U273, new_P1_R1105_U274, new_P1_R1105_U275,
    new_P1_R1105_U276, new_P1_R1105_U277, new_P1_R1105_U278,
    new_P1_R1105_U279, new_P1_R1105_U280, new_P1_R1105_U281,
    new_P1_R1105_U282, new_P1_R1105_U283, new_P1_R1105_U284,
    new_P1_R1105_U285, new_P1_R1105_U286, new_P1_R1105_U287,
    new_P1_R1105_U288, new_P1_R1105_U289, new_P1_R1105_U290,
    new_P1_R1105_U291, new_P1_R1105_U292, new_P1_R1105_U293,
    new_P1_R1105_U294, new_P1_R1105_U295, new_P1_R1105_U296,
    new_P1_R1105_U297, new_P1_R1105_U298, new_P1_R1105_U299,
    new_P1_R1105_U300, new_P1_R1105_U301, new_P1_R1105_U302,
    new_P1_R1105_U303, new_P1_R1105_U304, new_P1_R1105_U305,
    new_P1_R1105_U306, new_P1_R1105_U307, new_P1_R1105_U308,
    new_P1_SUB_88_U6, new_P1_SUB_88_U7, new_P1_SUB_88_U8, new_P1_SUB_88_U9,
    new_P1_SUB_88_U10, new_P1_SUB_88_U11, new_P1_SUB_88_U12,
    new_P1_SUB_88_U13, new_P1_SUB_88_U14, new_P1_SUB_88_U15,
    new_P1_SUB_88_U16, new_P1_SUB_88_U17, new_P1_SUB_88_U18,
    new_P1_SUB_88_U19, new_P1_SUB_88_U20, new_P1_SUB_88_U21,
    new_P1_SUB_88_U22, new_P1_SUB_88_U23, new_P1_SUB_88_U24,
    new_P1_SUB_88_U25, new_P1_SUB_88_U26, new_P1_SUB_88_U27,
    new_P1_SUB_88_U28, new_P1_SUB_88_U29, new_P1_SUB_88_U30,
    new_P1_SUB_88_U31, new_P1_SUB_88_U32, new_P1_SUB_88_U33,
    new_P1_SUB_88_U34, new_P1_SUB_88_U35, new_P1_SUB_88_U36,
    new_P1_SUB_88_U37, new_P1_SUB_88_U38, new_P1_SUB_88_U39,
    new_P1_SUB_88_U40, new_P1_SUB_88_U41, new_P1_SUB_88_U42,
    new_P1_SUB_88_U43, new_P1_SUB_88_U44, new_P1_SUB_88_U45,
    new_P1_SUB_88_U46, new_P1_SUB_88_U47, new_P1_SUB_88_U48,
    new_P1_SUB_88_U49, new_P1_SUB_88_U50, new_P1_SUB_88_U51,
    new_P1_SUB_88_U52, new_P1_SUB_88_U53, new_P1_SUB_88_U54,
    new_P1_SUB_88_U55, new_P1_SUB_88_U56, new_P1_SUB_88_U57,
    new_P1_SUB_88_U58, new_P1_SUB_88_U59, new_P1_SUB_88_U60,
    new_P1_SUB_88_U61, new_P1_SUB_88_U62, new_P1_SUB_88_U63,
    new_P1_SUB_88_U64, new_P1_SUB_88_U65, new_P1_SUB_88_U66,
    new_P1_SUB_88_U67, new_P1_SUB_88_U68, new_P1_SUB_88_U69,
    new_P1_SUB_88_U70, new_P1_SUB_88_U71, new_P1_SUB_88_U72,
    new_P1_SUB_88_U73, new_P1_SUB_88_U74, new_P1_SUB_88_U75,
    new_P1_SUB_88_U76, new_P1_SUB_88_U77, new_P1_SUB_88_U78,
    new_P1_SUB_88_U79, new_P1_SUB_88_U80, new_P1_SUB_88_U81,
    new_P1_SUB_88_U82, new_P1_SUB_88_U83, new_P1_SUB_88_U84,
    new_P1_SUB_88_U85, new_P1_SUB_88_U86, new_P1_SUB_88_U87,
    new_P1_SUB_88_U88, new_P1_SUB_88_U89, new_P1_SUB_88_U90,
    new_P1_SUB_88_U91, new_P1_SUB_88_U92, new_P1_SUB_88_U93,
    new_P1_SUB_88_U94, new_P1_SUB_88_U95, new_P1_SUB_88_U96,
    new_P1_SUB_88_U97, new_P1_SUB_88_U98, new_P1_SUB_88_U99,
    new_P1_SUB_88_U100, new_P1_SUB_88_U101, new_P1_SUB_88_U102,
    new_P1_SUB_88_U103, new_P1_SUB_88_U104, new_P1_SUB_88_U105,
    new_P1_SUB_88_U106, new_P1_SUB_88_U107, new_P1_SUB_88_U108,
    new_P1_SUB_88_U109, new_P1_SUB_88_U110, new_P1_SUB_88_U111,
    new_P1_SUB_88_U112, new_P1_SUB_88_U113, new_P1_SUB_88_U114,
    new_P1_SUB_88_U115, new_P1_SUB_88_U116, new_P1_SUB_88_U117,
    new_P1_SUB_88_U118, new_P1_SUB_88_U119, new_P1_SUB_88_U120,
    new_P1_SUB_88_U121, new_P1_SUB_88_U122, new_P1_SUB_88_U123,
    new_P1_SUB_88_U124, new_P1_SUB_88_U125, new_P1_SUB_88_U126,
    new_P1_SUB_88_U127, new_P1_SUB_88_U128, new_P1_SUB_88_U129,
    new_P1_SUB_88_U130, new_P1_SUB_88_U131, new_P1_SUB_88_U132,
    new_P1_SUB_88_U133, new_P1_SUB_88_U134, new_P1_SUB_88_U135,
    new_P1_SUB_88_U136, new_P1_SUB_88_U137, new_P1_SUB_88_U138,
    new_P1_SUB_88_U139, new_P1_SUB_88_U140, new_P1_SUB_88_U141,
    new_P1_SUB_88_U142, new_P1_SUB_88_U143, new_P1_SUB_88_U144,
    new_P1_SUB_88_U145, new_P1_SUB_88_U146, new_P1_SUB_88_U147,
    new_P1_SUB_88_U148, new_P1_SUB_88_U149, new_P1_SUB_88_U150,
    new_P1_SUB_88_U151, new_P1_SUB_88_U152, new_P1_SUB_88_U153,
    new_P1_SUB_88_U154, new_P1_SUB_88_U155, new_P1_SUB_88_U156,
    new_P1_SUB_88_U157, new_P1_SUB_88_U158, new_P1_SUB_88_U159,
    new_P1_SUB_88_U160, new_P1_SUB_88_U161, new_P1_SUB_88_U162,
    new_P1_SUB_88_U163, new_P1_SUB_88_U164, new_P1_SUB_88_U165,
    new_P1_SUB_88_U166, new_P1_SUB_88_U167, new_P1_SUB_88_U168,
    new_P1_SUB_88_U169, new_P1_SUB_88_U170, new_P1_SUB_88_U171,
    new_P1_SUB_88_U172, new_P1_SUB_88_U173, new_P1_SUB_88_U174,
    new_P1_SUB_88_U175, new_P1_SUB_88_U176, new_P1_SUB_88_U177,
    new_P1_SUB_88_U178, new_P1_SUB_88_U179, new_P1_SUB_88_U180,
    new_P1_SUB_88_U181, new_P1_SUB_88_U182, new_P1_SUB_88_U183,
    new_P1_SUB_88_U184, new_P1_SUB_88_U185, new_P1_SUB_88_U186,
    new_P1_SUB_88_U187, new_P1_SUB_88_U188, new_P1_SUB_88_U189,
    new_P1_SUB_88_U190, new_P1_SUB_88_U191, new_P1_SUB_88_U192,
    new_P1_SUB_88_U193, new_P1_SUB_88_U194, new_P1_SUB_88_U195,
    new_P1_SUB_88_U196, new_P1_SUB_88_U197, new_P1_SUB_88_U198,
    new_P1_SUB_88_U199, new_P1_SUB_88_U200, new_P1_SUB_88_U201,
    new_P1_SUB_88_U202, new_P1_SUB_88_U203, new_P1_SUB_88_U204,
    new_P1_SUB_88_U205, new_P1_SUB_88_U206, new_P1_SUB_88_U207,
    new_P1_SUB_88_U208, new_P1_SUB_88_U209, new_P1_SUB_88_U210,
    new_P1_SUB_88_U211, new_P1_SUB_88_U212, new_P1_SUB_88_U213,
    new_P1_SUB_88_U214, new_P1_SUB_88_U215, new_P1_SUB_88_U216,
    new_P1_SUB_88_U217, new_P1_SUB_88_U218, new_P1_SUB_88_U219,
    new_P1_SUB_88_U220, new_P1_SUB_88_U221, new_P1_SUB_88_U222,
    new_P1_SUB_88_U223, new_P1_SUB_88_U224, new_P1_SUB_88_U225,
    new_P1_SUB_88_U226, new_P1_SUB_88_U227, new_P1_SUB_88_U228,
    new_P1_SUB_88_U229, new_P1_SUB_88_U230, new_P1_SUB_88_U231,
    new_P1_SUB_88_U232, new_P1_SUB_88_U233, new_P1_SUB_88_U234,
    new_P1_SUB_88_U235, new_P1_SUB_88_U236, new_P1_SUB_88_U237,
    new_P1_SUB_88_U238, new_P1_SUB_88_U239, new_P1_SUB_88_U240,
    new_P1_SUB_88_U241, new_P1_SUB_88_U242, new_P1_SUB_88_U243,
    new_P1_SUB_88_U244, new_P1_SUB_88_U245, new_P1_SUB_88_U246,
    new_P1_SUB_88_U247, new_P1_SUB_88_U248, new_P1_SUB_88_U249,
    new_P1_SUB_88_U250, new_P1_SUB_88_U251, new_P1_R1309_U6,
    new_P1_R1309_U7, new_P1_R1309_U8, new_P1_R1309_U9, new_P1_R1309_U10,
    new_P1_R1282_U6, new_P1_R1282_U7, new_P1_R1282_U8, new_P1_R1282_U9,
    new_P1_R1282_U10, new_P1_R1282_U11, new_P1_R1282_U12, new_P1_R1282_U13,
    new_P1_R1282_U14, new_P1_R1282_U15, new_P1_R1282_U16, new_P1_R1282_U17,
    new_P1_R1282_U18, new_P1_R1282_U19, new_P1_R1282_U20, new_P1_R1282_U21,
    new_P1_R1282_U22, new_P1_R1282_U23, new_P1_R1282_U24, new_P1_R1282_U25,
    new_P1_R1282_U26, new_P1_R1282_U27, new_P1_R1282_U28, new_P1_R1282_U29,
    new_P1_R1282_U30, new_P1_R1282_U31, new_P1_R1282_U32, new_P1_R1282_U33,
    new_P1_R1282_U34, new_P1_R1282_U35, new_P1_R1282_U36, new_P1_R1282_U37,
    new_P1_R1282_U38, new_P1_R1282_U39, new_P1_R1282_U40, new_P1_R1282_U41,
    new_P1_R1282_U42, new_P1_R1282_U43, new_P1_R1282_U44, new_P1_R1282_U45,
    new_P1_R1282_U46, new_P1_R1282_U47, new_P1_R1282_U48, new_P1_R1282_U49,
    new_P1_R1282_U50, new_P1_R1282_U51, new_P1_R1282_U52, new_P1_R1282_U53,
    new_P1_R1282_U54, new_P1_R1282_U55, new_P1_R1282_U56, new_P1_R1282_U57,
    new_P1_R1282_U58, new_P1_R1282_U59, new_P1_R1282_U60, new_P1_R1282_U61,
    new_P1_R1282_U62, new_P1_R1282_U63, new_P1_R1282_U64, new_P1_R1282_U65,
    new_P1_R1282_U66, new_P1_R1282_U67, new_P1_R1282_U68, new_P1_R1282_U69,
    new_P1_R1282_U70, new_P1_R1282_U71, new_P1_R1282_U72, new_P1_R1282_U73,
    new_P1_R1282_U74, new_P1_R1282_U75, new_P1_R1282_U76, new_P1_R1282_U77,
    new_P1_R1282_U78, new_P1_R1282_U79, new_P1_R1282_U80, new_P1_R1282_U81,
    new_P1_R1282_U82, new_P1_R1282_U83, new_P1_R1282_U84, new_P1_R1282_U85,
    new_P1_R1282_U86, new_P1_R1282_U87, new_P1_R1282_U88, new_P1_R1282_U89,
    new_P1_R1282_U90, new_P1_R1282_U91, new_P1_R1282_U92, new_P1_R1282_U93,
    new_P1_R1282_U94, new_P1_R1282_U95, new_P1_R1282_U96, new_P1_R1282_U97,
    new_P1_R1282_U98, new_P1_R1282_U99, new_P1_R1282_U100,
    new_P1_R1282_U101, new_P1_R1282_U102, new_P1_R1282_U103,
    new_P1_R1282_U104, new_P1_R1282_U105, new_P1_R1282_U106,
    new_P1_R1282_U107, new_P1_R1282_U108, new_P1_R1282_U109,
    new_P1_R1282_U110, new_P1_R1282_U111, new_P1_R1282_U112,
    new_P1_R1282_U113, new_P1_R1282_U114, new_P1_R1282_U115,
    new_P1_R1282_U116, new_P1_R1282_U117, new_P1_R1282_U118,
    new_P1_R1282_U119, new_P1_R1282_U120, new_P1_R1282_U121,
    new_P1_R1282_U122, new_P1_R1282_U123, new_P1_R1282_U124,
    new_P1_R1282_U125, new_P1_R1282_U126, new_P1_R1282_U127,
    new_P1_R1282_U128, new_P1_R1282_U129, new_P1_R1282_U130,
    new_P1_R1282_U131, new_P1_R1282_U132, new_P1_R1282_U133,
    new_P1_R1282_U134, new_P1_R1282_U135, new_P1_R1282_U136,
    new_P1_R1282_U137, new_P1_R1282_U138, new_P1_R1282_U139,
    new_P1_R1282_U140, new_P1_R1282_U141, new_P1_R1282_U142,
    new_P1_R1282_U143, new_P1_R1282_U144, new_P1_R1282_U145,
    new_P1_R1282_U146, new_P1_R1282_U147, new_P1_R1282_U148,
    new_P1_R1282_U149, new_P1_R1282_U150, new_P1_R1282_U151,
    new_P1_R1282_U152, new_P1_R1282_U153, new_P1_R1282_U154,
    new_P1_R1282_U155, new_P1_R1282_U156, new_P1_R1282_U157,
    new_P1_R1282_U158, new_P1_R1282_U159, new_P1_R1240_U4, new_P1_R1240_U5,
    new_P1_R1240_U6, new_P1_R1240_U7, new_P1_R1240_U8, new_P1_R1240_U9,
    new_P1_R1240_U10, new_P1_R1240_U11, new_P1_R1240_U12, new_P1_R1240_U13,
    new_P1_R1240_U14, new_P1_R1240_U15, new_P1_R1240_U16, new_P1_R1240_U17,
    new_P1_R1240_U18, new_P1_R1240_U19, new_P1_R1240_U20, new_P1_R1240_U21,
    new_P1_R1240_U22, new_P1_R1240_U23, new_P1_R1240_U24, new_P1_R1240_U25,
    new_P1_R1240_U26, new_P1_R1240_U27, new_P1_R1240_U28, new_P1_R1240_U29,
    new_P1_R1240_U30, new_P1_R1240_U31, new_P1_R1240_U32, new_P1_R1240_U33,
    new_P1_R1240_U34, new_P1_R1240_U35, new_P1_R1240_U36, new_P1_R1240_U37,
    new_P1_R1240_U38, new_P1_R1240_U39, new_P1_R1240_U40, new_P1_R1240_U41,
    new_P1_R1240_U42, new_P1_R1240_U43, new_P1_R1240_U44, new_P1_R1240_U45,
    new_P1_R1240_U46, new_P1_R1240_U47, new_P1_R1240_U48, new_P1_R1240_U49,
    new_P1_R1240_U50, new_P1_R1240_U51, new_P1_R1240_U52, new_P1_R1240_U53,
    new_P1_R1240_U54, new_P1_R1240_U55, new_P1_R1240_U56, new_P1_R1240_U57,
    new_P1_R1240_U58, new_P1_R1240_U59, new_P1_R1240_U60, new_P1_R1240_U61,
    new_P1_R1240_U62, new_P1_R1240_U63, new_P1_R1240_U64, new_P1_R1240_U65,
    new_P1_R1240_U66, new_P1_R1240_U67, new_P1_R1240_U68, new_P1_R1240_U69,
    new_P1_R1240_U70, new_P1_R1240_U71, new_P1_R1240_U72, new_P1_R1240_U73,
    new_P1_R1240_U74, new_P1_R1240_U75, new_P1_R1240_U76, new_P1_R1240_U77,
    new_P1_R1240_U78, new_P1_R1240_U79, new_P1_R1240_U80, new_P1_R1240_U81,
    new_P1_R1240_U82, new_P1_R1240_U83, new_P1_R1240_U84, new_P1_R1240_U85,
    new_P1_R1240_U86, new_P1_R1240_U87, new_P1_R1240_U88, new_P1_R1240_U89,
    new_P1_R1240_U90, new_P1_R1240_U91, new_P1_R1240_U92, new_P1_R1240_U93,
    new_P1_R1240_U94, new_P1_R1240_U95, new_P1_R1240_U96, new_P1_R1240_U97,
    new_P1_R1240_U98, new_P1_R1240_U99, new_P1_R1240_U100,
    new_P1_R1240_U101, new_P1_R1240_U102, new_P1_R1240_U103,
    new_P1_R1240_U104, new_P1_R1240_U105, new_P1_R1240_U106,
    new_P1_R1240_U107, new_P1_R1240_U108, new_P1_R1240_U109,
    new_P1_R1240_U110, new_P1_R1240_U111, new_P1_R1240_U112,
    new_P1_R1240_U113, new_P1_R1240_U114, new_P1_R1240_U115,
    new_P1_R1240_U116, new_P1_R1240_U117, new_P1_R1240_U118,
    new_P1_R1240_U119, new_P1_R1240_U120, new_P1_R1240_U121,
    new_P1_R1240_U122, new_P1_R1240_U123, new_P1_R1240_U124,
    new_P1_R1240_U125, new_P1_R1240_U126, new_P1_R1240_U127,
    new_P1_R1240_U128, new_P1_R1240_U129, new_P1_R1240_U130,
    new_P1_R1240_U131, new_P1_R1240_U132, new_P1_R1240_U133,
    new_P1_R1240_U134, new_P1_R1240_U135, new_P1_R1240_U136,
    new_P1_R1240_U137, new_P1_R1240_U138, new_P1_R1240_U139,
    new_P1_R1240_U140, new_P1_R1240_U141, new_P1_R1240_U142,
    new_P1_R1240_U143, new_P1_R1240_U144, new_P1_R1240_U145,
    new_P1_R1240_U146, new_P1_R1240_U147, new_P1_R1240_U148,
    new_P1_R1240_U149, new_P1_R1240_U150, new_P1_R1240_U151,
    new_P1_R1240_U152, new_P1_R1240_U153, new_P1_R1240_U154,
    new_P1_R1240_U155, new_P1_R1240_U156, new_P1_R1240_U157,
    new_P1_R1240_U158, new_P1_R1240_U159, new_P1_R1240_U160,
    new_P1_R1240_U161, new_P1_R1240_U162, new_P1_R1240_U163,
    new_P1_R1240_U164, new_P1_R1240_U165, new_P1_R1240_U166,
    new_P1_R1240_U167, new_P1_R1240_U168, new_P1_R1240_U169,
    new_P1_R1240_U170, new_P1_R1240_U171, new_P1_R1240_U172,
    new_P1_R1240_U173, new_P1_R1240_U174, new_P1_R1240_U175,
    new_P1_R1240_U176, new_P1_R1240_U177, new_P1_R1240_U178,
    new_P1_R1240_U179, new_P1_R1240_U180, new_P1_R1240_U181,
    new_P1_R1240_U182, new_P1_R1240_U183, new_P1_R1240_U184,
    new_P1_R1240_U185, new_P1_R1240_U186, new_P1_R1240_U187,
    new_P1_R1240_U188, new_P1_R1240_U189, new_P1_R1240_U190,
    new_P1_R1240_U191, new_P1_R1240_U192, new_P1_R1240_U193,
    new_P1_R1240_U194, new_P1_R1240_U195, new_P1_R1240_U196,
    new_P1_R1240_U197, new_P1_R1240_U198, new_P1_R1240_U199,
    new_P1_R1240_U200, new_P1_R1240_U201, new_P1_R1240_U202,
    new_P1_R1240_U203, new_P1_R1240_U204, new_P1_R1240_U205,
    new_P1_R1240_U206, new_P1_R1240_U207, new_P1_R1240_U208,
    new_P1_R1240_U209, new_P1_R1240_U210, new_P1_R1240_U211,
    new_P1_R1240_U212, new_P1_R1240_U213, new_P1_R1240_U214,
    new_P1_R1240_U215, new_P1_R1240_U216, new_P1_R1240_U217,
    new_P1_R1240_U218, new_P1_R1240_U219, new_P1_R1240_U220,
    new_P1_R1240_U221, new_P1_R1240_U222, new_P1_R1240_U223,
    new_P1_R1240_U224, new_P1_R1240_U225, new_P1_R1240_U226,
    new_P1_R1240_U227, new_P1_R1240_U228, new_P1_R1240_U229,
    new_P1_R1240_U230, new_P1_R1240_U231, new_P1_R1240_U232,
    new_P1_R1240_U233, new_P1_R1240_U234, new_P1_R1240_U235,
    new_P1_R1240_U236, new_P1_R1240_U237, new_P1_R1240_U238,
    new_P1_R1240_U239, new_P1_R1240_U240, new_P1_R1240_U241,
    new_P1_R1240_U242, new_P1_R1240_U243, new_P1_R1240_U244,
    new_P1_R1240_U245, new_P1_R1240_U246, new_P1_R1240_U247,
    new_P1_R1240_U248, new_P1_R1240_U249, new_P1_R1240_U250,
    new_P1_R1240_U251, new_P1_R1240_U252, new_P1_R1240_U253,
    new_P1_R1240_U254, new_P1_R1240_U255, new_P1_R1240_U256,
    new_P1_R1240_U257, new_P1_R1240_U258, new_P1_R1240_U259,
    new_P1_R1240_U260, new_P1_R1240_U261, new_P1_R1240_U262,
    new_P1_R1240_U263, new_P1_R1240_U264, new_P1_R1240_U265,
    new_P1_R1240_U266, new_P1_R1240_U267, new_P1_R1240_U268,
    new_P1_R1240_U269, new_P1_R1240_U270, new_P1_R1240_U271,
    new_P1_R1240_U272, new_P1_R1240_U273, new_P1_R1240_U274,
    new_P1_R1240_U275, new_P1_R1240_U276, new_P1_R1240_U277,
    new_P1_R1240_U278, new_P1_R1240_U279, new_P1_R1240_U280,
    new_P1_R1240_U281, new_P1_R1240_U282, new_P1_R1240_U283,
    new_P1_R1240_U284, new_P1_R1240_U285, new_P1_R1240_U286,
    new_P1_R1240_U287, new_P1_R1240_U288, new_P1_R1240_U289,
    new_P1_R1240_U290, new_P1_R1240_U291, new_P1_R1240_U292,
    new_P1_R1240_U293, new_P1_R1240_U294, new_P1_R1240_U295,
    new_P1_R1240_U296, new_P1_R1240_U297, new_P1_R1240_U298,
    new_P1_R1240_U299, new_P1_R1240_U300, new_P1_R1240_U301,
    new_P1_R1240_U302, new_P1_R1240_U303, new_P1_R1240_U304,
    new_P1_R1240_U305, new_P1_R1240_U306, new_P1_R1240_U307,
    new_P1_R1240_U308, new_P1_R1240_U309, new_P1_R1240_U310,
    new_P1_R1240_U311, new_P1_R1240_U312, new_P1_R1240_U313,
    new_P1_R1240_U314, new_P1_R1240_U315, new_P1_R1240_U316,
    new_P1_R1240_U317, new_P1_R1240_U318, new_P1_R1240_U319,
    new_P1_R1240_U320, new_P1_R1240_U321, new_P1_R1240_U322,
    new_P1_R1240_U323, new_P1_R1240_U324, new_P1_R1240_U325,
    new_P1_R1240_U326, new_P1_R1240_U327, new_P1_R1240_U328,
    new_P1_R1240_U329, new_P1_R1240_U330, new_P1_R1240_U331,
    new_P1_R1240_U332, new_P1_R1240_U333, new_P1_R1240_U334,
    new_P1_R1240_U335, new_P1_R1240_U336, new_P1_R1240_U337,
    new_P1_R1240_U338, new_P1_R1240_U339, new_P1_R1240_U340,
    new_P1_R1240_U341, new_P1_R1240_U342, new_P1_R1240_U343,
    new_P1_R1240_U344, new_P1_R1240_U345, new_P1_R1240_U346,
    new_P1_R1240_U347, new_P1_R1240_U348, new_P1_R1240_U349,
    new_P1_R1240_U350, new_P1_R1240_U351, new_P1_R1240_U352,
    new_P1_R1240_U353, new_P1_R1240_U354, new_P1_R1240_U355,
    new_P1_R1240_U356, new_P1_R1240_U357, new_P1_R1240_U358,
    new_P1_R1240_U359, new_P1_R1240_U360, new_P1_R1240_U361,
    new_P1_R1240_U362, new_P1_R1240_U363, new_P1_R1240_U364,
    new_P1_R1240_U365, new_P1_R1240_U366, new_P1_R1240_U367,
    new_P1_R1240_U368, new_P1_R1240_U369, new_P1_R1240_U370,
    new_P1_R1240_U371, new_P1_R1240_U372, new_P1_R1240_U373,
    new_P1_R1240_U374, new_P1_R1240_U375, new_P1_R1240_U376,
    new_P1_R1240_U377, new_P1_R1240_U378, new_P1_R1240_U379,
    new_P1_R1240_U380, new_P1_R1240_U381, new_P1_R1240_U382,
    new_P1_R1240_U383, new_P1_R1240_U384, new_P1_R1240_U385,
    new_P1_R1240_U386, new_P1_R1240_U387, new_P1_R1240_U388,
    new_P1_R1240_U389, new_P1_R1240_U390, new_P1_R1240_U391,
    new_P1_R1240_U392, new_P1_R1240_U393, new_P1_R1240_U394,
    new_P1_R1240_U395, new_P1_R1240_U396, new_P1_R1240_U397,
    new_P1_R1240_U398, new_P1_R1240_U399, new_P1_R1240_U400,
    new_P1_R1240_U401, new_P1_R1240_U402, new_P1_R1240_U403,
    new_P1_R1240_U404, new_P1_R1240_U405, new_P1_R1240_U406,
    new_P1_R1240_U407, new_P1_R1240_U408, new_P1_R1240_U409,
    new_P1_R1240_U410, new_P1_R1240_U411, new_P1_R1240_U412,
    new_P1_R1240_U413, new_P1_R1240_U414, new_P1_R1240_U415,
    new_P1_R1240_U416, new_P1_R1240_U417, new_P1_R1240_U418,
    new_P1_R1240_U419, new_P1_R1240_U420, new_P1_R1240_U421,
    new_P1_R1240_U422, new_P1_R1240_U423, new_P1_R1240_U424,
    new_P1_R1240_U425, new_P1_R1240_U426, new_P1_R1240_U427,
    new_P1_R1240_U428, new_P1_R1240_U429, new_P1_R1240_U430,
    new_P1_R1240_U431, new_P1_R1240_U432, new_P1_R1240_U433,
    new_P1_R1240_U434, new_P1_R1240_U435, new_P1_R1240_U436,
    new_P1_R1240_U437, new_P1_R1240_U438, new_P1_R1240_U439,
    new_P1_R1240_U440, new_P1_R1240_U441, new_P1_R1240_U442,
    new_P1_R1240_U443, new_P1_R1240_U444, new_P1_R1240_U445,
    new_P1_R1240_U446, new_P1_R1240_U447, new_P1_R1240_U448,
    new_P1_R1240_U449, new_P1_R1240_U450, new_P1_R1240_U451,
    new_P1_R1240_U452, new_P1_R1240_U453, new_P1_R1240_U454,
    new_P1_R1240_U455, new_P1_R1240_U456, new_P1_R1240_U457,
    new_P1_R1240_U458, new_P1_R1240_U459, new_P1_R1240_U460,
    new_P1_R1240_U461, new_P1_R1240_U462, new_P1_R1240_U463,
    new_P1_R1240_U464, new_P1_R1240_U465, new_P1_R1240_U466,
    new_P1_R1240_U467, new_P1_R1240_U468, new_P1_R1240_U469,
    new_P1_R1240_U470, new_P1_R1240_U471, new_P1_R1240_U472,
    new_P1_R1240_U473, new_P1_R1240_U474, new_P1_R1240_U475,
    new_P1_R1240_U476, new_P1_R1240_U477, new_P1_R1240_U478,
    new_P1_R1240_U479, new_P1_R1240_U480, new_P1_R1240_U481,
    new_P1_R1240_U482, new_P1_R1240_U483, new_P1_R1240_U484,
    new_P1_R1240_U485, new_P1_R1240_U486, new_P1_R1240_U487,
    new_P1_R1240_U488, new_P1_R1240_U489, new_P1_R1240_U490,
    new_P1_R1240_U491, new_P1_R1240_U492, new_P1_R1240_U493,
    new_P1_R1240_U494, new_P1_R1240_U495, new_P1_R1240_U496,
    new_P1_R1240_U497, new_P1_R1240_U498, new_P1_R1240_U499,
    new_P1_R1240_U500, new_P1_R1240_U501, new_P1_R1162_U4, new_P1_R1162_U5,
    new_P1_R1162_U6, new_P1_R1162_U7, new_P1_R1162_U8, new_P1_R1162_U9,
    new_P1_R1162_U10, new_P1_R1162_U11, new_P1_R1162_U12, new_P1_R1162_U13,
    new_P1_R1162_U14, new_P1_R1162_U15, new_P1_R1162_U16, new_P1_R1162_U17,
    new_P1_R1162_U18, new_P1_R1162_U19, new_P1_R1162_U20, new_P1_R1162_U21,
    new_P1_R1162_U22, new_P1_R1162_U23, new_P1_R1162_U24, new_P1_R1162_U25,
    new_P1_R1162_U26, new_P1_R1162_U27, new_P1_R1162_U28, new_P1_R1162_U29,
    new_P1_R1162_U30, new_P1_R1162_U31, new_P1_R1162_U32, new_P1_R1162_U33,
    new_P1_R1162_U34, new_P1_R1162_U35, new_P1_R1162_U36, new_P1_R1162_U37,
    new_P1_R1162_U38, new_P1_R1162_U39, new_P1_R1162_U40, new_P1_R1162_U41,
    new_P1_R1162_U42, new_P1_R1162_U43, new_P1_R1162_U44, new_P1_R1162_U45,
    new_P1_R1162_U46, new_P1_R1162_U47, new_P1_R1162_U48, new_P1_R1162_U49,
    new_P1_R1162_U50, new_P1_R1162_U51, new_P1_R1162_U52, new_P1_R1162_U53,
    new_P1_R1162_U54, new_P1_R1162_U55, new_P1_R1162_U56, new_P1_R1162_U57,
    new_P1_R1162_U58, new_P1_R1162_U59, new_P1_R1162_U60, new_P1_R1162_U61,
    new_P1_R1162_U62, new_P1_R1162_U63, new_P1_R1162_U64, new_P1_R1162_U65,
    new_P1_R1162_U66, new_P1_R1162_U67, new_P1_R1162_U68, new_P1_R1162_U69,
    new_P1_R1162_U70, new_P1_R1162_U71, new_P1_R1162_U72, new_P1_R1162_U73,
    new_P1_R1162_U74, new_P1_R1162_U75, new_P1_R1162_U76, new_P1_R1162_U77,
    new_P1_R1162_U78, new_P1_R1162_U79, new_P1_R1162_U80, new_P1_R1162_U81,
    new_P1_R1162_U82, new_P1_R1162_U83, new_P1_R1162_U84, new_P1_R1162_U85,
    new_P1_R1162_U86, new_P1_R1162_U87, new_P1_R1162_U88, new_P1_R1162_U89,
    new_P1_R1162_U90, new_P1_R1162_U91, new_P1_R1162_U92, new_P1_R1162_U93,
    new_P1_R1162_U94, new_P1_R1162_U95, new_P1_R1162_U96, new_P1_R1162_U97,
    new_P1_R1162_U98, new_P1_R1162_U99, new_P1_R1162_U100,
    new_P1_R1162_U101, new_P1_R1162_U102, new_P1_R1162_U103,
    new_P1_R1162_U104, new_P1_R1162_U105, new_P1_R1162_U106,
    new_P1_R1162_U107, new_P1_R1162_U108, new_P1_R1162_U109,
    new_P1_R1162_U110, new_P1_R1162_U111, new_P1_R1162_U112,
    new_P1_R1162_U113, new_P1_R1162_U114, new_P1_R1162_U115,
    new_P1_R1162_U116, new_P1_R1162_U117, new_P1_R1162_U118,
    new_P1_R1162_U119, new_P1_R1162_U120, new_P1_R1162_U121,
    new_P1_R1162_U122, new_P1_R1162_U123, new_P1_R1162_U124,
    new_P1_R1162_U125, new_P1_R1162_U126, new_P1_R1162_U127,
    new_P1_R1162_U128, new_P1_R1162_U129, new_P1_R1162_U130,
    new_P1_R1162_U131, new_P1_R1162_U132, new_P1_R1162_U133,
    new_P1_R1162_U134, new_P1_R1162_U135, new_P1_R1162_U136,
    new_P1_R1162_U137, new_P1_R1162_U138, new_P1_R1162_U139,
    new_P1_R1162_U140, new_P1_R1162_U141, new_P1_R1162_U142,
    new_P1_R1162_U143, new_P1_R1162_U144, new_P1_R1162_U145,
    new_P1_R1162_U146, new_P1_R1162_U147, new_P1_R1162_U148,
    new_P1_R1162_U149, new_P1_R1162_U150, new_P1_R1162_U151,
    new_P1_R1162_U152, new_P1_R1162_U153, new_P1_R1162_U154,
    new_P1_R1162_U155, new_P1_R1162_U156, new_P1_R1162_U157,
    new_P1_R1162_U158, new_P1_R1162_U159, new_P1_R1162_U160,
    new_P1_R1162_U161, new_P1_R1162_U162, new_P1_R1162_U163,
    new_P1_R1162_U164, new_P1_R1162_U165, new_P1_R1162_U166,
    new_P1_R1162_U167, new_P1_R1162_U168, new_P1_R1162_U169,
    new_P1_R1162_U170, new_P1_R1162_U171, new_P1_R1162_U172,
    new_P1_R1162_U173, new_P1_R1162_U174, new_P1_R1162_U175,
    new_P1_R1162_U176, new_P1_R1162_U177, new_P1_R1162_U178,
    new_P1_R1162_U179, new_P1_R1162_U180, new_P1_R1162_U181,
    new_P1_R1162_U182, new_P1_R1162_U183, new_P1_R1162_U184,
    new_P1_R1162_U185, new_P1_R1162_U186, new_P1_R1162_U187,
    new_P1_R1162_U188, new_P1_R1162_U189, new_P1_R1162_U190,
    new_P1_R1162_U191, new_P1_R1162_U192, new_P1_R1162_U193,
    new_P1_R1162_U194, new_P1_R1162_U195, new_P1_R1162_U196,
    new_P1_R1162_U197, new_P1_R1162_U198, new_P1_R1162_U199,
    new_P1_R1162_U200, new_P1_R1162_U201, new_P1_R1162_U202,
    new_P1_R1162_U203, new_P1_R1162_U204, new_P1_R1162_U205,
    new_P1_R1162_U206, new_P1_R1162_U207, new_P1_R1162_U208,
    new_P1_R1162_U209, new_P1_R1162_U210, new_P1_R1162_U211,
    new_P1_R1162_U212, new_P1_R1162_U213, new_P1_R1162_U214,
    new_P1_R1162_U215, new_P1_R1162_U216, new_P1_R1162_U217,
    new_P1_R1162_U218, new_P1_R1162_U219, new_P1_R1162_U220,
    new_P1_R1162_U221, new_P1_R1162_U222, new_P1_R1162_U223,
    new_P1_R1162_U224, new_P1_R1162_U225, new_P1_R1162_U226,
    new_P1_R1162_U227, new_P1_R1162_U228, new_P1_R1162_U229,
    new_P1_R1162_U230, new_P1_R1162_U231, new_P1_R1162_U232,
    new_P1_R1162_U233, new_P1_R1162_U234, new_P1_R1162_U235,
    new_P1_R1162_U236, new_P1_R1162_U237, new_P1_R1162_U238,
    new_P1_R1162_U239, new_P1_R1162_U240, new_P1_R1162_U241,
    new_P1_R1162_U242, new_P1_R1162_U243, new_P1_R1162_U244,
    new_P1_R1162_U245, new_P1_R1162_U246, new_P1_R1162_U247,
    new_P1_R1162_U248, new_P1_R1162_U249, new_P1_R1162_U250,
    new_P1_R1162_U251, new_P1_R1162_U252, new_P1_R1162_U253,
    new_P1_R1162_U254, new_P1_R1162_U255, new_P1_R1162_U256,
    new_P1_R1162_U257, new_P1_R1162_U258, new_P1_R1162_U259,
    new_P1_R1162_U260, new_P1_R1162_U261, new_P1_R1162_U262,
    new_P1_R1162_U263, new_P1_R1162_U264, new_P1_R1162_U265,
    new_P1_R1162_U266, new_P1_R1162_U267, new_P1_R1162_U268,
    new_P1_R1162_U269, new_P1_R1162_U270, new_P1_R1162_U271,
    new_P1_R1162_U272, new_P1_R1162_U273, new_P1_R1162_U274,
    new_P1_R1162_U275, new_P1_R1162_U276, new_P1_R1162_U277,
    new_P1_R1162_U278, new_P1_R1162_U279, new_P1_R1162_U280,
    new_P1_R1162_U281, new_P1_R1162_U282, new_P1_R1162_U283,
    new_P1_R1162_U284, new_P1_R1162_U285, new_P1_R1162_U286,
    new_P1_R1162_U287, new_P1_R1162_U288, new_P1_R1162_U289,
    new_P1_R1162_U290, new_P1_R1162_U291, new_P1_R1162_U292,
    new_P1_R1162_U293, new_P1_R1162_U294, new_P1_R1162_U295,
    new_P1_R1162_U296, new_P1_R1162_U297, new_P1_R1162_U298,
    new_P1_R1162_U299, new_P1_R1162_U300, new_P1_R1162_U301,
    new_P1_R1162_U302, new_P1_R1162_U303, new_P1_R1162_U304,
    new_P1_R1162_U305, new_P1_R1162_U306, new_P1_R1162_U307,
    new_P1_R1162_U308, new_P1_R1117_U6, new_P1_R1117_U7, new_P1_R1117_U8,
    new_P1_R1117_U9, new_P1_R1117_U10, new_P1_R1117_U11, new_P1_R1117_U12,
    new_P1_R1117_U13, new_P1_R1117_U14, new_P1_R1117_U15, new_P1_R1117_U16,
    new_P1_R1117_U17, new_P1_R1117_U18, new_P1_R1117_U19, new_P1_R1117_U20,
    new_P1_R1117_U21, new_P1_R1117_U22, new_P1_R1117_U23, new_P1_R1117_U24,
    new_P1_R1117_U25, new_P1_R1117_U26, new_P1_R1117_U27, new_P1_R1117_U28,
    new_P1_R1117_U29, new_P1_R1117_U30, new_P1_R1117_U31, new_P1_R1117_U32,
    new_P1_R1117_U33, new_P1_R1117_U34, new_P1_R1117_U35, new_P1_R1117_U36,
    new_P1_R1117_U37, new_P1_R1117_U38, new_P1_R1117_U39, new_P1_R1117_U40,
    new_P1_R1117_U41, new_P1_R1117_U42, new_P1_R1117_U43, new_P1_R1117_U44,
    new_P1_R1117_U45, new_P1_R1117_U46, new_P1_R1117_U47, new_P1_R1117_U48,
    new_P1_R1117_U49, new_P1_R1117_U50, new_P1_R1117_U51, new_P1_R1117_U52,
    new_P1_R1117_U53, new_P1_R1117_U54, new_P1_R1117_U55, new_P1_R1117_U56,
    new_P1_R1117_U57, new_P1_R1117_U58, new_P1_R1117_U59, new_P1_R1117_U60,
    new_P1_R1117_U61, new_P1_R1117_U62, new_P1_R1117_U63, new_P1_R1117_U64,
    new_P1_R1117_U65, new_P1_R1117_U66, new_P1_R1117_U67, new_P1_R1117_U68,
    new_P1_R1117_U69, new_P1_R1117_U70, new_P1_R1117_U71, new_P1_R1117_U72,
    new_P1_R1117_U73, new_P1_R1117_U74, new_P1_R1117_U75, new_P1_R1117_U76,
    new_P1_R1117_U77, new_P1_R1117_U78, new_P1_R1117_U79, new_P1_R1117_U80,
    new_P1_R1117_U81, new_P1_R1117_U82, new_P1_R1117_U83, new_P1_R1117_U84,
    new_P1_R1117_U85, new_P1_R1117_U86, new_P1_R1117_U87, new_P1_R1117_U88,
    new_P1_R1117_U89, new_P1_R1117_U90, new_P1_R1117_U91, new_P1_R1117_U92,
    new_P1_R1117_U93, new_P1_R1117_U94, new_P1_R1117_U95, new_P1_R1117_U96,
    new_P1_R1117_U97, new_P1_R1117_U98, new_P1_R1117_U99,
    new_P1_R1117_U100, new_P1_R1117_U101, new_P1_R1117_U102,
    new_P1_R1117_U103, new_P1_R1117_U104, new_P1_R1117_U105,
    new_P1_R1117_U106, new_P1_R1117_U107, new_P1_R1117_U108,
    new_P1_R1117_U109, new_P1_R1117_U110, new_P1_R1117_U111,
    new_P1_R1117_U112, new_P1_R1117_U113, new_P1_R1117_U114,
    new_P1_R1117_U115, new_P1_R1117_U116, new_P1_R1117_U117,
    new_P1_R1117_U118, new_P1_R1117_U119, new_P1_R1117_U120,
    new_P1_R1117_U121, new_P1_R1117_U122, new_P1_R1117_U123,
    new_P1_R1117_U124, new_P1_R1117_U125, new_P1_R1117_U126,
    new_P1_R1117_U127, new_P1_R1117_U128, new_P1_R1117_U129,
    new_P1_R1117_U130, new_P1_R1117_U131, new_P1_R1117_U132,
    new_P1_R1117_U133, new_P1_R1117_U134, new_P1_R1117_U135,
    new_P1_R1117_U136, new_P1_R1117_U137, new_P1_R1117_U138,
    new_P1_R1117_U139, new_P1_R1117_U140, new_P1_R1117_U141,
    new_P1_R1117_U142, new_P1_R1117_U143, new_P1_R1117_U144,
    new_P1_R1117_U145, new_P1_R1117_U146, new_P1_R1117_U147,
    new_P1_R1117_U148, new_P1_R1117_U149, new_P1_R1117_U150,
    new_P1_R1117_U151, new_P1_R1117_U152, new_P1_R1117_U153,
    new_P1_R1117_U154, new_P1_R1117_U155, new_P1_R1117_U156,
    new_P1_R1117_U157, new_P1_R1117_U158, new_P1_R1117_U159,
    new_P1_R1117_U160, new_P1_R1117_U161, new_P1_R1117_U162,
    new_P1_R1117_U163, new_P1_R1117_U164, new_P1_R1117_U165,
    new_P1_R1117_U166, new_P1_R1117_U167, new_P1_R1117_U168,
    new_P1_R1117_U169, new_P1_R1117_U170, new_P1_R1117_U171,
    new_P1_R1117_U172, new_P1_R1117_U173, new_P1_R1117_U174,
    new_P1_R1117_U175, new_P1_R1117_U176, new_P1_R1117_U177,
    new_P1_R1117_U178, new_P1_R1117_U179, new_P1_R1117_U180,
    new_P1_R1117_U181, new_P1_R1117_U182, new_P1_R1117_U183,
    new_P1_R1117_U184, new_P1_R1117_U185, new_P1_R1117_U186,
    new_P1_R1117_U187, new_P1_R1117_U188, new_P1_R1117_U189,
    new_P1_R1117_U190, new_P1_R1117_U191, new_P1_R1117_U192,
    new_P1_R1117_U193, new_P1_R1117_U194, new_P1_R1117_U195,
    new_P1_R1117_U196, new_P1_R1117_U197, new_P1_R1117_U198,
    new_P1_R1117_U199, new_P1_R1117_U200, new_P1_R1117_U201,
    new_P1_R1117_U202, new_P1_R1117_U203, new_P1_R1117_U204,
    new_P1_R1117_U205, new_P1_R1117_U206, new_P1_R1117_U207,
    new_P1_R1117_U208, new_P1_R1117_U209, new_P1_R1117_U210,
    new_P1_R1117_U211, new_P1_R1117_U212, new_P1_R1117_U213,
    new_P1_R1117_U214, new_P1_R1117_U215, new_P1_R1117_U216,
    new_P1_R1117_U217, new_P1_R1117_U218, new_P1_R1117_U219,
    new_P1_R1117_U220, new_P1_R1117_U221, new_P1_R1117_U222,
    new_P1_R1117_U223, new_P1_R1117_U224, new_P1_R1117_U225,
    new_P1_R1117_U226, new_P1_R1117_U227, new_P1_R1117_U228,
    new_P1_R1117_U229, new_P1_R1117_U230, new_P1_R1117_U231,
    new_P1_R1117_U232, new_P1_R1117_U233, new_P1_R1117_U234,
    new_P1_R1117_U235, new_P1_R1117_U236, new_P1_R1117_U237,
    new_P1_R1117_U238, new_P1_R1117_U239, new_P1_R1117_U240,
    new_P1_R1117_U241, new_P1_R1117_U242, new_P1_R1117_U243,
    new_P1_R1117_U244, new_P1_R1117_U245, new_P1_R1117_U246,
    new_P1_R1117_U247, new_P1_R1117_U248, new_P1_R1117_U249,
    new_P1_R1117_U250, new_P1_R1117_U251, new_P1_R1117_U252,
    new_P1_R1117_U253, new_P1_R1117_U254, new_P1_R1117_U255,
    new_P1_R1117_U256, new_P1_R1117_U257, new_P1_R1117_U258,
    new_P1_R1117_U259, new_P1_R1117_U260, new_P1_R1117_U261,
    new_P1_R1117_U262, new_P1_R1117_U263, new_P1_R1117_U264,
    new_P1_R1117_U265, new_P1_R1117_U266, new_P1_R1117_U267,
    new_P1_R1117_U268, new_P1_R1117_U269, new_P1_R1117_U270,
    new_P1_R1117_U271, new_P1_R1117_U272, new_P1_R1117_U273,
    new_P1_R1117_U274, new_P1_R1117_U275, new_P1_R1117_U276,
    new_P1_R1117_U277, new_P1_R1117_U278, new_P1_R1117_U279,
    new_P1_R1117_U280, new_P1_R1117_U281, new_P1_R1117_U282,
    new_P1_R1117_U283, new_P1_R1117_U284, new_P1_R1117_U285,
    new_P1_R1117_U286, new_P1_R1117_U287, new_P1_R1117_U288,
    new_P1_R1117_U289, new_P1_R1117_U290, new_P1_R1117_U291,
    new_P1_R1117_U292, new_P1_R1117_U293, new_P1_R1117_U294,
    new_P1_R1117_U295, new_P1_R1117_U296, new_P1_R1117_U297,
    new_P1_R1117_U298, new_P1_R1117_U299, new_P1_R1117_U300,
    new_P1_R1117_U301, new_P1_R1117_U302, new_P1_R1117_U303,
    new_P1_R1117_U304, new_P1_R1117_U305, new_P1_R1117_U306,
    new_P1_R1117_U307, new_P1_R1117_U308, new_P1_R1117_U309,
    new_P1_R1117_U310, new_P1_R1117_U311, new_P1_R1117_U312,
    new_P1_R1117_U313, new_P1_R1117_U314, new_P1_R1117_U315,
    new_P1_R1117_U316, new_P1_R1117_U317, new_P1_R1117_U318,
    new_P1_R1117_U319, new_P1_R1117_U320, new_P1_R1117_U321,
    new_P1_R1117_U322, new_P1_R1117_U323, new_P1_R1117_U324,
    new_P1_R1117_U325, new_P1_R1117_U326, new_P1_R1117_U327,
    new_P1_R1117_U328, new_P1_R1117_U329, new_P1_R1117_U330,
    new_P1_R1117_U331, new_P1_R1117_U332, new_P1_R1117_U333,
    new_P1_R1117_U334, new_P1_R1117_U335, new_P1_R1117_U336,
    new_P1_R1117_U337, new_P1_R1117_U338, new_P1_R1117_U339,
    new_P1_R1117_U340, new_P1_R1117_U341, new_P1_R1117_U342,
    new_P1_R1117_U343, new_P1_R1117_U344, new_P1_R1117_U345,
    new_P1_R1117_U346, new_P1_R1117_U347, new_P1_R1117_U348,
    new_P1_R1117_U349, new_P1_R1117_U350, new_P1_R1117_U351,
    new_P1_R1117_U352, new_P1_R1117_U353, new_P1_R1117_U354,
    new_P1_R1117_U355, new_P1_R1117_U356, new_P1_R1117_U357,
    new_P1_R1117_U358, new_P1_R1117_U359, new_P1_R1117_U360,
    new_P1_R1117_U361, new_P1_R1117_U362, new_P1_R1117_U363,
    new_P1_R1117_U364, new_P1_R1117_U365, new_P1_R1117_U366,
    new_P1_R1117_U367, new_P1_R1117_U368, new_P1_R1117_U369,
    new_P1_R1117_U370, new_P1_R1117_U371, new_P1_R1117_U372,
    new_P1_R1117_U373, new_P1_R1117_U374, new_P1_R1117_U375,
    new_P1_R1117_U376, new_P1_R1117_U377, new_P1_R1117_U378,
    new_P1_R1117_U379, new_P1_R1117_U380, new_P1_R1117_U381,
    new_P1_R1117_U382, new_P1_R1117_U383, new_P1_R1117_U384,
    new_P1_R1117_U385, new_P1_R1117_U386, new_P1_R1117_U387,
    new_P1_R1117_U388, new_P1_R1117_U389, new_P1_R1117_U390,
    new_P1_R1117_U391, new_P1_R1117_U392, new_P1_R1117_U393,
    new_P1_R1117_U394, new_P1_R1117_U395, new_P1_R1117_U396,
    new_P1_R1117_U397, new_P1_R1117_U398, new_P1_R1117_U399,
    new_P1_R1117_U400, new_P1_R1117_U401, new_P1_R1117_U402,
    new_P1_R1117_U403, new_P1_R1117_U404, new_P1_R1117_U405,
    new_P1_R1117_U406, new_P1_R1117_U407, new_P1_R1117_U408,
    new_P1_R1117_U409, new_P1_R1117_U410, new_P1_R1117_U411,
    new_P1_R1117_U412, new_P1_R1117_U413, new_P1_R1117_U414,
    new_P1_R1117_U415, new_P1_R1117_U416, new_P1_R1117_U417,
    new_P1_R1117_U418, new_P1_R1117_U419, new_P1_R1117_U420,
    new_P1_R1117_U421, new_P1_R1117_U422, new_P1_R1117_U423,
    new_P1_R1117_U424, new_P1_R1117_U425, new_P1_R1117_U426,
    new_P1_R1117_U427, new_P1_R1117_U428, new_P1_R1117_U429,
    new_P1_R1117_U430, new_P1_R1117_U431, new_P1_R1117_U432,
    new_P1_R1117_U433, new_P1_R1117_U434, new_P1_R1117_U435,
    new_P1_R1117_U436, new_P1_R1117_U437, new_P1_R1117_U438,
    new_P1_R1117_U439, new_P1_R1117_U440, new_P1_R1117_U441,
    new_P1_R1117_U442, new_P1_R1117_U443, new_P1_R1117_U444,
    new_P1_R1117_U445, new_P1_R1117_U446, new_P1_R1117_U447,
    new_P1_R1117_U448, new_P1_R1117_U449, new_P1_R1117_U450,
    new_P1_R1117_U451, new_P1_R1117_U452, new_P1_R1117_U453,
    new_P1_R1117_U454, new_P1_R1117_U455, new_P1_R1117_U456,
    new_P1_R1117_U457, new_P1_R1117_U458, new_P1_R1117_U459,
    new_P1_R1117_U460, new_P1_R1117_U461, new_P1_R1117_U462,
    new_P1_R1117_U463, new_P1_R1117_U464, new_P1_R1117_U465,
    new_P1_R1117_U466, new_P1_R1117_U467, new_P1_R1117_U468,
    new_P1_R1117_U469, new_P1_R1117_U470, new_P1_R1117_U471,
    new_P1_R1117_U472, new_P1_R1117_U473, new_P1_R1117_U474,
    new_P1_R1117_U475, new_P1_R1117_U476, new_P1_R1375_U6, new_P1_R1375_U7,
    new_P1_R1375_U8, new_P1_R1375_U9, new_P1_R1375_U10, new_P1_R1375_U11,
    new_P1_R1375_U12, new_P1_R1375_U13, new_P1_R1375_U14, new_P1_R1375_U15,
    new_P1_R1375_U16, new_P1_R1375_U17, new_P1_R1375_U18, new_P1_R1375_U19,
    new_P1_R1375_U20, new_P1_R1375_U21, new_P1_R1375_U22, new_P1_R1375_U23,
    new_P1_R1375_U24, new_P1_R1375_U25, new_P1_R1375_U26, new_P1_R1375_U27,
    new_P1_R1375_U28, new_P1_R1375_U29, new_P1_R1375_U30, new_P1_R1375_U31,
    new_P1_R1375_U32, new_P1_R1375_U33, new_P1_R1375_U34, new_P1_R1375_U35,
    new_P1_R1375_U36, new_P1_R1375_U37, new_P1_R1375_U38, new_P1_R1375_U39,
    new_P1_R1375_U40, new_P1_R1375_U41, new_P1_R1375_U42, new_P1_R1375_U43,
    new_P1_R1375_U44, new_P1_R1375_U45, new_P1_R1375_U46, new_P1_R1375_U47,
    new_P1_R1375_U48, new_P1_R1375_U49, new_P1_R1375_U50, new_P1_R1375_U51,
    new_P1_R1375_U52, new_P1_R1375_U53, new_P1_R1375_U54, new_P1_R1375_U55,
    new_P1_R1375_U56, new_P1_R1375_U57, new_P1_R1375_U58, new_P1_R1375_U59,
    new_P1_R1375_U60, new_P1_R1375_U61, new_P1_R1375_U62, new_P1_R1375_U63,
    new_P1_R1375_U64, new_P1_R1375_U65, new_P1_R1375_U66, new_P1_R1375_U67,
    new_P1_R1375_U68, new_P1_R1375_U69, new_P1_R1375_U70, new_P1_R1375_U71,
    new_P1_R1375_U72, new_P1_R1375_U73, new_P1_R1375_U74, new_P1_R1375_U75,
    new_P1_R1375_U76, new_P1_R1375_U77, new_P1_R1375_U78, new_P1_R1375_U79,
    new_P1_R1375_U80, new_P1_R1375_U81, new_P1_R1375_U82, new_P1_R1375_U83,
    new_P1_R1375_U84, new_P1_R1375_U85, new_P1_R1375_U86, new_P1_R1375_U87,
    new_P1_R1375_U88, new_P1_R1375_U89, new_P1_R1375_U90, new_P1_R1375_U91,
    new_P1_R1375_U92, new_P1_R1375_U93, new_P1_R1375_U94, new_P1_R1375_U95,
    new_P1_R1375_U96, new_P1_R1375_U97, new_P1_R1375_U98, new_P1_R1375_U99,
    new_P1_R1375_U100, new_P1_R1375_U101, new_P1_R1375_U102,
    new_P1_R1375_U103, new_P1_R1375_U104, new_P1_R1375_U105,
    new_P1_R1375_U106, new_P1_R1375_U107, new_P1_R1375_U108,
    new_P1_R1375_U109, new_P1_R1375_U110, new_P1_R1375_U111,
    new_P1_R1375_U112, new_P1_R1375_U113, new_P1_R1375_U114,
    new_P1_R1375_U115, new_P1_R1375_U116, new_P1_R1375_U117,
    new_P1_R1375_U118, new_P1_R1375_U119, new_P1_R1375_U120,
    new_P1_R1375_U121, new_P1_R1375_U122, new_P1_R1375_U123,
    new_P1_R1375_U124, new_P1_R1375_U125, new_P1_R1375_U126,
    new_P1_R1375_U127, new_P1_R1375_U128, new_P1_R1375_U129,
    new_P1_R1375_U130, new_P1_R1375_U131, new_P1_R1375_U132,
    new_P1_R1375_U133, new_P1_R1375_U134, new_P1_R1375_U135,
    new_P1_R1375_U136, new_P1_R1375_U137, new_P1_R1375_U138,
    new_P1_R1375_U139, new_P1_R1375_U140, new_P1_R1375_U141,
    new_P1_R1375_U142, new_P1_R1375_U143, new_P1_R1375_U144,
    new_P1_R1375_U145, new_P1_R1375_U146, new_P1_R1375_U147,
    new_P1_R1375_U148, new_P1_R1375_U149, new_P1_R1375_U150,
    new_P1_R1375_U151, new_P1_R1375_U152, new_P1_R1375_U153,
    new_P1_R1375_U154, new_P1_R1375_U155, new_P1_R1375_U156,
    new_P1_R1375_U157, new_P1_R1375_U158, new_P1_R1375_U159,
    new_P1_R1375_U160, new_P1_R1375_U161, new_P1_R1375_U162,
    new_P1_R1375_U163, new_P1_R1375_U164, new_P1_R1375_U165,
    new_P1_R1375_U166, new_P1_R1375_U167, new_P1_R1375_U168,
    new_P1_R1375_U169, new_P1_R1375_U170, new_P1_R1375_U171,
    new_P1_R1375_U172, new_P1_R1375_U173, new_P1_R1375_U174,
    new_P1_R1375_U175, new_P1_R1375_U176, new_P1_R1375_U177,
    new_P1_R1375_U178, new_P1_R1375_U179, new_P1_R1375_U180,
    new_P1_R1375_U181, new_P1_R1375_U182, new_P1_R1375_U183,
    new_P1_R1375_U184, new_P1_R1375_U185, new_P1_R1375_U186,
    new_P1_R1375_U187, new_P1_R1375_U188, new_P1_R1375_U189,
    new_P1_R1375_U190, new_P1_R1375_U191, new_P1_R1375_U192,
    new_P1_R1375_U193, new_P1_R1375_U194, new_P1_R1375_U195,
    new_P1_R1375_U196, new_P1_R1375_U197, new_P1_R1352_U6, new_P1_R1352_U7,
    new_P1_R1207_U6, new_P1_R1207_U7, new_P1_R1207_U8, new_P1_R1207_U9,
    new_P1_R1207_U10, new_P1_R1207_U11, new_P1_R1207_U12, new_P1_R1207_U13,
    new_P1_R1207_U14, new_P1_R1207_U15, new_P1_R1207_U16, new_P1_R1207_U17,
    new_P1_R1207_U18, new_P1_R1207_U19, new_P1_R1207_U20, new_P1_R1207_U21,
    new_P1_R1207_U22, new_P1_R1207_U23, new_P1_R1207_U24, new_P1_R1207_U25,
    new_P1_R1207_U26, new_P1_R1207_U27, new_P1_R1207_U28, new_P1_R1207_U29,
    new_P1_R1207_U30, new_P1_R1207_U31, new_P1_R1207_U32, new_P1_R1207_U33,
    new_P1_R1207_U34, new_P1_R1207_U35, new_P1_R1207_U36, new_P1_R1207_U37,
    new_P1_R1207_U38, new_P1_R1207_U39, new_P1_R1207_U40, new_P1_R1207_U41,
    new_P1_R1207_U42, new_P1_R1207_U43, new_P1_R1207_U44, new_P1_R1207_U45,
    new_P1_R1207_U46, new_P1_R1207_U47, new_P1_R1207_U48, new_P1_R1207_U49,
    new_P1_R1207_U50, new_P1_R1207_U51, new_P1_R1207_U52, new_P1_R1207_U53,
    new_P1_R1207_U54, new_P1_R1207_U55, new_P1_R1207_U56, new_P1_R1207_U57,
    new_P1_R1207_U58, new_P1_R1207_U59, new_P1_R1207_U60, new_P1_R1207_U61,
    new_P1_R1207_U62, new_P1_R1207_U63, new_P1_R1207_U64, new_P1_R1207_U65,
    new_P1_R1207_U66, new_P1_R1207_U67, new_P1_R1207_U68, new_P1_R1207_U69,
    new_P1_R1207_U70, new_P1_R1207_U71, new_P1_R1207_U72, new_P1_R1207_U73,
    new_P1_R1207_U74, new_P1_R1207_U75, new_P1_R1207_U76, new_P1_R1207_U77,
    new_P1_R1207_U78, new_P1_R1207_U79, new_P1_R1207_U80, new_P1_R1207_U81,
    new_P1_R1207_U82, new_P1_R1207_U83, new_P1_R1207_U84, new_P1_R1207_U85,
    new_P1_R1207_U86, new_P1_R1207_U87, new_P1_R1207_U88, new_P1_R1207_U89,
    new_P1_R1207_U90, new_P1_R1207_U91, new_P1_R1207_U92, new_P1_R1207_U93,
    new_P1_R1207_U94, new_P1_R1207_U95, new_P1_R1207_U96, new_P1_R1207_U97,
    new_P1_R1207_U98, new_P1_R1207_U99, new_P1_R1207_U100,
    new_P1_R1207_U101, new_P1_R1207_U102, new_P1_R1207_U103,
    new_P1_R1207_U104, new_P1_R1207_U105, new_P1_R1207_U106,
    new_P1_R1207_U107, new_P1_R1207_U108, new_P1_R1207_U109,
    new_P1_R1207_U110, new_P1_R1207_U111, new_P1_R1207_U112,
    new_P1_R1207_U113, new_P1_R1207_U114, new_P1_R1207_U115,
    new_P1_R1207_U116, new_P1_R1207_U117, new_P1_R1207_U118,
    new_P1_R1207_U119, new_P1_R1207_U120, new_P1_R1207_U121,
    new_P1_R1207_U122, new_P1_R1207_U123, new_P1_R1207_U124,
    new_P1_R1207_U125, new_P1_R1207_U126, new_P1_R1207_U127,
    new_P1_R1207_U128, new_P1_R1207_U129, new_P1_R1207_U130,
    new_P1_R1207_U131, new_P1_R1207_U132, new_P1_R1207_U133,
    new_P1_R1207_U134, new_P1_R1207_U135, new_P1_R1207_U136,
    new_P1_R1207_U137, new_P1_R1207_U138, new_P1_R1207_U139,
    new_P1_R1207_U140, new_P1_R1207_U141, new_P1_R1207_U142,
    new_P1_R1207_U143, new_P1_R1207_U144, new_P1_R1207_U145,
    new_P1_R1207_U146, new_P1_R1207_U147, new_P1_R1207_U148,
    new_P1_R1207_U149, new_P1_R1207_U150, new_P1_R1207_U151,
    new_P1_R1207_U152, new_P1_R1207_U153, new_P1_R1207_U154,
    new_P1_R1207_U155, new_P1_R1207_U156, new_P1_R1207_U157,
    new_P1_R1207_U158, new_P1_R1207_U159, new_P1_R1207_U160,
    new_P1_R1207_U161, new_P1_R1207_U162, new_P1_R1207_U163,
    new_P1_R1207_U164, new_P1_R1207_U165, new_P1_R1207_U166,
    new_P1_R1207_U167, new_P1_R1207_U168, new_P1_R1207_U169,
    new_P1_R1207_U170, new_P1_R1207_U171, new_P1_R1207_U172,
    new_P1_R1207_U173, new_P1_R1207_U174, new_P1_R1207_U175,
    new_P1_R1207_U176, new_P1_R1207_U177, new_P1_R1207_U178,
    new_P1_R1207_U179, new_P1_R1207_U180, new_P1_R1207_U181,
    new_P1_R1207_U182, new_P1_R1207_U183, new_P1_R1207_U184,
    new_P1_R1207_U185, new_P1_R1207_U186, new_P1_R1207_U187,
    new_P1_R1207_U188, new_P1_R1207_U189, new_P1_R1207_U190,
    new_P1_R1207_U191, new_P1_R1207_U192, new_P1_R1207_U193,
    new_P1_R1207_U194, new_P1_R1207_U195, new_P1_R1207_U196,
    new_P1_R1207_U197, new_P1_R1207_U198, new_P1_R1207_U199,
    new_P1_R1207_U200, new_P1_R1207_U201, new_P1_R1207_U202,
    new_P1_R1207_U203, new_P1_R1207_U204, new_P1_R1207_U205,
    new_P1_R1207_U206, new_P1_R1207_U207, new_P1_R1207_U208,
    new_P1_R1207_U209, new_P1_R1207_U210, new_P1_R1207_U211,
    new_P1_R1207_U212, new_P1_R1207_U213, new_P1_R1207_U214,
    new_P1_R1207_U215, new_P1_R1207_U216, new_P1_R1207_U217,
    new_P1_R1207_U218, new_P1_R1207_U219, new_P1_R1207_U220,
    new_P1_R1207_U221, new_P1_R1207_U222, new_P1_R1207_U223,
    new_P1_R1207_U224, new_P1_R1207_U225, new_P1_R1207_U226,
    new_P1_R1207_U227, new_P1_R1207_U228, new_P1_R1207_U229,
    new_P1_R1207_U230, new_P1_R1207_U231, new_P1_R1207_U232,
    new_P1_R1207_U233, new_P1_R1207_U234, new_P1_R1207_U235,
    new_P1_R1207_U236, new_P1_R1207_U237, new_P1_R1207_U238,
    new_P1_R1207_U239, new_P1_R1207_U240, new_P1_R1207_U241,
    new_P1_R1207_U242, new_P1_R1207_U243, new_P1_R1207_U244,
    new_P1_R1207_U245, new_P1_R1207_U246, new_P1_R1207_U247,
    new_P1_R1207_U248, new_P1_R1207_U249, new_P1_R1207_U250,
    new_P1_R1207_U251, new_P1_R1207_U252, new_P1_R1207_U253,
    new_P1_R1207_U254, new_P1_R1207_U255, new_P1_R1207_U256,
    new_P1_R1207_U257, new_P1_R1207_U258, new_P1_R1207_U259,
    new_P1_R1207_U260, new_P1_R1207_U261, new_P1_R1207_U262,
    new_P1_R1207_U263, new_P1_R1207_U264, new_P1_R1207_U265,
    new_P1_R1207_U266, new_P1_R1207_U267, new_P1_R1207_U268,
    new_P1_R1207_U269, new_P1_R1207_U270, new_P1_R1207_U271,
    new_P1_R1207_U272, new_P1_R1207_U273, new_P1_R1207_U274,
    new_P1_R1207_U275, new_P1_R1207_U276, new_P1_R1207_U277,
    new_P1_R1207_U278, new_P1_R1207_U279, new_P1_R1207_U280,
    new_P1_R1207_U281, new_P1_R1207_U282, new_P1_R1207_U283,
    new_P1_R1207_U284, new_P1_R1207_U285, new_P1_R1207_U286,
    new_P1_R1207_U287, new_P1_R1207_U288, new_P1_R1207_U289,
    new_P1_R1207_U290, new_P1_R1207_U291, new_P1_R1207_U292,
    new_P1_R1207_U293, new_P1_R1207_U294, new_P1_R1207_U295,
    new_P1_R1207_U296, new_P1_R1207_U297, new_P1_R1207_U298,
    new_P1_R1207_U299, new_P1_R1207_U300, new_P1_R1207_U301,
    new_P1_R1207_U302, new_P1_R1207_U303, new_P1_R1207_U304,
    new_P1_R1207_U305, new_P1_R1207_U306, new_P1_R1207_U307,
    new_P1_R1207_U308, new_P1_R1207_U309, new_P1_R1207_U310,
    new_P1_R1207_U311, new_P1_R1207_U312, new_P1_R1207_U313,
    new_P1_R1207_U314, new_P1_R1207_U315, new_P1_R1207_U316,
    new_P1_R1207_U317, new_P1_R1207_U318, new_P1_R1207_U319,
    new_P1_R1207_U320, new_P1_R1207_U321, new_P1_R1207_U322,
    new_P1_R1207_U323, new_P1_R1207_U324, new_P1_R1207_U325,
    new_P1_R1207_U326, new_P1_R1207_U327, new_P1_R1207_U328,
    new_P1_R1207_U329, new_P1_R1207_U330, new_P1_R1207_U331,
    new_P1_R1207_U332, new_P1_R1207_U333, new_P1_R1207_U334,
    new_P1_R1207_U335, new_P1_R1207_U336, new_P1_R1207_U337,
    new_P1_R1207_U338, new_P1_R1207_U339, new_P1_R1207_U340,
    new_P1_R1207_U341, new_P1_R1207_U342, new_P1_R1207_U343,
    new_P1_R1207_U344, new_P1_R1207_U345, new_P1_R1207_U346,
    new_P1_R1207_U347, new_P1_R1207_U348, new_P1_R1207_U349,
    new_P1_R1207_U350, new_P1_R1207_U351, new_P1_R1207_U352,
    new_P1_R1207_U353, new_P1_R1207_U354, new_P1_R1207_U355,
    new_P1_R1207_U356, new_P1_R1207_U357, new_P1_R1207_U358,
    new_P1_R1207_U359, new_P1_R1207_U360, new_P1_R1207_U361,
    new_P1_R1207_U362, new_P1_R1207_U363, new_P1_R1207_U364,
    new_P1_R1207_U365, new_P1_R1207_U366, new_P1_R1207_U367,
    new_P1_R1207_U368, new_P1_R1207_U369, new_P1_R1207_U370,
    new_P1_R1207_U371, new_P1_R1207_U372, new_P1_R1207_U373,
    new_P1_R1207_U374, new_P1_R1207_U375, new_P1_R1207_U376,
    new_P1_R1207_U377, new_P1_R1207_U378, new_P1_R1207_U379,
    new_P1_R1207_U380, new_P1_R1207_U381, new_P1_R1207_U382,
    new_P1_R1207_U383, new_P1_R1207_U384, new_P1_R1207_U385,
    new_P1_R1207_U386, new_P1_R1207_U387, new_P1_R1207_U388,
    new_P1_R1207_U389, new_P1_R1207_U390, new_P1_R1207_U391,
    new_P1_R1207_U392, new_P1_R1207_U393, new_P1_R1207_U394,
    new_P1_R1207_U395, new_P1_R1207_U396, new_P1_R1207_U397,
    new_P1_R1207_U398, new_P1_R1207_U399, new_P1_R1207_U400,
    new_P1_R1207_U401, new_P1_R1207_U402, new_P1_R1207_U403,
    new_P1_R1207_U404, new_P1_R1207_U405, new_P1_R1207_U406,
    new_P1_R1207_U407, new_P1_R1207_U408, new_P1_R1207_U409,
    new_P1_R1207_U410, new_P1_R1207_U411, new_P1_R1207_U412,
    new_P1_R1207_U413, new_P1_R1207_U414, new_P1_R1207_U415,
    new_P1_R1207_U416, new_P1_R1207_U417, new_P1_R1207_U418,
    new_P1_R1207_U419, new_P1_R1207_U420, new_P1_R1207_U421,
    new_P1_R1207_U422, new_P1_R1207_U423, new_P1_R1207_U424,
    new_P1_R1207_U425, new_P1_R1207_U426, new_P1_R1207_U427,
    new_P1_R1207_U428, new_P1_R1207_U429, new_P1_R1207_U430,
    new_P1_R1207_U431, new_P1_R1207_U432, new_P1_R1207_U433,
    new_P1_R1207_U434, new_P1_R1207_U435, new_P1_R1207_U436,
    new_P1_R1207_U437, new_P1_R1207_U438, new_P1_R1207_U439,
    new_P1_R1207_U440, new_P1_R1207_U441, new_P1_R1207_U442,
    new_P1_R1207_U443, new_P1_R1207_U444, new_P1_R1207_U445,
    new_P1_R1207_U446, new_P1_R1207_U447, new_P1_R1207_U448,
    new_P1_R1207_U449, new_P1_R1207_U450, new_P1_R1207_U451,
    new_P1_R1207_U452, new_P1_R1207_U453, new_P1_R1207_U454,
    new_P1_R1207_U455, new_P1_R1207_U456, new_P1_R1207_U457,
    new_P1_R1207_U458, new_P1_R1207_U459, new_P1_R1207_U460,
    new_P1_R1207_U461, new_P1_R1207_U462, new_P1_R1207_U463,
    new_P1_R1207_U464, new_P1_R1207_U465, new_P1_R1207_U466,
    new_P1_R1207_U467, new_P1_R1207_U468, new_P1_R1207_U469,
    new_P1_R1207_U470, new_P1_R1207_U471, new_P1_R1207_U472,
    new_P1_R1207_U473, new_P1_R1207_U474, new_P1_R1207_U475,
    new_P1_R1207_U476, new_P1_R1165_U4, new_P1_R1165_U5, new_P1_R1165_U6,
    new_P1_R1165_U7, new_P1_R1165_U8, new_P1_R1165_U9, new_P1_R1165_U10,
    new_P1_R1165_U11, new_P1_R1165_U12, new_P1_R1165_U13, new_P1_R1165_U14,
    new_P1_R1165_U15, new_P1_R1165_U16, new_P1_R1165_U17, new_P1_R1165_U18,
    new_P1_R1165_U19, new_P1_R1165_U20, new_P1_R1165_U21, new_P1_R1165_U22,
    new_P1_R1165_U23, new_P1_R1165_U24, new_P1_R1165_U25, new_P1_R1165_U26,
    new_P1_R1165_U27, new_P1_R1165_U28, new_P1_R1165_U29, new_P1_R1165_U30,
    new_P1_R1165_U31, new_P1_R1165_U32, new_P1_R1165_U33, new_P1_R1165_U34,
    new_P1_R1165_U35, new_P1_R1165_U36, new_P1_R1165_U37, new_P1_R1165_U38,
    new_P1_R1165_U39, new_P1_R1165_U40, new_P1_R1165_U41, new_P1_R1165_U42,
    new_P1_R1165_U43, new_P1_R1165_U44, new_P1_R1165_U45, new_P1_R1165_U46,
    new_P1_R1165_U47, new_P1_R1165_U48, new_P1_R1165_U49, new_P1_R1165_U50,
    new_P1_R1165_U51, new_P1_R1165_U52, new_P1_R1165_U53, new_P1_R1165_U54,
    new_P1_R1165_U55, new_P1_R1165_U56, new_P1_R1165_U57, new_P1_R1165_U58,
    new_P1_R1165_U59, new_P1_R1165_U60, new_P1_R1165_U61, new_P1_R1165_U62,
    new_P1_R1165_U63, new_P1_R1165_U64, new_P1_R1165_U65, new_P1_R1165_U66,
    new_P1_R1165_U67, new_P1_R1165_U68, new_P1_R1165_U69, new_P1_R1165_U70,
    new_P1_R1165_U71, new_P1_R1165_U72, new_P1_R1165_U73, new_P1_R1165_U74,
    new_P1_R1165_U75, new_P1_R1165_U76, new_P1_R1165_U77, new_P1_R1165_U78,
    new_P1_R1165_U79, new_P1_R1165_U80, new_P1_R1165_U81, new_P1_R1165_U82,
    new_P1_R1165_U83, new_P1_R1165_U84, new_P1_R1165_U85, new_P1_R1165_U86,
    new_P1_R1165_U87, new_P1_R1165_U88, new_P1_R1165_U89, new_P1_R1165_U90,
    new_P1_R1165_U91, new_P1_R1165_U92, new_P1_R1165_U93, new_P1_R1165_U94,
    new_P1_R1165_U95, new_P1_R1165_U96, new_P1_R1165_U97, new_P1_R1165_U98,
    new_P1_R1165_U99, new_P1_R1165_U100, new_P1_R1165_U101,
    new_P1_R1165_U102, new_P1_R1165_U103, new_P1_R1165_U104,
    new_P1_R1165_U105, new_P1_R1165_U106, new_P1_R1165_U107,
    new_P1_R1165_U108, new_P1_R1165_U109, new_P1_R1165_U110,
    new_P1_R1165_U111, new_P1_R1165_U112, new_P1_R1165_U113,
    new_P1_R1165_U114, new_P1_R1165_U115, new_P1_R1165_U116,
    new_P1_R1165_U117, new_P1_R1165_U118, new_P1_R1165_U119,
    new_P1_R1165_U120, new_P1_R1165_U121, new_P1_R1165_U122,
    new_P1_R1165_U123, new_P1_R1165_U124, new_P1_R1165_U125,
    new_P1_R1165_U126, new_P1_R1165_U127, new_P1_R1165_U128,
    new_P1_R1165_U129, new_P1_R1165_U130, new_P1_R1165_U131,
    new_P1_R1165_U132, new_P1_R1165_U133, new_P1_R1165_U134,
    new_P1_R1165_U135, new_P1_R1165_U136, new_P1_R1165_U137,
    new_P1_R1165_U138, new_P1_R1165_U139, new_P1_R1165_U140,
    new_P1_R1165_U141, new_P1_R1165_U142, new_P1_R1165_U143,
    new_P1_R1165_U144, new_P1_R1165_U145, new_P1_R1165_U146,
    new_P1_R1165_U147, new_P1_R1165_U148, new_P1_R1165_U149,
    new_P1_R1165_U150, new_P1_R1165_U151, new_P1_R1165_U152,
    new_P1_R1165_U153, new_P1_R1165_U154, new_P1_R1165_U155,
    new_P1_R1165_U156, new_P1_R1165_U157, new_P1_R1165_U158,
    new_P1_R1165_U159, new_P1_R1165_U160, new_P1_R1165_U161,
    new_P1_R1165_U162, new_P1_R1165_U163, new_P1_R1165_U164,
    new_P1_R1165_U165, new_P1_R1165_U166, new_P1_R1165_U167,
    new_P1_R1165_U168, new_P1_R1165_U169, new_P1_R1165_U170,
    new_P1_R1165_U171, new_P1_R1165_U172, new_P1_R1165_U173,
    new_P1_R1165_U174, new_P1_R1165_U175, new_P1_R1165_U176,
    new_P1_R1165_U177, new_P1_R1165_U178, new_P1_R1165_U179,
    new_P1_R1165_U180, new_P1_R1165_U181, new_P1_R1165_U182,
    new_P1_R1165_U183, new_P1_R1165_U184, new_P1_R1165_U185,
    new_P1_R1165_U186, new_P1_R1165_U187, new_P1_R1165_U188,
    new_P1_R1165_U189, new_P1_R1165_U190, new_P1_R1165_U191,
    new_P1_R1165_U192, new_P1_R1165_U193, new_P1_R1165_U194,
    new_P1_R1165_U195, new_P1_R1165_U196, new_P1_R1165_U197,
    new_P1_R1165_U198, new_P1_R1165_U199, new_P1_R1165_U200,
    new_P1_R1165_U201, new_P1_R1165_U202, new_P1_R1165_U203,
    new_P1_R1165_U204, new_P1_R1165_U205, new_P1_R1165_U206,
    new_P1_R1165_U207, new_P1_R1165_U208, new_P1_R1165_U209,
    new_P1_R1165_U210, new_P1_R1165_U211, new_P1_R1165_U212,
    new_P1_R1165_U213, new_P1_R1165_U214, new_P1_R1165_U215,
    new_P1_R1165_U216, new_P1_R1165_U217, new_P1_R1165_U218,
    new_P1_R1165_U219, new_P1_R1165_U220, new_P1_R1165_U221,
    new_P1_R1165_U222, new_P1_R1165_U223, new_P1_R1165_U224,
    new_P1_R1165_U225, new_P1_R1165_U226, new_P1_R1165_U227,
    new_P1_R1165_U228, new_P1_R1165_U229, new_P1_R1165_U230,
    new_P1_R1165_U231, new_P1_R1165_U232, new_P1_R1165_U233,
    new_P1_R1165_U234, new_P1_R1165_U235, new_P1_R1165_U236,
    new_P1_R1165_U237, new_P1_R1165_U238, new_P1_R1165_U239,
    new_P1_R1165_U240, new_P1_R1165_U241, new_P1_R1165_U242,
    new_P1_R1165_U243, new_P1_R1165_U244, new_P1_R1165_U245,
    new_P1_R1165_U246, new_P1_R1165_U247, new_P1_R1165_U248,
    new_P1_R1165_U249, new_P1_R1165_U250, new_P1_R1165_U251,
    new_P1_R1165_U252, new_P1_R1165_U253, new_P1_R1165_U254,
    new_P1_R1165_U255, new_P1_R1165_U256, new_P1_R1165_U257,
    new_P1_R1165_U258, new_P1_R1165_U259, new_P1_R1165_U260,
    new_P1_R1165_U261, new_P1_R1165_U262, new_P1_R1165_U263,
    new_P1_R1165_U264, new_P1_R1165_U265, new_P1_R1165_U266,
    new_P1_R1165_U267, new_P1_R1165_U268, new_P1_R1165_U269,
    new_P1_R1165_U270, new_P1_R1165_U271, new_P1_R1165_U272,
    new_P1_R1165_U273, new_P1_R1165_U274, new_P1_R1165_U275,
    new_P1_R1165_U276, new_P1_R1165_U277, new_P1_R1165_U278,
    new_P1_R1165_U279, new_P1_R1165_U280, new_P1_R1165_U281,
    new_P1_R1165_U282, new_P1_R1165_U283, new_P1_R1165_U284,
    new_P1_R1165_U285, new_P1_R1165_U286, new_P1_R1165_U287,
    new_P1_R1165_U288, new_P1_R1165_U289, new_P1_R1165_U290,
    new_P1_R1165_U291, new_P1_R1165_U292, new_P1_R1165_U293,
    new_P1_R1165_U294, new_P1_R1165_U295, new_P1_R1165_U296,
    new_P1_R1165_U297, new_P1_R1165_U298, new_P1_R1165_U299,
    new_P1_R1165_U300, new_P1_R1165_U301, new_P1_R1165_U302,
    new_P1_R1165_U303, new_P1_R1165_U304, new_P1_R1165_U305,
    new_P1_R1165_U306, new_P1_R1165_U307, new_P1_R1165_U308,
    new_P1_R1165_U309, new_P1_R1165_U310, new_P1_R1165_U311,
    new_P1_R1165_U312, new_P1_R1165_U313, new_P1_R1165_U314,
    new_P1_R1165_U315, new_P1_R1165_U316, new_P1_R1165_U317,
    new_P1_R1165_U318, new_P1_R1165_U319, new_P1_R1165_U320,
    new_P1_R1165_U321, new_P1_R1165_U322, new_P1_R1165_U323,
    new_P1_R1165_U324, new_P1_R1165_U325, new_P1_R1165_U326,
    new_P1_R1165_U327, new_P1_R1165_U328, new_P1_R1165_U329,
    new_P1_R1165_U330, new_P1_R1165_U331, new_P1_R1165_U332,
    new_P1_R1165_U333, new_P1_R1165_U334, new_P1_R1165_U335,
    new_P1_R1165_U336, new_P1_R1165_U337, new_P1_R1165_U338,
    new_P1_R1165_U339, new_P1_R1165_U340, new_P1_R1165_U341,
    new_P1_R1165_U342, new_P1_R1165_U343, new_P1_R1165_U344,
    new_P1_R1165_U345, new_P1_R1165_U346, new_P1_R1165_U347,
    new_P1_R1165_U348, new_P1_R1165_U349, new_P1_R1165_U350,
    new_P1_R1165_U351, new_P1_R1165_U352, new_P1_R1165_U353,
    new_P1_R1165_U354, new_P1_R1165_U355, new_P1_R1165_U356,
    new_P1_R1165_U357, new_P1_R1165_U358, new_P1_R1165_U359,
    new_P1_R1165_U360, new_P1_R1165_U361, new_P1_R1165_U362,
    new_P1_R1165_U363, new_P1_R1165_U364, new_P1_R1165_U365,
    new_P1_R1165_U366, new_P1_R1165_U367, new_P1_R1165_U368,
    new_P1_R1165_U369, new_P1_R1165_U370, new_P1_R1165_U371,
    new_P1_R1165_U372, new_P1_R1165_U373, new_P1_R1165_U374,
    new_P1_R1165_U375, new_P1_R1165_U376, new_P1_R1165_U377,
    new_P1_R1165_U378, new_P1_R1165_U379, new_P1_R1165_U380,
    new_P1_R1165_U381, new_P1_R1165_U382, new_P1_R1165_U383,
    new_P1_R1165_U384, new_P1_R1165_U385, new_P1_R1165_U386,
    new_P1_R1165_U387, new_P1_R1165_U388, new_P1_R1165_U389,
    new_P1_R1165_U390, new_P1_R1165_U391, new_P1_R1165_U392,
    new_P1_R1165_U393, new_P1_R1165_U394, new_P1_R1165_U395,
    new_P1_R1165_U396, new_P1_R1165_U397, new_P1_R1165_U398,
    new_P1_R1165_U399, new_P1_R1165_U400, new_P1_R1165_U401,
    new_P1_R1165_U402, new_P1_R1165_U403, new_P1_R1165_U404,
    new_P1_R1165_U405, new_P1_R1165_U406, new_P1_R1165_U407,
    new_P1_R1165_U408, new_P1_R1165_U409, new_P1_R1165_U410,
    new_P1_R1165_U411, new_P1_R1165_U412, new_P1_R1165_U413,
    new_P1_R1165_U414, new_P1_R1165_U415, new_P1_R1165_U416,
    new_P1_R1165_U417, new_P1_R1165_U418, new_P1_R1165_U419,
    new_P1_R1165_U420, new_P1_R1165_U421, new_P1_R1165_U422,
    new_P1_R1165_U423, new_P1_R1165_U424, new_P1_R1165_U425,
    new_P1_R1165_U426, new_P1_R1165_U427, new_P1_R1165_U428,
    new_P1_R1165_U429, new_P1_R1165_U430, new_P1_R1165_U431,
    new_P1_R1165_U432, new_P1_R1165_U433, new_P1_R1165_U434,
    new_P1_R1165_U435, new_P1_R1165_U436, new_P1_R1165_U437,
    new_P1_R1165_U438, new_P1_R1165_U439, new_P1_R1165_U440,
    new_P1_R1165_U441, new_P1_R1165_U442, new_P1_R1165_U443,
    new_P1_R1165_U444, new_P1_R1165_U445, new_P1_R1165_U446,
    new_P1_R1165_U447, new_P1_R1165_U448, new_P1_R1165_U449,
    new_P1_R1165_U450, new_P1_R1165_U451, new_P1_R1165_U452,
    new_P1_R1165_U453, new_P1_R1165_U454, new_P1_R1165_U455,
    new_P1_R1165_U456, new_P1_R1165_U457, new_P1_R1165_U458,
    new_P1_R1165_U459, new_P1_R1165_U460, new_P1_R1165_U461,
    new_P1_R1165_U462, new_P1_R1165_U463, new_P1_R1165_U464,
    new_P1_R1165_U465, new_P1_R1165_U466, new_P1_R1165_U467,
    new_P1_R1165_U468, new_P1_R1165_U469, new_P1_R1165_U470,
    new_P1_R1165_U471, new_P1_R1165_U472, new_P1_R1165_U473,
    new_P1_R1165_U474, new_P1_R1165_U475, new_P1_R1165_U476,
    new_P1_R1165_U477, new_P1_R1165_U478, new_P1_R1165_U479,
    new_P1_R1165_U480, new_P1_R1165_U481, new_P1_R1165_U482,
    new_P1_R1165_U483, new_P1_R1165_U484, new_P1_R1165_U485,
    new_P1_R1165_U486, new_P1_R1165_U487, new_P1_R1165_U488,
    new_P1_R1165_U489, new_P1_R1165_U490, new_P1_R1165_U491,
    new_P1_R1165_U492, new_P1_R1165_U493, new_P1_R1165_U494,
    new_P1_R1165_U495, new_P1_R1165_U496, new_P1_R1165_U497,
    new_P1_R1165_U498, new_P1_R1165_U499, new_P1_R1165_U500,
    new_P1_R1165_U501, new_P1_R1165_U502, new_P1_R1165_U503,
    new_P1_R1165_U504, new_P1_R1165_U505, new_P1_R1165_U506,
    new_P1_R1165_U507, new_P1_R1165_U508, new_P1_R1165_U509,
    new_P1_R1165_U510, new_P1_R1165_U511, new_P1_R1165_U512,
    new_P1_R1165_U513, new_P1_R1165_U514, new_P1_R1165_U515,
    new_P1_R1165_U516, new_P1_R1165_U517, new_P1_R1165_U518,
    new_P1_R1165_U519, new_P1_R1165_U520, new_P1_R1165_U521,
    new_P1_R1165_U522, new_P1_R1165_U523, new_P1_R1165_U524,
    new_P1_R1165_U525, new_P1_R1165_U526, new_P1_R1165_U527,
    new_P1_R1165_U528, new_P1_R1165_U529, new_P1_R1165_U530,
    new_P1_R1165_U531, new_P1_R1165_U532, new_P1_R1165_U533,
    new_P1_R1165_U534, new_P1_R1165_U535, new_P1_R1165_U536,
    new_P1_R1165_U537, new_P1_R1165_U538, new_P1_R1165_U539,
    new_P1_R1165_U540, new_P1_R1165_U541, new_P1_R1165_U542,
    new_P1_R1165_U543, new_P1_R1165_U544, new_P1_R1165_U545,
    new_P1_R1165_U546, new_P1_R1165_U547, new_P1_R1165_U548,
    new_P1_R1165_U549, new_P1_R1165_U550, new_P1_R1165_U551,
    new_P1_R1165_U552, new_P1_R1165_U553, new_P1_R1165_U554,
    new_P1_R1165_U555, new_P1_R1165_U556, new_P1_R1165_U557,
    new_P1_R1165_U558, new_P1_R1165_U559, new_P1_R1165_U560,
    new_P1_R1165_U561, new_P1_R1165_U562, new_P1_R1165_U563,
    new_P1_R1165_U564, new_P1_R1165_U565, new_P1_R1165_U566,
    new_P1_R1165_U567, new_P1_R1165_U568, new_P1_R1165_U569,
    new_P1_R1165_U570, new_P1_R1165_U571, new_P1_R1165_U572,
    new_P1_R1165_U573, new_P1_R1165_U574, new_P1_R1165_U575,
    new_P1_R1165_U576, new_P1_R1165_U577, new_P1_R1165_U578,
    new_P1_R1165_U579, new_P1_R1165_U580, new_P1_R1165_U581,
    new_P1_R1165_U582, new_P1_R1165_U583, new_P1_R1165_U584,
    new_P1_R1165_U585, new_P1_R1165_U586, new_P1_R1165_U587,
    new_P1_R1165_U588, new_P1_R1165_U589, new_P1_R1165_U590,
    new_P1_R1165_U591, new_P1_R1165_U592, new_P1_R1165_U593,
    new_P1_R1165_U594, new_P1_R1165_U595, new_P1_R1150_U6, new_P1_R1150_U7,
    new_P1_R1150_U8, new_P1_R1150_U9, new_P1_R1150_U10, new_P1_R1150_U11,
    new_P1_R1150_U12, new_P1_R1150_U13, new_P1_R1150_U14, new_P1_R1150_U15,
    new_P1_R1150_U16, new_P1_R1150_U17, new_P1_R1150_U18, new_P1_R1150_U19,
    new_P1_R1150_U20, new_P1_R1150_U21, new_P1_R1150_U22, new_P1_R1150_U23,
    new_P1_R1150_U24, new_P1_R1150_U25, new_P1_R1150_U26, new_P1_R1150_U27,
    new_P1_R1150_U28, new_P1_R1150_U29, new_P1_R1150_U30, new_P1_R1150_U31,
    new_P1_R1150_U32, new_P1_R1150_U33, new_P1_R1150_U34, new_P1_R1150_U35,
    new_P1_R1150_U36, new_P1_R1150_U37, new_P1_R1150_U38, new_P1_R1150_U39,
    new_P1_R1150_U40, new_P1_R1150_U41, new_P1_R1150_U42, new_P1_R1150_U43,
    new_P1_R1150_U44, new_P1_R1150_U45, new_P1_R1150_U46, new_P1_R1150_U47,
    new_P1_R1150_U48, new_P1_R1150_U49, new_P1_R1150_U50, new_P1_R1150_U51,
    new_P1_R1150_U52, new_P1_R1150_U53, new_P1_R1150_U54, new_P1_R1150_U55,
    new_P1_R1150_U56, new_P1_R1150_U57, new_P1_R1150_U58, new_P1_R1150_U59,
    new_P1_R1150_U60, new_P1_R1150_U61, new_P1_R1150_U62, new_P1_R1150_U63,
    new_P1_R1150_U64, new_P1_R1150_U65, new_P1_R1150_U66, new_P1_R1150_U67,
    new_P1_R1150_U68, new_P1_R1150_U69, new_P1_R1150_U70, new_P1_R1150_U71,
    new_P1_R1150_U72, new_P1_R1150_U73, new_P1_R1150_U74, new_P1_R1150_U75,
    new_P1_R1150_U76, new_P1_R1150_U77, new_P1_R1150_U78, new_P1_R1150_U79,
    new_P1_R1150_U80, new_P1_R1150_U81, new_P1_R1150_U82, new_P1_R1150_U83,
    new_P1_R1150_U84, new_P1_R1150_U85, new_P1_R1150_U86, new_P1_R1150_U87,
    new_P1_R1150_U88, new_P1_R1150_U89, new_P1_R1150_U90, new_P1_R1150_U91,
    new_P1_R1150_U92, new_P1_R1150_U93, new_P1_R1150_U94, new_P1_R1150_U95,
    new_P1_R1150_U96, new_P1_R1150_U97, new_P1_R1150_U98, new_P1_R1150_U99,
    new_P1_R1150_U100, new_P1_R1150_U101, new_P1_R1150_U102,
    new_P1_R1150_U103, new_P1_R1150_U104, new_P1_R1150_U105,
    new_P1_R1150_U106, new_P1_R1150_U107, new_P1_R1150_U108,
    new_P1_R1150_U109, new_P1_R1150_U110, new_P1_R1150_U111,
    new_P1_R1150_U112, new_P1_R1150_U113, new_P1_R1150_U114,
    new_P1_R1150_U115, new_P1_R1150_U116, new_P1_R1150_U117,
    new_P1_R1150_U118, new_P1_R1150_U119, new_P1_R1150_U120,
    new_P1_R1150_U121, new_P1_R1150_U122, new_P1_R1150_U123,
    new_P1_R1150_U124, new_P1_R1150_U125, new_P1_R1150_U126,
    new_P1_R1150_U127, new_P1_R1150_U128, new_P1_R1150_U129,
    new_P1_R1150_U130, new_P1_R1150_U131, new_P1_R1150_U132,
    new_P1_R1150_U133, new_P1_R1150_U134, new_P1_R1150_U135,
    new_P1_R1150_U136, new_P1_R1150_U137, new_P1_R1150_U138,
    new_P1_R1150_U139, new_P1_R1150_U140, new_P1_R1150_U141,
    new_P1_R1150_U142, new_P1_R1150_U143, new_P1_R1150_U144,
    new_P1_R1150_U145, new_P1_R1150_U146, new_P1_R1150_U147,
    new_P1_R1150_U148, new_P1_R1150_U149, new_P1_R1150_U150,
    new_P1_R1150_U151, new_P1_R1150_U152, new_P1_R1150_U153,
    new_P1_R1150_U154, new_P1_R1150_U155, new_P1_R1150_U156,
    new_P1_R1150_U157, new_P1_R1150_U158, new_P1_R1150_U159,
    new_P1_R1150_U160, new_P1_R1150_U161, new_P1_R1150_U162,
    new_P1_R1150_U163, new_P1_R1150_U164, new_P1_R1150_U165,
    new_P1_R1150_U166, new_P1_R1150_U167, new_P1_R1150_U168,
    new_P1_R1150_U169, new_P1_R1150_U170, new_P1_R1150_U171,
    new_P1_R1150_U172, new_P1_R1150_U173, new_P1_R1150_U174,
    new_P1_R1150_U175, new_P1_R1150_U176, new_P1_R1150_U177,
    new_P1_R1150_U178, new_P1_R1150_U179, new_P1_R1150_U180,
    new_P1_R1150_U181, new_P1_R1150_U182, new_P1_R1150_U183,
    new_P1_R1150_U184, new_P1_R1150_U185, new_P1_R1150_U186,
    new_P1_R1150_U187, new_P1_R1150_U188, new_P1_R1150_U189,
    new_P1_R1150_U190, new_P1_R1150_U191, new_P1_R1150_U192,
    new_P1_R1150_U193, new_P1_R1150_U194, new_P1_R1150_U195,
    new_P1_R1150_U196, new_P1_R1150_U197, new_P1_R1150_U198,
    new_P1_R1150_U199, new_P1_R1150_U200, new_P1_R1150_U201,
    new_P1_R1150_U202, new_P1_R1150_U203, new_P1_R1150_U204,
    new_P1_R1150_U205, new_P1_R1150_U206, new_P1_R1150_U207,
    new_P1_R1150_U208, new_P1_R1150_U209, new_P1_R1150_U210,
    new_P1_R1150_U211, new_P1_R1150_U212, new_P1_R1150_U213,
    new_P1_R1150_U214, new_P1_R1150_U215, new_P1_R1150_U216,
    new_P1_R1150_U217, new_P1_R1150_U218, new_P1_R1150_U219,
    new_P1_R1150_U220, new_P1_R1150_U221, new_P1_R1150_U222,
    new_P1_R1150_U223, new_P1_R1150_U224, new_P1_R1150_U225,
    new_P1_R1150_U226, new_P1_R1150_U227, new_P1_R1150_U228,
    new_P1_R1150_U229, new_P1_R1150_U230, new_P1_R1150_U231,
    new_P1_R1150_U232, new_P1_R1150_U233, new_P1_R1150_U234,
    new_P1_R1150_U235, new_P1_R1150_U236, new_P1_R1150_U237,
    new_P1_R1150_U238, new_P1_R1150_U239, new_P1_R1150_U240,
    new_P1_R1150_U241, new_P1_R1150_U242, new_P1_R1150_U243,
    new_P1_R1150_U244, new_P1_R1150_U245, new_P1_R1150_U246,
    new_P1_R1150_U247, new_P1_R1150_U248, new_P1_R1150_U249,
    new_P1_R1150_U250, new_P1_R1150_U251, new_P1_R1150_U252,
    new_P1_R1150_U253, new_P1_R1150_U254, new_P1_R1150_U255,
    new_P1_R1150_U256, new_P1_R1150_U257, new_P1_R1150_U258,
    new_P1_R1150_U259, new_P1_R1150_U260, new_P1_R1150_U261,
    new_P1_R1150_U262, new_P1_R1150_U263, new_P1_R1150_U264,
    new_P1_R1150_U265, new_P1_R1150_U266, new_P1_R1150_U267,
    new_P1_R1150_U268, new_P1_R1150_U269, new_P1_R1150_U270,
    new_P1_R1150_U271, new_P1_R1150_U272, new_P1_R1150_U273,
    new_P1_R1150_U274, new_P1_R1150_U275, new_P1_R1150_U276,
    new_P1_R1150_U277, new_P1_R1150_U278, new_P1_R1150_U279,
    new_P1_R1150_U280, new_P1_R1150_U281, new_P1_R1150_U282,
    new_P1_R1150_U283, new_P1_R1150_U284, new_P1_R1150_U285,
    new_P1_R1150_U286, new_P1_R1150_U287, new_P1_R1150_U288,
    new_P1_R1150_U289, new_P1_R1150_U290, new_P1_R1150_U291,
    new_P1_R1150_U292, new_P1_R1150_U293, new_P1_R1150_U294,
    new_P1_R1150_U295, new_P1_R1150_U296, new_P1_R1150_U297,
    new_P1_R1150_U298, new_P1_R1150_U299, new_P1_R1150_U300,
    new_P1_R1150_U301, new_P1_R1150_U302, new_P1_R1150_U303,
    new_P1_R1150_U304, new_P1_R1150_U305, new_P1_R1150_U306,
    new_P1_R1150_U307, new_P1_R1150_U308, new_P1_R1150_U309,
    new_P1_R1150_U310, new_P1_R1150_U311, new_P1_R1150_U312,
    new_P1_R1150_U313, new_P1_R1150_U314, new_P1_R1150_U315,
    new_P1_R1150_U316, new_P1_R1150_U317, new_P1_R1150_U318,
    new_P1_R1150_U319, new_P1_R1150_U320, new_P1_R1150_U321,
    new_P1_R1150_U322, new_P1_R1150_U323, new_P1_R1150_U324,
    new_P1_R1150_U325, new_P1_R1150_U326, new_P1_R1150_U327,
    new_P1_R1150_U328, new_P1_R1150_U329, new_P1_R1150_U330,
    new_P1_R1150_U331, new_P1_R1150_U332, new_P1_R1150_U333,
    new_P1_R1150_U334, new_P1_R1150_U335, new_P1_R1150_U336,
    new_P1_R1150_U337, new_P1_R1150_U338, new_P1_R1150_U339,
    new_P1_R1150_U340, new_P1_R1150_U341, new_P1_R1150_U342,
    new_P1_R1150_U343, new_P1_R1150_U344, new_P1_R1150_U345,
    new_P1_R1150_U346, new_P1_R1150_U347, new_P1_R1150_U348,
    new_P1_R1150_U349, new_P1_R1150_U350, new_P1_R1150_U351,
    new_P1_R1150_U352, new_P1_R1150_U353, new_P1_R1150_U354,
    new_P1_R1150_U355, new_P1_R1150_U356, new_P1_R1150_U357,
    new_P1_R1150_U358, new_P1_R1150_U359, new_P1_R1150_U360,
    new_P1_R1150_U361, new_P1_R1150_U362, new_P1_R1150_U363,
    new_P1_R1150_U364, new_P1_R1150_U365, new_P1_R1150_U366,
    new_P1_R1150_U367, new_P1_R1150_U368, new_P1_R1150_U369,
    new_P1_R1150_U370, new_P1_R1150_U371, new_P1_R1150_U372,
    new_P1_R1150_U373, new_P1_R1150_U374, new_P1_R1150_U375,
    new_P1_R1150_U376, new_P1_R1150_U377, new_P1_R1150_U378,
    new_P1_R1150_U379, new_P1_R1150_U380, new_P1_R1150_U381,
    new_P1_R1150_U382, new_P1_R1150_U383, new_P1_R1150_U384,
    new_P1_R1150_U385, new_P1_R1150_U386, new_P1_R1150_U387,
    new_P1_R1150_U388, new_P1_R1150_U389, new_P1_R1150_U390,
    new_P1_R1150_U391, new_P1_R1150_U392, new_P1_R1150_U393,
    new_P1_R1150_U394, new_P1_R1150_U395, new_P1_R1150_U396,
    new_P1_R1150_U397, new_P1_R1150_U398, new_P1_R1150_U399,
    new_P1_R1150_U400, new_P1_R1150_U401, new_P1_R1150_U402,
    new_P1_R1150_U403, new_P1_R1150_U404, new_P1_R1150_U405,
    new_P1_R1150_U406, new_P1_R1150_U407, new_P1_R1150_U408,
    new_P1_R1150_U409, new_P1_R1150_U410, new_P1_R1150_U411,
    new_P1_R1150_U412, new_P1_R1150_U413, new_P1_R1150_U414,
    new_P1_R1150_U415, new_P1_R1150_U416, new_P1_R1150_U417,
    new_P1_R1150_U418, new_P1_R1150_U419, new_P1_R1150_U420,
    new_P1_R1150_U421, new_P1_R1150_U422, new_P1_R1150_U423,
    new_P1_R1150_U424, new_P1_R1150_U425, new_P1_R1150_U426,
    new_P1_R1150_U427, new_P1_R1150_U428, new_P1_R1150_U429,
    new_P1_R1150_U430, new_P1_R1150_U431, new_P1_R1150_U432,
    new_P1_R1150_U433, new_P1_R1150_U434, new_P1_R1150_U435,
    new_P1_R1150_U436, new_P1_R1150_U437, new_P1_R1150_U438,
    new_P1_R1150_U439, new_P1_R1150_U440, new_P1_R1150_U441,
    new_P1_R1150_U442, new_P1_R1150_U443, new_P1_R1150_U444,
    new_P1_R1150_U445, new_P1_R1150_U446, new_P1_R1150_U447,
    new_P1_R1150_U448, new_P1_R1150_U449, new_P1_R1150_U450,
    new_P1_R1150_U451, new_P1_R1150_U452, new_P1_R1150_U453,
    new_P1_R1150_U454, new_P1_R1150_U455, new_P1_R1150_U456,
    new_P1_R1150_U457, new_P1_R1150_U458, new_P1_R1150_U459,
    new_P1_R1150_U460, new_P1_R1150_U461, new_P1_R1150_U462,
    new_P1_R1150_U463, new_P1_R1150_U464, new_P1_R1150_U465,
    new_P1_R1150_U466, new_P1_R1150_U467, new_P1_R1150_U468,
    new_P1_R1150_U469, new_P1_R1150_U470, new_P1_R1150_U471,
    new_P1_R1150_U472, new_P1_R1150_U473, new_P1_R1150_U474,
    new_P1_R1150_U475, new_P1_R1150_U476, new_P1_R1192_U6, new_P1_R1192_U7,
    new_P1_R1192_U8, new_P1_R1192_U9, new_P1_R1192_U10, new_P1_R1192_U11,
    new_P1_R1192_U12, new_P1_R1192_U13, new_P1_R1192_U14, new_P1_R1192_U15,
    new_P1_R1192_U16, new_P1_R1192_U17, new_P1_R1192_U18, new_P1_R1192_U19,
    new_P1_R1192_U20, new_P1_R1192_U21, new_P1_R1192_U22, new_P1_R1192_U23,
    new_P1_R1192_U24, new_P1_R1192_U25, new_P1_R1192_U26, new_P1_R1192_U27,
    new_P1_R1192_U28, new_P1_R1192_U29, new_P1_R1192_U30, new_P1_R1192_U31,
    new_P1_R1192_U32, new_P1_R1192_U33, new_P1_R1192_U34, new_P1_R1192_U35,
    new_P1_R1192_U36, new_P1_R1192_U37, new_P1_R1192_U38, new_P1_R1192_U39,
    new_P1_R1192_U40, new_P1_R1192_U41, new_P1_R1192_U42, new_P1_R1192_U43,
    new_P1_R1192_U44, new_P1_R1192_U45, new_P1_R1192_U46, new_P1_R1192_U47,
    new_P1_R1192_U48, new_P1_R1192_U49, new_P1_R1192_U50, new_P1_R1192_U51,
    new_P1_R1192_U52, new_P1_R1192_U53, new_P1_R1192_U54, new_P1_R1192_U55,
    new_P1_R1192_U56, new_P1_R1192_U57, new_P1_R1192_U58, new_P1_R1192_U59,
    new_P1_R1192_U60, new_P1_R1192_U61, new_P1_R1192_U62, new_P1_R1192_U63,
    new_P1_R1192_U64, new_P1_R1192_U65, new_P1_R1192_U66, new_P1_R1192_U67,
    new_P1_R1192_U68, new_P1_R1192_U69, new_P1_R1192_U70, new_P1_R1192_U71,
    new_P1_R1192_U72, new_P1_R1192_U73, new_P1_R1192_U74, new_P1_R1192_U75,
    new_P1_R1192_U76, new_P1_R1192_U77, new_P1_R1192_U78, new_P1_R1192_U79,
    new_P1_R1192_U80, new_P1_R1192_U81, new_P1_R1192_U82, new_P1_R1192_U83,
    new_P1_R1192_U84, new_P1_R1192_U85, new_P1_R1192_U86, new_P1_R1192_U87,
    new_P1_R1192_U88, new_P1_R1192_U89, new_P1_R1192_U90, new_P1_R1192_U91,
    new_P1_R1192_U92, new_P1_R1192_U93, new_P1_R1192_U94, new_P1_R1192_U95,
    new_P1_R1192_U96, new_P1_R1192_U97, new_P1_R1192_U98, new_P1_R1192_U99,
    new_P1_R1192_U100, new_P1_R1192_U101, new_P1_R1192_U102,
    new_P1_R1192_U103, new_P1_R1192_U104, new_P1_R1192_U105,
    new_P1_R1192_U106, new_P1_R1192_U107, new_P1_R1192_U108,
    new_P1_R1192_U109, new_P1_R1192_U110, new_P1_R1192_U111,
    new_P1_R1192_U112, new_P1_R1192_U113, new_P1_R1192_U114,
    new_P1_R1192_U115, new_P1_R1192_U116, new_P1_R1192_U117,
    new_P1_R1192_U118, new_P1_R1192_U119, new_P1_R1192_U120,
    new_P1_R1192_U121, new_P1_R1192_U122, new_P1_R1192_U123,
    new_P1_R1192_U124, new_P1_R1192_U125, new_P1_R1192_U126,
    new_P1_R1192_U127, new_P1_R1192_U128, new_P1_R1192_U129,
    new_P1_R1192_U130, new_P1_R1192_U131, new_P1_R1192_U132,
    new_P1_R1192_U133, new_P1_R1192_U134, new_P1_R1192_U135,
    new_P1_R1192_U136, new_P1_R1192_U137, new_P1_R1192_U138,
    new_P1_R1192_U139, new_P1_R1192_U140, new_P1_R1192_U141,
    new_P1_R1192_U142, new_P1_R1192_U143, new_P1_R1192_U144,
    new_P1_R1192_U145, new_P1_R1192_U146, new_P1_R1192_U147,
    new_P1_R1192_U148, new_P1_R1192_U149, new_P1_R1192_U150,
    new_P1_R1192_U151, new_P1_R1192_U152, new_P1_R1192_U153,
    new_P1_R1192_U154, new_P1_R1192_U155, new_P1_R1192_U156,
    new_P1_R1192_U157, new_P1_R1192_U158, new_P1_R1192_U159,
    new_P1_R1192_U160, new_P1_R1192_U161, new_P1_R1192_U162,
    new_P1_R1192_U163, new_P1_R1192_U164, new_P1_R1192_U165,
    new_P1_R1192_U166, new_P1_R1192_U167, new_P1_R1192_U168,
    new_P1_R1192_U169, new_P1_R1192_U170, new_P1_R1192_U171,
    new_P1_R1192_U172, new_P1_R1192_U173, new_P1_R1192_U174,
    new_P1_R1192_U175, new_P1_R1192_U176, new_P1_R1192_U177,
    new_P1_R1192_U178, new_P1_R1192_U179, new_P1_R1192_U180,
    new_P1_R1192_U181, new_P1_R1192_U182, new_P1_R1192_U183,
    new_P1_R1192_U184, new_P1_R1192_U185, new_P1_R1192_U186,
    new_P1_R1192_U187, new_P1_R1192_U188, new_P1_R1192_U189,
    new_P1_R1192_U190, new_P1_R1192_U191, new_P1_R1192_U192,
    new_P1_R1192_U193, new_P1_R1192_U194, new_P1_R1192_U195,
    new_P1_R1192_U196, new_P1_R1192_U197, new_P1_R1192_U198,
    new_P1_R1192_U199, new_P1_R1192_U200, new_P1_R1192_U201,
    new_P1_R1192_U202, new_P1_R1192_U203, new_P1_R1192_U204,
    new_P1_R1192_U205, new_P1_R1192_U206, new_P1_R1192_U207,
    new_P1_R1192_U208, new_P1_R1192_U209, new_P1_R1192_U210,
    new_P1_R1192_U211, new_P1_R1192_U212, new_P1_R1192_U213,
    new_P1_R1192_U214, new_P1_R1192_U215, new_P1_R1192_U216,
    new_P1_R1192_U217, new_P1_R1192_U218, new_P1_R1192_U219,
    new_P1_R1192_U220, new_P1_R1192_U221, new_P1_R1192_U222,
    new_P1_R1192_U223, new_P1_R1192_U224, new_P1_R1192_U225,
    new_P1_R1192_U226, new_P1_R1192_U227, new_P1_R1192_U228,
    new_P1_R1192_U229, new_P1_R1192_U230, new_P1_R1192_U231,
    new_P1_R1192_U232, new_P1_R1192_U233, new_P1_R1192_U234,
    new_P1_R1192_U235, new_P1_R1192_U236, new_P1_R1192_U237,
    new_P1_R1192_U238, new_P1_R1192_U239, new_P1_R1192_U240,
    new_P1_R1192_U241, new_P1_R1192_U242, new_P1_R1192_U243,
    new_P1_R1192_U244, new_P1_R1192_U245, new_P1_R1192_U246,
    new_P1_R1192_U247, new_P1_R1192_U248, new_P1_R1192_U249,
    new_P1_R1192_U250, new_P1_R1192_U251, new_P1_R1192_U252,
    new_P1_R1192_U253, new_P1_R1192_U254, new_P1_R1192_U255,
    new_P1_R1192_U256, new_P1_R1192_U257, new_P1_R1192_U258,
    new_P1_R1192_U259, new_P1_R1192_U260, new_P1_R1192_U261,
    new_P1_R1192_U262, new_P1_R1192_U263, new_P1_R1192_U264,
    new_P1_R1192_U265, new_P1_R1192_U266, new_P1_R1192_U267,
    new_P1_R1192_U268, new_P1_R1192_U269, new_P1_R1192_U270,
    new_P1_R1192_U271, new_P1_R1192_U272, new_P1_R1192_U273,
    new_P1_R1192_U274, new_P1_R1192_U275, new_P1_R1192_U276,
    new_P1_R1192_U277, new_P1_R1192_U278, new_P1_R1192_U279,
    new_P1_R1192_U280, new_P1_R1192_U281, new_P1_R1192_U282,
    new_P1_R1192_U283, new_P1_R1192_U284, new_P1_R1192_U285,
    new_P1_R1192_U286, new_P1_R1192_U287, new_P1_R1192_U288,
    new_P1_R1192_U289, new_P1_R1192_U290, new_P1_R1192_U291,
    new_P1_R1192_U292, new_P1_R1192_U293, new_P1_R1192_U294,
    new_P1_R1192_U295, new_P1_R1192_U296, new_P1_R1192_U297,
    new_P1_R1192_U298, new_P1_R1192_U299, new_P1_R1192_U300,
    new_P1_R1192_U301, new_P1_R1192_U302, new_P1_R1192_U303,
    new_P1_R1192_U304, new_P1_R1192_U305, new_P1_R1192_U306,
    new_P1_R1192_U307, new_P1_R1192_U308, new_P1_R1192_U309,
    new_P1_R1192_U310, new_P1_R1192_U311, new_P1_R1192_U312,
    new_P1_R1192_U313, new_P1_R1192_U314, new_P1_R1192_U315,
    new_P1_R1192_U316, new_P1_R1192_U317, new_P1_R1192_U318,
    new_P1_R1192_U319, new_P1_R1192_U320, new_P1_R1192_U321,
    new_P1_R1192_U322, new_P1_R1192_U323, new_P1_R1192_U324,
    new_P1_R1192_U325, new_P1_R1192_U326, new_P1_R1192_U327,
    new_P1_R1192_U328, new_P1_R1192_U329, new_P1_R1192_U330,
    new_P1_R1192_U331, new_P1_R1192_U332, new_P1_R1192_U333,
    new_P1_R1192_U334, new_P1_R1192_U335, new_P1_R1192_U336,
    new_P1_R1192_U337, new_P1_R1192_U338, new_P1_R1192_U339,
    new_P1_R1192_U340, new_P1_R1192_U341, new_P1_R1192_U342,
    new_P1_R1192_U343, new_P1_R1192_U344, new_P1_R1192_U345,
    new_P1_R1192_U346, new_P1_R1192_U347, new_P1_R1192_U348,
    new_P1_R1192_U349, new_P1_R1192_U350, new_P1_R1192_U351,
    new_P1_R1192_U352, new_P1_R1192_U353, new_P1_R1192_U354,
    new_P1_R1192_U355, new_P1_R1192_U356, new_P1_R1192_U357,
    new_P1_R1192_U358, new_P1_R1192_U359, new_P1_R1192_U360,
    new_P1_R1192_U361, new_P1_R1192_U362, new_P1_R1192_U363,
    new_P1_R1192_U364, new_P1_R1192_U365, new_P1_R1192_U366,
    new_P1_R1192_U367, new_P1_R1192_U368, new_P1_R1192_U369,
    new_P1_R1192_U370, new_P1_R1192_U371, new_P1_R1192_U372,
    new_P1_R1192_U373, new_P1_R1192_U374, new_P1_R1192_U375,
    new_P1_R1192_U376, new_P1_R1192_U377, new_P1_R1192_U378,
    new_P1_R1192_U379, new_P1_R1192_U380, new_P1_R1192_U381,
    new_P1_R1192_U382, new_P1_R1192_U383, new_P1_R1192_U384,
    new_P1_R1192_U385, new_P1_R1192_U386, new_P1_R1192_U387,
    new_P1_R1192_U388, new_P1_R1192_U389, new_P1_R1192_U390,
    new_P1_R1192_U391, new_P1_R1192_U392, new_P1_R1192_U393,
    new_P1_R1192_U394, new_P1_R1192_U395, new_P1_R1192_U396,
    new_P1_R1192_U397, new_P1_R1192_U398, new_P1_R1192_U399,
    new_P1_R1192_U400, new_P1_R1192_U401, new_P1_R1192_U402,
    new_P1_R1192_U403, new_P1_R1192_U404, new_P1_R1192_U405,
    new_P1_R1192_U406, new_P1_R1192_U407, new_P1_R1192_U408,
    new_P1_R1192_U409, new_P1_R1192_U410, new_P1_R1192_U411,
    new_P1_R1192_U412, new_P1_R1192_U413, new_P1_R1192_U414,
    new_P1_R1192_U415, new_P1_R1192_U416, new_P1_R1192_U417,
    new_P1_R1192_U418, new_P1_R1192_U419, new_P1_R1192_U420,
    new_P1_R1192_U421, new_P1_R1192_U422, new_P1_R1192_U423,
    new_P1_R1192_U424, new_P1_R1192_U425, new_P1_R1192_U426,
    new_P1_R1192_U427, new_P1_R1192_U428, new_P1_R1192_U429,
    new_P1_R1192_U430, new_P1_R1192_U431, new_P1_R1192_U432,
    new_P1_R1192_U433, new_P1_R1192_U434, new_P1_R1192_U435,
    new_P1_R1192_U436, new_P1_R1192_U437, new_P1_R1192_U438,
    new_P1_R1192_U439, new_P1_R1192_U440, new_P1_R1192_U441,
    new_P1_R1192_U442, new_P1_R1192_U443, new_P1_R1192_U444,
    new_P1_R1192_U445, new_P1_R1192_U446, new_P1_R1192_U447,
    new_P1_R1192_U448, new_P1_R1192_U449, new_P1_R1192_U450,
    new_P1_R1192_U451, new_P1_R1192_U452, new_P1_R1192_U453,
    new_P1_R1192_U454, new_P1_R1192_U455, new_P1_R1192_U456,
    new_P1_R1192_U457, new_P1_R1192_U458, new_P1_R1192_U459,
    new_P1_R1192_U460, new_P1_R1192_U461, new_P1_R1192_U462,
    new_P1_R1192_U463, new_P1_R1192_U464, new_P1_R1192_U465,
    new_P1_R1192_U466, new_P1_R1192_U467, new_P1_R1192_U468,
    new_P1_R1192_U469, new_P1_R1192_U470, new_P1_R1192_U471,
    new_P1_R1192_U472, new_P1_R1192_U473, new_P1_R1192_U474,
    new_P1_R1192_U475, new_P1_R1192_U476, new_P1_R1171_U4, new_P1_R1171_U5,
    new_P1_R1171_U6, new_P1_R1171_U7, new_P1_R1171_U8, new_P1_R1171_U9,
    new_P1_R1171_U10, new_P1_R1171_U11, new_P1_R1171_U12, new_P1_R1171_U13,
    new_P1_R1171_U14, new_P1_R1171_U15, new_P1_R1171_U16, new_P1_R1171_U17,
    new_P1_R1171_U18, new_P1_R1171_U19, new_P1_R1171_U20, new_P1_R1171_U21,
    new_P1_R1171_U22, new_P1_R1171_U23, new_P1_R1171_U24, new_P1_R1171_U25,
    new_P1_R1171_U26, new_P1_R1171_U27, new_P1_R1171_U28, new_P1_R1171_U29,
    new_P1_R1171_U30, new_P1_R1171_U31, new_P1_R1171_U32, new_P1_R1171_U33,
    new_P1_R1171_U34, new_P1_R1171_U35, new_P1_R1171_U36, new_P1_R1171_U37,
    new_P1_R1171_U38, new_P1_R1171_U39, new_P1_R1171_U40, new_P1_R1171_U41,
    new_P1_R1171_U42, new_P1_R1171_U43, new_P1_R1171_U44, new_P1_R1171_U45,
    new_P1_R1171_U46, new_P1_R1171_U47, new_P1_R1171_U48, new_P1_R1171_U49,
    new_P1_R1171_U50, new_P1_R1171_U51, new_P1_R1171_U52, new_P1_R1171_U53,
    new_P1_R1171_U54, new_P1_R1171_U55, new_P1_R1171_U56, new_P1_R1171_U57,
    new_P1_R1171_U58, new_P1_R1171_U59, new_P1_R1171_U60, new_P1_R1171_U61,
    new_P1_R1171_U62, new_P1_R1171_U63, new_P1_R1171_U64, new_P1_R1171_U65,
    new_P1_R1171_U66, new_P1_R1171_U67, new_P1_R1171_U68, new_P1_R1171_U69,
    new_P1_R1171_U70, new_P1_R1171_U71, new_P1_R1171_U72, new_P1_R1171_U73,
    new_P1_R1171_U74, new_P1_R1171_U75, new_P1_R1171_U76, new_P1_R1171_U77,
    new_P1_R1171_U78, new_P1_R1171_U79, new_P1_R1171_U80, new_P1_R1171_U81,
    new_P1_R1171_U82, new_P1_R1171_U83, new_P1_R1171_U84, new_P1_R1171_U85,
    new_P1_R1171_U86, new_P1_R1171_U87, new_P1_R1171_U88, new_P1_R1171_U89,
    new_P1_R1171_U90, new_P1_R1171_U91, new_P1_R1171_U92, new_P1_R1171_U93,
    new_P1_R1171_U94, new_P1_R1171_U95, new_P1_R1171_U96, new_P1_R1171_U97,
    new_P1_R1171_U98, new_P1_R1171_U99, new_P1_R1171_U100,
    new_P1_R1171_U101, new_P1_R1171_U102, new_P1_R1171_U103,
    new_P1_R1171_U104, new_P1_R1171_U105, new_P1_R1171_U106,
    new_P1_R1171_U107, new_P1_R1171_U108, new_P1_R1171_U109,
    new_P1_R1171_U110, new_P1_R1171_U111, new_P1_R1171_U112,
    new_P1_R1171_U113, new_P1_R1171_U114, new_P1_R1171_U115,
    new_P1_R1171_U116, new_P1_R1171_U117, new_P1_R1171_U118,
    new_P1_R1171_U119, new_P1_R1171_U120, new_P1_R1171_U121,
    new_P1_R1171_U122, new_P1_R1171_U123, new_P1_R1171_U124,
    new_P1_R1171_U125, new_P1_R1171_U126, new_P1_R1171_U127,
    new_P1_R1171_U128, new_P1_R1171_U129, new_P1_R1171_U130,
    new_P1_R1171_U131, new_P1_R1171_U132, new_P1_R1171_U133,
    new_P1_R1171_U134, new_P1_R1171_U135, new_P1_R1171_U136,
    new_P1_R1171_U137, new_P1_R1171_U138, new_P1_R1171_U139,
    new_P1_R1171_U140, new_P1_R1171_U141, new_P1_R1171_U142,
    new_P1_R1171_U143, new_P1_R1171_U144, new_P1_R1171_U145,
    new_P1_R1171_U146, new_P1_R1171_U147, new_P1_R1171_U148,
    new_P1_R1171_U149, new_P1_R1171_U150, new_P1_R1171_U151,
    new_P1_R1171_U152, new_P1_R1171_U153, new_P1_R1171_U154,
    new_P1_R1171_U155, new_P1_R1171_U156, new_P1_R1171_U157,
    new_P1_R1171_U158, new_P1_R1171_U159, new_P1_R1171_U160,
    new_P1_R1171_U161, new_P1_R1171_U162, new_P1_R1171_U163,
    new_P1_R1171_U164, new_P1_R1171_U165, new_P1_R1171_U166,
    new_P1_R1171_U167, new_P1_R1171_U168, new_P1_R1171_U169,
    new_P1_R1171_U170, new_P1_R1171_U171, new_P1_R1171_U172,
    new_P1_R1171_U173, new_P1_R1171_U174, new_P1_R1171_U175,
    new_P1_R1171_U176, new_P1_R1171_U177, new_P1_R1171_U178,
    new_P1_R1171_U179, new_P1_R1171_U180, new_P1_R1171_U181,
    new_P1_R1171_U182, new_P1_R1171_U183, new_P1_R1171_U184,
    new_P1_R1171_U185, new_P1_R1171_U186, new_P1_R1171_U187,
    new_P1_R1171_U188, new_P1_R1171_U189, new_P1_R1171_U190,
    new_P1_R1171_U191, new_P1_R1171_U192, new_P1_R1171_U193,
    new_P1_R1171_U194, new_P1_R1171_U195, new_P1_R1171_U196,
    new_P1_R1171_U197, new_P1_R1171_U198, new_P1_R1171_U199,
    new_P1_R1171_U200, new_P1_R1171_U201, new_P1_R1171_U202,
    new_P1_R1171_U203, new_P1_R1171_U204, new_P1_R1171_U205,
    new_P1_R1171_U206, new_P1_R1171_U207, new_P1_R1171_U208,
    new_P1_R1171_U209, new_P1_R1171_U210, new_P1_R1171_U211,
    new_P1_R1171_U212, new_P1_R1171_U213, new_P1_R1171_U214,
    new_P1_R1171_U215, new_P1_R1171_U216, new_P1_R1171_U217,
    new_P1_R1171_U218, new_P1_R1171_U219, new_P1_R1171_U220,
    new_P1_R1171_U221, new_P1_R1171_U222, new_P1_R1171_U223,
    new_P1_R1171_U224, new_P1_R1171_U225, new_P1_R1171_U226,
    new_P1_R1171_U227, new_P1_R1171_U228, new_P1_R1171_U229,
    new_P1_R1171_U230, new_P1_R1171_U231, new_P1_R1171_U232,
    new_P1_R1171_U233, new_P1_R1171_U234, new_P1_R1171_U235,
    new_P1_R1171_U236, new_P1_R1171_U237, new_P1_R1171_U238,
    new_P1_R1171_U239, new_P1_R1171_U240, new_P1_R1171_U241,
    new_P1_R1171_U242, new_P1_R1171_U243, new_P1_R1171_U244,
    new_P1_R1171_U245, new_P1_R1171_U246, new_P1_R1171_U247,
    new_P1_R1171_U248, new_P1_R1171_U249, new_P1_R1171_U250,
    new_P1_R1171_U251, new_P1_R1171_U252, new_P1_R1171_U253,
    new_P1_R1171_U254, new_P1_R1171_U255, new_P1_R1171_U256,
    new_P1_R1171_U257, new_P1_R1171_U258, new_P1_R1171_U259,
    new_P1_R1171_U260, new_P1_R1171_U261, new_P1_R1171_U262,
    new_P1_R1171_U263, new_P1_R1171_U264, new_P1_R1171_U265,
    new_P1_R1171_U266, new_P1_R1171_U267, new_P1_R1171_U268,
    new_P1_R1171_U269, new_P1_R1171_U270, new_P1_R1171_U271,
    new_P1_R1171_U272, new_P1_R1171_U273, new_P1_R1171_U274,
    new_P1_R1171_U275, new_P1_R1171_U276, new_P1_R1171_U277,
    new_P1_R1171_U278, new_P1_R1171_U279, new_P1_R1171_U280,
    new_P1_R1171_U281, new_P1_R1171_U282, new_P1_R1171_U283,
    new_P1_R1171_U284, new_P1_R1171_U285, new_P1_R1171_U286,
    new_P1_R1171_U287, new_P1_R1171_U288, new_P1_R1171_U289,
    new_P1_R1171_U290, new_P1_R1171_U291, new_P1_R1171_U292,
    new_P1_R1171_U293, new_P1_R1171_U294, new_P1_R1171_U295,
    new_P1_R1171_U296, new_P1_R1171_U297, new_P1_R1171_U298,
    new_P1_R1171_U299, new_P1_R1171_U300, new_P1_R1171_U301,
    new_P1_R1171_U302, new_P1_R1171_U303, new_P1_R1171_U304,
    new_P1_R1171_U305, new_P1_R1171_U306, new_P1_R1171_U307,
    new_P1_R1171_U308, new_P1_R1171_U309, new_P1_R1171_U310,
    new_P1_R1171_U311, new_P1_R1171_U312, new_P1_R1171_U313,
    new_P1_R1171_U314, new_P1_R1171_U315, new_P1_R1171_U316,
    new_P1_R1171_U317, new_P1_R1171_U318, new_P1_R1171_U319,
    new_P1_R1171_U320, new_P1_R1171_U321, new_P1_R1171_U322,
    new_P1_R1171_U323, new_P1_R1171_U324, new_P1_R1171_U325,
    new_P1_R1171_U326, new_P1_R1171_U327, new_P1_R1171_U328,
    new_P1_R1171_U329, new_P1_R1171_U330, new_P1_R1171_U331,
    new_P1_R1171_U332, new_P1_R1171_U333, new_P1_R1171_U334,
    new_P1_R1171_U335, new_P1_R1171_U336, new_P1_R1171_U337,
    new_P1_R1171_U338, new_P1_R1171_U339, new_P1_R1171_U340,
    new_P1_R1171_U341, new_P1_R1171_U342, new_P1_R1171_U343,
    new_P1_R1171_U344, new_P1_R1171_U345, new_P1_R1171_U346,
    new_P1_R1171_U347, new_P1_R1171_U348, new_P1_R1171_U349,
    new_P1_R1171_U350, new_P1_R1171_U351, new_P1_R1171_U352,
    new_P1_R1171_U353, new_P1_R1171_U354, new_P1_R1171_U355,
    new_P1_R1171_U356, new_P1_R1171_U357, new_P1_R1171_U358,
    new_P1_R1171_U359, new_P1_R1171_U360, new_P1_R1171_U361,
    new_P1_R1171_U362, new_P1_R1171_U363, new_P1_R1171_U364,
    new_P1_R1171_U365, new_P1_R1171_U366, new_P1_R1171_U367,
    new_P1_R1171_U368, new_P1_R1171_U369, new_P1_R1171_U370,
    new_P1_R1171_U371, new_P1_R1171_U372, new_P1_R1171_U373,
    new_P1_R1171_U374, new_P1_R1171_U375, new_P1_R1171_U376,
    new_P1_R1171_U377, new_P1_R1171_U378, new_P1_R1171_U379,
    new_P1_R1171_U380, new_P1_R1171_U381, new_P1_R1171_U382,
    new_P1_R1171_U383, new_P1_R1171_U384, new_P1_R1171_U385,
    new_P1_R1171_U386, new_P1_R1171_U387, new_P1_R1171_U388,
    new_P1_R1171_U389, new_P1_R1171_U390, new_P1_R1171_U391,
    new_P1_R1171_U392, new_P1_R1171_U393, new_P1_R1171_U394,
    new_P1_R1171_U395, new_P1_R1171_U396, new_P1_R1171_U397,
    new_P1_R1171_U398, new_P1_R1171_U399, new_P1_R1171_U400,
    new_P1_R1171_U401, new_P1_R1171_U402, new_P1_R1171_U403,
    new_P1_R1171_U404, new_P1_R1171_U405, new_P1_R1171_U406,
    new_P1_R1171_U407, new_P1_R1171_U408, new_P1_R1171_U409,
    new_P1_R1171_U410, new_P1_R1171_U411, new_P1_R1171_U412,
    new_P1_R1171_U413, new_P1_R1171_U414, new_P1_R1171_U415,
    new_P1_R1171_U416, new_P1_R1171_U417, new_P1_R1171_U418,
    new_P1_R1171_U419, new_P1_R1171_U420, new_P1_R1171_U421,
    new_P1_R1171_U422, new_P1_R1171_U423, new_P1_R1171_U424,
    new_P1_R1171_U425, new_P1_R1171_U426, new_P1_R1171_U427,
    new_P1_R1171_U428, new_P1_R1171_U429, new_P1_R1171_U430,
    new_P1_R1171_U431, new_P1_R1171_U432, new_P1_R1171_U433,
    new_P1_R1171_U434, new_P1_R1171_U435, new_P1_R1171_U436,
    new_P1_R1171_U437, new_P1_R1171_U438, new_P1_R1171_U439,
    new_P1_R1171_U440, new_P1_R1171_U441, new_P1_R1171_U442,
    new_P1_R1171_U443, new_P1_R1171_U444, new_P1_R1171_U445,
    new_P1_R1171_U446, new_P1_R1171_U447, new_P1_R1171_U448,
    new_P1_R1171_U449, new_P1_R1171_U450, new_P1_R1171_U451,
    new_P1_R1171_U452, new_P1_R1171_U453, new_P1_R1171_U454,
    new_P1_R1171_U455, new_P1_R1171_U456, new_P1_R1171_U457,
    new_P1_R1171_U458, new_P1_R1171_U459, new_P1_R1171_U460,
    new_P1_R1171_U461, new_P1_R1171_U462, new_P1_R1171_U463,
    new_P1_R1171_U464, new_P1_R1171_U465, new_P1_R1171_U466,
    new_P1_R1171_U467, new_P1_R1171_U468, new_P1_R1171_U469,
    new_P1_R1171_U470, new_P1_R1171_U471, new_P1_R1171_U472,
    new_P1_R1171_U473, new_P1_R1171_U474, new_P1_R1171_U475,
    new_P1_R1171_U476, new_P1_R1171_U477, new_P1_R1171_U478,
    new_P1_R1171_U479, new_P1_R1171_U480, new_P1_R1171_U481,
    new_P1_R1171_U482, new_P1_R1171_U483, new_P1_R1171_U484,
    new_P1_R1171_U485, new_P1_R1171_U486, new_P1_R1171_U487,
    new_P1_R1171_U488, new_P1_R1171_U489, new_P1_R1171_U490,
    new_P1_R1171_U491, new_P1_R1171_U492, new_P1_R1171_U493,
    new_P1_R1171_U494, new_P1_R1171_U495, new_P1_R1171_U496,
    new_P1_R1171_U497, new_P1_R1171_U498, new_P1_R1171_U499,
    new_P1_R1171_U500, new_P1_R1171_U501, new_P1_R1138_U4, new_P1_R1138_U5,
    new_P1_R1138_U6, new_P1_R1138_U7, new_P1_R1138_U8, new_P1_R1138_U9,
    new_P1_R1138_U10, new_P1_R1138_U11, new_P1_R1138_U12, new_P1_R1138_U13,
    new_P1_R1138_U14, new_P1_R1138_U15, new_P1_R1138_U16, new_P1_R1138_U17,
    new_P1_R1138_U18, new_P1_R1138_U19, new_P1_R1138_U20, new_P1_R1138_U21,
    new_P1_R1138_U22, new_P1_R1138_U23, new_P1_R1138_U24, new_P1_R1138_U25,
    new_P1_R1138_U26, new_P1_R1138_U27, new_P1_R1138_U28, new_P1_R1138_U29,
    new_P1_R1138_U30, new_P1_R1138_U31, new_P1_R1138_U32, new_P1_R1138_U33,
    new_P1_R1138_U34, new_P1_R1138_U35, new_P1_R1138_U36, new_P1_R1138_U37,
    new_P1_R1138_U38, new_P1_R1138_U39, new_P1_R1138_U40, new_P1_R1138_U41,
    new_P1_R1138_U42, new_P1_R1138_U43, new_P1_R1138_U44, new_P1_R1138_U45,
    new_P1_R1138_U46, new_P1_R1138_U47, new_P1_R1138_U48, new_P1_R1138_U49,
    new_P1_R1138_U50, new_P1_R1138_U51, new_P1_R1138_U52, new_P1_R1138_U53,
    new_P1_R1138_U54, new_P1_R1138_U55, new_P1_R1138_U56, new_P1_R1138_U57,
    new_P1_R1138_U58, new_P1_R1138_U59, new_P1_R1138_U60, new_P1_R1138_U61,
    new_P1_R1138_U62, new_P1_R1138_U63, new_P1_R1138_U64, new_P1_R1138_U65,
    new_P1_R1138_U66, new_P1_R1138_U67, new_P1_R1138_U68, new_P1_R1138_U69,
    new_P1_R1138_U70, new_P1_R1138_U71, new_P1_R1138_U72, new_P1_R1138_U73,
    new_P1_R1138_U74, new_P1_R1138_U75, new_P1_R1138_U76, new_P1_R1138_U77,
    new_P1_R1138_U78, new_P1_R1138_U79, new_P1_R1138_U80, new_P1_R1138_U81,
    new_P1_R1138_U82, new_P1_R1138_U83, new_P1_R1138_U84, new_P1_R1138_U85,
    new_P1_R1138_U86, new_P1_R1138_U87, new_P1_R1138_U88, new_P1_R1138_U89,
    new_P1_R1138_U90, new_P1_R1138_U91, new_P1_R1138_U92, new_P1_R1138_U93,
    new_P1_R1138_U94, new_P1_R1138_U95, new_P1_R1138_U96, new_P1_R1138_U97,
    new_P1_R1138_U98, new_P1_R1138_U99, new_P1_R1138_U100,
    new_P1_R1138_U101, new_P1_R1138_U102, new_P1_R1138_U103,
    new_P1_R1138_U104, new_P1_R1138_U105, new_P1_R1138_U106,
    new_P1_R1138_U107, new_P1_R1138_U108, new_P1_R1138_U109,
    new_P1_R1138_U110, new_P1_R1138_U111, new_P1_R1138_U112,
    new_P1_R1138_U113, new_P1_R1138_U114, new_P1_R1138_U115,
    new_P1_R1138_U116, new_P1_R1138_U117, new_P1_R1138_U118,
    new_P1_R1138_U119, new_P1_R1138_U120, new_P1_R1138_U121,
    new_P1_R1138_U122, new_P1_R1138_U123, new_P1_R1138_U124,
    new_P1_R1138_U125, new_P1_R1138_U126, new_P1_R1138_U127,
    new_P1_R1138_U128, new_P1_R1138_U129, new_P1_R1138_U130,
    new_P1_R1138_U131, new_P1_R1138_U132, new_P1_R1138_U133,
    new_P1_R1138_U134, new_P1_R1138_U135, new_P1_R1138_U136,
    new_P1_R1138_U137, new_P1_R1138_U138, new_P1_R1138_U139,
    new_P1_R1138_U140, new_P1_R1138_U141, new_P1_R1138_U142,
    new_P1_R1138_U143, new_P1_R1138_U144, new_P1_R1138_U145,
    new_P1_R1138_U146, new_P1_R1138_U147, new_P1_R1138_U148,
    new_P1_R1138_U149, new_P1_R1138_U150, new_P1_R1138_U151,
    new_P1_R1138_U152, new_P1_R1138_U153, new_P1_R1138_U154,
    new_P1_R1138_U155, new_P1_R1138_U156, new_P1_R1138_U157,
    new_P1_R1138_U158, new_P1_R1138_U159, new_P1_R1138_U160,
    new_P1_R1138_U161, new_P1_R1138_U162, new_P1_R1138_U163,
    new_P1_R1138_U164, new_P1_R1138_U165, new_P1_R1138_U166,
    new_P1_R1138_U167, new_P1_R1138_U168, new_P1_R1138_U169,
    new_P1_R1138_U170, new_P1_R1138_U171, new_P1_R1138_U172,
    new_P1_R1138_U173, new_P1_R1138_U174, new_P1_R1138_U175,
    new_P1_R1138_U176, new_P1_R1138_U177, new_P1_R1138_U178,
    new_P1_R1138_U179, new_P1_R1138_U180, new_P1_R1138_U181,
    new_P1_R1138_U182, new_P1_R1138_U183, new_P1_R1138_U184,
    new_P1_R1138_U185, new_P1_R1138_U186, new_P1_R1138_U187,
    new_P1_R1138_U188, new_P1_R1138_U189, new_P1_R1138_U190,
    new_P1_R1138_U191, new_P1_R1138_U192, new_P1_R1138_U193,
    new_P1_R1138_U194, new_P1_R1138_U195, new_P1_R1138_U196,
    new_P1_R1138_U197, new_P1_R1138_U198, new_P1_R1138_U199,
    new_P1_R1138_U200, new_P1_R1138_U201, new_P1_R1138_U202,
    new_P1_R1138_U203, new_P1_R1138_U204, new_P1_R1138_U205,
    new_P1_R1138_U206, new_P1_R1138_U207, new_P1_R1138_U208,
    new_P1_R1138_U209, new_P1_R1138_U210, new_P1_R1138_U211,
    new_P1_R1138_U212, new_P1_R1138_U213, new_P1_R1138_U214,
    new_P1_R1138_U215, new_P1_R1138_U216, new_P1_R1138_U217,
    new_P1_R1138_U218, new_P1_R1138_U219, new_P1_R1138_U220,
    new_P1_R1138_U221, new_P1_R1138_U222, new_P1_R1138_U223,
    new_P1_R1138_U224, new_P1_R1138_U225, new_P1_R1138_U226,
    new_P1_R1138_U227, new_P1_R1138_U228, new_P1_R1138_U229,
    new_P1_R1138_U230, new_P1_R1138_U231, new_P1_R1138_U232,
    new_P1_R1138_U233, new_P1_R1138_U234, new_P1_R1138_U235,
    new_P1_R1138_U236, new_P1_R1138_U237, new_P1_R1138_U238,
    new_P1_R1138_U239, new_P1_R1138_U240, new_P1_R1138_U241,
    new_P1_R1138_U242, new_P1_R1138_U243, new_P1_R1138_U244,
    new_P1_R1138_U245, new_P1_R1138_U246, new_P1_R1138_U247,
    new_P1_R1138_U248, new_P1_R1138_U249, new_P1_R1138_U250,
    new_P1_R1138_U251, new_P1_R1138_U252, new_P1_R1138_U253,
    new_P1_R1138_U254, new_P1_R1138_U255, new_P1_R1138_U256,
    new_P1_R1138_U257, new_P1_R1138_U258, new_P1_R1138_U259,
    new_P1_R1138_U260, new_P1_R1138_U261, new_P1_R1138_U262,
    new_P1_R1138_U263, new_P1_R1138_U264, new_P1_R1138_U265,
    new_P1_R1138_U266, new_P1_R1138_U267, new_P1_R1138_U268,
    new_P1_R1138_U269, new_P1_R1138_U270, new_P1_R1138_U271,
    new_P1_R1138_U272, new_P1_R1138_U273, new_P1_R1138_U274,
    new_P1_R1138_U275, new_P1_R1138_U276, new_P1_R1138_U277,
    new_P1_R1138_U278, new_P1_R1138_U279, new_P1_R1138_U280,
    new_P1_R1138_U281, new_P1_R1138_U282, new_P1_R1138_U283,
    new_P1_R1138_U284, new_P1_R1138_U285, new_P1_R1138_U286,
    new_P1_R1138_U287, new_P1_R1138_U288, new_P1_R1138_U289,
    new_P1_R1138_U290, new_P1_R1138_U291, new_P1_R1138_U292,
    new_P1_R1138_U293, new_P1_R1138_U294, new_P1_R1138_U295,
    new_P1_R1138_U296, new_P1_R1138_U297, new_P1_R1138_U298,
    new_P1_R1138_U299, new_P1_R1138_U300, new_P1_R1138_U301,
    new_P1_R1138_U302, new_P1_R1138_U303, new_P1_R1138_U304,
    new_P1_R1138_U305, new_P1_R1138_U306, new_P1_R1138_U307,
    new_P1_R1138_U308, new_P1_R1138_U309, new_P1_R1138_U310,
    new_P1_R1138_U311, new_P1_R1138_U312, new_P1_R1138_U313,
    new_P1_R1138_U314, new_P1_R1138_U315, new_P1_R1138_U316,
    new_P1_R1138_U317, new_P1_R1138_U318, new_P1_R1138_U319,
    new_P1_R1138_U320, new_P1_R1138_U321, new_P1_R1138_U322,
    new_P1_R1138_U323, new_P1_R1138_U324, new_P1_R1138_U325,
    new_P1_R1138_U326, new_P1_R1138_U327, new_P1_R1138_U328,
    new_P1_R1138_U329, new_P1_R1138_U330, new_P1_R1138_U331,
    new_P1_R1138_U332, new_P1_R1138_U333, new_P1_R1138_U334,
    new_P1_R1138_U335, new_P1_R1138_U336, new_P1_R1138_U337,
    new_P1_R1138_U338, new_P1_R1138_U339, new_P1_R1138_U340,
    new_P1_R1138_U341, new_P1_R1138_U342, new_P1_R1138_U343,
    new_P1_R1138_U344, new_P1_R1138_U345, new_P1_R1138_U346,
    new_P1_R1138_U347, new_P1_R1138_U348, new_P1_R1138_U349,
    new_P1_R1138_U350, new_P1_R1138_U351, new_P1_R1138_U352,
    new_P1_R1138_U353, new_P1_R1138_U354, new_P1_R1138_U355,
    new_P1_R1138_U356, new_P1_R1138_U357, new_P1_R1138_U358,
    new_P1_R1138_U359, new_P1_R1138_U360, new_P1_R1138_U361,
    new_P1_R1138_U362, new_P1_R1138_U363, new_P1_R1138_U364,
    new_P1_R1138_U365, new_P1_R1138_U366, new_P1_R1138_U367,
    new_P1_R1138_U368, new_P1_R1138_U369, new_P1_R1138_U370,
    new_P1_R1138_U371, new_P1_R1138_U372, new_P1_R1138_U373,
    new_P1_R1138_U374, new_P1_R1138_U375, new_P1_R1138_U376,
    new_P1_R1138_U377, new_P1_R1138_U378, new_P1_R1138_U379,
    new_P1_R1138_U380, new_P1_R1138_U381, new_P1_R1138_U382,
    new_P1_R1138_U383, new_P1_R1138_U384, new_P1_R1138_U385,
    new_P1_R1138_U386, new_P1_R1138_U387, new_P1_R1138_U388,
    new_P1_R1138_U389, new_P1_R1138_U390, new_P1_R1138_U391,
    new_P1_R1138_U392, new_P1_R1138_U393, new_P1_R1138_U394,
    new_P1_R1138_U395, new_P1_R1138_U396, new_P1_R1138_U397,
    new_P1_R1138_U398, new_P1_R1138_U399, new_P1_R1138_U400,
    new_P1_R1138_U401, new_P1_R1138_U402, new_P1_R1138_U403,
    new_P1_R1138_U404, new_P1_R1138_U405, new_P1_R1138_U406,
    new_P1_R1138_U407, new_P1_R1138_U408, new_P1_R1138_U409,
    new_P1_R1138_U410, new_P1_R1138_U411, new_P1_R1138_U412,
    new_P1_R1138_U413, new_P1_R1138_U414, new_P1_R1138_U415,
    new_P1_R1138_U416, new_P1_R1138_U417, new_P1_R1138_U418,
    new_P1_R1138_U419, new_P1_R1138_U420, new_P1_R1138_U421,
    new_P1_R1138_U422, new_P1_R1138_U423, new_P1_R1138_U424,
    new_P1_R1138_U425, new_P1_R1138_U426, new_P1_R1138_U427,
    new_P1_R1138_U428, new_P1_R1138_U429, new_P1_R1138_U430,
    new_P1_R1138_U431, new_P1_R1138_U432, new_P1_R1138_U433,
    new_P1_R1138_U434, new_P1_R1138_U435, new_P1_R1138_U436,
    new_P1_R1138_U437, new_P1_R1138_U438, new_P1_R1138_U439,
    new_P1_R1138_U440, new_P1_R1138_U441, new_P1_R1138_U442,
    new_P1_R1138_U443, new_P1_R1138_U444, new_P1_R1138_U445,
    new_P1_R1138_U446, new_P1_R1138_U447, new_P1_R1138_U448,
    new_P1_R1138_U449, new_P1_R1138_U450, new_P1_R1138_U451,
    new_P1_R1138_U452, new_P1_R1138_U453, new_P1_R1138_U454,
    new_P1_R1138_U455, new_P1_R1138_U456, new_P1_R1138_U457,
    new_P1_R1138_U458, new_P1_R1138_U459, new_P1_R1138_U460,
    new_P1_R1138_U461, new_P1_R1138_U462, new_P1_R1138_U463,
    new_P1_R1138_U464, new_P1_R1138_U465, new_P1_R1138_U466,
    new_P1_R1138_U467, new_P1_R1138_U468, new_P1_R1138_U469,
    new_P1_R1138_U470, new_P1_R1138_U471, new_P1_R1138_U472,
    new_P1_R1138_U473, new_P1_R1138_U474, new_P1_R1138_U475,
    new_P1_R1138_U476, new_P1_R1138_U477, new_P1_R1138_U478,
    new_P1_R1138_U479, new_P1_R1138_U480, new_P1_R1138_U481,
    new_P1_R1138_U482, new_P1_R1138_U483, new_P1_R1138_U484,
    new_P1_R1138_U485, new_P1_R1138_U486, new_P1_R1138_U487,
    new_P1_R1138_U488, new_P1_R1138_U489, new_P1_R1138_U490,
    new_P1_R1138_U491, new_P1_R1138_U492, new_P1_R1138_U493,
    new_P1_R1138_U494, new_P1_R1138_U495, new_P1_R1138_U496,
    new_P1_R1138_U497, new_P1_R1138_U498, new_P1_R1138_U499,
    new_P1_R1138_U500, new_P1_R1138_U501, new_P1_R1222_U4, new_P1_R1222_U5,
    new_P1_R1222_U6, new_P1_R1222_U7, new_P1_R1222_U8, new_P1_R1222_U9,
    new_P1_R1222_U10, new_P1_R1222_U11, new_P1_R1222_U12, new_P1_R1222_U13,
    new_P1_R1222_U14, new_P1_R1222_U15, new_P1_R1222_U16, new_P1_R1222_U17,
    new_P1_R1222_U18, new_P1_R1222_U19, new_P1_R1222_U20, new_P1_R1222_U21,
    new_P1_R1222_U22, new_P1_R1222_U23, new_P1_R1222_U24, new_P1_R1222_U25,
    new_P1_R1222_U26, new_P1_R1222_U27, new_P1_R1222_U28, new_P1_R1222_U29,
    new_P1_R1222_U30, new_P1_R1222_U31, new_P1_R1222_U32, new_P1_R1222_U33,
    new_P1_R1222_U34, new_P1_R1222_U35, new_P1_R1222_U36, new_P1_R1222_U37,
    new_P1_R1222_U38, new_P1_R1222_U39, new_P1_R1222_U40, new_P1_R1222_U41,
    new_P1_R1222_U42, new_P1_R1222_U43, new_P1_R1222_U44, new_P1_R1222_U45,
    new_P1_R1222_U46, new_P1_R1222_U47, new_P1_R1222_U48, new_P1_R1222_U49,
    new_P1_R1222_U50, new_P1_R1222_U51, new_P1_R1222_U52, new_P1_R1222_U53,
    new_P1_R1222_U54, new_P1_R1222_U55, new_P1_R1222_U56, new_P1_R1222_U57,
    new_P1_R1222_U58, new_P1_R1222_U59, new_P1_R1222_U60, new_P1_R1222_U61,
    new_P1_R1222_U62, new_P1_R1222_U63, new_P1_R1222_U64, new_P1_R1222_U65,
    new_P1_R1222_U66, new_P1_R1222_U67, new_P1_R1222_U68, new_P1_R1222_U69,
    new_P1_R1222_U70, new_P1_R1222_U71, new_P1_R1222_U72, new_P1_R1222_U73,
    new_P1_R1222_U74, new_P1_R1222_U75, new_P1_R1222_U76, new_P1_R1222_U77,
    new_P1_R1222_U78, new_P1_R1222_U79, new_P1_R1222_U80, new_P1_R1222_U81,
    new_P1_R1222_U82, new_P1_R1222_U83, new_P1_R1222_U84, new_P1_R1222_U85,
    new_P1_R1222_U86, new_P1_R1222_U87, new_P1_R1222_U88, new_P1_R1222_U89,
    new_P1_R1222_U90, new_P1_R1222_U91, new_P1_R1222_U92, new_P1_R1222_U93,
    new_P1_R1222_U94, new_P1_R1222_U95, new_P1_R1222_U96, new_P1_R1222_U97,
    new_P1_R1222_U98, new_P1_R1222_U99, new_P1_R1222_U100,
    new_P1_R1222_U101, new_P1_R1222_U102, new_P1_R1222_U103,
    new_P1_R1222_U104, new_P1_R1222_U105, new_P1_R1222_U106,
    new_P1_R1222_U107, new_P1_R1222_U108, new_P1_R1222_U109,
    new_P1_R1222_U110, new_P1_R1222_U111, new_P1_R1222_U112,
    new_P1_R1222_U113, new_P1_R1222_U114, new_P1_R1222_U115,
    new_P1_R1222_U116, new_P1_R1222_U117, new_P1_R1222_U118,
    new_P1_R1222_U119, new_P1_R1222_U120, new_P1_R1222_U121,
    new_P1_R1222_U122, new_P1_R1222_U123, new_P1_R1222_U124,
    new_P1_R1222_U125, new_P1_R1222_U126, new_P1_R1222_U127,
    new_P1_R1222_U128, new_P1_R1222_U129, new_P1_R1222_U130,
    new_P1_R1222_U131, new_P1_R1222_U132, new_P1_R1222_U133,
    new_P1_R1222_U134, new_P1_R1222_U135, new_P1_R1222_U136,
    new_P1_R1222_U137, new_P1_R1222_U138, new_P1_R1222_U139,
    new_P1_R1222_U140, new_P1_R1222_U141, new_P1_R1222_U142,
    new_P1_R1222_U143, new_P1_R1222_U144, new_P1_R1222_U145,
    new_P1_R1222_U146, new_P1_R1222_U147, new_P1_R1222_U148,
    new_P1_R1222_U149, new_P1_R1222_U150, new_P1_R1222_U151,
    new_P1_R1222_U152, new_P1_R1222_U153, new_P1_R1222_U154,
    new_P1_R1222_U155, new_P1_R1222_U156, new_P1_R1222_U157,
    new_P1_R1222_U158, new_P1_R1222_U159, new_P1_R1222_U160,
    new_P1_R1222_U161, new_P1_R1222_U162, new_P1_R1222_U163,
    new_P1_R1222_U164, new_P1_R1222_U165, new_P1_R1222_U166,
    new_P1_R1222_U167, new_P1_R1222_U168, new_P1_R1222_U169,
    new_P1_R1222_U170, new_P1_R1222_U171, new_P1_R1222_U172,
    new_P1_R1222_U173, new_P1_R1222_U174, new_P1_R1222_U175,
    new_P1_R1222_U176, new_P1_R1222_U177, new_P1_R1222_U178,
    new_P1_R1222_U179, new_P1_R1222_U180, new_P1_R1222_U181,
    new_P1_R1222_U182, new_P1_R1222_U183, new_P1_R1222_U184,
    new_P1_R1222_U185, new_P1_R1222_U186, new_P1_R1222_U187,
    new_P1_R1222_U188, new_P1_R1222_U189, new_P1_R1222_U190,
    new_P1_R1222_U191, new_P1_R1222_U192, new_P1_R1222_U193,
    new_P1_R1222_U194, new_P1_R1222_U195, new_P1_R1222_U196,
    new_P1_R1222_U197, new_P1_R1222_U198, new_P1_R1222_U199,
    new_P1_R1222_U200, new_P1_R1222_U201, new_P1_R1222_U202,
    new_P1_R1222_U203, new_P1_R1222_U204, new_P1_R1222_U205,
    new_P1_R1222_U206, new_P1_R1222_U207, new_P1_R1222_U208,
    new_P1_R1222_U209, new_P1_R1222_U210, new_P1_R1222_U211,
    new_P1_R1222_U212, new_P1_R1222_U213, new_P1_R1222_U214,
    new_P1_R1222_U215, new_P1_R1222_U216, new_P1_R1222_U217,
    new_P1_R1222_U218, new_P1_R1222_U219, new_P1_R1222_U220,
    new_P1_R1222_U221, new_P1_R1222_U222, new_P1_R1222_U223,
    new_P1_R1222_U224, new_P1_R1222_U225, new_P1_R1222_U226,
    new_P1_R1222_U227, new_P1_R1222_U228, new_P1_R1222_U229,
    new_P1_R1222_U230, new_P1_R1222_U231, new_P1_R1222_U232,
    new_P1_R1222_U233, new_P1_R1222_U234, new_P1_R1222_U235,
    new_P1_R1222_U236, new_P1_R1222_U237, new_P1_R1222_U238,
    new_P1_R1222_U239, new_P1_R1222_U240, new_P1_R1222_U241,
    new_P1_R1222_U242, new_P1_R1222_U243, new_P1_R1222_U244,
    new_P1_R1222_U245, new_P1_R1222_U246, new_P1_R1222_U247,
    new_P1_R1222_U248, new_P1_R1222_U249, new_P1_R1222_U250,
    new_P1_R1222_U251, new_P1_R1222_U252, new_P1_R1222_U253,
    new_P1_R1222_U254, new_P1_R1222_U255, new_P1_R1222_U256,
    new_P1_R1222_U257, new_P1_R1222_U258, new_P1_R1222_U259,
    new_P1_R1222_U260, new_P1_R1222_U261, new_P1_R1222_U262,
    new_P1_R1222_U263, new_P1_R1222_U264, new_P1_R1222_U265,
    new_P1_R1222_U266, new_P1_R1222_U267, new_P1_R1222_U268,
    new_P1_R1222_U269, new_P1_R1222_U270, new_P1_R1222_U271,
    new_P1_R1222_U272, new_P1_R1222_U273, new_P1_R1222_U274,
    new_P1_R1222_U275, new_P1_R1222_U276, new_P1_R1222_U277,
    new_P1_R1222_U278, new_P1_R1222_U279, new_P1_R1222_U280,
    new_P1_R1222_U281, new_P1_R1222_U282, new_P1_R1222_U283,
    new_P1_R1222_U284, new_P1_R1222_U285, new_P1_R1222_U286,
    new_P1_R1222_U287, new_P1_R1222_U288, new_P1_R1222_U289,
    new_P1_R1222_U290, new_P1_R1222_U291, new_P1_R1222_U292,
    new_P1_R1222_U293, new_P1_R1222_U294, new_P1_R1222_U295,
    new_P1_R1222_U296, new_P1_R1222_U297, new_P1_R1222_U298,
    new_P1_R1222_U299, new_P1_R1222_U300, new_P1_R1222_U301,
    new_P1_R1222_U302, new_P1_R1222_U303, new_P1_R1222_U304,
    new_P1_R1222_U305, new_P1_R1222_U306, new_P1_R1222_U307,
    new_P1_R1222_U308, new_P1_R1222_U309, new_P1_R1222_U310,
    new_P1_R1222_U311, new_P1_R1222_U312, new_P1_R1222_U313,
    new_P1_R1222_U314, new_P1_R1222_U315, new_P1_R1222_U316,
    new_P1_R1222_U317, new_P1_R1222_U318, new_P1_R1222_U319,
    new_P1_R1222_U320, new_P1_R1222_U321, new_P1_R1222_U322,
    new_P1_R1222_U323, new_P1_R1222_U324, new_P1_R1222_U325,
    new_P1_R1222_U326, new_P1_R1222_U327, new_P1_R1222_U328,
    new_P1_R1222_U329, new_P1_R1222_U330, new_P1_R1222_U331,
    new_P1_R1222_U332, new_P1_R1222_U333, new_P1_R1222_U334,
    new_P1_R1222_U335, new_P1_R1222_U336, new_P1_R1222_U337,
    new_P1_R1222_U338, new_P1_R1222_U339, new_P1_R1222_U340,
    new_P1_R1222_U341, new_P1_R1222_U342, new_P1_R1222_U343,
    new_P1_R1222_U344, new_P1_R1222_U345, new_P1_R1222_U346,
    new_P1_R1222_U347, new_P1_R1222_U348, new_P1_R1222_U349,
    new_P1_R1222_U350, new_P1_R1222_U351, new_P1_R1222_U352,
    new_P1_R1222_U353, new_P1_R1222_U354, new_P1_R1222_U355,
    new_P1_R1222_U356, new_P1_R1222_U357, new_P1_R1222_U358,
    new_P1_R1222_U359, new_P1_R1222_U360, new_P1_R1222_U361,
    new_P1_R1222_U362, new_P1_R1222_U363, new_P1_R1222_U364,
    new_P1_R1222_U365, new_P1_R1222_U366, new_P1_R1222_U367,
    new_P1_R1222_U368, new_P1_R1222_U369, new_P1_R1222_U370,
    new_P1_R1222_U371, new_P1_R1222_U372, new_P1_R1222_U373,
    new_P1_R1222_U374, new_P1_R1222_U375, new_P1_R1222_U376,
    new_P1_R1222_U377, new_P1_R1222_U378, new_P1_R1222_U379,
    new_P1_R1222_U380, new_P1_R1222_U381, new_P1_R1222_U382,
    new_P1_R1222_U383, new_P1_R1222_U384, new_P1_R1222_U385,
    new_P1_R1222_U386, new_P1_R1222_U387, new_P1_R1222_U388,
    new_P1_R1222_U389, new_P1_R1222_U390, new_P1_R1222_U391,
    new_P1_R1222_U392, new_P1_R1222_U393, new_P1_R1222_U394,
    new_P1_R1222_U395, new_P1_R1222_U396, new_P1_R1222_U397,
    new_P1_R1222_U398, new_P1_R1222_U399, new_P1_R1222_U400,
    new_P1_R1222_U401, new_P1_R1222_U402, new_P1_R1222_U403,
    new_P1_R1222_U404, new_P1_R1222_U405, new_P1_R1222_U406,
    new_P1_R1222_U407, new_P1_R1222_U408, new_P1_R1222_U409,
    new_P1_R1222_U410, new_P1_R1222_U411, new_P1_R1222_U412,
    new_P1_R1222_U413, new_P1_R1222_U414, new_P1_R1222_U415,
    new_P1_R1222_U416, new_P1_R1222_U417, new_P1_R1222_U418,
    new_P1_R1222_U419, new_P1_R1222_U420, new_P1_R1222_U421,
    new_P1_R1222_U422, new_P1_R1222_U423, new_P1_R1222_U424,
    new_P1_R1222_U425, new_P1_R1222_U426, new_P1_R1222_U427,
    new_P1_R1222_U428, new_P1_R1222_U429, new_P1_R1222_U430,
    new_P1_R1222_U431, new_P1_R1222_U432, new_P1_R1222_U433,
    new_P1_R1222_U434, new_P1_R1222_U435, new_P1_R1222_U436,
    new_P1_R1222_U437, new_P1_R1222_U438, new_P1_R1222_U439,
    new_P1_R1222_U440, new_P1_R1222_U441, new_P1_R1222_U442,
    new_P1_R1222_U443, new_P1_R1222_U444, new_P1_R1222_U445,
    new_P1_R1222_U446, new_P1_R1222_U447, new_P1_R1222_U448,
    new_P1_R1222_U449, new_P1_R1222_U450, new_P1_R1222_U451,
    new_P1_R1222_U452, new_P1_R1222_U453, new_P1_R1222_U454,
    new_P1_R1222_U455, new_P1_R1222_U456, new_P1_R1222_U457,
    new_P1_R1222_U458, new_P1_R1222_U459, new_P1_R1222_U460,
    new_P1_R1222_U461, new_P1_R1222_U462, new_P1_R1222_U463,
    new_P1_R1222_U464, new_P1_R1222_U465, new_P1_R1222_U466,
    new_P1_R1222_U467, new_P1_R1222_U468, new_P1_R1222_U469,
    new_P1_R1222_U470, new_P1_R1222_U471, new_P1_R1222_U472,
    new_P1_R1222_U473, new_P1_R1222_U474, new_P1_R1222_U475,
    new_P1_R1222_U476, new_P1_R1222_U477, new_P1_R1222_U478,
    new_P1_R1222_U479, new_P1_R1222_U480, new_P1_R1222_U481,
    new_P1_R1222_U482, new_P1_R1222_U483, new_P1_R1222_U484,
    new_P1_R1222_U485, new_P1_R1222_U486, new_P1_R1222_U487,
    new_P1_R1222_U488, new_P1_R1222_U489, new_P1_R1222_U490,
    new_P1_R1222_U491, new_P1_R1222_U492, new_P1_R1222_U493,
    new_P1_R1222_U494, new_P1_R1222_U495, new_P1_R1222_U496,
    new_P1_R1222_U497, new_P1_R1222_U498, new_P1_R1222_U499,
    new_P1_R1222_U500, new_P1_R1222_U501, new_P2_ADD_1119_U4,
    new_P2_ADD_1119_U5, new_P2_ADD_1119_U6, new_P2_ADD_1119_U7,
    new_P2_ADD_1119_U8, new_P2_ADD_1119_U9, new_P2_ADD_1119_U10,
    new_P2_ADD_1119_U11, new_P2_ADD_1119_U12, new_P2_ADD_1119_U13,
    new_P2_ADD_1119_U14, new_P2_ADD_1119_U15, new_P2_ADD_1119_U16,
    new_P2_ADD_1119_U17, new_P2_ADD_1119_U18, new_P2_ADD_1119_U19,
    new_P2_ADD_1119_U20, new_P2_ADD_1119_U21, new_P2_ADD_1119_U22,
    new_P2_ADD_1119_U23, new_P2_ADD_1119_U24, new_P2_ADD_1119_U25,
    new_P2_ADD_1119_U26, new_P2_ADD_1119_U27, new_P2_ADD_1119_U28,
    new_P2_ADD_1119_U29, new_P2_ADD_1119_U30, new_P2_ADD_1119_U31,
    new_P2_ADD_1119_U32, new_P2_ADD_1119_U33, new_P2_ADD_1119_U34,
    new_P2_ADD_1119_U35, new_P2_ADD_1119_U36, new_P2_ADD_1119_U37,
    new_P2_ADD_1119_U38, new_P2_ADD_1119_U39, new_P2_ADD_1119_U40,
    new_P2_ADD_1119_U41, new_P2_ADD_1119_U42, new_P2_ADD_1119_U43,
    new_P2_ADD_1119_U44, new_P2_ADD_1119_U45, new_P2_ADD_1119_U46,
    new_P2_ADD_1119_U47, new_P2_ADD_1119_U48, new_P2_ADD_1119_U49,
    new_P2_ADD_1119_U50, new_P2_ADD_1119_U51, new_P2_ADD_1119_U52,
    new_P2_ADD_1119_U53, new_P2_ADD_1119_U54, new_P2_ADD_1119_U55,
    new_P2_ADD_1119_U56, new_P2_ADD_1119_U57, new_P2_ADD_1119_U58,
    new_P2_ADD_1119_U59, new_P2_ADD_1119_U60, new_P2_ADD_1119_U61,
    new_P2_ADD_1119_U62, new_P2_ADD_1119_U63, new_P2_ADD_1119_U64,
    new_P2_ADD_1119_U65, new_P2_ADD_1119_U66, new_P2_ADD_1119_U67,
    new_P2_ADD_1119_U68, new_P2_ADD_1119_U69, new_P2_ADD_1119_U70,
    new_P2_ADD_1119_U71, new_P2_ADD_1119_U72, new_P2_ADD_1119_U73,
    new_P2_ADD_1119_U74, new_P2_ADD_1119_U75, new_P2_ADD_1119_U76,
    new_P2_ADD_1119_U77, new_P2_ADD_1119_U78, new_P2_ADD_1119_U79,
    new_P2_ADD_1119_U80, new_P2_ADD_1119_U81, new_P2_ADD_1119_U82,
    new_P2_ADD_1119_U83, new_P2_ADD_1119_U84, new_P2_ADD_1119_U85,
    new_P2_ADD_1119_U86, new_P2_ADD_1119_U87, new_P2_ADD_1119_U88,
    new_P2_ADD_1119_U89, new_P2_ADD_1119_U90, new_P2_ADD_1119_U91,
    new_P2_ADD_1119_U92, new_P2_ADD_1119_U93, new_P2_ADD_1119_U94,
    new_P2_ADD_1119_U95, new_P2_ADD_1119_U96, new_P2_ADD_1119_U97,
    new_P2_ADD_1119_U98, new_P2_ADD_1119_U99, new_P2_ADD_1119_U100,
    new_P2_ADD_1119_U101, new_P2_ADD_1119_U102, new_P2_ADD_1119_U103,
    new_P2_ADD_1119_U104, new_P2_ADD_1119_U105, new_P2_ADD_1119_U106,
    new_P2_ADD_1119_U107, new_P2_ADD_1119_U108, new_P2_ADD_1119_U109,
    new_P2_ADD_1119_U110, new_P2_ADD_1119_U111, new_P2_ADD_1119_U112,
    new_P2_ADD_1119_U113, new_P2_ADD_1119_U114, new_P2_ADD_1119_U115,
    new_P2_ADD_1119_U116, new_P2_ADD_1119_U117, new_P2_ADD_1119_U118,
    new_P2_ADD_1119_U119, new_P2_ADD_1119_U120, new_P2_ADD_1119_U121,
    new_P2_ADD_1119_U122, new_P2_ADD_1119_U123, new_P2_ADD_1119_U124,
    new_P2_ADD_1119_U125, new_P2_ADD_1119_U126, new_P2_ADD_1119_U127,
    new_P2_ADD_1119_U128, new_P2_ADD_1119_U129, new_P2_ADD_1119_U130,
    new_P2_ADD_1119_U131, new_P2_ADD_1119_U132, new_P2_ADD_1119_U133,
    new_P2_ADD_1119_U134, new_P2_ADD_1119_U135, new_P2_ADD_1119_U136,
    new_P2_ADD_1119_U137, new_P2_ADD_1119_U138, new_P2_ADD_1119_U139,
    new_P2_ADD_1119_U140, new_P2_ADD_1119_U141, new_P2_ADD_1119_U142,
    new_P2_ADD_1119_U143, new_P2_ADD_1119_U144, new_P2_ADD_1119_U145,
    new_P2_ADD_1119_U146, new_P2_ADD_1119_U147, new_P2_ADD_1119_U148,
    new_P2_ADD_1119_U149, new_P2_ADD_1119_U150, new_P2_ADD_1119_U151,
    new_P2_ADD_1119_U152, new_P2_ADD_1119_U153, new_P2_ADD_1119_U154,
    new_P2_ADD_1119_U155, new_P2_ADD_1119_U156, new_P2_ADD_1119_U157,
    new_P2_SUB_1108_U6, new_P2_SUB_1108_U7, new_P2_SUB_1108_U8,
    new_P2_SUB_1108_U9, new_P2_SUB_1108_U10, new_P2_SUB_1108_U11,
    new_P2_SUB_1108_U12, new_P2_SUB_1108_U13, new_P2_SUB_1108_U14,
    new_P2_SUB_1108_U15, new_P2_SUB_1108_U16, new_P2_SUB_1108_U17,
    new_P2_SUB_1108_U18, new_P2_SUB_1108_U19, new_P2_SUB_1108_U20,
    new_P2_SUB_1108_U21, new_P2_SUB_1108_U22, new_P2_SUB_1108_U23,
    new_P2_SUB_1108_U24, new_P2_SUB_1108_U25, new_P2_SUB_1108_U26,
    new_P2_SUB_1108_U27, new_P2_SUB_1108_U28, new_P2_SUB_1108_U29,
    new_P2_SUB_1108_U30, new_P2_SUB_1108_U31, new_P2_SUB_1108_U32,
    new_P2_SUB_1108_U33, new_P2_SUB_1108_U34, new_P2_SUB_1108_U35,
    new_P2_SUB_1108_U36, new_P2_SUB_1108_U37, new_P2_SUB_1108_U38,
    new_P2_SUB_1108_U39, new_P2_SUB_1108_U40, new_P2_SUB_1108_U41,
    new_P2_SUB_1108_U42, new_P2_SUB_1108_U43, new_P2_SUB_1108_U44,
    new_P2_SUB_1108_U45, new_P2_SUB_1108_U46, new_P2_SUB_1108_U47,
    new_P2_SUB_1108_U48, new_P2_SUB_1108_U49, new_P2_SUB_1108_U50,
    new_P2_SUB_1108_U51, new_P2_SUB_1108_U52, new_P2_SUB_1108_U53,
    new_P2_SUB_1108_U54, new_P2_SUB_1108_U55, new_P2_SUB_1108_U56,
    new_P2_SUB_1108_U57, new_P2_SUB_1108_U58, new_P2_SUB_1108_U59,
    new_P2_SUB_1108_U60, new_P2_SUB_1108_U61, new_P2_SUB_1108_U62,
    new_P2_SUB_1108_U63, new_P2_SUB_1108_U64, new_P2_SUB_1108_U65,
    new_P2_SUB_1108_U66, new_P2_SUB_1108_U67, new_P2_SUB_1108_U68,
    new_P2_SUB_1108_U69, new_P2_SUB_1108_U70, new_P2_SUB_1108_U71,
    new_P2_SUB_1108_U72, new_P2_SUB_1108_U73, new_P2_SUB_1108_U74,
    new_P2_SUB_1108_U75, new_P2_SUB_1108_U76, new_P2_SUB_1108_U77,
    new_P2_SUB_1108_U78, new_P2_SUB_1108_U79, new_P2_SUB_1108_U80,
    new_P2_SUB_1108_U81, new_P2_SUB_1108_U82, new_P2_SUB_1108_U83,
    new_P2_SUB_1108_U84, new_P2_SUB_1108_U85, new_P2_SUB_1108_U86,
    new_P2_SUB_1108_U87, new_P2_SUB_1108_U88, new_P2_SUB_1108_U89,
    new_P2_SUB_1108_U90, new_P2_SUB_1108_U91, new_P2_SUB_1108_U92,
    new_P2_SUB_1108_U93, new_P2_SUB_1108_U94, new_P2_SUB_1108_U95,
    new_P2_SUB_1108_U96, new_P2_SUB_1108_U97, new_P2_SUB_1108_U98,
    new_P2_SUB_1108_U99, new_P2_SUB_1108_U100, new_P2_SUB_1108_U101,
    new_P2_SUB_1108_U102, new_P2_SUB_1108_U103, new_P2_SUB_1108_U104,
    new_P2_SUB_1108_U105, new_P2_SUB_1108_U106, new_P2_SUB_1108_U107,
    new_P2_SUB_1108_U108, new_P2_SUB_1108_U109, new_P2_SUB_1108_U110,
    new_P2_SUB_1108_U111, new_P2_SUB_1108_U112, new_P2_SUB_1108_U113,
    new_P2_SUB_1108_U114, new_P2_SUB_1108_U115, new_P2_SUB_1108_U116,
    new_P2_SUB_1108_U117, new_P2_SUB_1108_U118, new_P2_SUB_1108_U119,
    new_P2_SUB_1108_U120, new_P2_SUB_1108_U121, new_P2_SUB_1108_U122,
    new_P2_SUB_1108_U123, new_P2_SUB_1108_U124, new_P2_SUB_1108_U125,
    new_P2_SUB_1108_U126, new_P2_SUB_1108_U127, new_P2_SUB_1108_U128,
    new_P2_SUB_1108_U129, new_P2_SUB_1108_U130, new_P2_SUB_1108_U131,
    new_P2_SUB_1108_U132, new_P2_SUB_1108_U133, new_P2_SUB_1108_U134,
    new_P2_SUB_1108_U135, new_P2_SUB_1108_U136, new_P2_SUB_1108_U137,
    new_P2_SUB_1108_U138, new_P2_SUB_1108_U139, new_P2_SUB_1108_U140,
    new_P2_SUB_1108_U141, new_P2_SUB_1108_U142, new_P2_SUB_1108_U143,
    new_P2_SUB_1108_U144, new_P2_SUB_1108_U145, new_P2_SUB_1108_U146,
    new_P2_SUB_1108_U147, new_P2_SUB_1108_U148, new_P2_SUB_1108_U149,
    new_P2_SUB_1108_U150, new_P2_SUB_1108_U151, new_P2_SUB_1108_U152,
    new_P2_SUB_1108_U153, new_P2_SUB_1108_U154, new_P2_SUB_1108_U155,
    new_P2_SUB_1108_U156, new_P2_SUB_1108_U157, new_P2_SUB_1108_U158,
    new_P2_SUB_1108_U159, new_P2_SUB_1108_U160, new_P2_SUB_1108_U161,
    new_P2_SUB_1108_U162, new_P2_SUB_1108_U163, new_P2_SUB_1108_U164,
    new_P2_SUB_1108_U165, new_P2_SUB_1108_U166, new_P2_SUB_1108_U167,
    new_P2_SUB_1108_U168, new_P2_SUB_1108_U169, new_P2_SUB_1108_U170,
    new_P2_SUB_1108_U171, new_P2_SUB_1108_U172, new_P2_SUB_1108_U173,
    new_P2_SUB_1108_U174, new_P2_SUB_1108_U175, new_P2_SUB_1108_U176,
    new_P2_SUB_1108_U177, new_P2_SUB_1108_U178, new_P2_SUB_1108_U179,
    new_P2_SUB_1108_U180, new_P2_SUB_1108_U181, new_P2_SUB_1108_U182,
    new_P2_SUB_1108_U183, new_P2_SUB_1108_U184, new_P2_SUB_1108_U185,
    new_P2_SUB_1108_U186, new_P2_SUB_1108_U187, new_P2_SUB_1108_U188,
    new_P2_SUB_1108_U189, new_P2_SUB_1108_U190, new_P2_SUB_1108_U191,
    new_P2_SUB_1108_U192, new_P2_SUB_1108_U193, new_P2_SUB_1108_U194,
    new_P2_SUB_1108_U195, new_P2_SUB_1108_U196, new_P2_SUB_1108_U197,
    new_P2_SUB_1108_U198, new_P2_SUB_1108_U199, new_P2_SUB_1108_U200,
    new_P2_SUB_1108_U201, new_P2_SUB_1108_U202, new_P2_R1299_U6,
    new_P2_R1299_U7, new_P2_R1312_U6, new_P2_R1312_U7, new_P2_R1312_U8,
    new_P2_R1312_U9, new_P2_R1312_U10, new_P2_R1312_U11, new_P2_R1312_U12,
    new_P2_R1312_U13, new_P2_R1312_U14, new_P2_R1312_U15, new_P2_R1312_U16,
    new_P2_R1312_U17, new_P2_R1312_U18, new_P2_R1312_U19, new_P2_R1312_U20,
    new_P2_R1312_U21, new_P2_R1312_U22, new_P2_R1312_U23, new_P2_R1312_U24,
    new_P2_R1312_U25, new_P2_R1312_U26, new_P2_R1312_U27, new_P2_R1312_U28,
    new_P2_R1312_U29, new_P2_R1312_U30, new_P2_R1312_U31, new_P2_R1312_U32,
    new_P2_R1312_U33, new_P2_R1312_U34, new_P2_R1312_U35, new_P2_R1312_U36,
    new_P2_R1312_U37, new_P2_R1312_U38, new_P2_R1312_U39, new_P2_R1312_U40,
    new_P2_R1312_U41, new_P2_R1312_U42, new_P2_R1312_U43, new_P2_R1312_U44,
    new_P2_R1312_U45, new_P2_R1312_U46, new_P2_R1312_U47, new_P2_R1312_U48,
    new_P2_R1312_U49, new_P2_R1312_U50, new_P2_R1312_U51, new_P2_R1312_U52,
    new_P2_R1312_U53, new_P2_R1312_U54, new_P2_R1312_U55, new_P2_R1312_U56,
    new_P2_R1312_U57, new_P2_R1312_U58, new_P2_R1312_U59, new_P2_R1312_U60,
    new_P2_R1312_U61, new_P2_R1312_U62, new_P2_R1312_U63, new_P2_R1312_U64,
    new_P2_R1312_U65, new_P2_R1312_U66, new_P2_R1312_U67, new_P2_R1312_U68,
    new_P2_R1312_U69, new_P2_R1312_U70, new_P2_R1312_U71, new_P2_R1312_U72,
    new_P2_R1312_U73, new_P2_R1312_U74, new_P2_R1312_U75, new_P2_R1312_U76,
    new_P2_R1312_U77, new_P2_R1312_U78, new_P2_R1312_U79, new_P2_R1312_U80,
    new_P2_R1312_U81, new_P2_R1312_U82, new_P2_R1312_U83, new_P2_R1312_U84,
    new_P2_R1312_U85, new_P2_R1312_U86, new_P2_R1312_U87, new_P2_R1312_U88,
    new_P2_R1312_U89, new_P2_R1312_U90, new_P2_R1312_U91, new_P2_R1312_U92,
    new_P2_R1312_U93, new_P2_R1312_U94, new_P2_R1312_U95, new_P2_R1312_U96,
    new_P2_R1312_U97, new_P2_R1312_U98, new_P2_R1312_U99,
    new_P2_R1312_U100, new_P2_R1312_U101, new_P2_R1312_U102,
    new_P2_R1312_U103, new_P2_R1312_U104, new_P2_R1312_U105,
    new_P2_R1312_U106, new_P2_R1312_U107, new_P2_R1312_U108,
    new_P2_R1312_U109, new_P2_R1312_U110, new_P2_R1312_U111,
    new_P2_R1312_U112, new_P2_R1312_U113, new_P2_R1312_U114,
    new_P2_R1312_U115, new_P2_R1312_U116, new_P2_R1312_U117,
    new_P2_R1312_U118, new_P2_R1312_U119, new_P2_R1312_U120,
    new_P2_R1312_U121, new_P2_R1312_U122, new_P2_R1312_U123,
    new_P2_R1312_U124, new_P2_R1312_U125, new_P2_R1312_U126,
    new_P2_R1312_U127, new_P2_R1312_U128, new_P2_R1312_U129,
    new_P2_R1312_U130, new_P2_R1312_U131, new_P2_R1312_U132,
    new_P2_R1312_U133, new_P2_R1312_U134, new_P2_R1312_U135,
    new_P2_R1312_U136, new_P2_R1312_U137, new_P2_R1312_U138,
    new_P2_R1312_U139, new_P2_R1312_U140, new_P2_R1312_U141,
    new_P2_R1312_U142, new_P2_R1312_U143, new_P2_R1312_U144,
    new_P2_R1312_U145, new_P2_R1312_U146, new_P2_R1312_U147,
    new_P2_R1312_U148, new_P2_R1312_U149, new_P2_R1312_U150,
    new_P2_R1312_U151, new_P2_R1312_U152, new_P2_R1312_U153,
    new_P2_R1312_U154, new_P2_R1312_U155, new_P2_R1312_U156,
    new_P2_R1312_U157, new_P2_R1312_U158, new_P2_R1312_U159,
    new_P2_R1312_U160, new_P2_R1312_U161, new_P2_R1312_U162,
    new_P2_R1312_U163, new_P2_R1312_U164, new_P2_R1312_U165,
    new_P2_R1312_U166, new_P2_R1312_U167, new_P2_R1312_U168,
    new_P2_R1312_U169, new_P2_R1312_U170, new_P2_R1312_U171,
    new_P2_R1312_U172, new_P2_R1312_U173, new_P2_R1312_U174,
    new_P2_R1312_U175, new_P2_R1312_U176, new_P2_R1312_U177,
    new_P2_R1312_U178, new_P2_R1312_U179, new_P2_R1312_U180,
    new_P2_R1312_U181, new_P2_R1312_U182, new_P2_R1312_U183,
    new_P2_R1312_U184, new_P2_R1312_U185, new_P2_R1312_U186,
    new_P2_R1312_U187, new_P2_R1312_U188, new_P2_R1312_U189,
    new_P2_R1312_U190, new_P2_R1312_U191, new_P2_R1312_U192,
    new_P2_R1312_U193, new_P2_R1312_U194, new_P2_R1312_U195,
    new_P2_R1312_U196, new_P2_R1312_U197, new_P2_R1312_U198,
    new_P2_R1312_U199, new_P2_R1312_U200, new_P2_R1312_U201,
    new_P2_R1312_U202, new_P2_R1312_U203, new_P2_R1312_U204,
    new_P2_R1312_U205, new_P2_R1312_U206, new_P2_R1312_U207,
    new_P2_R1312_U208, new_P2_R1312_U209, new_P2_R1312_U210,
    new_P2_R1312_U211, new_P2_R1312_U212, new_P2_R1312_U213,
    new_P2_R1312_U214, new_P2_R1312_U215, new_P2_R1312_U216,
    new_P2_R1312_U217, new_P2_R1312_U218, new_P2_R1312_U219,
    new_P2_R1312_U220, new_P2_R1312_U221, new_P2_R1312_U222,
    new_P2_R1312_U223, new_P2_R1312_U224, new_P2_R1312_U225,
    new_P2_R1312_U226, new_P2_R1312_U227, new_P2_R1335_U6, new_P2_R1335_U7,
    new_P2_R1335_U8, new_P2_R1335_U9, new_P2_R1335_U10, new_P2_R1209_U4,
    new_P2_R1209_U5, new_P2_R1209_U6, new_P2_R1209_U7, new_P2_R1209_U8,
    new_P2_R1209_U9, new_P2_R1209_U10, new_P2_R1209_U11, new_P2_R1209_U12,
    new_P2_R1209_U13, new_P2_R1209_U14, new_P2_R1209_U15, new_P2_R1209_U16,
    new_P2_R1209_U17, new_P2_R1209_U18, new_P2_R1209_U19, new_P2_R1209_U20,
    new_P2_R1209_U21, new_P2_R1209_U22, new_P2_R1209_U23, new_P2_R1209_U24,
    new_P2_R1209_U25, new_P2_R1209_U26, new_P2_R1209_U27, new_P2_R1209_U28,
    new_P2_R1209_U29, new_P2_R1209_U30, new_P2_R1209_U31, new_P2_R1209_U32,
    new_P2_R1209_U33, new_P2_R1209_U34, new_P2_R1209_U35, new_P2_R1209_U36,
    new_P2_R1209_U37, new_P2_R1209_U38, new_P2_R1209_U39, new_P2_R1209_U40,
    new_P2_R1209_U41, new_P2_R1209_U42, new_P2_R1209_U43, new_P2_R1209_U44,
    new_P2_R1209_U45, new_P2_R1209_U46, new_P2_R1209_U47, new_P2_R1209_U48,
    new_P2_R1209_U49, new_P2_R1209_U50, new_P2_R1209_U51, new_P2_R1209_U52,
    new_P2_R1209_U53, new_P2_R1209_U54, new_P2_R1209_U55, new_P2_R1209_U56,
    new_P2_R1209_U57, new_P2_R1209_U58, new_P2_R1209_U59, new_P2_R1209_U60,
    new_P2_R1209_U61, new_P2_R1209_U62, new_P2_R1209_U63, new_P2_R1209_U64,
    new_P2_R1209_U65, new_P2_R1209_U66, new_P2_R1209_U67, new_P2_R1209_U68,
    new_P2_R1209_U69, new_P2_R1209_U70, new_P2_R1209_U71, new_P2_R1209_U72,
    new_P2_R1209_U73, new_P2_R1209_U74, new_P2_R1209_U75, new_P2_R1209_U76,
    new_P2_R1209_U77, new_P2_R1209_U78, new_P2_R1209_U79, new_P2_R1209_U80,
    new_P2_R1209_U81, new_P2_R1209_U82, new_P2_R1209_U83, new_P2_R1209_U84,
    new_P2_R1209_U85, new_P2_R1209_U86, new_P2_R1209_U87, new_P2_R1209_U88,
    new_P2_R1209_U89, new_P2_R1209_U90, new_P2_R1209_U91, new_P2_R1209_U92,
    new_P2_R1209_U93, new_P2_R1209_U94, new_P2_R1209_U95, new_P2_R1209_U96,
    new_P2_R1209_U97, new_P2_R1209_U98, new_P2_R1209_U99,
    new_P2_R1209_U100, new_P2_R1209_U101, new_P2_R1209_U102,
    new_P2_R1209_U103, new_P2_R1209_U104, new_P2_R1209_U105,
    new_P2_R1209_U106, new_P2_R1209_U107, new_P2_R1209_U108,
    new_P2_R1209_U109, new_P2_R1209_U110, new_P2_R1209_U111,
    new_P2_R1209_U112, new_P2_R1209_U113, new_P2_R1209_U114,
    new_P2_R1209_U115, new_P2_R1209_U116, new_P2_R1209_U117,
    new_P2_R1209_U118, new_P2_R1209_U119, new_P2_R1209_U120,
    new_P2_R1209_U121, new_P2_R1209_U122, new_P2_R1209_U123,
    new_P2_R1209_U124, new_P2_R1209_U125, new_P2_R1209_U126,
    new_P2_R1209_U127, new_P2_R1209_U128, new_P2_R1209_U129,
    new_P2_R1209_U130, new_P2_R1209_U131, new_P2_R1209_U132,
    new_P2_R1209_U133, new_P2_R1209_U134, new_P2_R1209_U135,
    new_P2_R1209_U136, new_P2_R1209_U137, new_P2_R1209_U138,
    new_P2_R1209_U139, new_P2_R1209_U140, new_P2_R1209_U141,
    new_P2_R1209_U142, new_P2_R1209_U143, new_P2_R1209_U144,
    new_P2_R1209_U145, new_P2_R1209_U146, new_P2_R1209_U147,
    new_P2_R1209_U148, new_P2_R1209_U149, new_P2_R1209_U150,
    new_P2_R1209_U151, new_P2_R1209_U152, new_P2_R1209_U153,
    new_P2_R1209_U154, new_P2_R1209_U155, new_P2_R1209_U156,
    new_P2_R1209_U157, new_P2_R1209_U158, new_P2_R1209_U159,
    new_P2_R1209_U160, new_P2_R1209_U161, new_P2_R1209_U162,
    new_P2_R1209_U163, new_P2_R1209_U164, new_P2_R1209_U165,
    new_P2_R1209_U166, new_P2_R1209_U167, new_P2_R1209_U168,
    new_P2_R1209_U169, new_P2_R1209_U170, new_P2_R1209_U171,
    new_P2_R1209_U172, new_P2_R1209_U173, new_P2_R1209_U174,
    new_P2_R1209_U175, new_P2_R1209_U176, new_P2_R1209_U177,
    new_P2_R1209_U178, new_P2_R1209_U179, new_P2_R1209_U180,
    new_P2_R1209_U181, new_P2_R1209_U182, new_P2_R1209_U183,
    new_P2_R1209_U184, new_P2_R1209_U185, new_P2_R1209_U186,
    new_P2_R1209_U187, new_P2_R1209_U188, new_P2_R1209_U189,
    new_P2_R1209_U190, new_P2_R1209_U191, new_P2_R1209_U192,
    new_P2_R1209_U193, new_P2_R1209_U194, new_P2_R1209_U195,
    new_P2_R1209_U196, new_P2_R1209_U197, new_P2_R1209_U198,
    new_P2_R1209_U199, new_P2_R1209_U200, new_P2_R1209_U201,
    new_P2_R1209_U202, new_P2_R1209_U203, new_P2_R1209_U204,
    new_P2_R1209_U205, new_P2_R1209_U206, new_P2_R1209_U207,
    new_P2_R1209_U208, new_P2_R1209_U209, new_P2_R1209_U210,
    new_P2_R1209_U211, new_P2_R1209_U212, new_P2_R1209_U213,
    new_P2_R1209_U214, new_P2_R1209_U215, new_P2_R1209_U216,
    new_P2_R1209_U217, new_P2_R1209_U218, new_P2_R1209_U219,
    new_P2_R1209_U220, new_P2_R1209_U221, new_P2_R1209_U222,
    new_P2_R1209_U223, new_P2_R1209_U224, new_P2_R1209_U225,
    new_P2_R1209_U226, new_P2_R1209_U227, new_P2_R1209_U228,
    new_P2_R1209_U229, new_P2_R1209_U230, new_P2_R1209_U231,
    new_P2_R1209_U232, new_P2_R1209_U233, new_P2_R1209_U234,
    new_P2_R1209_U235, new_P2_R1209_U236, new_P2_R1209_U237,
    new_P2_R1209_U238, new_P2_R1209_U239, new_P2_R1209_U240,
    new_P2_R1209_U241, new_P2_R1209_U242, new_P2_R1209_U243,
    new_P2_R1209_U244, new_P2_R1209_U245, new_P2_R1209_U246,
    new_P2_R1209_U247, new_P2_R1209_U248, new_P2_R1209_U249,
    new_P2_R1209_U250, new_P2_R1209_U251, new_P2_R1209_U252,
    new_P2_R1209_U253, new_P2_R1209_U254, new_P2_R1209_U255,
    new_P2_R1209_U256, new_P2_R1209_U257, new_P2_R1209_U258,
    new_P2_R1209_U259, new_P2_R1209_U260, new_P2_R1209_U261,
    new_P2_R1209_U262, new_P2_R1209_U263, new_P2_R1209_U264,
    new_P2_R1209_U265, new_P2_R1209_U266, new_P2_R1209_U267,
    new_P2_R1209_U268, new_P2_R1209_U269, new_P2_R1209_U270,
    new_P2_R1209_U271, new_P2_R1209_U272, new_P2_R1209_U273,
    new_P2_R1209_U274, new_P2_R1209_U275, new_P2_R1209_U276,
    new_P2_R1209_U277, new_P2_R1209_U278, new_P2_R1209_U279,
    new_P2_R1209_U280, new_P2_R1209_U281, new_P2_R1209_U282,
    new_P2_R1209_U283, new_P2_R1209_U284, new_P2_R1209_U285,
    new_P2_R1209_U286, new_P2_R1209_U287, new_P2_R1209_U288,
    new_P2_R1209_U289, new_P2_R1209_U290, new_P2_R1209_U291,
    new_P2_R1209_U292, new_P2_R1209_U293, new_P2_R1209_U294,
    new_P2_R1209_U295, new_P2_R1209_U296, new_P2_R1209_U297,
    new_P2_R1209_U298, new_P2_R1209_U299, new_P2_R1209_U300,
    new_P2_R1209_U301, new_P2_R1209_U302, new_P2_R1209_U303,
    new_P2_R1209_U304, new_P2_R1209_U305, new_P2_R1209_U306,
    new_P2_R1209_U307, new_P2_R1209_U308, new_P2_R1170_U4, new_P2_R1170_U5,
    new_P2_R1170_U6, new_P2_R1170_U7, new_P2_R1170_U8, new_P2_R1170_U9,
    new_P2_R1170_U10, new_P2_R1170_U11, new_P2_R1170_U12, new_P2_R1170_U13,
    new_P2_R1170_U14, new_P2_R1170_U15, new_P2_R1170_U16, new_P2_R1170_U17,
    new_P2_R1170_U18, new_P2_R1170_U19, new_P2_R1170_U20, new_P2_R1170_U21,
    new_P2_R1170_U22, new_P2_R1170_U23, new_P2_R1170_U24, new_P2_R1170_U25,
    new_P2_R1170_U26, new_P2_R1170_U27, new_P2_R1170_U28, new_P2_R1170_U29,
    new_P2_R1170_U30, new_P2_R1170_U31, new_P2_R1170_U32, new_P2_R1170_U33,
    new_P2_R1170_U34, new_P2_R1170_U35, new_P2_R1170_U36, new_P2_R1170_U37,
    new_P2_R1170_U38, new_P2_R1170_U39, new_P2_R1170_U40, new_P2_R1170_U41,
    new_P2_R1170_U42, new_P2_R1170_U43, new_P2_R1170_U44, new_P2_R1170_U45,
    new_P2_R1170_U46, new_P2_R1170_U47, new_P2_R1170_U48, new_P2_R1170_U49,
    new_P2_R1170_U50, new_P2_R1170_U51, new_P2_R1170_U52, new_P2_R1170_U53,
    new_P2_R1170_U54, new_P2_R1170_U55, new_P2_R1170_U56, new_P2_R1170_U57,
    new_P2_R1170_U58, new_P2_R1170_U59, new_P2_R1170_U60, new_P2_R1170_U61,
    new_P2_R1170_U62, new_P2_R1170_U63, new_P2_R1170_U64, new_P2_R1170_U65,
    new_P2_R1170_U66, new_P2_R1170_U67, new_P2_R1170_U68, new_P2_R1170_U69,
    new_P2_R1170_U70, new_P2_R1170_U71, new_P2_R1170_U72, new_P2_R1170_U73,
    new_P2_R1170_U74, new_P2_R1170_U75, new_P2_R1170_U76, new_P2_R1170_U77,
    new_P2_R1170_U78, new_P2_R1170_U79, new_P2_R1170_U80, new_P2_R1170_U81,
    new_P2_R1170_U82, new_P2_R1170_U83, new_P2_R1170_U84, new_P2_R1170_U85,
    new_P2_R1170_U86, new_P2_R1170_U87, new_P2_R1170_U88, new_P2_R1170_U89,
    new_P2_R1170_U90, new_P2_R1170_U91, new_P2_R1170_U92, new_P2_R1170_U93,
    new_P2_R1170_U94, new_P2_R1170_U95, new_P2_R1170_U96, new_P2_R1170_U97,
    new_P2_R1170_U98, new_P2_R1170_U99, new_P2_R1170_U100,
    new_P2_R1170_U101, new_P2_R1170_U102, new_P2_R1170_U103,
    new_P2_R1170_U104, new_P2_R1170_U105, new_P2_R1170_U106,
    new_P2_R1170_U107, new_P2_R1170_U108, new_P2_R1170_U109,
    new_P2_R1170_U110, new_P2_R1170_U111, new_P2_R1170_U112,
    new_P2_R1170_U113, new_P2_R1170_U114, new_P2_R1170_U115,
    new_P2_R1170_U116, new_P2_R1170_U117, new_P2_R1170_U118,
    new_P2_R1170_U119, new_P2_R1170_U120, new_P2_R1170_U121,
    new_P2_R1170_U122, new_P2_R1170_U123, new_P2_R1170_U124,
    new_P2_R1170_U125, new_P2_R1170_U126, new_P2_R1170_U127,
    new_P2_R1170_U128, new_P2_R1170_U129, new_P2_R1170_U130,
    new_P2_R1170_U131, new_P2_R1170_U132, new_P2_R1170_U133,
    new_P2_R1170_U134, new_P2_R1170_U135, new_P2_R1170_U136,
    new_P2_R1170_U137, new_P2_R1170_U138, new_P2_R1170_U139,
    new_P2_R1170_U140, new_P2_R1170_U141, new_P2_R1170_U142,
    new_P2_R1170_U143, new_P2_R1170_U144, new_P2_R1170_U145,
    new_P2_R1170_U146, new_P2_R1170_U147, new_P2_R1170_U148,
    new_P2_R1170_U149, new_P2_R1170_U150, new_P2_R1170_U151,
    new_P2_R1170_U152, new_P2_R1170_U153, new_P2_R1170_U154,
    new_P2_R1170_U155, new_P2_R1170_U156, new_P2_R1170_U157,
    new_P2_R1170_U158, new_P2_R1170_U159, new_P2_R1170_U160,
    new_P2_R1170_U161, new_P2_R1170_U162, new_P2_R1170_U163,
    new_P2_R1170_U164, new_P2_R1170_U165, new_P2_R1170_U166,
    new_P2_R1170_U167, new_P2_R1170_U168, new_P2_R1170_U169,
    new_P2_R1170_U170, new_P2_R1170_U171, new_P2_R1170_U172,
    new_P2_R1170_U173, new_P2_R1170_U174, new_P2_R1170_U175,
    new_P2_R1170_U176, new_P2_R1170_U177, new_P2_R1170_U178,
    new_P2_R1170_U179, new_P2_R1170_U180, new_P2_R1170_U181,
    new_P2_R1170_U182, new_P2_R1170_U183, new_P2_R1170_U184,
    new_P2_R1170_U185, new_P2_R1170_U186, new_P2_R1170_U187,
    new_P2_R1170_U188, new_P2_R1170_U189, new_P2_R1170_U190,
    new_P2_R1170_U191, new_P2_R1170_U192, new_P2_R1170_U193,
    new_P2_R1170_U194, new_P2_R1170_U195, new_P2_R1170_U196,
    new_P2_R1170_U197, new_P2_R1170_U198, new_P2_R1170_U199,
    new_P2_R1170_U200, new_P2_R1170_U201, new_P2_R1170_U202,
    new_P2_R1170_U203, new_P2_R1170_U204, new_P2_R1170_U205,
    new_P2_R1170_U206, new_P2_R1170_U207, new_P2_R1170_U208,
    new_P2_R1170_U209, new_P2_R1170_U210, new_P2_R1170_U211,
    new_P2_R1170_U212, new_P2_R1170_U213, new_P2_R1170_U214,
    new_P2_R1170_U215, new_P2_R1170_U216, new_P2_R1170_U217,
    new_P2_R1170_U218, new_P2_R1170_U219, new_P2_R1170_U220,
    new_P2_R1170_U221, new_P2_R1170_U222, new_P2_R1170_U223,
    new_P2_R1170_U224, new_P2_R1170_U225, new_P2_R1170_U226,
    new_P2_R1170_U227, new_P2_R1170_U228, new_P2_R1170_U229,
    new_P2_R1170_U230, new_P2_R1170_U231, new_P2_R1170_U232,
    new_P2_R1170_U233, new_P2_R1170_U234, new_P2_R1170_U235,
    new_P2_R1170_U236, new_P2_R1170_U237, new_P2_R1170_U238,
    new_P2_R1170_U239, new_P2_R1170_U240, new_P2_R1170_U241,
    new_P2_R1170_U242, new_P2_R1170_U243, new_P2_R1170_U244,
    new_P2_R1170_U245, new_P2_R1170_U246, new_P2_R1170_U247,
    new_P2_R1170_U248, new_P2_R1170_U249, new_P2_R1170_U250,
    new_P2_R1170_U251, new_P2_R1170_U252, new_P2_R1170_U253,
    new_P2_R1170_U254, new_P2_R1170_U255, new_P2_R1170_U256,
    new_P2_R1170_U257, new_P2_R1170_U258, new_P2_R1170_U259,
    new_P2_R1170_U260, new_P2_R1170_U261, new_P2_R1170_U262,
    new_P2_R1170_U263, new_P2_R1170_U264, new_P2_R1170_U265,
    new_P2_R1170_U266, new_P2_R1170_U267, new_P2_R1170_U268,
    new_P2_R1170_U269, new_P2_R1170_U270, new_P2_R1170_U271,
    new_P2_R1170_U272, new_P2_R1170_U273, new_P2_R1170_U274,
    new_P2_R1170_U275, new_P2_R1170_U276, new_P2_R1170_U277,
    new_P2_R1170_U278, new_P2_R1170_U279, new_P2_R1170_U280,
    new_P2_R1170_U281, new_P2_R1170_U282, new_P2_R1170_U283,
    new_P2_R1170_U284, new_P2_R1170_U285, new_P2_R1170_U286,
    new_P2_R1170_U287, new_P2_R1170_U288, new_P2_R1170_U289,
    new_P2_R1170_U290, new_P2_R1170_U291, new_P2_R1170_U292,
    new_P2_R1170_U293, new_P2_R1170_U294, new_P2_R1170_U295,
    new_P2_R1170_U296, new_P2_R1170_U297, new_P2_R1170_U298,
    new_P2_R1170_U299, new_P2_R1170_U300, new_P2_R1170_U301,
    new_P2_R1170_U302, new_P2_R1170_U303, new_P2_R1170_U304,
    new_P2_R1170_U305, new_P2_R1170_U306, new_P2_R1170_U307,
    new_P2_R1170_U308, new_P2_R1275_U6, new_P2_R1275_U7, new_P2_R1275_U8,
    new_P2_R1275_U9, new_P2_R1275_U10, new_P2_R1275_U11, new_P2_R1275_U12,
    new_P2_R1275_U13, new_P2_R1275_U14, new_P2_R1275_U15, new_P2_R1275_U16,
    new_P2_R1275_U17, new_P2_R1275_U18, new_P2_R1275_U19, new_P2_R1275_U20,
    new_P2_R1275_U21, new_P2_R1275_U22, new_P2_R1275_U23, new_P2_R1275_U24,
    new_P2_R1275_U25, new_P2_R1275_U26, new_P2_R1275_U27, new_P2_R1275_U28,
    new_P2_R1275_U29, new_P2_R1275_U30, new_P2_R1275_U31, new_P2_R1275_U32,
    new_P2_R1275_U33, new_P2_R1275_U34, new_P2_R1275_U35, new_P2_R1275_U36,
    new_P2_R1275_U37, new_P2_R1275_U38, new_P2_R1275_U39, new_P2_R1275_U40,
    new_P2_R1275_U41, new_P2_R1275_U42, new_P2_R1275_U43, new_P2_R1275_U44,
    new_P2_R1275_U45, new_P2_R1275_U46, new_P2_R1275_U47, new_P2_R1275_U48,
    new_P2_R1275_U49, new_P2_R1275_U50, new_P2_R1275_U51, new_P2_R1275_U52,
    new_P2_R1275_U53, new_P2_R1275_U54, new_P2_R1275_U55, new_P2_R1275_U56,
    new_P2_R1275_U57, new_P2_R1275_U58, new_P2_R1275_U59, new_P2_R1275_U60,
    new_P2_R1275_U61, new_P2_R1275_U62, new_P2_R1275_U63, new_P2_R1275_U64,
    new_P2_R1275_U65, new_P2_R1275_U66, new_P2_R1275_U67, new_P2_R1275_U68,
    new_P2_R1275_U69, new_P2_R1275_U70, new_P2_R1275_U71, new_P2_R1275_U72,
    new_P2_R1275_U73, new_P2_R1275_U74, new_P2_R1275_U75, new_P2_R1275_U76,
    new_P2_R1275_U77, new_P2_R1275_U78, new_P2_R1275_U79, new_P2_R1275_U80,
    new_P2_R1275_U81, new_P2_R1275_U82, new_P2_R1275_U83, new_P2_R1275_U84,
    new_P2_R1275_U85, new_P2_R1275_U86, new_P2_R1275_U87, new_P2_R1275_U88,
    new_P2_R1275_U89, new_P2_R1275_U90, new_P2_R1275_U91, new_P2_R1275_U92,
    new_P2_R1275_U93, new_P2_R1275_U94, new_P2_R1275_U95, new_P2_R1275_U96,
    new_P2_R1275_U97, new_P2_R1275_U98, new_P2_R1275_U99,
    new_P2_R1275_U100, new_P2_R1275_U101, new_P2_R1275_U102,
    new_P2_R1275_U103, new_P2_R1275_U104, new_P2_R1275_U105,
    new_P2_R1275_U106, new_P2_R1275_U107, new_P2_R1275_U108,
    new_P2_R1275_U109, new_P2_R1275_U110, new_P2_R1275_U111,
    new_P2_R1275_U112, new_P2_R1275_U113, new_P2_R1275_U114,
    new_P2_R1275_U115, new_P2_R1275_U116, new_P2_R1275_U117,
    new_P2_R1275_U118, new_P2_R1275_U119, new_P2_R1275_U120,
    new_P2_R1275_U121, new_P2_R1275_U122, new_P2_R1275_U123,
    new_P2_R1275_U124, new_P2_R1275_U125, new_P2_R1275_U126,
    new_P2_R1275_U127, new_P2_R1275_U128, new_P2_R1275_U129,
    new_P2_R1275_U130, new_P2_R1275_U131, new_P2_R1275_U132,
    new_P2_R1275_U133, new_P2_R1275_U134, new_P2_R1275_U135,
    new_P2_R1275_U136, new_P2_R1275_U137, new_P2_R1275_U138,
    new_P2_R1275_U139, new_P2_R1275_U140, new_P2_R1275_U141,
    new_P2_R1275_U142, new_P2_R1275_U143, new_P2_R1275_U144,
    new_P2_R1275_U145, new_P2_R1275_U146, new_P2_R1275_U147,
    new_P2_R1275_U148, new_P2_R1275_U149, new_P2_R1275_U150,
    new_P2_R1275_U151, new_P2_R1275_U152, new_P2_R1275_U153,
    new_P2_R1275_U154, new_P2_R1275_U155, new_P2_R1275_U156,
    new_P2_R1275_U157, new_P2_R1275_U158, new_P2_R1275_U159,
    new_P2_R1179_U6, new_P2_R1179_U7, new_P2_R1179_U8, new_P2_R1179_U9,
    new_P2_R1179_U10, new_P2_R1179_U11, new_P2_R1179_U12, new_P2_R1179_U13,
    new_P2_R1179_U14, new_P2_R1179_U15, new_P2_R1179_U16, new_P2_R1179_U17,
    new_P2_R1179_U18, new_P2_R1179_U19, new_P2_R1179_U20, new_P2_R1179_U21,
    new_P2_R1179_U22, new_P2_R1179_U23, new_P2_R1179_U24, new_P2_R1179_U25,
    new_P2_R1179_U26, new_P2_R1179_U27, new_P2_R1179_U28, new_P2_R1179_U29,
    new_P2_R1179_U30, new_P2_R1179_U31, new_P2_R1179_U32, new_P2_R1179_U33,
    new_P2_R1179_U34, new_P2_R1179_U35, new_P2_R1179_U36, new_P2_R1179_U37,
    new_P2_R1179_U38, new_P2_R1179_U39, new_P2_R1179_U40, new_P2_R1179_U41,
    new_P2_R1179_U42, new_P2_R1179_U43, new_P2_R1179_U44, new_P2_R1179_U45,
    new_P2_R1179_U46, new_P2_R1179_U47, new_P2_R1179_U48, new_P2_R1179_U49,
    new_P2_R1179_U50, new_P2_R1179_U51, new_P2_R1179_U52, new_P2_R1179_U53,
    new_P2_R1179_U54, new_P2_R1179_U55, new_P2_R1179_U56, new_P2_R1179_U57,
    new_P2_R1179_U58, new_P2_R1179_U59, new_P2_R1179_U60, new_P2_R1179_U61,
    new_P2_R1179_U62, new_P2_R1179_U63, new_P2_R1179_U64, new_P2_R1179_U65,
    new_P2_R1179_U66, new_P2_R1179_U67, new_P2_R1179_U68, new_P2_R1179_U69,
    new_P2_R1179_U70, new_P2_R1179_U71, new_P2_R1179_U72, new_P2_R1179_U73,
    new_P2_R1179_U74, new_P2_R1179_U75, new_P2_R1179_U76, new_P2_R1179_U77,
    new_P2_R1179_U78, new_P2_R1179_U79, new_P2_R1179_U80, new_P2_R1179_U81,
    new_P2_R1179_U82, new_P2_R1179_U83, new_P2_R1179_U84, new_P2_R1179_U85,
    new_P2_R1179_U86, new_P2_R1179_U87, new_P2_R1179_U88, new_P2_R1179_U89,
    new_P2_R1179_U90, new_P2_R1179_U91, new_P2_R1179_U92, new_P2_R1179_U93,
    new_P2_R1179_U94, new_P2_R1179_U95, new_P2_R1179_U96, new_P2_R1179_U97,
    new_P2_R1179_U98, new_P2_R1179_U99, new_P2_R1179_U100,
    new_P2_R1179_U101, new_P2_R1179_U102, new_P2_R1179_U103,
    new_P2_R1179_U104, new_P2_R1179_U105, new_P2_R1179_U106,
    new_P2_R1179_U107, new_P2_R1179_U108, new_P2_R1179_U109,
    new_P2_R1179_U110, new_P2_R1179_U111, new_P2_R1179_U112,
    new_P2_R1179_U113, new_P2_R1179_U114, new_P2_R1179_U115,
    new_P2_R1179_U116, new_P2_R1179_U117, new_P2_R1179_U118,
    new_P2_R1179_U119, new_P2_R1179_U120, new_P2_R1179_U121,
    new_P2_R1179_U122, new_P2_R1179_U123, new_P2_R1179_U124,
    new_P2_R1179_U125, new_P2_R1179_U126, new_P2_R1179_U127,
    new_P2_R1179_U128, new_P2_R1179_U129, new_P2_R1179_U130,
    new_P2_R1179_U131, new_P2_R1179_U132, new_P2_R1179_U133,
    new_P2_R1179_U134, new_P2_R1179_U135, new_P2_R1179_U136,
    new_P2_R1179_U137, new_P2_R1179_U138, new_P2_R1179_U139,
    new_P2_R1179_U140, new_P2_R1179_U141, new_P2_R1179_U142,
    new_P2_R1179_U143, new_P2_R1179_U144, new_P2_R1179_U145,
    new_P2_R1179_U146, new_P2_R1179_U147, new_P2_R1179_U148,
    new_P2_R1179_U149, new_P2_R1179_U150, new_P2_R1179_U151,
    new_P2_R1179_U152, new_P2_R1179_U153, new_P2_R1179_U154,
    new_P2_R1179_U155, new_P2_R1179_U156, new_P2_R1179_U157,
    new_P2_R1179_U158, new_P2_R1179_U159, new_P2_R1179_U160,
    new_P2_R1179_U161, new_P2_R1179_U162, new_P2_R1179_U163,
    new_P2_R1179_U164, new_P2_R1179_U165, new_P2_R1179_U166,
    new_P2_R1179_U167, new_P2_R1179_U168, new_P2_R1179_U169,
    new_P2_R1179_U170, new_P2_R1179_U171, new_P2_R1179_U172,
    new_P2_R1179_U173, new_P2_R1179_U174, new_P2_R1179_U175,
    new_P2_R1179_U176, new_P2_R1179_U177, new_P2_R1179_U178,
    new_P2_R1179_U179, new_P2_R1179_U180, new_P2_R1179_U181,
    new_P2_R1179_U182, new_P2_R1179_U183, new_P2_R1179_U184,
    new_P2_R1179_U185, new_P2_R1179_U186, new_P2_R1179_U187,
    new_P2_R1179_U188, new_P2_R1179_U189, new_P2_R1179_U190,
    new_P2_R1179_U191, new_P2_R1179_U192, new_P2_R1179_U193,
    new_P2_R1179_U194, new_P2_R1179_U195, new_P2_R1179_U196,
    new_P2_R1179_U197, new_P2_R1179_U198, new_P2_R1179_U199,
    new_P2_R1179_U200, new_P2_R1179_U201, new_P2_R1179_U202,
    new_P2_R1179_U203, new_P2_R1179_U204, new_P2_R1179_U205,
    new_P2_R1179_U206, new_P2_R1179_U207, new_P2_R1179_U208,
    new_P2_R1179_U209, new_P2_R1179_U210, new_P2_R1179_U211,
    new_P2_R1179_U212, new_P2_R1179_U213, new_P2_R1179_U214,
    new_P2_R1179_U215, new_P2_R1179_U216, new_P2_R1179_U217,
    new_P2_R1179_U218, new_P2_R1179_U219, new_P2_R1179_U220,
    new_P2_R1179_U221, new_P2_R1179_U222, new_P2_R1179_U223,
    new_P2_R1179_U224, new_P2_R1179_U225, new_P2_R1179_U226,
    new_P2_R1179_U227, new_P2_R1179_U228, new_P2_R1179_U229,
    new_P2_R1179_U230, new_P2_R1179_U231, new_P2_R1179_U232,
    new_P2_R1179_U233, new_P2_R1179_U234, new_P2_R1179_U235,
    new_P2_R1179_U236, new_P2_R1179_U237, new_P2_R1179_U238,
    new_P2_R1179_U239, new_P2_R1179_U240, new_P2_R1179_U241,
    new_P2_R1179_U242, new_P2_R1179_U243, new_P2_R1179_U244,
    new_P2_R1179_U245, new_P2_R1179_U246, new_P2_R1179_U247,
    new_P2_R1179_U248, new_P2_R1179_U249, new_P2_R1179_U250,
    new_P2_R1179_U251, new_P2_R1179_U252, new_P2_R1179_U253,
    new_P2_R1179_U254, new_P2_R1179_U255, new_P2_R1179_U256,
    new_P2_R1179_U257, new_P2_R1179_U258, new_P2_R1179_U259,
    new_P2_R1179_U260, new_P2_R1179_U261, new_P2_R1179_U262,
    new_P2_R1179_U263, new_P2_R1179_U264, new_P2_R1179_U265,
    new_P2_R1179_U266, new_P2_R1179_U267, new_P2_R1179_U268,
    new_P2_R1179_U269, new_P2_R1179_U270, new_P2_R1179_U271,
    new_P2_R1179_U272, new_P2_R1179_U273, new_P2_R1179_U274,
    new_P2_R1179_U275, new_P2_R1179_U276, new_P2_R1179_U277,
    new_P2_R1179_U278, new_P2_R1179_U279, new_P2_R1179_U280,
    new_P2_R1179_U281, new_P2_R1179_U282, new_P2_R1179_U283,
    new_P2_R1179_U284, new_P2_R1179_U285, new_P2_R1179_U286,
    new_P2_R1179_U287, new_P2_R1179_U288, new_P2_R1179_U289,
    new_P2_R1179_U290, new_P2_R1179_U291, new_P2_R1179_U292,
    new_P2_R1179_U293, new_P2_R1179_U294, new_P2_R1179_U295,
    new_P2_R1179_U296, new_P2_R1179_U297, new_P2_R1179_U298,
    new_P2_R1179_U299, new_P2_R1179_U300, new_P2_R1179_U301,
    new_P2_R1179_U302, new_P2_R1179_U303, new_P2_R1179_U304,
    new_P2_R1179_U305, new_P2_R1179_U306, new_P2_R1179_U307,
    new_P2_R1179_U308, new_P2_R1179_U309, new_P2_R1179_U310,
    new_P2_R1179_U311, new_P2_R1179_U312, new_P2_R1179_U313,
    new_P2_R1179_U314, new_P2_R1179_U315, new_P2_R1179_U316,
    new_P2_R1179_U317, new_P2_R1179_U318, new_P2_R1179_U319,
    new_P2_R1179_U320, new_P2_R1179_U321, new_P2_R1179_U322,
    new_P2_R1179_U323, new_P2_R1179_U324, new_P2_R1179_U325,
    new_P2_R1179_U326, new_P2_R1179_U327, new_P2_R1179_U328,
    new_P2_R1179_U329, new_P2_R1179_U330, new_P2_R1179_U331,
    new_P2_R1179_U332, new_P2_R1179_U333, new_P2_R1179_U334,
    new_P2_R1179_U335, new_P2_R1179_U336, new_P2_R1179_U337,
    new_P2_R1179_U338, new_P2_R1179_U339, new_P2_R1179_U340,
    new_P2_R1179_U341, new_P2_R1179_U342, new_P2_R1179_U343,
    new_P2_R1179_U344, new_P2_R1179_U345, new_P2_R1179_U346,
    new_P2_R1179_U347, new_P2_R1179_U348, new_P2_R1179_U349,
    new_P2_R1179_U350, new_P2_R1179_U351, new_P2_R1179_U352,
    new_P2_R1179_U353, new_P2_R1179_U354, new_P2_R1179_U355,
    new_P2_R1179_U356, new_P2_R1179_U357, new_P2_R1179_U358,
    new_P2_R1179_U359, new_P2_R1179_U360, new_P2_R1179_U361,
    new_P2_R1179_U362, new_P2_R1179_U363, new_P2_R1179_U364,
    new_P2_R1179_U365, new_P2_R1179_U366, new_P2_R1179_U367,
    new_P2_R1179_U368, new_P2_R1179_U369, new_P2_R1179_U370,
    new_P2_R1179_U371, new_P2_R1179_U372, new_P2_R1179_U373,
    new_P2_R1179_U374, new_P2_R1179_U375, new_P2_R1179_U376,
    new_P2_R1179_U377, new_P2_R1179_U378, new_P2_R1179_U379,
    new_P2_R1179_U380, new_P2_R1179_U381, new_P2_R1179_U382,
    new_P2_R1179_U383, new_P2_R1179_U384, new_P2_R1179_U385,
    new_P2_R1179_U386, new_P2_R1179_U387, new_P2_R1179_U388,
    new_P2_R1179_U389, new_P2_R1179_U390, new_P2_R1179_U391,
    new_P2_R1179_U392, new_P2_R1179_U393, new_P2_R1179_U394,
    new_P2_R1179_U395, new_P2_R1179_U396, new_P2_R1179_U397,
    new_P2_R1179_U398, new_P2_R1179_U399, new_P2_R1179_U400,
    new_P2_R1179_U401, new_P2_R1179_U402, new_P2_R1179_U403,
    new_P2_R1179_U404, new_P2_R1179_U405, new_P2_R1179_U406,
    new_P2_R1179_U407, new_P2_R1179_U408, new_P2_R1179_U409,
    new_P2_R1179_U410, new_P2_R1179_U411, new_P2_R1179_U412,
    new_P2_R1179_U413, new_P2_R1179_U414, new_P2_R1179_U415,
    new_P2_R1179_U416, new_P2_R1179_U417, new_P2_R1179_U418,
    new_P2_R1179_U419, new_P2_R1179_U420, new_P2_R1179_U421,
    new_P2_R1179_U422, new_P2_R1179_U423, new_P2_R1179_U424,
    new_P2_R1179_U425, new_P2_R1179_U426, new_P2_R1179_U427,
    new_P2_R1179_U428, new_P2_R1179_U429, new_P2_R1179_U430,
    new_P2_R1179_U431, new_P2_R1179_U432, new_P2_R1179_U433,
    new_P2_R1179_U434, new_P2_R1179_U435, new_P2_R1179_U436,
    new_P2_R1179_U437, new_P2_R1179_U438, new_P2_R1179_U439,
    new_P2_R1179_U440, new_P2_R1179_U441, new_P2_R1179_U442,
    new_P2_R1179_U443, new_P2_R1179_U444, new_P2_R1179_U445,
    new_P2_R1179_U446, new_P2_R1179_U447, new_P2_R1179_U448,
    new_P2_R1179_U449, new_P2_R1179_U450, new_P2_R1179_U451,
    new_P2_R1179_U452, new_P2_R1179_U453, new_P2_R1179_U454,
    new_P2_R1179_U455, new_P2_R1179_U456, new_P2_R1179_U457,
    new_P2_R1179_U458, new_P2_R1179_U459, new_P2_R1179_U460,
    new_P2_R1179_U461, new_P2_R1179_U462, new_P2_R1179_U463,
    new_P2_R1179_U464, new_P2_R1179_U465, new_P2_R1179_U466,
    new_P2_R1179_U467, new_P2_R1179_U468, new_P2_R1179_U469,
    new_P2_R1179_U470, new_P2_R1179_U471, new_P2_R1179_U472,
    new_P2_R1179_U473, new_P2_R1179_U474, new_P2_R1179_U475,
    new_P2_R1179_U476, new_P2_R1179_U477, new_P2_R1179_U478,
    new_P2_R1215_U4, new_P2_R1215_U5, new_P2_R1215_U6, new_P2_R1215_U7,
    new_P2_R1215_U8, new_P2_R1215_U9, new_P2_R1215_U10, new_P2_R1215_U11,
    new_P2_R1215_U12, new_P2_R1215_U13, new_P2_R1215_U14, new_P2_R1215_U15,
    new_P2_R1215_U16, new_P2_R1215_U17, new_P2_R1215_U18, new_P2_R1215_U19,
    new_P2_R1215_U20, new_P2_R1215_U21, new_P2_R1215_U22, new_P2_R1215_U23,
    new_P2_R1215_U24, new_P2_R1215_U25, new_P2_R1215_U26, new_P2_R1215_U27,
    new_P2_R1215_U28, new_P2_R1215_U29, new_P2_R1215_U30, new_P2_R1215_U31,
    new_P2_R1215_U32, new_P2_R1215_U33, new_P2_R1215_U34, new_P2_R1215_U35,
    new_P2_R1215_U36, new_P2_R1215_U37, new_P2_R1215_U38, new_P2_R1215_U39,
    new_P2_R1215_U40, new_P2_R1215_U41, new_P2_R1215_U42, new_P2_R1215_U43,
    new_P2_R1215_U44, new_P2_R1215_U45, new_P2_R1215_U46, new_P2_R1215_U47,
    new_P2_R1215_U48, new_P2_R1215_U49, new_P2_R1215_U50, new_P2_R1215_U51,
    new_P2_R1215_U52, new_P2_R1215_U53, new_P2_R1215_U54, new_P2_R1215_U55,
    new_P2_R1215_U56, new_P2_R1215_U57, new_P2_R1215_U58, new_P2_R1215_U59,
    new_P2_R1215_U60, new_P2_R1215_U61, new_P2_R1215_U62, new_P2_R1215_U63,
    new_P2_R1215_U64, new_P2_R1215_U65, new_P2_R1215_U66, new_P2_R1215_U67,
    new_P2_R1215_U68, new_P2_R1215_U69, new_P2_R1215_U70, new_P2_R1215_U71,
    new_P2_R1215_U72, new_P2_R1215_U73, new_P2_R1215_U74, new_P2_R1215_U75,
    new_P2_R1215_U76, new_P2_R1215_U77, new_P2_R1215_U78, new_P2_R1215_U79,
    new_P2_R1215_U80, new_P2_R1215_U81, new_P2_R1215_U82, new_P2_R1215_U83,
    new_P2_R1215_U84, new_P2_R1215_U85, new_P2_R1215_U86, new_P2_R1215_U87,
    new_P2_R1215_U88, new_P2_R1215_U89, new_P2_R1215_U90, new_P2_R1215_U91,
    new_P2_R1215_U92, new_P2_R1215_U93, new_P2_R1215_U94, new_P2_R1215_U95,
    new_P2_R1215_U96, new_P2_R1215_U97, new_P2_R1215_U98, new_P2_R1215_U99,
    new_P2_R1215_U100, new_P2_R1215_U101, new_P2_R1215_U102,
    new_P2_R1215_U103, new_P2_R1215_U104, new_P2_R1215_U105,
    new_P2_R1215_U106, new_P2_R1215_U107, new_P2_R1215_U108,
    new_P2_R1215_U109, new_P2_R1215_U110, new_P2_R1215_U111,
    new_P2_R1215_U112, new_P2_R1215_U113, new_P2_R1215_U114,
    new_P2_R1215_U115, new_P2_R1215_U116, new_P2_R1215_U117,
    new_P2_R1215_U118, new_P2_R1215_U119, new_P2_R1215_U120,
    new_P2_R1215_U121, new_P2_R1215_U122, new_P2_R1215_U123,
    new_P2_R1215_U124, new_P2_R1215_U125, new_P2_R1215_U126,
    new_P2_R1215_U127, new_P2_R1215_U128, new_P2_R1215_U129,
    new_P2_R1215_U130, new_P2_R1215_U131, new_P2_R1215_U132,
    new_P2_R1215_U133, new_P2_R1215_U134, new_P2_R1215_U135,
    new_P2_R1215_U136, new_P2_R1215_U137, new_P2_R1215_U138,
    new_P2_R1215_U139, new_P2_R1215_U140, new_P2_R1215_U141,
    new_P2_R1215_U142, new_P2_R1215_U143, new_P2_R1215_U144,
    new_P2_R1215_U145, new_P2_R1215_U146, new_P2_R1215_U147,
    new_P2_R1215_U148, new_P2_R1215_U149, new_P2_R1215_U150,
    new_P2_R1215_U151, new_P2_R1215_U152, new_P2_R1215_U153,
    new_P2_R1215_U154, new_P2_R1215_U155, new_P2_R1215_U156,
    new_P2_R1215_U157, new_P2_R1215_U158, new_P2_R1215_U159,
    new_P2_R1215_U160, new_P2_R1215_U161, new_P2_R1215_U162,
    new_P2_R1215_U163, new_P2_R1215_U164, new_P2_R1215_U165,
    new_P2_R1215_U166, new_P2_R1215_U167, new_P2_R1215_U168,
    new_P2_R1215_U169, new_P2_R1215_U170, new_P2_R1215_U171,
    new_P2_R1215_U172, new_P2_R1215_U173, new_P2_R1215_U174,
    new_P2_R1215_U175, new_P2_R1215_U176, new_P2_R1215_U177,
    new_P2_R1215_U178, new_P2_R1215_U179, new_P2_R1215_U180,
    new_P2_R1215_U181, new_P2_R1215_U182, new_P2_R1215_U183,
    new_P2_R1215_U184, new_P2_R1215_U185, new_P2_R1215_U186,
    new_P2_R1215_U187, new_P2_R1215_U188, new_P2_R1215_U189,
    new_P2_R1215_U190, new_P2_R1215_U191, new_P2_R1215_U192,
    new_P2_R1215_U193, new_P2_R1215_U194, new_P2_R1215_U195,
    new_P2_R1215_U196, new_P2_R1215_U197, new_P2_R1215_U198,
    new_P2_R1215_U199, new_P2_R1215_U200, new_P2_R1215_U201,
    new_P2_R1215_U202, new_P2_R1215_U203, new_P2_R1215_U204,
    new_P2_R1215_U205, new_P2_R1215_U206, new_P2_R1215_U207,
    new_P2_R1215_U208, new_P2_R1215_U209, new_P2_R1215_U210,
    new_P2_R1215_U211, new_P2_R1215_U212, new_P2_R1215_U213,
    new_P2_R1215_U214, new_P2_R1215_U215, new_P2_R1215_U216,
    new_P2_R1215_U217, new_P2_R1215_U218, new_P2_R1215_U219,
    new_P2_R1215_U220, new_P2_R1215_U221, new_P2_R1215_U222,
    new_P2_R1215_U223, new_P2_R1215_U224, new_P2_R1215_U225,
    new_P2_R1215_U226, new_P2_R1215_U227, new_P2_R1215_U228,
    new_P2_R1215_U229, new_P2_R1215_U230, new_P2_R1215_U231,
    new_P2_R1215_U232, new_P2_R1215_U233, new_P2_R1215_U234,
    new_P2_R1215_U235, new_P2_R1215_U236, new_P2_R1215_U237,
    new_P2_R1215_U238, new_P2_R1215_U239, new_P2_R1215_U240,
    new_P2_R1215_U241, new_P2_R1215_U242, new_P2_R1215_U243,
    new_P2_R1215_U244, new_P2_R1215_U245, new_P2_R1215_U246,
    new_P2_R1215_U247, new_P2_R1215_U248, new_P2_R1215_U249,
    new_P2_R1215_U250, new_P2_R1215_U251, new_P2_R1215_U252,
    new_P2_R1215_U253, new_P2_R1215_U254, new_P2_R1215_U255,
    new_P2_R1215_U256, new_P2_R1215_U257, new_P2_R1215_U258,
    new_P2_R1215_U259, new_P2_R1215_U260, new_P2_R1215_U261,
    new_P2_R1215_U262, new_P2_R1215_U263, new_P2_R1215_U264,
    new_P2_R1215_U265, new_P2_R1215_U266, new_P2_R1215_U267,
    new_P2_R1215_U268, new_P2_R1215_U269, new_P2_R1215_U270,
    new_P2_R1215_U271, new_P2_R1215_U272, new_P2_R1215_U273,
    new_P2_R1215_U274, new_P2_R1215_U275, new_P2_R1215_U276,
    new_P2_R1215_U277, new_P2_R1215_U278, new_P2_R1215_U279,
    new_P2_R1215_U280, new_P2_R1215_U281, new_P2_R1215_U282,
    new_P2_R1215_U283, new_P2_R1215_U284, new_P2_R1215_U285,
    new_P2_R1215_U286, new_P2_R1215_U287, new_P2_R1215_U288,
    new_P2_R1215_U289, new_P2_R1215_U290, new_P2_R1215_U291,
    new_P2_R1215_U292, new_P2_R1215_U293, new_P2_R1215_U294,
    new_P2_R1215_U295, new_P2_R1215_U296, new_P2_R1215_U297,
    new_P2_R1215_U298, new_P2_R1215_U299, new_P2_R1215_U300,
    new_P2_R1215_U301, new_P2_R1215_U302, new_P2_R1215_U303,
    new_P2_R1215_U304, new_P2_R1215_U305, new_P2_R1215_U306,
    new_P2_R1215_U307, new_P2_R1215_U308, new_P2_R1215_U309,
    new_P2_R1215_U310, new_P2_R1215_U311, new_P2_R1215_U312,
    new_P2_R1215_U313, new_P2_R1215_U314, new_P2_R1215_U315,
    new_P2_R1215_U316, new_P2_R1215_U317, new_P2_R1215_U318,
    new_P2_R1215_U319, new_P2_R1215_U320, new_P2_R1215_U321,
    new_P2_R1215_U322, new_P2_R1215_U323, new_P2_R1215_U324,
    new_P2_R1215_U325, new_P2_R1215_U326, new_P2_R1215_U327,
    new_P2_R1215_U328, new_P2_R1215_U329, new_P2_R1215_U330,
    new_P2_R1215_U331, new_P2_R1215_U332, new_P2_R1215_U333,
    new_P2_R1215_U334, new_P2_R1215_U335, new_P2_R1215_U336,
    new_P2_R1215_U337, new_P2_R1215_U338, new_P2_R1215_U339,
    new_P2_R1215_U340, new_P2_R1215_U341, new_P2_R1215_U342,
    new_P2_R1215_U343, new_P2_R1215_U344, new_P2_R1215_U345,
    new_P2_R1215_U346, new_P2_R1215_U347, new_P2_R1215_U348,
    new_P2_R1215_U349, new_P2_R1215_U350, new_P2_R1215_U351,
    new_P2_R1215_U352, new_P2_R1215_U353, new_P2_R1215_U354,
    new_P2_R1215_U355, new_P2_R1215_U356, new_P2_R1215_U357,
    new_P2_R1215_U358, new_P2_R1215_U359, new_P2_R1215_U360,
    new_P2_R1215_U361, new_P2_R1215_U362, new_P2_R1215_U363,
    new_P2_R1215_U364, new_P2_R1215_U365, new_P2_R1215_U366,
    new_P2_R1215_U367, new_P2_R1215_U368, new_P2_R1215_U369,
    new_P2_R1215_U370, new_P2_R1215_U371, new_P2_R1215_U372,
    new_P2_R1215_U373, new_P2_R1215_U374, new_P2_R1215_U375,
    new_P2_R1215_U376, new_P2_R1215_U377, new_P2_R1215_U378,
    new_P2_R1215_U379, new_P2_R1215_U380, new_P2_R1215_U381,
    new_P2_R1215_U382, new_P2_R1215_U383, new_P2_R1215_U384,
    new_P2_R1215_U385, new_P2_R1215_U386, new_P2_R1215_U387,
    new_P2_R1215_U388, new_P2_R1215_U389, new_P2_R1215_U390,
    new_P2_R1215_U391, new_P2_R1215_U392, new_P2_R1215_U393,
    new_P2_R1215_U394, new_P2_R1215_U395, new_P2_R1215_U396,
    new_P2_R1215_U397, new_P2_R1215_U398, new_P2_R1215_U399,
    new_P2_R1215_U400, new_P2_R1215_U401, new_P2_R1215_U402,
    new_P2_R1215_U403, new_P2_R1215_U404, new_P2_R1215_U405,
    new_P2_R1215_U406, new_P2_R1215_U407, new_P2_R1215_U408,
    new_P2_R1215_U409, new_P2_R1215_U410, new_P2_R1215_U411,
    new_P2_R1215_U412, new_P2_R1215_U413, new_P2_R1215_U414,
    new_P2_R1215_U415, new_P2_R1215_U416, new_P2_R1215_U417,
    new_P2_R1215_U418, new_P2_R1215_U419, new_P2_R1215_U420,
    new_P2_R1215_U421, new_P2_R1215_U422, new_P2_R1215_U423,
    new_P2_R1215_U424, new_P2_R1215_U425, new_P2_R1215_U426,
    new_P2_R1215_U427, new_P2_R1215_U428, new_P2_R1215_U429,
    new_P2_R1215_U430, new_P2_R1215_U431, new_P2_R1215_U432,
    new_P2_R1215_U433, new_P2_R1215_U434, new_P2_R1215_U435,
    new_P2_R1215_U436, new_P2_R1215_U437, new_P2_R1215_U438,
    new_P2_R1215_U439, new_P2_R1215_U440, new_P2_R1215_U441,
    new_P2_R1215_U442, new_P2_R1215_U443, new_P2_R1215_U444,
    new_P2_R1215_U445, new_P2_R1215_U446, new_P2_R1215_U447,
    new_P2_R1215_U448, new_P2_R1215_U449, new_P2_R1215_U450,
    new_P2_R1215_U451, new_P2_R1215_U452, new_P2_R1215_U453,
    new_P2_R1215_U454, new_P2_R1215_U455, new_P2_R1215_U456,
    new_P2_R1215_U457, new_P2_R1215_U458, new_P2_R1215_U459,
    new_P2_R1215_U460, new_P2_R1215_U461, new_P2_R1215_U462,
    new_P2_R1215_U463, new_P2_R1215_U464, new_P2_R1215_U465,
    new_P2_R1215_U466, new_P2_R1215_U467, new_P2_R1215_U468,
    new_P2_R1215_U469, new_P2_R1215_U470, new_P2_R1215_U471,
    new_P2_R1215_U472, new_P2_R1215_U473, new_P2_R1215_U474,
    new_P2_R1215_U475, new_P2_R1215_U476, new_P2_R1215_U477,
    new_P2_R1215_U478, new_P2_R1215_U479, new_P2_R1215_U480,
    new_P2_R1215_U481, new_P2_R1215_U482, new_P2_R1215_U483,
    new_P2_R1215_U484, new_P2_R1215_U485, new_P2_R1215_U486,
    new_P2_R1215_U487, new_P2_R1215_U488, new_P2_R1215_U489,
    new_P2_R1215_U490, new_P2_R1215_U491, new_P2_R1215_U492,
    new_P2_R1215_U493, new_P2_R1215_U494, new_P2_R1215_U495,
    new_P2_R1215_U496, new_P2_R1215_U497, new_P2_R1215_U498,
    new_P2_R1215_U499, new_P2_R1215_U500, new_P2_R1215_U501,
    new_P2_R1215_U502, new_P2_R1215_U503, new_P2_R1215_U504,
    new_P2_R1164_U4, new_P2_R1164_U5, new_P2_R1164_U6, new_P2_R1164_U7,
    new_P2_R1164_U8, new_P2_R1164_U9, new_P2_R1164_U10, new_P2_R1164_U11,
    new_P2_R1164_U12, new_P2_R1164_U13, new_P2_R1164_U14, new_P2_R1164_U15,
    new_P2_R1164_U16, new_P2_R1164_U17, new_P2_R1164_U18, new_P2_R1164_U19,
    new_P2_R1164_U20, new_P2_R1164_U21, new_P2_R1164_U22, new_P2_R1164_U23,
    new_P2_R1164_U24, new_P2_R1164_U25, new_P2_R1164_U26, new_P2_R1164_U27,
    new_P2_R1164_U28, new_P2_R1164_U29, new_P2_R1164_U30, new_P2_R1164_U31,
    new_P2_R1164_U32, new_P2_R1164_U33, new_P2_R1164_U34, new_P2_R1164_U35,
    new_P2_R1164_U36, new_P2_R1164_U37, new_P2_R1164_U38, new_P2_R1164_U39,
    new_P2_R1164_U40, new_P2_R1164_U41, new_P2_R1164_U42, new_P2_R1164_U43,
    new_P2_R1164_U44, new_P2_R1164_U45, new_P2_R1164_U46, new_P2_R1164_U47,
    new_P2_R1164_U48, new_P2_R1164_U49, new_P2_R1164_U50, new_P2_R1164_U51,
    new_P2_R1164_U52, new_P2_R1164_U53, new_P2_R1164_U54, new_P2_R1164_U55,
    new_P2_R1164_U56, new_P2_R1164_U57, new_P2_R1164_U58, new_P2_R1164_U59,
    new_P2_R1164_U60, new_P2_R1164_U61, new_P2_R1164_U62, new_P2_R1164_U63,
    new_P2_R1164_U64, new_P2_R1164_U65, new_P2_R1164_U66, new_P2_R1164_U67,
    new_P2_R1164_U68, new_P2_R1164_U69, new_P2_R1164_U70, new_P2_R1164_U71,
    new_P2_R1164_U72, new_P2_R1164_U73, new_P2_R1164_U74, new_P2_R1164_U75,
    new_P2_R1164_U76, new_P2_R1164_U77, new_P2_R1164_U78, new_P2_R1164_U79,
    new_P2_R1164_U80, new_P2_R1164_U81, new_P2_R1164_U82, new_P2_R1164_U83,
    new_P2_R1164_U84, new_P2_R1164_U85, new_P2_R1164_U86, new_P2_R1164_U87,
    new_P2_R1164_U88, new_P2_R1164_U89, new_P2_R1164_U90, new_P2_R1164_U91,
    new_P2_R1164_U92, new_P2_R1164_U93, new_P2_R1164_U94, new_P2_R1164_U95,
    new_P2_R1164_U96, new_P2_R1164_U97, new_P2_R1164_U98, new_P2_R1164_U99,
    new_P2_R1164_U100, new_P2_R1164_U101, new_P2_R1164_U102,
    new_P2_R1164_U103, new_P2_R1164_U104, new_P2_R1164_U105,
    new_P2_R1164_U106, new_P2_R1164_U107, new_P2_R1164_U108,
    new_P2_R1164_U109, new_P2_R1164_U110, new_P2_R1164_U111,
    new_P2_R1164_U112, new_P2_R1164_U113, new_P2_R1164_U114,
    new_P2_R1164_U115, new_P2_R1164_U116, new_P2_R1164_U117,
    new_P2_R1164_U118, new_P2_R1164_U119, new_P2_R1164_U120,
    new_P2_R1164_U121, new_P2_R1164_U122, new_P2_R1164_U123,
    new_P2_R1164_U124, new_P2_R1164_U125, new_P2_R1164_U126,
    new_P2_R1164_U127, new_P2_R1164_U128, new_P2_R1164_U129,
    new_P2_R1164_U130, new_P2_R1164_U131, new_P2_R1164_U132,
    new_P2_R1164_U133, new_P2_R1164_U134, new_P2_R1164_U135,
    new_P2_R1164_U136, new_P2_R1164_U137, new_P2_R1164_U138,
    new_P2_R1164_U139, new_P2_R1164_U140, new_P2_R1164_U141,
    new_P2_R1164_U142, new_P2_R1164_U143, new_P2_R1164_U144,
    new_P2_R1164_U145, new_P2_R1164_U146, new_P2_R1164_U147,
    new_P2_R1164_U148, new_P2_R1164_U149, new_P2_R1164_U150,
    new_P2_R1164_U151, new_P2_R1164_U152, new_P2_R1164_U153,
    new_P2_R1164_U154, new_P2_R1164_U155, new_P2_R1164_U156,
    new_P2_R1164_U157, new_P2_R1164_U158, new_P2_R1164_U159,
    new_P2_R1164_U160, new_P2_R1164_U161, new_P2_R1164_U162,
    new_P2_R1164_U163, new_P2_R1164_U164, new_P2_R1164_U165,
    new_P2_R1164_U166, new_P2_R1164_U167, new_P2_R1164_U168,
    new_P2_R1164_U169, new_P2_R1164_U170, new_P2_R1164_U171,
    new_P2_R1164_U172, new_P2_R1164_U173, new_P2_R1164_U174,
    new_P2_R1164_U175, new_P2_R1164_U176, new_P2_R1164_U177,
    new_P2_R1164_U178, new_P2_R1164_U179, new_P2_R1164_U180,
    new_P2_R1164_U181, new_P2_R1164_U182, new_P2_R1164_U183,
    new_P2_R1164_U184, new_P2_R1164_U185, new_P2_R1164_U186,
    new_P2_R1164_U187, new_P2_R1164_U188, new_P2_R1164_U189,
    new_P2_R1164_U190, new_P2_R1164_U191, new_P2_R1164_U192,
    new_P2_R1164_U193, new_P2_R1164_U194, new_P2_R1164_U195,
    new_P2_R1164_U196, new_P2_R1164_U197, new_P2_R1164_U198,
    new_P2_R1164_U199, new_P2_R1164_U200, new_P2_R1164_U201,
    new_P2_R1164_U202, new_P2_R1164_U203, new_P2_R1164_U204,
    new_P2_R1164_U205, new_P2_R1164_U206, new_P2_R1164_U207,
    new_P2_R1164_U208, new_P2_R1164_U209, new_P2_R1164_U210,
    new_P2_R1164_U211, new_P2_R1164_U212, new_P2_R1164_U213,
    new_P2_R1164_U214, new_P2_R1164_U215, new_P2_R1164_U216,
    new_P2_R1164_U217, new_P2_R1164_U218, new_P2_R1164_U219,
    new_P2_R1164_U220, new_P2_R1164_U221, new_P2_R1164_U222,
    new_P2_R1164_U223, new_P2_R1164_U224, new_P2_R1164_U225,
    new_P2_R1164_U226, new_P2_R1164_U227, new_P2_R1164_U228,
    new_P2_R1164_U229, new_P2_R1164_U230, new_P2_R1164_U231,
    new_P2_R1164_U232, new_P2_R1164_U233, new_P2_R1164_U234,
    new_P2_R1164_U235, new_P2_R1164_U236, new_P2_R1164_U237,
    new_P2_R1164_U238, new_P2_R1164_U239, new_P2_R1164_U240,
    new_P2_R1164_U241, new_P2_R1164_U242, new_P2_R1164_U243,
    new_P2_R1164_U244, new_P2_R1164_U245, new_P2_R1164_U246,
    new_P2_R1164_U247, new_P2_R1164_U248, new_P2_R1164_U249,
    new_P2_R1164_U250, new_P2_R1164_U251, new_P2_R1164_U252,
    new_P2_R1164_U253, new_P2_R1164_U254, new_P2_R1164_U255,
    new_P2_R1164_U256, new_P2_R1164_U257, new_P2_R1164_U258,
    new_P2_R1164_U259, new_P2_R1164_U260, new_P2_R1164_U261,
    new_P2_R1164_U262, new_P2_R1164_U263, new_P2_R1164_U264,
    new_P2_R1164_U265, new_P2_R1164_U266, new_P2_R1164_U267,
    new_P2_R1164_U268, new_P2_R1164_U269, new_P2_R1164_U270,
    new_P2_R1164_U271, new_P2_R1164_U272, new_P2_R1164_U273,
    new_P2_R1164_U274, new_P2_R1164_U275, new_P2_R1164_U276,
    new_P2_R1164_U277, new_P2_R1164_U278, new_P2_R1164_U279,
    new_P2_R1164_U280, new_P2_R1164_U281, new_P2_R1164_U282,
    new_P2_R1164_U283, new_P2_R1164_U284, new_P2_R1164_U285,
    new_P2_R1164_U286, new_P2_R1164_U287, new_P2_R1164_U288,
    new_P2_R1164_U289, new_P2_R1164_U290, new_P2_R1164_U291,
    new_P2_R1164_U292, new_P2_R1164_U293, new_P2_R1164_U294,
    new_P2_R1164_U295, new_P2_R1164_U296, new_P2_R1164_U297,
    new_P2_R1164_U298, new_P2_R1164_U299, new_P2_R1164_U300,
    new_P2_R1164_U301, new_P2_R1164_U302, new_P2_R1164_U303,
    new_P2_R1164_U304, new_P2_R1164_U305, new_P2_R1164_U306,
    new_P2_R1164_U307, new_P2_R1164_U308, new_P2_R1164_U309,
    new_P2_R1164_U310, new_P2_R1164_U311, new_P2_R1164_U312,
    new_P2_R1164_U313, new_P2_R1164_U314, new_P2_R1164_U315,
    new_P2_R1164_U316, new_P2_R1164_U317, new_P2_R1164_U318,
    new_P2_R1164_U319, new_P2_R1164_U320, new_P2_R1164_U321,
    new_P2_R1164_U322, new_P2_R1164_U323, new_P2_R1164_U324,
    new_P2_R1164_U325, new_P2_R1164_U326, new_P2_R1164_U327,
    new_P2_R1164_U328, new_P2_R1164_U329, new_P2_R1164_U330,
    new_P2_R1164_U331, new_P2_R1164_U332, new_P2_R1164_U333,
    new_P2_R1164_U334, new_P2_R1164_U335, new_P2_R1164_U336,
    new_P2_R1164_U337, new_P2_R1164_U338, new_P2_R1164_U339,
    new_P2_R1164_U340, new_P2_R1164_U341, new_P2_R1164_U342,
    new_P2_R1164_U343, new_P2_R1164_U344, new_P2_R1164_U345,
    new_P2_R1164_U346, new_P2_R1164_U347, new_P2_R1164_U348,
    new_P2_R1164_U349, new_P2_R1164_U350, new_P2_R1164_U351,
    new_P2_R1164_U352, new_P2_R1164_U353, new_P2_R1164_U354,
    new_P2_R1164_U355, new_P2_R1164_U356, new_P2_R1164_U357,
    new_P2_R1164_U358, new_P2_R1164_U359, new_P2_R1164_U360,
    new_P2_R1164_U361, new_P2_R1164_U362, new_P2_R1164_U363,
    new_P2_R1164_U364, new_P2_R1164_U365, new_P2_R1164_U366,
    new_P2_R1164_U367, new_P2_R1164_U368, new_P2_R1164_U369,
    new_P2_R1164_U370, new_P2_R1164_U371, new_P2_R1164_U372,
    new_P2_R1164_U373, new_P2_R1164_U374, new_P2_R1164_U375,
    new_P2_R1164_U376, new_P2_R1164_U377, new_P2_R1164_U378,
    new_P2_R1164_U379, new_P2_R1164_U380, new_P2_R1164_U381,
    new_P2_R1164_U382, new_P2_R1164_U383, new_P2_R1164_U384,
    new_P2_R1164_U385, new_P2_R1164_U386, new_P2_R1164_U387,
    new_P2_R1164_U388, new_P2_R1164_U389, new_P2_R1164_U390,
    new_P2_R1164_U391, new_P2_R1164_U392, new_P2_R1164_U393,
    new_P2_R1164_U394, new_P2_R1164_U395, new_P2_R1164_U396,
    new_P2_R1164_U397, new_P2_R1164_U398, new_P2_R1164_U399,
    new_P2_R1164_U400, new_P2_R1164_U401, new_P2_R1164_U402,
    new_P2_R1164_U403, new_P2_R1164_U404, new_P2_R1164_U405,
    new_P2_R1164_U406, new_P2_R1164_U407, new_P2_R1164_U408,
    new_P2_R1164_U409, new_P2_R1164_U410, new_P2_R1164_U411,
    new_P2_R1164_U412, new_P2_R1164_U413, new_P2_R1164_U414,
    new_P2_R1164_U415, new_P2_R1164_U416, new_P2_R1164_U417,
    new_P2_R1164_U418, new_P2_R1164_U419, new_P2_R1164_U420,
    new_P2_R1164_U421, new_P2_R1164_U422, new_P2_R1164_U423,
    new_P2_R1164_U424, new_P2_R1164_U425, new_P2_R1164_U426,
    new_P2_R1164_U427, new_P2_R1164_U428, new_P2_R1164_U429,
    new_P2_R1164_U430, new_P2_R1164_U431, new_P2_R1164_U432,
    new_P2_R1164_U433, new_P2_R1164_U434, new_P2_R1164_U435,
    new_P2_R1164_U436, new_P2_R1164_U437, new_P2_R1164_U438,
    new_P2_R1164_U439, new_P2_R1164_U440, new_P2_R1164_U441,
    new_P2_R1164_U442, new_P2_R1164_U443, new_P2_R1164_U444,
    new_P2_R1164_U445, new_P2_R1164_U446, new_P2_R1164_U447,
    new_P2_R1164_U448, new_P2_R1164_U449, new_P2_R1164_U450,
    new_P2_R1164_U451, new_P2_R1164_U452, new_P2_R1164_U453,
    new_P2_R1164_U454, new_P2_R1164_U455, new_P2_R1164_U456,
    new_P2_R1164_U457, new_P2_R1164_U458, new_P2_R1164_U459,
    new_P2_R1164_U460, new_P2_R1164_U461, new_P2_R1164_U462,
    new_P2_R1164_U463, new_P2_R1164_U464, new_P2_R1164_U465,
    new_P2_R1164_U466, new_P2_R1164_U467, new_P2_R1164_U468,
    new_P2_R1164_U469, new_P2_R1164_U470, new_P2_R1164_U471,
    new_P2_R1164_U472, new_P2_R1164_U473, new_P2_R1164_U474,
    new_P2_R1164_U475, new_P2_R1164_U476, new_P2_R1164_U477,
    new_P2_R1164_U478, new_P2_R1164_U479, new_P2_R1164_U480,
    new_P2_R1164_U481, new_P2_R1164_U482, new_P2_R1164_U483,
    new_P2_R1164_U484, new_P2_R1164_U485, new_P2_R1164_U486,
    new_P2_R1164_U487, new_P2_R1164_U488, new_P2_R1164_U489,
    new_P2_R1164_U490, new_P2_R1164_U491, new_P2_R1164_U492,
    new_P2_R1164_U493, new_P2_R1164_U494, new_P2_R1164_U495,
    new_P2_R1164_U496, new_P2_R1164_U497, new_P2_R1164_U498,
    new_P2_R1164_U499, new_P2_R1164_U500, new_P2_R1164_U501,
    new_P2_R1164_U502, new_P2_R1164_U503, new_P2_R1164_U504,
    new_P2_R1233_U4, new_P2_R1233_U5, new_P2_R1233_U6, new_P2_R1233_U7,
    new_P2_R1233_U8, new_P2_R1233_U9, new_P2_R1233_U10, new_P2_R1233_U11,
    new_P2_R1233_U12, new_P2_R1233_U13, new_P2_R1233_U14, new_P2_R1233_U15,
    new_P2_R1233_U16, new_P2_R1233_U17, new_P2_R1233_U18, new_P2_R1233_U19,
    new_P2_R1233_U20, new_P2_R1233_U21, new_P2_R1233_U22, new_P2_R1233_U23,
    new_P2_R1233_U24, new_P2_R1233_U25, new_P2_R1233_U26, new_P2_R1233_U27,
    new_P2_R1233_U28, new_P2_R1233_U29, new_P2_R1233_U30, new_P2_R1233_U31,
    new_P2_R1233_U32, new_P2_R1233_U33, new_P2_R1233_U34, new_P2_R1233_U35,
    new_P2_R1233_U36, new_P2_R1233_U37, new_P2_R1233_U38, new_P2_R1233_U39,
    new_P2_R1233_U40, new_P2_R1233_U41, new_P2_R1233_U42, new_P2_R1233_U43,
    new_P2_R1233_U44, new_P2_R1233_U45, new_P2_R1233_U46, new_P2_R1233_U47,
    new_P2_R1233_U48, new_P2_R1233_U49, new_P2_R1233_U50, new_P2_R1233_U51,
    new_P2_R1233_U52, new_P2_R1233_U53, new_P2_R1233_U54, new_P2_R1233_U55,
    new_P2_R1233_U56, new_P2_R1233_U57, new_P2_R1233_U58, new_P2_R1233_U59,
    new_P2_R1233_U60, new_P2_R1233_U61, new_P2_R1233_U62, new_P2_R1233_U63,
    new_P2_R1233_U64, new_P2_R1233_U65, new_P2_R1233_U66, new_P2_R1233_U67,
    new_P2_R1233_U68, new_P2_R1233_U69, new_P2_R1233_U70, new_P2_R1233_U71,
    new_P2_R1233_U72, new_P2_R1233_U73, new_P2_R1233_U74, new_P2_R1233_U75,
    new_P2_R1233_U76, new_P2_R1233_U77, new_P2_R1233_U78, new_P2_R1233_U79,
    new_P2_R1233_U80, new_P2_R1233_U81, new_P2_R1233_U82, new_P2_R1233_U83,
    new_P2_R1233_U84, new_P2_R1233_U85, new_P2_R1233_U86, new_P2_R1233_U87,
    new_P2_R1233_U88, new_P2_R1233_U89, new_P2_R1233_U90, new_P2_R1233_U91,
    new_P2_R1233_U92, new_P2_R1233_U93, new_P2_R1233_U94, new_P2_R1233_U95,
    new_P2_R1233_U96, new_P2_R1233_U97, new_P2_R1233_U98, new_P2_R1233_U99,
    new_P2_R1233_U100, new_P2_R1233_U101, new_P2_R1233_U102,
    new_P2_R1233_U103, new_P2_R1233_U104, new_P2_R1233_U105,
    new_P2_R1233_U106, new_P2_R1233_U107, new_P2_R1233_U108,
    new_P2_R1233_U109, new_P2_R1233_U110, new_P2_R1233_U111,
    new_P2_R1233_U112, new_P2_R1233_U113, new_P2_R1233_U114,
    new_P2_R1233_U115, new_P2_R1233_U116, new_P2_R1233_U117,
    new_P2_R1233_U118, new_P2_R1233_U119, new_P2_R1233_U120,
    new_P2_R1233_U121, new_P2_R1233_U122, new_P2_R1233_U123,
    new_P2_R1233_U124, new_P2_R1233_U125, new_P2_R1233_U126,
    new_P2_R1233_U127, new_P2_R1233_U128, new_P2_R1233_U129,
    new_P2_R1233_U130, new_P2_R1233_U131, new_P2_R1233_U132,
    new_P2_R1233_U133, new_P2_R1233_U134, new_P2_R1233_U135,
    new_P2_R1233_U136, new_P2_R1233_U137, new_P2_R1233_U138,
    new_P2_R1233_U139, new_P2_R1233_U140, new_P2_R1233_U141,
    new_P2_R1233_U142, new_P2_R1233_U143, new_P2_R1233_U144,
    new_P2_R1233_U145, new_P2_R1233_U146, new_P2_R1233_U147,
    new_P2_R1233_U148, new_P2_R1233_U149, new_P2_R1233_U150,
    new_P2_R1233_U151, new_P2_R1233_U152, new_P2_R1233_U153,
    new_P2_R1233_U154, new_P2_R1233_U155, new_P2_R1233_U156,
    new_P2_R1233_U157, new_P2_R1233_U158, new_P2_R1233_U159,
    new_P2_R1233_U160, new_P2_R1233_U161, new_P2_R1233_U162,
    new_P2_R1233_U163, new_P2_R1233_U164, new_P2_R1233_U165,
    new_P2_R1233_U166, new_P2_R1233_U167, new_P2_R1233_U168,
    new_P2_R1233_U169, new_P2_R1233_U170, new_P2_R1233_U171,
    new_P2_R1233_U172, new_P2_R1233_U173, new_P2_R1233_U174,
    new_P2_R1233_U175, new_P2_R1233_U176, new_P2_R1233_U177,
    new_P2_R1233_U178, new_P2_R1233_U179, new_P2_R1233_U180,
    new_P2_R1233_U181, new_P2_R1233_U182, new_P2_R1233_U183,
    new_P2_R1233_U184, new_P2_R1233_U185, new_P2_R1233_U186,
    new_P2_R1233_U187, new_P2_R1233_U188, new_P2_R1233_U189,
    new_P2_R1233_U190, new_P2_R1233_U191, new_P2_R1233_U192,
    new_P2_R1233_U193, new_P2_R1233_U194, new_P2_R1233_U195,
    new_P2_R1233_U196, new_P2_R1233_U197, new_P2_R1233_U198,
    new_P2_R1233_U199, new_P2_R1233_U200, new_P2_R1233_U201,
    new_P2_R1233_U202, new_P2_R1233_U203, new_P2_R1233_U204,
    new_P2_R1233_U205, new_P2_R1233_U206, new_P2_R1233_U207,
    new_P2_R1233_U208, new_P2_R1233_U209, new_P2_R1233_U210,
    new_P2_R1233_U211, new_P2_R1233_U212, new_P2_R1233_U213,
    new_P2_R1233_U214, new_P2_R1233_U215, new_P2_R1233_U216,
    new_P2_R1233_U217, new_P2_R1233_U218, new_P2_R1233_U219,
    new_P2_R1233_U220, new_P2_R1233_U221, new_P2_R1233_U222,
    new_P2_R1233_U223, new_P2_R1233_U224, new_P2_R1233_U225,
    new_P2_R1233_U226, new_P2_R1233_U227, new_P2_R1233_U228,
    new_P2_R1233_U229, new_P2_R1233_U230, new_P2_R1233_U231,
    new_P2_R1233_U232, new_P2_R1233_U233, new_P2_R1233_U234,
    new_P2_R1233_U235, new_P2_R1233_U236, new_P2_R1233_U237,
    new_P2_R1233_U238, new_P2_R1233_U239, new_P2_R1233_U240,
    new_P2_R1233_U241, new_P2_R1233_U242, new_P2_R1233_U243,
    new_P2_R1233_U244, new_P2_R1233_U245, new_P2_R1233_U246,
    new_P2_R1233_U247, new_P2_R1233_U248, new_P2_R1233_U249,
    new_P2_R1233_U250, new_P2_R1233_U251, new_P2_R1233_U252,
    new_P2_R1233_U253, new_P2_R1233_U254, new_P2_R1233_U255,
    new_P2_R1233_U256, new_P2_R1233_U257, new_P2_R1233_U258,
    new_P2_R1233_U259, new_P2_R1233_U260, new_P2_R1233_U261,
    new_P2_R1233_U262, new_P2_R1233_U263, new_P2_R1233_U264,
    new_P2_R1233_U265, new_P2_R1233_U266, new_P2_R1233_U267,
    new_P2_R1233_U268, new_P2_R1233_U269, new_P2_R1233_U270,
    new_P2_R1233_U271, new_P2_R1233_U272, new_P2_R1233_U273,
    new_P2_R1233_U274, new_P2_R1233_U275, new_P2_R1233_U276,
    new_P2_R1233_U277, new_P2_R1233_U278, new_P2_R1233_U279,
    new_P2_R1233_U280, new_P2_R1233_U281, new_P2_R1233_U282,
    new_P2_R1233_U283, new_P2_R1233_U284, new_P2_R1233_U285,
    new_P2_R1233_U286, new_P2_R1233_U287, new_P2_R1233_U288,
    new_P2_R1233_U289, new_P2_R1233_U290, new_P2_R1233_U291,
    new_P2_R1233_U292, new_P2_R1233_U293, new_P2_R1233_U294,
    new_P2_R1233_U295, new_P2_R1233_U296, new_P2_R1233_U297,
    new_P2_R1233_U298, new_P2_R1233_U299, new_P2_R1233_U300,
    new_P2_R1233_U301, new_P2_R1233_U302, new_P2_R1233_U303,
    new_P2_R1233_U304, new_P2_R1233_U305, new_P2_R1233_U306,
    new_P2_R1233_U307, new_P2_R1233_U308, new_P2_R1233_U309,
    new_P2_R1233_U310, new_P2_R1233_U311, new_P2_R1233_U312,
    new_P2_R1233_U313, new_P2_R1233_U314, new_P2_R1233_U315,
    new_P2_R1233_U316, new_P2_R1233_U317, new_P2_R1233_U318,
    new_P2_R1233_U319, new_P2_R1233_U320, new_P2_R1233_U321,
    new_P2_R1233_U322, new_P2_R1233_U323, new_P2_R1233_U324,
    new_P2_R1233_U325, new_P2_R1233_U326, new_P2_R1233_U327,
    new_P2_R1233_U328, new_P2_R1233_U329, new_P2_R1233_U330,
    new_P2_R1233_U331, new_P2_R1233_U332, new_P2_R1233_U333,
    new_P2_R1233_U334, new_P2_R1233_U335, new_P2_R1233_U336,
    new_P2_R1233_U337, new_P2_R1233_U338, new_P2_R1233_U339,
    new_P2_R1233_U340, new_P2_R1233_U341, new_P2_R1233_U342,
    new_P2_R1233_U343, new_P2_R1233_U344, new_P2_R1233_U345,
    new_P2_R1233_U346, new_P2_R1233_U347, new_P2_R1233_U348,
    new_P2_R1233_U349, new_P2_R1233_U350, new_P2_R1233_U351,
    new_P2_R1233_U352, new_P2_R1233_U353, new_P2_R1233_U354,
    new_P2_R1233_U355, new_P2_R1233_U356, new_P2_R1233_U357,
    new_P2_R1233_U358, new_P2_R1233_U359, new_P2_R1233_U360,
    new_P2_R1233_U361, new_P2_R1233_U362, new_P2_R1233_U363,
    new_P2_R1233_U364, new_P2_R1233_U365, new_P2_R1233_U366,
    new_P2_R1233_U367, new_P2_R1233_U368, new_P2_R1233_U369,
    new_P2_R1233_U370, new_P2_R1233_U371, new_P2_R1233_U372,
    new_P2_R1233_U373, new_P2_R1233_U374, new_P2_R1233_U375,
    new_P2_R1233_U376, new_P2_R1233_U377, new_P2_R1233_U378,
    new_P2_R1233_U379, new_P2_R1233_U380, new_P2_R1233_U381,
    new_P2_R1233_U382, new_P2_R1233_U383, new_P2_R1233_U384,
    new_P2_R1233_U385, new_P2_R1233_U386, new_P2_R1233_U387,
    new_P2_R1233_U388, new_P2_R1233_U389, new_P2_R1233_U390,
    new_P2_R1233_U391, new_P2_R1233_U392, new_P2_R1233_U393,
    new_P2_R1233_U394, new_P2_R1233_U395, new_P2_R1233_U396,
    new_P2_R1233_U397, new_P2_R1233_U398, new_P2_R1233_U399,
    new_P2_R1233_U400, new_P2_R1233_U401, new_P2_R1233_U402,
    new_P2_R1233_U403, new_P2_R1233_U404, new_P2_R1233_U405,
    new_P2_R1233_U406, new_P2_R1233_U407, new_P2_R1233_U408,
    new_P2_R1233_U409, new_P2_R1233_U410, new_P2_R1233_U411,
    new_P2_R1233_U412, new_P2_R1233_U413, new_P2_R1233_U414,
    new_P2_R1233_U415, new_P2_R1233_U416, new_P2_R1233_U417,
    new_P2_R1233_U418, new_P2_R1233_U419, new_P2_R1233_U420,
    new_P2_R1233_U421, new_P2_R1233_U422, new_P2_R1233_U423,
    new_P2_R1233_U424, new_P2_R1233_U425, new_P2_R1233_U426,
    new_P2_R1233_U427, new_P2_R1233_U428, new_P2_R1233_U429,
    new_P2_R1233_U430, new_P2_R1233_U431, new_P2_R1233_U432,
    new_P2_R1233_U433, new_P2_R1233_U434, new_P2_R1233_U435,
    new_P2_R1233_U436, new_P2_R1233_U437, new_P2_R1233_U438,
    new_P2_R1233_U439, new_P2_R1233_U440, new_P2_R1233_U441,
    new_P2_R1233_U442, new_P2_R1233_U443, new_P2_R1233_U444,
    new_P2_R1233_U445, new_P2_R1233_U446, new_P2_R1233_U447,
    new_P2_R1233_U448, new_P2_R1233_U449, new_P2_R1233_U450,
    new_P2_R1233_U451, new_P2_R1233_U452, new_P2_R1233_U453,
    new_P2_R1233_U454, new_P2_R1233_U455, new_P2_R1233_U456,
    new_P2_R1233_U457, new_P2_R1233_U458, new_P2_R1233_U459,
    new_P2_R1233_U460, new_P2_R1233_U461, new_P2_R1233_U462,
    new_P2_R1233_U463, new_P2_R1233_U464, new_P2_R1233_U465,
    new_P2_R1233_U466, new_P2_R1233_U467, new_P2_R1233_U468,
    new_P2_R1233_U469, new_P2_R1233_U470, new_P2_R1233_U471,
    new_P2_R1233_U472, new_P2_R1233_U473, new_P2_R1233_U474,
    new_P2_R1233_U475, new_P2_R1233_U476, new_P2_R1233_U477,
    new_P2_R1233_U478, new_P2_R1233_U479, new_P2_R1233_U480,
    new_P2_R1233_U481, new_P2_R1233_U482, new_P2_R1233_U483,
    new_P2_R1233_U484, new_P2_R1233_U485, new_P2_R1233_U486,
    new_P2_R1233_U487, new_P2_R1233_U488, new_P2_R1233_U489,
    new_P2_R1233_U490, new_P2_R1233_U491, new_P2_R1233_U492,
    new_P2_R1233_U493, new_P2_R1233_U494, new_P2_R1233_U495,
    new_P2_R1233_U496, new_P2_R1233_U497, new_P2_R1233_U498,
    new_P2_R1233_U499, new_P2_R1233_U500, new_P2_R1233_U501,
    new_P2_R1233_U502, new_P2_R1233_U503, new_P2_R1233_U504,
    new_P2_R1176_U4, new_P2_R1176_U5, new_P2_R1176_U6, new_P2_R1176_U7,
    new_P2_R1176_U8, new_P2_R1176_U9, new_P2_R1176_U10, new_P2_R1176_U11,
    new_P2_R1176_U12, new_P2_R1176_U13, new_P2_R1176_U14, new_P2_R1176_U15,
    new_P2_R1176_U16, new_P2_R1176_U17, new_P2_R1176_U18, new_P2_R1176_U19,
    new_P2_R1176_U20, new_P2_R1176_U21, new_P2_R1176_U22, new_P2_R1176_U23,
    new_P2_R1176_U24, new_P2_R1176_U25, new_P2_R1176_U26, new_P2_R1176_U27,
    new_P2_R1176_U28, new_P2_R1176_U29, new_P2_R1176_U30, new_P2_R1176_U31,
    new_P2_R1176_U32, new_P2_R1176_U33, new_P2_R1176_U34, new_P2_R1176_U35,
    new_P2_R1176_U36, new_P2_R1176_U37, new_P2_R1176_U38, new_P2_R1176_U39,
    new_P2_R1176_U40, new_P2_R1176_U41, new_P2_R1176_U42, new_P2_R1176_U43,
    new_P2_R1176_U44, new_P2_R1176_U45, new_P2_R1176_U46, new_P2_R1176_U47,
    new_P2_R1176_U48, new_P2_R1176_U49, new_P2_R1176_U50, new_P2_R1176_U51,
    new_P2_R1176_U52, new_P2_R1176_U53, new_P2_R1176_U54, new_P2_R1176_U55,
    new_P2_R1176_U56, new_P2_R1176_U57, new_P2_R1176_U58, new_P2_R1176_U59,
    new_P2_R1176_U60, new_P2_R1176_U61, new_P2_R1176_U62, new_P2_R1176_U63,
    new_P2_R1176_U64, new_P2_R1176_U65, new_P2_R1176_U66, new_P2_R1176_U67,
    new_P2_R1176_U68, new_P2_R1176_U69, new_P2_R1176_U70, new_P2_R1176_U71,
    new_P2_R1176_U72, new_P2_R1176_U73, new_P2_R1176_U74, new_P2_R1176_U75,
    new_P2_R1176_U76, new_P2_R1176_U77, new_P2_R1176_U78, new_P2_R1176_U79,
    new_P2_R1176_U80, new_P2_R1176_U81, new_P2_R1176_U82, new_P2_R1176_U83,
    new_P2_R1176_U84, new_P2_R1176_U85, new_P2_R1176_U86, new_P2_R1176_U87,
    new_P2_R1176_U88, new_P2_R1176_U89, new_P2_R1176_U90, new_P2_R1176_U91,
    new_P2_R1176_U92, new_P2_R1176_U93, new_P2_R1176_U94, new_P2_R1176_U95,
    new_P2_R1176_U96, new_P2_R1176_U97, new_P2_R1176_U98, new_P2_R1176_U99,
    new_P2_R1176_U100, new_P2_R1176_U101, new_P2_R1176_U102,
    new_P2_R1176_U103, new_P2_R1176_U104, new_P2_R1176_U105,
    new_P2_R1176_U106, new_P2_R1176_U107, new_P2_R1176_U108,
    new_P2_R1176_U109, new_P2_R1176_U110, new_P2_R1176_U111,
    new_P2_R1176_U112, new_P2_R1176_U113, new_P2_R1176_U114,
    new_P2_R1176_U115, new_P2_R1176_U116, new_P2_R1176_U117,
    new_P2_R1176_U118, new_P2_R1176_U119, new_P2_R1176_U120,
    new_P2_R1176_U121, new_P2_R1176_U122, new_P2_R1176_U123,
    new_P2_R1176_U124, new_P2_R1176_U125, new_P2_R1176_U126,
    new_P2_R1176_U127, new_P2_R1176_U128, new_P2_R1176_U129,
    new_P2_R1176_U130, new_P2_R1176_U131, new_P2_R1176_U132,
    new_P2_R1176_U133, new_P2_R1176_U134, new_P2_R1176_U135,
    new_P2_R1176_U136, new_P2_R1176_U137, new_P2_R1176_U138,
    new_P2_R1176_U139, new_P2_R1176_U140, new_P2_R1176_U141,
    new_P2_R1176_U142, new_P2_R1176_U143, new_P2_R1176_U144,
    new_P2_R1176_U145, new_P2_R1176_U146, new_P2_R1176_U147,
    new_P2_R1176_U148, new_P2_R1176_U149, new_P2_R1176_U150,
    new_P2_R1176_U151, new_P2_R1176_U152, new_P2_R1176_U153,
    new_P2_R1176_U154, new_P2_R1176_U155, new_P2_R1176_U156,
    new_P2_R1176_U157, new_P2_R1176_U158, new_P2_R1176_U159,
    new_P2_R1176_U160, new_P2_R1176_U161, new_P2_R1176_U162,
    new_P2_R1176_U163, new_P2_R1176_U164, new_P2_R1176_U165,
    new_P2_R1176_U166, new_P2_R1176_U167, new_P2_R1176_U168,
    new_P2_R1176_U169, new_P2_R1176_U170, new_P2_R1176_U171,
    new_P2_R1176_U172, new_P2_R1176_U173, new_P2_R1176_U174,
    new_P2_R1176_U175, new_P2_R1176_U176, new_P2_R1176_U177,
    new_P2_R1176_U178, new_P2_R1176_U179, new_P2_R1176_U180,
    new_P2_R1176_U181, new_P2_R1176_U182, new_P2_R1176_U183,
    new_P2_R1176_U184, new_P2_R1176_U185, new_P2_R1176_U186,
    new_P2_R1176_U187, new_P2_R1176_U188, new_P2_R1176_U189,
    new_P2_R1176_U190, new_P2_R1176_U191, new_P2_R1176_U192,
    new_P2_R1176_U193, new_P2_R1176_U194, new_P2_R1176_U195,
    new_P2_R1176_U196, new_P2_R1176_U197, new_P2_R1176_U198,
    new_P2_R1176_U199, new_P2_R1176_U200, new_P2_R1176_U201,
    new_P2_R1176_U202, new_P2_R1176_U203, new_P2_R1176_U204,
    new_P2_R1176_U205, new_P2_R1176_U206, new_P2_R1176_U207,
    new_P2_R1176_U208, new_P2_R1176_U209, new_P2_R1176_U210,
    new_P2_R1176_U211, new_P2_R1176_U212, new_P2_R1176_U213,
    new_P2_R1176_U214, new_P2_R1176_U215, new_P2_R1176_U216,
    new_P2_R1176_U217, new_P2_R1176_U218, new_P2_R1176_U219,
    new_P2_R1176_U220, new_P2_R1176_U221, new_P2_R1176_U222,
    new_P2_R1176_U223, new_P2_R1176_U224, new_P2_R1176_U225,
    new_P2_R1176_U226, new_P2_R1176_U227, new_P2_R1176_U228,
    new_P2_R1176_U229, new_P2_R1176_U230, new_P2_R1176_U231,
    new_P2_R1176_U232, new_P2_R1176_U233, new_P2_R1176_U234,
    new_P2_R1176_U235, new_P2_R1176_U236, new_P2_R1176_U237,
    new_P2_R1176_U238, new_P2_R1176_U239, new_P2_R1176_U240,
    new_P2_R1176_U241, new_P2_R1176_U242, new_P2_R1176_U243,
    new_P2_R1176_U244, new_P2_R1176_U245, new_P2_R1176_U246,
    new_P2_R1176_U247, new_P2_R1176_U248, new_P2_R1176_U249,
    new_P2_R1176_U250, new_P2_R1176_U251, new_P2_R1176_U252,
    new_P2_R1176_U253, new_P2_R1176_U254, new_P2_R1176_U255,
    new_P2_R1176_U256, new_P2_R1176_U257, new_P2_R1176_U258,
    new_P2_R1176_U259, new_P2_R1176_U260, new_P2_R1176_U261,
    new_P2_R1176_U262, new_P2_R1176_U263, new_P2_R1176_U264,
    new_P2_R1176_U265, new_P2_R1176_U266, new_P2_R1176_U267,
    new_P2_R1176_U268, new_P2_R1176_U269, new_P2_R1176_U270,
    new_P2_R1176_U271, new_P2_R1176_U272, new_P2_R1176_U273,
    new_P2_R1176_U274, new_P2_R1176_U275, new_P2_R1176_U276,
    new_P2_R1176_U277, new_P2_R1176_U278, new_P2_R1176_U279,
    new_P2_R1176_U280, new_P2_R1176_U281, new_P2_R1176_U282,
    new_P2_R1176_U283, new_P2_R1176_U284, new_P2_R1176_U285,
    new_P2_R1176_U286, new_P2_R1176_U287, new_P2_R1176_U288,
    new_P2_R1176_U289, new_P2_R1176_U290, new_P2_R1176_U291,
    new_P2_R1176_U292, new_P2_R1176_U293, new_P2_R1176_U294,
    new_P2_R1176_U295, new_P2_R1176_U296, new_P2_R1176_U297,
    new_P2_R1176_U298, new_P2_R1176_U299, new_P2_R1176_U300,
    new_P2_R1176_U301, new_P2_R1176_U302, new_P2_R1176_U303,
    new_P2_R1176_U304, new_P2_R1176_U305, new_P2_R1176_U306,
    new_P2_R1176_U307, new_P2_R1176_U308, new_P2_R1176_U309,
    new_P2_R1176_U310, new_P2_R1176_U311, new_P2_R1176_U312,
    new_P2_R1176_U313, new_P2_R1176_U314, new_P2_R1176_U315,
    new_P2_R1176_U316, new_P2_R1176_U317, new_P2_R1176_U318,
    new_P2_R1176_U319, new_P2_R1176_U320, new_P2_R1176_U321,
    new_P2_R1176_U322, new_P2_R1176_U323, new_P2_R1176_U324,
    new_P2_R1176_U325, new_P2_R1176_U326, new_P2_R1176_U327,
    new_P2_R1176_U328, new_P2_R1176_U329, new_P2_R1176_U330,
    new_P2_R1176_U331, new_P2_R1176_U332, new_P2_R1176_U333,
    new_P2_R1176_U334, new_P2_R1176_U335, new_P2_R1176_U336,
    new_P2_R1176_U337, new_P2_R1176_U338, new_P2_R1176_U339,
    new_P2_R1176_U340, new_P2_R1176_U341, new_P2_R1176_U342,
    new_P2_R1176_U343, new_P2_R1176_U344, new_P2_R1176_U345,
    new_P2_R1176_U346, new_P2_R1176_U347, new_P2_R1176_U348,
    new_P2_R1176_U349, new_P2_R1176_U350, new_P2_R1176_U351,
    new_P2_R1176_U352, new_P2_R1176_U353, new_P2_R1176_U354,
    new_P2_R1176_U355, new_P2_R1176_U356, new_P2_R1176_U357,
    new_P2_R1176_U358, new_P2_R1176_U359, new_P2_R1176_U360,
    new_P2_R1176_U361, new_P2_R1176_U362, new_P2_R1176_U363,
    new_P2_R1176_U364, new_P2_R1176_U365, new_P2_R1176_U366,
    new_P2_R1176_U367, new_P2_R1176_U368, new_P2_R1176_U369,
    new_P2_R1176_U370, new_P2_R1176_U371, new_P2_R1176_U372,
    new_P2_R1176_U373, new_P2_R1176_U374, new_P2_R1176_U375,
    new_P2_R1176_U376, new_P2_R1176_U377, new_P2_R1176_U378,
    new_P2_R1176_U379, new_P2_R1176_U380, new_P2_R1176_U381,
    new_P2_R1176_U382, new_P2_R1176_U383, new_P2_R1176_U384,
    new_P2_R1176_U385, new_P2_R1176_U386, new_P2_R1176_U387,
    new_P2_R1176_U388, new_P2_R1176_U389, new_P2_R1176_U390,
    new_P2_R1176_U391, new_P2_R1176_U392, new_P2_R1176_U393,
    new_P2_R1176_U394, new_P2_R1176_U395, new_P2_R1176_U396,
    new_P2_R1176_U397, new_P2_R1176_U398, new_P2_R1176_U399,
    new_P2_R1176_U400, new_P2_R1176_U401, new_P2_R1176_U402,
    new_P2_R1176_U403, new_P2_R1176_U404, new_P2_R1176_U405,
    new_P2_R1176_U406, new_P2_R1176_U407, new_P2_R1176_U408,
    new_P2_R1176_U409, new_P2_R1176_U410, new_P2_R1176_U411,
    new_P2_R1176_U412, new_P2_R1176_U413, new_P2_R1176_U414,
    new_P2_R1176_U415, new_P2_R1176_U416, new_P2_R1176_U417,
    new_P2_R1176_U418, new_P2_R1176_U419, new_P2_R1176_U420,
    new_P2_R1176_U421, new_P2_R1176_U422, new_P2_R1176_U423,
    new_P2_R1176_U424, new_P2_R1176_U425, new_P2_R1176_U426,
    new_P2_R1176_U427, new_P2_R1176_U428, new_P2_R1176_U429,
    new_P2_R1176_U430, new_P2_R1176_U431, new_P2_R1176_U432,
    new_P2_R1176_U433, new_P2_R1176_U434, new_P2_R1176_U435,
    new_P2_R1176_U436, new_P2_R1176_U437, new_P2_R1176_U438,
    new_P2_R1176_U439, new_P2_R1176_U440, new_P2_R1176_U441,
    new_P2_R1176_U442, new_P2_R1176_U443, new_P2_R1176_U444,
    new_P2_R1176_U445, new_P2_R1176_U446, new_P2_R1176_U447,
    new_P2_R1176_U448, new_P2_R1176_U449, new_P2_R1176_U450,
    new_P2_R1176_U451, new_P2_R1176_U452, new_P2_R1176_U453,
    new_P2_R1176_U454, new_P2_R1176_U455, new_P2_R1176_U456,
    new_P2_R1176_U457, new_P2_R1176_U458, new_P2_R1176_U459,
    new_P2_R1176_U460, new_P2_R1176_U461, new_P2_R1176_U462,
    new_P2_R1176_U463, new_P2_R1176_U464, new_P2_R1176_U465,
    new_P2_R1176_U466, new_P2_R1176_U467, new_P2_R1176_U468,
    new_P2_R1176_U469, new_P2_R1176_U470, new_P2_R1176_U471,
    new_P2_R1176_U472, new_P2_R1176_U473, new_P2_R1176_U474,
    new_P2_R1176_U475, new_P2_R1176_U476, new_P2_R1176_U477,
    new_P2_R1176_U478, new_P2_R1176_U479, new_P2_R1176_U480,
    new_P2_R1176_U481, new_P2_R1176_U482, new_P2_R1176_U483,
    new_P2_R1176_U484, new_P2_R1176_U485, new_P2_R1176_U486,
    new_P2_R1176_U487, new_P2_R1176_U488, new_P2_R1176_U489,
    new_P2_R1176_U490, new_P2_R1176_U491, new_P2_R1176_U492,
    new_P2_R1176_U493, new_P2_R1176_U494, new_P2_R1176_U495,
    new_P2_R1176_U496, new_P2_R1176_U497, new_P2_R1176_U498,
    new_P2_R1176_U499, new_P2_R1176_U500, new_P2_R1176_U501,
    new_P2_R1176_U502, new_P2_R1176_U503, new_P2_R1176_U504,
    new_P2_R1176_U505, new_P2_R1176_U506, new_P2_R1176_U507,
    new_P2_R1176_U508, new_P2_R1176_U509, new_P2_R1176_U510,
    new_P2_R1176_U511, new_P2_R1176_U512, new_P2_R1176_U513,
    new_P2_R1176_U514, new_P2_R1176_U515, new_P2_R1176_U516,
    new_P2_R1176_U517, new_P2_R1176_U518, new_P2_R1176_U519,
    new_P2_R1176_U520, new_P2_R1176_U521, new_P2_R1176_U522,
    new_P2_R1176_U523, new_P2_R1176_U524, new_P2_R1176_U525,
    new_P2_R1176_U526, new_P2_R1176_U527, new_P2_R1176_U528,
    new_P2_R1176_U529, new_P2_R1176_U530, new_P2_R1176_U531,
    new_P2_R1176_U532, new_P2_R1176_U533, new_P2_R1176_U534,
    new_P2_R1176_U535, new_P2_R1176_U536, new_P2_R1176_U537,
    new_P2_R1176_U538, new_P2_R1176_U539, new_P2_R1176_U540,
    new_P2_R1176_U541, new_P2_R1176_U542, new_P2_R1176_U543,
    new_P2_R1176_U544, new_P2_R1176_U545, new_P2_R1176_U546,
    new_P2_R1176_U547, new_P2_R1176_U548, new_P2_R1176_U549,
    new_P2_R1176_U550, new_P2_R1176_U551, new_P2_R1176_U552,
    new_P2_R1176_U553, new_P2_R1176_U554, new_P2_R1176_U555,
    new_P2_R1176_U556, new_P2_R1176_U557, new_P2_R1176_U558,
    new_P2_R1176_U559, new_P2_R1176_U560, new_P2_R1176_U561,
    new_P2_R1176_U562, new_P2_R1176_U563, new_P2_R1176_U564,
    new_P2_R1176_U565, new_P2_R1176_U566, new_P2_R1176_U567,
    new_P2_R1176_U568, new_P2_R1176_U569, new_P2_R1176_U570,
    new_P2_R1176_U571, new_P2_R1176_U572, new_P2_R1176_U573,
    new_P2_R1176_U574, new_P2_R1176_U575, new_P2_R1176_U576,
    new_P2_R1176_U577, new_P2_R1176_U578, new_P2_R1176_U579,
    new_P2_R1176_U580, new_P2_R1176_U581, new_P2_R1176_U582,
    new_P2_R1176_U583, new_P2_R1176_U584, new_P2_R1176_U585,
    new_P2_R1176_U586, new_P2_R1176_U587, new_P2_R1176_U588,
    new_P2_R1176_U589, new_P2_R1176_U590, new_P2_R1176_U591,
    new_P2_R1176_U592, new_P2_R1176_U593, new_P2_R1176_U594,
    new_P2_R1176_U595, new_P2_R1176_U596, new_P2_R1176_U597,
    new_P2_R1176_U598, new_P2_R1176_U599, new_P2_R1176_U600,
    new_P2_R1176_U601, new_P2_R1176_U602, new_P2_R1176_U603,
    new_P2_R1176_U604, new_P2_R1176_U605, new_P2_R1176_U606,
    new_P2_R1176_U607, new_P2_R1176_U608, new_P2_R1176_U609,
    new_P2_R1176_U610, new_P2_R1176_U611, new_P2_R1176_U612,
    new_P2_R1176_U613, new_P2_R1176_U614, new_P2_R1176_U615,
    new_P2_R1176_U616, new_P2_R1176_U617, new_P2_R1176_U618,
    new_P2_R1176_U619, new_P2_R1176_U620, new_P2_R1176_U621,
    new_P2_R1176_U622, new_P2_R1176_U623, new_P2_R1131_U4, new_P2_R1131_U5,
    new_P2_R1131_U6, new_P2_R1131_U7, new_P2_R1131_U8, new_P2_R1131_U9,
    new_P2_R1131_U10, new_P2_R1131_U11, new_P2_R1131_U12, new_P2_R1131_U13,
    new_P2_R1131_U14, new_P2_R1131_U15, new_P2_R1131_U16, new_P2_R1131_U17,
    new_P2_R1131_U18, new_P2_R1131_U19, new_P2_R1131_U20, new_P2_R1131_U21,
    new_P2_R1131_U22, new_P2_R1131_U23, new_P2_R1131_U24, new_P2_R1131_U25,
    new_P2_R1131_U26, new_P2_R1131_U27, new_P2_R1131_U28, new_P2_R1131_U29,
    new_P2_R1131_U30, new_P2_R1131_U31, new_P2_R1131_U32, new_P2_R1131_U33,
    new_P2_R1131_U34, new_P2_R1131_U35, new_P2_R1131_U36, new_P2_R1131_U37,
    new_P2_R1131_U38, new_P2_R1131_U39, new_P2_R1131_U40, new_P2_R1131_U41,
    new_P2_R1131_U42, new_P2_R1131_U43, new_P2_R1131_U44, new_P2_R1131_U45,
    new_P2_R1131_U46, new_P2_R1131_U47, new_P2_R1131_U48, new_P2_R1131_U49,
    new_P2_R1131_U50, new_P2_R1131_U51, new_P2_R1131_U52, new_P2_R1131_U53,
    new_P2_R1131_U54, new_P2_R1131_U55, new_P2_R1131_U56, new_P2_R1131_U57,
    new_P2_R1131_U58, new_P2_R1131_U59, new_P2_R1131_U60, new_P2_R1131_U61,
    new_P2_R1131_U62, new_P2_R1131_U63, new_P2_R1131_U64, new_P2_R1131_U65,
    new_P2_R1131_U66, new_P2_R1131_U67, new_P2_R1131_U68, new_P2_R1131_U69,
    new_P2_R1131_U70, new_P2_R1131_U71, new_P2_R1131_U72, new_P2_R1131_U73,
    new_P2_R1131_U74, new_P2_R1131_U75, new_P2_R1131_U76, new_P2_R1131_U77,
    new_P2_R1131_U78, new_P2_R1131_U79, new_P2_R1131_U80, new_P2_R1131_U81,
    new_P2_R1131_U82, new_P2_R1131_U83, new_P2_R1131_U84, new_P2_R1131_U85,
    new_P2_R1131_U86, new_P2_R1131_U87, new_P2_R1131_U88, new_P2_R1131_U89,
    new_P2_R1131_U90, new_P2_R1131_U91, new_P2_R1131_U92, new_P2_R1131_U93,
    new_P2_R1131_U94, new_P2_R1131_U95, new_P2_R1131_U96, new_P2_R1131_U97,
    new_P2_R1131_U98, new_P2_R1131_U99, new_P2_R1131_U100,
    new_P2_R1131_U101, new_P2_R1131_U102, new_P2_R1131_U103,
    new_P2_R1131_U104, new_P2_R1131_U105, new_P2_R1131_U106,
    new_P2_R1131_U107, new_P2_R1131_U108, new_P2_R1131_U109,
    new_P2_R1131_U110, new_P2_R1131_U111, new_P2_R1131_U112,
    new_P2_R1131_U113, new_P2_R1131_U114, new_P2_R1131_U115,
    new_P2_R1131_U116, new_P2_R1131_U117, new_P2_R1131_U118,
    new_P2_R1131_U119, new_P2_R1131_U120, new_P2_R1131_U121,
    new_P2_R1131_U122, new_P2_R1131_U123, new_P2_R1131_U124,
    new_P2_R1131_U125, new_P2_R1131_U126, new_P2_R1131_U127,
    new_P2_R1131_U128, new_P2_R1131_U129, new_P2_R1131_U130,
    new_P2_R1131_U131, new_P2_R1131_U132, new_P2_R1131_U133,
    new_P2_R1131_U134, new_P2_R1131_U135, new_P2_R1131_U136,
    new_P2_R1131_U137, new_P2_R1131_U138, new_P2_R1131_U139,
    new_P2_R1131_U140, new_P2_R1131_U141, new_P2_R1131_U142,
    new_P2_R1131_U143, new_P2_R1131_U144, new_P2_R1131_U145,
    new_P2_R1131_U146, new_P2_R1131_U147, new_P2_R1131_U148,
    new_P2_R1131_U149, new_P2_R1131_U150, new_P2_R1131_U151,
    new_P2_R1131_U152, new_P2_R1131_U153, new_P2_R1131_U154,
    new_P2_R1131_U155, new_P2_R1131_U156, new_P2_R1131_U157,
    new_P2_R1131_U158, new_P2_R1131_U159, new_P2_R1131_U160,
    new_P2_R1131_U161, new_P2_R1131_U162, new_P2_R1131_U163,
    new_P2_R1131_U164, new_P2_R1131_U165, new_P2_R1131_U166,
    new_P2_R1131_U167, new_P2_R1131_U168, new_P2_R1131_U169,
    new_P2_R1131_U170, new_P2_R1131_U171, new_P2_R1131_U172,
    new_P2_R1131_U173, new_P2_R1131_U174, new_P2_R1131_U175,
    new_P2_R1131_U176, new_P2_R1131_U177, new_P2_R1131_U178,
    new_P2_R1131_U179, new_P2_R1131_U180, new_P2_R1131_U181,
    new_P2_R1131_U182, new_P2_R1131_U183, new_P2_R1131_U184,
    new_P2_R1131_U185, new_P2_R1131_U186, new_P2_R1131_U187,
    new_P2_R1131_U188, new_P2_R1131_U189, new_P2_R1131_U190,
    new_P2_R1131_U191, new_P2_R1131_U192, new_P2_R1131_U193,
    new_P2_R1131_U194, new_P2_R1131_U195, new_P2_R1131_U196,
    new_P2_R1131_U197, new_P2_R1131_U198, new_P2_R1131_U199,
    new_P2_R1131_U200, new_P2_R1131_U201, new_P2_R1131_U202,
    new_P2_R1131_U203, new_P2_R1131_U204, new_P2_R1131_U205,
    new_P2_R1131_U206, new_P2_R1131_U207, new_P2_R1131_U208,
    new_P2_R1131_U209, new_P2_R1131_U210, new_P2_R1131_U211,
    new_P2_R1131_U212, new_P2_R1131_U213, new_P2_R1131_U214,
    new_P2_R1131_U215, new_P2_R1131_U216, new_P2_R1131_U217,
    new_P2_R1131_U218, new_P2_R1131_U219, new_P2_R1131_U220,
    new_P2_R1131_U221, new_P2_R1131_U222, new_P2_R1131_U223,
    new_P2_R1131_U224, new_P2_R1131_U225, new_P2_R1131_U226,
    new_P2_R1131_U227, new_P2_R1131_U228, new_P2_R1131_U229,
    new_P2_R1131_U230, new_P2_R1131_U231, new_P2_R1131_U232,
    new_P2_R1131_U233, new_P2_R1131_U234, new_P2_R1131_U235,
    new_P2_R1131_U236, new_P2_R1131_U237, new_P2_R1131_U238,
    new_P2_R1131_U239, new_P2_R1131_U240, new_P2_R1131_U241,
    new_P2_R1131_U242, new_P2_R1131_U243, new_P2_R1131_U244,
    new_P2_R1131_U245, new_P2_R1131_U246, new_P2_R1131_U247,
    new_P2_R1131_U248, new_P2_R1131_U249, new_P2_R1131_U250,
    new_P2_R1131_U251, new_P2_R1131_U252, new_P2_R1131_U253,
    new_P2_R1131_U254, new_P2_R1131_U255, new_P2_R1131_U256,
    new_P2_R1131_U257, new_P2_R1131_U258, new_P2_R1131_U259,
    new_P2_R1131_U260, new_P2_R1131_U261, new_P2_R1131_U262,
    new_P2_R1131_U263, new_P2_R1131_U264, new_P2_R1131_U265,
    new_P2_R1131_U266, new_P2_R1131_U267, new_P2_R1131_U268,
    new_P2_R1131_U269, new_P2_R1131_U270, new_P2_R1131_U271,
    new_P2_R1131_U272, new_P2_R1131_U273, new_P2_R1131_U274,
    new_P2_R1131_U275, new_P2_R1131_U276, new_P2_R1131_U277,
    new_P2_R1131_U278, new_P2_R1131_U279, new_P2_R1131_U280,
    new_P2_R1131_U281, new_P2_R1131_U282, new_P2_R1131_U283,
    new_P2_R1131_U284, new_P2_R1131_U285, new_P2_R1131_U286,
    new_P2_R1131_U287, new_P2_R1131_U288, new_P2_R1131_U289,
    new_P2_R1131_U290, new_P2_R1131_U291, new_P2_R1131_U292,
    new_P2_R1131_U293, new_P2_R1131_U294, new_P2_R1131_U295,
    new_P2_R1131_U296, new_P2_R1131_U297, new_P2_R1131_U298,
    new_P2_R1131_U299, new_P2_R1131_U300, new_P2_R1131_U301,
    new_P2_R1131_U302, new_P2_R1131_U303, new_P2_R1131_U304,
    new_P2_R1131_U305, new_P2_R1131_U306, new_P2_R1131_U307,
    new_P2_R1131_U308, new_P2_R1131_U309, new_P2_R1131_U310,
    new_P2_R1131_U311, new_P2_R1131_U312, new_P2_R1131_U313,
    new_P2_R1131_U314, new_P2_R1131_U315, new_P2_R1131_U316,
    new_P2_R1131_U317, new_P2_R1131_U318, new_P2_R1131_U319,
    new_P2_R1131_U320, new_P2_R1131_U321, new_P2_R1131_U322,
    new_P2_R1131_U323, new_P2_R1131_U324, new_P2_R1131_U325,
    new_P2_R1131_U326, new_P2_R1131_U327, new_P2_R1131_U328,
    new_P2_R1131_U329, new_P2_R1131_U330, new_P2_R1131_U331,
    new_P2_R1131_U332, new_P2_R1131_U333, new_P2_R1131_U334,
    new_P2_R1131_U335, new_P2_R1131_U336, new_P2_R1131_U337,
    new_P2_R1131_U338, new_P2_R1131_U339, new_P2_R1131_U340,
    new_P2_R1131_U341, new_P2_R1131_U342, new_P2_R1131_U343,
    new_P2_R1131_U344, new_P2_R1131_U345, new_P2_R1131_U346,
    new_P2_R1131_U347, new_P2_R1131_U348, new_P2_R1131_U349,
    new_P2_R1131_U350, new_P2_R1131_U351, new_P2_R1131_U352,
    new_P2_R1131_U353, new_P2_R1131_U354, new_P2_R1131_U355,
    new_P2_R1131_U356, new_P2_R1131_U357, new_P2_R1131_U358,
    new_P2_R1131_U359, new_P2_R1131_U360, new_P2_R1131_U361,
    new_P2_R1131_U362, new_P2_R1131_U363, new_P2_R1131_U364,
    new_P2_R1131_U365, new_P2_R1131_U366, new_P2_R1131_U367,
    new_P2_R1131_U368, new_P2_R1131_U369, new_P2_R1131_U370,
    new_P2_R1131_U371, new_P2_R1131_U372, new_P2_R1131_U373,
    new_P2_R1131_U374, new_P2_R1131_U375, new_P2_R1131_U376,
    new_P2_R1131_U377, new_P2_R1131_U378, new_P2_R1131_U379,
    new_P2_R1131_U380, new_P2_R1131_U381, new_P2_R1131_U382,
    new_P2_R1131_U383, new_P2_R1131_U384, new_P2_R1131_U385,
    new_P2_R1131_U386, new_P2_R1131_U387, new_P2_R1131_U388,
    new_P2_R1131_U389, new_P2_R1131_U390, new_P2_R1131_U391,
    new_P2_R1131_U392, new_P2_R1131_U393, new_P2_R1131_U394,
    new_P2_R1131_U395, new_P2_R1131_U396, new_P2_R1131_U397,
    new_P2_R1131_U398, new_P2_R1131_U399, new_P2_R1131_U400,
    new_P2_R1131_U401, new_P2_R1131_U402, new_P2_R1131_U403,
    new_P2_R1131_U404, new_P2_R1131_U405, new_P2_R1131_U406,
    new_P2_R1131_U407, new_P2_R1131_U408, new_P2_R1131_U409,
    new_P2_R1131_U410, new_P2_R1131_U411, new_P2_R1131_U412,
    new_P2_R1131_U413, new_P2_R1131_U414, new_P2_R1131_U415,
    new_P2_R1131_U416, new_P2_R1131_U417, new_P2_R1131_U418,
    new_P2_R1131_U419, new_P2_R1131_U420, new_P2_R1131_U421,
    new_P2_R1131_U422, new_P2_R1131_U423, new_P2_R1131_U424,
    new_P2_R1131_U425, new_P2_R1131_U426, new_P2_R1131_U427,
    new_P2_R1131_U428, new_P2_R1131_U429, new_P2_R1131_U430,
    new_P2_R1131_U431, new_P2_R1131_U432, new_P2_R1131_U433,
    new_P2_R1131_U434, new_P2_R1131_U435, new_P2_R1131_U436,
    new_P2_R1131_U437, new_P2_R1131_U438, new_P2_R1131_U439,
    new_P2_R1131_U440, new_P2_R1131_U441, new_P2_R1131_U442,
    new_P2_R1131_U443, new_P2_R1131_U444, new_P2_R1131_U445,
    new_P2_R1131_U446, new_P2_R1131_U447, new_P2_R1131_U448,
    new_P2_R1131_U449, new_P2_R1131_U450, new_P2_R1131_U451,
    new_P2_R1131_U452, new_P2_R1131_U453, new_P2_R1131_U454,
    new_P2_R1131_U455, new_P2_R1131_U456, new_P2_R1131_U457,
    new_P2_R1131_U458, new_P2_R1131_U459, new_P2_R1131_U460,
    new_P2_R1131_U461, new_P2_R1131_U462, new_P2_R1131_U463,
    new_P2_R1131_U464, new_P2_R1131_U465, new_P2_R1131_U466,
    new_P2_R1131_U467, new_P2_R1131_U468, new_P2_R1131_U469,
    new_P2_R1131_U470, new_P2_R1131_U471, new_P2_R1131_U472,
    new_P2_R1131_U473, new_P2_R1131_U474, new_P2_R1131_U475,
    new_P2_R1131_U476, new_P2_R1131_U477, new_P2_R1131_U478,
    new_P2_R1131_U479, new_P2_R1131_U480, new_P2_R1131_U481,
    new_P2_R1131_U482, new_P2_R1131_U483, new_P2_R1131_U484,
    new_P2_R1131_U485, new_P2_R1131_U486, new_P2_R1131_U487,
    new_P2_R1131_U488, new_P2_R1131_U489, new_P2_R1131_U490,
    new_P2_R1131_U491, new_P2_R1131_U492, new_P2_R1131_U493,
    new_P2_R1131_U494, new_P2_R1131_U495, new_P2_R1131_U496,
    new_P2_R1131_U497, new_P2_R1131_U498, new_P2_R1131_U499,
    new_P2_R1131_U500, new_P2_R1131_U501, new_P2_R1131_U502,
    new_P2_R1131_U503, new_P2_R1131_U504, new_P2_R1146_U6, new_P2_R1146_U7,
    new_P2_R1146_U8, new_P2_R1146_U9, new_P2_R1146_U10, new_P2_R1146_U11,
    new_P2_R1146_U12, new_P2_R1146_U13, new_P2_R1146_U14, new_P2_R1146_U15,
    new_P2_R1146_U16, new_P2_R1146_U17, new_P2_R1146_U18, new_P2_R1146_U19,
    new_P2_R1146_U20, new_P2_R1146_U21, new_P2_R1146_U22, new_P2_R1146_U23,
    new_P2_R1146_U24, new_P2_R1146_U25, new_P2_R1146_U26, new_P2_R1146_U27,
    new_P2_R1146_U28, new_P2_R1146_U29, new_P2_R1146_U30, new_P2_R1146_U31,
    new_P2_R1146_U32, new_P2_R1146_U33, new_P2_R1146_U34, new_P2_R1146_U35,
    new_P2_R1146_U36, new_P2_R1146_U37, new_P2_R1146_U38, new_P2_R1146_U39,
    new_P2_R1146_U40, new_P2_R1146_U41, new_P2_R1146_U42, new_P2_R1146_U43,
    new_P2_R1146_U44, new_P2_R1146_U45, new_P2_R1146_U46, new_P2_R1146_U47,
    new_P2_R1146_U48, new_P2_R1146_U49, new_P2_R1146_U50, new_P2_R1146_U51,
    new_P2_R1146_U52, new_P2_R1146_U53, new_P2_R1146_U54, new_P2_R1146_U55,
    new_P2_R1146_U56, new_P2_R1146_U57, new_P2_R1146_U58, new_P2_R1146_U59,
    new_P2_R1146_U60, new_P2_R1146_U61, new_P2_R1146_U62, new_P2_R1146_U63,
    new_P2_R1146_U64, new_P2_R1146_U65, new_P2_R1146_U66, new_P2_R1146_U67,
    new_P2_R1146_U68, new_P2_R1146_U69, new_P2_R1146_U70, new_P2_R1146_U71,
    new_P2_R1146_U72, new_P2_R1146_U73, new_P2_R1146_U74, new_P2_R1146_U75,
    new_P2_R1146_U76, new_P2_R1146_U77, new_P2_R1146_U78, new_P2_R1146_U79,
    new_P2_R1146_U80, new_P2_R1146_U81, new_P2_R1146_U82, new_P2_R1146_U83,
    new_P2_R1146_U84, new_P2_R1146_U85, new_P2_R1146_U86, new_P2_R1146_U87,
    new_P2_R1146_U88, new_P2_R1146_U89, new_P2_R1146_U90, new_P2_R1146_U91,
    new_P2_R1146_U92, new_P2_R1146_U93, new_P2_R1146_U94, new_P2_R1146_U95,
    new_P2_R1146_U96, new_P2_R1146_U97, new_P2_R1146_U98, new_P2_R1146_U99,
    new_P2_R1146_U100, new_P2_R1146_U101, new_P2_R1146_U102,
    new_P2_R1146_U103, new_P2_R1146_U104, new_P2_R1146_U105,
    new_P2_R1146_U106, new_P2_R1146_U107, new_P2_R1146_U108,
    new_P2_R1146_U109, new_P2_R1146_U110, new_P2_R1146_U111,
    new_P2_R1146_U112, new_P2_R1146_U113, new_P2_R1146_U114,
    new_P2_R1146_U115, new_P2_R1146_U116, new_P2_R1146_U117,
    new_P2_R1146_U118, new_P2_R1146_U119, new_P2_R1146_U120,
    new_P2_R1146_U121, new_P2_R1146_U122, new_P2_R1146_U123,
    new_P2_R1146_U124, new_P2_R1146_U125, new_P2_R1146_U126,
    new_P2_R1146_U127, new_P2_R1146_U128, new_P2_R1146_U129,
    new_P2_R1146_U130, new_P2_R1146_U131, new_P2_R1146_U132,
    new_P2_R1146_U133, new_P2_R1146_U134, new_P2_R1146_U135,
    new_P2_R1146_U136, new_P2_R1146_U137, new_P2_R1146_U138,
    new_P2_R1146_U139, new_P2_R1146_U140, new_P2_R1146_U141,
    new_P2_R1146_U142, new_P2_R1146_U143, new_P2_R1146_U144,
    new_P2_R1146_U145, new_P2_R1146_U146, new_P2_R1146_U147,
    new_P2_R1146_U148, new_P2_R1146_U149, new_P2_R1146_U150,
    new_P2_R1146_U151, new_P2_R1146_U152, new_P2_R1146_U153,
    new_P2_R1146_U154, new_P2_R1146_U155, new_P2_R1146_U156,
    new_P2_R1146_U157, new_P2_R1146_U158, new_P2_R1146_U159,
    new_P2_R1146_U160, new_P2_R1146_U161, new_P2_R1146_U162,
    new_P2_R1146_U163, new_P2_R1146_U164, new_P2_R1146_U165,
    new_P2_R1146_U166, new_P2_R1146_U167, new_P2_R1146_U168,
    new_P2_R1146_U169, new_P2_R1146_U170, new_P2_R1146_U171,
    new_P2_R1146_U172, new_P2_R1146_U173, new_P2_R1146_U174,
    new_P2_R1146_U175, new_P2_R1146_U176, new_P2_R1146_U177,
    new_P2_R1146_U178, new_P2_R1146_U179, new_P2_R1146_U180,
    new_P2_R1146_U181, new_P2_R1146_U182, new_P2_R1146_U183,
    new_P2_R1146_U184, new_P2_R1146_U185, new_P2_R1146_U186,
    new_P2_R1146_U187, new_P2_R1146_U188, new_P2_R1146_U189,
    new_P2_R1146_U190, new_P2_R1146_U191, new_P2_R1146_U192,
    new_P2_R1146_U193, new_P2_R1146_U194, new_P2_R1146_U195,
    new_P2_R1146_U196, new_P2_R1146_U197, new_P2_R1146_U198,
    new_P2_R1146_U199, new_P2_R1146_U200, new_P2_R1146_U201,
    new_P2_R1146_U202, new_P2_R1146_U203, new_P2_R1146_U204,
    new_P2_R1146_U205, new_P2_R1146_U206, new_P2_R1146_U207,
    new_P2_R1146_U208, new_P2_R1146_U209, new_P2_R1146_U210,
    new_P2_R1146_U211, new_P2_R1146_U212, new_P2_R1146_U213,
    new_P2_R1146_U214, new_P2_R1146_U215, new_P2_R1146_U216,
    new_P2_R1146_U217, new_P2_R1146_U218, new_P2_R1146_U219,
    new_P2_R1146_U220, new_P2_R1146_U221, new_P2_R1146_U222,
    new_P2_R1146_U223, new_P2_R1146_U224, new_P2_R1146_U225,
    new_P2_R1146_U226, new_P2_R1146_U227, new_P2_R1146_U228,
    new_P2_R1146_U229, new_P2_R1146_U230, new_P2_R1146_U231,
    new_P2_R1146_U232, new_P2_R1146_U233, new_P2_R1146_U234,
    new_P2_R1146_U235, new_P2_R1146_U236, new_P2_R1146_U237,
    new_P2_R1146_U238, new_P2_R1146_U239, new_P2_R1146_U240,
    new_P2_R1146_U241, new_P2_R1146_U242, new_P2_R1146_U243,
    new_P2_R1146_U244, new_P2_R1146_U245, new_P2_R1146_U246,
    new_P2_R1146_U247, new_P2_R1146_U248, new_P2_R1146_U249,
    new_P2_R1146_U250, new_P2_R1146_U251, new_P2_R1146_U252,
    new_P2_R1146_U253, new_P2_R1146_U254, new_P2_R1146_U255,
    new_P2_R1146_U256, new_P2_R1146_U257, new_P2_R1146_U258,
    new_P2_R1146_U259, new_P2_R1146_U260, new_P2_R1146_U261,
    new_P2_R1146_U262, new_P2_R1146_U263, new_P2_R1146_U264,
    new_P2_R1146_U265, new_P2_R1146_U266, new_P2_R1146_U267,
    new_P2_R1146_U268, new_P2_R1146_U269, new_P2_R1146_U270,
    new_P2_R1146_U271, new_P2_R1146_U272, new_P2_R1146_U273,
    new_P2_R1146_U274, new_P2_R1146_U275, new_P2_R1146_U276,
    new_P2_R1146_U277, new_P2_R1146_U278, new_P2_R1146_U279,
    new_P2_R1146_U280, new_P2_R1146_U281, new_P2_R1146_U282,
    new_P2_R1146_U283, new_P2_R1146_U284, new_P2_R1146_U285,
    new_P2_R1146_U286, new_P2_R1146_U287, new_P2_R1146_U288,
    new_P2_R1146_U289, new_P2_R1146_U290, new_P2_R1146_U291,
    new_P2_R1146_U292, new_P2_R1146_U293, new_P2_R1146_U294,
    new_P2_R1146_U295, new_P2_R1146_U296, new_P2_R1146_U297,
    new_P2_R1146_U298, new_P2_R1146_U299, new_P2_R1146_U300,
    new_P2_R1146_U301, new_P2_R1146_U302, new_P2_R1146_U303,
    new_P2_R1146_U304, new_P2_R1146_U305, new_P2_R1146_U306,
    new_P2_R1146_U307, new_P2_R1146_U308, new_P2_R1146_U309,
    new_P2_R1146_U310, new_P2_R1146_U311, new_P2_R1146_U312,
    new_P2_R1146_U313, new_P2_R1146_U314, new_P2_R1146_U315,
    new_P2_R1146_U316, new_P2_R1146_U317, new_P2_R1146_U318,
    new_P2_R1146_U319, new_P2_R1146_U320, new_P2_R1146_U321,
    new_P2_R1146_U322, new_P2_R1146_U323, new_P2_R1146_U324,
    new_P2_R1146_U325, new_P2_R1146_U326, new_P2_R1146_U327,
    new_P2_R1146_U328, new_P2_R1146_U329, new_P2_R1146_U330,
    new_P2_R1146_U331, new_P2_R1146_U332, new_P2_R1146_U333,
    new_P2_R1146_U334, new_P2_R1146_U335, new_P2_R1146_U336,
    new_P2_R1146_U337, new_P2_R1146_U338, new_P2_R1146_U339,
    new_P2_R1146_U340, new_P2_R1146_U341, new_P2_R1146_U342,
    new_P2_R1146_U343, new_P2_R1146_U344, new_P2_R1146_U345,
    new_P2_R1146_U346, new_P2_R1146_U347, new_P2_R1146_U348,
    new_P2_R1146_U349, new_P2_R1146_U350, new_P2_R1146_U351,
    new_P2_R1146_U352, new_P2_R1146_U353, new_P2_R1146_U354,
    new_P2_R1146_U355, new_P2_R1146_U356, new_P2_R1146_U357,
    new_P2_R1146_U358, new_P2_R1146_U359, new_P2_R1146_U360,
    new_P2_R1146_U361, new_P2_R1146_U362, new_P2_R1146_U363,
    new_P2_R1146_U364, new_P2_R1146_U365, new_P2_R1146_U366,
    new_P2_R1146_U367, new_P2_R1146_U368, new_P2_R1146_U369,
    new_P2_R1146_U370, new_P2_R1146_U371, new_P2_R1146_U372,
    new_P2_R1146_U373, new_P2_R1146_U374, new_P2_R1146_U375,
    new_P2_R1146_U376, new_P2_R1146_U377, new_P2_R1146_U378,
    new_P2_R1146_U379, new_P2_R1146_U380, new_P2_R1146_U381,
    new_P2_R1146_U382, new_P2_R1146_U383, new_P2_R1146_U384,
    new_P2_R1146_U385, new_P2_R1146_U386, new_P2_R1146_U387,
    new_P2_R1146_U388, new_P2_R1146_U389, new_P2_R1146_U390,
    new_P2_R1146_U391, new_P2_R1146_U392, new_P2_R1146_U393,
    new_P2_R1146_U394, new_P2_R1146_U395, new_P2_R1146_U396,
    new_P2_R1146_U397, new_P2_R1146_U398, new_P2_R1146_U399,
    new_P2_R1146_U400, new_P2_R1146_U401, new_P2_R1146_U402,
    new_P2_R1146_U403, new_P2_R1146_U404, new_P2_R1146_U405,
    new_P2_R1146_U406, new_P2_R1146_U407, new_P2_R1146_U408,
    new_P2_R1146_U409, new_P2_R1146_U410, new_P2_R1146_U411,
    new_P2_R1146_U412, new_P2_R1146_U413, new_P2_R1146_U414,
    new_P2_R1146_U415, new_P2_R1146_U416, new_P2_R1146_U417,
    new_P2_R1146_U418, new_P2_R1146_U419, new_P2_R1146_U420,
    new_P2_R1146_U421, new_P2_R1146_U422, new_P2_R1146_U423,
    new_P2_R1146_U424, new_P2_R1146_U425, new_P2_R1146_U426,
    new_P2_R1146_U427, new_P2_R1146_U428, new_P2_R1146_U429,
    new_P2_R1146_U430, new_P2_R1146_U431, new_P2_R1146_U432,
    new_P2_R1146_U433, new_P2_R1146_U434, new_P2_R1146_U435,
    new_P2_R1146_U436, new_P2_R1146_U437, new_P2_R1146_U438,
    new_P2_R1146_U439, new_P2_R1146_U440, new_P2_R1146_U441,
    new_P2_R1146_U442, new_P2_R1146_U443, new_P2_R1146_U444,
    new_P2_R1146_U445, new_P2_R1146_U446, new_P2_R1146_U447,
    new_P2_R1146_U448, new_P2_R1146_U449, new_P2_R1146_U450,
    new_P2_R1146_U451, new_P2_R1146_U452, new_P2_R1146_U453,
    new_P2_R1146_U454, new_P2_R1146_U455, new_P2_R1146_U456,
    new_P2_R1146_U457, new_P2_R1146_U458, new_P2_R1146_U459,
    new_P2_R1146_U460, new_P2_R1146_U461, new_P2_R1146_U462,
    new_P2_R1146_U463, new_P2_R1146_U464, new_P2_R1146_U465,
    new_P2_R1146_U466, new_P2_R1146_U467, new_P2_R1146_U468,
    new_P2_R1146_U469, new_P2_R1146_U470, new_P2_R1146_U471,
    new_P2_R1146_U472, new_P2_R1146_U473, new_P2_R1146_U474,
    new_P2_R1146_U475, new_P2_R1146_U476, new_P2_R1146_U477,
    new_P2_R1146_U478, new_P2_R1203_U6, new_P2_R1203_U7, new_P2_R1203_U8,
    new_P2_R1203_U9, new_P2_R1203_U10, new_P2_R1203_U11, new_P2_R1203_U12,
    new_P2_R1203_U13, new_P2_R1203_U14, new_P2_R1203_U15, new_P2_R1203_U16,
    new_P2_R1203_U17, new_P2_R1203_U18, new_P2_R1203_U19, new_P2_R1203_U20,
    new_P2_R1203_U21, new_P2_R1203_U22, new_P2_R1203_U23, new_P2_R1203_U24,
    new_P2_R1203_U25, new_P2_R1203_U26, new_P2_R1203_U27, new_P2_R1203_U28,
    new_P2_R1203_U29, new_P2_R1203_U30, new_P2_R1203_U31, new_P2_R1203_U32,
    new_P2_R1203_U33, new_P2_R1203_U34, new_P2_R1203_U35, new_P2_R1203_U36,
    new_P2_R1203_U37, new_P2_R1203_U38, new_P2_R1203_U39, new_P2_R1203_U40,
    new_P2_R1203_U41, new_P2_R1203_U42, new_P2_R1203_U43, new_P2_R1203_U44,
    new_P2_R1203_U45, new_P2_R1203_U46, new_P2_R1203_U47, new_P2_R1203_U48,
    new_P2_R1203_U49, new_P2_R1203_U50, new_P2_R1203_U51, new_P2_R1203_U52,
    new_P2_R1203_U53, new_P2_R1203_U54, new_P2_R1203_U55, new_P2_R1203_U56,
    new_P2_R1203_U57, new_P2_R1203_U58, new_P2_R1203_U59, new_P2_R1203_U60,
    new_P2_R1203_U61, new_P2_R1203_U62, new_P2_R1203_U63, new_P2_R1203_U64,
    new_P2_R1203_U65, new_P2_R1203_U66, new_P2_R1203_U67, new_P2_R1203_U68,
    new_P2_R1203_U69, new_P2_R1203_U70, new_P2_R1203_U71, new_P2_R1203_U72,
    new_P2_R1203_U73, new_P2_R1203_U74, new_P2_R1203_U75, new_P2_R1203_U76,
    new_P2_R1203_U77, new_P2_R1203_U78, new_P2_R1203_U79, new_P2_R1203_U80,
    new_P2_R1203_U81, new_P2_R1203_U82, new_P2_R1203_U83, new_P2_R1203_U84,
    new_P2_R1203_U85, new_P2_R1203_U86, new_P2_R1203_U87, new_P2_R1203_U88,
    new_P2_R1203_U89, new_P2_R1203_U90, new_P2_R1203_U91, new_P2_R1203_U92,
    new_P2_R1203_U93, new_P2_R1203_U94, new_P2_R1203_U95, new_P2_R1203_U96,
    new_P2_R1203_U97, new_P2_R1203_U98, new_P2_R1203_U99,
    new_P2_R1203_U100, new_P2_R1203_U101, new_P2_R1203_U102,
    new_P2_R1203_U103, new_P2_R1203_U104, new_P2_R1203_U105,
    new_P2_R1203_U106, new_P2_R1203_U107, new_P2_R1203_U108,
    new_P2_R1203_U109, new_P2_R1203_U110, new_P2_R1203_U111,
    new_P2_R1203_U112, new_P2_R1203_U113, new_P2_R1203_U114,
    new_P2_R1203_U115, new_P2_R1203_U116, new_P2_R1203_U117,
    new_P2_R1203_U118, new_P2_R1203_U119, new_P2_R1203_U120,
    new_P2_R1203_U121, new_P2_R1203_U122, new_P2_R1203_U123,
    new_P2_R1203_U124, new_P2_R1203_U125, new_P2_R1203_U126,
    new_P2_R1203_U127, new_P2_R1203_U128, new_P2_R1203_U129,
    new_P2_R1203_U130, new_P2_R1203_U131, new_P2_R1203_U132,
    new_P2_R1203_U133, new_P2_R1203_U134, new_P2_R1203_U135,
    new_P2_R1203_U136, new_P2_R1203_U137, new_P2_R1203_U138,
    new_P2_R1203_U139, new_P2_R1203_U140, new_P2_R1203_U141,
    new_P2_R1203_U142, new_P2_R1203_U143, new_P2_R1203_U144,
    new_P2_R1203_U145, new_P2_R1203_U146, new_P2_R1203_U147,
    new_P2_R1203_U148, new_P2_R1203_U149, new_P2_R1203_U150,
    new_P2_R1203_U151, new_P2_R1203_U152, new_P2_R1203_U153,
    new_P2_R1203_U154, new_P2_R1203_U155, new_P2_R1203_U156,
    new_P2_R1203_U157, new_P2_R1203_U158, new_P2_R1203_U159,
    new_P2_R1203_U160, new_P2_R1203_U161, new_P2_R1203_U162,
    new_P2_R1203_U163, new_P2_R1203_U164, new_P2_R1203_U165,
    new_P2_R1203_U166, new_P2_R1203_U167, new_P2_R1203_U168,
    new_P2_R1203_U169, new_P2_R1203_U170, new_P2_R1203_U171,
    new_P2_R1203_U172, new_P2_R1203_U173, new_P2_R1203_U174,
    new_P2_R1203_U175, new_P2_R1203_U176, new_P2_R1203_U177,
    new_P2_R1203_U178, new_P2_R1203_U179, new_P2_R1203_U180,
    new_P2_R1203_U181, new_P2_R1203_U182, new_P2_R1203_U183,
    new_P2_R1203_U184, new_P2_R1203_U185, new_P2_R1203_U186,
    new_P2_R1203_U187, new_P2_R1203_U188, new_P2_R1203_U189,
    new_P2_R1203_U190, new_P2_R1203_U191, new_P2_R1203_U192,
    new_P2_R1203_U193, new_P2_R1203_U194, new_P2_R1203_U195,
    new_P2_R1203_U196, new_P2_R1203_U197, new_P2_R1203_U198,
    new_P2_R1203_U199, new_P2_R1203_U200, new_P2_R1203_U201,
    new_P2_R1203_U202, new_P2_R1203_U203, new_P2_R1203_U204,
    new_P2_R1203_U205, new_P2_R1203_U206, new_P2_R1203_U207,
    new_P2_R1203_U208, new_P2_R1203_U209, new_P2_R1203_U210,
    new_P2_R1203_U211, new_P2_R1203_U212, new_P2_R1203_U213,
    new_P2_R1203_U214, new_P2_R1203_U215, new_P2_R1203_U216,
    new_P2_R1203_U217, new_P2_R1203_U218, new_P2_R1203_U219,
    new_P2_R1203_U220, new_P2_R1203_U221, new_P2_R1203_U222,
    new_P2_R1203_U223, new_P2_R1203_U224, new_P2_R1203_U225,
    new_P2_R1203_U226, new_P2_R1203_U227, new_P2_R1203_U228,
    new_P2_R1203_U229, new_P2_R1203_U230, new_P2_R1203_U231,
    new_P2_R1203_U232, new_P2_R1203_U233, new_P2_R1203_U234,
    new_P2_R1203_U235, new_P2_R1203_U236, new_P2_R1203_U237,
    new_P2_R1203_U238, new_P2_R1203_U239, new_P2_R1203_U240,
    new_P2_R1203_U241, new_P2_R1203_U242, new_P2_R1203_U243,
    new_P2_R1203_U244, new_P2_R1203_U245, new_P2_R1203_U246,
    new_P2_R1203_U247, new_P2_R1203_U248, new_P2_R1203_U249,
    new_P2_R1203_U250, new_P2_R1203_U251, new_P2_R1203_U252,
    new_P2_R1203_U253, new_P2_R1203_U254, new_P2_R1203_U255,
    new_P2_R1203_U256, new_P2_R1203_U257, new_P2_R1203_U258,
    new_P2_R1203_U259, new_P2_R1203_U260, new_P2_R1203_U261,
    new_P2_R1203_U262, new_P2_R1203_U263, new_P2_R1203_U264,
    new_P2_R1203_U265, new_P2_R1203_U266, new_P2_R1203_U267,
    new_P2_R1203_U268, new_P2_R1203_U269, new_P2_R1203_U270,
    new_P2_R1203_U271, new_P2_R1203_U272, new_P2_R1203_U273,
    new_P2_R1203_U274, new_P2_R1203_U275, new_P2_R1203_U276,
    new_P2_R1203_U277, new_P2_R1203_U278, new_P2_R1203_U279,
    new_P2_R1203_U280, new_P2_R1203_U281, new_P2_R1203_U282,
    new_P2_R1203_U283, new_P2_R1203_U284, new_P2_R1203_U285,
    new_P2_R1203_U286, new_P2_R1203_U287, new_P2_R1203_U288,
    new_P2_R1203_U289, new_P2_R1203_U290, new_P2_R1203_U291,
    new_P2_R1203_U292, new_P2_R1203_U293, new_P2_R1203_U294,
    new_P2_R1203_U295, new_P2_R1203_U296, new_P2_R1203_U297,
    new_P2_R1203_U298, new_P2_R1203_U299, new_P2_R1203_U300,
    new_P2_R1203_U301, new_P2_R1203_U302, new_P2_R1203_U303,
    new_P2_R1203_U304, new_P2_R1203_U305, new_P2_R1203_U306,
    new_P2_R1203_U307, new_P2_R1203_U308, new_P2_R1203_U309,
    new_P2_R1203_U310, new_P2_R1203_U311, new_P2_R1203_U312,
    new_P2_R1203_U313, new_P2_R1203_U314, new_P2_R1203_U315,
    new_P2_R1203_U316, new_P2_R1203_U317, new_P2_R1203_U318,
    new_P2_R1203_U319, new_P2_R1203_U320, new_P2_R1203_U321,
    new_P2_R1203_U322, new_P2_R1203_U323, new_P2_R1203_U324,
    new_P2_R1203_U325, new_P2_R1203_U326, new_P2_R1203_U327,
    new_P2_R1203_U328, new_P2_R1203_U329, new_P2_R1203_U330,
    new_P2_R1203_U331, new_P2_R1203_U332, new_P2_R1203_U333,
    new_P2_R1203_U334, new_P2_R1203_U335, new_P2_R1203_U336,
    new_P2_R1203_U337, new_P2_R1203_U338, new_P2_R1203_U339,
    new_P2_R1203_U340, new_P2_R1203_U341, new_P2_R1203_U342,
    new_P2_R1203_U343, new_P2_R1203_U344, new_P2_R1203_U345,
    new_P2_R1203_U346, new_P2_R1203_U347, new_P2_R1203_U348,
    new_P2_R1203_U349, new_P2_R1203_U350, new_P2_R1203_U351,
    new_P2_R1203_U352, new_P2_R1203_U353, new_P2_R1203_U354,
    new_P2_R1203_U355, new_P2_R1203_U356, new_P2_R1203_U357,
    new_P2_R1203_U358, new_P2_R1203_U359, new_P2_R1203_U360,
    new_P2_R1203_U361, new_P2_R1203_U362, new_P2_R1203_U363,
    new_P2_R1203_U364, new_P2_R1203_U365, new_P2_R1203_U366,
    new_P2_R1203_U367, new_P2_R1203_U368, new_P2_R1203_U369,
    new_P2_R1203_U370, new_P2_R1203_U371, new_P2_R1203_U372,
    new_P2_R1203_U373, new_P2_R1203_U374, new_P2_R1203_U375,
    new_P2_R1203_U376, new_P2_R1203_U377, new_P2_R1203_U378,
    new_P2_R1203_U379, new_P2_R1203_U380, new_P2_R1203_U381,
    new_P2_R1203_U382, new_P2_R1203_U383, new_P2_R1203_U384,
    new_P2_R1203_U385, new_P2_R1203_U386, new_P2_R1203_U387,
    new_P2_R1203_U388, new_P2_R1203_U389, new_P2_R1203_U390,
    new_P2_R1203_U391, new_P2_R1203_U392, new_P2_R1203_U393,
    new_P2_R1203_U394, new_P2_R1203_U395, new_P2_R1203_U396,
    new_P2_R1203_U397, new_P2_R1203_U398, new_P2_R1203_U399,
    new_P2_R1203_U400, new_P2_R1203_U401, new_P2_R1203_U402,
    new_P2_R1203_U403, new_P2_R1203_U404, new_P2_R1203_U405,
    new_P2_R1203_U406, new_P2_R1203_U407, new_P2_R1203_U408,
    new_P2_R1203_U409, new_P2_R1203_U410, new_P2_R1203_U411,
    new_P2_R1203_U412, new_P2_R1203_U413, new_P2_R1203_U414,
    new_P2_R1203_U415, new_P2_R1203_U416, new_P2_R1203_U417,
    new_P2_R1203_U418, new_P2_R1203_U419, new_P2_R1203_U420,
    new_P2_R1203_U421, new_P2_R1203_U422, new_P2_R1203_U423,
    new_P2_R1203_U424, new_P2_R1203_U425, new_P2_R1203_U426,
    new_P2_R1203_U427, new_P2_R1203_U428, new_P2_R1203_U429,
    new_P2_R1203_U430, new_P2_R1203_U431, new_P2_R1203_U432,
    new_P2_R1203_U433, new_P2_R1203_U434, new_P2_R1203_U435,
    new_P2_R1203_U436, new_P2_R1203_U437, new_P2_R1203_U438,
    new_P2_R1203_U439, new_P2_R1203_U440, new_P2_R1203_U441,
    new_P2_R1203_U442, new_P2_R1203_U443, new_P2_R1203_U444,
    new_P2_R1203_U445, new_P2_R1203_U446, new_P2_R1203_U447,
    new_P2_R1203_U448, new_P2_R1203_U449, new_P2_R1203_U450,
    new_P2_R1203_U451, new_P2_R1203_U452, new_P2_R1203_U453,
    new_P2_R1203_U454, new_P2_R1203_U455, new_P2_R1203_U456,
    new_P2_R1203_U457, new_P2_R1203_U458, new_P2_R1203_U459,
    new_P2_R1203_U460, new_P2_R1203_U461, new_P2_R1203_U462,
    new_P2_R1203_U463, new_P2_R1203_U464, new_P2_R1203_U465,
    new_P2_R1203_U466, new_P2_R1203_U467, new_P2_R1203_U468,
    new_P2_R1203_U469, new_P2_R1203_U470, new_P2_R1203_U471,
    new_P2_R1203_U472, new_P2_R1203_U473, new_P2_R1203_U474,
    new_P2_R1203_U475, new_P2_R1203_U476, new_P2_R1203_U477,
    new_P2_R1203_U478, new_P2_R1113_U6, new_P2_R1113_U7, new_P2_R1113_U8,
    new_P2_R1113_U9, new_P2_R1113_U10, new_P2_R1113_U11, new_P2_R1113_U12,
    new_P2_R1113_U13, new_P2_R1113_U14, new_P2_R1113_U15, new_P2_R1113_U16,
    new_P2_R1113_U17, new_P2_R1113_U18, new_P2_R1113_U19, new_P2_R1113_U20,
    new_P2_R1113_U21, new_P2_R1113_U22, new_P2_R1113_U23, new_P2_R1113_U24,
    new_P2_R1113_U25, new_P2_R1113_U26, new_P2_R1113_U27, new_P2_R1113_U28,
    new_P2_R1113_U29, new_P2_R1113_U30, new_P2_R1113_U31, new_P2_R1113_U32,
    new_P2_R1113_U33, new_P2_R1113_U34, new_P2_R1113_U35, new_P2_R1113_U36,
    new_P2_R1113_U37, new_P2_R1113_U38, new_P2_R1113_U39, new_P2_R1113_U40,
    new_P2_R1113_U41, new_P2_R1113_U42, new_P2_R1113_U43, new_P2_R1113_U44,
    new_P2_R1113_U45, new_P2_R1113_U46, new_P2_R1113_U47, new_P2_R1113_U48,
    new_P2_R1113_U49, new_P2_R1113_U50, new_P2_R1113_U51, new_P2_R1113_U52,
    new_P2_R1113_U53, new_P2_R1113_U54, new_P2_R1113_U55, new_P2_R1113_U56,
    new_P2_R1113_U57, new_P2_R1113_U58, new_P2_R1113_U59, new_P2_R1113_U60,
    new_P2_R1113_U61, new_P2_R1113_U62, new_P2_R1113_U63, new_P2_R1113_U64,
    new_P2_R1113_U65, new_P2_R1113_U66, new_P2_R1113_U67, new_P2_R1113_U68,
    new_P2_R1113_U69, new_P2_R1113_U70, new_P2_R1113_U71, new_P2_R1113_U72,
    new_P2_R1113_U73, new_P2_R1113_U74, new_P2_R1113_U75, new_P2_R1113_U76,
    new_P2_R1113_U77, new_P2_R1113_U78, new_P2_R1113_U79, new_P2_R1113_U80,
    new_P2_R1113_U81, new_P2_R1113_U82, new_P2_R1113_U83, new_P2_R1113_U84,
    new_P2_R1113_U85, new_P2_R1113_U86, new_P2_R1113_U87, new_P2_R1113_U88,
    new_P2_R1113_U89, new_P2_R1113_U90, new_P2_R1113_U91, new_P2_R1113_U92,
    new_P2_R1113_U93, new_P2_R1113_U94, new_P2_R1113_U95, new_P2_R1113_U96,
    new_P2_R1113_U97, new_P2_R1113_U98, new_P2_R1113_U99,
    new_P2_R1113_U100, new_P2_R1113_U101, new_P2_R1113_U102,
    new_P2_R1113_U103, new_P2_R1113_U104, new_P2_R1113_U105,
    new_P2_R1113_U106, new_P2_R1113_U107, new_P2_R1113_U108,
    new_P2_R1113_U109, new_P2_R1113_U110, new_P2_R1113_U111,
    new_P2_R1113_U112, new_P2_R1113_U113, new_P2_R1113_U114,
    new_P2_R1113_U115, new_P2_R1113_U116, new_P2_R1113_U117,
    new_P2_R1113_U118, new_P2_R1113_U119, new_P2_R1113_U120,
    new_P2_R1113_U121, new_P2_R1113_U122, new_P2_R1113_U123,
    new_P2_R1113_U124, new_P2_R1113_U125, new_P2_R1113_U126,
    new_P2_R1113_U127, new_P2_R1113_U128, new_P2_R1113_U129,
    new_P2_R1113_U130, new_P2_R1113_U131, new_P2_R1113_U132,
    new_P2_R1113_U133, new_P2_R1113_U134, new_P2_R1113_U135,
    new_P2_R1113_U136, new_P2_R1113_U137, new_P2_R1113_U138,
    new_P2_R1113_U139, new_P2_R1113_U140, new_P2_R1113_U141,
    new_P2_R1113_U142, new_P2_R1113_U143, new_P2_R1113_U144,
    new_P2_R1113_U145, new_P2_R1113_U146, new_P2_R1113_U147,
    new_P2_R1113_U148, new_P2_R1113_U149, new_P2_R1113_U150,
    new_P2_R1113_U151, new_P2_R1113_U152, new_P2_R1113_U153,
    new_P2_R1113_U154, new_P2_R1113_U155, new_P2_R1113_U156,
    new_P2_R1113_U157, new_P2_R1113_U158, new_P2_R1113_U159,
    new_P2_R1113_U160, new_P2_R1113_U161, new_P2_R1113_U162,
    new_P2_R1113_U163, new_P2_R1113_U164, new_P2_R1113_U165,
    new_P2_R1113_U166, new_P2_R1113_U167, new_P2_R1113_U168,
    new_P2_R1113_U169, new_P2_R1113_U170, new_P2_R1113_U171,
    new_P2_R1113_U172, new_P2_R1113_U173, new_P2_R1113_U174,
    new_P2_R1113_U175, new_P2_R1113_U176, new_P2_R1113_U177,
    new_P2_R1113_U178, new_P2_R1113_U179, new_P2_R1113_U180,
    new_P2_R1113_U181, new_P2_R1113_U182, new_P2_R1113_U183,
    new_P2_R1113_U184, new_P2_R1113_U185, new_P2_R1113_U186,
    new_P2_R1113_U187, new_P2_R1113_U188, new_P2_R1113_U189,
    new_P2_R1113_U190, new_P2_R1113_U191, new_P2_R1113_U192,
    new_P2_R1113_U193, new_P2_R1113_U194, new_P2_R1113_U195,
    new_P2_R1113_U196, new_P2_R1113_U197, new_P2_R1113_U198,
    new_P2_R1113_U199, new_P2_R1113_U200, new_P2_R1113_U201,
    new_P2_R1113_U202, new_P2_R1113_U203, new_P2_R1113_U204,
    new_P2_R1113_U205, new_P2_R1113_U206, new_P2_R1113_U207,
    new_P2_R1113_U208, new_P2_R1113_U209, new_P2_R1113_U210,
    new_P2_R1113_U211, new_P2_R1113_U212, new_P2_R1113_U213,
    new_P2_R1113_U214, new_P2_R1113_U215, new_P2_R1113_U216,
    new_P2_R1113_U217, new_P2_R1113_U218, new_P2_R1113_U219,
    new_P2_R1113_U220, new_P2_R1113_U221, new_P2_R1113_U222,
    new_P2_R1113_U223, new_P2_R1113_U224, new_P2_R1113_U225,
    new_P2_R1113_U226, new_P2_R1113_U227, new_P2_R1113_U228,
    new_P2_R1113_U229, new_P2_R1113_U230, new_P2_R1113_U231,
    new_P2_R1113_U232, new_P2_R1113_U233, new_P2_R1113_U234,
    new_P2_R1113_U235, new_P2_R1113_U236, new_P2_R1113_U237,
    new_P2_R1113_U238, new_P2_R1113_U239, new_P2_R1113_U240,
    new_P2_R1113_U241, new_P2_R1113_U242, new_P2_R1113_U243,
    new_P2_R1113_U244, new_P2_R1113_U245, new_P2_R1113_U246,
    new_P2_R1113_U247, new_P2_R1113_U248, new_P2_R1113_U249,
    new_P2_R1113_U250, new_P2_R1113_U251, new_P2_R1113_U252,
    new_P2_R1113_U253, new_P2_R1113_U254, new_P2_R1113_U255,
    new_P2_R1113_U256, new_P2_R1113_U257, new_P2_R1113_U258,
    new_P2_R1113_U259, new_P2_R1113_U260, new_P2_R1113_U261,
    new_P2_R1113_U262, new_P2_R1113_U263, new_P2_R1113_U264,
    new_P2_R1113_U265, new_P2_R1113_U266, new_P2_R1113_U267,
    new_P2_R1113_U268, new_P2_R1113_U269, new_P2_R1113_U270,
    new_P2_R1113_U271, new_P2_R1113_U272, new_P2_R1113_U273,
    new_P2_R1113_U274, new_P2_R1113_U275, new_P2_R1113_U276,
    new_P2_R1113_U277, new_P2_R1113_U278, new_P2_R1113_U279,
    new_P2_R1113_U280, new_P2_R1113_U281, new_P2_R1113_U282,
    new_P2_R1113_U283, new_P2_R1113_U284, new_P2_R1113_U285,
    new_P2_R1113_U286, new_P2_R1113_U287, new_P2_R1113_U288,
    new_P2_R1113_U289, new_P2_R1113_U290, new_P2_R1113_U291,
    new_P2_R1113_U292, new_P2_R1113_U293, new_P2_R1113_U294,
    new_P2_R1113_U295, new_P2_R1113_U296, new_P2_R1113_U297,
    new_P2_R1113_U298, new_P2_R1113_U299, new_P2_R1113_U300,
    new_P2_R1113_U301, new_P2_R1113_U302, new_P2_R1113_U303,
    new_P2_R1113_U304, new_P2_R1113_U305, new_P2_R1113_U306,
    new_P2_R1113_U307, new_P2_R1113_U308, new_P2_R1113_U309,
    new_P2_R1113_U310, new_P2_R1113_U311, new_P2_R1113_U312,
    new_P2_R1113_U313, new_P2_R1113_U314, new_P2_R1113_U315,
    new_P2_R1113_U316, new_P2_R1113_U317, new_P2_R1113_U318,
    new_P2_R1113_U319, new_P2_R1113_U320, new_P2_R1113_U321,
    new_P2_R1113_U322, new_P2_R1113_U323, new_P2_R1113_U324,
    new_P2_R1113_U325, new_P2_R1113_U326, new_P2_R1113_U327,
    new_P2_R1113_U328, new_P2_R1113_U329, new_P2_R1113_U330,
    new_P2_R1113_U331, new_P2_R1113_U332, new_P2_R1113_U333,
    new_P2_R1113_U334, new_P2_R1113_U335, new_P2_R1113_U336,
    new_P2_R1113_U337, new_P2_R1113_U338, new_P2_R1113_U339,
    new_P2_R1113_U340, new_P2_R1113_U341, new_P2_R1113_U342,
    new_P2_R1113_U343, new_P2_R1113_U344, new_P2_R1113_U345,
    new_P2_R1113_U346, new_P2_R1113_U347, new_P2_R1113_U348,
    new_P2_R1113_U349, new_P2_R1113_U350, new_P2_R1113_U351,
    new_P2_R1113_U352, new_P2_R1113_U353, new_P2_R1113_U354,
    new_P2_R1113_U355, new_P2_R1113_U356, new_P2_R1113_U357,
    new_P2_R1113_U358, new_P2_R1113_U359, new_P2_R1113_U360,
    new_P2_R1113_U361, new_P2_R1113_U362, new_P2_R1113_U363,
    new_P2_R1113_U364, new_P2_R1113_U365, new_P2_R1113_U366,
    new_P2_R1113_U367, new_P2_R1113_U368, new_P2_R1113_U369,
    new_P2_R1113_U370, new_P2_R1113_U371, new_P2_R1113_U372,
    new_P2_R1113_U373, new_P2_R1113_U374, new_P2_R1113_U375,
    new_P2_R1113_U376, new_P2_R1113_U377, new_P2_R1113_U378,
    new_P2_R1113_U379, new_P2_R1113_U380, new_P2_R1113_U381,
    new_P2_R1113_U382, new_P2_R1113_U383, new_P2_R1113_U384,
    new_P2_R1113_U385, new_P2_R1113_U386, new_P2_R1113_U387,
    new_P2_R1113_U388, new_P2_R1113_U389, new_P2_R1113_U390,
    new_P2_R1113_U391, new_P2_R1113_U392, new_P2_R1113_U393,
    new_P2_R1113_U394, new_P2_R1113_U395, new_P2_R1113_U396,
    new_P2_R1113_U397, new_P2_R1113_U398, new_P2_R1113_U399,
    new_P2_R1113_U400, new_P2_R1113_U401, new_P2_R1113_U402,
    new_P2_R1113_U403, new_P2_R1113_U404, new_P2_R1113_U405,
    new_P2_R1113_U406, new_P2_R1113_U407, new_P2_R1113_U408,
    new_P2_R1113_U409, new_P2_R1113_U410, new_P2_R1113_U411,
    new_P2_R1113_U412, new_P2_R1113_U413, new_P2_R1113_U414,
    new_P2_R1113_U415, new_P2_R1113_U416, new_P2_R1113_U417,
    new_P2_R1113_U418, new_P2_R1113_U419, new_P2_R1113_U420,
    new_P2_R1113_U421, new_P2_R1113_U422, new_P2_R1113_U423,
    new_P2_R1113_U424, new_P2_R1113_U425, new_P2_R1113_U426,
    new_P2_R1113_U427, new_P2_R1113_U428, new_P2_R1113_U429,
    new_P2_R1113_U430, new_P2_R1113_U431, new_P2_R1113_U432,
    new_P2_R1113_U433, new_P2_R1113_U434, new_P2_R1113_U435,
    new_P2_R1113_U436, new_P2_R1113_U437, new_P2_R1113_U438,
    new_P2_R1113_U439, new_P2_R1113_U440, new_P2_R1113_U441,
    new_P2_R1113_U442, new_P2_R1113_U443, new_P2_R1113_U444,
    new_P2_R1113_U445, new_P2_R1113_U446, new_P2_R1113_U447,
    new_P2_R1113_U448, new_P2_R1113_U449, new_P2_R1113_U450,
    new_P2_R1113_U451, new_P2_R1113_U452, new_P2_R1113_U453,
    new_P2_R1113_U454, new_P2_R1113_U455, new_P2_R1113_U456,
    new_P2_R1113_U457, new_P2_R1113_U458, new_P2_R1113_U459,
    new_P2_R1113_U460, new_P2_R1113_U461, new_P2_R1113_U462,
    new_P2_R1113_U463, new_P2_R1113_U464, new_P2_R1113_U465,
    new_P2_R1113_U466, new_P2_R1113_U467, new_P2_R1113_U468,
    new_P2_R1113_U469, new_P2_R1113_U470, new_P2_R1113_U471,
    new_P2_R1113_U472, new_P2_R1113_U473, new_P2_R1113_U474,
    new_P2_R1113_U475, new_P2_R1113_U476, new_P2_R1113_U477,
    new_P2_R1113_U478, new_P3_SUB_598_U6, new_P3_SUB_598_U7,
    new_P3_SUB_598_U8, new_P3_SUB_598_U9, new_P3_SUB_598_U10,
    new_P3_SUB_598_U11, new_P3_SUB_598_U12, new_P3_SUB_598_U13,
    new_P3_SUB_598_U14, new_P3_SUB_598_U15, new_P3_SUB_598_U16,
    new_P3_SUB_598_U17, new_P3_SUB_598_U18, new_P3_SUB_598_U19,
    new_P3_SUB_598_U20, new_P3_SUB_598_U21, new_P3_SUB_598_U22,
    new_P3_SUB_598_U23, new_P3_SUB_598_U24, new_P3_SUB_598_U25,
    new_P3_SUB_598_U26, new_P3_SUB_598_U27, new_P3_SUB_598_U28,
    new_P3_SUB_598_U29, new_P3_SUB_598_U30, new_P3_SUB_598_U31,
    new_P3_SUB_598_U32, new_P3_SUB_598_U33, new_P3_SUB_598_U34,
    new_P3_SUB_598_U35, new_P3_SUB_598_U36, new_P3_SUB_598_U37,
    new_P3_SUB_598_U38, new_P3_SUB_598_U39, new_P3_SUB_598_U40,
    new_P3_SUB_598_U41, new_P3_SUB_598_U42, new_P3_SUB_598_U43,
    new_P3_SUB_598_U44, new_P3_SUB_598_U45, new_P3_SUB_598_U46,
    new_P3_SUB_598_U47, new_P3_SUB_598_U48, new_P3_SUB_598_U49,
    new_P3_SUB_598_U50, new_P3_SUB_598_U51, new_P3_SUB_598_U52,
    new_P3_SUB_598_U53, new_P3_SUB_598_U54, new_P3_SUB_598_U55,
    new_P3_SUB_598_U56, new_P3_SUB_598_U57, new_P3_SUB_598_U58,
    new_P3_SUB_598_U59, new_P3_SUB_598_U60, new_P3_SUB_598_U61,
    new_P3_SUB_598_U62, new_P3_SUB_598_U63, new_P3_SUB_598_U64,
    new_P3_SUB_598_U65, new_P3_SUB_598_U66, new_P3_SUB_598_U67,
    new_P3_SUB_598_U68, new_P3_SUB_598_U69, new_P3_SUB_598_U70,
    new_P3_SUB_598_U71, new_P3_SUB_598_U72, new_P3_SUB_598_U73,
    new_P3_SUB_598_U74, new_P3_SUB_598_U75, new_P3_SUB_598_U76,
    new_P3_SUB_598_U77, new_P3_SUB_598_U78, new_P3_SUB_598_U79,
    new_P3_SUB_598_U80, new_P3_SUB_598_U81, new_P3_SUB_598_U82,
    new_P3_SUB_598_U83, new_P3_SUB_598_U84, new_P3_SUB_598_U85,
    new_P3_SUB_598_U86, new_P3_SUB_598_U87, new_P3_SUB_598_U88,
    new_P3_SUB_598_U89, new_P3_SUB_598_U90, new_P3_SUB_598_U91,
    new_P3_SUB_598_U92, new_P3_SUB_598_U93, new_P3_SUB_598_U94,
    new_P3_SUB_598_U95, new_P3_SUB_598_U96, new_P3_SUB_598_U97,
    new_P3_SUB_598_U98, new_P3_SUB_598_U99, new_P3_SUB_598_U100,
    new_P3_SUB_598_U101, new_P3_SUB_598_U102, new_P3_SUB_598_U103,
    new_P3_SUB_598_U104, new_P3_SUB_598_U105, new_P3_SUB_598_U106,
    new_P3_SUB_598_U107, new_P3_SUB_598_U108, new_P3_SUB_598_U109,
    new_P3_SUB_598_U110, new_P3_SUB_598_U111, new_P3_SUB_598_U112,
    new_P3_SUB_598_U113, new_P3_SUB_598_U114, new_P3_SUB_598_U115,
    new_P3_SUB_598_U116, new_P3_SUB_598_U117, new_P3_SUB_598_U118,
    new_P3_SUB_598_U119, new_P3_SUB_598_U120, new_P3_SUB_598_U121,
    new_P3_SUB_598_U122, new_P3_SUB_598_U123, new_P3_SUB_598_U124,
    new_P3_SUB_598_U125, new_P3_SUB_598_U126, new_P3_SUB_598_U127,
    new_P3_SUB_598_U128, new_P3_SUB_598_U129, new_P3_SUB_598_U130,
    new_P3_SUB_598_U131, new_P3_SUB_598_U132, new_P3_SUB_598_U133,
    new_P3_SUB_598_U134, new_P3_SUB_598_U135, new_P3_SUB_598_U136,
    new_P3_SUB_598_U137, new_P3_SUB_598_U138, new_P3_SUB_598_U139,
    new_P3_SUB_598_U140, new_P3_SUB_598_U141, new_P3_SUB_598_U142,
    new_P3_SUB_598_U143, new_P3_SUB_598_U144, new_P3_SUB_598_U145,
    new_P3_SUB_598_U146, new_P3_SUB_598_U147, new_P3_SUB_598_U148,
    new_P3_SUB_598_U149, new_P3_SUB_598_U150, new_P3_SUB_598_U151,
    new_P3_SUB_598_U152, new_P3_SUB_598_U153, new_P3_SUB_598_U154,
    new_P3_SUB_598_U155, new_P3_SUB_598_U156, new_P3_SUB_598_U157,
    new_P3_SUB_598_U158, new_P3_SUB_598_U159, new_P3_SUB_598_U160,
    new_P3_R693_U6, new_P3_R693_U7, new_P3_R693_U8, new_P3_R693_U9,
    new_P3_R693_U10, new_P3_R693_U11, new_P3_R693_U12, new_P3_R693_U13,
    new_P3_R693_U14, new_P3_R693_U15, new_P3_R693_U16, new_P3_R693_U17,
    new_P3_R693_U18, new_P3_R693_U19, new_P3_R693_U20, new_P3_R693_U21,
    new_P3_R693_U22, new_P3_R693_U23, new_P3_R693_U24, new_P3_R693_U25,
    new_P3_R693_U26, new_P3_R693_U27, new_P3_R693_U28, new_P3_R693_U29,
    new_P3_R693_U30, new_P3_R693_U31, new_P3_R693_U32, new_P3_R693_U33,
    new_P3_R693_U34, new_P3_R693_U35, new_P3_R693_U36, new_P3_R693_U37,
    new_P3_R693_U38, new_P3_R693_U39, new_P3_R693_U40, new_P3_R693_U41,
    new_P3_R693_U42, new_P3_R693_U43, new_P3_R693_U44, new_P3_R693_U45,
    new_P3_R693_U46, new_P3_R693_U47, new_P3_R693_U48, new_P3_R693_U49,
    new_P3_R693_U50, new_P3_R693_U51, new_P3_R693_U52, new_P3_R693_U53,
    new_P3_R693_U54, new_P3_R693_U55, new_P3_R693_U56, new_P3_R693_U57,
    new_P3_R693_U58, new_P3_R693_U59, new_P3_R693_U60, new_P3_R693_U61,
    new_P3_R693_U62, new_P3_R693_U63, new_P3_R693_U64, new_P3_R693_U65,
    new_P3_R693_U66, new_P3_R693_U67, new_P3_R693_U68, new_P3_R693_U69,
    new_P3_R693_U70, new_P3_R693_U71, new_P3_R693_U72, new_P3_R693_U73,
    new_P3_R693_U74, new_P3_R693_U75, new_P3_R693_U76, new_P3_R693_U77,
    new_P3_R693_U78, new_P3_R693_U79, new_P3_R693_U80, new_P3_R693_U81,
    new_P3_R693_U82, new_P3_R693_U83, new_P3_R693_U84, new_P3_R693_U85,
    new_P3_R693_U86, new_P3_R693_U87, new_P3_R693_U88, new_P3_R693_U89,
    new_P3_R693_U90, new_P3_R693_U91, new_P3_R693_U92, new_P3_R693_U93,
    new_P3_R693_U94, new_P3_R693_U95, new_P3_R693_U96, new_P3_R693_U97,
    new_P3_R693_U98, new_P3_R693_U99, new_P3_R693_U100, new_P3_R693_U101,
    new_P3_R693_U102, new_P3_R693_U103, new_P3_R693_U104, new_P3_R693_U105,
    new_P3_R693_U106, new_P3_R693_U107, new_P3_R693_U108, new_P3_R693_U109,
    new_P3_R693_U110, new_P3_R693_U111, new_P3_R693_U112, new_P3_R693_U113,
    new_P3_R693_U114, new_P3_R693_U115, new_P3_R693_U116, new_P3_R693_U117,
    new_P3_R693_U118, new_P3_R693_U119, new_P3_R693_U120, new_P3_R693_U121,
    new_P3_R693_U122, new_P3_R693_U123, new_P3_R693_U124, new_P3_R693_U125,
    new_P3_R693_U126, new_P3_R693_U127, new_P3_R693_U128, new_P3_R693_U129,
    new_P3_R693_U130, new_P3_R693_U131, new_P3_R693_U132, new_P3_R693_U133,
    new_P3_R693_U134, new_P3_R693_U135, new_P3_R693_U136, new_P3_R693_U137,
    new_P3_R693_U138, new_P3_R693_U139, new_P3_R693_U140, new_P3_R693_U141,
    new_P3_R693_U142, new_P3_R693_U143, new_P3_R693_U144, new_P3_R693_U145,
    new_P3_R693_U146, new_P3_R693_U147, new_P3_R693_U148, new_P3_R693_U149,
    new_P3_R693_U150, new_P3_R693_U151, new_P3_R693_U152, new_P3_R693_U153,
    new_P3_R693_U154, new_P3_R693_U155, new_P3_R693_U156, new_P3_R693_U157,
    new_P3_R693_U158, new_P3_R693_U159, new_P3_R693_U160, new_P3_R693_U161,
    new_P3_R693_U162, new_P3_R693_U163, new_P3_R693_U164, new_P3_R693_U165,
    new_P3_R693_U166, new_P3_R693_U167, new_P3_R693_U168, new_P3_R693_U169,
    new_P3_R693_U170, new_P3_R693_U171, new_P3_R693_U172, new_P3_R693_U173,
    new_P3_R693_U174, new_P3_R693_U175, new_P3_R693_U176, new_P3_R693_U177,
    new_P3_R693_U178, new_P3_R693_U179, new_P3_R693_U180, new_P3_R693_U181,
    new_P3_R693_U182, new_P3_R693_U183, new_P3_R693_U184, new_P3_R693_U185,
    new_P3_R693_U186, new_P3_R693_U187, new_P3_R693_U188, new_P3_R693_U189,
    new_P3_R693_U190, new_P3_R693_U191, new_P3_R693_U192, new_P3_R693_U193,
    new_P3_R693_U194, new_P3_R693_U195, new_P3_R693_U196,
    new_P3_SUB_609_U6, new_P3_SUB_609_U7, new_P3_SUB_609_U8,
    new_P3_SUB_609_U9, new_P3_SUB_609_U10, new_P3_SUB_609_U11,
    new_P3_SUB_609_U12, new_P3_SUB_609_U13, new_P3_SUB_609_U14,
    new_P3_SUB_609_U15, new_P3_SUB_609_U16, new_P3_SUB_609_U17,
    new_P3_SUB_609_U18, new_P3_SUB_609_U19, new_P3_SUB_609_U20,
    new_P3_SUB_609_U21, new_P3_SUB_609_U22, new_P3_SUB_609_U23,
    new_P3_SUB_609_U24, new_P3_SUB_609_U25, new_P3_SUB_609_U26,
    new_P3_SUB_609_U27, new_P3_SUB_609_U28, new_P3_SUB_609_U29,
    new_P3_SUB_609_U30, new_P3_SUB_609_U31, new_P3_SUB_609_U32,
    new_P3_SUB_609_U33, new_P3_SUB_609_U34, new_P3_SUB_609_U35,
    new_P3_SUB_609_U36, new_P3_SUB_609_U37, new_P3_SUB_609_U38,
    new_P3_SUB_609_U39, new_P3_SUB_609_U40, new_P3_SUB_609_U41,
    new_P3_SUB_609_U42, new_P3_SUB_609_U43, new_P3_SUB_609_U44,
    new_P3_SUB_609_U45, new_P3_SUB_609_U46, new_P3_SUB_609_U47,
    new_P3_SUB_609_U48, new_P3_SUB_609_U49, new_P3_SUB_609_U50,
    new_P3_SUB_609_U51, new_P3_SUB_609_U52, new_P3_SUB_609_U53,
    new_P3_SUB_609_U54, new_P3_SUB_609_U55, new_P3_SUB_609_U56,
    new_P3_SUB_609_U57, new_P3_SUB_609_U58, new_P3_SUB_609_U59,
    new_P3_SUB_609_U60, new_P3_SUB_609_U61, new_P3_SUB_609_U62,
    new_P3_SUB_609_U63, new_P3_SUB_609_U64, new_P3_SUB_609_U65,
    new_P3_SUB_609_U66, new_P3_SUB_609_U67, new_P3_SUB_609_U68,
    new_P3_SUB_609_U69, new_P3_SUB_609_U70, new_P3_SUB_609_U71,
    new_P3_SUB_609_U72, new_P3_SUB_609_U73, new_P3_SUB_609_U74,
    new_P3_SUB_609_U75, new_P3_SUB_609_U76, new_P3_SUB_609_U77,
    new_P3_SUB_609_U78, new_P3_SUB_609_U79, new_P3_SUB_609_U80,
    new_P3_SUB_609_U81, new_P3_SUB_609_U82, new_P3_SUB_609_U83,
    new_P3_SUB_609_U84, new_P3_SUB_609_U85, new_P3_SUB_609_U86,
    new_P3_SUB_609_U87, new_P3_SUB_609_U88, new_P3_SUB_609_U89,
    new_P3_SUB_609_U90, new_P3_SUB_609_U91, new_P3_SUB_609_U92,
    new_P3_SUB_609_U93, new_P3_SUB_609_U94, new_P3_SUB_609_U95,
    new_P3_SUB_609_U96, new_P3_SUB_609_U97, new_P3_SUB_609_U98,
    new_P3_SUB_609_U99, new_P3_SUB_609_U100, new_P3_SUB_609_U101,
    new_P3_SUB_609_U102, new_P3_SUB_609_U103, new_P3_SUB_609_U104,
    new_P3_SUB_609_U105, new_P3_SUB_609_U106, new_P3_SUB_609_U107,
    new_P3_SUB_609_U108, new_P3_SUB_609_U109, new_P3_SUB_609_U110,
    new_P3_SUB_609_U111, new_P3_SUB_609_U112, new_P3_SUB_609_U113,
    new_P3_SUB_609_U114, new_P3_SUB_609_U115, new_P3_R1095_U6,
    new_P3_R1095_U7, new_P3_R1095_U8, new_P3_R1095_U9, new_P3_R1095_U10,
    new_P3_R1095_U11, new_P3_R1095_U12, new_P3_R1095_U13, new_P3_R1095_U14,
    new_P3_R1095_U15, new_P3_R1095_U16, new_P3_R1095_U17, new_P3_R1095_U18,
    new_P3_R1095_U19, new_P3_R1095_U20, new_P3_R1095_U21, new_P3_R1095_U22,
    new_P3_R1095_U23, new_P3_R1095_U24, new_P3_R1095_U25, new_P3_R1095_U26,
    new_P3_R1095_U27, new_P3_R1095_U28, new_P3_R1095_U29, new_P3_R1095_U30,
    new_P3_R1095_U31, new_P3_R1095_U32, new_P3_R1095_U33, new_P3_R1095_U34,
    new_P3_R1095_U35, new_P3_R1095_U36, new_P3_R1095_U37, new_P3_R1095_U38,
    new_P3_R1095_U39, new_P3_R1095_U40, new_P3_R1095_U41, new_P3_R1095_U42,
    new_P3_R1095_U43, new_P3_R1095_U44, new_P3_R1095_U45, new_P3_R1095_U46,
    new_P3_R1095_U47, new_P3_R1095_U48, new_P3_R1095_U49, new_P3_R1095_U50,
    new_P3_R1095_U51, new_P3_R1095_U52, new_P3_R1095_U53, new_P3_R1095_U54,
    new_P3_R1095_U55, new_P3_R1095_U56, new_P3_R1095_U57, new_P3_R1095_U58,
    new_P3_R1095_U59, new_P3_R1095_U60, new_P3_R1095_U61, new_P3_R1095_U62,
    new_P3_R1095_U63, new_P3_R1095_U64, new_P3_R1095_U65, new_P3_R1095_U66,
    new_P3_R1095_U67, new_P3_R1095_U68, new_P3_R1095_U69, new_P3_R1095_U70,
    new_P3_R1095_U71, new_P3_R1095_U72, new_P3_R1095_U73, new_P3_R1095_U74,
    new_P3_R1095_U75, new_P3_R1095_U76, new_P3_R1095_U77, new_P3_R1095_U78,
    new_P3_R1095_U79, new_P3_R1095_U80, new_P3_R1095_U81, new_P3_R1095_U82,
    new_P3_R1095_U83, new_P3_R1095_U84, new_P3_R1095_U85, new_P3_R1095_U86,
    new_P3_R1095_U87, new_P3_R1095_U88, new_P3_R1095_U89, new_P3_R1095_U90,
    new_P3_R1095_U91, new_P3_R1095_U92, new_P3_R1095_U93, new_P3_R1095_U94,
    new_P3_R1095_U95, new_P3_R1095_U96, new_P3_R1095_U97, new_P3_R1095_U98,
    new_P3_R1095_U99, new_P3_R1095_U100, new_P3_R1095_U101,
    new_P3_R1095_U102, new_P3_R1095_U103, new_P3_R1095_U104,
    new_P3_R1095_U105, new_P3_R1095_U106, new_P3_R1095_U107,
    new_P3_R1095_U108, new_P3_R1095_U109, new_P3_R1095_U110,
    new_P3_R1095_U111, new_P3_R1095_U112, new_P3_R1095_U113,
    new_P3_R1095_U114, new_P3_R1095_U115, new_P3_R1095_U116,
    new_P3_R1095_U117, new_P3_R1095_U118, new_P3_R1095_U119,
    new_P3_R1095_U120, new_P3_R1095_U121, new_P3_R1095_U122,
    new_P3_R1095_U123, new_P3_R1095_U124, new_P3_R1095_U125,
    new_P3_R1095_U126, new_P3_R1095_U127, new_P3_R1095_U128,
    new_P3_R1095_U129, new_P3_R1095_U130, new_P3_R1095_U131,
    new_P3_R1095_U132, new_P3_R1095_U133, new_P3_R1095_U134,
    new_P3_R1095_U135, new_P3_R1095_U136, new_P3_R1095_U137,
    new_P3_R1095_U138, new_P3_R1095_U139, new_P3_R1095_U140,
    new_P3_R1095_U141, new_P3_R1095_U142, new_P3_R1095_U143,
    new_P3_R1095_U144, new_P3_R1095_U145, new_P3_R1095_U146,
    new_P3_R1095_U147, new_P3_R1095_U148, new_P3_R1095_U149,
    new_P3_R1095_U150, new_P3_R1095_U151, new_P3_R1095_U152,
    new_P3_R1095_U153, new_P3_R1095_U154, new_P3_R1095_U155,
    new_P3_R1095_U156, new_P3_R1095_U157, new_P3_R1095_U158,
    new_P3_R1095_U159, new_P3_R1095_U160, new_P3_R1095_U161,
    new_P3_R1095_U162, new_P3_R1095_U163, new_P3_R1095_U164,
    new_P3_R1095_U165, new_P3_R1095_U166, new_P3_R1095_U167,
    new_P3_R1095_U168, new_P3_R1095_U169, new_P3_R1095_U170,
    new_P3_R1095_U171, new_P3_R1095_U172, new_P3_R1095_U173,
    new_P3_R1095_U174, new_P3_R1095_U175, new_P3_R1095_U176,
    new_P3_R1095_U177, new_P3_R1095_U178, new_P3_R1095_U179,
    new_P3_R1095_U180, new_P3_R1095_U181, new_P3_R1095_U182,
    new_P3_R1095_U183, new_P3_R1095_U184, new_P3_R1095_U185,
    new_P3_R1095_U186, new_P3_R1095_U187, new_P3_R1095_U188,
    new_P3_R1095_U189, new_P3_R1095_U190, new_P3_R1095_U191,
    new_P3_R1095_U192, new_P3_R1095_U193, new_P3_R1095_U194,
    new_P3_R1095_U195, new_P3_R1095_U196, new_P3_R1095_U197,
    new_P3_R1095_U198, new_P3_R1095_U199, new_P3_R1095_U200,
    new_P3_R1095_U201, new_P3_R1095_U202, new_P3_R1095_U203,
    new_P3_R1095_U204, new_P3_R1095_U205, new_P3_R1095_U206,
    new_P3_R1095_U207, new_P3_R1095_U208, new_P3_R1095_U209,
    new_P3_R1095_U210, new_P3_R1095_U211, new_P3_R1095_U212,
    new_P3_R1095_U213, new_P3_R1095_U214, new_P3_R1095_U215,
    new_P3_R1095_U216, new_P3_R1095_U217, new_P3_R1095_U218,
    new_P3_R1095_U219, new_P3_R1095_U220, new_P3_R1095_U221,
    new_P3_R1095_U222, new_P3_R1095_U223, new_P3_R1095_U224,
    new_P3_R1095_U225, new_P3_R1095_U226, new_P3_R1095_U227,
    new_P3_R1095_U228, new_P3_R1095_U229, new_P3_R1095_U230,
    new_P3_R1095_U231, new_P3_R1095_U232, new_P3_R1095_U233,
    new_P3_R1095_U234, new_P3_R1095_U235, new_P3_R1095_U236,
    new_P3_R1095_U237, new_P3_R1095_U238, new_P3_R1095_U239,
    new_P3_R1095_U240, new_P3_R1095_U241, new_P3_R1095_U242,
    new_P3_R1095_U243, new_P3_R1095_U244, new_P3_R1095_U245,
    new_P3_R1095_U246, new_P3_R1095_U247, new_P3_R1095_U248,
    new_P3_R1095_U249, new_P3_R1095_U250, new_P3_R1095_U251,
    new_P3_R1095_U252, new_P3_R1095_U253, new_P3_R1095_U254,
    new_P3_R1095_U255, new_P3_R1095_U256, new_P3_R1095_U257,
    new_P3_R1095_U258, new_P3_R1095_U259, new_P3_R1095_U260,
    new_P3_R1095_U261, new_P3_R1095_U262, new_P3_R1095_U263,
    new_P3_R1095_U264, new_P3_R1095_U265, new_P3_R1095_U266,
    new_P3_R1095_U267, new_P3_R1095_U268, new_P3_R1095_U269,
    new_P3_R1095_U270, new_P3_R1095_U271, new_P3_R1095_U272,
    new_P3_R1095_U273, new_P3_R1095_U274, new_P3_R1095_U275,
    new_P3_R1095_U276, new_P3_R1095_U277, new_P3_R1095_U278,
    new_P3_R1095_U279, new_P3_R1095_U280, new_P3_R1095_U281,
    new_P3_R1095_U282, new_P3_R1095_U283, new_P3_R1095_U284,
    new_P3_R1095_U285, new_P3_R1095_U286, new_P3_R1095_U287,
    new_P3_R1095_U288, new_P3_R1095_U289, new_P3_R1095_U290,
    new_P3_R1095_U291, new_P3_R1095_U292, new_P3_R1095_U293,
    new_P3_R1095_U294, new_P3_R1095_U295, new_P3_R1095_U296,
    new_P3_R1095_U297, new_P3_R1095_U298, new_P3_R1095_U299,
    new_P3_R1095_U300, new_P3_R1095_U301, new_P3_R1095_U302,
    new_P3_R1095_U303, new_P3_R1095_U304, new_P3_R1095_U305,
    new_P3_R1095_U306, new_P3_R1095_U307, new_P3_R1095_U308,
    new_P3_R1095_U309, new_P3_R1095_U310, new_P3_R1095_U311,
    new_P3_R1095_U312, new_P3_R1095_U313, new_P3_R1095_U314,
    new_P3_R1095_U315, new_P3_R1095_U316, new_P3_R1095_U317,
    new_P3_R1095_U318, new_P3_R1095_U319, new_P3_R1095_U320,
    new_P3_R1095_U321, new_P3_R1095_U322, new_P3_R1095_U323,
    new_P3_R1095_U324, new_P3_R1095_U325, new_P3_R1095_U326,
    new_P3_R1095_U327, new_P3_R1095_U328, new_P3_R1095_U329,
    new_P3_R1095_U330, new_P3_R1095_U331, new_P3_R1095_U332,
    new_P3_R1095_U333, new_P3_R1095_U334, new_P3_R1095_U335,
    new_P3_R1095_U336, new_P3_R1095_U337, new_P3_R1095_U338,
    new_P3_R1095_U339, new_P3_R1095_U340, new_P3_R1095_U341,
    new_P3_R1095_U342, new_P3_R1095_U343, new_P3_R1095_U344,
    new_P3_R1095_U345, new_P3_R1095_U346, new_P3_R1095_U347,
    new_P3_R1095_U348, new_P3_R1095_U349, new_P3_R1095_U350,
    new_P3_R1095_U351, new_P3_R1095_U352, new_P3_R1095_U353,
    new_P3_R1095_U354, new_P3_R1095_U355, new_P3_R1095_U356,
    new_P3_R1095_U357, new_P3_R1095_U358, new_P3_R1095_U359,
    new_P3_R1095_U360, new_P3_R1095_U361, new_P3_R1095_U362,
    new_P3_R1095_U363, new_P3_R1095_U364, new_P3_R1095_U365,
    new_P3_R1095_U366, new_P3_R1095_U367, new_P3_R1095_U368,
    new_P3_R1095_U369, new_P3_R1095_U370, new_P3_R1095_U371,
    new_P3_R1095_U372, new_P3_R1095_U373, new_P3_R1095_U374,
    new_P3_R1095_U375, new_P3_R1095_U376, new_P3_R1095_U377,
    new_P3_R1095_U378, new_P3_R1095_U379, new_P3_R1095_U380,
    new_P3_R1095_U381, new_P3_R1095_U382, new_P3_R1095_U383,
    new_P3_R1095_U384, new_P3_R1095_U385, new_P3_R1095_U386,
    new_P3_R1095_U387, new_P3_R1095_U388, new_P3_R1095_U389,
    new_P3_R1095_U390, new_P3_R1095_U391, new_P3_R1095_U392,
    new_P3_R1095_U393, new_P3_R1095_U394, new_P3_R1095_U395,
    new_P3_R1095_U396, new_P3_R1095_U397, new_P3_R1095_U398,
    new_P3_R1095_U399, new_P3_R1095_U400, new_P3_R1095_U401,
    new_P3_R1095_U402, new_P3_R1095_U403, new_P3_R1095_U404,
    new_P3_R1095_U405, new_P3_R1095_U406, new_P3_R1095_U407,
    new_P3_R1095_U408, new_P3_R1095_U409, new_P3_R1095_U410,
    new_P3_R1095_U411, new_P3_R1095_U412, new_P3_R1095_U413,
    new_P3_R1095_U414, new_P3_R1095_U415, new_P3_R1095_U416,
    new_P3_R1095_U417, new_P3_R1095_U418, new_P3_R1095_U419,
    new_P3_R1095_U420, new_P3_R1095_U421, new_P3_R1095_U422,
    new_P3_R1095_U423, new_P3_R1095_U424, new_P3_R1095_U425,
    new_P3_R1095_U426, new_P3_R1095_U427, new_P3_R1095_U428,
    new_P3_R1095_U429, new_P3_R1095_U430, new_P3_R1095_U431,
    new_P3_R1095_U432, new_P3_R1095_U433, new_P3_R1095_U434,
    new_P3_R1095_U435, new_P3_R1095_U436, new_P3_R1095_U437,
    new_P3_R1095_U438, new_P3_R1095_U439, new_P3_R1095_U440,
    new_P3_R1095_U441, new_P3_R1095_U442, new_P3_R1095_U443,
    new_P3_R1095_U444, new_P3_R1095_U445, new_P3_R1095_U446,
    new_P3_R1095_U447, new_P3_R1095_U448, new_P3_R1095_U449,
    new_P3_R1095_U450, new_P3_R1095_U451, new_P3_R1095_U452,
    new_P3_R1095_U453, new_P3_R1095_U454, new_P3_R1095_U455,
    new_P3_R1095_U456, new_P3_R1095_U457, new_P3_R1095_U458,
    new_P3_R1095_U459, new_P3_R1095_U460, new_P3_R1095_U461,
    new_P3_R1095_U462, new_P3_R1095_U463, new_P3_R1095_U464,
    new_P3_R1095_U465, new_P3_R1095_U466, new_P3_R1095_U467,
    new_P3_R1095_U468, new_P3_R1095_U469, new_P3_R1095_U470,
    new_P3_R1095_U471, new_P3_R1095_U472, new_P3_R1095_U473,
    new_P3_R1095_U474, new_P3_R1095_U475, new_P3_R1095_U476,
    new_P3_R1095_U477, new_P3_R1095_U478, new_P3_R1095_U479,
    new_P3_R1095_U480, new_P3_R1095_U481, new_P3_R1095_U482,
    new_P3_R1095_U483, new_P3_R1095_U484, new_P3_R1095_U485,
    new_P3_R1212_U6, new_P3_R1212_U7, new_P3_R1212_U8, new_P3_R1212_U9,
    new_P3_R1212_U10, new_P3_R1212_U11, new_P3_R1212_U12, new_P3_R1212_U13,
    new_P3_R1212_U14, new_P3_R1212_U15, new_P3_R1212_U16, new_P3_R1212_U17,
    new_P3_R1212_U18, new_P3_R1212_U19, new_P3_R1212_U20, new_P3_R1212_U21,
    new_P3_R1212_U22, new_P3_R1212_U23, new_P3_R1212_U24, new_P3_R1212_U25,
    new_P3_R1212_U26, new_P3_R1212_U27, new_P3_R1212_U28, new_P3_R1212_U29,
    new_P3_R1212_U30, new_P3_R1212_U31, new_P3_R1212_U32, new_P3_R1212_U33,
    new_P3_R1212_U34, new_P3_R1212_U35, new_P3_R1212_U36, new_P3_R1212_U37,
    new_P3_R1212_U38, new_P3_R1212_U39, new_P3_R1212_U40, new_P3_R1212_U41,
    new_P3_R1212_U42, new_P3_R1212_U43, new_P3_R1212_U44, new_P3_R1212_U45,
    new_P3_R1212_U46, new_P3_R1212_U47, new_P3_R1212_U48, new_P3_R1212_U49,
    new_P3_R1212_U50, new_P3_R1212_U51, new_P3_R1212_U52, new_P3_R1212_U53,
    new_P3_R1212_U54, new_P3_R1212_U55, new_P3_R1212_U56, new_P3_R1212_U57,
    new_P3_R1212_U58, new_P3_R1212_U59, new_P3_R1212_U60, new_P3_R1212_U61,
    new_P3_R1212_U62, new_P3_R1212_U63, new_P3_R1212_U64, new_P3_R1212_U65,
    new_P3_R1212_U66, new_P3_R1212_U67, new_P3_R1212_U68, new_P3_R1212_U69,
    new_P3_R1212_U70, new_P3_R1212_U71, new_P3_R1212_U72, new_P3_R1212_U73,
    new_P3_R1212_U74, new_P3_R1212_U75, new_P3_R1212_U76, new_P3_R1212_U77,
    new_P3_R1212_U78, new_P3_R1212_U79, new_P3_R1212_U80, new_P3_R1212_U81,
    new_P3_R1212_U82, new_P3_R1212_U83, new_P3_R1212_U84, new_P3_R1212_U85,
    new_P3_R1212_U86, new_P3_R1212_U87, new_P3_R1212_U88, new_P3_R1212_U89,
    new_P3_R1212_U90, new_P3_R1212_U91, new_P3_R1212_U92, new_P3_R1212_U93,
    new_P3_R1212_U94, new_P3_R1212_U95, new_P3_R1212_U96, new_P3_R1212_U97,
    new_P3_R1212_U98, new_P3_R1212_U99, new_P3_R1212_U100,
    new_P3_R1212_U101, new_P3_R1212_U102, new_P3_R1212_U103,
    new_P3_R1212_U104, new_P3_R1212_U105, new_P3_R1212_U106,
    new_P3_R1212_U107, new_P3_R1212_U108, new_P3_R1212_U109,
    new_P3_R1212_U110, new_P3_R1212_U111, new_P3_R1212_U112,
    new_P3_R1212_U113, new_P3_R1212_U114, new_P3_R1212_U115,
    new_P3_R1212_U116, new_P3_R1212_U117, new_P3_R1212_U118,
    new_P3_R1212_U119, new_P3_R1212_U120, new_P3_R1212_U121,
    new_P3_R1212_U122, new_P3_R1212_U123, new_P3_R1212_U124,
    new_P3_R1212_U125, new_P3_R1212_U126, new_P3_R1212_U127,
    new_P3_R1212_U128, new_P3_R1212_U129, new_P3_R1212_U130,
    new_P3_R1212_U131, new_P3_R1212_U132, new_P3_R1212_U133,
    new_P3_R1212_U134, new_P3_R1212_U135, new_P3_R1212_U136,
    new_P3_R1212_U137, new_P3_R1212_U138, new_P3_R1212_U139,
    new_P3_R1212_U140, new_P3_R1212_U141, new_P3_R1212_U142,
    new_P3_R1212_U143, new_P3_R1212_U144, new_P3_R1212_U145,
    new_P3_R1212_U146, new_P3_R1212_U147, new_P3_R1212_U148,
    new_P3_R1212_U149, new_P3_R1212_U150, new_P3_R1212_U151,
    new_P3_R1212_U152, new_P3_R1212_U153, new_P3_R1212_U154,
    new_P3_R1212_U155, new_P3_R1212_U156, new_P3_R1212_U157,
    new_P3_R1212_U158, new_P3_R1212_U159, new_P3_R1212_U160,
    new_P3_R1212_U161, new_P3_R1212_U162, new_P3_R1212_U163,
    new_P3_R1212_U164, new_P3_R1212_U165, new_P3_R1212_U166,
    new_P3_R1212_U167, new_P3_R1212_U168, new_P3_R1212_U169,
    new_P3_R1212_U170, new_P3_R1212_U171, new_P3_R1212_U172,
    new_P3_R1212_U173, new_P3_R1212_U174, new_P3_R1212_U175,
    new_P3_R1212_U176, new_P3_R1212_U177, new_P3_R1212_U178,
    new_P3_R1212_U179, new_P3_R1212_U180, new_P3_R1212_U181,
    new_P3_R1212_U182, new_P3_R1212_U183, new_P3_R1212_U184,
    new_P3_R1212_U185, new_P3_R1212_U186, new_P3_R1212_U187,
    new_P3_R1212_U188, new_P3_R1212_U189, new_P3_R1212_U190,
    new_P3_R1212_U191, new_P3_R1212_U192, new_P3_R1212_U193,
    new_P3_R1212_U194, new_P3_R1212_U195, new_P3_R1212_U196,
    new_P3_R1212_U197, new_P3_R1212_U198, new_P3_R1212_U199,
    new_P3_R1212_U200, new_P3_R1212_U201, new_P3_R1212_U202,
    new_P3_R1212_U203, new_P3_R1212_U204, new_P3_R1212_U205,
    new_P3_R1212_U206, new_P3_R1212_U207, new_P3_R1212_U208,
    new_P3_R1212_U209, new_P3_R1212_U210, new_P3_R1212_U211,
    new_P3_R1212_U212, new_P3_R1212_U213, new_P3_R1212_U214,
    new_P3_R1212_U215, new_P3_R1212_U216, new_P3_R1212_U217,
    new_P3_R1212_U218, new_P3_R1212_U219, new_P3_R1212_U220,
    new_P3_R1212_U221, new_P3_R1212_U222, new_P3_R1212_U223,
    new_P3_R1212_U224, new_P3_R1212_U225, new_P3_R1212_U226,
    new_P3_R1212_U227, new_P3_R1212_U228, new_P3_R1212_U229,
    new_P3_R1212_U230, new_P3_R1212_U231, new_P3_R1212_U232,
    new_P3_R1212_U233, new_P3_R1212_U234, new_P3_R1212_U235,
    new_P3_R1212_U236, new_P3_R1212_U237, new_P3_R1212_U238,
    new_P3_R1212_U239, new_P3_R1212_U240, new_P3_R1212_U241,
    new_P3_R1212_U242, new_P3_R1212_U243, new_P3_R1212_U244,
    new_P3_R1212_U245, new_P3_R1212_U246, new_P3_R1212_U247,
    new_P3_R1212_U248, new_P3_R1212_U249, new_P3_R1212_U250,
    new_P3_R1212_U251, new_P3_R1212_U252, new_P3_R1212_U253,
    new_P3_R1212_U254, new_P3_R1212_U255, new_P3_R1212_U256,
    new_P3_R1212_U257, new_P3_R1212_U258, new_P3_R1212_U259,
    new_P3_R1212_U260, new_P3_R1212_U261, new_P3_R1212_U262,
    new_P3_R1212_U263, new_P3_R1212_U264, new_P3_R1212_U265,
    new_P3_R1212_U266, new_P3_R1212_U267, new_P3_R1212_U268,
    new_P3_R1212_U269, new_P3_R1212_U270, new_P3_R1212_U271,
    new_P3_R1212_U272, new_P3_R1212_U273, new_P3_R1212_U274,
    new_P3_R1212_U275, new_P3_R1212_U276, new_P3_R1209_U6, new_P3_R1209_U7,
    new_P3_R1209_U8, new_P3_R1209_U9, new_P3_R1209_U10, new_P3_R1209_U11,
    new_P3_R1209_U12, new_P3_R1209_U13, new_P3_R1209_U14, new_P3_R1209_U15,
    new_P3_R1209_U16, new_P3_R1209_U17, new_P3_R1209_U18, new_P3_R1209_U19,
    new_P3_R1209_U20, new_P3_R1209_U21, new_P3_R1209_U22, new_P3_R1209_U23,
    new_P3_R1209_U24, new_P3_R1209_U25, new_P3_R1209_U26, new_P3_R1209_U27,
    new_P3_R1209_U28, new_P3_R1209_U29, new_P3_R1209_U30, new_P3_R1209_U31,
    new_P3_R1209_U32, new_P3_R1209_U33, new_P3_R1209_U34, new_P3_R1209_U35,
    new_P3_R1209_U36, new_P3_R1209_U37, new_P3_R1209_U38, new_P3_R1209_U39,
    new_P3_R1209_U40, new_P3_R1209_U41, new_P3_R1209_U42, new_P3_R1209_U43,
    new_P3_R1209_U44, new_P3_R1209_U45, new_P3_R1209_U46, new_P3_R1209_U47,
    new_P3_R1209_U48, new_P3_R1209_U49, new_P3_R1209_U50, new_P3_R1209_U51,
    new_P3_R1209_U52, new_P3_R1209_U53, new_P3_R1209_U54, new_P3_R1209_U55,
    new_P3_R1209_U56, new_P3_R1209_U57, new_P3_R1209_U58, new_P3_R1209_U59,
    new_P3_R1209_U60, new_P3_R1209_U61, new_P3_R1209_U62, new_P3_R1209_U63,
    new_P3_R1209_U64, new_P3_R1209_U65, new_P3_R1209_U66, new_P3_R1209_U67,
    new_P3_R1209_U68, new_P3_R1209_U69, new_P3_R1209_U70, new_P3_R1209_U71,
    new_P3_R1209_U72, new_P3_R1209_U73, new_P3_R1209_U74, new_P3_R1209_U75,
    new_P3_R1209_U76, new_P3_R1209_U77, new_P3_R1209_U78, new_P3_R1209_U79,
    new_P3_R1209_U80, new_P3_R1209_U81, new_P3_R1209_U82, new_P3_R1209_U83,
    new_P3_R1209_U84, new_P3_R1209_U85, new_P3_R1209_U86, new_P3_R1209_U87,
    new_P3_R1209_U88, new_P3_R1209_U89, new_P3_R1209_U90, new_P3_R1209_U91,
    new_P3_R1209_U92, new_P3_R1209_U93, new_P3_R1209_U94, new_P3_R1209_U95,
    new_P3_R1209_U96, new_P3_R1209_U97, new_P3_R1209_U98, new_P3_R1209_U99,
    new_P3_R1209_U100, new_P3_R1209_U101, new_P3_R1209_U102,
    new_P3_R1209_U103, new_P3_R1209_U104, new_P3_R1209_U105,
    new_P3_R1209_U106, new_P3_R1209_U107, new_P3_R1209_U108,
    new_P3_R1209_U109, new_P3_R1209_U110, new_P3_R1209_U111,
    new_P3_R1209_U112, new_P3_R1209_U113, new_P3_R1209_U114,
    new_P3_R1209_U115, new_P3_R1209_U116, new_P3_R1209_U117,
    new_P3_R1209_U118, new_P3_R1209_U119, new_P3_R1209_U120,
    new_P3_R1209_U121, new_P3_R1209_U122, new_P3_R1209_U123,
    new_P3_R1209_U124, new_P3_R1209_U125, new_P3_R1209_U126,
    new_P3_R1209_U127, new_P3_R1209_U128, new_P3_R1209_U129,
    new_P3_R1209_U130, new_P3_R1209_U131, new_P3_R1209_U132,
    new_P3_R1209_U133, new_P3_R1209_U134, new_P3_R1209_U135,
    new_P3_R1209_U136, new_P3_R1209_U137, new_P3_R1209_U138,
    new_P3_R1209_U139, new_P3_R1209_U140, new_P3_R1209_U141,
    new_P3_R1209_U142, new_P3_R1209_U143, new_P3_R1209_U144,
    new_P3_R1209_U145, new_P3_R1209_U146, new_P3_R1209_U147,
    new_P3_R1209_U148, new_P3_R1209_U149, new_P3_R1209_U150,
    new_P3_R1209_U151, new_P3_R1209_U152, new_P3_R1209_U153,
    new_P3_R1209_U154, new_P3_R1209_U155, new_P3_R1209_U156,
    new_P3_R1209_U157, new_P3_R1209_U158, new_P3_R1209_U159,
    new_P3_R1209_U160, new_P3_R1209_U161, new_P3_R1209_U162,
    new_P3_R1209_U163, new_P3_R1209_U164, new_P3_R1209_U165,
    new_P3_R1209_U166, new_P3_R1209_U167, new_P3_R1209_U168,
    new_P3_R1209_U169, new_P3_R1209_U170, new_P3_R1209_U171,
    new_P3_R1209_U172, new_P3_R1209_U173, new_P3_R1209_U174,
    new_P3_R1209_U175, new_P3_R1209_U176, new_P3_R1209_U177,
    new_P3_R1209_U178, new_P3_R1209_U179, new_P3_R1209_U180,
    new_P3_R1209_U181, new_P3_R1209_U182, new_P3_R1209_U183,
    new_P3_R1209_U184, new_P3_R1209_U185, new_P3_R1209_U186,
    new_P3_R1209_U187, new_P3_R1209_U188, new_P3_R1209_U189,
    new_P3_R1209_U190, new_P3_R1209_U191, new_P3_R1209_U192,
    new_P3_R1209_U193, new_P3_R1209_U194, new_P3_R1209_U195,
    new_P3_R1209_U196, new_P3_R1209_U197, new_P3_R1209_U198,
    new_P3_R1209_U199, new_P3_R1209_U200, new_P3_R1209_U201,
    new_P3_R1209_U202, new_P3_R1209_U203, new_P3_R1209_U204,
    new_P3_R1209_U205, new_P3_R1209_U206, new_P3_R1209_U207,
    new_P3_R1209_U208, new_P3_R1209_U209, new_P3_R1209_U210,
    new_P3_R1209_U211, new_P3_R1209_U212, new_P3_R1209_U213,
    new_P3_R1209_U214, new_P3_R1209_U215, new_P3_R1209_U216,
    new_P3_R1209_U217, new_P3_R1209_U218, new_P3_R1209_U219,
    new_P3_R1209_U220, new_P3_R1209_U221, new_P3_R1209_U222,
    new_P3_R1209_U223, new_P3_R1209_U224, new_P3_R1209_U225,
    new_P3_R1209_U226, new_P3_R1209_U227, new_P3_R1209_U228,
    new_P3_R1209_U229, new_P3_R1209_U230, new_P3_R1209_U231,
    new_P3_R1209_U232, new_P3_R1209_U233, new_P3_R1209_U234,
    new_P3_R1209_U235, new_P3_R1209_U236, new_P3_R1209_U237,
    new_P3_R1209_U238, new_P3_R1209_U239, new_P3_R1209_U240,
    new_P3_R1209_U241, new_P3_R1209_U242, new_P3_R1209_U243,
    new_P3_R1209_U244, new_P3_R1209_U245, new_P3_R1209_U246,
    new_P3_R1209_U247, new_P3_R1209_U248, new_P3_R1209_U249,
    new_P3_R1209_U250, new_P3_R1209_U251, new_P3_R1209_U252,
    new_P3_R1209_U253, new_P3_R1209_U254, new_P3_R1209_U255,
    new_P3_R1209_U256, new_P3_R1209_U257, new_P3_R1209_U258,
    new_P3_R1209_U259, new_P3_R1209_U260, new_P3_R1209_U261,
    new_P3_R1209_U262, new_P3_R1209_U263, new_P3_R1209_U264,
    new_P3_R1209_U265, new_P3_R1209_U266, new_P3_R1209_U267,
    new_P3_R1209_U268, new_P3_R1209_U269, new_P3_R1209_U270,
    new_P3_R1209_U271, new_P3_R1209_U272, new_P3_R1209_U273,
    new_P3_R1209_U274, new_P3_R1209_U275, new_P3_R1209_U276,
    new_P3_R1300_U6, new_P3_R1300_U7, new_P3_R1300_U8, new_P3_R1300_U9,
    new_P3_R1300_U10, new_P3_R1200_U6, new_P3_R1200_U7, new_P3_R1200_U8,
    new_P3_R1200_U9, new_P3_R1200_U10, new_P3_R1200_U11, new_P3_R1200_U12,
    new_P3_R1200_U13, new_P3_R1200_U14, new_P3_R1200_U15, new_P3_R1200_U16,
    new_P3_R1200_U17, new_P3_R1200_U18, new_P3_R1200_U19, new_P3_R1200_U20,
    new_P3_R1200_U21, new_P3_R1200_U22, new_P3_R1200_U23, new_P3_R1200_U24,
    new_P3_R1200_U25, new_P3_R1200_U26, new_P3_R1200_U27, new_P3_R1200_U28,
    new_P3_R1200_U29, new_P3_R1200_U30, new_P3_R1200_U31, new_P3_R1200_U32,
    new_P3_R1200_U33, new_P3_R1200_U34, new_P3_R1200_U35, new_P3_R1200_U36,
    new_P3_R1200_U37, new_P3_R1200_U38, new_P3_R1200_U39, new_P3_R1200_U40,
    new_P3_R1200_U41, new_P3_R1200_U42, new_P3_R1200_U43, new_P3_R1200_U44,
    new_P3_R1200_U45, new_P3_R1200_U46, new_P3_R1200_U47, new_P3_R1200_U48,
    new_P3_R1200_U49, new_P3_R1200_U50, new_P3_R1200_U51, new_P3_R1200_U52,
    new_P3_R1200_U53, new_P3_R1200_U54, new_P3_R1200_U55, new_P3_R1200_U56,
    new_P3_R1200_U57, new_P3_R1200_U58, new_P3_R1200_U59, new_P3_R1200_U60,
    new_P3_R1200_U61, new_P3_R1200_U62, new_P3_R1200_U63, new_P3_R1200_U64,
    new_P3_R1200_U65, new_P3_R1200_U66, new_P3_R1200_U67, new_P3_R1200_U68,
    new_P3_R1200_U69, new_P3_R1200_U70, new_P3_R1200_U71, new_P3_R1200_U72,
    new_P3_R1200_U73, new_P3_R1200_U74, new_P3_R1200_U75, new_P3_R1200_U76,
    new_P3_R1200_U77, new_P3_R1200_U78, new_P3_R1200_U79, new_P3_R1200_U80,
    new_P3_R1200_U81, new_P3_R1200_U82, new_P3_R1200_U83, new_P3_R1200_U84,
    new_P3_R1200_U85, new_P3_R1200_U86, new_P3_R1200_U87, new_P3_R1200_U88,
    new_P3_R1200_U89, new_P3_R1200_U90, new_P3_R1200_U91, new_P3_R1200_U92,
    new_P3_R1200_U93, new_P3_R1200_U94, new_P3_R1200_U95, new_P3_R1200_U96,
    new_P3_R1200_U97, new_P3_R1200_U98, new_P3_R1200_U99,
    new_P3_R1200_U100, new_P3_R1200_U101, new_P3_R1200_U102,
    new_P3_R1200_U103, new_P3_R1200_U104, new_P3_R1200_U105,
    new_P3_R1200_U106, new_P3_R1200_U107, new_P3_R1200_U108,
    new_P3_R1200_U109, new_P3_R1200_U110, new_P3_R1200_U111,
    new_P3_R1200_U112, new_P3_R1200_U113, new_P3_R1200_U114,
    new_P3_R1200_U115, new_P3_R1200_U116, new_P3_R1200_U117,
    new_P3_R1200_U118, new_P3_R1200_U119, new_P3_R1200_U120,
    new_P3_R1200_U121, new_P3_R1200_U122, new_P3_R1200_U123,
    new_P3_R1200_U124, new_P3_R1200_U125, new_P3_R1200_U126,
    new_P3_R1200_U127, new_P3_R1200_U128, new_P3_R1200_U129,
    new_P3_R1200_U130, new_P3_R1200_U131, new_P3_R1200_U132,
    new_P3_R1200_U133, new_P3_R1200_U134, new_P3_R1200_U135,
    new_P3_R1200_U136, new_P3_R1200_U137, new_P3_R1200_U138,
    new_P3_R1200_U139, new_P3_R1200_U140, new_P3_R1200_U141,
    new_P3_R1200_U142, new_P3_R1200_U143, new_P3_R1200_U144,
    new_P3_R1200_U145, new_P3_R1200_U146, new_P3_R1200_U147,
    new_P3_R1200_U148, new_P3_R1200_U149, new_P3_R1200_U150,
    new_P3_R1200_U151, new_P3_R1200_U152, new_P3_R1200_U153,
    new_P3_R1200_U154, new_P3_R1200_U155, new_P3_R1200_U156,
    new_P3_R1200_U157, new_P3_R1200_U158, new_P3_R1200_U159,
    new_P3_R1200_U160, new_P3_R1200_U161, new_P3_R1200_U162,
    new_P3_R1200_U163, new_P3_R1200_U164, new_P3_R1200_U165,
    new_P3_R1200_U166, new_P3_R1200_U167, new_P3_R1200_U168,
    new_P3_R1200_U169, new_P3_R1200_U170, new_P3_R1200_U171,
    new_P3_R1200_U172, new_P3_R1200_U173, new_P3_R1200_U174,
    new_P3_R1200_U175, new_P3_R1200_U176, new_P3_R1200_U177,
    new_P3_R1200_U178, new_P3_R1200_U179, new_P3_R1200_U180,
    new_P3_R1200_U181, new_P3_R1200_U182, new_P3_R1200_U183,
    new_P3_R1200_U184, new_P3_R1200_U185, new_P3_R1200_U186,
    new_P3_R1200_U187, new_P3_R1200_U188, new_P3_R1200_U189,
    new_P3_R1200_U190, new_P3_R1200_U191, new_P3_R1200_U192,
    new_P3_R1200_U193, new_P3_R1200_U194, new_P3_R1200_U195,
    new_P3_R1200_U196, new_P3_R1200_U197, new_P3_R1200_U198,
    new_P3_R1200_U199, new_P3_R1200_U200, new_P3_R1200_U201,
    new_P3_R1200_U202, new_P3_R1200_U203, new_P3_R1200_U204,
    new_P3_R1200_U205, new_P3_R1200_U206, new_P3_R1200_U207,
    new_P3_R1200_U208, new_P3_R1200_U209, new_P3_R1200_U210,
    new_P3_R1200_U211, new_P3_R1200_U212, new_P3_R1200_U213,
    new_P3_R1200_U214, new_P3_R1200_U215, new_P3_R1200_U216,
    new_P3_R1200_U217, new_P3_R1200_U218, new_P3_R1200_U219,
    new_P3_R1200_U220, new_P3_R1200_U221, new_P3_R1200_U222,
    new_P3_R1200_U223, new_P3_R1200_U224, new_P3_R1200_U225,
    new_P3_R1200_U226, new_P3_R1200_U227, new_P3_R1200_U228,
    new_P3_R1200_U229, new_P3_R1200_U230, new_P3_R1200_U231,
    new_P3_R1200_U232, new_P3_R1200_U233, new_P3_R1200_U234,
    new_P3_R1200_U235, new_P3_R1200_U236, new_P3_R1200_U237,
    new_P3_R1200_U238, new_P3_R1200_U239, new_P3_R1200_U240,
    new_P3_R1200_U241, new_P3_R1200_U242, new_P3_R1200_U243,
    new_P3_R1200_U244, new_P3_R1200_U245, new_P3_R1200_U246,
    new_P3_R1200_U247, new_P3_R1200_U248, new_P3_R1200_U249,
    new_P3_R1200_U250, new_P3_R1200_U251, new_P3_R1200_U252,
    new_P3_R1200_U253, new_P3_R1200_U254, new_P3_R1200_U255,
    new_P3_R1200_U256, new_P3_R1200_U257, new_P3_R1200_U258,
    new_P3_R1200_U259, new_P3_R1200_U260, new_P3_R1200_U261,
    new_P3_R1200_U262, new_P3_R1200_U263, new_P3_R1200_U264,
    new_P3_R1200_U265, new_P3_R1200_U266, new_P3_R1200_U267,
    new_P3_R1200_U268, new_P3_R1200_U269, new_P3_R1200_U270,
    new_P3_R1200_U271, new_P3_R1200_U272, new_P3_R1200_U273,
    new_P3_R1200_U274, new_P3_R1200_U275, new_P3_R1200_U276,
    new_P3_R1200_U277, new_P3_R1200_U278, new_P3_R1200_U279,
    new_P3_R1200_U280, new_P3_R1200_U281, new_P3_R1200_U282,
    new_P3_R1200_U283, new_P3_R1200_U284, new_P3_R1200_U285,
    new_P3_R1200_U286, new_P3_R1200_U287, new_P3_R1200_U288,
    new_P3_R1200_U289, new_P3_R1200_U290, new_P3_R1200_U291,
    new_P3_R1200_U292, new_P3_R1200_U293, new_P3_R1200_U294,
    new_P3_R1200_U295, new_P3_R1200_U296, new_P3_R1200_U297,
    new_P3_R1200_U298, new_P3_R1200_U299, new_P3_R1200_U300,
    new_P3_R1200_U301, new_P3_R1200_U302, new_P3_R1200_U303,
    new_P3_R1200_U304, new_P3_R1200_U305, new_P3_R1200_U306,
    new_P3_R1200_U307, new_P3_R1200_U308, new_P3_R1200_U309,
    new_P3_R1200_U310, new_P3_R1200_U311, new_P3_R1200_U312,
    new_P3_R1200_U313, new_P3_R1200_U314, new_P3_R1200_U315,
    new_P3_R1200_U316, new_P3_R1200_U317, new_P3_R1200_U318,
    new_P3_R1200_U319, new_P3_R1200_U320, new_P3_R1200_U321,
    new_P3_R1200_U322, new_P3_R1200_U323, new_P3_R1200_U324,
    new_P3_R1200_U325, new_P3_R1200_U326, new_P3_R1200_U327,
    new_P3_R1200_U328, new_P3_R1200_U329, new_P3_R1200_U330,
    new_P3_R1200_U331, new_P3_R1200_U332, new_P3_R1200_U333,
    new_P3_R1200_U334, new_P3_R1200_U335, new_P3_R1200_U336,
    new_P3_R1200_U337, new_P3_R1200_U338, new_P3_R1200_U339,
    new_P3_R1200_U340, new_P3_R1200_U341, new_P3_R1200_U342,
    new_P3_R1200_U343, new_P3_R1200_U344, new_P3_R1200_U345,
    new_P3_R1200_U346, new_P3_R1200_U347, new_P3_R1200_U348,
    new_P3_R1200_U349, new_P3_R1200_U350, new_P3_R1200_U351,
    new_P3_R1200_U352, new_P3_R1200_U353, new_P3_R1200_U354,
    new_P3_R1200_U355, new_P3_R1200_U356, new_P3_R1200_U357,
    new_P3_R1200_U358, new_P3_R1200_U359, new_P3_R1200_U360,
    new_P3_R1200_U361, new_P3_R1200_U362, new_P3_R1200_U363,
    new_P3_R1200_U364, new_P3_R1200_U365, new_P3_R1200_U366,
    new_P3_R1200_U367, new_P3_R1200_U368, new_P3_R1200_U369,
    new_P3_R1200_U370, new_P3_R1200_U371, new_P3_R1200_U372,
    new_P3_R1200_U373, new_P3_R1200_U374, new_P3_R1200_U375,
    new_P3_R1200_U376, new_P3_R1200_U377, new_P3_R1200_U378,
    new_P3_R1200_U379, new_P3_R1200_U380, new_P3_R1200_U381,
    new_P3_R1200_U382, new_P3_R1200_U383, new_P3_R1200_U384,
    new_P3_R1200_U385, new_P3_R1200_U386, new_P3_R1200_U387,
    new_P3_R1200_U388, new_P3_R1200_U389, new_P3_R1200_U390,
    new_P3_R1200_U391, new_P3_R1200_U392, new_P3_R1200_U393,
    new_P3_R1200_U394, new_P3_R1200_U395, new_P3_R1200_U396,
    new_P3_R1200_U397, new_P3_R1200_U398, new_P3_R1200_U399,
    new_P3_R1200_U400, new_P3_R1200_U401, new_P3_R1200_U402,
    new_P3_R1200_U403, new_P3_R1200_U404, new_P3_R1200_U405,
    new_P3_R1200_U406, new_P3_R1200_U407, new_P3_R1200_U408,
    new_P3_R1200_U409, new_P3_R1200_U410, new_P3_R1200_U411,
    new_P3_R1200_U412, new_P3_R1200_U413, new_P3_R1200_U414,
    new_P3_R1200_U415, new_P3_R1200_U416, new_P3_R1200_U417,
    new_P3_R1200_U418, new_P3_R1200_U419, new_P3_R1200_U420,
    new_P3_R1200_U421, new_P3_R1200_U422, new_P3_R1200_U423,
    new_P3_R1200_U424, new_P3_R1200_U425, new_P3_R1200_U426,
    new_P3_R1200_U427, new_P3_R1200_U428, new_P3_R1200_U429,
    new_P3_R1200_U430, new_P3_R1200_U431, new_P3_R1200_U432,
    new_P3_R1200_U433, new_P3_R1200_U434, new_P3_R1200_U435,
    new_P3_R1200_U436, new_P3_R1200_U437, new_P3_R1200_U438,
    new_P3_R1200_U439, new_P3_R1200_U440, new_P3_R1200_U441,
    new_P3_R1200_U442, new_P3_R1200_U443, new_P3_R1200_U444,
    new_P3_R1200_U445, new_P3_R1200_U446, new_P3_R1200_U447,
    new_P3_R1200_U448, new_P3_R1200_U449, new_P3_R1200_U450,
    new_P3_R1200_U451, new_P3_R1200_U452, new_P3_R1200_U453,
    new_P3_R1200_U454, new_P3_R1200_U455, new_P3_R1200_U456,
    new_P3_R1200_U457, new_P3_R1200_U458, new_P3_R1200_U459,
    new_P3_R1200_U460, new_P3_R1200_U461, new_P3_R1200_U462,
    new_P3_R1200_U463, new_P3_R1200_U464, new_P3_R1200_U465,
    new_P3_R1200_U466, new_P3_R1200_U467, new_P3_R1200_U468,
    new_P3_R1200_U469, new_P3_R1200_U470, new_P3_R1200_U471,
    new_P3_R1200_U472, new_P3_R1200_U473, new_P3_R1200_U474,
    new_P3_R1200_U475, new_P3_R1200_U476, new_P3_R1200_U477,
    new_P3_R1200_U478, new_P3_R1200_U479, new_P3_R1200_U480,
    new_P3_R1200_U481, new_P3_R1200_U482, new_P3_R1200_U483,
    new_P3_R1200_U484, new_P3_R1200_U485, new_P3_R1179_U6, new_P3_R1179_U7,
    new_P3_R1179_U8, new_P3_R1179_U9, new_P3_R1179_U10, new_P3_R1179_U11,
    new_P3_R1179_U12, new_P3_R1179_U13, new_P3_R1179_U14, new_P3_R1179_U15,
    new_P3_R1179_U16, new_P3_R1179_U17, new_P3_R1179_U18, new_P3_R1179_U19,
    new_P3_R1179_U20, new_P3_R1179_U21, new_P3_R1179_U22, new_P3_R1179_U23,
    new_P3_R1179_U24, new_P3_R1179_U25, new_P3_R1179_U26, new_P3_R1179_U27,
    new_P3_R1179_U28, new_P3_R1179_U29, new_P3_R1179_U30, new_P3_R1179_U31,
    new_P3_R1179_U32, new_P3_R1179_U33, new_P3_R1179_U34, new_P3_R1179_U35,
    new_P3_R1179_U36, new_P3_R1179_U37, new_P3_R1179_U38, new_P3_R1179_U39,
    new_P3_R1179_U40, new_P3_R1179_U41, new_P3_R1179_U42, new_P3_R1179_U43,
    new_P3_R1179_U44, new_P3_R1179_U45, new_P3_R1179_U46, new_P3_R1179_U47,
    new_P3_R1179_U48, new_P3_R1179_U49, new_P3_R1179_U50, new_P3_R1179_U51,
    new_P3_R1179_U52, new_P3_R1179_U53, new_P3_R1179_U54, new_P3_R1179_U55,
    new_P3_R1179_U56, new_P3_R1179_U57, new_P3_R1179_U58, new_P3_R1179_U59,
    new_P3_R1179_U60, new_P3_R1179_U61, new_P3_R1179_U62, new_P3_R1179_U63,
    new_P3_R1179_U64, new_P3_R1179_U65, new_P3_R1179_U66, new_P3_R1179_U67,
    new_P3_R1179_U68, new_P3_R1179_U69, new_P3_R1179_U70, new_P3_R1179_U71,
    new_P3_R1179_U72, new_P3_R1179_U73, new_P3_R1179_U74, new_P3_R1179_U75,
    new_P3_R1179_U76, new_P3_R1179_U77, new_P3_R1179_U78, new_P3_R1179_U79,
    new_P3_R1179_U80, new_P3_R1179_U81, new_P3_R1179_U82, new_P3_R1179_U83,
    new_P3_R1179_U84, new_P3_R1179_U85, new_P3_R1179_U86, new_P3_R1179_U87,
    new_P3_R1179_U88, new_P3_R1179_U89, new_P3_R1179_U90, new_P3_R1179_U91,
    new_P3_R1179_U92, new_P3_R1179_U93, new_P3_R1179_U94, new_P3_R1179_U95,
    new_P3_R1179_U96, new_P3_R1179_U97, new_P3_R1179_U98, new_P3_R1179_U99,
    new_P3_R1179_U100, new_P3_R1179_U101, new_P3_R1179_U102,
    new_P3_R1179_U103, new_P3_R1179_U104, new_P3_R1179_U105,
    new_P3_R1179_U106, new_P3_R1179_U107, new_P3_R1179_U108,
    new_P3_R1179_U109, new_P3_R1179_U110, new_P3_R1179_U111,
    new_P3_R1179_U112, new_P3_R1179_U113, new_P3_R1179_U114,
    new_P3_R1179_U115, new_P3_R1179_U116, new_P3_R1179_U117,
    new_P3_R1179_U118, new_P3_R1179_U119, new_P3_R1179_U120,
    new_P3_R1179_U121, new_P3_R1179_U122, new_P3_R1179_U123,
    new_P3_R1179_U124, new_P3_R1179_U125, new_P3_R1179_U126,
    new_P3_R1179_U127, new_P3_R1179_U128, new_P3_R1179_U129,
    new_P3_R1179_U130, new_P3_R1179_U131, new_P3_R1179_U132,
    new_P3_R1179_U133, new_P3_R1179_U134, new_P3_R1179_U135,
    new_P3_R1179_U136, new_P3_R1179_U137, new_P3_R1179_U138,
    new_P3_R1179_U139, new_P3_R1179_U140, new_P3_R1179_U141,
    new_P3_R1179_U142, new_P3_R1179_U143, new_P3_R1179_U144,
    new_P3_R1179_U145, new_P3_R1179_U146, new_P3_R1179_U147,
    new_P3_R1179_U148, new_P3_R1179_U149, new_P3_R1179_U150,
    new_P3_R1179_U151, new_P3_R1179_U152, new_P3_R1179_U153,
    new_P3_R1179_U154, new_P3_R1179_U155, new_P3_R1179_U156,
    new_P3_R1179_U157, new_P3_R1179_U158, new_P3_R1179_U159,
    new_P3_R1179_U160, new_P3_R1179_U161, new_P3_R1179_U162,
    new_P3_R1179_U163, new_P3_R1179_U164, new_P3_R1179_U165,
    new_P3_R1179_U166, new_P3_R1179_U167, new_P3_R1179_U168,
    new_P3_R1179_U169, new_P3_R1179_U170, new_P3_R1179_U171,
    new_P3_R1179_U172, new_P3_R1179_U173, new_P3_R1179_U174,
    new_P3_R1179_U175, new_P3_R1179_U176, new_P3_R1179_U177,
    new_P3_R1179_U178, new_P3_R1179_U179, new_P3_R1179_U180,
    new_P3_R1179_U181, new_P3_R1179_U182, new_P3_R1179_U183,
    new_P3_R1179_U184, new_P3_R1179_U185, new_P3_R1179_U186,
    new_P3_R1179_U187, new_P3_R1179_U188, new_P3_R1179_U189,
    new_P3_R1179_U190, new_P3_R1179_U191, new_P3_R1179_U192,
    new_P3_R1179_U193, new_P3_R1179_U194, new_P3_R1179_U195,
    new_P3_R1179_U196, new_P3_R1179_U197, new_P3_R1179_U198,
    new_P3_R1179_U199, new_P3_R1179_U200, new_P3_R1179_U201,
    new_P3_R1179_U202, new_P3_R1179_U203, new_P3_R1179_U204,
    new_P3_R1179_U205, new_P3_R1179_U206, new_P3_R1179_U207,
    new_P3_R1179_U208, new_P3_R1179_U209, new_P3_R1179_U210,
    new_P3_R1179_U211, new_P3_R1179_U212, new_P3_R1179_U213,
    new_P3_R1179_U214, new_P3_R1179_U215, new_P3_R1179_U216,
    new_P3_R1179_U217, new_P3_R1179_U218, new_P3_R1179_U219,
    new_P3_R1179_U220, new_P3_R1179_U221, new_P3_R1179_U222,
    new_P3_R1179_U223, new_P3_R1179_U224, new_P3_R1179_U225,
    new_P3_R1179_U226, new_P3_R1179_U227, new_P3_R1179_U228,
    new_P3_R1179_U229, new_P3_R1179_U230, new_P3_R1179_U231,
    new_P3_R1179_U232, new_P3_R1179_U233, new_P3_R1179_U234,
    new_P3_R1179_U235, new_P3_R1179_U236, new_P3_R1179_U237,
    new_P3_R1179_U238, new_P3_R1179_U239, new_P3_R1179_U240,
    new_P3_R1179_U241, new_P3_R1179_U242, new_P3_R1179_U243,
    new_P3_R1179_U244, new_P3_R1179_U245, new_P3_R1179_U246,
    new_P3_R1179_U247, new_P3_R1179_U248, new_P3_R1179_U249,
    new_P3_R1179_U250, new_P3_R1179_U251, new_P3_R1179_U252,
    new_P3_R1179_U253, new_P3_R1179_U254, new_P3_R1179_U255,
    new_P3_R1179_U256, new_P3_R1179_U257, new_P3_R1179_U258,
    new_P3_R1179_U259, new_P3_R1179_U260, new_P3_R1179_U261,
    new_P3_R1179_U262, new_P3_R1179_U263, new_P3_R1179_U264,
    new_P3_R1179_U265, new_P3_R1179_U266, new_P3_R1179_U267,
    new_P3_R1179_U268, new_P3_R1179_U269, new_P3_R1179_U270,
    new_P3_R1179_U271, new_P3_R1179_U272, new_P3_R1179_U273,
    new_P3_R1179_U274, new_P3_R1179_U275, new_P3_R1179_U276,
    new_P3_R1179_U277, new_P3_R1179_U278, new_P3_R1179_U279,
    new_P3_R1179_U280, new_P3_R1179_U281, new_P3_R1179_U282,
    new_P3_R1179_U283, new_P3_R1179_U284, new_P3_R1179_U285,
    new_P3_R1179_U286, new_P3_R1179_U287, new_P3_R1179_U288,
    new_P3_R1179_U289, new_P3_R1179_U290, new_P3_R1179_U291,
    new_P3_R1179_U292, new_P3_R1179_U293, new_P3_R1179_U294,
    new_P3_R1179_U295, new_P3_R1179_U296, new_P3_R1179_U297,
    new_P3_R1179_U298, new_P3_R1179_U299, new_P3_R1179_U300,
    new_P3_R1179_U301, new_P3_R1179_U302, new_P3_R1179_U303,
    new_P3_R1179_U304, new_P3_R1179_U305, new_P3_R1179_U306,
    new_P3_R1179_U307, new_P3_R1179_U308, new_P3_R1179_U309,
    new_P3_R1179_U310, new_P3_R1179_U311, new_P3_R1179_U312,
    new_P3_R1179_U313, new_P3_R1179_U314, new_P3_R1179_U315,
    new_P3_R1179_U316, new_P3_R1179_U317, new_P3_R1179_U318,
    new_P3_R1179_U319, new_P3_R1179_U320, new_P3_R1179_U321,
    new_P3_R1179_U322, new_P3_R1179_U323, new_P3_R1179_U324,
    new_P3_R1179_U325, new_P3_R1179_U326, new_P3_R1179_U327,
    new_P3_R1179_U328, new_P3_R1179_U329, new_P3_R1179_U330,
    new_P3_R1179_U331, new_P3_R1179_U332, new_P3_R1179_U333,
    new_P3_R1179_U334, new_P3_R1179_U335, new_P3_R1179_U336,
    new_P3_R1179_U337, new_P3_R1179_U338, new_P3_R1179_U339,
    new_P3_R1179_U340, new_P3_R1179_U341, new_P3_R1179_U342,
    new_P3_R1179_U343, new_P3_R1179_U344, new_P3_R1179_U345,
    new_P3_R1179_U346, new_P3_R1179_U347, new_P3_R1179_U348,
    new_P3_R1179_U349, new_P3_R1179_U350, new_P3_R1179_U351,
    new_P3_R1179_U352, new_P3_R1179_U353, new_P3_R1179_U354,
    new_P3_R1179_U355, new_P3_R1179_U356, new_P3_R1179_U357,
    new_P3_R1179_U358, new_P3_R1179_U359, new_P3_R1179_U360,
    new_P3_R1179_U361, new_P3_R1179_U362, new_P3_R1179_U363,
    new_P3_R1179_U364, new_P3_R1179_U365, new_P3_R1179_U366,
    new_P3_R1179_U367, new_P3_R1179_U368, new_P3_R1179_U369,
    new_P3_R1179_U370, new_P3_R1179_U371, new_P3_R1179_U372,
    new_P3_R1179_U373, new_P3_R1179_U374, new_P3_R1179_U375,
    new_P3_R1179_U376, new_P3_R1179_U377, new_P3_R1179_U378,
    new_P3_R1179_U379, new_P3_R1179_U380, new_P3_R1179_U381,
    new_P3_R1179_U382, new_P3_R1179_U383, new_P3_R1179_U384,
    new_P3_R1179_U385, new_P3_R1179_U386, new_P3_R1179_U387,
    new_P3_R1179_U388, new_P3_R1179_U389, new_P3_R1179_U390,
    new_P3_R1179_U391, new_P3_R1179_U392, new_P3_R1179_U393,
    new_P3_R1179_U394, new_P3_R1179_U395, new_P3_R1179_U396,
    new_P3_R1179_U397, new_P3_R1179_U398, new_P3_R1179_U399,
    new_P3_R1179_U400, new_P3_R1179_U401, new_P3_R1179_U402,
    new_P3_R1179_U403, new_P3_R1179_U404, new_P3_R1179_U405,
    new_P3_R1179_U406, new_P3_R1179_U407, new_P3_R1179_U408,
    new_P3_R1179_U409, new_P3_R1179_U410, new_P3_R1179_U411,
    new_P3_R1179_U412, new_P3_R1179_U413, new_P3_R1179_U414,
    new_P3_R1179_U415, new_P3_R1179_U416, new_P3_R1179_U417,
    new_P3_R1179_U418, new_P3_R1179_U419, new_P3_R1179_U420,
    new_P3_R1179_U421, new_P3_R1179_U422, new_P3_R1179_U423,
    new_P3_R1179_U424, new_P3_R1179_U425, new_P3_R1179_U426,
    new_P3_R1179_U427, new_P3_R1179_U428, new_P3_R1179_U429,
    new_P3_R1179_U430, new_P3_R1179_U431, new_P3_R1179_U432,
    new_P3_R1179_U433, new_P3_R1179_U434, new_P3_R1179_U435,
    new_P3_R1179_U436, new_P3_R1179_U437, new_P3_R1179_U438,
    new_P3_R1179_U439, new_P3_R1179_U440, new_P3_R1179_U441,
    new_P3_R1179_U442, new_P3_R1179_U443, new_P3_R1179_U444,
    new_P3_R1179_U445, new_P3_R1179_U446, new_P3_R1179_U447,
    new_P3_R1179_U448, new_P3_R1179_U449, new_P3_R1179_U450,
    new_P3_R1179_U451, new_P3_R1179_U452, new_P3_R1179_U453,
    new_P3_R1179_U454, new_P3_R1179_U455, new_P3_R1179_U456,
    new_P3_R1179_U457, new_P3_R1179_U458, new_P3_R1179_U459,
    new_P3_R1179_U460, new_P3_R1179_U461, new_P3_R1179_U462,
    new_P3_R1179_U463, new_P3_R1179_U464, new_P3_R1179_U465,
    new_P3_R1179_U466, new_P3_R1179_U467, new_P3_R1179_U468,
    new_P3_R1179_U469, new_P3_R1179_U470, new_P3_R1179_U471,
    new_P3_R1179_U472, new_P3_R1179_U473, new_P3_R1179_U474,
    new_P3_R1179_U475, new_P3_R1179_U476, new_P3_R1179_U477,
    new_P3_R1179_U478, new_P3_R1179_U479, new_P3_R1179_U480,
    new_P3_R1179_U481, new_P3_R1179_U482, new_P3_R1179_U483,
    new_P3_R1179_U484, new_P3_R1179_U485, new_P3_R1269_U6, new_P3_R1269_U7,
    new_P3_R1269_U8, new_P3_R1269_U9, new_P3_R1269_U10, new_P3_R1269_U11,
    new_P3_R1269_U12, new_P3_R1269_U13, new_P3_R1269_U14, new_P3_R1269_U15,
    new_P3_R1269_U16, new_P3_R1269_U17, new_P3_R1269_U18, new_P3_R1269_U19,
    new_P3_R1269_U20, new_P3_R1269_U21, new_P3_R1269_U22, new_P3_R1269_U23,
    new_P3_R1269_U24, new_P3_R1269_U25, new_P3_R1269_U26, new_P3_R1269_U27,
    new_P3_R1269_U28, new_P3_R1269_U29, new_P3_R1269_U30, new_P3_R1269_U31,
    new_P3_R1269_U32, new_P3_R1269_U33, new_P3_R1269_U34, new_P3_R1269_U35,
    new_P3_R1269_U36, new_P3_R1269_U37, new_P3_R1269_U38, new_P3_R1269_U39,
    new_P3_R1269_U40, new_P3_R1269_U41, new_P3_R1269_U42, new_P3_R1269_U43,
    new_P3_R1269_U44, new_P3_R1269_U45, new_P3_R1269_U46, new_P3_R1269_U47,
    new_P3_R1269_U48, new_P3_R1269_U49, new_P3_R1269_U50, new_P3_R1269_U51,
    new_P3_R1269_U52, new_P3_R1269_U53, new_P3_R1269_U54, new_P3_R1269_U55,
    new_P3_R1269_U56, new_P3_R1269_U57, new_P3_R1269_U58, new_P3_R1269_U59,
    new_P3_R1269_U60, new_P3_R1269_U61, new_P3_R1269_U62, new_P3_R1269_U63,
    new_P3_R1269_U64, new_P3_R1269_U65, new_P3_R1269_U66, new_P3_R1269_U67,
    new_P3_R1269_U68, new_P3_R1269_U69, new_P3_R1269_U70, new_P3_R1269_U71,
    new_P3_R1269_U72, new_P3_R1269_U73, new_P3_R1269_U74, new_P3_R1269_U75,
    new_P3_R1269_U76, new_P3_R1269_U77, new_P3_R1269_U78, new_P3_R1269_U79,
    new_P3_R1269_U80, new_P3_R1269_U81, new_P3_R1269_U82, new_P3_R1269_U83,
    new_P3_R1269_U84, new_P3_R1269_U85, new_P3_R1269_U86, new_P3_R1269_U87,
    new_P3_R1269_U88, new_P3_R1269_U89, new_P3_R1269_U90, new_P3_R1269_U91,
    new_P3_R1269_U92, new_P3_R1269_U93, new_P3_R1269_U94, new_P3_R1269_U95,
    new_P3_R1269_U96, new_P3_R1269_U97, new_P3_R1269_U98, new_P3_R1269_U99,
    new_P3_R1269_U100, new_P3_R1269_U101, new_P3_R1269_U102,
    new_P3_R1269_U103, new_P3_R1269_U104, new_P3_R1269_U105,
    new_P3_R1269_U106, new_P3_R1269_U107, new_P3_R1269_U108,
    new_P3_R1269_U109, new_P3_R1269_U110, new_P3_R1269_U111,
    new_P3_R1269_U112, new_P3_R1269_U113, new_P3_R1269_U114,
    new_P3_R1269_U115, new_P3_R1269_U116, new_P3_R1269_U117,
    new_P3_R1269_U118, new_P3_R1269_U119, new_P3_R1269_U120,
    new_P3_R1269_U121, new_P3_R1269_U122, new_P3_R1269_U123,
    new_P3_R1269_U124, new_P3_R1269_U125, new_P3_R1269_U126,
    new_P3_R1269_U127, new_P3_R1269_U128, new_P3_R1269_U129,
    new_P3_R1269_U130, new_P3_R1269_U131, new_P3_R1269_U132,
    new_P3_R1269_U133, new_P3_R1269_U134, new_P3_R1269_U135,
    new_P3_R1269_U136, new_P3_R1269_U137, new_P3_R1269_U138,
    new_P3_R1269_U139, new_P3_R1269_U140, new_P3_R1269_U141,
    new_P3_R1269_U142, new_P3_R1269_U143, new_P3_R1269_U144,
    new_P3_R1269_U145, new_P3_R1269_U146, new_P3_R1269_U147,
    new_P3_R1269_U148, new_P3_R1269_U149, new_P3_R1269_U150,
    new_P3_R1269_U151, new_P3_R1269_U152, new_P3_R1269_U153,
    new_P3_R1269_U154, new_P3_R1269_U155, new_P3_R1269_U156,
    new_P3_R1269_U157, new_P3_R1269_U158, new_P3_R1269_U159,
    new_P3_R1269_U160, new_P3_R1269_U161, new_P3_R1269_U162,
    new_P3_R1269_U163, new_P3_R1269_U164, new_P3_R1269_U165,
    new_P3_R1269_U166, new_P3_R1269_U167, new_P3_R1269_U168,
    new_P3_R1269_U169, new_P3_R1269_U170, new_P3_R1269_U171,
    new_P3_R1269_U172, new_P3_R1269_U173, new_P3_R1269_U174,
    new_P3_R1269_U175, new_P3_R1269_U176, new_P3_R1269_U177,
    new_P3_R1269_U178, new_P3_R1269_U179, new_P3_R1269_U180,
    new_P3_R1269_U181, new_P3_R1269_U182, new_P3_R1269_U183,
    new_P3_R1269_U184, new_P3_R1269_U185, new_P3_R1269_U186,
    new_P3_R1269_U187, new_P3_R1269_U188, new_P3_R1269_U189,
    new_P3_R1269_U190, new_P3_R1269_U191, new_P3_R1269_U192,
    new_P3_R1269_U193, new_P3_R1269_U194, new_P3_R1269_U195,
    new_P3_R1269_U196, new_P3_R1269_U197, new_P3_R1269_U198,
    new_P3_R1269_U199, new_P3_R1269_U200, new_P3_R1269_U201,
    new_P3_R1269_U202, new_P3_R1110_U4, new_P3_R1110_U5, new_P3_R1110_U6,
    new_P3_R1110_U7, new_P3_R1110_U8, new_P3_R1110_U9, new_P3_R1110_U10,
    new_P3_R1110_U11, new_P3_R1110_U12, new_P3_R1110_U13, new_P3_R1110_U14,
    new_P3_R1110_U15, new_P3_R1110_U16, new_P3_R1110_U17, new_P3_R1110_U18,
    new_P3_R1110_U19, new_P3_R1110_U20, new_P3_R1110_U21, new_P3_R1110_U22,
    new_P3_R1110_U23, new_P3_R1110_U24, new_P3_R1110_U25, new_P3_R1110_U26,
    new_P3_R1110_U27, new_P3_R1110_U28, new_P3_R1110_U29, new_P3_R1110_U30,
    new_P3_R1110_U31, new_P3_R1110_U32, new_P3_R1110_U33, new_P3_R1110_U34,
    new_P3_R1110_U35, new_P3_R1110_U36, new_P3_R1110_U37, new_P3_R1110_U38,
    new_P3_R1110_U39, new_P3_R1110_U40, new_P3_R1110_U41, new_P3_R1110_U42,
    new_P3_R1110_U43, new_P3_R1110_U44, new_P3_R1110_U45, new_P3_R1110_U46,
    new_P3_R1110_U47, new_P3_R1110_U48, new_P3_R1110_U49, new_P3_R1110_U50,
    new_P3_R1110_U51, new_P3_R1110_U52, new_P3_R1110_U53, new_P3_R1110_U54,
    new_P3_R1110_U55, new_P3_R1110_U56, new_P3_R1110_U57, new_P3_R1110_U58,
    new_P3_R1110_U59, new_P3_R1110_U60, new_P3_R1110_U61, new_P3_R1110_U62,
    new_P3_R1110_U63, new_P3_R1110_U64, new_P3_R1110_U65, new_P3_R1110_U66,
    new_P3_R1110_U67, new_P3_R1110_U68, new_P3_R1110_U69, new_P3_R1110_U70,
    new_P3_R1110_U71, new_P3_R1110_U72, new_P3_R1110_U73, new_P3_R1110_U74,
    new_P3_R1110_U75, new_P3_R1110_U76, new_P3_R1110_U77, new_P3_R1110_U78,
    new_P3_R1110_U79, new_P3_R1110_U80, new_P3_R1110_U81, new_P3_R1110_U82,
    new_P3_R1110_U83, new_P3_R1110_U84, new_P3_R1110_U85, new_P3_R1110_U86,
    new_P3_R1110_U87, new_P3_R1110_U88, new_P3_R1110_U89, new_P3_R1110_U90,
    new_P3_R1110_U91, new_P3_R1110_U92, new_P3_R1110_U93, new_P3_R1110_U94,
    new_P3_R1110_U95, new_P3_R1110_U96, new_P3_R1110_U97, new_P3_R1110_U98,
    new_P3_R1110_U99, new_P3_R1110_U100, new_P3_R1110_U101,
    new_P3_R1110_U102, new_P3_R1110_U103, new_P3_R1110_U104,
    new_P3_R1110_U105, new_P3_R1110_U106, new_P3_R1110_U107,
    new_P3_R1110_U108, new_P3_R1110_U109, new_P3_R1110_U110,
    new_P3_R1110_U111, new_P3_R1110_U112, new_P3_R1110_U113,
    new_P3_R1110_U114, new_P3_R1110_U115, new_P3_R1110_U116,
    new_P3_R1110_U117, new_P3_R1110_U118, new_P3_R1110_U119,
    new_P3_R1110_U120, new_P3_R1110_U121, new_P3_R1110_U122,
    new_P3_R1110_U123, new_P3_R1110_U124, new_P3_R1110_U125,
    new_P3_R1110_U126, new_P3_R1110_U127, new_P3_R1110_U128,
    new_P3_R1110_U129, new_P3_R1110_U130, new_P3_R1110_U131,
    new_P3_R1110_U132, new_P3_R1110_U133, new_P3_R1110_U134,
    new_P3_R1110_U135, new_P3_R1110_U136, new_P3_R1110_U137,
    new_P3_R1110_U138, new_P3_R1110_U139, new_P3_R1110_U140,
    new_P3_R1110_U141, new_P3_R1110_U142, new_P3_R1110_U143,
    new_P3_R1110_U144, new_P3_R1110_U145, new_P3_R1110_U146,
    new_P3_R1110_U147, new_P3_R1110_U148, new_P3_R1110_U149,
    new_P3_R1110_U150, new_P3_R1110_U151, new_P3_R1110_U152,
    new_P3_R1110_U153, new_P3_R1110_U154, new_P3_R1110_U155,
    new_P3_R1110_U156, new_P3_R1110_U157, new_P3_R1110_U158,
    new_P3_R1110_U159, new_P3_R1110_U160, new_P3_R1110_U161,
    new_P3_R1110_U162, new_P3_R1110_U163, new_P3_R1110_U164,
    new_P3_R1110_U165, new_P3_R1110_U166, new_P3_R1110_U167,
    new_P3_R1110_U168, new_P3_R1110_U169, new_P3_R1110_U170,
    new_P3_R1110_U171, new_P3_R1110_U172, new_P3_R1110_U173,
    new_P3_R1110_U174, new_P3_R1110_U175, new_P3_R1110_U176,
    new_P3_R1110_U177, new_P3_R1110_U178, new_P3_R1110_U179,
    new_P3_R1110_U180, new_P3_R1110_U181, new_P3_R1110_U182,
    new_P3_R1110_U183, new_P3_R1110_U184, new_P3_R1110_U185,
    new_P3_R1110_U186, new_P3_R1110_U187, new_P3_R1110_U188,
    new_P3_R1110_U189, new_P3_R1110_U190, new_P3_R1110_U191,
    new_P3_R1110_U192, new_P3_R1110_U193, new_P3_R1110_U194,
    new_P3_R1110_U195, new_P3_R1110_U196, new_P3_R1110_U197,
    new_P3_R1110_U198, new_P3_R1110_U199, new_P3_R1110_U200,
    new_P3_R1110_U201, new_P3_R1110_U202, new_P3_R1110_U203,
    new_P3_R1110_U204, new_P3_R1110_U205, new_P3_R1110_U206,
    new_P3_R1110_U207, new_P3_R1110_U208, new_P3_R1110_U209,
    new_P3_R1110_U210, new_P3_R1110_U211, new_P3_R1110_U212,
    new_P3_R1110_U213, new_P3_R1110_U214, new_P3_R1110_U215,
    new_P3_R1110_U216, new_P3_R1110_U217, new_P3_R1110_U218,
    new_P3_R1110_U219, new_P3_R1110_U220, new_P3_R1110_U221,
    new_P3_R1110_U222, new_P3_R1110_U223, new_P3_R1110_U224,
    new_P3_R1110_U225, new_P3_R1110_U226, new_P3_R1110_U227,
    new_P3_R1110_U228, new_P3_R1110_U229, new_P3_R1110_U230,
    new_P3_R1110_U231, new_P3_R1110_U232, new_P3_R1110_U233,
    new_P3_R1110_U234, new_P3_R1110_U235, new_P3_R1110_U236,
    new_P3_R1110_U237, new_P3_R1110_U238, new_P3_R1110_U239,
    new_P3_R1110_U240, new_P3_R1110_U241, new_P3_R1110_U242,
    new_P3_R1110_U243, new_P3_R1110_U244, new_P3_R1110_U245,
    new_P3_R1110_U246, new_P3_R1110_U247, new_P3_R1110_U248,
    new_P3_R1110_U249, new_P3_R1110_U250, new_P3_R1110_U251,
    new_P3_R1110_U252, new_P3_R1110_U253, new_P3_R1110_U254,
    new_P3_R1110_U255, new_P3_R1110_U256, new_P3_R1110_U257,
    new_P3_R1110_U258, new_P3_R1110_U259, new_P3_R1110_U260,
    new_P3_R1110_U261, new_P3_R1110_U262, new_P3_R1110_U263,
    new_P3_R1110_U264, new_P3_R1110_U265, new_P3_R1110_U266,
    new_P3_R1110_U267, new_P3_R1110_U268, new_P3_R1110_U269,
    new_P3_R1110_U270, new_P3_R1110_U271, new_P3_R1110_U272,
    new_P3_R1110_U273, new_P3_R1110_U274, new_P3_R1110_U275,
    new_P3_R1110_U276, new_P3_R1110_U277, new_P3_R1110_U278,
    new_P3_R1110_U279, new_P3_R1110_U280, new_P3_R1110_U281,
    new_P3_R1110_U282, new_P3_R1110_U283, new_P3_R1110_U284,
    new_P3_R1110_U285, new_P3_R1110_U286, new_P3_R1110_U287,
    new_P3_R1110_U288, new_P3_R1110_U289, new_P3_R1110_U290,
    new_P3_R1110_U291, new_P3_R1110_U292, new_P3_R1110_U293,
    new_P3_R1110_U294, new_P3_R1110_U295, new_P3_R1110_U296,
    new_P3_R1110_U297, new_P3_R1110_U298, new_P3_R1110_U299,
    new_P3_R1110_U300, new_P3_R1110_U301, new_P3_R1110_U302,
    new_P3_R1110_U303, new_P3_R1110_U304, new_P3_R1110_U305,
    new_P3_R1110_U306, new_P3_R1110_U307, new_P3_R1110_U308,
    new_P3_R1110_U309, new_P3_R1110_U310, new_P3_R1110_U311,
    new_P3_R1110_U312, new_P3_R1110_U313, new_P3_R1110_U314,
    new_P3_R1110_U315, new_P3_R1110_U316, new_P3_R1110_U317,
    new_P3_R1110_U318, new_P3_R1110_U319, new_P3_R1110_U320,
    new_P3_R1110_U321, new_P3_R1110_U322, new_P3_R1110_U323,
    new_P3_R1110_U324, new_P3_R1110_U325, new_P3_R1110_U326,
    new_P3_R1110_U327, new_P3_R1110_U328, new_P3_R1110_U329,
    new_P3_R1110_U330, new_P3_R1110_U331, new_P3_R1110_U332,
    new_P3_R1110_U333, new_P3_R1110_U334, new_P3_R1110_U335,
    new_P3_R1110_U336, new_P3_R1110_U337, new_P3_R1110_U338,
    new_P3_R1110_U339, new_P3_R1110_U340, new_P3_R1110_U341,
    new_P3_R1110_U342, new_P3_R1110_U343, new_P3_R1110_U344,
    new_P3_R1110_U345, new_P3_R1110_U346, new_P3_R1110_U347,
    new_P3_R1110_U348, new_P3_R1110_U349, new_P3_R1110_U350,
    new_P3_R1110_U351, new_P3_R1110_U352, new_P3_R1110_U353,
    new_P3_R1110_U354, new_P3_R1110_U355, new_P3_R1110_U356,
    new_P3_R1110_U357, new_P3_R1110_U358, new_P3_R1110_U359,
    new_P3_R1110_U360, new_P3_R1110_U361, new_P3_R1110_U362,
    new_P3_R1110_U363, new_P3_R1110_U364, new_P3_R1110_U365,
    new_P3_R1110_U366, new_P3_R1110_U367, new_P3_R1110_U368,
    new_P3_R1110_U369, new_P3_R1110_U370, new_P3_R1110_U371,
    new_P3_R1110_U372, new_P3_R1110_U373, new_P3_R1110_U374,
    new_P3_R1110_U375, new_P3_R1110_U376, new_P3_R1110_U377,
    new_P3_R1110_U378, new_P3_R1110_U379, new_P3_R1110_U380,
    new_P3_R1110_U381, new_P3_R1110_U382, new_P3_R1110_U383,
    new_P3_R1110_U384, new_P3_R1110_U385, new_P3_R1110_U386,
    new_P3_R1110_U387, new_P3_R1110_U388, new_P3_R1110_U389,
    new_P3_R1110_U390, new_P3_R1110_U391, new_P3_R1110_U392,
    new_P3_R1110_U393, new_P3_R1110_U394, new_P3_R1110_U395,
    new_P3_R1110_U396, new_P3_R1110_U397, new_P3_R1110_U398,
    new_P3_R1110_U399, new_P3_R1110_U400, new_P3_R1110_U401,
    new_P3_R1110_U402, new_P3_R1110_U403, new_P3_R1110_U404,
    new_P3_R1110_U405, new_P3_R1110_U406, new_P3_R1110_U407,
    new_P3_R1110_U408, new_P3_R1110_U409, new_P3_R1110_U410,
    new_P3_R1110_U411, new_P3_R1110_U412, new_P3_R1110_U413,
    new_P3_R1110_U414, new_P3_R1110_U415, new_P3_R1110_U416,
    new_P3_R1110_U417, new_P3_R1110_U418, new_P3_R1110_U419,
    new_P3_R1110_U420, new_P3_R1110_U421, new_P3_R1110_U422,
    new_P3_R1110_U423, new_P3_R1110_U424, new_P3_R1110_U425,
    new_P3_R1110_U426, new_P3_R1110_U427, new_P3_R1110_U428,
    new_P3_R1110_U429, new_P3_R1110_U430, new_P3_R1110_U431,
    new_P3_R1110_U432, new_P3_R1110_U433, new_P3_R1110_U434,
    new_P3_R1110_U435, new_P3_R1110_U436, new_P3_R1110_U437,
    new_P3_R1110_U438, new_P3_R1110_U439, new_P3_R1110_U440,
    new_P3_R1110_U441, new_P3_R1110_U442, new_P3_R1110_U443,
    new_P3_R1110_U444, new_P3_R1110_U445, new_P3_R1110_U446,
    new_P3_R1110_U447, new_P3_R1110_U448, new_P3_R1110_U449,
    new_P3_R1110_U450, new_P3_R1110_U451, new_P3_R1110_U452,
    new_P3_R1110_U453, new_P3_R1110_U454, new_P3_R1110_U455,
    new_P3_R1110_U456, new_P3_R1110_U457, new_P3_R1110_U458,
    new_P3_R1110_U459, new_P3_R1110_U460, new_P3_R1110_U461,
    new_P3_R1110_U462, new_P3_R1110_U463, new_P3_R1110_U464,
    new_P3_R1110_U465, new_P3_R1110_U466, new_P3_R1110_U467,
    new_P3_R1110_U468, new_P3_R1110_U469, new_P3_R1110_U470,
    new_P3_R1110_U471, new_P3_R1110_U472, new_P3_R1110_U473,
    new_P3_R1110_U474, new_P3_R1110_U475, new_P3_R1110_U476,
    new_P3_R1110_U477, new_P3_R1110_U478, new_P3_R1110_U479,
    new_P3_R1110_U480, new_P3_R1110_U481, new_P3_R1110_U482,
    new_P3_R1110_U483, new_P3_R1110_U484, new_P3_R1110_U485,
    new_P3_R1110_U486, new_P3_R1110_U487, new_P3_R1110_U488,
    new_P3_R1110_U489, new_P3_R1110_U490, new_P3_R1110_U491,
    new_P3_R1110_U492, new_P3_R1110_U493, new_P3_R1110_U494,
    new_P3_R1110_U495, new_P3_R1110_U496, new_P3_R1110_U497,
    new_P3_R1110_U498, new_P3_R1110_U499, new_P3_R1110_U500,
    new_P3_R1110_U501, new_P3_R1110_U502, new_P3_R1110_U503,
    new_P3_R1110_U504, new_P3_R1297_U6, new_P3_R1297_U7, new_P3_R1077_U4,
    new_P3_R1077_U5, new_P3_R1077_U6, new_P3_R1077_U7, new_P3_R1077_U8,
    new_P3_R1077_U9, new_P3_R1077_U10, new_P3_R1077_U11, new_P3_R1077_U12,
    new_P3_R1077_U13, new_P3_R1077_U14, new_P3_R1077_U15, new_P3_R1077_U16,
    new_P3_R1077_U17, new_P3_R1077_U18, new_P3_R1077_U19, new_P3_R1077_U20,
    new_P3_R1077_U21, new_P3_R1077_U22, new_P3_R1077_U23, new_P3_R1077_U24,
    new_P3_R1077_U25, new_P3_R1077_U26, new_P3_R1077_U27, new_P3_R1077_U28,
    new_P3_R1077_U29, new_P3_R1077_U30, new_P3_R1077_U31, new_P3_R1077_U32,
    new_P3_R1077_U33, new_P3_R1077_U34, new_P3_R1077_U35, new_P3_R1077_U36,
    new_P3_R1077_U37, new_P3_R1077_U38, new_P3_R1077_U39, new_P3_R1077_U40,
    new_P3_R1077_U41, new_P3_R1077_U42, new_P3_R1077_U43, new_P3_R1077_U44,
    new_P3_R1077_U45, new_P3_R1077_U46, new_P3_R1077_U47, new_P3_R1077_U48,
    new_P3_R1077_U49, new_P3_R1077_U50, new_P3_R1077_U51, new_P3_R1077_U52,
    new_P3_R1077_U53, new_P3_R1077_U54, new_P3_R1077_U55, new_P3_R1077_U56,
    new_P3_R1077_U57, new_P3_R1077_U58, new_P3_R1077_U59, new_P3_R1077_U60,
    new_P3_R1077_U61, new_P3_R1077_U62, new_P3_R1077_U63, new_P3_R1077_U64,
    new_P3_R1077_U65, new_P3_R1077_U66, new_P3_R1077_U67, new_P3_R1077_U68,
    new_P3_R1077_U69, new_P3_R1077_U70, new_P3_R1077_U71, new_P3_R1077_U72,
    new_P3_R1077_U73, new_P3_R1077_U74, new_P3_R1077_U75, new_P3_R1077_U76,
    new_P3_R1077_U77, new_P3_R1077_U78, new_P3_R1077_U79, new_P3_R1077_U80,
    new_P3_R1077_U81, new_P3_R1077_U82, new_P3_R1077_U83, new_P3_R1077_U84,
    new_P3_R1077_U85, new_P3_R1077_U86, new_P3_R1077_U87, new_P3_R1077_U88,
    new_P3_R1077_U89, new_P3_R1077_U90, new_P3_R1077_U91, new_P3_R1077_U92,
    new_P3_R1077_U93, new_P3_R1077_U94, new_P3_R1077_U95, new_P3_R1077_U96,
    new_P3_R1077_U97, new_P3_R1077_U98, new_P3_R1077_U99,
    new_P3_R1077_U100, new_P3_R1077_U101, new_P3_R1077_U102,
    new_P3_R1077_U103, new_P3_R1077_U104, new_P3_R1077_U105,
    new_P3_R1077_U106, new_P3_R1077_U107, new_P3_R1077_U108,
    new_P3_R1077_U109, new_P3_R1077_U110, new_P3_R1077_U111,
    new_P3_R1077_U112, new_P3_R1077_U113, new_P3_R1077_U114,
    new_P3_R1077_U115, new_P3_R1077_U116, new_P3_R1077_U117,
    new_P3_R1077_U118, new_P3_R1077_U119, new_P3_R1077_U120,
    new_P3_R1077_U121, new_P3_R1077_U122, new_P3_R1077_U123,
    new_P3_R1077_U124, new_P3_R1077_U125, new_P3_R1077_U126,
    new_P3_R1077_U127, new_P3_R1077_U128, new_P3_R1077_U129,
    new_P3_R1077_U130, new_P3_R1077_U131, new_P3_R1077_U132,
    new_P3_R1077_U133, new_P3_R1077_U134, new_P3_R1077_U135,
    new_P3_R1077_U136, new_P3_R1077_U137, new_P3_R1077_U138,
    new_P3_R1077_U139, new_P3_R1077_U140, new_P3_R1077_U141,
    new_P3_R1077_U142, new_P3_R1077_U143, new_P3_R1077_U144,
    new_P3_R1077_U145, new_P3_R1077_U146, new_P3_R1077_U147,
    new_P3_R1077_U148, new_P3_R1077_U149, new_P3_R1077_U150,
    new_P3_R1077_U151, new_P3_R1077_U152, new_P3_R1077_U153,
    new_P3_R1077_U154, new_P3_R1077_U155, new_P3_R1077_U156,
    new_P3_R1077_U157, new_P3_R1077_U158, new_P3_R1077_U159,
    new_P3_R1077_U160, new_P3_R1077_U161, new_P3_R1077_U162,
    new_P3_R1077_U163, new_P3_R1077_U164, new_P3_R1077_U165,
    new_P3_R1077_U166, new_P3_R1077_U167, new_P3_R1077_U168,
    new_P3_R1077_U169, new_P3_R1077_U170, new_P3_R1077_U171,
    new_P3_R1077_U172, new_P3_R1077_U173, new_P3_R1077_U174,
    new_P3_R1077_U175, new_P3_R1077_U176, new_P3_R1077_U177,
    new_P3_R1077_U178, new_P3_R1077_U179, new_P3_R1077_U180,
    new_P3_R1077_U181, new_P3_R1077_U182, new_P3_R1077_U183,
    new_P3_R1077_U184, new_P3_R1077_U185, new_P3_R1077_U186,
    new_P3_R1077_U187, new_P3_R1077_U188, new_P3_R1077_U189,
    new_P3_R1077_U190, new_P3_R1077_U191, new_P3_R1077_U192,
    new_P3_R1077_U193, new_P3_R1077_U194, new_P3_R1077_U195,
    new_P3_R1077_U196, new_P3_R1077_U197, new_P3_R1077_U198,
    new_P3_R1077_U199, new_P3_R1077_U200, new_P3_R1077_U201,
    new_P3_R1077_U202, new_P3_R1077_U203, new_P3_R1077_U204,
    new_P3_R1077_U205, new_P3_R1077_U206, new_P3_R1077_U207,
    new_P3_R1077_U208, new_P3_R1077_U209, new_P3_R1077_U210,
    new_P3_R1077_U211, new_P3_R1077_U212, new_P3_R1077_U213,
    new_P3_R1077_U214, new_P3_R1077_U215, new_P3_R1077_U216,
    new_P3_R1077_U217, new_P3_R1077_U218, new_P3_R1077_U219,
    new_P3_R1077_U220, new_P3_R1077_U221, new_P3_R1077_U222,
    new_P3_R1077_U223, new_P3_R1077_U224, new_P3_R1077_U225,
    new_P3_R1077_U226, new_P3_R1077_U227, new_P3_R1077_U228,
    new_P3_R1077_U229, new_P3_R1077_U230, new_P3_R1077_U231,
    new_P3_R1077_U232, new_P3_R1077_U233, new_P3_R1077_U234,
    new_P3_R1077_U235, new_P3_R1077_U236, new_P3_R1077_U237,
    new_P3_R1077_U238, new_P3_R1077_U239, new_P3_R1077_U240,
    new_P3_R1077_U241, new_P3_R1077_U242, new_P3_R1077_U243,
    new_P3_R1077_U244, new_P3_R1077_U245, new_P3_R1077_U246,
    new_P3_R1077_U247, new_P3_R1077_U248, new_P3_R1077_U249,
    new_P3_R1077_U250, new_P3_R1077_U251, new_P3_R1077_U252,
    new_P3_R1077_U253, new_P3_R1077_U254, new_P3_R1077_U255,
    new_P3_R1077_U256, new_P3_R1077_U257, new_P3_R1077_U258,
    new_P3_R1077_U259, new_P3_R1077_U260, new_P3_R1077_U261,
    new_P3_R1077_U262, new_P3_R1077_U263, new_P3_R1077_U264,
    new_P3_R1077_U265, new_P3_R1077_U266, new_P3_R1077_U267,
    new_P3_R1077_U268, new_P3_R1077_U269, new_P3_R1077_U270,
    new_P3_R1077_U271, new_P3_R1077_U272, new_P3_R1077_U273,
    new_P3_R1077_U274, new_P3_R1077_U275, new_P3_R1077_U276,
    new_P3_R1077_U277, new_P3_R1077_U278, new_P3_R1077_U279,
    new_P3_R1077_U280, new_P3_R1077_U281, new_P3_R1077_U282,
    new_P3_R1077_U283, new_P3_R1077_U284, new_P3_R1077_U285,
    new_P3_R1077_U286, new_P3_R1077_U287, new_P3_R1077_U288,
    new_P3_R1077_U289, new_P3_R1077_U290, new_P3_R1077_U291,
    new_P3_R1077_U292, new_P3_R1077_U293, new_P3_R1077_U294,
    new_P3_R1077_U295, new_P3_R1077_U296, new_P3_R1077_U297,
    new_P3_R1077_U298, new_P3_R1077_U299, new_P3_R1077_U300,
    new_P3_R1077_U301, new_P3_R1077_U302, new_P3_R1077_U303,
    new_P3_R1077_U304, new_P3_R1077_U305, new_P3_R1077_U306,
    new_P3_R1077_U307, new_P3_R1077_U308, new_P3_R1077_U309,
    new_P3_R1077_U310, new_P3_R1077_U311, new_P3_R1077_U312,
    new_P3_R1077_U313, new_P3_R1077_U314, new_P3_R1077_U315,
    new_P3_R1077_U316, new_P3_R1077_U317, new_P3_R1077_U318,
    new_P3_R1077_U319, new_P3_R1077_U320, new_P3_R1077_U321,
    new_P3_R1077_U322, new_P3_R1077_U323, new_P3_R1077_U324,
    new_P3_R1077_U325, new_P3_R1077_U326, new_P3_R1077_U327,
    new_P3_R1077_U328, new_P3_R1077_U329, new_P3_R1077_U330,
    new_P3_R1077_U331, new_P3_R1077_U332, new_P3_R1077_U333,
    new_P3_R1077_U334, new_P3_R1077_U335, new_P3_R1077_U336,
    new_P3_R1077_U337, new_P3_R1077_U338, new_P3_R1077_U339,
    new_P3_R1077_U340, new_P3_R1077_U341, new_P3_R1077_U342,
    new_P3_R1077_U343, new_P3_R1077_U344, new_P3_R1077_U345,
    new_P3_R1077_U346, new_P3_R1077_U347, new_P3_R1077_U348,
    new_P3_R1077_U349, new_P3_R1077_U350, new_P3_R1077_U351,
    new_P3_R1077_U352, new_P3_R1077_U353, new_P3_R1077_U354,
    new_P3_R1077_U355, new_P3_R1077_U356, new_P3_R1077_U357,
    new_P3_R1077_U358, new_P3_R1077_U359, new_P3_R1077_U360,
    new_P3_R1077_U361, new_P3_R1077_U362, new_P3_R1077_U363,
    new_P3_R1077_U364, new_P3_R1077_U365, new_P3_R1077_U366,
    new_P3_R1077_U367, new_P3_R1077_U368, new_P3_R1077_U369,
    new_P3_R1077_U370, new_P3_R1077_U371, new_P3_R1077_U372,
    new_P3_R1077_U373, new_P3_R1077_U374, new_P3_R1077_U375,
    new_P3_R1077_U376, new_P3_R1077_U377, new_P3_R1077_U378,
    new_P3_R1077_U379, new_P3_R1077_U380, new_P3_R1077_U381,
    new_P3_R1077_U382, new_P3_R1077_U383, new_P3_R1077_U384,
    new_P3_R1077_U385, new_P3_R1077_U386, new_P3_R1077_U387,
    new_P3_R1077_U388, new_P3_R1077_U389, new_P3_R1077_U390,
    new_P3_R1077_U391, new_P3_R1077_U392, new_P3_R1077_U393,
    new_P3_R1077_U394, new_P3_R1077_U395, new_P3_R1077_U396,
    new_P3_R1077_U397, new_P3_R1077_U398, new_P3_R1077_U399,
    new_P3_R1077_U400, new_P3_R1077_U401, new_P3_R1077_U402,
    new_P3_R1077_U403, new_P3_R1077_U404, new_P3_R1077_U405,
    new_P3_R1077_U406, new_P3_R1077_U407, new_P3_R1077_U408,
    new_P3_R1077_U409, new_P3_R1077_U410, new_P3_R1077_U411,
    new_P3_R1077_U412, new_P3_R1077_U413, new_P3_R1077_U414,
    new_P3_R1077_U415, new_P3_R1077_U416, new_P3_R1077_U417,
    new_P3_R1077_U418, new_P3_R1077_U419, new_P3_R1077_U420,
    new_P3_R1077_U421, new_P3_R1077_U422, new_P3_R1077_U423,
    new_P3_R1077_U424, new_P3_R1077_U425, new_P3_R1077_U426,
    new_P3_R1077_U427, new_P3_R1077_U428, new_P3_R1077_U429,
    new_P3_R1077_U430, new_P3_R1077_U431, new_P3_R1077_U432,
    new_P3_R1077_U433, new_P3_R1077_U434, new_P3_R1077_U435,
    new_P3_R1077_U436, new_P3_R1077_U437, new_P3_R1077_U438,
    new_P3_R1077_U439, new_P3_R1077_U440, new_P3_R1077_U441,
    new_P3_R1077_U442, new_P3_R1077_U443, new_P3_R1077_U444,
    new_P3_R1077_U445, new_P3_R1077_U446, new_P3_R1077_U447,
    new_P3_R1077_U448, new_P3_R1077_U449, new_P3_R1077_U450,
    new_P3_R1077_U451, new_P3_R1077_U452, new_P3_R1077_U453,
    new_P3_R1077_U454, new_P3_R1077_U455, new_P3_R1077_U456,
    new_P3_R1077_U457, new_P3_R1077_U458, new_P3_R1077_U459,
    new_P3_R1077_U460, new_P3_R1077_U461, new_P3_R1077_U462,
    new_P3_R1077_U463, new_P3_R1077_U464, new_P3_R1077_U465,
    new_P3_R1077_U466, new_P3_R1077_U467, new_P3_R1077_U468,
    new_P3_R1077_U469, new_P3_R1077_U470, new_P3_R1077_U471,
    new_P3_R1077_U472, new_P3_R1077_U473, new_P3_R1077_U474,
    new_P3_R1077_U475, new_P3_R1077_U476, new_P3_R1077_U477,
    new_P3_R1077_U478, new_P3_R1077_U479, new_P3_R1077_U480,
    new_P3_R1077_U481, new_P3_R1077_U482, new_P3_R1077_U483,
    new_P3_R1077_U484, new_P3_R1077_U485, new_P3_R1077_U486,
    new_P3_R1077_U487, new_P3_R1077_U488, new_P3_R1077_U489,
    new_P3_R1077_U490, new_P3_R1077_U491, new_P3_R1077_U492,
    new_P3_R1077_U493, new_P3_R1077_U494, new_P3_R1077_U495,
    new_P3_R1077_U496, new_P3_R1077_U497, new_P3_R1077_U498,
    new_P3_R1077_U499, new_P3_R1077_U500, new_P3_R1077_U501,
    new_P3_R1077_U502, new_P3_R1077_U503, new_P3_R1077_U504,
    new_P3_R1143_U4, new_P3_R1143_U5, new_P3_R1143_U6, new_P3_R1143_U7,
    new_P3_R1143_U8, new_P3_R1143_U9, new_P3_R1143_U10, new_P3_R1143_U11,
    new_P3_R1143_U12, new_P3_R1143_U13, new_P3_R1143_U14, new_P3_R1143_U15,
    new_P3_R1143_U16, new_P3_R1143_U17, new_P3_R1143_U18, new_P3_R1143_U19,
    new_P3_R1143_U20, new_P3_R1143_U21, new_P3_R1143_U22, new_P3_R1143_U23,
    new_P3_R1143_U24, new_P3_R1143_U25, new_P3_R1143_U26, new_P3_R1143_U27,
    new_P3_R1143_U28, new_P3_R1143_U29, new_P3_R1143_U30, new_P3_R1143_U31,
    new_P3_R1143_U32, new_P3_R1143_U33, new_P3_R1143_U34, new_P3_R1143_U35,
    new_P3_R1143_U36, new_P3_R1143_U37, new_P3_R1143_U38, new_P3_R1143_U39,
    new_P3_R1143_U40, new_P3_R1143_U41, new_P3_R1143_U42, new_P3_R1143_U43,
    new_P3_R1143_U44, new_P3_R1143_U45, new_P3_R1143_U46, new_P3_R1143_U47,
    new_P3_R1143_U48, new_P3_R1143_U49, new_P3_R1143_U50, new_P3_R1143_U51,
    new_P3_R1143_U52, new_P3_R1143_U53, new_P3_R1143_U54, new_P3_R1143_U55,
    new_P3_R1143_U56, new_P3_R1143_U57, new_P3_R1143_U58, new_P3_R1143_U59,
    new_P3_R1143_U60, new_P3_R1143_U61, new_P3_R1143_U62, new_P3_R1143_U63,
    new_P3_R1143_U64, new_P3_R1143_U65, new_P3_R1143_U66, new_P3_R1143_U67,
    new_P3_R1143_U68, new_P3_R1143_U69, new_P3_R1143_U70, new_P3_R1143_U71,
    new_P3_R1143_U72, new_P3_R1143_U73, new_P3_R1143_U74, new_P3_R1143_U75,
    new_P3_R1143_U76, new_P3_R1143_U77, new_P3_R1143_U78, new_P3_R1143_U79,
    new_P3_R1143_U80, new_P3_R1143_U81, new_P3_R1143_U82, new_P3_R1143_U83,
    new_P3_R1143_U84, new_P3_R1143_U85, new_P3_R1143_U86, new_P3_R1143_U87,
    new_P3_R1143_U88, new_P3_R1143_U89, new_P3_R1143_U90, new_P3_R1143_U91,
    new_P3_R1143_U92, new_P3_R1143_U93, new_P3_R1143_U94, new_P3_R1143_U95,
    new_P3_R1143_U96, new_P3_R1143_U97, new_P3_R1143_U98, new_P3_R1143_U99,
    new_P3_R1143_U100, new_P3_R1143_U101, new_P3_R1143_U102,
    new_P3_R1143_U103, new_P3_R1143_U104, new_P3_R1143_U105,
    new_P3_R1143_U106, new_P3_R1143_U107, new_P3_R1143_U108,
    new_P3_R1143_U109, new_P3_R1143_U110, new_P3_R1143_U111,
    new_P3_R1143_U112, new_P3_R1143_U113, new_P3_R1143_U114,
    new_P3_R1143_U115, new_P3_R1143_U116, new_P3_R1143_U117,
    new_P3_R1143_U118, new_P3_R1143_U119, new_P3_R1143_U120,
    new_P3_R1143_U121, new_P3_R1143_U122, new_P3_R1143_U123,
    new_P3_R1143_U124, new_P3_R1143_U125, new_P3_R1143_U126,
    new_P3_R1143_U127, new_P3_R1143_U128, new_P3_R1143_U129,
    new_P3_R1143_U130, new_P3_R1143_U131, new_P3_R1143_U132,
    new_P3_R1143_U133, new_P3_R1143_U134, new_P3_R1143_U135,
    new_P3_R1143_U136, new_P3_R1143_U137, new_P3_R1143_U138,
    new_P3_R1143_U139, new_P3_R1143_U140, new_P3_R1143_U141,
    new_P3_R1143_U142, new_P3_R1143_U143, new_P3_R1143_U144,
    new_P3_R1143_U145, new_P3_R1143_U146, new_P3_R1143_U147,
    new_P3_R1143_U148, new_P3_R1143_U149, new_P3_R1143_U150,
    new_P3_R1143_U151, new_P3_R1143_U152, new_P3_R1143_U153,
    new_P3_R1143_U154, new_P3_R1143_U155, new_P3_R1143_U156,
    new_P3_R1143_U157, new_P3_R1143_U158, new_P3_R1143_U159,
    new_P3_R1143_U160, new_P3_R1143_U161, new_P3_R1143_U162,
    new_P3_R1143_U163, new_P3_R1143_U164, new_P3_R1143_U165,
    new_P3_R1143_U166, new_P3_R1143_U167, new_P3_R1143_U168,
    new_P3_R1143_U169, new_P3_R1143_U170, new_P3_R1143_U171,
    new_P3_R1143_U172, new_P3_R1143_U173, new_P3_R1143_U174,
    new_P3_R1143_U175, new_P3_R1143_U176, new_P3_R1143_U177,
    new_P3_R1143_U178, new_P3_R1143_U179, new_P3_R1143_U180,
    new_P3_R1143_U181, new_P3_R1143_U182, new_P3_R1143_U183,
    new_P3_R1143_U184, new_P3_R1143_U185, new_P3_R1143_U186,
    new_P3_R1143_U187, new_P3_R1143_U188, new_P3_R1143_U189,
    new_P3_R1143_U190, new_P3_R1143_U191, new_P3_R1143_U192,
    new_P3_R1143_U193, new_P3_R1143_U194, new_P3_R1143_U195,
    new_P3_R1143_U196, new_P3_R1143_U197, new_P3_R1143_U198,
    new_P3_R1143_U199, new_P3_R1143_U200, new_P3_R1143_U201,
    new_P3_R1143_U202, new_P3_R1143_U203, new_P3_R1143_U204,
    new_P3_R1143_U205, new_P3_R1143_U206, new_P3_R1143_U207,
    new_P3_R1143_U208, new_P3_R1143_U209, new_P3_R1143_U210,
    new_P3_R1143_U211, new_P3_R1143_U212, new_P3_R1143_U213,
    new_P3_R1143_U214, new_P3_R1143_U215, new_P3_R1143_U216,
    new_P3_R1143_U217, new_P3_R1143_U218, new_P3_R1143_U219,
    new_P3_R1143_U220, new_P3_R1143_U221, new_P3_R1143_U222,
    new_P3_R1143_U223, new_P3_R1143_U224, new_P3_R1143_U225,
    new_P3_R1143_U226, new_P3_R1143_U227, new_P3_R1143_U228,
    new_P3_R1143_U229, new_P3_R1143_U230, new_P3_R1143_U231,
    new_P3_R1143_U232, new_P3_R1143_U233, new_P3_R1143_U234,
    new_P3_R1143_U235, new_P3_R1143_U236, new_P3_R1143_U237,
    new_P3_R1143_U238, new_P3_R1143_U239, new_P3_R1143_U240,
    new_P3_R1143_U241, new_P3_R1143_U242, new_P3_R1143_U243,
    new_P3_R1143_U244, new_P3_R1143_U245, new_P3_R1143_U246,
    new_P3_R1143_U247, new_P3_R1143_U248, new_P3_R1143_U249,
    new_P3_R1143_U250, new_P3_R1143_U251, new_P3_R1143_U252,
    new_P3_R1143_U253, new_P3_R1143_U254, new_P3_R1143_U255,
    new_P3_R1143_U256, new_P3_R1143_U257, new_P3_R1143_U258,
    new_P3_R1143_U259, new_P3_R1143_U260, new_P3_R1143_U261,
    new_P3_R1143_U262, new_P3_R1143_U263, new_P3_R1143_U264,
    new_P3_R1143_U265, new_P3_R1143_U266, new_P3_R1143_U267,
    new_P3_R1143_U268, new_P3_R1143_U269, new_P3_R1143_U270,
    new_P3_R1143_U271, new_P3_R1143_U272, new_P3_R1143_U273,
    new_P3_R1143_U274, new_P3_R1143_U275, new_P3_R1143_U276,
    new_P3_R1143_U277, new_P3_R1143_U278, new_P3_R1143_U279,
    new_P3_R1143_U280, new_P3_R1143_U281, new_P3_R1143_U282,
    new_P3_R1143_U283, new_P3_R1143_U284, new_P3_R1143_U285,
    new_P3_R1143_U286, new_P3_R1143_U287, new_P3_R1143_U288,
    new_P3_R1143_U289, new_P3_R1143_U290, new_P3_R1143_U291,
    new_P3_R1143_U292, new_P3_R1143_U293, new_P3_R1143_U294,
    new_P3_R1143_U295, new_P3_R1143_U296, new_P3_R1143_U297,
    new_P3_R1143_U298, new_P3_R1143_U299, new_P3_R1143_U300,
    new_P3_R1143_U301, new_P3_R1143_U302, new_P3_R1143_U303,
    new_P3_R1143_U304, new_P3_R1143_U305, new_P3_R1143_U306,
    new_P3_R1143_U307, new_P3_R1143_U308, new_P3_R1143_U309,
    new_P3_R1143_U310, new_P3_R1143_U311, new_P3_R1143_U312,
    new_P3_R1143_U313, new_P3_R1143_U314, new_P3_R1143_U315,
    new_P3_R1143_U316, new_P3_R1143_U317, new_P3_R1143_U318,
    new_P3_R1143_U319, new_P3_R1143_U320, new_P3_R1143_U321,
    new_P3_R1143_U322, new_P3_R1143_U323, new_P3_R1143_U324,
    new_P3_R1143_U325, new_P3_R1143_U326, new_P3_R1143_U327,
    new_P3_R1143_U328, new_P3_R1143_U329, new_P3_R1143_U330,
    new_P3_R1143_U331, new_P3_R1143_U332, new_P3_R1143_U333,
    new_P3_R1143_U334, new_P3_R1143_U335, new_P3_R1143_U336,
    new_P3_R1143_U337, new_P3_R1143_U338, new_P3_R1143_U339,
    new_P3_R1143_U340, new_P3_R1143_U341, new_P3_R1143_U342,
    new_P3_R1143_U343, new_P3_R1143_U344, new_P3_R1143_U345,
    new_P3_R1143_U346, new_P3_R1143_U347, new_P3_R1143_U348,
    new_P3_R1143_U349, new_P3_R1143_U350, new_P3_R1143_U351,
    new_P3_R1143_U352, new_P3_R1143_U353, new_P3_R1143_U354,
    new_P3_R1143_U355, new_P3_R1143_U356, new_P3_R1143_U357,
    new_P3_R1143_U358, new_P3_R1143_U359, new_P3_R1143_U360,
    new_P3_R1143_U361, new_P3_R1143_U362, new_P3_R1143_U363,
    new_P3_R1143_U364, new_P3_R1143_U365, new_P3_R1143_U366,
    new_P3_R1143_U367, new_P3_R1143_U368, new_P3_R1143_U369,
    new_P3_R1143_U370, new_P3_R1143_U371, new_P3_R1143_U372,
    new_P3_R1143_U373, new_P3_R1143_U374, new_P3_R1143_U375,
    new_P3_R1143_U376, new_P3_R1143_U377, new_P3_R1143_U378,
    new_P3_R1143_U379, new_P3_R1143_U380, new_P3_R1143_U381,
    new_P3_R1143_U382, new_P3_R1143_U383, new_P3_R1143_U384,
    new_P3_R1143_U385, new_P3_R1143_U386, new_P3_R1143_U387,
    new_P3_R1143_U388, new_P3_R1143_U389, new_P3_R1143_U390,
    new_P3_R1143_U391, new_P3_R1143_U392, new_P3_R1143_U393,
    new_P3_R1143_U394, new_P3_R1143_U395, new_P3_R1143_U396,
    new_P3_R1143_U397, new_P3_R1143_U398, new_P3_R1143_U399,
    new_P3_R1143_U400, new_P3_R1143_U401, new_P3_R1143_U402,
    new_P3_R1143_U403, new_P3_R1143_U404, new_P3_R1143_U405,
    new_P3_R1143_U406, new_P3_R1143_U407, new_P3_R1143_U408,
    new_P3_R1143_U409, new_P3_R1143_U410, new_P3_R1143_U411,
    new_P3_R1143_U412, new_P3_R1143_U413, new_P3_R1143_U414,
    new_P3_R1143_U415, new_P3_R1143_U416, new_P3_R1143_U417,
    new_P3_R1143_U418, new_P3_R1143_U419, new_P3_R1143_U420,
    new_P3_R1143_U421, new_P3_R1143_U422, new_P3_R1143_U423,
    new_P3_R1143_U424, new_P3_R1143_U425, new_P3_R1143_U426,
    new_P3_R1143_U427, new_P3_R1143_U428, new_P3_R1143_U429,
    new_P3_R1143_U430, new_P3_R1143_U431, new_P3_R1143_U432,
    new_P3_R1143_U433, new_P3_R1143_U434, new_P3_R1143_U435,
    new_P3_R1143_U436, new_P3_R1143_U437, new_P3_R1143_U438,
    new_P3_R1143_U439, new_P3_R1143_U440, new_P3_R1143_U441,
    new_P3_R1143_U442, new_P3_R1143_U443, new_P3_R1143_U444,
    new_P3_R1143_U445, new_P3_R1143_U446, new_P3_R1143_U447,
    new_P3_R1143_U448, new_P3_R1143_U449, new_P3_R1143_U450,
    new_P3_R1143_U451, new_P3_R1143_U452, new_P3_R1143_U453,
    new_P3_R1143_U454, new_P3_R1143_U455, new_P3_R1143_U456,
    new_P3_R1143_U457, new_P3_R1143_U458, new_P3_R1143_U459,
    new_P3_R1143_U460, new_P3_R1143_U461, new_P3_R1143_U462,
    new_P3_R1143_U463, new_P3_R1143_U464, new_P3_R1143_U465,
    new_P3_R1143_U466, new_P3_R1143_U467, new_P3_R1143_U468,
    new_P3_R1143_U469, new_P3_R1143_U470, new_P3_R1143_U471,
    new_P3_R1143_U472, new_P3_R1143_U473, new_P3_R1143_U474,
    new_P3_R1143_U475, new_P3_R1143_U476, new_P3_R1143_U477,
    new_P3_R1143_U478, new_P3_R1143_U479, new_P3_R1143_U480,
    new_P3_R1143_U481, new_P3_R1143_U482, new_P3_R1143_U483,
    new_P3_R1143_U484, new_P3_R1143_U485, new_P3_R1143_U486,
    new_P3_R1143_U487, new_P3_R1143_U488, new_P3_R1143_U489,
    new_P3_R1143_U490, new_P3_R1143_U491, new_P3_R1143_U492,
    new_P3_R1143_U493, new_P3_R1143_U494, new_P3_R1143_U495,
    new_P3_R1143_U496, new_P3_R1143_U497, new_P3_R1143_U498,
    new_P3_R1143_U499, new_P3_R1143_U500, new_P3_R1143_U501,
    new_P3_R1143_U502, new_P3_R1143_U503, new_P3_R1143_U504,
    new_P3_R1158_U4, new_P3_R1158_U5, new_P3_R1158_U6, new_P3_R1158_U7,
    new_P3_R1158_U8, new_P3_R1158_U9, new_P3_R1158_U10, new_P3_R1158_U11,
    new_P3_R1158_U12, new_P3_R1158_U13, new_P3_R1158_U14, new_P3_R1158_U15,
    new_P3_R1158_U16, new_P3_R1158_U17, new_P3_R1158_U18, new_P3_R1158_U19,
    new_P3_R1158_U20, new_P3_R1158_U21, new_P3_R1158_U22, new_P3_R1158_U23,
    new_P3_R1158_U24, new_P3_R1158_U25, new_P3_R1158_U26, new_P3_R1158_U27,
    new_P3_R1158_U28, new_P3_R1158_U29, new_P3_R1158_U30, new_P3_R1158_U31,
    new_P3_R1158_U32, new_P3_R1158_U33, new_P3_R1158_U34, new_P3_R1158_U35,
    new_P3_R1158_U36, new_P3_R1158_U37, new_P3_R1158_U38, new_P3_R1158_U39,
    new_P3_R1158_U40, new_P3_R1158_U41, new_P3_R1158_U42, new_P3_R1158_U43,
    new_P3_R1158_U44, new_P3_R1158_U45, new_P3_R1158_U46, new_P3_R1158_U47,
    new_P3_R1158_U48, new_P3_R1158_U49, new_P3_R1158_U50, new_P3_R1158_U51,
    new_P3_R1158_U52, new_P3_R1158_U53, new_P3_R1158_U54, new_P3_R1158_U55,
    new_P3_R1158_U56, new_P3_R1158_U57, new_P3_R1158_U58, new_P3_R1158_U59,
    new_P3_R1158_U60, new_P3_R1158_U61, new_P3_R1158_U62, new_P3_R1158_U63,
    new_P3_R1158_U64, new_P3_R1158_U65, new_P3_R1158_U66, new_P3_R1158_U67,
    new_P3_R1158_U68, new_P3_R1158_U69, new_P3_R1158_U70, new_P3_R1158_U71,
    new_P3_R1158_U72, new_P3_R1158_U73, new_P3_R1158_U74, new_P3_R1158_U75,
    new_P3_R1158_U76, new_P3_R1158_U77, new_P3_R1158_U78, new_P3_R1158_U79,
    new_P3_R1158_U80, new_P3_R1158_U81, new_P3_R1158_U82, new_P3_R1158_U83,
    new_P3_R1158_U84, new_P3_R1158_U85, new_P3_R1158_U86, new_P3_R1158_U87,
    new_P3_R1158_U88, new_P3_R1158_U89, new_P3_R1158_U90, new_P3_R1158_U91,
    new_P3_R1158_U92, new_P3_R1158_U93, new_P3_R1158_U94, new_P3_R1158_U95,
    new_P3_R1158_U96, new_P3_R1158_U97, new_P3_R1158_U98, new_P3_R1158_U99,
    new_P3_R1158_U100, new_P3_R1158_U101, new_P3_R1158_U102,
    new_P3_R1158_U103, new_P3_R1158_U104, new_P3_R1158_U105,
    new_P3_R1158_U106, new_P3_R1158_U107, new_P3_R1158_U108,
    new_P3_R1158_U109, new_P3_R1158_U110, new_P3_R1158_U111,
    new_P3_R1158_U112, new_P3_R1158_U113, new_P3_R1158_U114,
    new_P3_R1158_U115, new_P3_R1158_U116, new_P3_R1158_U117,
    new_P3_R1158_U118, new_P3_R1158_U119, new_P3_R1158_U120,
    new_P3_R1158_U121, new_P3_R1158_U122, new_P3_R1158_U123,
    new_P3_R1158_U124, new_P3_R1158_U125, new_P3_R1158_U126,
    new_P3_R1158_U127, new_P3_R1158_U128, new_P3_R1158_U129,
    new_P3_R1158_U130, new_P3_R1158_U131, new_P3_R1158_U132,
    new_P3_R1158_U133, new_P3_R1158_U134, new_P3_R1158_U135,
    new_P3_R1158_U136, new_P3_R1158_U137, new_P3_R1158_U138,
    new_P3_R1158_U139, new_P3_R1158_U140, new_P3_R1158_U141,
    new_P3_R1158_U142, new_P3_R1158_U143, new_P3_R1158_U144,
    new_P3_R1158_U145, new_P3_R1158_U146, new_P3_R1158_U147,
    new_P3_R1158_U148, new_P3_R1158_U149, new_P3_R1158_U150,
    new_P3_R1158_U151, new_P3_R1158_U152, new_P3_R1158_U153,
    new_P3_R1158_U154, new_P3_R1158_U155, new_P3_R1158_U156,
    new_P3_R1158_U157, new_P3_R1158_U158, new_P3_R1158_U159,
    new_P3_R1158_U160, new_P3_R1158_U161, new_P3_R1158_U162,
    new_P3_R1158_U163, new_P3_R1158_U164, new_P3_R1158_U165,
    new_P3_R1158_U166, new_P3_R1158_U167, new_P3_R1158_U168,
    new_P3_R1158_U169, new_P3_R1158_U170, new_P3_R1158_U171,
    new_P3_R1158_U172, new_P3_R1158_U173, new_P3_R1158_U174,
    new_P3_R1158_U175, new_P3_R1158_U176, new_P3_R1158_U177,
    new_P3_R1158_U178, new_P3_R1158_U179, new_P3_R1158_U180,
    new_P3_R1158_U181, new_P3_R1158_U182, new_P3_R1158_U183,
    new_P3_R1158_U184, new_P3_R1158_U185, new_P3_R1158_U186,
    new_P3_R1158_U187, new_P3_R1158_U188, new_P3_R1158_U189,
    new_P3_R1158_U190, new_P3_R1158_U191, new_P3_R1158_U192,
    new_P3_R1158_U193, new_P3_R1158_U194, new_P3_R1158_U195,
    new_P3_R1158_U196, new_P3_R1158_U197, new_P3_R1158_U198,
    new_P3_R1158_U199, new_P3_R1158_U200, new_P3_R1158_U201,
    new_P3_R1158_U202, new_P3_R1158_U203, new_P3_R1158_U204,
    new_P3_R1158_U205, new_P3_R1158_U206, new_P3_R1158_U207,
    new_P3_R1158_U208, new_P3_R1158_U209, new_P3_R1158_U210,
    new_P3_R1158_U211, new_P3_R1158_U212, new_P3_R1158_U213,
    new_P3_R1158_U214, new_P3_R1158_U215, new_P3_R1158_U216,
    new_P3_R1158_U217, new_P3_R1158_U218, new_P3_R1158_U219,
    new_P3_R1158_U220, new_P3_R1158_U221, new_P3_R1158_U222,
    new_P3_R1158_U223, new_P3_R1158_U224, new_P3_R1158_U225,
    new_P3_R1158_U226, new_P3_R1158_U227, new_P3_R1158_U228,
    new_P3_R1158_U229, new_P3_R1158_U230, new_P3_R1158_U231,
    new_P3_R1158_U232, new_P3_R1158_U233, new_P3_R1158_U234,
    new_P3_R1158_U235, new_P3_R1158_U236, new_P3_R1158_U237,
    new_P3_R1158_U238, new_P3_R1158_U239, new_P3_R1158_U240,
    new_P3_R1158_U241, new_P3_R1158_U242, new_P3_R1158_U243,
    new_P3_R1158_U244, new_P3_R1158_U245, new_P3_R1158_U246,
    new_P3_R1158_U247, new_P3_R1158_U248, new_P3_R1158_U249,
    new_P3_R1158_U250, new_P3_R1158_U251, new_P3_R1158_U252,
    new_P3_R1158_U253, new_P3_R1158_U254, new_P3_R1158_U255,
    new_P3_R1158_U256, new_P3_R1158_U257, new_P3_R1158_U258,
    new_P3_R1158_U259, new_P3_R1158_U260, new_P3_R1158_U261,
    new_P3_R1158_U262, new_P3_R1158_U263, new_P3_R1158_U264,
    new_P3_R1158_U265, new_P3_R1158_U266, new_P3_R1158_U267,
    new_P3_R1158_U268, new_P3_R1158_U269, new_P3_R1158_U270,
    new_P3_R1158_U271, new_P3_R1158_U272, new_P3_R1158_U273,
    new_P3_R1158_U274, new_P3_R1158_U275, new_P3_R1158_U276,
    new_P3_R1158_U277, new_P3_R1158_U278, new_P3_R1158_U279,
    new_P3_R1158_U280, new_P3_R1158_U281, new_P3_R1158_U282,
    new_P3_R1158_U283, new_P3_R1158_U284, new_P3_R1158_U285,
    new_P3_R1158_U286, new_P3_R1158_U287, new_P3_R1158_U288,
    new_P3_R1158_U289, new_P3_R1158_U290, new_P3_R1158_U291,
    new_P3_R1158_U292, new_P3_R1158_U293, new_P3_R1158_U294,
    new_P3_R1158_U295, new_P3_R1158_U296, new_P3_R1158_U297,
    new_P3_R1158_U298, new_P3_R1158_U299, new_P3_R1158_U300,
    new_P3_R1158_U301, new_P3_R1158_U302, new_P3_R1158_U303,
    new_P3_R1158_U304, new_P3_R1158_U305, new_P3_R1158_U306,
    new_P3_R1158_U307, new_P3_R1158_U308, new_P3_R1158_U309,
    new_P3_R1158_U310, new_P3_R1158_U311, new_P3_R1158_U312,
    new_P3_R1158_U313, new_P3_R1158_U314, new_P3_R1158_U315,
    new_P3_R1158_U316, new_P3_R1158_U317, new_P3_R1158_U318,
    new_P3_R1158_U319, new_P3_R1158_U320, new_P3_R1158_U321,
    new_P3_R1158_U322, new_P3_R1158_U323, new_P3_R1158_U324,
    new_P3_R1158_U325, new_P3_R1158_U326, new_P3_R1158_U327,
    new_P3_R1158_U328, new_P3_R1158_U329, new_P3_R1158_U330,
    new_P3_R1158_U331, new_P3_R1158_U332, new_P3_R1158_U333,
    new_P3_R1158_U334, new_P3_R1158_U335, new_P3_R1158_U336,
    new_P3_R1158_U337, new_P3_R1158_U338, new_P3_R1158_U339,
    new_P3_R1158_U340, new_P3_R1158_U341, new_P3_R1158_U342,
    new_P3_R1158_U343, new_P3_R1158_U344, new_P3_R1158_U345,
    new_P3_R1158_U346, new_P3_R1158_U347, new_P3_R1158_U348,
    new_P3_R1158_U349, new_P3_R1158_U350, new_P3_R1158_U351,
    new_P3_R1158_U352, new_P3_R1158_U353, new_P3_R1158_U354,
    new_P3_R1158_U355, new_P3_R1158_U356, new_P3_R1158_U357,
    new_P3_R1158_U358, new_P3_R1158_U359, new_P3_R1158_U360,
    new_P3_R1158_U361, new_P3_R1158_U362, new_P3_R1158_U363,
    new_P3_R1158_U364, new_P3_R1158_U365, new_P3_R1158_U366,
    new_P3_R1158_U367, new_P3_R1158_U368, new_P3_R1158_U369,
    new_P3_R1158_U370, new_P3_R1158_U371, new_P3_R1158_U372,
    new_P3_R1158_U373, new_P3_R1158_U374, new_P3_R1158_U375,
    new_P3_R1158_U376, new_P3_R1158_U377, new_P3_R1158_U378,
    new_P3_R1158_U379, new_P3_R1158_U380, new_P3_R1158_U381,
    new_P3_R1158_U382, new_P3_R1158_U383, new_P3_R1158_U384,
    new_P3_R1158_U385, new_P3_R1158_U386, new_P3_R1158_U387,
    new_P3_R1158_U388, new_P3_R1158_U389, new_P3_R1158_U390,
    new_P3_R1158_U391, new_P3_R1158_U392, new_P3_R1158_U393,
    new_P3_R1158_U394, new_P3_R1158_U395, new_P3_R1158_U396,
    new_P3_R1158_U397, new_P3_R1158_U398, new_P3_R1158_U399,
    new_P3_R1158_U400, new_P3_R1158_U401, new_P3_R1158_U402,
    new_P3_R1158_U403, new_P3_R1158_U404, new_P3_R1158_U405,
    new_P3_R1158_U406, new_P3_R1158_U407, new_P3_R1158_U408,
    new_P3_R1158_U409, new_P3_R1158_U410, new_P3_R1158_U411,
    new_P3_R1158_U412, new_P3_R1158_U413, new_P3_R1158_U414,
    new_P3_R1158_U415, new_P3_R1158_U416, new_P3_R1158_U417,
    new_P3_R1158_U418, new_P3_R1158_U419, new_P3_R1158_U420,
    new_P3_R1158_U421, new_P3_R1158_U422, new_P3_R1158_U423,
    new_P3_R1158_U424, new_P3_R1158_U425, new_P3_R1158_U426,
    new_P3_R1158_U427, new_P3_R1158_U428, new_P3_R1158_U429,
    new_P3_R1158_U430, new_P3_R1158_U431, new_P3_R1158_U432,
    new_P3_R1158_U433, new_P3_R1158_U434, new_P3_R1158_U435,
    new_P3_R1158_U436, new_P3_R1158_U437, new_P3_R1158_U438,
    new_P3_R1158_U439, new_P3_R1158_U440, new_P3_R1158_U441,
    new_P3_R1158_U442, new_P3_R1158_U443, new_P3_R1158_U444,
    new_P3_R1158_U445, new_P3_R1158_U446, new_P3_R1158_U447,
    new_P3_R1158_U448, new_P3_R1158_U449, new_P3_R1158_U450,
    new_P3_R1158_U451, new_P3_R1158_U452, new_P3_R1158_U453,
    new_P3_R1158_U454, new_P3_R1158_U455, new_P3_R1158_U456,
    new_P3_R1158_U457, new_P3_R1158_U458, new_P3_R1158_U459,
    new_P3_R1158_U460, new_P3_R1158_U461, new_P3_R1158_U462,
    new_P3_R1158_U463, new_P3_R1158_U464, new_P3_R1158_U465,
    new_P3_R1158_U466, new_P3_R1158_U467, new_P3_R1158_U468,
    new_P3_R1158_U469, new_P3_R1158_U470, new_P3_R1158_U471,
    new_P3_R1158_U472, new_P3_R1158_U473, new_P3_R1158_U474,
    new_P3_R1158_U475, new_P3_R1158_U476, new_P3_R1158_U477,
    new_P3_R1158_U478, new_P3_R1158_U479, new_P3_R1158_U480,
    new_P3_R1158_U481, new_P3_R1158_U482, new_P3_R1158_U483,
    new_P3_R1158_U484, new_P3_R1158_U485, new_P3_R1158_U486,
    new_P3_R1158_U487, new_P3_R1158_U488, new_P3_R1158_U489,
    new_P3_R1158_U490, new_P3_R1158_U491, new_P3_R1158_U492,
    new_P3_R1158_U493, new_P3_R1158_U494, new_P3_R1158_U495,
    new_P3_R1158_U496, new_P3_R1158_U497, new_P3_R1158_U498,
    new_P3_R1158_U499, new_P3_R1158_U500, new_P3_R1158_U501,
    new_P3_R1158_U502, new_P3_R1158_U503, new_P3_R1158_U504,
    new_P3_R1158_U505, new_P3_R1158_U506, new_P3_R1158_U507,
    new_P3_R1158_U508, new_P3_R1158_U509, new_P3_R1158_U510,
    new_P3_R1158_U511, new_P3_R1158_U512, new_P3_R1158_U513,
    new_P3_R1158_U514, new_P3_R1158_U515, new_P3_R1158_U516,
    new_P3_R1158_U517, new_P3_R1158_U518, new_P3_R1158_U519,
    new_P3_R1158_U520, new_P3_R1158_U521, new_P3_R1158_U522,
    new_P3_R1158_U523, new_P3_R1158_U524, new_P3_R1158_U525,
    new_P3_R1158_U526, new_P3_R1158_U527, new_P3_R1158_U528,
    new_P3_R1158_U529, new_P3_R1158_U530, new_P3_R1158_U531,
    new_P3_R1158_U532, new_P3_R1158_U533, new_P3_R1158_U534,
    new_P3_R1158_U535, new_P3_R1158_U536, new_P3_R1158_U537,
    new_P3_R1158_U538, new_P3_R1158_U539, new_P3_R1158_U540,
    new_P3_R1158_U541, new_P3_R1158_U542, new_P3_R1158_U543,
    new_P3_R1158_U544, new_P3_R1158_U545, new_P3_R1158_U546,
    new_P3_R1158_U547, new_P3_R1158_U548, new_P3_R1158_U549,
    new_P3_R1158_U550, new_P3_R1158_U551, new_P3_R1158_U552,
    new_P3_R1158_U553, new_P3_R1158_U554, new_P3_R1158_U555,
    new_P3_R1158_U556, new_P3_R1158_U557, new_P3_R1158_U558,
    new_P3_R1158_U559, new_P3_R1158_U560, new_P3_R1158_U561,
    new_P3_R1158_U562, new_P3_R1158_U563, new_P3_R1158_U564,
    new_P3_R1158_U565, new_P3_R1158_U566, new_P3_R1158_U567,
    new_P3_R1158_U568, new_P3_R1158_U569, new_P3_R1158_U570,
    new_P3_R1158_U571, new_P3_R1158_U572, new_P3_R1158_U573,
    new_P3_R1158_U574, new_P3_R1158_U575, new_P3_R1158_U576,
    new_P3_R1158_U577, new_P3_R1158_U578, new_P3_R1158_U579,
    new_P3_R1158_U580, new_P3_R1158_U581, new_P3_R1158_U582,
    new_P3_R1158_U583, new_P3_R1158_U584, new_P3_R1158_U585,
    new_P3_R1158_U586, new_P3_R1158_U587, new_P3_R1158_U588,
    new_P3_R1158_U589, new_P3_R1158_U590, new_P3_R1158_U591,
    new_P3_R1158_U592, new_P3_R1158_U593, new_P3_R1158_U594,
    new_P3_R1158_U595, new_P3_R1158_U596, new_P3_R1158_U597,
    new_P3_R1158_U598, new_P3_R1158_U599, new_P3_R1158_U600,
    new_P3_R1158_U601, new_P3_R1158_U602, new_P3_R1158_U603,
    new_P3_R1158_U604, new_P3_R1158_U605, new_P3_R1158_U606,
    new_P3_R1158_U607, new_P3_R1158_U608, new_P3_R1158_U609,
    new_P3_R1158_U610, new_P3_R1158_U611, new_P3_R1158_U612,
    new_P3_R1158_U613, new_P3_R1158_U614, new_P3_R1158_U615,
    new_P3_R1158_U616, new_P3_R1158_U617, new_P3_R1158_U618,
    new_P3_R1158_U619, new_P3_R1158_U620, new_P3_R1158_U621,
    new_P3_R1158_U622, new_P3_R1158_U623, new_P3_R1158_U624,
    new_P3_R1158_U625, new_P3_R1158_U626, new_P3_R1158_U627,
    new_P3_R1158_U628, new_P3_R1158_U629, new_P3_R1158_U630,
    new_P3_R1158_U631, new_P3_R1158_U632, new_P3_R1131_U6, new_P3_R1131_U7,
    new_P3_R1131_U8, new_P3_R1131_U9, new_P3_R1131_U10, new_P3_R1131_U11,
    new_P3_R1131_U12, new_P3_R1131_U13, new_P3_R1131_U14, new_P3_R1131_U15,
    new_P3_R1131_U16, new_P3_R1131_U17, new_P3_R1131_U18, new_P3_R1131_U19,
    new_P3_R1131_U20, new_P3_R1131_U21, new_P3_R1131_U22, new_P3_R1131_U23,
    new_P3_R1131_U24, new_P3_R1131_U25, new_P3_R1131_U26, new_P3_R1131_U27,
    new_P3_R1131_U28, new_P3_R1131_U29, new_P3_R1131_U30, new_P3_R1131_U31,
    new_P3_R1131_U32, new_P3_R1131_U33, new_P3_R1131_U34, new_P3_R1131_U35,
    new_P3_R1131_U36, new_P3_R1131_U37, new_P3_R1131_U38, new_P3_R1131_U39,
    new_P3_R1131_U40, new_P3_R1131_U41, new_P3_R1131_U42, new_P3_R1131_U43,
    new_P3_R1131_U44, new_P3_R1131_U45, new_P3_R1131_U46, new_P3_R1131_U47,
    new_P3_R1131_U48, new_P3_R1131_U49, new_P3_R1131_U50, new_P3_R1131_U51,
    new_P3_R1131_U52, new_P3_R1131_U53, new_P3_R1131_U54, new_P3_R1131_U55,
    new_P3_R1131_U56, new_P3_R1131_U57, new_P3_R1131_U58, new_P3_R1131_U59,
    new_P3_R1131_U60, new_P3_R1131_U61, new_P3_R1131_U62, new_P3_R1131_U63,
    new_P3_R1131_U64, new_P3_R1131_U65, new_P3_R1131_U66, new_P3_R1131_U67,
    new_P3_R1131_U68, new_P3_R1131_U69, new_P3_R1131_U70, new_P3_R1131_U71,
    new_P3_R1131_U72, new_P3_R1131_U73, new_P3_R1131_U74, new_P3_R1131_U75,
    new_P3_R1131_U76, new_P3_R1131_U77, new_P3_R1131_U78, new_P3_R1131_U79,
    new_P3_R1131_U80, new_P3_R1131_U81, new_P3_R1131_U82, new_P3_R1131_U83,
    new_P3_R1131_U84, new_P3_R1131_U85, new_P3_R1131_U86, new_P3_R1131_U87,
    new_P3_R1131_U88, new_P3_R1131_U89, new_P3_R1131_U90, new_P3_R1131_U91,
    new_P3_R1131_U92, new_P3_R1131_U93, new_P3_R1131_U94, new_P3_R1131_U95,
    new_P3_R1131_U96, new_P3_R1131_U97, new_P3_R1131_U98, new_P3_R1131_U99,
    new_P3_R1131_U100, new_P3_R1131_U101, new_P3_R1131_U102,
    new_P3_R1131_U103, new_P3_R1131_U104, new_P3_R1131_U105,
    new_P3_R1131_U106, new_P3_R1131_U107, new_P3_R1131_U108,
    new_P3_R1131_U109, new_P3_R1131_U110, new_P3_R1131_U111,
    new_P3_R1131_U112, new_P3_R1131_U113, new_P3_R1131_U114,
    new_P3_R1131_U115, new_P3_R1131_U116, new_P3_R1131_U117,
    new_P3_R1131_U118, new_P3_R1131_U119, new_P3_R1131_U120,
    new_P3_R1131_U121, new_P3_R1131_U122, new_P3_R1131_U123,
    new_P3_R1131_U124, new_P3_R1131_U125, new_P3_R1131_U126,
    new_P3_R1131_U127, new_P3_R1131_U128, new_P3_R1131_U129,
    new_P3_R1131_U130, new_P3_R1131_U131, new_P3_R1131_U132,
    new_P3_R1131_U133, new_P3_R1131_U134, new_P3_R1131_U135,
    new_P3_R1131_U136, new_P3_R1131_U137, new_P3_R1131_U138,
    new_P3_R1131_U139, new_P3_R1131_U140, new_P3_R1131_U141,
    new_P3_R1131_U142, new_P3_R1131_U143, new_P3_R1131_U144,
    new_P3_R1131_U145, new_P3_R1131_U146, new_P3_R1131_U147,
    new_P3_R1131_U148, new_P3_R1131_U149, new_P3_R1131_U150,
    new_P3_R1131_U151, new_P3_R1131_U152, new_P3_R1131_U153,
    new_P3_R1131_U154, new_P3_R1131_U155, new_P3_R1131_U156,
    new_P3_R1131_U157, new_P3_R1131_U158, new_P3_R1131_U159,
    new_P3_R1131_U160, new_P3_R1131_U161, new_P3_R1131_U162,
    new_P3_R1131_U163, new_P3_R1131_U164, new_P3_R1131_U165,
    new_P3_R1131_U166, new_P3_R1131_U167, new_P3_R1131_U168,
    new_P3_R1131_U169, new_P3_R1131_U170, new_P3_R1131_U171,
    new_P3_R1131_U172, new_P3_R1131_U173, new_P3_R1131_U174,
    new_P3_R1131_U175, new_P3_R1131_U176, new_P3_R1131_U177,
    new_P3_R1131_U178, new_P3_R1131_U179, new_P3_R1131_U180,
    new_P3_R1131_U181, new_P3_R1131_U182, new_P3_R1131_U183,
    new_P3_R1131_U184, new_P3_R1131_U185, new_P3_R1131_U186,
    new_P3_R1131_U187, new_P3_R1131_U188, new_P3_R1131_U189,
    new_P3_R1131_U190, new_P3_R1131_U191, new_P3_R1131_U192,
    new_P3_R1131_U193, new_P3_R1131_U194, new_P3_R1131_U195,
    new_P3_R1131_U196, new_P3_R1131_U197, new_P3_R1131_U198,
    new_P3_R1131_U199, new_P3_R1131_U200, new_P3_R1131_U201,
    new_P3_R1131_U202, new_P3_R1131_U203, new_P3_R1131_U204,
    new_P3_R1131_U205, new_P3_R1131_U206, new_P3_R1131_U207,
    new_P3_R1131_U208, new_P3_R1131_U209, new_P3_R1131_U210,
    new_P3_R1131_U211, new_P3_R1131_U212, new_P3_R1131_U213,
    new_P3_R1131_U214, new_P3_R1131_U215, new_P3_R1131_U216,
    new_P3_R1131_U217, new_P3_R1131_U218, new_P3_R1131_U219,
    new_P3_R1131_U220, new_P3_R1131_U221, new_P3_R1131_U222,
    new_P3_R1131_U223, new_P3_R1131_U224, new_P3_R1131_U225,
    new_P3_R1131_U226, new_P3_R1131_U227, new_P3_R1131_U228,
    new_P3_R1131_U229, new_P3_R1131_U230, new_P3_R1131_U231,
    new_P3_R1131_U232, new_P3_R1131_U233, new_P3_R1131_U234,
    new_P3_R1131_U235, new_P3_R1131_U236, new_P3_R1131_U237,
    new_P3_R1131_U238, new_P3_R1131_U239, new_P3_R1131_U240,
    new_P3_R1131_U241, new_P3_R1131_U242, new_P3_R1131_U243,
    new_P3_R1131_U244, new_P3_R1131_U245, new_P3_R1131_U246,
    new_P3_R1131_U247, new_P3_R1131_U248, new_P3_R1131_U249,
    new_P3_R1131_U250, new_P3_R1131_U251, new_P3_R1131_U252,
    new_P3_R1131_U253, new_P3_R1131_U254, new_P3_R1131_U255,
    new_P3_R1131_U256, new_P3_R1131_U257, new_P3_R1131_U258,
    new_P3_R1131_U259, new_P3_R1131_U260, new_P3_R1131_U261,
    new_P3_R1131_U262, new_P3_R1131_U263, new_P3_R1131_U264,
    new_P3_R1131_U265, new_P3_R1131_U266, new_P3_R1131_U267,
    new_P3_R1131_U268, new_P3_R1131_U269, new_P3_R1131_U270,
    new_P3_R1131_U271, new_P3_R1131_U272, new_P3_R1131_U273,
    new_P3_R1131_U274, new_P3_R1131_U275, new_P3_R1131_U276,
    new_P3_R1131_U277, new_P3_R1131_U278, new_P3_R1131_U279,
    new_P3_R1131_U280, new_P3_R1131_U281, new_P3_R1131_U282,
    new_P3_R1131_U283, new_P3_R1131_U284, new_P3_R1131_U285,
    new_P3_R1131_U286, new_P3_R1131_U287, new_P3_R1131_U288,
    new_P3_R1131_U289, new_P3_R1131_U290, new_P3_R1131_U291,
    new_P3_R1131_U292, new_P3_R1131_U293, new_P3_R1131_U294,
    new_P3_R1131_U295, new_P3_R1131_U296, new_P3_R1131_U297,
    new_P3_R1131_U298, new_P3_R1131_U299, new_P3_R1131_U300,
    new_P3_R1131_U301, new_P3_R1131_U302, new_P3_R1131_U303,
    new_P3_R1131_U304, new_P3_R1131_U305, new_P3_R1131_U306,
    new_P3_R1131_U307, new_P3_R1131_U308, new_P3_R1131_U309,
    new_P3_R1131_U310, new_P3_R1131_U311, new_P3_R1131_U312,
    new_P3_R1131_U313, new_P3_R1131_U314, new_P3_R1131_U315,
    new_P3_R1131_U316, new_P3_R1131_U317, new_P3_R1131_U318,
    new_P3_R1131_U319, new_P3_R1131_U320, new_P3_R1131_U321,
    new_P3_R1131_U322, new_P3_R1131_U323, new_P3_R1131_U324,
    new_P3_R1131_U325, new_P3_R1131_U326, new_P3_R1131_U327,
    new_P3_R1131_U328, new_P3_R1131_U329, new_P3_R1131_U330,
    new_P3_R1131_U331, new_P3_R1131_U332, new_P3_R1131_U333,
    new_P3_R1131_U334, new_P3_R1131_U335, new_P3_R1131_U336,
    new_P3_R1131_U337, new_P3_R1131_U338, new_P3_R1131_U339,
    new_P3_R1131_U340, new_P3_R1131_U341, new_P3_R1131_U342,
    new_P3_R1131_U343, new_P3_R1131_U344, new_P3_R1131_U345,
    new_P3_R1131_U346, new_P3_R1131_U347, new_P3_R1131_U348,
    new_P3_R1131_U349, new_P3_R1131_U350, new_P3_R1131_U351,
    new_P3_R1131_U352, new_P3_R1131_U353, new_P3_R1131_U354,
    new_P3_R1131_U355, new_P3_R1131_U356, new_P3_R1131_U357,
    new_P3_R1131_U358, new_P3_R1131_U359, new_P3_R1131_U360,
    new_P3_R1131_U361, new_P3_R1131_U362, new_P3_R1131_U363,
    new_P3_R1131_U364, new_P3_R1131_U365, new_P3_R1131_U366,
    new_P3_R1131_U367, new_P3_R1131_U368, new_P3_R1131_U369,
    new_P3_R1131_U370, new_P3_R1131_U371, new_P3_R1131_U372,
    new_P3_R1131_U373, new_P3_R1131_U374, new_P3_R1131_U375,
    new_P3_R1131_U376, new_P3_R1131_U377, new_P3_R1131_U378,
    new_P3_R1131_U379, new_P3_R1131_U380, new_P3_R1131_U381,
    new_P3_R1131_U382, new_P3_R1131_U383, new_P3_R1131_U384,
    new_P3_R1131_U385, new_P3_R1131_U386, new_P3_R1131_U387,
    new_P3_R1131_U388, new_P3_R1131_U389, new_P3_R1131_U390,
    new_P3_R1131_U391, new_P3_R1131_U392, new_P3_R1131_U393,
    new_P3_R1131_U394, new_P3_R1131_U395, new_P3_R1131_U396,
    new_P3_R1131_U397, new_P3_R1131_U398, new_P3_R1131_U399,
    new_P3_R1131_U400, new_P3_R1131_U401, new_P3_R1131_U402,
    new_P3_R1131_U403, new_P3_R1131_U404, new_P3_R1131_U405,
    new_P3_R1131_U406, new_P3_R1131_U407, new_P3_R1131_U408,
    new_P3_R1131_U409, new_P3_R1131_U410, new_P3_R1131_U411,
    new_P3_R1131_U412, new_P3_R1131_U413, new_P3_R1131_U414,
    new_P3_R1131_U415, new_P3_R1131_U416, new_P3_R1131_U417,
    new_P3_R1131_U418, new_P3_R1131_U419, new_P3_R1131_U420,
    new_P3_R1131_U421, new_P3_R1131_U422, new_P3_R1131_U423,
    new_P3_R1131_U424, new_P3_R1131_U425, new_P3_R1131_U426,
    new_P3_R1131_U427, new_P3_R1131_U428, new_P3_R1131_U429,
    new_P3_R1131_U430, new_P3_R1131_U431, new_P3_R1131_U432,
    new_P3_R1131_U433, new_P3_R1131_U434, new_P3_R1131_U435,
    new_P3_R1131_U436, new_P3_R1131_U437, new_P3_R1131_U438,
    new_P3_R1131_U439, new_P3_R1131_U440, new_P3_R1131_U441,
    new_P3_R1131_U442, new_P3_R1131_U443, new_P3_R1131_U444,
    new_P3_R1131_U445, new_P3_R1131_U446, new_P3_R1131_U447,
    new_P3_R1131_U448, new_P3_R1131_U449, new_P3_R1131_U450,
    new_P3_R1131_U451, new_P3_R1131_U452, new_P3_R1131_U453,
    new_P3_R1131_U454, new_P3_R1131_U455, new_P3_R1131_U456,
    new_P3_R1131_U457, new_P3_R1131_U458, new_P3_R1131_U459,
    new_P3_R1131_U460, new_P3_R1131_U461, new_P3_R1131_U462,
    new_P3_R1131_U463, new_P3_R1131_U464, new_P3_R1131_U465,
    new_P3_R1131_U466, new_P3_R1131_U467, new_P3_R1131_U468,
    new_P3_R1131_U469, new_P3_R1131_U470, new_P3_R1131_U471,
    new_P3_R1131_U472, new_P3_R1131_U473, new_P3_R1131_U474,
    new_P3_R1131_U475, new_P3_R1131_U476, new_P3_R1131_U477,
    new_P3_R1131_U478, new_P3_R1131_U479, new_P3_R1131_U480,
    new_P3_R1131_U481, new_P3_R1131_U482, new_P3_R1131_U483,
    new_P3_R1131_U484, new_P3_R1131_U485, new_P3_R1054_U6, new_P3_R1054_U7,
    new_P3_R1054_U8, new_P3_R1054_U9, new_P3_R1054_U10, new_P3_R1054_U11,
    new_P3_R1054_U12, new_P3_R1054_U13, new_P3_R1054_U14, new_P3_R1054_U15,
    new_P3_R1054_U16, new_P3_R1054_U17, new_P3_R1054_U18, new_P3_R1054_U19,
    new_P3_R1054_U20, new_P3_R1054_U21, new_P3_R1054_U22, new_P3_R1054_U23,
    new_P3_R1054_U24, new_P3_R1054_U25, new_P3_R1054_U26, new_P3_R1054_U27,
    new_P3_R1054_U28, new_P3_R1054_U29, new_P3_R1054_U30, new_P3_R1054_U31,
    new_P3_R1054_U32, new_P3_R1054_U33, new_P3_R1054_U34, new_P3_R1054_U35,
    new_P3_R1054_U36, new_P3_R1054_U37, new_P3_R1054_U38, new_P3_R1054_U39,
    new_P3_R1054_U40, new_P3_R1054_U41, new_P3_R1054_U42, new_P3_R1054_U43,
    new_P3_R1054_U44, new_P3_R1054_U45, new_P3_R1054_U46, new_P3_R1054_U47,
    new_P3_R1054_U48, new_P3_R1054_U49, new_P3_R1054_U50, new_P3_R1054_U51,
    new_P3_R1054_U52, new_P3_R1054_U53, new_P3_R1054_U54, new_P3_R1054_U55,
    new_P3_R1054_U56, new_P3_R1054_U57, new_P3_R1054_U58, new_P3_R1054_U59,
    new_P3_R1054_U60, new_P3_R1054_U61, new_P3_R1054_U62, new_P3_R1054_U63,
    new_P3_R1054_U64, new_P3_R1054_U65, new_P3_R1054_U66, new_P3_R1054_U67,
    new_P3_R1054_U68, new_P3_R1054_U69, new_P3_R1054_U70, new_P3_R1054_U71,
    new_P3_R1054_U72, new_P3_R1054_U73, new_P3_R1054_U74, new_P3_R1054_U75,
    new_P3_R1054_U76, new_P3_R1054_U77, new_P3_R1054_U78, new_P3_R1054_U79,
    new_P3_R1054_U80, new_P3_R1054_U81, new_P3_R1054_U82, new_P3_R1054_U83,
    new_P3_R1054_U84, new_P3_R1054_U85, new_P3_R1054_U86, new_P3_R1054_U87,
    new_P3_R1054_U88, new_P3_R1054_U89, new_P3_R1054_U90, new_P3_R1054_U91,
    new_P3_R1054_U92, new_P3_R1054_U93, new_P3_R1054_U94, new_P3_R1054_U95,
    new_P3_R1054_U96, new_P3_R1054_U97, new_P3_R1054_U98, new_P3_R1054_U99,
    new_P3_R1054_U100, new_P3_R1054_U101, new_P3_R1054_U102,
    new_P3_R1054_U103, new_P3_R1054_U104, new_P3_R1054_U105,
    new_P3_R1054_U106, new_P3_R1054_U107, new_P3_R1054_U108,
    new_P3_R1054_U109, new_P3_R1054_U110, new_P3_R1054_U111,
    new_P3_R1054_U112, new_P3_R1054_U113, new_P3_R1054_U114,
    new_P3_R1054_U115, new_P3_R1054_U116, new_P3_R1054_U117,
    new_P3_R1054_U118, new_P3_R1054_U119, new_P3_R1054_U120,
    new_P3_R1054_U121, new_P3_R1054_U122, new_P3_R1054_U123,
    new_P3_R1054_U124, new_P3_R1054_U125, new_P3_R1054_U126,
    new_P3_R1054_U127, new_P3_R1054_U128, new_P3_R1054_U129,
    new_P3_R1054_U130, new_P3_R1054_U131, new_P3_R1054_U132,
    new_P3_R1054_U133, new_P3_R1054_U134, new_P3_R1054_U135,
    new_P3_R1054_U136, new_P3_R1054_U137, new_P3_R1054_U138,
    new_P3_R1054_U139, new_P3_R1054_U140, new_P3_R1054_U141,
    new_P3_R1054_U142, new_P3_R1054_U143, new_P3_R1054_U144,
    new_P3_R1054_U145, new_P3_R1054_U146, new_P3_R1054_U147,
    new_P3_R1054_U148, new_P3_R1054_U149, new_P3_R1054_U150,
    new_P3_R1054_U151, new_P3_R1054_U152, new_P3_R1054_U153,
    new_P3_R1054_U154, new_P3_R1054_U155, new_P3_R1054_U156,
    new_P3_R1054_U157, new_P3_R1054_U158, new_P3_R1054_U159,
    new_P3_R1054_U160, new_P3_R1054_U161, new_P3_R1054_U162,
    new_P3_R1054_U163, new_P3_R1054_U164, new_P3_R1054_U165,
    new_P3_R1054_U166, new_P3_R1054_U167, new_P3_R1054_U168,
    new_P3_R1054_U169, new_P3_R1054_U170, new_P3_R1054_U171,
    new_P3_R1054_U172, new_P3_R1054_U173, new_P3_R1054_U174,
    new_P3_R1054_U175, new_P3_R1054_U176, new_P3_R1054_U177,
    new_P3_R1054_U178, new_P3_R1054_U179, new_P3_R1054_U180,
    new_P3_R1054_U181, new_P3_R1054_U182, new_P3_R1054_U183,
    new_P3_R1054_U184, new_P3_R1054_U185, new_P3_R1054_U186,
    new_P3_R1054_U187, new_P3_R1054_U188, new_P3_R1054_U189,
    new_P3_R1054_U190, new_P3_R1054_U191, new_P3_R1054_U192,
    new_P3_R1054_U193, new_P3_R1054_U194, new_P3_R1054_U195,
    new_P3_R1054_U196, new_P3_R1054_U197, new_P3_R1054_U198,
    new_P3_R1054_U199, new_P3_R1054_U200, new_P3_R1054_U201,
    new_P3_R1054_U202, new_P3_R1054_U203, new_P3_R1054_U204,
    new_P3_R1054_U205, new_P3_R1054_U206, new_P3_R1054_U207,
    new_P3_R1054_U208, new_P3_R1054_U209, new_P3_R1054_U210,
    new_P3_R1054_U211, new_P3_R1054_U212, new_P3_R1054_U213,
    new_P3_R1054_U214, new_P3_R1054_U215, new_P3_R1054_U216,
    new_P3_R1054_U217, new_P3_R1054_U218, new_P3_R1054_U219,
    new_P3_R1054_U220, new_P3_R1054_U221, new_P3_R1054_U222,
    new_P3_R1054_U223, new_P3_R1054_U224, new_P3_R1054_U225,
    new_P3_R1054_U226, new_P3_R1054_U227, new_P3_R1054_U228,
    new_P3_R1054_U229, new_P3_R1054_U230, new_P3_R1054_U231,
    new_P3_R1054_U232, new_P3_R1054_U233, new_P3_R1054_U234,
    new_P3_R1054_U235, new_P3_R1054_U236, new_P3_R1054_U237,
    new_P3_R1054_U238, new_P3_R1054_U239, new_P3_R1054_U240,
    new_P3_R1054_U241, new_P3_R1054_U242, new_P3_R1054_U243,
    new_P3_R1054_U244, new_P3_R1054_U245, new_P3_R1054_U246,
    new_P3_R1054_U247, new_P3_R1054_U248, new_P3_R1054_U249,
    new_P3_R1054_U250, new_P3_R1054_U251, new_P3_R1054_U252,
    new_P3_R1054_U253, new_P3_R1054_U254, new_P3_R1054_U255,
    new_P3_R1054_U256, new_P3_R1054_U257, new_P3_R1054_U258,
    new_P3_R1054_U259, new_P3_R1054_U260, new_P3_R1054_U261,
    new_P3_R1054_U262, new_P3_R1054_U263, new_P3_R1054_U264,
    new_P3_R1054_U265, new_P3_R1054_U266, new_P3_R1054_U267,
    new_P3_R1054_U268, new_P3_R1054_U269, new_P3_R1054_U270,
    new_P3_R1054_U271, new_P3_R1054_U272, new_P3_R1054_U273,
    new_P3_R1054_U274, new_P3_R1054_U275, new_P3_R1054_U276,
    new_P3_R1054_U277, new_P3_R1054_U278, new_P3_R1054_U279,
    new_P3_R1054_U280, new_P3_R1054_U281, new_P3_R1054_U282,
    new_P3_R1054_U283, new_P3_R1054_U284, new_P3_R1054_U285,
    new_P3_R1054_U286, new_P3_R1054_U287, new_P3_R1054_U288,
    new_P3_R1054_U289, new_P3_R1054_U290, new_P3_R1054_U291,
    new_P3_R1054_U292, new_P3_R1054_U293, new_P3_R1054_U294,
    new_P3_R1161_U4, new_P3_R1161_U5, new_P3_R1161_U6, new_P3_R1161_U7,
    new_P3_R1161_U8, new_P3_R1161_U9, new_P3_R1161_U10, new_P3_R1161_U11,
    new_P3_R1161_U12, new_P3_R1161_U13, new_P3_R1161_U14, new_P3_R1161_U15,
    new_P3_R1161_U16, new_P3_R1161_U17, new_P3_R1161_U18, new_P3_R1161_U19,
    new_P3_R1161_U20, new_P3_R1161_U21, new_P3_R1161_U22, new_P3_R1161_U23,
    new_P3_R1161_U24, new_P3_R1161_U25, new_P3_R1161_U26, new_P3_R1161_U27,
    new_P3_R1161_U28, new_P3_R1161_U29, new_P3_R1161_U30, new_P3_R1161_U31,
    new_P3_R1161_U32, new_P3_R1161_U33, new_P3_R1161_U34, new_P3_R1161_U35,
    new_P3_R1161_U36, new_P3_R1161_U37, new_P3_R1161_U38, new_P3_R1161_U39,
    new_P3_R1161_U40, new_P3_R1161_U41, new_P3_R1161_U42, new_P3_R1161_U43,
    new_P3_R1161_U44, new_P3_R1161_U45, new_P3_R1161_U46, new_P3_R1161_U47,
    new_P3_R1161_U48, new_P3_R1161_U49, new_P3_R1161_U50, new_P3_R1161_U51,
    new_P3_R1161_U52, new_P3_R1161_U53, new_P3_R1161_U54, new_P3_R1161_U55,
    new_P3_R1161_U56, new_P3_R1161_U57, new_P3_R1161_U58, new_P3_R1161_U59,
    new_P3_R1161_U60, new_P3_R1161_U61, new_P3_R1161_U62, new_P3_R1161_U63,
    new_P3_R1161_U64, new_P3_R1161_U65, new_P3_R1161_U66, new_P3_R1161_U67,
    new_P3_R1161_U68, new_P3_R1161_U69, new_P3_R1161_U70, new_P3_R1161_U71,
    new_P3_R1161_U72, new_P3_R1161_U73, new_P3_R1161_U74, new_P3_R1161_U75,
    new_P3_R1161_U76, new_P3_R1161_U77, new_P3_R1161_U78, new_P3_R1161_U79,
    new_P3_R1161_U80, new_P3_R1161_U81, new_P3_R1161_U82, new_P3_R1161_U83,
    new_P3_R1161_U84, new_P3_R1161_U85, new_P3_R1161_U86, new_P3_R1161_U87,
    new_P3_R1161_U88, new_P3_R1161_U89, new_P3_R1161_U90, new_P3_R1161_U91,
    new_P3_R1161_U92, new_P3_R1161_U93, new_P3_R1161_U94, new_P3_R1161_U95,
    new_P3_R1161_U96, new_P3_R1161_U97, new_P3_R1161_U98, new_P3_R1161_U99,
    new_P3_R1161_U100, new_P3_R1161_U101, new_P3_R1161_U102,
    new_P3_R1161_U103, new_P3_R1161_U104, new_P3_R1161_U105,
    new_P3_R1161_U106, new_P3_R1161_U107, new_P3_R1161_U108,
    new_P3_R1161_U109, new_P3_R1161_U110, new_P3_R1161_U111,
    new_P3_R1161_U112, new_P3_R1161_U113, new_P3_R1161_U114,
    new_P3_R1161_U115, new_P3_R1161_U116, new_P3_R1161_U117,
    new_P3_R1161_U118, new_P3_R1161_U119, new_P3_R1161_U120,
    new_P3_R1161_U121, new_P3_R1161_U122, new_P3_R1161_U123,
    new_P3_R1161_U124, new_P3_R1161_U125, new_P3_R1161_U126,
    new_P3_R1161_U127, new_P3_R1161_U128, new_P3_R1161_U129,
    new_P3_R1161_U130, new_P3_R1161_U131, new_P3_R1161_U132,
    new_P3_R1161_U133, new_P3_R1161_U134, new_P3_R1161_U135,
    new_P3_R1161_U136, new_P3_R1161_U137, new_P3_R1161_U138,
    new_P3_R1161_U139, new_P3_R1161_U140, new_P3_R1161_U141,
    new_P3_R1161_U142, new_P3_R1161_U143, new_P3_R1161_U144,
    new_P3_R1161_U145, new_P3_R1161_U146, new_P3_R1161_U147,
    new_P3_R1161_U148, new_P3_R1161_U149, new_P3_R1161_U150,
    new_P3_R1161_U151, new_P3_R1161_U152, new_P3_R1161_U153,
    new_P3_R1161_U154, new_P3_R1161_U155, new_P3_R1161_U156,
    new_P3_R1161_U157, new_P3_R1161_U158, new_P3_R1161_U159,
    new_P3_R1161_U160, new_P3_R1161_U161, new_P3_R1161_U162,
    new_P3_R1161_U163, new_P3_R1161_U164, new_P3_R1161_U165,
    new_P3_R1161_U166, new_P3_R1161_U167, new_P3_R1161_U168,
    new_P3_R1161_U169, new_P3_R1161_U170, new_P3_R1161_U171,
    new_P3_R1161_U172, new_P3_R1161_U173, new_P3_R1161_U174,
    new_P3_R1161_U175, new_P3_R1161_U176, new_P3_R1161_U177,
    new_P3_R1161_U178, new_P3_R1161_U179, new_P3_R1161_U180,
    new_P3_R1161_U181, new_P3_R1161_U182, new_P3_R1161_U183,
    new_P3_R1161_U184, new_P3_R1161_U185, new_P3_R1161_U186,
    new_P3_R1161_U187, new_P3_R1161_U188, new_P3_R1161_U189,
    new_P3_R1161_U190, new_P3_R1161_U191, new_P3_R1161_U192,
    new_P3_R1161_U193, new_P3_R1161_U194, new_P3_R1161_U195,
    new_P3_R1161_U196, new_P3_R1161_U197, new_P3_R1161_U198,
    new_P3_R1161_U199, new_P3_R1161_U200, new_P3_R1161_U201,
    new_P3_R1161_U202, new_P3_R1161_U203, new_P3_R1161_U204,
    new_P3_R1161_U205, new_P3_R1161_U206, new_P3_R1161_U207,
    new_P3_R1161_U208, new_P3_R1161_U209, new_P3_R1161_U210,
    new_P3_R1161_U211, new_P3_R1161_U212, new_P3_R1161_U213,
    new_P3_R1161_U214, new_P3_R1161_U215, new_P3_R1161_U216,
    new_P3_R1161_U217, new_P3_R1161_U218, new_P3_R1161_U219,
    new_P3_R1161_U220, new_P3_R1161_U221, new_P3_R1161_U222,
    new_P3_R1161_U223, new_P3_R1161_U224, new_P3_R1161_U225,
    new_P3_R1161_U226, new_P3_R1161_U227, new_P3_R1161_U228,
    new_P3_R1161_U229, new_P3_R1161_U230, new_P3_R1161_U231,
    new_P3_R1161_U232, new_P3_R1161_U233, new_P3_R1161_U234,
    new_P3_R1161_U235, new_P3_R1161_U236, new_P3_R1161_U237,
    new_P3_R1161_U238, new_P3_R1161_U239, new_P3_R1161_U240,
    new_P3_R1161_U241, new_P3_R1161_U242, new_P3_R1161_U243,
    new_P3_R1161_U244, new_P3_R1161_U245, new_P3_R1161_U246,
    new_P3_R1161_U247, new_P3_R1161_U248, new_P3_R1161_U249,
    new_P3_R1161_U250, new_P3_R1161_U251, new_P3_R1161_U252,
    new_P3_R1161_U253, new_P3_R1161_U254, new_P3_R1161_U255,
    new_P3_R1161_U256, new_P3_R1161_U257, new_P3_R1161_U258,
    new_P3_R1161_U259, new_P3_R1161_U260, new_P3_R1161_U261,
    new_P3_R1161_U262, new_P3_R1161_U263, new_P3_R1161_U264,
    new_P3_R1161_U265, new_P3_R1161_U266, new_P3_R1161_U267,
    new_P3_R1161_U268, new_P3_R1161_U269, new_P3_R1161_U270,
    new_P3_R1161_U271, new_P3_R1161_U272, new_P3_R1161_U273,
    new_P3_R1161_U274, new_P3_R1161_U275, new_P3_R1161_U276,
    new_P3_R1161_U277, new_P3_R1161_U278, new_P3_R1161_U279,
    new_P3_R1161_U280, new_P3_R1161_U281, new_P3_R1161_U282,
    new_P3_R1161_U283, new_P3_R1161_U284, new_P3_R1161_U285,
    new_P3_R1161_U286, new_P3_R1161_U287, new_P3_R1161_U288,
    new_P3_R1161_U289, new_P3_R1161_U290, new_P3_R1161_U291,
    new_P3_R1161_U292, new_P3_R1161_U293, new_P3_R1161_U294,
    new_P3_R1161_U295, new_P3_R1161_U296, new_P3_R1161_U297,
    new_P3_R1161_U298, new_P3_R1161_U299, new_P3_R1161_U300,
    new_P3_R1161_U301, new_P3_R1161_U302, new_P3_R1161_U303,
    new_P3_R1161_U304, new_P3_R1161_U305, new_P3_R1161_U306,
    new_P3_R1161_U307, new_P3_R1161_U308, new_P3_R1161_U309,
    new_P3_R1161_U310, new_P3_R1161_U311, new_P3_R1161_U312,
    new_P3_R1161_U313, new_P3_R1161_U314, new_P3_R1161_U315,
    new_P3_R1161_U316, new_P3_R1161_U317, new_P3_R1161_U318,
    new_P3_R1161_U319, new_P3_R1161_U320, new_P3_R1161_U321,
    new_P3_R1161_U322, new_P3_R1161_U323, new_P3_R1161_U324,
    new_P3_R1161_U325, new_P3_R1161_U326, new_P3_R1161_U327,
    new_P3_R1161_U328, new_P3_R1161_U329, new_P3_R1161_U330,
    new_P3_R1161_U331, new_P3_R1161_U332, new_P3_R1161_U333,
    new_P3_R1161_U334, new_P3_R1161_U335, new_P3_R1161_U336,
    new_P3_R1161_U337, new_P3_R1161_U338, new_P3_R1161_U339,
    new_P3_R1161_U340, new_P3_R1161_U341, new_P3_R1161_U342,
    new_P3_R1161_U343, new_P3_R1161_U344, new_P3_R1161_U345,
    new_P3_R1161_U346, new_P3_R1161_U347, new_P3_R1161_U348,
    new_P3_R1161_U349, new_P3_R1161_U350, new_P3_R1161_U351,
    new_P3_R1161_U352, new_P3_R1161_U353, new_P3_R1161_U354,
    new_P3_R1161_U355, new_P3_R1161_U356, new_P3_R1161_U357,
    new_P3_R1161_U358, new_P3_R1161_U359, new_P3_R1161_U360,
    new_P3_R1161_U361, new_P3_R1161_U362, new_P3_R1161_U363,
    new_P3_R1161_U364, new_P3_R1161_U365, new_P3_R1161_U366,
    new_P3_R1161_U367, new_P3_R1161_U368, new_P3_R1161_U369,
    new_P3_R1161_U370, new_P3_R1161_U371, new_P3_R1161_U372,
    new_P3_R1161_U373, new_P3_R1161_U374, new_P3_R1161_U375,
    new_P3_R1161_U376, new_P3_R1161_U377, new_P3_R1161_U378,
    new_P3_R1161_U379, new_P3_R1161_U380, new_P3_R1161_U381,
    new_P3_R1161_U382, new_P3_R1161_U383, new_P3_R1161_U384,
    new_P3_R1161_U385, new_P3_R1161_U386, new_P3_R1161_U387,
    new_P3_R1161_U388, new_P3_R1161_U389, new_P3_R1161_U390,
    new_P3_R1161_U391, new_P3_R1161_U392, new_P3_R1161_U393,
    new_P3_R1161_U394, new_P3_R1161_U395, new_P3_R1161_U396,
    new_P3_R1161_U397, new_P3_R1161_U398, new_P3_R1161_U399,
    new_P3_R1161_U400, new_P3_R1161_U401, new_P3_R1161_U402,
    new_P3_R1161_U403, new_P3_R1161_U404, new_P3_R1161_U405,
    new_P3_R1161_U406, new_P3_R1161_U407, new_P3_R1161_U408,
    new_P3_R1161_U409, new_P3_R1161_U410, new_P3_R1161_U411,
    new_P3_R1161_U412, new_P3_R1161_U413, new_P3_R1161_U414,
    new_P3_R1161_U415, new_P3_R1161_U416, new_P3_R1161_U417,
    new_P3_R1161_U418, new_P3_R1161_U419, new_P3_R1161_U420,
    new_P3_R1161_U421, new_P3_R1161_U422, new_P3_R1161_U423,
    new_P3_R1161_U424, new_P3_R1161_U425, new_P3_R1161_U426,
    new_P3_R1161_U427, new_P3_R1161_U428, new_P3_R1161_U429,
    new_not_keyinput0, new_not_keyinput1, new_not_keyinput2,
    new_not_keyinput3, new_not_keyinput4, new_not_keyinput5,
    new_not_keyinput6, new_not_keyinput7, new_not_keyinput8,
    new_not_keyinput9, new_not_keyinput10, new_not_keyinput11,
    new_not_keyinput12, new_not_keyinput13, new_not_keyinput14,
    new_not_keyinput15, new_not_keyinput16, new_not_keyinput17,
    new_not_keyinput18, new_not_keyinput19, new_not_keyinput20,
    new_not_keyinput21, new_not_keyinput22, new_not_keyinput23,
    new_not_keyinput24, new_not_keyinput25, new_not_keyinput26,
    new_not_keyinput27, new_not_keyinput28, new_not_keyinput29,
    new_not_keyinput30, new_not_keyinput31, new_not_0, new_and_1,
    new_not_2, new_and_3, new_not_4, new_and_5, new_not_6, new_and_7,
    new_not_8, new_and_9, new_not_11, new_and_12, new_not_13, new_and_14,
    new_not_15, new_and_16, new_not_17, new_and_18, new_not_20, new_and_21,
    new_not_22, new_and_23, new_not_24, new_and_25, new_not_27, new_and_28,
    new_not_29, new_and_30, new_not_Q_0, new_not_Q_1, new_not_Q_2,
    new_not_Q_3, new_not_Q_4, new_count_state_1, new_count_state_2,
    new_count_state_3, new_count_state_4, new_count_state_5,
    new_count_state_6, new_count_state_7, new_count_state_8,
    new_count_state_9, new_count_state_10, new_count_state_11,
    new_count_state_12, new_count_state_13, new_count_state_14,
    new_count_state_15, new_count_state_16, new_count_state_17,
    new_count_state_18, new_count_state_19, new_count_state_20,
    new_count_state_21, new_count_state_22, new_count_state_23,
    new_count_state_24, new_count_state_25, new_count_state_26,
    new_count_state_27, new_count_state_28, new_count_state_29,
    new_count_state_30, new_count_state_31, new_y_mux_key0_and_0,
    new_y_mux_key0_and_1, new_y_mux_key0_and_2, new_y_mux_key0_and_3,
    new_y_mux_key0_and_4, new_y_mux_key0_and_5, new_y_mux_key0_and_6,
    new_y_mux_key0_and_7, new_y_mux_key0_and_8, new_y_mux_key0_and_9,
    new_y_mux_key0_and_10, new_y_mux_key0_and_11, new_y_mux_key0_and_12,
    new_y_mux_key0_and_13, new_y_mux_key0_and_14, new_y_mux_key0_and_15,
    new_y_mux_key0, new_y_mux_key1_and_0, new_y_mux_key1_and_1,
    new_y_mux_key1_and_2, new_y_mux_key1_and_3, new_y_mux_key1_and_4,
    new_y_mux_key1_and_5, new_y_mux_key1_and_6, new_y_mux_key1_and_7,
    new_y_mux_key1_and_8, new_y_mux_key1_and_9, new_y_mux_key1_and_10,
    new_y_mux_key1_and_11, new_y_mux_key1_and_12, new_y_mux_key1_and_13,
    new_y_mux_key1_and_14, new_y_mux_key1_and_15, new_y_mux_key1,
    new_y_mux_key2_and_0, new_y_mux_key2_and_1, new_y_mux_key2_and_2,
    new_y_mux_key2_and_3, new_y_mux_key2_and_4, new_y_mux_key2_and_5,
    new_y_mux_key2_and_6, new_y_mux_key2_and_7, new_y_mux_key2_and_8,
    new_y_mux_key2_and_9, new_y_mux_key2_and_10, new_y_mux_key2_and_11,
    new_y_mux_key2_and_12, new_y_mux_key2_and_13, new_y_mux_key2_and_14,
    new_y_mux_key2_and_15, new_y_mux_key2, new_y_mux_key3_and_0,
    new_y_mux_key3_and_1, new_y_mux_key3_and_2, new_y_mux_key3_and_3,
    new_y_mux_key3_and_4, new_y_mux_key3_and_5, new_y_mux_key3_and_6,
    new_y_mux_key3_and_7, new_y_mux_key3_and_8, new_y_mux_key3_and_9,
    new_y_mux_key3_and_10, new_y_mux_key3_and_11, new_y_mux_key3_and_12,
    new_y_mux_key3_and_13, new_y_mux_key3_and_14, new_y_mux_key3_and_15,
    new_y_mux_key3, new_y_mux_key4_and_0, new_y_mux_key4_and_1,
    new_y_mux_key4_and_2, new_y_mux_key4_and_3, new_y_mux_key4_and_4,
    new_y_mux_key4_and_5, new_y_mux_key4_and_6, new_y_mux_key4_and_7,
    new_y_mux_key4_and_8, new_y_mux_key4_and_9, new_y_mux_key4_and_10,
    new_y_mux_key4_and_11, new_y_mux_key4_and_12, new_y_mux_key4_and_13,
    new_y_mux_key4_and_14, new_y_mux_key4_and_15, new_y_mux_key4,
    new_y_mux_key5_and_0, new_y_mux_key5_and_1, new_y_mux_key5_and_2,
    new_y_mux_key5_and_3, new_y_mux_key5_and_4, new_y_mux_key5_and_5,
    new_y_mux_key5_and_6, new_y_mux_key5_and_7, new_y_mux_key5_and_8,
    new_y_mux_key5_and_9, new_y_mux_key5_and_10, new_y_mux_key5_and_11,
    new_y_mux_key5_and_12, new_y_mux_key5_and_13, new_y_mux_key5_and_14,
    new_y_mux_key5_and_15, new_y_mux_key5, new_y_mux_key6_and_0,
    new_y_mux_key6_and_1, new_y_mux_key6_and_2, new_y_mux_key6_and_3,
    new_y_mux_key6_and_4, new_y_mux_key6_and_5, new_y_mux_key6_and_6,
    new_y_mux_key6_and_7, new_y_mux_key6_and_8, new_y_mux_key6_and_9,
    new_y_mux_key6_and_10, new_y_mux_key6_and_11, new_y_mux_key6_and_12,
    new_y_mux_key6_and_13, new_y_mux_key6_and_14, new_y_mux_key6_and_15,
    new_y_mux_key6, new_y_mux_key7_and_0, new_y_mux_key7_and_1,
    new_y_mux_key7_and_2, new_y_mux_key7_and_3, new_y_mux_key7_and_4,
    new_y_mux_key7_and_5, new_y_mux_key7_and_6, new_y_mux_key7_and_7,
    new_y_mux_key7_and_8, new_y_mux_key7_and_9, new_y_mux_key7_and_10,
    new_y_mux_key7_and_11, new_y_mux_key7_and_12, new_y_mux_key7_and_13,
    new_y_mux_key7_and_14, new_y_mux_key7_and_15, new_y_mux_key7,
    new_y_mux_key8_and_0, new_y_mux_key8_and_1, new_y_mux_key8_and_2,
    new_y_mux_key8_and_3, new_y_mux_key8_and_4, new_y_mux_key8_and_5,
    new_y_mux_key8_and_6, new_y_mux_key8_and_7, new_y_mux_key8_and_8,
    new_y_mux_key8_and_9, new_y_mux_key8_and_10, new_y_mux_key8_and_11,
    new_y_mux_key8_and_12, new_y_mux_key8_and_13, new_y_mux_key8_and_14,
    new_y_mux_key8_and_15, new_y_mux_key8, new_y_mux_key9_and_0,
    new_y_mux_key9_and_1, new_y_mux_key9_and_2, new_y_mux_key9_and_3,
    new_y_mux_key9_and_4, new_y_mux_key9_and_5, new_y_mux_key9_and_6,
    new_y_mux_key9_and_7, new_y_mux_key9_and_8, new_y_mux_key9_and_9,
    new_y_mux_key9_and_10, new_y_mux_key9_and_11, new_y_mux_key9_and_12,
    new_y_mux_key9_and_13, new_y_mux_key9_and_14, new_y_mux_key9_and_15,
    new_y_mux_key9, new_y_mux_key10_and_0, new_y_mux_key10_and_1,
    new_y_mux_key10_and_2, new_y_mux_key10_and_3, new_y_mux_key10_and_4,
    new_y_mux_key10_and_5, new_y_mux_key10_and_6, new_y_mux_key10_and_7,
    new_y_mux_key10_and_8, new_y_mux_key10_and_9, new_y_mux_key10_and_10,
    new_y_mux_key10_and_11, new_y_mux_key10_and_12, new_y_mux_key10_and_13,
    new_y_mux_key10_and_14, new_y_mux_key10_and_15, new_y_mux_key10,
    new_y_mux_key11_and_0, new_y_mux_key11_and_1, new_y_mux_key11_and_2,
    new_y_mux_key11_and_3, new_y_mux_key11_and_4, new_y_mux_key11_and_5,
    new_y_mux_key11_and_6, new_y_mux_key11_and_7, new_y_mux_key11_and_8,
    new_y_mux_key11_and_9, new_y_mux_key11_and_10, new_y_mux_key11_and_11,
    new_y_mux_key11_and_12, new_y_mux_key11_and_13, new_y_mux_key11_and_14,
    new_y_mux_key11_and_15, new_y_mux_key11, new_y_mux_key12_and_0,
    new_y_mux_key12_and_1, new_y_mux_key12_and_2, new_y_mux_key12_and_3,
    new_y_mux_key12_and_4, new_y_mux_key12_and_5, new_y_mux_key12_and_6,
    new_y_mux_key12_and_7, new_y_mux_key12_and_8, new_y_mux_key12_and_9,
    new_y_mux_key12_and_10, new_y_mux_key12_and_11, new_y_mux_key12_and_12,
    new_y_mux_key12_and_13, new_y_mux_key12_and_14, new_y_mux_key12_and_15,
    new_y_mux_key12, new_y_mux_key13_and_0, new_y_mux_key13_and_1,
    new_y_mux_key13_and_2, new_y_mux_key13_and_3, new_y_mux_key13_and_4,
    new_y_mux_key13_and_5, new_y_mux_key13_and_6, new_y_mux_key13_and_7,
    new_y_mux_key13_and_8, new_y_mux_key13_and_9, new_y_mux_key13_and_10,
    new_y_mux_key13_and_11, new_y_mux_key13_and_12, new_y_mux_key13_and_13,
    new_y_mux_key13_and_14, new_y_mux_key13_and_15, new_y_mux_key13,
    new_y_mux_key14_and_0, new_y_mux_key14_and_1, new_y_mux_key14_and_2,
    new_y_mux_key14_and_3, new_y_mux_key14_and_4, new_y_mux_key14_and_5,
    new_y_mux_key14_and_6, new_y_mux_key14_and_7, new_y_mux_key14_and_8,
    new_y_mux_key14_and_9, new_y_mux_key14_and_10, new_y_mux_key14_and_11,
    new_y_mux_key14_and_12, new_y_mux_key14_and_13, new_y_mux_key14_and_14,
    new_y_mux_key14_and_15, new_y_mux_key14, new_y_mux_key15_and_0,
    new_y_mux_key15_and_1, new_y_mux_key15_and_2, new_y_mux_key15_and_3,
    new_y_mux_key15_and_4, new_y_mux_key15_and_5, new_y_mux_key15_and_6,
    new_y_mux_key15_and_7, new_y_mux_key15_and_8, new_y_mux_key15_and_9,
    new_y_mux_key15_and_10, new_y_mux_key15_and_11, new_y_mux_key15_and_12,
    new_y_mux_key15_and_13, new_y_mux_key15_and_14, new_y_mux_key15_and_15,
    new_y_mux_key15, new_y_mux_key16_and_0, new_y_mux_key16_and_1,
    new_y_mux_key16_and_2, new_y_mux_key16_and_3, new_y_mux_key16_and_4,
    new_y_mux_key16_and_5, new_y_mux_key16_and_6, new_y_mux_key16_and_7,
    new_y_mux_key16_and_8, new_y_mux_key16_and_9, new_y_mux_key16_and_10,
    new_y_mux_key16_and_11, new_y_mux_key16_and_12, new_y_mux_key16_and_13,
    new_y_mux_key16_and_14, new_y_mux_key16_and_15, new_y_mux_key16,
    new_y_mux_key17_and_0, new_y_mux_key17_and_1, new_y_mux_key17_and_2,
    new_y_mux_key17_and_3, new_y_mux_key17_and_4, new_y_mux_key17_and_5,
    new_y_mux_key17_and_6, new_y_mux_key17_and_7, new_y_mux_key17_and_8,
    new_y_mux_key17_and_9, new_y_mux_key17_and_10, new_y_mux_key17_and_11,
    new_y_mux_key17_and_12, new_y_mux_key17_and_13, new_y_mux_key17_and_14,
    new_y_mux_key17_and_15, new_y_mux_key17, new_y_mux_key18_and_0,
    new_y_mux_key18_and_1, new_y_mux_key18_and_2, new_y_mux_key18_and_3,
    new_y_mux_key18_and_4, new_y_mux_key18_and_5, new_y_mux_key18_and_6,
    new_y_mux_key18_and_7, new_y_mux_key18_and_8, new_y_mux_key18_and_9,
    new_y_mux_key18_and_10, new_y_mux_key18_and_11, new_y_mux_key18_and_12,
    new_y_mux_key18_and_13, new_y_mux_key18_and_14, new_y_mux_key18_and_15,
    new_y_mux_key18, new_y_mux_key19_and_0, new_y_mux_key19_and_1,
    new_y_mux_key19_and_2, new_y_mux_key19_and_3, new_y_mux_key19_and_4,
    new_y_mux_key19_and_5, new_y_mux_key19_and_6, new_y_mux_key19_and_7,
    new_y_mux_key19_and_8, new_y_mux_key19_and_9, new_y_mux_key19_and_10,
    new_y_mux_key19_and_11, new_y_mux_key19_and_12, new_y_mux_key19_and_13,
    new_y_mux_key19_and_14, new_y_mux_key19_and_15, new_y_mux_key19,
    new_y_mux_key20_and_0, new_y_mux_key20_and_1, new_y_mux_key20_and_2,
    new_y_mux_key20_and_3, new_y_mux_key20_and_4, new_y_mux_key20_and_5,
    new_y_mux_key20_and_6, new_y_mux_key20_and_7, new_y_mux_key20_and_8,
    new_y_mux_key20_and_9, new_y_mux_key20_and_10, new_y_mux_key20_and_11,
    new_y_mux_key20_and_12, new_y_mux_key20_and_13, new_y_mux_key20_and_14,
    new_y_mux_key20_and_15, new_y_mux_key20, new_y_mux_key21_and_0,
    new_y_mux_key21_and_1, new_y_mux_key21_and_2, new_y_mux_key21_and_3,
    new_y_mux_key21_and_4, new_y_mux_key21_and_5, new_y_mux_key21_and_6,
    new_y_mux_key21_and_7, new_y_mux_key21_and_8, new_y_mux_key21_and_9,
    new_y_mux_key21_and_10, new_y_mux_key21_and_11, new_y_mux_key21_and_12,
    new_y_mux_key21_and_13, new_y_mux_key21_and_14, new_y_mux_key21_and_15,
    new_y_mux_key21, new_y_mux_key22_and_0, new_y_mux_key22_and_1,
    new_y_mux_key22_and_2, new_y_mux_key22_and_3, new_y_mux_key22_and_4,
    new_y_mux_key22_and_5, new_y_mux_key22_and_6, new_y_mux_key22_and_7,
    new_y_mux_key22_and_8, new_y_mux_key22_and_9, new_y_mux_key22_and_10,
    new_y_mux_key22_and_11, new_y_mux_key22_and_12, new_y_mux_key22_and_13,
    new_y_mux_key22_and_14, new_y_mux_key22_and_15, new_y_mux_key22,
    new_y_mux_key23_and_0, new_y_mux_key23_and_1, new_y_mux_key23_and_2,
    new_y_mux_key23_and_3, new_y_mux_key23_and_4, new_y_mux_key23_and_5,
    new_y_mux_key23_and_6, new_y_mux_key23_and_7, new_y_mux_key23_and_8,
    new_y_mux_key23_and_9, new_y_mux_key23_and_10, new_y_mux_key23_and_11,
    new_y_mux_key23_and_12, new_y_mux_key23_and_13, new_y_mux_key23_and_14,
    new_y_mux_key23_and_15, new_y_mux_key23, new_y_mux_key24_and_0,
    new_y_mux_key24_and_1, new_y_mux_key24_and_2, new_y_mux_key24_and_3,
    new_y_mux_key24_and_4, new_y_mux_key24_and_5, new_y_mux_key24_and_6,
    new_y_mux_key24_and_7, new_y_mux_key24_and_8, new_y_mux_key24_and_9,
    new_y_mux_key24_and_10, new_y_mux_key24_and_11, new_y_mux_key24_and_12,
    new_y_mux_key24_and_13, new_y_mux_key24_and_14, new_y_mux_key24_and_15,
    new_y_mux_key24, new_y_mux_key25_and_0, new_y_mux_key25_and_1,
    new_y_mux_key25_and_2, new_y_mux_key25_and_3, new_y_mux_key25_and_4,
    new_y_mux_key25_and_5, new_y_mux_key25_and_6, new_y_mux_key25_and_7,
    new_y_mux_key25_and_8, new_y_mux_key25_and_9, new_y_mux_key25_and_10,
    new_y_mux_key25_and_11, new_y_mux_key25_and_12, new_y_mux_key25_and_13,
    new_y_mux_key25_and_14, new_y_mux_key25_and_15, new_y_mux_key25,
    new_y_mux_key26_and_0, new_y_mux_key26_and_1, new_y_mux_key26_and_2,
    new_y_mux_key26_and_3, new_y_mux_key26_and_4, new_y_mux_key26_and_5,
    new_y_mux_key26_and_6, new_y_mux_key26_and_7, new_y_mux_key26_and_8,
    new_y_mux_key26_and_9, new_y_mux_key26_and_10, new_y_mux_key26_and_11,
    new_y_mux_key26_and_12, new_y_mux_key26_and_13, new_y_mux_key26_and_14,
    new_y_mux_key26_and_15, new_y_mux_key26, new_y_mux_key27_and_0,
    new_y_mux_key27_and_1, new_y_mux_key27_and_2, new_y_mux_key27_and_3,
    new_y_mux_key27_and_4, new_y_mux_key27_and_5, new_y_mux_key27_and_6,
    new_y_mux_key27_and_7, new_y_mux_key27_and_8, new_y_mux_key27_and_9,
    new_y_mux_key27_and_10, new_y_mux_key27_and_11, new_y_mux_key27_and_12,
    new_y_mux_key27_and_13, new_y_mux_key27_and_14, new_y_mux_key27_and_15,
    new_y_mux_key27, new_y_mux_key28_and_0, new_y_mux_key28_and_1,
    new_y_mux_key28_and_2, new_y_mux_key28_and_3, new_y_mux_key28_and_4,
    new_y_mux_key28_and_5, new_y_mux_key28_and_6, new_y_mux_key28_and_7,
    new_y_mux_key28_and_8, new_y_mux_key28_and_9, new_y_mux_key28_and_10,
    new_y_mux_key28_and_11, new_y_mux_key28_and_12, new_y_mux_key28_and_13,
    new_y_mux_key28_and_14, new_y_mux_key28_and_15, new_y_mux_key28,
    new_y_mux_key29_and_0, new_y_mux_key29_and_1, new_y_mux_key29_and_2,
    new_y_mux_key29_and_3, new_y_mux_key29_and_4, new_y_mux_key29_and_5,
    new_y_mux_key29_and_6, new_y_mux_key29_and_7, new_y_mux_key29_and_8,
    new_y_mux_key29_and_9, new_y_mux_key29_and_10, new_y_mux_key29_and_11,
    new_y_mux_key29_and_12, new_y_mux_key29_and_13, new_y_mux_key29_and_14,
    new_y_mux_key29_and_15, new_y_mux_key29, new_y_mux_key30_and_0,
    new_y_mux_key30_and_1, new_y_mux_key30_and_2, new_y_mux_key30_and_3,
    new_y_mux_key30_and_4, new_y_mux_key30_and_5, new_y_mux_key30_and_6,
    new_y_mux_key30_and_7, new_y_mux_key30_and_8, new_y_mux_key30_and_9,
    new_y_mux_key30_and_10, new_y_mux_key30_and_11, new_y_mux_key30_and_12,
    new_y_mux_key30_and_13, new_y_mux_key30_and_14, new_y_mux_key30_and_15,
    new_y_mux_key30, new_y_mux_key31_and_0, new_y_mux_key31_and_1,
    new_y_mux_key31_and_2, new_y_mux_key31_and_3, new_y_mux_key31_and_4,
    new_y_mux_key31_and_5, new_y_mux_key31_and_6, new_y_mux_key31_and_7,
    new_y_mux_key31_and_8, new_y_mux_key31_and_9, new_y_mux_key31_and_10,
    new_y_mux_key31_and_11, new_y_mux_key31_and_12, new_y_mux_key31_and_13,
    new_y_mux_key31_and_14, new_y_mux_key31_and_15, new_y_mux_key31,
    new__state_1, new__state_2, new__state_3, new__state_4, new__state_5,
    new__state_6, new__state_7, new__state_8, new__state_9, new__state_10,
    new__state_11, new__state_12, new__state_13, new__state_14,
    new__state_15, new__state_16, new__state_17, new__state_18,
    new__state_19, new__state_20, new__state_21, new__state_22,
    new__state_23, new__state_24, new__state_25, new__state_26,
    new__state_27, new__state_28, new__state_29, new__state_30,
    new__state_31, new__state_33, new__state_34, new__state_35,
    new__state_36, new__state_37, new__state_38, new__state_39,
    new__state_40, new__state_41, new__state_42, new__state_43,
    new__state_44, new__state_45, new__state_46, new__state_47,
    new__state_49, new__state_50, new__state_51, new__state_52,
    new__state_53, new__state_54, new__state_55, new__state_57,
    new__state_58, new__state_59, new__state_61, new_s__state_1,
    new_not_s__state_1, new_I0__state_1, new_I1__state_1,
    new_and_mux__state_1, new_and_mux__state_1_2, new_y_mux_32,
    new_s__state_3, new_not_s__state_3, new_I0__state_3, new_I1__state_3,
    new_and_mux__state_3, new_and_mux__state_3_2, new_y_mux_33,
    new_s__state_5, new_not_s__state_5, new_I0__state_5, new_I1__state_5,
    new_and_mux__state_5, new_and_mux__state_5_2, new_y_mux_34,
    new_s__state_7, new_not_s__state_7, new_I0__state_7, new_I1__state_7,
    new_and_mux__state_7, new_and_mux__state_7_2, new_y_mux_35,
    new_s__state_9, new_not_s__state_9, new_I0__state_9, new_I1__state_9,
    new_and_mux__state_9, new_and_mux__state_9_2, new_y_mux_36,
    new_s__state_11, new_not_s__state_11, new_I0__state_11,
    new_I1__state_11, new_and_mux__state_11, new_and_mux__state_11_2,
    new_y_mux_37, new_s__state_13, new_not_s__state_13, new_I0__state_13,
    new_I1__state_13, new_and_mux__state_13, new_and_mux__state_13_2,
    new_y_mux_38, new_s__state_15, new_not_s__state_15, new_I0__state_15,
    new_I1__state_15, new_and_mux__state_15, new_and_mux__state_15_2,
    new_y_mux_39, new_s__state_17, new_not_s__state_17, new_I0__state_17,
    new_I1__state_17, new_and_mux__state_17, new_and_mux__state_17_2,
    new_y_mux_40, new_s__state_19, new_not_s__state_19, new_I0__state_19,
    new_I1__state_19, new_and_mux__state_19, new_and_mux__state_19_2,
    new_y_mux_41, new_s__state_21, new_not_s__state_21, new_I0__state_21,
    new_I1__state_21, new_and_mux__state_21, new_and_mux__state_21_2,
    new_y_mux_42, new_s__state_23, new_not_s__state_23, new_I0__state_23,
    new_I1__state_23, new_and_mux__state_23, new_and_mux__state_23_2,
    new_y_mux_43, new_s__state_25, new_not_s__state_25, new_I0__state_25,
    new_I1__state_25, new_and_mux__state_25, new_and_mux__state_25_2,
    new_y_mux_44, new_s__state_27, new_not_s__state_27, new_I0__state_27,
    new_I1__state_27, new_and_mux__state_27, new_and_mux__state_27_2,
    new_y_mux_45, new_s__state_29, new_not_s__state_29, new_I0__state_29,
    new_I1__state_29, new_and_mux__state_29, new_and_mux__state_29_2,
    new_y_mux_46, new_s__state_31, new_not_s__state_31, new_I0__state_31,
    new_I1__state_31, new_and_mux__state_31, new_and_mux__state_31_2,
    new_y_mux_47, new_s__state_33, new_not_s__state_33, new_I0__state_33,
    new_I1__state_33, new_and_mux__state_33, new_and_mux__state_33_2,
    new_y_mux_48, new_s__state_35, new_not_s__state_35, new_I0__state_35,
    new_I1__state_35, new_and_mux__state_35, new_and_mux__state_35_2,
    new_y_mux_49, new_s__state_37, new_not_s__state_37, new_I0__state_37,
    new_I1__state_37, new_and_mux__state_37, new_and_mux__state_37_2,
    new_y_mux_50, new_s__state_39, new_not_s__state_39, new_I0__state_39,
    new_I1__state_39, new_and_mux__state_39, new_and_mux__state_39_2,
    new_y_mux_51, new_s__state_41, new_not_s__state_41, new_I0__state_41,
    new_I1__state_41, new_and_mux__state_41, new_and_mux__state_41_2,
    new_y_mux_52, new_s__state_43, new_not_s__state_43, new_I0__state_43,
    new_I1__state_43, new_and_mux__state_43, new_and_mux__state_43_2,
    new_y_mux_53, new_s__state_45, new_not_s__state_45, new_I0__state_45,
    new_I1__state_45, new_and_mux__state_45, new_and_mux__state_45_2,
    new_y_mux_54, new_s__state_47, new_not_s__state_47, new_I0__state_47,
    new_I1__state_47, new_and_mux__state_47, new_and_mux__state_47_2,
    new_y_mux_55, new_s__state_49, new_not_s__state_49, new_I0__state_49,
    new_I1__state_49, new_and_mux__state_49, new_and_mux__state_49_2,
    new_y_mux_56, new_s__state_51, new_not_s__state_51, new_I0__state_51,
    new_I1__state_51, new_and_mux__state_51, new_and_mux__state_51_2,
    new_y_mux_57, new_s__state_53, new_not_s__state_53, new_I0__state_53,
    new_I1__state_53, new_and_mux__state_53, new_and_mux__state_53_2,
    new_y_mux_58, new_s__state_55, new_not_s__state_55, new_I0__state_55,
    new_I1__state_55, new_and_mux__state_55, new_and_mux__state_55_2,
    new_y_mux_59, new_s__state_57, new_not_s__state_57, new_I0__state_57,
    new_I1__state_57, new_and_mux__state_57, new_and_mux__state_57_2,
    new_y_mux_60, new_s__state_59, new_not_s__state_59, new_I0__state_59,
    new_I1__state_59, new_and_mux__state_59, new_and_mux__state_59_2,
    new_y_mux_61, new_s__state_61, new_not_s__state_61, new_I0__state_61,
    new_I1__state_61, new_and_mux__state_61, new_and_mux__state_61_2, n174,
    n179, n184, n189, n194, n199, n204, n209, n214, n219, n224, n229, n234,
    n239, n244, n249, n254, n259, n264, n269, n274, n279, n284, n289, n294,
    n299, n304, n309, n314, n319, n324, n329, n334, n339, n344, n349, n354,
    n359, n364, n369, n374, n379, n384, n389, n394, n399, n404, n409, n414,
    n419, n424, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474,
    n479, n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534,
    n539, n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594,
    n599, n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654,
    n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714,
    n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774,
    n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834,
    n839, n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894,
    n899, n904, n909, n914, n919, n924, n929, n934, n939, n944, n949, n954,
    n959, n964, n969, n974, n979, n984, n989, n994, n999, n1004, n1009,
    n1014, n1019, n1024, n1029, n1034, n1039, n1044, n1049, n1054, n1059,
    n1064, n1069, n1074, n1079, n1084, n1089, n1094, n1099, n1104, n1109,
    n1114, n1119, n1124, n1129, n1134, n1139, n1144, n1149, n1154, n1159,
    n1164, n1169, n1174, n1179, n1184, n1189, n1194, n1199, n1204, n1209,
    n1214, n1219, n1224, n1229, n1234, n1239, n1244, n1249, n1254, n1259,
    n1264, n1269, n1274, n1279, n1284, n1289, n1294, n1299, n1304, n1309,
    n1314, n1319, n1324, n1329, n1334, n1339, n1344, n1349, n1354, n1359,
    n1364, n1369, n1374, n1379, n1384, n1389, n1394, n1399, n1404, n1409,
    n1414, n1419, n1424, n1429, n1434, n1439, n1444, n1449, n1454, n1459,
    n1464, n1469, n1474, n1479, n1484, n1489, n1494, n1499, n1504, n1509,
    n1514, n1519, n1524, n1529, n1534, n1539, n1544, n1549, n1554, n1559,
    n1564, n1569, n1574, n1579, n1584, n1589, n1594, n1599, n1604, n1609,
    n1614, n1619, n1624, n1629, n1634, n1639, n1644, n1649, n1654, n1659,
    n1664, n1669, n1674, n1679, n1684, n1689, n1694, n1699, n1704, n1709,
    n1714, n1719, n1724, n1729, n1734, n1739, n1744, n1749, n1754, n1759,
    n1764, n1769, n1774, n1779, n1784, n1789, n1794, n1799, n1804, n1809,
    n1814, n1819, n1824, n1829, n1834, n1839, n1844, n1849, n1854, n1859,
    n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899, n1904, n1909,
    n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949, n1954, n1959,
    n1964, n1969, n1974, n1979, n1984, n1989, n1994, n1999, n2004, n2009,
    n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049, n2054, n2059,
    n2064, n2069, n2074, n2079, n2084, n2089, n2094, n2099, n2104, n2109,
    n2114, n2119, n2124, n2129, n2134, n2139, n2144, n2149, n2154, n2159,
    n2164, n2169, n2174, n2179, n2184, n2189, n2194, n2199, n2204, n2209,
    n2214, n2219, n2224, n2229, n2234, n2239, n2244, n2249, n2254, n2259,
    n2264, n2269, n2274, n2279, n2284, n2289, n2294, n2299, n2304, n2309,
    n2314, n2319, n2324, n2329, n2334, n2339, n2344, n2349, n2354, n2359,
    n2364, n2369, n2374, n2379, n2384, n2389, n2394, n2399, n2404, n2409,
    n2414, n2419, n2424, n2429, n2434, n2439, n2444, n2449, n2454, n2459,
    n2464, n2469, n2474, n2479, n2484, n2489, n2494, n2499, n2504, n2509,
    n2514, n2519, n2524, n2529, n2534, n2539, n2544, n2549, n2554, n2559,
    n2564, n2569, n2574, n2579, n2584, n2589, n2594, n2599, n2604, n2609,
    n2614, n2619, n2624, n2629, n2634, n2639, n2644, n2649, n2654, n2659,
    n2664, n2669, n2674, n2679, n2684, n2689, n2694, n2699, n2704, n2709,
    n2714, n2719, n2724, n2729, n2734, n2739, n2744, n2749, n2754, n2759,
    n2764, n2769, n2774, n2779, n2784, n2789, n2794, n2799, n2804, n2809,
    n2814, n2819, n2824, n2829, n2834, n2839, n2844, n2849, n2854, n2859,
    n2864, n2869, n2874, n2879, n2884, n2889, n2894, n2899, n2904, n2909,
    n2914, n2919, n2924, n2929, n2934, n2939, n2944, n2949, n2954, n2959,
    n2964, n2969, n2974, n2979, n2984, n2989, n2994, n2999, n3004, n3009,
    n3014, n3019, n3024, n3029, n3034, n3039, n3044, n3049, n3054, n3059,
    n3064, n3069, n3074, n3079, n3084, n3089, n3094, n3099, n3104, n3109,
    n3114, n3119, n3124, n3129, n3134, n3139, n3144, n3149, n3154, n3159,
    n3164, n3169, n3174, n3179, n3184, n3189, n3194, n3199, n3204, n3209,
    n3214, n3219, n3224, n3229, n3234, n3239, n3244, n3249, n3254, n3259,
    n3264, n3269, n3274, n3279, n3284, n3289, n3294, n3299, n3304, n3309,
    n3314, n3319, n3324, n3329, n3334, n3339, n3344, n3349, n3354, n3359,
    n3364, n3369, n3374, n3379, n3384, n3389, n3394, n3399, n3404, n3409,
    n3414, n3419, n3424, n3429, n3434, n3439, n3444, n3449, n3454, n3459,
    n3464, n3469, n3474, n3479, n3484, n3489, n3494, n3499, n3504, n3509,
    n3514, n3519, n3524, n3529, n3534, n3539, n3544, n3549, n3554, n3559,
    n3564, n3569, n3574, n3579, n3584, n3589, n3594, n3599, n3604, n3609,
    n3614, n3619, n3624, n3629, n3634, n3639, n3644, n3649, n3654, n3659,
    n3664, n3669, n3674, n3679, n3684, n3689, n3694, n3699, n3704, n3709,
    n3714, n3719, n3724, n3729, n3734, n3739, n3744, n3749, n3754, n3759,
    n3764, n3769, n3774, n3779, n3784, n3789, n3794, n3799, n3804, n3809,
    n3814, n3819, n3824, n3829, n3834, n3839, n3844, n61551, n61554,
    n61557, n61560, n61563;
  assign new_P3_R1161_U504 = ~new_P3_U3387 | ~new_P3_R1161_U30;
  assign new_P3_R1161_U503 = ~new_P3_U3076 | ~new_P3_R1161_U29;
  assign new_P3_R1161_U502 = ~new_P3_U3419 | ~new_P3_R1161_U62;
  assign U28 = P3_WR_REG | new_U160;
  assign U29 = P3_RD_REG | new_U163;
  assign new_U30 = ~new_U173 | ~new_U172;
  assign new_U31 = ~new_U175 | ~new_U174;
  assign new_U32 = ~new_U177 | ~new_U176;
  assign new_U33 = ~new_U179 | ~new_U178;
  assign new_U34 = ~new_U181 | ~new_U180;
  assign new_U35 = ~new_U183 | ~new_U182;
  assign new_U36 = ~new_U185 | ~new_U184;
  assign new_U37 = ~new_U187 | ~new_U186;
  assign new_U38 = ~new_U189 | ~new_U188;
  assign new_U39 = ~new_U191 | ~new_U190;
  assign new_U40 = ~new_U193 | ~new_U192;
  assign new_U41 = ~new_U195 | ~new_U194;
  assign new_U42 = ~new_U197 | ~new_U196;
  assign new_U43 = ~new_U199 | ~new_U198;
  assign new_U44 = ~new_U201 | ~new_U200;
  assign new_U45 = ~new_U203 | ~new_U202;
  assign new_U46 = ~new_U205 | ~new_U204;
  assign new_U47 = ~new_U207 | ~new_U206;
  assign new_U48 = ~new_U209 | ~new_U208;
  assign new_U49 = ~new_U211 | ~new_U210;
  assign new_U50 = ~new_U213 | ~new_U212;
  assign new_U51 = ~new_U215 | ~new_U214;
  assign new_U52 = ~new_U217 | ~new_U216;
  assign new_U53 = ~new_U219 | ~new_U218;
  assign new_U54 = ~new_U221 | ~new_U220;
  assign new_U55 = ~new_U223 | ~new_U222;
  assign new_U56 = ~new_U225 | ~new_U224;
  assign new_U57 = ~new_U227 | ~new_U226;
  assign new_U58 = ~new_U229 | ~new_U228;
  assign new_U59 = ~new_U231 | ~new_U230;
  assign new_U60 = ~new_U233 | ~new_U232;
  assign new_U61 = ~new_U235 | ~new_U234;
  assign new_U62 = ~new_U237 | ~new_U236;
  assign new_U63 = ~new_U239 | ~new_U238;
  assign new_U64 = ~new_U241 | ~new_U240;
  assign new_U65 = ~new_U243 | ~new_U242;
  assign new_U66 = ~new_U245 | ~new_U244;
  assign new_U67 = ~new_U247 | ~new_U246;
  assign new_U68 = ~new_U249 | ~new_U248;
  assign new_U69 = ~new_U251 | ~new_U250;
  assign new_U70 = ~new_U253 | ~new_U252;
  assign new_U71 = ~new_U255 | ~new_U254;
  assign new_U72 = ~new_U257 | ~new_U256;
  assign new_U73 = ~new_U259 | ~new_U258;
  assign new_U74 = ~new_U261 | ~new_U260;
  assign new_U75 = ~new_U263 | ~new_U262;
  assign new_U76 = ~new_U265 | ~new_U264;
  assign new_U77 = ~new_U267 | ~new_U266;
  assign new_U78 = ~new_U269 | ~new_U268;
  assign new_U79 = ~new_U271 | ~new_U270;
  assign new_U80 = ~new_U273 | ~new_U272;
  assign new_U81 = ~new_U275 | ~new_U274;
  assign new_U82 = ~new_U277 | ~new_U276;
  assign new_U83 = ~new_U279 | ~new_U278;
  assign new_U84 = ~new_U281 | ~new_U280;
  assign new_U85 = ~new_U283 | ~new_U282;
  assign new_U86 = ~new_U285 | ~new_U284;
  assign new_U87 = ~new_U287 | ~new_U286;
  assign new_U88 = ~new_U289 | ~new_U288;
  assign new_U89 = ~new_U291 | ~new_U290;
  assign new_U90 = ~new_U293 | ~new_U292;
  assign new_U91 = ~new_U295 | ~new_U294;
  assign new_U92 = ~new_U297 | ~new_U296;
  assign new_U93 = ~new_U299 | ~new_U298;
  assign new_U94 = ~new_U301 | ~new_U300;
  assign new_U95 = ~new_U303 | ~new_U302;
  assign new_U96 = ~new_U305 | ~new_U304;
  assign new_U97 = ~new_U307 | ~new_U306;
  assign new_U98 = ~new_U309 | ~new_U308;
  assign new_U99 = ~new_U311 | ~new_U310;
  assign new_U100 = ~new_U313 | ~new_U312;
  assign new_U101 = ~new_U315 | ~new_U314;
  assign new_U102 = ~new_U317 | ~new_U316;
  assign new_U103 = ~new_U319 | ~new_U318;
  assign new_U104 = ~new_U321 | ~new_U320;
  assign new_U105 = ~new_U323 | ~new_U322;
  assign new_U106 = ~new_U325 | ~new_U324;
  assign new_U107 = ~new_U327 | ~new_U326;
  assign new_U108 = ~new_U329 | ~new_U328;
  assign new_U109 = ~new_U331 | ~new_U330;
  assign new_U110 = ~new_U333 | ~new_U332;
  assign new_U111 = ~new_U335 | ~new_U334;
  assign new_U112 = ~new_U337 | ~new_U336;
  assign new_U113 = ~new_U339 | ~new_U338;
  assign new_U114 = ~new_U341 | ~new_U340;
  assign new_U115 = ~new_U343 | ~new_U342;
  assign new_U116 = ~new_U345 | ~new_U344;
  assign new_U117 = ~new_U347 | ~new_U346;
  assign new_U118 = ~new_U349 | ~new_U348;
  assign new_U119 = ~new_U351 | ~new_U350;
  assign new_U120 = ~new_U353 | ~new_U352;
  assign new_U121 = ~new_U355 | ~new_U354;
  assign new_U122 = ~new_U357 | ~new_U356;
  assign new_U123 = ~new_U359 | ~new_U358;
  assign new_U124 = ~new_U361 | ~new_U360;
  assign new_U125 = ~new_U363 | ~new_U362;
  assign new_U126 = ~new_U365 | ~new_U364;
  assign new_U127 = ~new_U367 | ~new_U366;
  assign new_U128 = ~new_U369 | ~new_U368;
  assign new_U129 = ~new_U371 | ~new_U370;
  assign new_U130 = ~new_U373 | ~new_U372;
  assign new_U131 = ~new_U375 | ~new_U374;
  assign new_U132 = ~new_U377 | ~new_U376;
  assign new_U133 = ~new_U379 | ~new_U378;
  assign new_U134 = ~new_U381 | ~new_U380;
  assign new_U135 = ~new_U383 | ~new_U382;
  assign new_U136 = ~new_U385 | ~new_U384;
  assign new_U137 = ~new_U387 | ~new_U386;
  assign new_U138 = ~new_U389 | ~new_U388;
  assign new_U139 = ~new_U391 | ~new_U390;
  assign new_U140 = ~new_U393 | ~new_U392;
  assign new_U141 = ~new_U395 | ~new_U394;
  assign new_U142 = ~new_U397 | ~new_U396;
  assign new_U143 = ~new_U399 | ~new_U398;
  assign new_U144 = ~new_U401 | ~new_U400;
  assign new_U145 = ~new_U403 | ~new_U402;
  assign new_U146 = ~new_U405 | ~new_U404;
  assign new_U147 = ~new_U407 | ~new_U406;
  assign new_U148 = ~new_U409 | ~new_U408;
  assign new_U149 = ~new_U411 | ~new_U410;
  assign new_U150 = ~new_U413 | ~new_U412;
  assign new_U151 = ~new_U415 | ~new_U414;
  assign new_U152 = ~new_U417 | ~new_U416;
  assign new_U153 = ~new_U419 | ~new_U418;
  assign new_U154 = ~new_U421 | ~new_U420;
  assign new_U155 = ~new_U423 | ~new_U422;
  assign new_U156 = ~new_U425 | ~new_U424;
  assign new_U157 = ~new_U427 | ~new_U426;
  assign new_U158 = ~P2_WR_REG;
  assign new_U159 = ~P1_WR_REG;
  assign new_U160 = new_U169 & new_U168;
  assign new_U161 = ~P2_RD_REG;
  assign new_U162 = ~P1_RD_REG;
  assign new_U163 = new_U171 & new_U170;
  assign new_U164 = ~new_U166 | ~new_U165;
  assign new_U165 = ~new_U161 | ~new_LT_1602_U6 | ~P1_ADDR_REG_19_ | ~P2_ADDR_REG_19_;
  assign new_U166 = ~new_U162 | ~P3_ADDR_REG_19_ | ~new_LT_1601_U6 | ~new_LT_1601_21_U6;
  assign new_U167 = ~new_U164;
  assign new_U168 = ~P2_WR_REG | ~new_U159;
  assign new_U169 = ~P1_WR_REG | ~new_U158;
  assign new_U170 = ~P2_RD_REG | ~new_U162;
  assign new_U171 = ~P1_RD_REG | ~new_U161;
  assign new_U172 = ~new_SUB_1605_U79 | ~new_U164;
  assign new_U173 = ~SI_9_ | ~new_U167;
  assign new_U174 = ~new_SUB_1605_U80 | ~new_U164;
  assign new_U175 = ~SI_8_ | ~new_U167;
  assign new_U176 = ~new_SUB_1605_U81 | ~new_U164;
  assign new_U177 = ~SI_7_ | ~new_U167;
  assign new_U178 = ~new_SUB_1605_U82 | ~new_U164;
  assign new_U179 = ~SI_6_ | ~new_U167;
  assign new_U180 = ~new_SUB_1605_U83 | ~new_U164;
  assign new_U181 = ~SI_5_ | ~new_U167;
  assign new_U182 = ~new_SUB_1605_U84 | ~new_U164;
  assign new_U183 = ~SI_4_ | ~new_U167;
  assign new_U184 = ~new_SUB_1605_U85 | ~new_U164;
  assign new_U185 = ~SI_3_ | ~new_U167;
  assign new_U186 = ~new_SUB_1605_U12 | ~new_U164;
  assign new_U187 = ~SI_31_ | ~new_U167;
  assign new_U188 = ~new_SUB_1605_U86 | ~new_U164;
  assign new_U189 = ~SI_30_ | ~new_U167;
  assign new_U190 = ~new_SUB_1605_U87 | ~new_U164;
  assign new_U191 = ~SI_2_ | ~new_U167;
  assign new_U192 = ~new_SUB_1605_U88 | ~new_U164;
  assign new_U193 = ~SI_29_ | ~new_U167;
  assign new_U194 = ~new_SUB_1605_U89 | ~new_U164;
  assign new_U195 = ~SI_28_ | ~new_U167;
  assign new_U196 = ~new_SUB_1605_U90 | ~new_U164;
  assign new_U197 = ~SI_27_ | ~new_U167;
  assign new_U198 = ~new_SUB_1605_U91 | ~new_U164;
  assign new_U199 = ~SI_26_ | ~new_U167;
  assign new_U200 = ~new_SUB_1605_U92 | ~new_U164;
  assign new_U201 = ~SI_25_ | ~new_U167;
  assign new_U202 = ~new_SUB_1605_U93 | ~new_U164;
  assign new_U203 = ~SI_24_ | ~new_U167;
  assign new_U204 = ~new_SUB_1605_U94 | ~new_U164;
  assign new_U205 = ~SI_23_ | ~new_U167;
  assign new_U206 = ~new_SUB_1605_U95 | ~new_U164;
  assign new_U207 = ~SI_22_ | ~new_U167;
  assign new_U208 = ~new_SUB_1605_U96 | ~new_U164;
  assign new_U209 = ~SI_21_ | ~new_U167;
  assign new_U210 = ~new_SUB_1605_U97 | ~new_U164;
  assign new_U211 = ~SI_20_ | ~new_U167;
  assign new_U212 = ~new_SUB_1605_U98 | ~new_U164;
  assign new_U213 = ~SI_1_ | ~new_U167;
  assign new_U214 = ~new_SUB_1605_U99 | ~new_U164;
  assign new_U215 = ~SI_19_ | ~new_U167;
  assign new_U216 = ~new_SUB_1605_U100 | ~new_U164;
  assign new_U217 = ~SI_18_ | ~new_U167;
  assign new_U218 = ~new_SUB_1605_U101 | ~new_U164;
  assign new_U219 = ~SI_17_ | ~new_U167;
  assign new_U220 = ~new_SUB_1605_U102 | ~new_U164;
  assign new_U221 = ~SI_16_ | ~new_U167;
  assign new_U222 = ~new_SUB_1605_U103 | ~new_U164;
  assign new_U223 = ~SI_15_ | ~new_U167;
  assign new_U224 = ~new_SUB_1605_U104 | ~new_U164;
  assign new_U225 = ~SI_14_ | ~new_U167;
  assign new_U226 = ~new_SUB_1605_U105 | ~new_U164;
  assign new_U227 = ~SI_13_ | ~new_U167;
  assign new_U228 = ~new_SUB_1605_U106 | ~new_U164;
  assign new_U229 = ~SI_12_ | ~new_U167;
  assign new_U230 = ~new_SUB_1605_U107 | ~new_U164;
  assign new_U231 = ~SI_11_ | ~new_U167;
  assign new_U232 = ~new_SUB_1605_U108 | ~new_U164;
  assign new_U233 = ~SI_10_ | ~new_U167;
  assign new_U234 = ~new_SUB_1605_U13 | ~new_U164;
  assign new_U235 = ~SI_0_ | ~new_U167;
  assign new_U236 = ~P1_DATAO_REG_9_ | ~new_U164;
  assign new_U237 = ~new_R152_U85 | ~new_U167;
  assign new_U238 = ~P1_DATAO_REG_8_ | ~new_U164;
  assign new_U239 = ~new_R152_U86 | ~new_U167;
  assign new_U240 = ~P1_DATAO_REG_7_ | ~new_U164;
  assign new_U241 = ~new_R152_U87 | ~new_U167;
  assign new_U242 = ~P1_DATAO_REG_6_ | ~new_U164;
  assign new_U243 = ~new_R152_U88 | ~new_U167;
  assign new_U244 = ~P1_DATAO_REG_5_ | ~new_U164;
  assign new_U245 = ~new_R152_U89 | ~new_U167;
  assign new_U246 = ~P1_DATAO_REG_4_ | ~new_U164;
  assign new_U247 = ~new_R152_U90 | ~new_U167;
  assign new_U248 = ~P1_DATAO_REG_3_ | ~new_U164;
  assign new_U249 = ~new_R152_U91 | ~new_U167;
  assign new_U250 = ~P1_DATAO_REG_31_ | ~new_U164;
  assign new_U251 = ~new_R152_U12 | ~new_U167;
  assign new_U252 = ~P1_DATAO_REG_30_ | ~new_U164;
  assign new_U253 = ~new_R152_U92 | ~new_U167;
  assign new_U254 = ~P1_DATAO_REG_2_ | ~new_U164;
  assign new_U255 = ~new_R152_U93 | ~new_U167;
  assign new_U256 = ~P1_DATAO_REG_29_ | ~new_U164;
  assign new_U257 = ~new_R152_U94 | ~new_U167;
  assign new_U258 = ~P1_DATAO_REG_28_ | ~new_U164;
  assign new_U259 = ~new_R152_U95 | ~new_U167;
  assign new_U260 = ~P1_DATAO_REG_27_ | ~new_U164;
  assign new_U261 = ~new_R152_U96 | ~new_U167;
  assign new_U262 = ~P1_DATAO_REG_26_ | ~new_U164;
  assign new_U263 = ~new_R152_U97 | ~new_U167;
  assign new_U264 = ~P1_DATAO_REG_25_ | ~new_U164;
  assign new_U265 = ~new_R152_U98 | ~new_U167;
  assign new_U266 = ~P1_DATAO_REG_24_ | ~new_U164;
  assign new_U267 = ~new_R152_U99 | ~new_U167;
  assign new_U268 = ~P1_DATAO_REG_23_ | ~new_U164;
  assign new_U269 = ~new_R152_U100 | ~new_U167;
  assign new_U270 = ~P1_DATAO_REG_22_ | ~new_U164;
  assign new_U271 = ~new_R152_U101 | ~new_U167;
  assign new_U272 = ~P1_DATAO_REG_21_ | ~new_U164;
  assign new_U273 = ~new_R152_U102 | ~new_U167;
  assign new_U274 = ~P1_DATAO_REG_20_ | ~new_U164;
  assign new_U275 = ~new_R152_U103 | ~new_U167;
  assign new_U276 = ~P1_DATAO_REG_1_ | ~new_U164;
  assign new_U277 = ~new_R152_U13 | ~new_U167;
  assign new_U278 = ~P1_DATAO_REG_19_ | ~new_U164;
  assign new_U279 = ~new_R152_U104 | ~new_U167;
  assign new_U280 = ~P1_DATAO_REG_18_ | ~new_U164;
  assign new_U281 = ~new_R152_U105 | ~new_U167;
  assign new_U282 = ~P1_DATAO_REG_17_ | ~new_U164;
  assign new_U283 = ~new_R152_U106 | ~new_U167;
  assign new_U284 = ~P1_DATAO_REG_16_ | ~new_U164;
  assign new_U285 = ~new_R152_U107 | ~new_U167;
  assign new_U286 = ~P1_DATAO_REG_15_ | ~new_U164;
  assign new_U287 = ~new_R152_U108 | ~new_U167;
  assign new_U288 = ~P1_DATAO_REG_14_ | ~new_U164;
  assign new_U289 = ~new_R152_U109 | ~new_U167;
  assign new_U290 = ~P1_DATAO_REG_13_ | ~new_U164;
  assign new_U291 = ~new_R152_U110 | ~new_U167;
  assign new_U292 = ~P1_DATAO_REG_12_ | ~new_U164;
  assign new_U293 = ~new_R152_U111 | ~new_U167;
  assign new_U294 = ~P1_DATAO_REG_11_ | ~new_U164;
  assign new_U295 = ~new_R152_U112 | ~new_U167;
  assign new_U296 = ~P1_DATAO_REG_10_ | ~new_U164;
  assign new_U297 = ~new_R152_U113 | ~new_U167;
  assign new_U298 = ~P1_DATAO_REG_0_ | ~new_U164;
  assign new_U299 = ~new_R152_U84 | ~new_U167;
  assign new_U300 = ~new_R152_U85 | ~new_U164;
  assign new_U301 = ~P2_DATAO_REG_9_ | ~new_U167;
  assign new_U302 = ~new_R152_U86 | ~new_U164;
  assign new_U303 = ~P2_DATAO_REG_8_ | ~new_U167;
  assign new_U304 = ~new_R152_U87 | ~new_U164;
  assign new_U305 = ~P2_DATAO_REG_7_ | ~new_U167;
  assign new_U306 = ~new_R152_U88 | ~new_U164;
  assign new_U307 = ~P2_DATAO_REG_6_ | ~new_U167;
  assign new_U308 = ~new_R152_U89 | ~new_U164;
  assign new_U309 = ~P2_DATAO_REG_5_ | ~new_U167;
  assign new_U310 = ~new_R152_U90 | ~new_U164;
  assign new_U311 = ~P2_DATAO_REG_4_ | ~new_U167;
  assign new_U312 = ~new_R152_U91 | ~new_U164;
  assign new_U313 = ~P2_DATAO_REG_3_ | ~new_U167;
  assign new_U314 = ~new_R152_U12 | ~new_U164;
  assign new_U315 = ~P2_DATAO_REG_31_ | ~new_U167;
  assign new_U316 = ~new_R152_U92 | ~new_U164;
  assign new_U317 = ~P2_DATAO_REG_30_ | ~new_U167;
  assign new_U318 = ~new_R152_U93 | ~new_U164;
  assign new_U319 = ~P2_DATAO_REG_2_ | ~new_U167;
  assign new_U320 = ~new_R152_U94 | ~new_U164;
  assign new_U321 = ~P2_DATAO_REG_29_ | ~new_U167;
  assign new_U322 = ~new_R152_U95 | ~new_U164;
  assign new_U323 = ~P2_DATAO_REG_28_ | ~new_U167;
  assign new_U324 = ~new_R152_U96 | ~new_U164;
  assign new_U325 = ~P2_DATAO_REG_27_ | ~new_U167;
  assign new_U326 = ~new_R152_U97 | ~new_U164;
  assign new_U327 = ~P2_DATAO_REG_26_ | ~new_U167;
  assign new_U328 = ~new_R152_U98 | ~new_U164;
  assign new_U329 = ~P2_DATAO_REG_25_ | ~new_U167;
  assign new_U330 = ~new_R152_U99 | ~new_U164;
  assign new_U331 = ~P2_DATAO_REG_24_ | ~new_U167;
  assign new_U332 = ~new_R152_U100 | ~new_U164;
  assign new_U333 = ~P2_DATAO_REG_23_ | ~new_U167;
  assign new_U334 = ~new_R152_U101 | ~new_U164;
  assign new_U335 = ~P2_DATAO_REG_22_ | ~new_U167;
  assign new_U336 = ~new_R152_U102 | ~new_U164;
  assign new_U337 = ~P2_DATAO_REG_21_ | ~new_U167;
  assign new_U338 = ~new_R152_U103 | ~new_U164;
  assign new_U339 = ~P2_DATAO_REG_20_ | ~new_U167;
  assign new_U340 = ~new_R152_U13 | ~new_U164;
  assign new_U341 = ~P2_DATAO_REG_1_ | ~new_U167;
  assign new_U342 = ~new_R152_U104 | ~new_U164;
  assign new_U343 = ~P2_DATAO_REG_19_ | ~new_U167;
  assign new_U344 = ~new_R152_U105 | ~new_U164;
  assign new_U345 = ~P2_DATAO_REG_18_ | ~new_U167;
  assign new_U346 = ~new_R152_U106 | ~new_U164;
  assign new_U347 = ~P2_DATAO_REG_17_ | ~new_U167;
  assign new_U348 = ~new_R152_U107 | ~new_U164;
  assign new_U349 = ~P2_DATAO_REG_16_ | ~new_U167;
  assign new_U350 = ~new_R152_U108 | ~new_U164;
  assign new_U351 = ~P2_DATAO_REG_15_ | ~new_U167;
  assign new_U352 = ~new_R152_U109 | ~new_U164;
  assign new_U353 = ~P2_DATAO_REG_14_ | ~new_U167;
  assign new_U354 = ~new_R152_U110 | ~new_U164;
  assign new_U355 = ~P2_DATAO_REG_13_ | ~new_U167;
  assign new_U356 = ~new_R152_U111 | ~new_U164;
  assign new_U357 = ~P2_DATAO_REG_12_ | ~new_U167;
  assign new_U358 = ~new_R152_U112 | ~new_U164;
  assign new_U359 = ~P2_DATAO_REG_11_ | ~new_U167;
  assign new_U360 = ~new_R152_U113 | ~new_U164;
  assign new_U361 = ~P2_DATAO_REG_10_ | ~new_U167;
  assign new_U362 = ~new_R152_U84 | ~new_U164;
  assign new_U363 = ~P2_DATAO_REG_0_ | ~new_U167;
  assign new_U364 = ~P2_DATAO_REG_9_ | ~new_U164;
  assign new_U365 = ~P1_DATAO_REG_9_ | ~new_U167;
  assign new_U366 = ~P2_DATAO_REG_8_ | ~new_U164;
  assign new_U367 = ~P1_DATAO_REG_8_ | ~new_U167;
  assign new_U368 = ~P2_DATAO_REG_7_ | ~new_U164;
  assign new_U369 = ~P1_DATAO_REG_7_ | ~new_U167;
  assign new_U370 = ~P2_DATAO_REG_6_ | ~new_U164;
  assign new_U371 = ~P1_DATAO_REG_6_ | ~new_U167;
  assign new_U372 = ~P2_DATAO_REG_5_ | ~new_U164;
  assign new_U373 = ~P1_DATAO_REG_5_ | ~new_U167;
  assign new_U374 = ~P2_DATAO_REG_4_ | ~new_U164;
  assign new_U375 = ~P1_DATAO_REG_4_ | ~new_U167;
  assign new_U376 = ~P2_DATAO_REG_31_ | ~new_U164;
  assign new_U377 = ~P1_DATAO_REG_31_ | ~new_U167;
  assign new_U378 = ~P2_DATAO_REG_30_ | ~new_U164;
  assign new_U379 = ~P1_DATAO_REG_30_ | ~new_U167;
  assign new_U380 = ~P2_DATAO_REG_3_ | ~new_U164;
  assign new_U381 = ~P1_DATAO_REG_3_ | ~new_U167;
  assign new_U382 = ~P2_DATAO_REG_29_ | ~new_U164;
  assign new_U383 = ~P1_DATAO_REG_29_ | ~new_U167;
  assign new_U384 = ~P2_DATAO_REG_28_ | ~new_U164;
  assign new_U385 = ~P1_DATAO_REG_28_ | ~new_U167;
  assign new_U386 = ~P2_DATAO_REG_27_ | ~new_U164;
  assign new_U387 = ~P1_DATAO_REG_27_ | ~new_U167;
  assign new_U388 = ~P2_DATAO_REG_26_ | ~new_U164;
  assign new_U389 = ~P1_DATAO_REG_26_ | ~new_U167;
  assign new_U390 = ~P2_DATAO_REG_25_ | ~new_U164;
  assign new_U391 = ~P1_DATAO_REG_25_ | ~new_U167;
  assign new_U392 = ~P2_DATAO_REG_24_ | ~new_U164;
  assign new_U393 = ~P1_DATAO_REG_24_ | ~new_U167;
  assign new_U394 = ~P2_DATAO_REG_23_ | ~new_U164;
  assign new_U395 = ~P1_DATAO_REG_23_ | ~new_U167;
  assign new_U396 = ~P2_DATAO_REG_22_ | ~new_U164;
  assign new_U397 = ~P1_DATAO_REG_22_ | ~new_U167;
  assign new_U398 = ~P2_DATAO_REG_21_ | ~new_U164;
  assign new_U399 = ~P1_DATAO_REG_21_ | ~new_U167;
  assign new_U400 = ~P2_DATAO_REG_20_ | ~new_U164;
  assign new_U401 = ~P1_DATAO_REG_20_ | ~new_U167;
  assign new_U402 = ~P2_DATAO_REG_2_ | ~new_U164;
  assign new_U403 = ~P1_DATAO_REG_2_ | ~new_U167;
  assign new_U404 = ~P2_DATAO_REG_19_ | ~new_U164;
  assign new_U405 = ~P1_DATAO_REG_19_ | ~new_U167;
  assign new_U406 = ~P2_DATAO_REG_18_ | ~new_U164;
  assign new_U407 = ~P1_DATAO_REG_18_ | ~new_U167;
  assign new_U408 = ~P2_DATAO_REG_17_ | ~new_U164;
  assign new_U409 = ~P1_DATAO_REG_17_ | ~new_U167;
  assign new_U410 = ~P2_DATAO_REG_16_ | ~new_U164;
  assign new_U411 = ~P1_DATAO_REG_16_ | ~new_U167;
  assign new_U412 = ~P2_DATAO_REG_15_ | ~new_U164;
  assign new_U413 = ~P1_DATAO_REG_15_ | ~new_U167;
  assign new_U414 = ~P2_DATAO_REG_14_ | ~new_U164;
  assign new_U415 = ~P1_DATAO_REG_14_ | ~new_U167;
  assign new_U416 = ~P2_DATAO_REG_13_ | ~new_U164;
  assign new_U417 = ~P1_DATAO_REG_13_ | ~new_U167;
  assign new_U418 = ~P2_DATAO_REG_12_ | ~new_U164;
  assign new_U419 = ~P1_DATAO_REG_12_ | ~new_U167;
  assign new_U420 = ~P2_DATAO_REG_11_ | ~new_U164;
  assign new_U421 = ~P1_DATAO_REG_11_ | ~new_U167;
  assign new_U422 = ~P2_DATAO_REG_10_ | ~new_U164;
  assign new_U423 = ~P1_DATAO_REG_10_ | ~new_U167;
  assign new_U424 = ~P2_DATAO_REG_1_ | ~new_U164;
  assign new_U425 = ~P1_DATAO_REG_1_ | ~new_U167;
  assign new_U426 = ~P2_DATAO_REG_0_ | ~new_U164;
  assign new_U427 = ~P1_DATAO_REG_0_ | ~new_U167;
  assign new_P3_R1161_U501 = ~new_P3_U3061 | ~new_P3_R1161_U61;
  assign new_P3_R1161_U500 = ~new_P3_R1161_U244 | ~new_P3_R1161_U498;
  assign new_P3_R1161_U499 = ~new_P3_R1161_U363 | ~new_P3_R1161_U167;
  assign new_P3_R1161_U498 = ~new_P3_R1161_U497 | ~new_P3_R1161_U496;
  assign new_P3_R1161_U497 = ~new_P3_U3422 | ~new_P3_R1161_U67;
  assign new_P3_R1161_U496 = ~new_P3_U3062 | ~new_P3_R1161_U66;
  assign new_P3_R1161_U495 = ~new_P3_R1161_U493 | ~new_P3_R1161_U338;
  assign new_P3_R1161_U494 = ~new_P3_R1161_U362 | ~new_P3_R1161_U93;
  assign new_P3_R1161_U493 = ~new_P3_R1161_U492 | ~new_P3_R1161_U491;
  assign new_P3_R1161_U492 = ~new_P3_U3425 | ~new_P3_R1161_U65;
  assign new_P3_R1161_U491 = ~new_P3_U3071 | ~new_P3_R1161_U64;
  assign new_P3_R1161_U490 = ~new_P3_U3428 | ~new_P3_R1161_U70;
  assign new_P1_U3014 = new_P1_U4002 & new_P1_U3451;
  assign new_P1_U3015 = new_P1_U3455 & new_P1_U3449;
  assign new_P1_U3016 = new_P1_U3605 & new_P1_U3600;
  assign new_P1_U3017 = new_P1_U3447 & new_P1_U3448;
  assign new_P1_U3018 = new_P1_U5808 & new_P1_U3447;
  assign new_P1_U3019 = new_P1_U5805 & new_P1_U3448;
  assign new_P1_U3020 = new_P1_U5805 & new_P1_U5808;
  assign new_P1_U3021 = new_P1_U5412 & new_P1_U3425;
  assign new_P1_U3022 = new_P1_U3592 & new_P1_U3425;
  assign new_P1_U3023 = new_P1_U4043 & new_P1_U3428;
  assign new_P1_U3024 = new_P1_U3048 & new_P1_U5793;
  assign new_P1_U3025 = new_P1_U4030 & new_P1_U5811;
  assign new_P1_U3026 = new_P1_U3851 & new_P1_U4015;
  assign new_P1_U3027 = new_P1_R1352_U6 & new_P1_U3437;
  assign new_P1_U3028 = new_P1_R1352_U6 & new_P1_U3440;
  assign new_P1_U3029 = new_P1_U3357 & P1_STATE_REG;
  assign new_P1_U3030 = new_P1_U4008 & new_P1_U4031;
  assign new_P1_U3031 = new_P1_U4031 & new_P1_U3426;
  assign new_P1_U3032 = new_P1_U4003 & new_P1_U4031;
  assign new_P1_U3033 = new_P1_U4009 & new_P1_U4031;
  assign new_P1_U3034 = new_P1_U4030 & new_P1_U3449;
  assign new_P1_U3035 = new_P1_U4015 & new_P1_U5811;
  assign new_P1_U3036 = new_P1_U4031 & new_P1_U3025;
  assign new_P1_U3037 = new_P1_U4015 & new_P1_U3449;
  assign new_P1_U3038 = new_P1_U5817 & new_P1_U4923;
  assign new_P1_U3039 = new_P1_U3023 & new_P1_U5817;
  assign new_P1_U3040 = new_P1_U5811 & new_P1_U4923;
  assign new_P1_U3041 = new_P1_U3023 & new_P1_U5811;
  assign new_P1_U3042 = new_P1_U3015 & new_P1_U4923;
  assign new_P1_U3043 = new_P1_U3023 & new_P1_U3015;
  assign new_P1_U3044 = new_P1_U3022 & new_P1_U3428;
  assign new_P1_U3045 = new_P1_U3022 & new_P1_U5159;
  assign new_P1_U3046 = new_P1_U3606 & new_P1_U3016;
  assign new_P1_U3047 = new_P1_U3452 & new_P1_U3453;
  assign new_P1_U3048 = new_P1_U5799 & new_P1_U3452;
  assign new_P1_U3049 = new_P1_U5802 & new_P1_U5796;
  assign new_P1_U3050 = new_P1_U3850 & new_P1_U5148;
  assign new_P1_U3051 = new_P1_U3419 & new_P1_U3367;
  assign new_P1_U3052 = new_P1_U3879 & new_P1_U5541 & new_P1_U3422;
  assign new_P1_U3053 = ~new_P1_U4682 | ~new_P1_U4679 | ~new_P1_U4680 | ~new_P1_U4681;
  assign new_P1_U3054 = ~new_P1_U4701 | ~new_P1_U4698 | ~new_P1_U4699 | ~new_P1_U4700;
  assign new_P1_U3055 = ~new_P1_U4717 | ~new_P1_U4718 | ~new_P1_U4720 | ~new_P1_U4719;
  assign new_P1_U3056 = ~new_P1_U4756 | ~new_P1_U4757 | ~new_P1_U4758;
  assign new_P1_U3057 = ~new_P1_U4663 | ~new_P1_U4660 | ~new_P1_U4661 | ~new_P1_U4662;
  assign new_P1_U3058 = ~new_P1_U4644 | ~new_P1_U4641 | ~new_P1_U4642 | ~new_P1_U4643;
  assign new_P1_U3059 = ~new_P1_U4736 | ~new_P1_U4737 | ~new_P1_U4738;
  assign new_P1_U3060 = ~new_P1_U4242 | ~new_P1_U4243 | ~new_P1_U4245 | ~new_P1_U4244;
  assign new_P1_U3061 = ~new_P1_U4587 | ~new_P1_U4584 | ~new_P1_U4585 | ~new_P1_U4586;
  assign new_P1_U3062 = ~new_P1_U4359 | ~new_P1_U4356 | ~new_P1_U4357 | ~new_P1_U4358;
  assign new_P1_U3063 = ~new_P1_U4378 | ~new_P1_U4375 | ~new_P1_U4376 | ~new_P1_U4377;
  assign new_P1_U3064 = ~new_P1_U4223 | ~new_P1_U4224 | ~new_P1_U4226 | ~new_P1_U4225;
  assign new_P1_U3065 = ~new_P1_U4625 | ~new_P1_U4622 | ~new_P1_U4623 | ~new_P1_U4624;
  assign new_P1_U3066 = ~new_P1_U4606 | ~new_P1_U4603 | ~new_P1_U4604 | ~new_P1_U4605;
  assign new_P1_U3067 = ~new_P1_U4261 | ~new_P1_U4262 | ~new_P1_U4264 | ~new_P1_U4263;
  assign new_P1_U3068 = ~new_P1_U4199 | ~new_P1_U4200 | ~new_P1_U4202 | ~new_P1_U4201;
  assign new_P1_U3069 = ~new_P1_U4492 | ~new_P1_U4489 | ~new_P1_U4490 | ~new_P1_U4491;
  assign new_P1_U3070 = ~new_P1_U4299 | ~new_P1_U4300 | ~new_P1_U4302 | ~new_P1_U4301;
  assign new_P1_U3071 = ~new_P1_U4280 | ~new_P1_U4281 | ~new_P1_U4283 | ~new_P1_U4282;
  assign new_P1_U3072 = ~new_P1_U4397 | ~new_P1_U4394 | ~new_P1_U4395 | ~new_P1_U4396;
  assign new_P1_U3073 = ~new_P1_U4473 | ~new_P1_U4470 | ~new_P1_U4471 | ~new_P1_U4472;
  assign new_P1_U3074 = ~new_P1_U4454 | ~new_P1_U4451 | ~new_P1_U4452 | ~new_P1_U4453;
  assign new_P1_U3075 = ~new_P1_U4568 | ~new_P1_U4565 | ~new_P1_U4566 | ~new_P1_U4567;
  assign new_P1_U3076 = ~new_P1_U4549 | ~new_P1_U4546 | ~new_P1_U4547 | ~new_P1_U4548;
  assign new_P1_U3077 = ~new_P1_U4204 | ~new_P1_U4205 | ~new_P1_U4207 | ~new_P1_U4206;
  assign new_P1_U3078 = ~new_P1_U4180 | ~new_P1_U4181 | ~new_P1_U4183 | ~new_P1_U4182;
  assign new_P1_U3079 = ~new_P1_U4435 | ~new_P1_U4432 | ~new_P1_U4433 | ~new_P1_U4434;
  assign new_P1_U3080 = ~new_P1_U4416 | ~new_P1_U4413 | ~new_P1_U4414 | ~new_P1_U4415;
  assign new_P1_U3081 = ~new_P1_U4530 | ~new_P1_U4527 | ~new_P1_U4528 | ~new_P1_U4529;
  assign new_P1_U3082 = ~new_P1_U4511 | ~new_P1_U4508 | ~new_P1_U4509 | ~new_P1_U4510;
  assign new_P1_U3083 = ~new_P1_U4340 | ~new_P1_U4337 | ~new_P1_U4338 | ~new_P1_U4339;
  assign new_P1_U3084 = ~new_P1_U4318 | ~new_P1_U4319 | ~new_P1_U4321 | ~new_P1_U4320;
  assign n1389 = ~new_P1_U4930 | ~P1_STATE_REG;
  assign n1384 = ~P1_STATE_REG;
  assign new_P1_U3087 = ~new_P1_U5667 | ~new_P1_U5668 | ~new_P1_U5666;
  assign new_P1_U3088 = ~new_P1_U5670 | ~new_P1_U5671 | ~new_P1_U5669;
  assign new_P1_U3089 = ~new_P1_U5679 | ~new_P1_U3929 | ~new_P1_U5678;
  assign new_P1_U3090 = ~new_P1_U3930 | ~new_P1_U5683 | ~new_P1_U5682;
  assign new_P1_U3091 = ~new_P1_U3931 | ~new_P1_U5687 | ~new_P1_U5686;
  assign new_P1_U3092 = ~new_P1_U3932 | ~new_P1_U5691 | ~new_P1_U5690;
  assign new_P1_U3093 = ~new_P1_U3933 | ~new_P1_U5695 | ~new_P1_U5694;
  assign new_P1_U3094 = ~new_P1_U3934 | ~new_P1_U5699 | ~new_P1_U5698;
  assign new_P1_U3095 = ~new_P1_U3935 | ~new_P1_U5703 | ~new_P1_U5702;
  assign new_P1_U3096 = ~new_P1_U3936 | ~new_P1_U5707 | ~new_P1_U5706;
  assign new_P1_U3097 = ~new_P1_U3937 | ~new_P1_U5711 | ~new_P1_U5710;
  assign new_P1_U3098 = ~new_P1_U3938 | ~new_P1_U5715 | ~new_P1_U5714;
  assign new_P1_U3099 = ~new_P1_U3940 | ~new_P1_U5723 | ~new_P1_U5722;
  assign new_P1_U3100 = ~new_P1_U3941 | ~new_P1_U5727 | ~new_P1_U5726;
  assign new_P1_U3101 = ~new_P1_U3942 | ~new_P1_U5731 | ~new_P1_U5730;
  assign new_P1_U3102 = ~new_P1_U3943 | ~new_P1_U5735 | ~new_P1_U5734;
  assign new_P1_U3103 = ~new_P1_U3944 | ~new_P1_U5739 | ~new_P1_U5738;
  assign new_P1_U3104 = ~new_P1_U3945 | ~new_P1_U5743 | ~new_P1_U5742;
  assign new_P1_U3105 = ~new_P1_U3946 | ~new_P1_U5747 | ~new_P1_U5746;
  assign new_P1_U3106 = ~new_P1_U3947 | ~new_P1_U5751 | ~new_P1_U5750;
  assign new_P1_U3107 = ~new_P1_U3948 | ~new_P1_U5755 | ~new_P1_U5754;
  assign new_P1_U3108 = ~new_P1_U3949 | ~new_P1_U5759 | ~new_P1_U5758;
  assign new_P1_U3109 = ~new_P1_U5643 | ~new_P1_U3922 | ~new_P1_U5644;
  assign new_P1_U3110 = ~new_P1_U5647 | ~new_P1_U3923 | ~new_P1_U5648;
  assign new_P1_U3111 = ~new_P1_U3924 | ~new_P1_U5653 | ~new_P1_U5652;
  assign new_P1_U3112 = ~new_P1_U3925 | ~new_P1_U5657 | ~new_P1_U5656;
  assign new_P1_U3113 = ~new_P1_U3926 | ~new_P1_U5661 | ~new_P1_U5660;
  assign new_P1_U3114 = ~new_P1_U3927 | ~new_P1_U5665 | ~new_P1_U5664;
  assign new_P1_U3115 = ~new_P1_U3928 | ~new_P1_U5674;
  assign new_P1_U3116 = ~new_P1_U3939 | ~new_P1_U5718;
  assign new_P1_U3117 = ~new_P1_U3950 | ~new_P1_U5762;
  assign new_P1_U3118 = ~new_P1_U3951 | ~new_P1_U5766;
  assign new_P1_U3119 = ~new_P1_U3892 | ~new_P1_U5563;
  assign new_P1_U3120 = ~new_P1_U3893 | ~new_P1_U5566;
  assign new_P1_U3121 = ~new_P1_U3896 | ~new_P1_U5572 | ~new_P1_U5571;
  assign new_P1_U3122 = ~new_P1_U3897 | ~new_P1_U5575 | ~new_P1_U5574;
  assign new_P1_U3123 = ~new_P1_U3898 | ~new_P1_U5578 | ~new_P1_U5577;
  assign new_P1_U3124 = ~new_P1_U3899 | ~new_P1_U5581 | ~new_P1_U5580;
  assign new_P1_U3125 = ~new_P1_U3900 | ~new_P1_U5584 | ~new_P1_U5583;
  assign new_P1_U3126 = ~new_P1_U3901 | ~new_P1_U5587 | ~new_P1_U5586;
  assign new_P1_U3127 = ~new_P1_U3902 | ~new_P1_U5590 | ~new_P1_U5589;
  assign new_P1_U3128 = ~new_P1_U3903 | ~new_P1_U5593 | ~new_P1_U5592;
  assign new_P1_U3129 = ~new_P1_U3904 | ~new_P1_U5596 | ~new_P1_U5595;
  assign new_P1_U3130 = ~new_P1_U3905 | ~new_P1_U5599 | ~new_P1_U5598;
  assign new_P1_U3131 = ~new_P1_U3908 | ~new_P1_U5605 | ~new_P1_U5604;
  assign new_P1_U3132 = ~new_P1_U3909 | ~new_P1_U5608 | ~new_P1_U5607;
  assign new_P1_U3133 = ~new_P1_U3910 | ~new_P1_U5611 | ~new_P1_U5610;
  assign new_P1_U3134 = ~new_P1_U3911 | ~new_P1_U5614 | ~new_P1_U5613;
  assign new_P1_U3135 = ~new_P1_U3912 | ~new_P1_U5617 | ~new_P1_U5616;
  assign new_P1_U3136 = ~new_P1_U3913 | ~new_P1_U5620 | ~new_P1_U5619;
  assign new_P1_U3137 = ~new_P1_U3914 | ~new_P1_U5623 | ~new_P1_U5622;
  assign new_P1_U3138 = ~new_P1_U3915 | ~new_P1_U5626 | ~new_P1_U5625;
  assign new_P1_U3139 = ~new_P1_U3916 | ~new_P1_U5629 | ~new_P1_U5628;
  assign new_P1_U3140 = ~new_P1_U3917 | ~new_P1_U5632 | ~new_P1_U5631;
  assign new_P1_U3141 = ~new_P1_U5545 | ~new_P1_U3880;
  assign new_P1_U3142 = ~new_P1_U5548 | ~new_P1_U3882;
  assign new_P1_U3143 = ~new_P1_U5551 | ~new_P1_U3884;
  assign new_P1_U3144 = ~new_P1_U5554 | ~new_P1_U3886;
  assign new_P1_U3145 = ~new_P1_U5557 | ~new_P1_U3888;
  assign new_P1_U3146 = ~new_P1_U5560 | ~new_P1_U3890;
  assign new_P1_U3147 = ~new_P1_U5569 | ~new_P1_U3894;
  assign new_P1_U3148 = ~new_P1_U5602 | ~new_P1_U3906;
  assign new_P1_U3149 = ~new_P1_U5635 | ~new_P1_U3918;
  assign new_P1_U3150 = ~new_P1_U5638 | ~new_P1_U3920;
  assign new_P1_U3151 = ~new_P1_U3877 | ~new_P1_U5537;
  assign new_P1_U3152 = ~new_P1_U3014 | ~new_P1_U5786;
  assign new_P1_U3153 = ~new_P1_U5492 | ~new_P1_U5491;
  assign new_P1_U3154 = ~new_P1_U5494 | ~new_P1_U5493;
  assign new_P1_U3155 = ~new_P1_U5496 | ~new_P1_U5495;
  assign new_P1_U3156 = ~new_P1_U5498 | ~new_P1_U5497;
  assign new_P1_U3157 = ~new_P1_U5500 | ~new_P1_U5499;
  assign new_P1_U3158 = ~new_P1_U5502 | ~new_P1_U5501;
  assign new_P1_U3159 = ~new_P1_U5504 | ~new_P1_U5503;
  assign new_P1_U3160 = ~new_P1_U5506 | ~new_P1_U5505;
  assign new_P1_U3161 = ~new_P1_U5508 | ~new_P1_U5507;
  assign new_P1_U3162 = ~new_P1_U5512 | ~new_P1_U5511;
  assign new_P1_U3163 = ~new_P1_U5514 | ~new_P1_U5513;
  assign new_P1_U3164 = ~new_P1_U5516 | ~new_P1_U5515;
  assign new_P1_U3165 = ~new_P1_U5518 | ~new_P1_U5517;
  assign new_P1_U3166 = ~new_P1_U5520 | ~new_P1_U5519;
  assign new_P1_U3167 = ~new_P1_U5522 | ~new_P1_U5521;
  assign new_P1_U3168 = ~new_P1_U5524 | ~new_P1_U5523;
  assign new_P1_U3169 = ~new_P1_U5526 | ~new_P1_U5525;
  assign new_P1_U3170 = ~new_P1_U5528 | ~new_P1_U5527;
  assign new_P1_U3171 = ~new_P1_U5530 | ~new_P1_U5529;
  assign new_P1_U3172 = ~new_P1_U5478 | ~new_P1_U5477;
  assign new_P1_U3173 = ~new_P1_U5480 | ~new_P1_U5479;
  assign new_P1_U3174 = ~new_P1_U5482 | ~new_P1_U5481;
  assign new_P1_U3175 = ~new_P1_U5484 | ~new_P1_U5483;
  assign new_P1_U3176 = ~new_P1_U5486 | ~new_P1_U5485;
  assign new_P1_U3177 = ~new_P1_U5488 | ~new_P1_U5487;
  assign new_P1_U3178 = ~new_P1_U5490 | ~new_P1_U5489;
  assign new_P1_U3179 = ~new_P1_U5510 | ~new_P1_U5509;
  assign new_P1_U3180 = ~new_P1_U5532 | ~new_P1_U5531;
  assign new_P1_U3181 = ~new_P1_U3876 | ~new_P1_U5534;
  assign new_P1_U3182 = ~new_P1_U5433 | ~new_P1_U5432;
  assign new_P1_U3183 = ~new_P1_U5435 | ~new_P1_U5434;
  assign new_P1_U3184 = ~new_P1_U5437 | ~new_P1_U5436;
  assign new_P1_U3185 = ~new_P1_U5439 | ~new_P1_U5438;
  assign new_P1_U3186 = ~new_P1_U5441 | ~new_P1_U5440;
  assign new_P1_U3187 = ~new_P1_U5443 | ~new_P1_U5442;
  assign new_P1_U3188 = ~new_P1_U5445 | ~new_P1_U5444;
  assign new_P1_U3189 = ~new_P1_U5447 | ~new_P1_U5446;
  assign new_P1_U3190 = ~new_P1_U5449 | ~new_P1_U5448;
  assign new_P1_U3191 = ~new_P1_U5453 | ~new_P1_U5452;
  assign new_P1_U3192 = ~new_P1_U5455 | ~new_P1_U5454;
  assign new_P1_U3193 = ~new_P1_U5457 | ~new_P1_U5456;
  assign new_P1_U3194 = ~new_P1_U5459 | ~new_P1_U5458;
  assign new_P1_U3195 = ~new_P1_U5461 | ~new_P1_U5460;
  assign new_P1_U3196 = ~new_P1_U5463 | ~new_P1_U5462;
  assign new_P1_U3197 = ~new_P1_U5465 | ~new_P1_U5464;
  assign new_P1_U3198 = ~new_P1_U5467 | ~new_P1_U5466;
  assign new_P1_U3199 = ~new_P1_U5469 | ~new_P1_U5468;
  assign new_P1_U3200 = ~new_P1_U5471 | ~new_P1_U5470;
  assign new_P1_U3201 = ~new_P1_U5419 | ~new_P1_U5418;
  assign new_P1_U3202 = ~new_P1_U5421 | ~new_P1_U5420;
  assign new_P1_U3203 = ~new_P1_U5423 | ~new_P1_U5422;
  assign new_P1_U3204 = ~new_P1_U5425 | ~new_P1_U5424;
  assign new_P1_U3205 = ~new_P1_U5427 | ~new_P1_U5426;
  assign new_P1_U3206 = ~new_P1_U5429 | ~new_P1_U5428;
  assign new_P1_U3207 = ~new_P1_U5431 | ~new_P1_U5430;
  assign new_P1_U3208 = ~new_P1_U5451 | ~new_P1_U5450;
  assign new_P1_U3209 = ~new_P1_U5473 | ~new_P1_U5472;
  assign new_P1_U3210 = ~new_P1_U3875 | ~new_P1_U5474;
  assign new_P1_U3211 = new_P1_U5411 & new_P1_U3425;
  assign new_P1_U3212 = ~new_P1_U5409 | ~new_P1_U6285 | ~new_P1_U6284;
  assign n1379 = ~new_P1_U5404 | ~new_P1_U3872 | ~new_P1_U5403 | ~new_P1_U5402;
  assign n1374 = ~new_P1_U5395 | ~new_P1_U5396 | ~new_P1_U5397 | ~new_P1_U5394 | ~new_P1_U5393;
  assign n1369 = ~new_P1_U5386 | ~new_P1_U5387 | ~new_P1_U5388 | ~new_P1_U5385 | ~new_P1_U5384;
  assign n1364 = ~new_P1_U5377 | ~new_P1_U5378 | ~new_P1_U5379 | ~new_P1_U5376 | ~new_P1_U5375;
  assign n1359 = ~new_P1_U5368 | ~new_P1_U3871 | ~new_P1_U5367 | ~new_P1_U5366;
  assign n1354 = ~new_P1_U3870 | ~new_P1_U3869 | ~new_P1_U5358;
  assign n1349 = ~new_P1_U5350 | ~new_P1_U5351 | ~new_P1_U5352 | ~new_P1_U5349 | ~new_P1_U5348;
  assign n1344 = ~new_P1_U5341 | ~new_P1_U5342 | ~new_P1_U5343 | ~new_P1_U5340 | ~new_P1_U5339;
  assign n1339 = ~new_P1_U5332 | ~new_P1_U3868 | ~new_P1_U5331 | ~new_P1_U5330;
  assign n1334 = ~new_P1_U3867 | ~new_P1_U3866 | ~new_P1_U5322;
  assign n1329 = ~new_P1_U5314 | ~new_P1_U5315 | ~new_P1_U5316 | ~new_P1_U5313 | ~new_P1_U5312;
  assign n1324 = ~new_P1_U5305 | ~new_P1_U3865 | ~new_P1_U5304 | ~new_P1_U5303;
  assign n1319 = ~new_P1_U5296 | ~new_P1_U5297 | ~new_P1_U5298 | ~new_P1_U5295 | ~new_P1_U5294;
  assign n1314 = ~new_P1_U5287 | ~new_P1_U5288 | ~new_P1_U5289 | ~new_P1_U5286 | ~new_P1_U5285;
  assign n1309 = ~new_P1_U3864 | ~new_P1_U5278 | ~new_P1_U5277 | ~new_P1_U5276;
  assign n1304 = ~new_P1_U5269 | ~new_P1_U5270 | ~new_P1_U5271 | ~new_P1_U5268 | ~new_P1_U5267;
  assign n1299 = ~new_P1_U5260 | ~new_P1_U5261 | ~new_P1_U5262 | ~new_P1_U5259 | ~new_P1_U5258;
  assign n1294 = ~new_P1_U3863 | ~new_P1_U3862 | ~new_P1_U5250;
  assign n1289 = ~new_P1_U5242 | ~new_P1_U3861 | ~new_P1_U5241 | ~new_P1_U5240;
  assign n1284 = ~new_P1_U5233 | ~new_P1_U3859;
  assign n1279 = ~new_P1_U5225 | ~new_P1_U5226 | ~new_P1_U5227 | ~new_P1_U5224 | ~new_P1_U5223;
  assign n1274 = ~new_P1_U5216 | ~new_P1_U3857 | ~new_P1_U5215 | ~new_P1_U5214;
  assign n1269 = ~new_P1_U5207 | ~new_P1_U5208 | ~new_P1_U5209 | ~new_P1_U5206 | ~new_P1_U5205;
  assign n1264 = ~new_P1_U5198 | ~new_P1_U3856 | ~new_P1_U5197 | ~new_P1_U5196;
  assign n1259 = ~new_P1_U3855 | ~new_P1_U3854 | ~new_P1_U5188;
  assign n1254 = ~new_P1_U5180 | ~new_P1_U5181 | ~new_P1_U5182 | ~new_P1_U5179 | ~new_P1_U5178;
  assign n1249 = ~new_P1_U5171 | ~new_P1_U3853 | ~new_P1_U5170 | ~new_P1_U5169;
  assign n1244 = ~new_P1_U5162 | ~new_P1_U5163 | ~new_P1_U5164 | ~new_P1_U5161 | ~new_P1_U5160;
  assign n1239 = ~new_P1_U5151 | ~new_P1_U5152 | ~new_P1_U5153 | ~new_P1_U5150 | ~new_P1_U5149;
  assign n1234 = ~new_P1_U3846 | ~new_P1_U5137;
  assign n1069 = ~new_P1_U3831 | ~new_P1_U3830 | ~new_P1_U5123;
  assign n1064 = ~new_P1_U3829 | ~new_P1_U3828 | ~new_P1_U5113;
  assign n1059 = ~new_P1_U3827 | ~new_P1_U5103 | ~new_P1_U3825;
  assign n1054 = ~new_P1_U3824 | ~new_P1_U3823 | ~new_P1_U5093;
  assign n1049 = ~new_P1_U3822 | ~new_P1_U5083 | ~new_P1_U3820;
  assign n1044 = ~new_P1_U3819 | ~new_P1_U3818 | ~new_P1_U5073;
  assign n1039 = ~new_P1_U5063 | ~new_P1_U3816 | ~new_P1_U3817;
  assign n1034 = ~new_P1_U5053 | ~new_P1_U3814 | ~new_P1_U3815;
  assign n1029 = ~new_P1_U5043 | ~new_P1_U3812 | ~new_P1_U3813;
  assign n1024 = ~new_P1_U5033 | ~new_P1_U3810 | ~new_P1_U3811;
  assign n1019 = ~new_P1_U5023 | ~new_P1_U3808 | ~new_P1_U3809;
  assign n1014 = ~new_P1_U5013 | ~new_P1_U3806 | ~new_P1_U3807;
  assign n1009 = ~new_P1_U5003 | ~new_P1_U3804 | ~new_P1_U3805;
  assign n1004 = ~new_P1_U4993 | ~new_P1_U3802 | ~new_P1_U3803;
  assign n999 = ~new_P1_U4983 | ~new_P1_U3800 | ~new_P1_U3801;
  assign n994 = ~new_P1_U4973 | ~new_P1_U3798 | ~new_P1_U3799;
  assign n989 = ~new_P1_U4963 | ~new_P1_U3796 | ~new_P1_U3797;
  assign n984 = ~new_P1_U4953 | ~new_P1_U3794 | ~new_P1_U3795;
  assign n979 = ~new_P1_U4943 | ~new_P1_U3792 | ~new_P1_U3793;
  assign n974 = ~new_P1_U4933 | ~new_P1_U3790 | ~new_P1_U3791;
  assign n969 = ~new_P1_U4922 | ~new_P1_U3989 | ~new_P1_U4921;
  assign n964 = ~new_P1_U4920 | ~new_P1_U3988 | ~new_P1_U4919;
  assign n954 = ~new_P1_U3985 | ~new_P1_U4912 | ~new_P1_U3784 | ~new_P1_U3785;
  assign n949 = ~new_P1_U3984 | ~new_P1_U4907 | ~new_P1_U3782 | ~new_P1_U3783;
  assign n944 = ~new_P1_U3983 | ~new_P1_U4902 | ~new_P1_U3780 | ~new_P1_U3781;
  assign n939 = ~new_P1_U3982 | ~new_P1_U4897 | ~new_P1_U3778 | ~new_P1_U3779;
  assign n934 = ~new_P1_U3981 | ~new_P1_U4892 | ~new_P1_U3776 | ~new_P1_U3777;
  assign n929 = ~new_P1_U3980 | ~new_P1_U4887 | ~new_P1_U3774 | ~new_P1_U3775;
  assign n924 = ~new_P1_U3979 | ~new_P1_U4882 | ~new_P1_U3772 | ~new_P1_U3773;
  assign n919 = ~new_P1_U3978 | ~new_P1_U4877 | ~new_P1_U3770 | ~new_P1_U3771;
  assign n914 = ~new_P1_U3977 | ~new_P1_U4872 | ~new_P1_U3768 | ~new_P1_U3769;
  assign n909 = ~new_P1_U3976 | ~new_P1_U4867 | ~new_P1_U3766 | ~new_P1_U3767;
  assign n904 = ~new_P1_U3975 | ~new_P1_U3765 | ~new_P1_U3764;
  assign n899 = ~new_P1_U3974 | ~new_P1_U3763 | ~new_P1_U3762;
  assign n894 = ~new_P1_U3973 | ~new_P1_U4852 | ~new_P1_U3760 | ~new_P1_U3761;
  assign n889 = ~new_P1_U3972 | ~new_P1_U4847 | ~new_P1_U3758 | ~new_P1_U3759;
  assign n884 = ~new_P1_U3971 | ~new_P1_U3757 | ~new_P1_U3756;
  assign n879 = ~new_P1_U3970 | ~new_P1_U3755 | ~new_P1_U3754;
  assign n874 = ~new_P1_U3969 | ~new_P1_U3753 | ~new_P1_U3752;
  assign n869 = ~new_P1_U3968 | ~new_P1_U3751 | ~new_P1_U3750;
  assign n864 = ~new_P1_U3967 | ~new_P1_U4822 | ~new_P1_U3748 | ~new_P1_U3749;
  assign n859 = ~new_P1_U3966 | ~new_P1_U4817 | ~new_P1_U3746 | ~new_P1_U3747;
  assign n854 = ~new_P1_U3965 | ~new_P1_U3745 | ~new_P1_U3744;
  assign n849 = ~new_P1_U3964 | ~new_P1_U3743 | ~new_P1_U3742;
  assign n844 = ~new_P1_U3963 | ~new_P1_U3741 | ~new_P1_U3740;
  assign n839 = ~new_P1_U3962 | ~new_P1_U3739 | ~new_P1_U3738;
  assign n834 = ~new_P1_U3737 | ~new_P1_U3736;
  assign n829 = ~new_P1_U3735 | ~new_P1_U3734;
  assign n824 = ~new_P1_U3733 | ~new_P1_U3732;
  assign n819 = ~new_P1_U3731 | ~new_P1_U3730;
  assign n814 = ~new_P1_U3729 | ~new_P1_U3728;
  assign n489 = P1_D_REG_31_ & new_P1_U3953;
  assign n484 = P1_D_REG_30_ & new_P1_U3953;
  assign n479 = P1_D_REG_29_ & new_P1_U3953;
  assign n474 = P1_D_REG_28_ & new_P1_U3953;
  assign n469 = P1_D_REG_27_ & new_P1_U3953;
  assign n464 = P1_D_REG_26_ & new_P1_U3953;
  assign n459 = P1_D_REG_25_ & new_P1_U3953;
  assign n454 = P1_D_REG_24_ & new_P1_U3953;
  assign n449 = P1_D_REG_23_ & new_P1_U3953;
  assign n444 = P1_D_REG_22_ & new_P1_U3953;
  assign n439 = P1_D_REG_21_ & new_P1_U3953;
  assign n434 = P1_D_REG_20_ & new_P1_U3953;
  assign n429 = P1_D_REG_19_ & new_P1_U3953;
  assign n424 = P1_D_REG_18_ & new_P1_U3953;
  assign n419 = P1_D_REG_17_ & new_P1_U3953;
  assign n414 = P1_D_REG_16_ & new_P1_U3953;
  assign n409 = P1_D_REG_15_ & new_P1_U3953;
  assign n404 = P1_D_REG_14_ & new_P1_U3953;
  assign n399 = P1_D_REG_13_ & new_P1_U3953;
  assign n394 = P1_D_REG_12_ & new_P1_U3953;
  assign n389 = P1_D_REG_11_ & new_P1_U3953;
  assign n384 = P1_D_REG_10_ & new_P1_U3953;
  assign n379 = P1_D_REG_9_ & new_P1_U3953;
  assign n374 = P1_D_REG_8_ & new_P1_U3953;
  assign n369 = P1_D_REG_7_ & new_P1_U3953;
  assign n364 = P1_D_REG_6_ & new_P1_U3953;
  assign n359 = P1_D_REG_5_ & new_P1_U3953;
  assign n354 = P1_D_REG_4_ & new_P1_U3953;
  assign n349 = P1_D_REG_3_ & new_P1_U3953;
  assign n344 = P1_D_REG_2_ & new_P1_U3953;
  assign n329 = ~new_P1_U4141 | ~new_P1_U4142 | ~new_P1_U4143;
  assign n324 = ~new_P1_U4138 | ~new_P1_U4139 | ~new_P1_U4140;
  assign n319 = ~new_P1_U4135 | ~new_P1_U4136 | ~new_P1_U4137;
  assign n314 = ~new_P1_U4132 | ~new_P1_U4133 | ~new_P1_U4134;
  assign n309 = ~new_P1_U4129 | ~new_P1_U4130 | ~new_P1_U4131;
  assign n304 = ~new_P1_U4126 | ~new_P1_U4127 | ~new_P1_U4128;
  assign n299 = ~new_P1_U4123 | ~new_P1_U4124 | ~new_P1_U4125;
  assign n294 = ~new_P1_U4120 | ~new_P1_U4121 | ~new_P1_U4122;
  assign n289 = ~new_P1_U4117 | ~new_P1_U4118 | ~new_P1_U4119;
  assign n284 = ~new_P1_U4114 | ~new_P1_U4115 | ~new_P1_U4116;
  assign n279 = ~new_P1_U4111 | ~new_P1_U4112 | ~new_P1_U4113;
  assign n274 = ~new_P1_U4108 | ~new_P1_U4109 | ~new_P1_U4110;
  assign n269 = ~new_P1_U4105 | ~new_P1_U4106 | ~new_P1_U4107;
  assign n264 = ~new_P1_U4102 | ~new_P1_U4103 | ~new_P1_U4104;
  assign n259 = ~new_P1_U4099 | ~new_P1_U4100 | ~new_P1_U4101;
  assign n254 = ~new_P1_U4096 | ~new_P1_U4097 | ~new_P1_U4098;
  assign n249 = ~new_P1_U4093 | ~new_P1_U4094 | ~new_P1_U4095;
  assign n244 = ~new_P1_U4090 | ~new_P1_U4091 | ~new_P1_U4092;
  assign n239 = ~new_P1_U4087 | ~new_P1_U4088 | ~new_P1_U4089;
  assign n234 = ~new_P1_U4084 | ~new_P1_U4085 | ~new_P1_U4086;
  assign n229 = ~new_P1_U4081 | ~new_P1_U4082 | ~new_P1_U4083;
  assign n224 = ~new_P1_U4078 | ~new_P1_U4079 | ~new_P1_U4080;
  assign n219 = ~new_P1_U4075 | ~new_P1_U4076 | ~new_P1_U4077;
  assign n214 = ~new_P1_U4072 | ~new_P1_U4073 | ~new_P1_U4074;
  assign n209 = ~new_P1_U4069 | ~new_P1_U4070 | ~new_P1_U4071;
  assign n204 = ~new_P1_U4066 | ~new_P1_U4067 | ~new_P1_U4068;
  assign n199 = ~new_P1_U4063 | ~new_P1_U4064 | ~new_P1_U4065;
  assign n194 = ~new_P1_U4060 | ~new_P1_U4061 | ~new_P1_U4062;
  assign n189 = ~new_P1_U4057 | ~new_P1_U4058 | ~new_P1_U4059;
  assign n184 = ~new_P1_U4054 | ~new_P1_U4055 | ~new_P1_U4056;
  assign n179 = ~new_P1_U4051 | ~new_P1_U4052 | ~new_P1_U4053;
  assign new_P1_U3355 = ~new_P1_U4048 | ~new_P1_U4049 | ~new_P1_U4050;
  assign n959 = ~new_P1_U3986 | ~new_P1_U4916 | ~new_P1_U4918 | ~new_P1_U4917 | ~new_P1_U4915;
  assign new_P1_U3357 = ~P1_STATE_REG | ~new_P1_U3952;
  assign new_P1_U3358 = ~new_P1_U3443 | ~new_P1_U5778;
  assign new_P1_U3359 = ~P1_B_REG;
  assign new_P1_U3360 = ~new_P1_U3443 | ~new_P1_U5783 | ~new_P1_U5782;
  assign new_P1_U3361 = ~new_P1_U3048 | ~new_P1_U3451;
  assign new_P1_U3362 = ~new_P1_U3047 | ~new_P1_U3451;
  assign new_P1_U3363 = ~new_P1_U3453 | ~new_P1_U5796;
  assign new_P1_U3364 = ~new_P1_U4042 | ~new_P1_U3451;
  assign new_P1_U3365 = ~new_P1_U3047 | ~new_P1_U3450;
  assign new_P1_U3366 = ~new_P1_U4042 | ~new_P1_U3450;
  assign new_P1_U3367 = ~new_P1_U3049 | ~new_P1_U3451;
  assign new_P1_U3368 = ~new_P1_U4001 | ~new_P1_U5799;
  assign new_P1_U3369 = ~new_P1_U5799 | ~new_P1_U5796;
  assign new_P1_U3370 = ~new_P1_U4044 | ~new_P1_U3450;
  assign new_P1_U3371 = ~new_P1_U4002 | ~new_P1_U5793;
  assign new_P1_U3372 = ~new_P1_U3451 | ~new_P1_U3450;
  assign new_P1_U3373 = ~new_P1_U5802 | ~new_P1_U5799 | ~new_P1_U5793;
  assign new_P1_U3374 = ~new_P1_U3049 | ~new_P1_U5793;
  assign new_P1_U3375 = ~new_P1_U5802 | ~new_P1_U3452;
  assign new_P1_U3376 = ~new_P1_U3593 | ~new_P1_U3594 | ~new_P1_U4192 | ~new_P1_U4191 | ~new_P1_U4190;
  assign new_P1_U3377 = ~P1_REG2_REG_0_;
  assign new_P1_U3378 = ~new_P1_U3610 | ~new_P1_U3608 | ~new_P1_U4210 | ~new_P1_U4209;
  assign new_P1_U3379 = ~new_P1_U3614 | ~new_P1_U3612 | ~new_P1_U4229 | ~new_P1_U4228;
  assign new_P1_U3380 = ~new_P1_U3618 | ~new_P1_U3616 | ~new_P1_U4248 | ~new_P1_U4247;
  assign new_P1_U3381 = ~new_P1_U3622 | ~new_P1_U3620 | ~new_P1_U4267 | ~new_P1_U4266;
  assign new_P1_U3382 = ~new_P1_U3626 | ~new_P1_U3624 | ~new_P1_U4286 | ~new_P1_U4285;
  assign new_P1_U3383 = ~new_P1_U3630 | ~new_P1_U3628 | ~new_P1_U4305 | ~new_P1_U4304;
  assign new_P1_U3384 = ~new_P1_U3634 | ~new_P1_U3632 | ~new_P1_U4324 | ~new_P1_U4323;
  assign new_P1_U3385 = ~new_P1_U3638 | ~new_P1_U3636 | ~new_P1_U4343 | ~new_P1_U4342;
  assign new_P1_U3386 = ~new_P1_U3642 | ~new_P1_U3640 | ~new_P1_U4362 | ~new_P1_U4361;
  assign new_P1_U3387 = ~new_P1_U3646 | ~new_P1_U3644 | ~new_P1_U4381 | ~new_P1_U4380;
  assign new_P1_U3388 = ~new_P1_U3650 | ~new_P1_U3648 | ~new_P1_U4400 | ~new_P1_U4399;
  assign new_P1_U3389 = ~new_P1_U3654 | ~new_P1_U3652 | ~new_P1_U4419 | ~new_P1_U4418;
  assign new_P1_U3390 = ~new_P1_U3658 | ~new_P1_U3656 | ~new_P1_U4438 | ~new_P1_U4437;
  assign new_P1_U3391 = ~new_P1_U3662 | ~new_P1_U3660 | ~new_P1_U4457 | ~new_P1_U4456;
  assign new_P1_U3392 = ~new_P1_U3666 | ~new_P1_U3664 | ~new_P1_U4476 | ~new_P1_U4475;
  assign new_P1_U3393 = ~new_P1_U3670 | ~new_P1_U3668 | ~new_P1_U4495 | ~new_P1_U4494;
  assign new_P1_U3394 = ~new_P1_U3674 | ~new_P1_U3672 | ~new_P1_U4514 | ~new_P1_U4513;
  assign new_P1_U3395 = ~new_P1_U3678 | ~new_P1_U3676 | ~new_P1_U4533 | ~new_P1_U4532;
  assign new_P1_U3396 = ~new_P1_U3682 | ~new_P1_U3680 | ~new_P1_U4552 | ~new_P1_U4551;
  assign new_P1_U3397 = ~new_U113 | ~new_P1_U3954;
  assign new_P1_U3398 = ~new_P1_U3686 | ~new_P1_U3684 | ~new_P1_U4571 | ~new_P1_U4570;
  assign new_P1_U3399 = ~new_U112 | ~new_P1_U3954;
  assign new_P1_U3400 = ~new_P1_U3690 | ~new_P1_U3688 | ~new_P1_U4590 | ~new_P1_U4589;
  assign new_P1_U3401 = ~new_U111 | ~new_P1_U3954;
  assign new_P1_U3402 = ~new_P1_U3694 | ~new_P1_U3692 | ~new_P1_U4609 | ~new_P1_U4608;
  assign new_P1_U3403 = ~new_U110 | ~new_P1_U3954;
  assign new_P1_U3404 = ~new_P1_U3698 | ~new_P1_U3696 | ~new_P1_U4628 | ~new_P1_U4627;
  assign new_P1_U3405 = ~new_U109 | ~new_P1_U3954;
  assign new_P1_U3406 = ~new_P1_U3702 | ~new_P1_U3700 | ~new_P1_U4647 | ~new_P1_U4646;
  assign new_P1_U3407 = ~new_U108 | ~new_P1_U3954;
  assign new_P1_U3408 = ~new_P1_U3706 | ~new_P1_U3704 | ~new_P1_U4666 | ~new_P1_U4665;
  assign new_P1_U3409 = ~new_U107 | ~new_P1_U3954;
  assign new_P1_U3410 = ~new_P1_U3710 | ~new_P1_U3708 | ~new_P1_U4685 | ~new_P1_U4684;
  assign new_P1_U3411 = ~new_U106 | ~new_P1_U3954;
  assign new_P1_U3412 = ~new_P1_U3714 | ~new_P1_U3712 | ~new_P1_U4704 | ~new_P1_U4703;
  assign new_P1_U3413 = ~new_U105 | ~new_P1_U3954;
  assign new_P1_U3414 = ~new_P1_U3718 | ~new_P1_U3716 | ~new_P1_U4723 | ~new_P1_U4722;
  assign new_P1_U3415 = ~new_U104 | ~new_P1_U3954;
  assign new_P1_U3416 = ~new_P1_U3723 | ~new_P1_U3721;
  assign new_P1_U3417 = ~new_U102 | ~new_P1_U3954;
  assign new_P1_U3418 = ~new_U101 | ~new_P1_U3954;
  assign new_P1_U3419 = ~new_P1_U4041 | ~new_P1_U5793;
  assign new_P1_U3420 = ~new_P1_U3022 | ~new_P1_U4767;
  assign new_P1_U3421 = ~new_P1_U3998 | ~new_P1_U5799;
  assign new_P1_U3422 = ~new_P1_U3048 | ~new_P1_U3450;
  assign new_P1_U3423 = ~new_P1_U3047 | ~new_P1_U5793;
  assign new_P1_U3424 = ~new_P1_U3993 | ~new_P1_U5799;
  assign new_P1_U3425 = ~new_P1_U3442 | ~new_P1_U3441 | ~new_P1_U3443;
  assign new_P1_U3426 = ~new_P1_U4010 | ~new_P1_U4768;
  assign new_P1_U3427 = ~new_P1_U3444 | ~P1_STATE_REG;
  assign new_P1_U3428 = ~new_P1_U3429 | ~new_P1_U4931;
  assign new_P1_U3429 = ~new_P1_U4145 | ~new_P1_U5786;
  assign new_P1_U3430 = ~new_P1_U4045 | ~P1_STATE_REG;
  assign new_P1_U3431 = ~new_P1_U3014 | ~new_P1_U3015;
  assign new_P1_U3432 = ~new_P1_R1375_U9;
  assign new_P1_U3433 = ~new_P1_U3022 | ~new_P1_U3426;
  assign new_P1_U3434 = ~new_P1_U3847 | ~new_P1_U3016;
  assign new_P1_U3435 = ~new_P1_U3852 | ~new_P1_U5143;
  assign new_P1_U3436 = ~new_P1_U5415 | ~new_P1_U5414;
  assign new_P1_U3437 = ~new_P1_U3999 | ~new_P1_U3362;
  assign new_P1_U3438 = ~new_P1_U5536 | ~new_P1_U3051;
  assign new_P1_U3439 = ~new_P1_R1352_U6;
  assign new_P1_U3440 = ~new_P1_U3364 | ~new_P1_U3423;
  assign new_P1_U3441 = ~new_P1_U5774 | ~new_P1_U5773;
  assign new_P1_U3442 = ~new_P1_U5777 | ~new_P1_U5776;
  assign new_P1_U3443 = ~new_P1_U5780 | ~new_P1_U5779;
  assign new_P1_U3444 = ~new_P1_U5785 | ~new_P1_U5784;
  assign n334 = ~new_P1_U5788 | ~new_P1_U5787;
  assign n339 = ~new_P1_U5790 | ~new_P1_U5789;
  assign new_P1_U3447 = ~new_P1_U5804 | ~new_P1_U5803;
  assign new_P1_U3448 = ~new_P1_U5807 | ~new_P1_U5806;
  assign new_P1_U3449 = ~new_P1_U5810 | ~new_P1_U5809;
  assign new_P1_U3450 = ~new_P1_U5801 | ~new_P1_U5800;
  assign new_P1_U3451 = ~new_P1_U5792 | ~new_P1_U5791;
  assign new_P1_U3452 = ~new_P1_U5795 | ~new_P1_U5794;
  assign new_P1_U3453 = ~new_P1_U5798 | ~new_P1_U5797;
  assign new_P1_U3454 = ~new_P1_U5813 | ~new_P1_U5812;
  assign new_P1_U3455 = ~new_P1_U5816 | ~new_P1_U5815;
  assign new_P1_U3456 = ~new_P1_U5819 | ~new_P1_U5818;
  assign new_P1_U3457 = ~new_P1_U5827 | ~new_P1_U5826;
  assign new_P1_U3458 = ~new_P1_U5824 | ~new_P1_U5823;
  assign n494 = ~new_P1_U5830 | ~new_P1_U5829;
  assign new_P1_U3460 = ~new_P1_U5832 | ~new_P1_U5831;
  assign new_P1_U3461 = ~new_P1_U5834 | ~new_P1_U5833;
  assign n499 = ~new_P1_U5837 | ~new_P1_U5836;
  assign new_P1_U3463 = ~new_P1_U5839 | ~new_P1_U5838;
  assign new_P1_U3464 = ~new_P1_U5841 | ~new_P1_U5840;
  assign n504 = ~new_P1_U5844 | ~new_P1_U5843;
  assign new_P1_U3466 = ~new_P1_U5846 | ~new_P1_U5845;
  assign new_P1_U3467 = ~new_P1_U5848 | ~new_P1_U5847;
  assign n509 = ~new_P1_U5851 | ~new_P1_U5850;
  assign new_P1_U3469 = ~new_P1_U5853 | ~new_P1_U5852;
  assign new_P1_U3470 = ~new_P1_U5855 | ~new_P1_U5854;
  assign n514 = ~new_P1_U5858 | ~new_P1_U5857;
  assign new_P1_U3472 = ~new_P1_U5860 | ~new_P1_U5859;
  assign new_P1_U3473 = ~new_P1_U5862 | ~new_P1_U5861;
  assign n519 = ~new_P1_U5865 | ~new_P1_U5864;
  assign new_P1_U3475 = ~new_P1_U5867 | ~new_P1_U5866;
  assign new_P1_U3476 = ~new_P1_U5869 | ~new_P1_U5868;
  assign n524 = ~new_P1_U5872 | ~new_P1_U5871;
  assign new_P1_U3478 = ~new_P1_U5874 | ~new_P1_U5873;
  assign new_P1_U3479 = ~new_P1_U5876 | ~new_P1_U5875;
  assign n529 = ~new_P1_U5879 | ~new_P1_U5878;
  assign new_P1_U3481 = ~new_P1_U5881 | ~new_P1_U5880;
  assign new_P1_U3482 = ~new_P1_U5883 | ~new_P1_U5882;
  assign n534 = ~new_P1_U5886 | ~new_P1_U5885;
  assign new_P1_U3484 = ~new_P1_U5888 | ~new_P1_U5887;
  assign new_P1_U3485 = ~new_P1_U5890 | ~new_P1_U5889;
  assign n539 = ~new_P1_U5893 | ~new_P1_U5892;
  assign new_P1_U3487 = ~new_P1_U5895 | ~new_P1_U5894;
  assign new_P1_U3488 = ~new_P1_U5897 | ~new_P1_U5896;
  assign n544 = ~new_P1_U5900 | ~new_P1_U5899;
  assign new_P1_U3490 = ~new_P1_U5902 | ~new_P1_U5901;
  assign new_P1_U3491 = ~new_P1_U5904 | ~new_P1_U5903;
  assign n549 = ~new_P1_U5907 | ~new_P1_U5906;
  assign new_P1_U3493 = ~new_P1_U5909 | ~new_P1_U5908;
  assign new_P1_U3494 = ~new_P1_U5911 | ~new_P1_U5910;
  assign n554 = ~new_P1_U5914 | ~new_P1_U5913;
  assign new_P1_U3496 = ~new_P1_U5916 | ~new_P1_U5915;
  assign new_P1_U3497 = ~new_P1_U5918 | ~new_P1_U5917;
  assign n559 = ~new_P1_U5921 | ~new_P1_U5920;
  assign new_P1_U3499 = ~new_P1_U5923 | ~new_P1_U5922;
  assign new_P1_U3500 = ~new_P1_U5925 | ~new_P1_U5924;
  assign n564 = ~new_P1_U5928 | ~new_P1_U5927;
  assign new_P1_U3502 = ~new_P1_U5930 | ~new_P1_U5929;
  assign new_P1_U3503 = ~new_P1_U5932 | ~new_P1_U5931;
  assign n569 = ~new_P1_U5935 | ~new_P1_U5934;
  assign new_P1_U3505 = ~new_P1_U5937 | ~new_P1_U5936;
  assign new_P1_U3506 = ~new_P1_U5939 | ~new_P1_U5938;
  assign n574 = ~new_P1_U5942 | ~new_P1_U5941;
  assign new_P1_U3508 = ~new_P1_U5944 | ~new_P1_U5943;
  assign new_P1_U3509 = ~new_P1_U5946 | ~new_P1_U5945;
  assign n579 = ~new_P1_U5949 | ~new_P1_U5948;
  assign new_P1_U3511 = ~new_P1_U5951 | ~new_P1_U5950;
  assign new_P1_U3512 = ~new_P1_U5953 | ~new_P1_U5952;
  assign n584 = ~new_P1_U5956 | ~new_P1_U5955;
  assign new_P1_U3514 = ~new_P1_U5958 | ~new_P1_U5957;
  assign n589 = ~new_P1_U5961 | ~new_P1_U5960;
  assign n594 = ~new_P1_U5963 | ~new_P1_U5962;
  assign n599 = ~new_P1_U5965 | ~new_P1_U5964;
  assign n604 = ~new_P1_U5967 | ~new_P1_U5966;
  assign n609 = ~new_P1_U5969 | ~new_P1_U5968;
  assign n614 = ~new_P1_U5971 | ~new_P1_U5970;
  assign n619 = ~new_P1_U5973 | ~new_P1_U5972;
  assign n624 = ~new_P1_U5975 | ~new_P1_U5974;
  assign n629 = ~new_P1_U5977 | ~new_P1_U5976;
  assign n634 = ~new_P1_U5979 | ~new_P1_U5978;
  assign n639 = ~new_P1_U5981 | ~new_P1_U5980;
  assign n644 = ~new_P1_U5983 | ~new_P1_U5982;
  assign n649 = ~new_P1_U5985 | ~new_P1_U5984;
  assign n654 = ~new_P1_U5987 | ~new_P1_U5986;
  assign n659 = ~new_P1_U5989 | ~new_P1_U5988;
  assign n664 = ~new_P1_U5991 | ~new_P1_U5990;
  assign n669 = ~new_P1_U5993 | ~new_P1_U5992;
  assign n674 = ~new_P1_U5995 | ~new_P1_U5994;
  assign n679 = ~new_P1_U5997 | ~new_P1_U5996;
  assign n684 = ~new_P1_U5999 | ~new_P1_U5998;
  assign n689 = ~new_P1_U6001 | ~new_P1_U6000;
  assign n694 = ~new_P1_U6003 | ~new_P1_U6002;
  assign n699 = ~new_P1_U6005 | ~new_P1_U6004;
  assign n704 = ~new_P1_U6007 | ~new_P1_U6006;
  assign n709 = ~new_P1_U6009 | ~new_P1_U6008;
  assign n714 = ~new_P1_U6011 | ~new_P1_U6010;
  assign n719 = ~new_P1_U6013 | ~new_P1_U6012;
  assign n724 = ~new_P1_U6015 | ~new_P1_U6014;
  assign n729 = ~new_P1_U6017 | ~new_P1_U6016;
  assign n734 = ~new_P1_U6019 | ~new_P1_U6018;
  assign n739 = ~new_P1_U6021 | ~new_P1_U6020;
  assign n744 = ~new_P1_U6023 | ~new_P1_U6022;
  assign n749 = ~new_P1_U6025 | ~new_P1_U6024;
  assign n754 = ~new_P1_U6027 | ~new_P1_U6026;
  assign n759 = ~new_P1_U6029 | ~new_P1_U6028;
  assign n764 = ~new_P1_U6031 | ~new_P1_U6030;
  assign n769 = ~new_P1_U6033 | ~new_P1_U6032;
  assign n774 = ~new_P1_U6035 | ~new_P1_U6034;
  assign n779 = ~new_P1_U6037 | ~new_P1_U6036;
  assign n784 = ~new_P1_U6039 | ~new_P1_U6038;
  assign n789 = ~new_P1_U6041 | ~new_P1_U6040;
  assign n794 = ~new_P1_U6043 | ~new_P1_U6042;
  assign n799 = ~new_P1_U6045 | ~new_P1_U6044;
  assign n804 = ~new_P1_U6047 | ~new_P1_U6046;
  assign n809 = ~new_P1_U6049 | ~new_P1_U6048;
  assign n1074 = ~new_P1_U6115 | ~new_P1_U6114;
  assign n1079 = ~new_P1_U6117 | ~new_P1_U6116;
  assign n1084 = ~new_P1_U6119 | ~new_P1_U6118;
  assign n1089 = ~new_P1_U6121 | ~new_P1_U6120;
  assign n1094 = ~new_P1_U6123 | ~new_P1_U6122;
  assign n1099 = ~new_P1_U6125 | ~new_P1_U6124;
  assign n1104 = ~new_P1_U6127 | ~new_P1_U6126;
  assign n1109 = ~new_P1_U6129 | ~new_P1_U6128;
  assign n1114 = ~new_P1_U6131 | ~new_P1_U6130;
  assign n1119 = ~new_P1_U6133 | ~new_P1_U6132;
  assign n1124 = ~new_P1_U6135 | ~new_P1_U6134;
  assign n1129 = ~new_P1_U6137 | ~new_P1_U6136;
  assign n1134 = ~new_P1_U6139 | ~new_P1_U6138;
  assign n1139 = ~new_P1_U6141 | ~new_P1_U6140;
  assign n1144 = ~new_P1_U6143 | ~new_P1_U6142;
  assign n1149 = ~new_P1_U6145 | ~new_P1_U6144;
  assign n1154 = ~new_P1_U6147 | ~new_P1_U6146;
  assign n1159 = ~new_P1_U6149 | ~new_P1_U6148;
  assign n1164 = ~new_P1_U6151 | ~new_P1_U6150;
  assign n1169 = ~new_P1_U6153 | ~new_P1_U6152;
  assign n1174 = ~new_P1_U6155 | ~new_P1_U6154;
  assign n1179 = ~new_P1_U6157 | ~new_P1_U6156;
  assign n1184 = ~new_P1_U6159 | ~new_P1_U6158;
  assign n1189 = ~new_P1_U6161 | ~new_P1_U6160;
  assign n1194 = ~new_P1_U6163 | ~new_P1_U6162;
  assign n1199 = ~new_P1_U6165 | ~new_P1_U6164;
  assign n1204 = ~new_P1_U6167 | ~new_P1_U6166;
  assign n1209 = ~new_P1_U6169 | ~new_P1_U6168;
  assign n1214 = ~new_P1_U6171 | ~new_P1_U6170;
  assign n1219 = ~new_P1_U6173 | ~new_P1_U6172;
  assign n1224 = ~new_P1_U6175 | ~new_P1_U6174;
  assign n1229 = ~new_P1_U6177 | ~new_P1_U6176;
  assign new_P1_U3592 = new_P1_U5786 & P1_STATE_REG;
  assign new_P1_U3593 = new_P1_U4187 & new_P1_U4186;
  assign new_P1_U3594 = new_P1_U4189 & new_P1_U4188;
  assign new_P1_U3595 = new_P1_U4195 & new_P1_U4196;
  assign new_P1_U3596 = new_P1_U4148 & new_P1_U4149 & new_P1_U4151 & new_P1_U4150;
  assign new_P1_U3597 = new_P1_U4152 & new_P1_U4153 & new_P1_U4155 & new_P1_U4154;
  assign new_P1_U3598 = new_P1_U4156 & new_P1_U4157 & new_P1_U4159 & new_P1_U4158;
  assign new_P1_U3599 = new_P1_U4162 & new_P1_U4161 & new_P1_U4160;
  assign new_P1_U3600 = new_P1_U3596 & new_P1_U3597 & new_P1_U3599 & new_P1_U3598;
  assign new_P1_U3601 = new_P1_U4163 & new_P1_U4164 & new_P1_U4166 & new_P1_U4165;
  assign new_P1_U3602 = new_P1_U4167 & new_P1_U4168 & new_P1_U4170 & new_P1_U4169;
  assign new_P1_U3603 = new_P1_U4171 & new_P1_U4172 & new_P1_U4174 & new_P1_U4173;
  assign new_P1_U3604 = new_P1_U4177 & new_P1_U4176 & new_P1_U4175;
  assign new_P1_U3605 = new_P1_U3601 & new_P1_U3602 & new_P1_U3604 & new_P1_U3603;
  assign new_P1_U3606 = new_P1_U5825 & new_P1_U4179;
  assign new_P1_U3607 = new_P1_U5828 & new_P1_U3022;
  assign new_P1_U3608 = new_P1_U4212 & new_P1_U4211;
  assign new_P1_U3609 = new_P1_U4214 & new_P1_U4213;
  assign new_P1_U3610 = new_P1_U3609 & new_P1_U4216 & new_P1_U4215;
  assign new_P1_U3611 = new_P1_U4219 & new_P1_U4221 & new_P1_U4220 & new_P1_U4218;
  assign new_P1_U3612 = new_P1_U4231 & new_P1_U4230;
  assign new_P1_U3613 = new_P1_U4233 & new_P1_U4232;
  assign new_P1_U3614 = new_P1_U3613 & new_P1_U4235 & new_P1_U4234;
  assign new_P1_U3615 = new_P1_U4238 & new_P1_U4240 & new_P1_U4239 & new_P1_U4237;
  assign new_P1_U3616 = new_P1_U4250 & new_P1_U4249;
  assign new_P1_U3617 = new_P1_U4252 & new_P1_U4251;
  assign new_P1_U3618 = new_P1_U3617 & new_P1_U4254 & new_P1_U4253;
  assign new_P1_U3619 = new_P1_U4257 & new_P1_U4259 & new_P1_U4258 & new_P1_U4256;
  assign new_P1_U3620 = new_P1_U4269 & new_P1_U4268;
  assign new_P1_U3621 = new_P1_U4271 & new_P1_U4270;
  assign new_P1_U3622 = new_P1_U3621 & new_P1_U4273 & new_P1_U4272;
  assign new_P1_U3623 = new_P1_U4276 & new_P1_U4278 & new_P1_U4277 & new_P1_U4275;
  assign new_P1_U3624 = new_P1_U4288 & new_P1_U4287;
  assign new_P1_U3625 = new_P1_U4290 & new_P1_U4289;
  assign new_P1_U3626 = new_P1_U3625 & new_P1_U4292 & new_P1_U4291;
  assign new_P1_U3627 = new_P1_U4295 & new_P1_U4297 & new_P1_U4296 & new_P1_U4294;
  assign new_P1_U3628 = new_P1_U4307 & new_P1_U4306;
  assign new_P1_U3629 = new_P1_U4309 & new_P1_U4308;
  assign new_P1_U3630 = new_P1_U3629 & new_P1_U4311 & new_P1_U4310;
  assign new_P1_U3631 = new_P1_U4314 & new_P1_U4316 & new_P1_U4315 & new_P1_U4313;
  assign new_P1_U3632 = new_P1_U4326 & new_P1_U4325;
  assign new_P1_U3633 = new_P1_U4328 & new_P1_U4327;
  assign new_P1_U3634 = new_P1_U3633 & new_P1_U4330 & new_P1_U4329;
  assign new_P1_U3635 = new_P1_U4333 & new_P1_U4335 & new_P1_U4334 & new_P1_U4332;
  assign new_P1_U3636 = new_P1_U4345 & new_P1_U4344;
  assign new_P1_U3637 = new_P1_U4347 & new_P1_U4346;
  assign new_P1_U3638 = new_P1_U3637 & new_P1_U4349 & new_P1_U4348;
  assign new_P1_U3639 = new_P1_U4352 & new_P1_U4354 & new_P1_U4353 & new_P1_U4351;
  assign new_P1_U3640 = new_P1_U4364 & new_P1_U4363;
  assign new_P1_U3641 = new_P1_U4366 & new_P1_U4365;
  assign new_P1_U3642 = new_P1_U3641 & new_P1_U4368 & new_P1_U4367;
  assign new_P1_U3643 = new_P1_U4371 & new_P1_U4373 & new_P1_U4372 & new_P1_U4370;
  assign new_P1_U3644 = new_P1_U4383 & new_P1_U4382;
  assign new_P1_U3645 = new_P1_U4385 & new_P1_U4384;
  assign new_P1_U3646 = new_P1_U3645 & new_P1_U4387 & new_P1_U4386;
  assign new_P1_U3647 = new_P1_U4390 & new_P1_U4392 & new_P1_U4391 & new_P1_U4389;
  assign new_P1_U3648 = new_P1_U4402 & new_P1_U4401;
  assign new_P1_U3649 = new_P1_U4404 & new_P1_U4403;
  assign new_P1_U3650 = new_P1_U3649 & new_P1_U4406 & new_P1_U4405;
  assign new_P1_U3651 = new_P1_U4408 & new_P1_U4409 & new_P1_U4411 & new_P1_U4410;
  assign new_P1_U3652 = new_P1_U4421 & new_P1_U4420;
  assign new_P1_U3653 = new_P1_U4423 & new_P1_U4422;
  assign new_P1_U3654 = new_P1_U3653 & new_P1_U4425 & new_P1_U4424;
  assign new_P1_U3655 = new_P1_U4427 & new_P1_U4429 & new_P1_U4430 & new_P1_U4428;
  assign new_P1_U3656 = new_P1_U4440 & new_P1_U4439;
  assign new_P1_U3657 = new_P1_U4442 & new_P1_U4441;
  assign new_P1_U3658 = new_P1_U3657 & new_P1_U4444 & new_P1_U4443;
  assign new_P1_U3659 = new_P1_U4446 & new_P1_U4447 & new_P1_U4449 & new_P1_U4448;
  assign new_P1_U3660 = new_P1_U4459 & new_P1_U4458;
  assign new_P1_U3661 = new_P1_U4461 & new_P1_U4460;
  assign new_P1_U3662 = new_P1_U3661 & new_P1_U4463 & new_P1_U4462;
  assign new_P1_U3663 = new_P1_U4465 & new_P1_U4467 & new_P1_U4468 & new_P1_U4466;
  assign new_P1_U3664 = new_P1_U4478 & new_P1_U4477;
  assign new_P1_U3665 = new_P1_U4480 & new_P1_U4479;
  assign new_P1_U3666 = new_P1_U3665 & new_P1_U4482 & new_P1_U4481;
  assign new_P1_U3667 = new_P1_U4485 & new_P1_U4487 & new_P1_U4486 & new_P1_U4484;
  assign new_P1_U3668 = new_P1_U4497 & new_P1_U4496;
  assign new_P1_U3669 = new_P1_U4499 & new_P1_U4498;
  assign new_P1_U3670 = new_P1_U3669 & new_P1_U4501 & new_P1_U4500;
  assign new_P1_U3671 = new_P1_U4504 & new_P1_U4506 & new_P1_U4505 & new_P1_U4503;
  assign new_P1_U3672 = new_P1_U4516 & new_P1_U4515;
  assign new_P1_U3673 = new_P1_U4518 & new_P1_U4517;
  assign new_P1_U3674 = new_P1_U3673 & new_P1_U4520 & new_P1_U4519;
  assign new_P1_U3675 = new_P1_U4522 & new_P1_U4524 & new_P1_U4525 & new_P1_U4523;
  assign new_P1_U3676 = new_P1_U4535 & new_P1_U4534;
  assign new_P1_U3677 = new_P1_U4537 & new_P1_U4536;
  assign new_P1_U3678 = new_P1_U3677 & new_P1_U4539 & new_P1_U4538;
  assign new_P1_U3679 = new_P1_U4541 & new_P1_U4543 & new_P1_U4544 & new_P1_U4542;
  assign new_P1_U3680 = new_P1_U4554 & new_P1_U4553;
  assign new_P1_U3681 = new_P1_U4556 & new_P1_U4555;
  assign new_P1_U3682 = new_P1_U3681 & new_P1_U4558 & new_P1_U4557;
  assign new_P1_U3683 = new_P1_U4561 & new_P1_U4563 & new_P1_U4562 & new_P1_U4560;
  assign new_P1_U3684 = new_P1_U4573 & new_P1_U4572;
  assign new_P1_U3685 = new_P1_U4575 & new_P1_U4574;
  assign new_P1_U3686 = new_P1_U3685 & new_P1_U4577 & new_P1_U4576;
  assign new_P1_U3687 = new_P1_U4580 & new_P1_U4582 & new_P1_U4581 & new_P1_U4579;
  assign new_P1_U3688 = new_P1_U4592 & new_P1_U4591;
  assign new_P1_U3689 = new_P1_U4594 & new_P1_U4593;
  assign new_P1_U3690 = new_P1_U3689 & new_P1_U4596 & new_P1_U4595;
  assign new_P1_U3691 = new_P1_U4599 & new_P1_U4601 & new_P1_U4600 & new_P1_U4598;
  assign new_P1_U3692 = new_P1_U4611 & new_P1_U4610;
  assign new_P1_U3693 = new_P1_U4613 & new_P1_U4612;
  assign new_P1_U3694 = new_P1_U3693 & new_P1_U4615 & new_P1_U4614;
  assign new_P1_U3695 = new_P1_U4618 & new_P1_U4620 & new_P1_U4619 & new_P1_U4617;
  assign new_P1_U3696 = new_P1_U4630 & new_P1_U4629;
  assign new_P1_U3697 = new_P1_U4632 & new_P1_U4631;
  assign new_P1_U3698 = new_P1_U3697 & new_P1_U4634 & new_P1_U4633;
  assign new_P1_U3699 = new_P1_U4637 & new_P1_U4639 & new_P1_U4638 & new_P1_U4636;
  assign new_P1_U3700 = new_P1_U4649 & new_P1_U4648;
  assign new_P1_U3701 = new_P1_U4651 & new_P1_U4650;
  assign new_P1_U3702 = new_P1_U3701 & new_P1_U4653 & new_P1_U4652;
  assign new_P1_U3703 = new_P1_U4656 & new_P1_U4658 & new_P1_U4657 & new_P1_U4655;
  assign new_P1_U3704 = new_P1_U4668 & new_P1_U4667;
  assign new_P1_U3705 = new_P1_U4670 & new_P1_U4669;
  assign new_P1_U3706 = new_P1_U3705 & new_P1_U4672 & new_P1_U4671;
  assign new_P1_U3707 = new_P1_U4675 & new_P1_U4677 & new_P1_U4676 & new_P1_U4674;
  assign new_P1_U3708 = new_P1_U4687 & new_P1_U4686;
  assign new_P1_U3709 = new_P1_U4689 & new_P1_U4688;
  assign new_P1_U3710 = new_P1_U3709 & new_P1_U4691 & new_P1_U4690;
  assign new_P1_U3711 = new_P1_U4694 & new_P1_U4696 & new_P1_U4695 & new_P1_U4693;
  assign new_P1_U3712 = new_P1_U4706 & new_P1_U4705;
  assign new_P1_U3713 = new_P1_U4708 & new_P1_U4707;
  assign new_P1_U3714 = new_P1_U3713 & new_P1_U4710 & new_P1_U4709;
  assign new_P1_U3715 = new_P1_U4713 & new_P1_U4715 & new_P1_U4714 & new_P1_U4712;
  assign new_P1_U3716 = new_P1_U4725 & new_P1_U4724;
  assign new_P1_U3717 = new_P1_U4727 & new_P1_U4726;
  assign new_P1_U3718 = new_P1_U3717 & new_P1_U4729 & new_P1_U4728;
  assign new_P1_U3719 = new_P1_U4732 & new_P1_U4734 & new_P1_U4733 & new_P1_U4731;
  assign new_P1_U3720 = new_P1_U4741 & new_P1_U4030;
  assign new_P1_U3721 = new_P1_U4746 & new_P1_U4745 & new_P1_U4744 & new_P1_U4743 & new_P1_U4742;
  assign new_P1_U3722 = new_P1_U4748 & new_P1_U4747;
  assign new_P1_U3723 = new_P1_U3722 & new_P1_U4750 & new_P1_U4749;
  assign new_P1_U3724 = new_P1_U4752 & new_P1_U4753 & new_P1_U4754;
  assign new_P1_U3725 = new_P1_U4030 & new_P1_U4741;
  assign new_P1_U3726 = new_P1_U3022 & new_P1_U3457;
  assign new_P1_U3727 = new_P1_U3458 & new_P1_U5828 & new_P1_U4012;
  assign new_P1_U3728 = new_P1_U4772 & new_P1_U4771 & new_P1_U4770;
  assign new_P1_U3729 = new_P1_U3957 & new_P1_U4774 & new_P1_U4773;
  assign new_P1_U3730 = new_P1_U4777 & new_P1_U4776 & new_P1_U4775;
  assign new_P1_U3731 = new_P1_U3958 & new_P1_U4779 & new_P1_U4778;
  assign new_P1_U3732 = new_P1_U4782 & new_P1_U4781 & new_P1_U4780;
  assign new_P1_U3733 = new_P1_U3959 & new_P1_U4784 & new_P1_U4783;
  assign new_P1_U3734 = new_P1_U4787 & new_P1_U4786 & new_P1_U4785;
  assign new_P1_U3735 = new_P1_U3960 & new_P1_U4789 & new_P1_U4788;
  assign new_P1_U3736 = new_P1_U4792 & new_P1_U4791 & new_P1_U4790;
  assign new_P1_U3737 = new_P1_U3961 & new_P1_U4794 & new_P1_U4793;
  assign new_P1_U3738 = new_P1_U4797 & new_P1_U4796 & new_P1_U4795;
  assign new_P1_U3739 = new_P1_U4799 & new_P1_U4798;
  assign new_P1_U3740 = new_P1_U4802 & new_P1_U4801 & new_P1_U4800;
  assign new_P1_U3741 = new_P1_U4804 & new_P1_U4803;
  assign new_P1_U3742 = new_P1_U4807 & new_P1_U4806 & new_P1_U4805;
  assign new_P1_U3743 = new_P1_U4809 & new_P1_U4808;
  assign new_P1_U3744 = new_P1_U4812 & new_P1_U4811 & new_P1_U4810;
  assign new_P1_U3745 = new_P1_U4814 & new_P1_U4813;
  assign new_P1_U3746 = new_P1_U4816 & new_P1_U4815;
  assign new_P1_U3747 = new_P1_U4819 & new_P1_U4818;
  assign new_P1_U3748 = new_P1_U4821 & new_P1_U4820;
  assign new_P1_U3749 = new_P1_U4824 & new_P1_U4823;
  assign new_P1_U3750 = new_P1_U4827 & new_P1_U4826 & new_P1_U4825;
  assign new_P1_U3751 = new_P1_U4829 & new_P1_U4828;
  assign new_P1_U3752 = new_P1_U4832 & new_P1_U4831 & new_P1_U4830;
  assign new_P1_U3753 = new_P1_U4834 & new_P1_U4833;
  assign new_P1_U3754 = new_P1_U4837 & new_P1_U4836 & new_P1_U4835;
  assign new_P1_U3755 = new_P1_U4839 & new_P1_U4838;
  assign new_P1_U3756 = new_P1_U4842 & new_P1_U4841 & new_P1_U4840;
  assign new_P1_U3757 = new_P1_U4844 & new_P1_U4843;
  assign new_P1_U3758 = new_P1_U4846 & new_P1_U4845;
  assign new_P1_U3759 = new_P1_U4849 & new_P1_U4848;
  assign new_P1_U3760 = new_P1_U4851 & new_P1_U4850;
  assign new_P1_U3761 = new_P1_U4854 & new_P1_U4853;
  assign new_P1_U3762 = new_P1_U4857 & new_P1_U4856 & new_P1_U4855;
  assign new_P1_U3763 = new_P1_U4859 & new_P1_U4858;
  assign new_P1_U3764 = new_P1_U4862 & new_P1_U4861 & new_P1_U4860;
  assign new_P1_U3765 = new_P1_U4864 & new_P1_U4863;
  assign new_P1_U3766 = new_P1_U4866 & new_P1_U4865;
  assign new_P1_U3767 = new_P1_U4869 & new_P1_U4868;
  assign new_P1_U3768 = new_P1_U4871 & new_P1_U4870;
  assign new_P1_U3769 = new_P1_U4874 & new_P1_U4873;
  assign new_P1_U3770 = new_P1_U4876 & new_P1_U4875;
  assign new_P1_U3771 = new_P1_U4879 & new_P1_U4878;
  assign new_P1_U3772 = new_P1_U4881 & new_P1_U4880;
  assign new_P1_U3773 = new_P1_U4884 & new_P1_U4883;
  assign new_P1_U3774 = new_P1_U4886 & new_P1_U4885;
  assign new_P1_U3775 = new_P1_U4889 & new_P1_U4888;
  assign new_P1_U3776 = new_P1_U4891 & new_P1_U4890;
  assign new_P1_U3777 = new_P1_U4894 & new_P1_U4893;
  assign new_P1_U3778 = new_P1_U4896 & new_P1_U4895;
  assign new_P1_U3779 = new_P1_U4899 & new_P1_U4898;
  assign new_P1_U3780 = new_P1_U4901 & new_P1_U4900;
  assign new_P1_U3781 = new_P1_U4904 & new_P1_U4903;
  assign new_P1_U3782 = new_P1_U4906 & new_P1_U4905;
  assign new_P1_U3783 = new_P1_U4909 & new_P1_U4908;
  assign new_P1_U3784 = new_P1_U4911 & new_P1_U4910;
  assign new_P1_U3785 = new_P1_U4914 & new_P1_U4913;
  assign new_P1_U3786 = new_P1_U3370 & new_P1_U3362 & new_P1_U3364;
  assign new_P1_U3787 = new_P1_U3365 & new_P1_U3366 & new_P1_U3422;
  assign new_P1_U3788 = new_P1_U3361 & new_P1_U4006;
  assign new_P1_U3789 = new_P1_U3788 & new_P1_U3424;
  assign new_P1_U3790 = new_P1_U4934 & new_P1_U4935;
  assign new_P1_U3791 = new_P1_U4937 & new_P1_U4938 & new_P1_U4936;
  assign new_P1_U3792 = new_P1_U4944 & new_P1_U4945;
  assign new_P1_U3793 = new_P1_U4947 & new_P1_U4948 & new_P1_U4946;
  assign new_P1_U3794 = new_P1_U4954 & new_P1_U4955;
  assign new_P1_U3795 = new_P1_U4957 & new_P1_U4958 & new_P1_U4956;
  assign new_P1_U3796 = new_P1_U4964 & new_P1_U4965;
  assign new_P1_U3797 = new_P1_U4967 & new_P1_U4968 & new_P1_U4966;
  assign new_P1_U3798 = new_P1_U4974 & new_P1_U4975;
  assign new_P1_U3799 = new_P1_U4977 & new_P1_U4978 & new_P1_U4976;
  assign new_P1_U3800 = new_P1_U4984 & new_P1_U4985;
  assign new_P1_U3801 = new_P1_U4987 & new_P1_U4988 & new_P1_U4986;
  assign new_P1_U3802 = new_P1_U4994 & new_P1_U4995;
  assign new_P1_U3803 = new_P1_U4997 & new_P1_U4998 & new_P1_U4996;
  assign new_P1_U3804 = new_P1_U5004 & new_P1_U5005;
  assign new_P1_U3805 = new_P1_U5007 & new_P1_U5008 & new_P1_U5006;
  assign new_P1_U3806 = new_P1_U5014 & new_P1_U5015;
  assign new_P1_U3807 = new_P1_U5017 & new_P1_U5018 & new_P1_U5016;
  assign new_P1_U3808 = new_P1_U5024 & new_P1_U5025;
  assign new_P1_U3809 = new_P1_U5027 & new_P1_U5028 & new_P1_U5026;
  assign new_P1_U3810 = new_P1_U5034 & new_P1_U5035;
  assign new_P1_U3811 = new_P1_U5037 & new_P1_U5038 & new_P1_U5036;
  assign new_P1_U3812 = new_P1_U5044 & new_P1_U5045;
  assign new_P1_U3813 = new_P1_U5047 & new_P1_U5048 & new_P1_U5046;
  assign new_P1_U3814 = new_P1_U5054 & new_P1_U5055;
  assign new_P1_U3815 = new_P1_U5057 & new_P1_U5058 & new_P1_U5056;
  assign new_P1_U3816 = new_P1_U5064 & new_P1_U5065;
  assign new_P1_U3817 = new_P1_U5068 & new_P1_U5067 & new_P1_U5066;
  assign new_P1_U3818 = new_P1_U5074 & new_P1_U5075;
  assign new_P1_U3819 = new_P1_U5078 & new_P1_U5077 & new_P1_U5076;
  assign new_P1_U3820 = new_P1_U3821 & new_P1_U5084;
  assign new_P1_U3821 = new_P1_U5085 & new_P1_U4040;
  assign new_P1_U3822 = new_P1_U5088 & new_P1_U5087 & new_P1_U5086;
  assign new_P1_U3823 = new_P1_U5094 & new_P1_U5095;
  assign new_P1_U3824 = new_P1_U5098 & new_P1_U5097 & new_P1_U5096;
  assign new_P1_U3825 = new_P1_U3826 & new_P1_U5104;
  assign new_P1_U3826 = new_P1_U5105 & new_P1_U4040;
  assign new_P1_U3827 = new_P1_U5108 & new_P1_U5107 & new_P1_U5106;
  assign new_P1_U3828 = new_P1_U5114 & new_P1_U5115;
  assign new_P1_U3829 = new_P1_U5118 & new_P1_U5117 & new_P1_U5116;
  assign new_P1_U3830 = new_P1_U5124 & new_P1_U5125;
  assign new_P1_U3831 = new_P1_U5128 & new_P1_U5127 & new_P1_U5126;
  assign new_P1_U3832 = new_P1_U6221 & new_P1_U6218 & new_P1_U6215;
  assign new_P1_U3833 = new_P1_U6233 & new_P1_U3834 & new_P1_U3832;
  assign new_P1_U3834 = new_P1_U6224 & new_P1_U6230 & new_P1_U6227;
  assign new_P1_U3835 = new_P1_U6245 & new_P1_U6242 & new_P1_U6239;
  assign new_P1_U3836 = new_P1_U6254 & new_P1_U6251 & new_P1_U6248;
  assign new_P1_U3837 = new_P1_U6236 & new_P1_U3836 & new_P1_U3835;
  assign new_P1_U3838 = new_P1_U6191 & new_P1_U6188 & new_P1_U6185;
  assign new_P1_U3839 = new_P1_U6206 & new_P1_U6194 & new_P1_U6197 & new_P1_U6203 & new_P1_U6200;
  assign new_P1_U3840 = new_P1_U6260 & new_P1_U6263 & new_P1_U6269 & new_P1_U6266;
  assign new_P1_U3841 = new_P1_U6275 & new_P1_U6272;
  assign new_P1_U3842 = new_P1_U3841 & new_P1_U3840;
  assign new_P1_U3843 = new_P1_U6209 & new_P1_U6257 & new_P1_U6212 & new_P1_U3837 & new_P1_U3833;
  assign new_P1_U3844 = new_P1_U6182 & new_P1_U3839 & new_P1_U3838;
  assign new_P1_U3845 = new_P1_U3429 & P1_STATE_REG;
  assign new_P1_U3846 = new_P1_U5138 & new_P1_U5136;
  assign new_P1_U3847 = new_P1_U3457 & new_P1_U3458;
  assign new_P1_U3848 = new_P1_U3996 & new_P1_U3997 & new_P1_U3371;
  assign new_P1_U3849 = new_P1_U3368 & new_P1_U3424;
  assign new_P1_U3850 = new_P1_U3427 & new_P1_U3430;
  assign new_P1_U3851 = new_P1_U3022 & new_P1_U5145;
  assign new_P1_U3852 = new_P1_U3425 & P1_STATE_REG;
  assign new_P1_U3853 = new_P1_U5173 & new_P1_U5172;
  assign new_P1_U3854 = new_P1_U5189 & new_P1_U5187;
  assign new_P1_U3855 = new_P1_U5191 & new_P1_U5190;
  assign new_P1_U3856 = new_P1_U5200 & new_P1_U5199;
  assign new_P1_U3857 = new_P1_U5218 & new_P1_U5217;
  assign new_P1_U3858 = new_P1_U4037 & new_P1_U3078;
  assign new_P1_U3859 = new_P1_U3860 & new_P1_U5232 & new_P1_U5231;
  assign new_P1_U3860 = new_P1_U5235 & new_P1_U5234;
  assign new_P1_U3861 = new_P1_U5244 & new_P1_U5243;
  assign new_P1_U3862 = new_P1_U5251 & new_P1_U5249;
  assign new_P1_U3863 = new_P1_U5253 & new_P1_U5252;
  assign new_P1_U3864 = new_P1_U5280 & new_P1_U5279;
  assign new_P1_U3865 = new_P1_U5307 & new_P1_U5306;
  assign new_P1_U3866 = new_P1_U5323 & new_P1_U5321;
  assign new_P1_U3867 = new_P1_U5325 & new_P1_U5324;
  assign new_P1_U3868 = new_P1_U5334 & new_P1_U5333;
  assign new_P1_U3869 = new_P1_U5359 & new_P1_U5357;
  assign new_P1_U3870 = new_P1_U5361 & new_P1_U5360;
  assign new_P1_U3871 = new_P1_U5370 & new_P1_U5369;
  assign new_P1_U3872 = new_P1_U5406 & new_P1_U5405;
  assign new_P1_U3873 = new_P1_U5802 & new_P1_U5793;
  assign new_P1_U3874 = new_P1_U3375 & new_P1_U5410;
  assign new_P1_U3875 = new_P1_U5475 & new_P1_U5476;
  assign new_P1_U3876 = new_P1_U5535 & new_P1_U5533;
  assign new_P1_U3877 = new_P1_U3444 & new_P1_U5538;
  assign new_P1_U3878 = new_P1_U3374 & new_P1_U3997;
  assign new_P1_U3879 = new_P1_U3878 & new_P1_U3371;
  assign new_P1_U3880 = new_P1_U3881 & new_P1_U5546;
  assign new_P1_U3881 = new_P1_U3444 & new_P1_U5544;
  assign new_P1_U3882 = new_P1_U3883 & new_P1_U5549;
  assign new_P1_U3883 = new_P1_U3444 & new_P1_U5547;
  assign new_P1_U3884 = new_P1_U3885 & new_P1_U5552;
  assign new_P1_U3885 = new_P1_U3444 & new_P1_U5550;
  assign new_P1_U3886 = new_P1_U3887 & new_P1_U5555;
  assign new_P1_U3887 = new_P1_U3444 & new_P1_U5553;
  assign new_P1_U3888 = new_P1_U3889 & new_P1_U5558;
  assign new_P1_U3889 = new_P1_U3444 & new_P1_U5556;
  assign new_P1_U3890 = new_P1_U3891 & new_P1_U5561;
  assign new_P1_U3891 = new_P1_U3444 & new_P1_U5559;
  assign new_P1_U3892 = new_P1_U5564 & new_P1_U5562;
  assign new_P1_U3893 = new_P1_U5567 & new_P1_U5565;
  assign new_P1_U3894 = new_P1_U3895 & new_P1_U5570;
  assign new_P1_U3895 = new_P1_U3444 & new_P1_U5568;
  assign new_P1_U3896 = new_P1_U3444 & new_P1_U5573;
  assign new_P1_U3897 = new_P1_U3444 & new_P1_U5576;
  assign new_P1_U3898 = new_P1_U3444 & new_P1_U5579;
  assign new_P1_U3899 = new_P1_U3444 & new_P1_U5582;
  assign new_P1_U3900 = new_P1_U3444 & new_P1_U5585;
  assign new_P1_U3901 = new_P1_U3444 & new_P1_U5588;
  assign new_P1_U3902 = new_P1_U3444 & new_P1_U5591;
  assign new_P1_U3903 = new_P1_U3444 & new_P1_U5594;
  assign new_P1_U3904 = new_P1_U3444 & new_P1_U5597;
  assign new_P1_U3905 = new_P1_U3444 & new_P1_U5600;
  assign new_P1_U3906 = new_P1_U3907 & new_P1_U5603;
  assign new_P1_U3907 = new_P1_U3444 & new_P1_U5601;
  assign new_P1_U3908 = new_P1_U3444 & new_P1_U5606;
  assign new_P1_U3909 = new_P1_U3444 & new_P1_U5609;
  assign new_P1_U3910 = new_P1_U3444 & new_P1_U5612;
  assign new_P1_U3911 = new_P1_U3444 & new_P1_U5615;
  assign new_P1_U3912 = new_P1_U3444 & new_P1_U5618;
  assign new_P1_U3913 = new_P1_U3444 & new_P1_U5621;
  assign new_P1_U3914 = new_P1_U3444 & new_P1_U5624;
  assign new_P1_U3915 = new_P1_U3444 & new_P1_U5627;
  assign new_P1_U3916 = new_P1_U3444 & new_P1_U5630;
  assign new_P1_U3917 = new_P1_U3444 & new_P1_U5633;
  assign new_P1_U3918 = new_P1_U3919 & new_P1_U5636;
  assign new_P1_U3919 = new_P1_U3444 & new_P1_U5634;
  assign new_P1_U3920 = new_P1_U3921 & new_P1_U5639;
  assign new_P1_U3921 = new_P1_U3444 & new_P1_U5637;
  assign new_P1_U3922 = new_P1_U5645 & new_P1_U5642;
  assign new_P1_U3923 = new_P1_U5649 & new_P1_U5646;
  assign new_P1_U3924 = new_P1_U5651 & new_P1_U5650;
  assign new_P1_U3925 = new_P1_U5655 & new_P1_U5654;
  assign new_P1_U3926 = new_P1_U5659 & new_P1_U5658;
  assign new_P1_U3927 = new_P1_U5663 & new_P1_U5662;
  assign new_P1_U3928 = new_P1_U5675 & new_P1_U5673 & new_P1_U5672;
  assign new_P1_U3929 = new_P1_U5677 & new_P1_U5676;
  assign new_P1_U3930 = new_P1_U5681 & new_P1_U5680;
  assign new_P1_U3931 = new_P1_U5685 & new_P1_U5684;
  assign new_P1_U3932 = new_P1_U5689 & new_P1_U5688;
  assign new_P1_U3933 = new_P1_U5693 & new_P1_U5692;
  assign new_P1_U3934 = new_P1_U5697 & new_P1_U5696;
  assign new_P1_U3935 = new_P1_U5701 & new_P1_U5700;
  assign new_P1_U3936 = new_P1_U5705 & new_P1_U5704;
  assign new_P1_U3937 = new_P1_U5709 & new_P1_U5708;
  assign new_P1_U3938 = new_P1_U5713 & new_P1_U5712;
  assign new_P1_U3939 = new_P1_U5719 & new_P1_U5717 & new_P1_U5716;
  assign new_P1_U3940 = new_P1_U5721 & new_P1_U5720;
  assign new_P1_U3941 = new_P1_U5725 & new_P1_U5724;
  assign new_P1_U3942 = new_P1_U5729 & new_P1_U5728;
  assign new_P1_U3943 = new_P1_U5733 & new_P1_U5732;
  assign new_P1_U3944 = new_P1_U5737 & new_P1_U5736;
  assign new_P1_U3945 = new_P1_U5741 & new_P1_U5740;
  assign new_P1_U3946 = new_P1_U5745 & new_P1_U5744;
  assign new_P1_U3947 = new_P1_U5749 & new_P1_U5748;
  assign new_P1_U3948 = new_P1_U5753 & new_P1_U5752;
  assign new_P1_U3949 = new_P1_U5757 & new_P1_U5756;
  assign new_P1_U3950 = new_P1_U5763 & new_P1_U5761 & new_P1_U5760;
  assign new_P1_U3951 = new_P1_U5765 & new_P1_U5764;
  assign new_P1_U3952 = ~P1_IR_REG_31_;
  assign new_P1_U3953 = ~new_P1_U3022 | ~new_P1_U3360;
  assign new_P1_U3954 = ~new_P1_U5817 | ~new_P1_U5811;
  assign new_P1_U3955 = ~new_P1_U3607 | ~new_P1_U3046;
  assign new_P1_U3956 = ~new_P1_U3726 | ~new_P1_U3046;
  assign new_P1_U3957 = new_P1_U6051 & new_P1_U6050;
  assign new_P1_U3958 = new_P1_U6053 & new_P1_U6052;
  assign new_P1_U3959 = new_P1_U6055 & new_P1_U6054;
  assign new_P1_U3960 = new_P1_U6057 & new_P1_U6056;
  assign new_P1_U3961 = new_P1_U6059 & new_P1_U6058;
  assign new_P1_U3962 = new_P1_U6061 & new_P1_U6060;
  assign new_P1_U3963 = new_P1_U6063 & new_P1_U6062;
  assign new_P1_U3964 = new_P1_U6065 & new_P1_U6064;
  assign new_P1_U3965 = new_P1_U6067 & new_P1_U6066;
  assign new_P1_U3966 = new_P1_U6069 & new_P1_U6068;
  assign new_P1_U3967 = new_P1_U6071 & new_P1_U6070;
  assign new_P1_U3968 = new_P1_U6073 & new_P1_U6072;
  assign new_P1_U3969 = new_P1_U6075 & new_P1_U6074;
  assign new_P1_U3970 = new_P1_U6077 & new_P1_U6076;
  assign new_P1_U3971 = new_P1_U6079 & new_P1_U6078;
  assign new_P1_U3972 = new_P1_U6081 & new_P1_U6080;
  assign new_P1_U3973 = new_P1_U6083 & new_P1_U6082;
  assign new_P1_U3974 = new_P1_U6085 & new_P1_U6084;
  assign new_P1_U3975 = new_P1_U6087 & new_P1_U6086;
  assign new_P1_U3976 = new_P1_U6089 & new_P1_U6088;
  assign new_P1_U3977 = new_P1_U6091 & new_P1_U6090;
  assign new_P1_U3978 = new_P1_U6093 & new_P1_U6092;
  assign new_P1_U3979 = new_P1_U6095 & new_P1_U6094;
  assign new_P1_U3980 = new_P1_U6097 & new_P1_U6096;
  assign new_P1_U3981 = new_P1_U6099 & new_P1_U6098;
  assign new_P1_U3982 = new_P1_U6101 & new_P1_U6100;
  assign new_P1_U3983 = new_P1_U6103 & new_P1_U6102;
  assign new_P1_U3984 = new_P1_U6105 & new_P1_U6104;
  assign new_P1_U3985 = new_P1_U6107 & new_P1_U6106;
  assign new_P1_U3986 = new_P1_U6109 & new_P1_U6108;
  assign new_P1_U3987 = ~new_P1_U3725 | ~new_P1_U3056;
  assign new_P1_U3988 = new_P1_U6111 & new_P1_U6110;
  assign new_P1_U3989 = new_P1_U6113 & new_P1_U6112;
  assign new_P1_U3990 = new_P1_U6179 & new_P1_U6178;
  assign new_P1_U3991 = ~new_P1_U3844 | ~new_P1_U3842 | ~new_P1_U3843;
  assign new_P1_U3992 = ~new_P1_U3371;
  assign new_P1_U3993 = ~new_P1_U3374;
  assign new_P1_U3994 = ~new_P1_U3364;
  assign new_P1_U3995 = ~new_P1_U3423;
  assign new_P1_U3996 = ~new_P1_U4003 | ~new_P1_U5793;
  assign new_P1_U3997 = ~new_P1_U4041 | ~new_P1_U3451;
  assign new_P1_U3998 = ~new_P1_U3419;
  assign new_P1_U3999 = ~new_P1_U4042 | ~new_P1_U5793;
  assign new_P1_U4000 = ~new_P1_U3362;
  assign new_P1_U4001 = ~new_P1_U3367;
  assign new_P1_U4002 = ~new_P1_U3370;
  assign new_P1_U4003 = ~new_P1_U3422;
  assign new_P1_U4004 = ~new_P1_U3366;
  assign new_P1_U4005 = ~new_P1_U3365;
  assign new_P1_U4006 = ~new_P1_U4044 | ~new_P1_U3451;
  assign new_P1_U4007 = ~new_P1_U3361;
  assign new_P1_U4008 = ~new_P1_U3424;
  assign new_P1_U4009 = ~new_P1_U3421;
  assign new_P1_U4010 = ~new_P1_U3993 | ~new_P1_U3453;
  assign new_P1_U4011 = ~new_P1_U3368;
  assign new_P1_U4012 = ~new_P1_U4030 | ~new_P1_U3369;
  assign new_P1_U4013 = ~new_P1_U3873 | ~new_P1_U3425;
  assign new_P1_U4014 = ~new_P1_U3954;
  assign new_P1_U4015 = ~new_P1_U3434;
  assign n1394 = ~new_P1_U3430;
  assign new_P1_U4017 = ~new_P1_U3413;
  assign new_P1_U4018 = ~new_P1_U3411;
  assign new_P1_U4019 = ~new_P1_U3409;
  assign new_P1_U4020 = ~new_P1_U3407;
  assign new_P1_U4021 = ~new_P1_U3405;
  assign new_P1_U4022 = ~new_P1_U3403;
  assign new_P1_U4023 = ~new_P1_U3401;
  assign new_P1_U4024 = ~new_P1_U3399;
  assign new_P1_U4025 = ~new_P1_U3397;
  assign new_P1_U4026 = ~new_P1_U3418;
  assign new_P1_U4027 = ~new_P1_U3417;
  assign new_P1_U4028 = ~new_P1_U3415;
  assign new_P1_U4029 = ~new_P1_U3431;
  assign new_P1_U4030 = ~new_P1_U3372;
  assign new_P1_U4031 = ~new_P1_U3420;
  assign new_P1_U4032 = ~new_P1_U3956;
  assign new_P1_U4033 = ~new_P1_U3955;
  assign new_P1_U4034 = ~new_P1_U3953;
  assign new_P1_U4035 = ~new_P1_U3987;
  assign new_P1_U4036 = ~new_P1_U3373;
  assign new_P1_U4037 = ~new_P1_U3435;
  assign new_P1_U4038 = ~new_P1_U3433;
  assign new_P1_U4039 = ~new_P1_U4009 | ~new_P1_U3022;
  assign new_P1_U4040 = ~n1394 | ~new_P1_U3212;
  assign new_P1_U4041 = ~new_P1_U3375;
  assign new_P1_U4042 = ~new_P1_U3363;
  assign new_P1_U4043 = ~new_P1_U3427;
  assign new_P1_U4044 = ~new_P1_U3369;
  assign new_P1_U4045 = ~new_P1_U3429;
  assign new_P1_U4046 = ~new_P1_U3358;
  assign new_P1_U4047 = ~new_P1_U3357;
  assign new_P1_U4048 = ~new_U125 | ~n1384;
  assign new_P1_U4049 = ~P1_IR_REG_0_ | ~new_P1_U3029;
  assign new_P1_U4050 = ~P1_IR_REG_0_ | ~new_P1_U4047;
  assign new_P1_U4051 = ~new_U114 | ~n1384;
  assign new_P1_U4052 = ~new_P1_SUB_88_U40 | ~new_P1_U3029;
  assign new_P1_U4053 = ~P1_IR_REG_1_ | ~new_P1_U4047;
  assign new_P1_U4054 = ~new_U103 | ~n1384;
  assign new_P1_U4055 = ~new_P1_SUB_88_U21 | ~new_P1_U3029;
  assign new_P1_U4056 = ~P1_IR_REG_2_ | ~new_P1_U4047;
  assign new_P1_U4057 = ~new_U100 | ~n1384;
  assign new_P1_U4058 = ~new_P1_SUB_88_U22 | ~new_P1_U3029;
  assign new_P1_U4059 = ~P1_IR_REG_3_ | ~new_P1_U4047;
  assign new_P1_U4060 = ~new_U99 | ~n1384;
  assign new_P1_U4061 = ~new_P1_SUB_88_U23 | ~new_P1_U3029;
  assign new_P1_U4062 = ~P1_IR_REG_4_ | ~new_P1_U4047;
  assign new_P1_U4063 = ~new_U98 | ~n1384;
  assign new_P1_U4064 = ~new_P1_SUB_88_U162 | ~new_P1_U3029;
  assign new_P1_U4065 = ~P1_IR_REG_5_ | ~new_P1_U4047;
  assign new_P1_U4066 = ~new_U97 | ~n1384;
  assign new_P1_U4067 = ~new_P1_SUB_88_U24 | ~new_P1_U3029;
  assign new_P1_U4068 = ~P1_IR_REG_6_ | ~new_P1_U4047;
  assign new_P1_U4069 = ~new_U96 | ~n1384;
  assign new_P1_U4070 = ~new_P1_SUB_88_U25 | ~new_P1_U3029;
  assign new_P1_U4071 = ~P1_IR_REG_7_ | ~new_P1_U4047;
  assign new_P1_U4072 = ~new_U95 | ~n1384;
  assign new_P1_U4073 = ~new_P1_SUB_88_U26 | ~new_P1_U3029;
  assign new_P1_U4074 = ~P1_IR_REG_8_ | ~new_P1_U4047;
  assign new_P1_U4075 = ~new_U94 | ~n1384;
  assign new_P1_U4076 = ~new_P1_SUB_88_U160 | ~new_P1_U3029;
  assign new_P1_U4077 = ~P1_IR_REG_9_ | ~new_P1_U4047;
  assign new_P1_U4078 = ~new_U124 | ~n1384;
  assign new_P1_U4079 = ~new_P1_SUB_88_U6 | ~new_P1_U3029;
  assign new_P1_U4080 = ~P1_IR_REG_10_ | ~new_P1_U4047;
  assign new_P1_U4081 = ~new_U123 | ~n1384;
  assign new_P1_U4082 = ~new_P1_SUB_88_U7 | ~new_P1_U3029;
  assign new_P1_U4083 = ~P1_IR_REG_11_ | ~new_P1_U4047;
  assign new_P1_U4084 = ~new_U122 | ~n1384;
  assign new_P1_U4085 = ~new_P1_SUB_88_U8 | ~new_P1_U3029;
  assign new_P1_U4086 = ~P1_IR_REG_12_ | ~new_P1_U4047;
  assign new_P1_U4087 = ~new_U121 | ~n1384;
  assign new_P1_U4088 = ~new_P1_SUB_88_U179 | ~new_P1_U3029;
  assign new_P1_U4089 = ~P1_IR_REG_13_ | ~new_P1_U4047;
  assign new_P1_U4090 = ~new_U120 | ~n1384;
  assign new_P1_U4091 = ~new_P1_SUB_88_U9 | ~new_P1_U3029;
  assign new_P1_U4092 = ~P1_IR_REG_14_ | ~new_P1_U4047;
  assign new_P1_U4093 = ~new_U119 | ~n1384;
  assign new_P1_U4094 = ~new_P1_SUB_88_U10 | ~new_P1_U3029;
  assign new_P1_U4095 = ~P1_IR_REG_15_ | ~new_P1_U4047;
  assign new_P1_U4096 = ~new_U118 | ~n1384;
  assign new_P1_U4097 = ~new_P1_SUB_88_U11 | ~new_P1_U3029;
  assign new_P1_U4098 = ~P1_IR_REG_16_ | ~new_P1_U4047;
  assign new_P1_U4099 = ~new_U117 | ~n1384;
  assign new_P1_U4100 = ~new_P1_SUB_88_U177 | ~new_P1_U3029;
  assign new_P1_U4101 = ~P1_IR_REG_17_ | ~new_P1_U4047;
  assign new_P1_U4102 = ~new_U116 | ~n1384;
  assign new_P1_U4103 = ~new_P1_SUB_88_U12 | ~new_P1_U3029;
  assign new_P1_U4104 = ~P1_IR_REG_18_ | ~new_P1_U4047;
  assign new_P1_U4105 = ~new_U115 | ~n1384;
  assign new_P1_U4106 = ~new_P1_SUB_88_U13 | ~new_P1_U3029;
  assign new_P1_U4107 = ~P1_IR_REG_19_ | ~new_P1_U4047;
  assign new_P1_U4108 = ~new_U113 | ~n1384;
  assign new_P1_U4109 = ~new_P1_SUB_88_U14 | ~new_P1_U3029;
  assign new_P1_U4110 = ~P1_IR_REG_20_ | ~new_P1_U4047;
  assign new_P1_U4111 = ~new_U112 | ~n1384;
  assign new_P1_U4112 = ~new_P1_SUB_88_U173 | ~new_P1_U3029;
  assign new_P1_U4113 = ~P1_IR_REG_21_ | ~new_P1_U4047;
  assign new_P1_U4114 = ~new_U111 | ~n1384;
  assign new_P1_U4115 = ~new_P1_SUB_88_U15 | ~new_P1_U3029;
  assign new_P1_U4116 = ~P1_IR_REG_22_ | ~new_P1_U4047;
  assign new_P1_U4117 = ~new_U110 | ~n1384;
  assign new_P1_U4118 = ~new_P1_SUB_88_U16 | ~new_P1_U3029;
  assign new_P1_U4119 = ~P1_IR_REG_23_ | ~new_P1_U4047;
  assign new_P1_U4120 = ~new_U109 | ~n1384;
  assign new_P1_U4121 = ~new_P1_SUB_88_U17 | ~new_P1_U3029;
  assign new_P1_U4122 = ~P1_IR_REG_24_ | ~new_P1_U4047;
  assign new_P1_U4123 = ~new_U108 | ~n1384;
  assign new_P1_U4124 = ~new_P1_SUB_88_U170 | ~new_P1_U3029;
  assign new_P1_U4125 = ~P1_IR_REG_25_ | ~new_P1_U4047;
  assign new_P1_U4126 = ~new_U107 | ~n1384;
  assign new_P1_U4127 = ~new_P1_SUB_88_U18 | ~new_P1_U3029;
  assign new_P1_U4128 = ~P1_IR_REG_26_ | ~new_P1_U4047;
  assign new_P1_U4129 = ~new_U106 | ~n1384;
  assign new_P1_U4130 = ~new_P1_SUB_88_U42 | ~new_P1_U3029;
  assign new_P1_U4131 = ~P1_IR_REG_27_ | ~new_P1_U4047;
  assign new_P1_U4132 = ~new_U105 | ~n1384;
  assign new_P1_U4133 = ~new_P1_SUB_88_U19 | ~new_P1_U3029;
  assign new_P1_U4134 = ~P1_IR_REG_28_ | ~new_P1_U4047;
  assign new_P1_U4135 = ~new_U104 | ~n1384;
  assign new_P1_U4136 = ~new_P1_SUB_88_U20 | ~new_P1_U3029;
  assign new_P1_U4137 = ~P1_IR_REG_29_ | ~new_P1_U4047;
  assign new_P1_U4138 = ~new_U102 | ~n1384;
  assign new_P1_U4139 = ~new_P1_SUB_88_U165 | ~new_P1_U3029;
  assign new_P1_U4140 = ~P1_IR_REG_30_ | ~new_P1_U4047;
  assign new_P1_U4141 = ~new_U101 | ~n1384;
  assign new_P1_U4142 = ~new_P1_SUB_88_U41 | ~new_P1_U3029;
  assign new_P1_U4143 = ~P1_IR_REG_31_ | ~new_P1_U4047;
  assign new_P1_U4144 = ~new_P1_U3360;
  assign new_P1_U4145 = ~new_P1_U3425;
  assign new_P1_U4146 = ~new_P1_U3358 | ~new_P1_U5775;
  assign new_P1_U4147 = ~new_P1_U3358 | ~new_P1_U5778;
  assign new_P1_U4148 = ~new_P1_U4144 | ~P1_D_REG_10_;
  assign new_P1_U4149 = ~new_P1_U4144 | ~P1_D_REG_11_;
  assign new_P1_U4150 = ~new_P1_U4144 | ~P1_D_REG_12_;
  assign new_P1_U4151 = ~new_P1_U4144 | ~P1_D_REG_13_;
  assign new_P1_U4152 = ~new_P1_U4144 | ~P1_D_REG_14_;
  assign new_P1_U4153 = ~new_P1_U4144 | ~P1_D_REG_15_;
  assign new_P1_U4154 = ~new_P1_U4144 | ~P1_D_REG_16_;
  assign new_P1_U4155 = ~new_P1_U4144 | ~P1_D_REG_17_;
  assign new_P1_U4156 = ~new_P1_U4144 | ~P1_D_REG_18_;
  assign new_P1_U4157 = ~new_P1_U4144 | ~P1_D_REG_19_;
  assign new_P1_U4158 = ~new_P1_U4144 | ~P1_D_REG_20_;
  assign new_P1_U4159 = ~new_P1_U4144 | ~P1_D_REG_21_;
  assign new_P1_U4160 = ~new_P1_U4144 | ~P1_D_REG_22_;
  assign new_P1_U4161 = ~new_P1_U4144 | ~P1_D_REG_23_;
  assign new_P1_U4162 = ~new_P1_U4144 | ~P1_D_REG_24_;
  assign new_P1_U4163 = ~new_P1_U4144 | ~P1_D_REG_25_;
  assign new_P1_U4164 = ~new_P1_U4144 | ~P1_D_REG_26_;
  assign new_P1_U4165 = ~new_P1_U4144 | ~P1_D_REG_27_;
  assign new_P1_U4166 = ~new_P1_U4144 | ~P1_D_REG_28_;
  assign new_P1_U4167 = ~new_P1_U4144 | ~P1_D_REG_29_;
  assign new_P1_U4168 = ~new_P1_U4144 | ~P1_D_REG_2_;
  assign new_P1_U4169 = ~new_P1_U4144 | ~P1_D_REG_30_;
  assign new_P1_U4170 = ~new_P1_U4144 | ~P1_D_REG_31_;
  assign new_P1_U4171 = ~new_P1_U4144 | ~P1_D_REG_3_;
  assign new_P1_U4172 = ~new_P1_U4144 | ~P1_D_REG_4_;
  assign new_P1_U4173 = ~new_P1_U4144 | ~P1_D_REG_5_;
  assign new_P1_U4174 = ~new_P1_U4144 | ~P1_D_REG_6_;
  assign new_P1_U4175 = ~new_P1_U4144 | ~P1_D_REG_7_;
  assign new_P1_U4176 = ~new_P1_U4144 | ~P1_D_REG_8_;
  assign new_P1_U4177 = ~new_P1_U4144 | ~P1_D_REG_9_;
  assign new_P1_U4178 = ~new_P1_U5802 | ~new_P1_U5799;
  assign new_P1_U4179 = ~new_P1_U3369 | ~new_P1_U5822 | ~new_P1_U5821;
  assign new_P1_U4180 = ~new_P1_U3018 | ~P1_REG2_REG_1_;
  assign new_P1_U4181 = ~new_P1_U3019 | ~P1_REG1_REG_1_;
  assign new_P1_U4182 = ~new_P1_U3020 | ~P1_REG0_REG_1_;
  assign new_P1_U4183 = ~P1_REG3_REG_1_ | ~new_P1_U3017;
  assign new_P1_U4184 = ~new_P1_U3078;
  assign new_P1_U4185 = ~new_P1_U3419 | ~new_P1_U4010;
  assign new_P1_U4186 = ~new_P1_U4007 | ~new_P1_R1150_U21;
  assign new_P1_U4187 = ~new_P1_U4000 | ~new_P1_R1117_U21;
  assign new_P1_U4188 = ~new_P1_U3994 | ~new_P1_R1138_U96;
  assign new_P1_U4189 = ~new_P1_U4005 | ~new_P1_R1192_U21;
  assign new_P1_U4190 = ~new_P1_U4004 | ~new_P1_R1207_U21;
  assign new_P1_U4191 = ~new_P1_U4011 | ~new_P1_R1171_U96;
  assign new_P1_U4192 = ~new_P1_U3992 | ~new_P1_R1240_U96;
  assign new_P1_U4193 = ~new_P1_U3376;
  assign new_P1_U4194 = ~new_P1_U3025 | ~new_P1_U3078;
  assign new_P1_U4195 = ~new_P1_R1222_U96 | ~new_P1_U3024;
  assign new_P1_U4196 = ~new_P1_U3456 | ~new_P1_U4036;
  assign new_P1_U4197 = ~new_P1_U3456 | ~new_P1_U4185;
  assign new_P1_U4198 = ~new_P1_U4193 | ~new_P1_U3595 | ~new_P1_U4197 | ~new_P1_U4194;
  assign new_P1_U4199 = ~P1_REG2_REG_2_ | ~new_P1_U3018;
  assign new_P1_U4200 = ~P1_REG1_REG_2_ | ~new_P1_U3019;
  assign new_P1_U4201 = ~P1_REG0_REG_2_ | ~new_P1_U3020;
  assign new_P1_U4202 = ~P1_REG3_REG_2_ | ~new_P1_U3017;
  assign new_P1_U4203 = ~new_P1_U3068;
  assign new_P1_U4204 = ~P1_REG0_REG_0_ | ~new_P1_U3020;
  assign new_P1_U4205 = ~P1_REG1_REG_0_ | ~new_P1_U3019;
  assign new_P1_U4206 = ~P1_REG2_REG_0_ | ~new_P1_U3018;
  assign new_P1_U4207 = ~P1_REG3_REG_0_ | ~new_P1_U3017;
  assign new_P1_U4208 = ~new_P1_U3077;
  assign new_P1_U4209 = ~new_P1_U3034 | ~new_P1_U3077;
  assign new_P1_U4210 = ~new_P1_R1150_U98 | ~new_P1_U4007;
  assign new_P1_U4211 = ~new_P1_R1117_U98 | ~new_P1_U4000;
  assign new_P1_U4212 = ~new_P1_R1138_U95 | ~new_P1_U3994;
  assign new_P1_U4213 = ~new_P1_R1192_U98 | ~new_P1_U4005;
  assign new_P1_U4214 = ~new_P1_R1207_U98 | ~new_P1_U4004;
  assign new_P1_U4215 = ~new_P1_R1171_U95 | ~new_P1_U4011;
  assign new_P1_U4216 = ~new_P1_R1240_U95 | ~new_P1_U3992;
  assign new_P1_U4217 = ~new_P1_U3378;
  assign new_P1_U4218 = ~new_P1_U3025 | ~new_P1_U3068;
  assign new_P1_U4219 = ~new_P1_R1222_U95 | ~new_P1_U3024;
  assign new_P1_U4220 = ~new_P1_R1282_U56 | ~new_P1_U4036;
  assign new_P1_U4221 = ~new_P1_U3461 | ~new_P1_U4185;
  assign new_P1_U4222 = ~new_P1_U3611 | ~new_P1_U4217;
  assign new_P1_U4223 = ~P1_REG2_REG_3_ | ~new_P1_U3018;
  assign new_P1_U4224 = ~P1_REG1_REG_3_ | ~new_P1_U3019;
  assign new_P1_U4225 = ~P1_REG0_REG_3_ | ~new_P1_U3020;
  assign new_P1_U4226 = ~new_P1_ADD_99_U4 | ~new_P1_U3017;
  assign new_P1_U4227 = ~new_P1_U3064;
  assign new_P1_U4228 = ~new_P1_U3034 | ~new_P1_U3078;
  assign new_P1_U4229 = ~new_P1_R1150_U108 | ~new_P1_U4007;
  assign new_P1_U4230 = ~new_P1_R1117_U108 | ~new_P1_U4000;
  assign new_P1_U4231 = ~new_P1_R1138_U17 | ~new_P1_U3994;
  assign new_P1_U4232 = ~new_P1_R1192_U108 | ~new_P1_U4005;
  assign new_P1_U4233 = ~new_P1_R1207_U108 | ~new_P1_U4004;
  assign new_P1_U4234 = ~new_P1_R1171_U17 | ~new_P1_U4011;
  assign new_P1_U4235 = ~new_P1_R1240_U17 | ~new_P1_U3992;
  assign new_P1_U4236 = ~new_P1_U3379;
  assign new_P1_U4237 = ~new_P1_U3025 | ~new_P1_U3064;
  assign new_P1_U4238 = ~new_P1_R1222_U17 | ~new_P1_U3024;
  assign new_P1_U4239 = ~new_P1_R1282_U18 | ~new_P1_U4036;
  assign new_P1_U4240 = ~new_P1_U3464 | ~new_P1_U4185;
  assign new_P1_U4241 = ~new_P1_U3615 | ~new_P1_U4236;
  assign new_P1_U4242 = ~P1_REG2_REG_4_ | ~new_P1_U3018;
  assign new_P1_U4243 = ~P1_REG1_REG_4_ | ~new_P1_U3019;
  assign new_P1_U4244 = ~P1_REG0_REG_4_ | ~new_P1_U3020;
  assign new_P1_U4245 = ~new_P1_ADD_99_U59 | ~new_P1_U3017;
  assign new_P1_U4246 = ~new_P1_U3060;
  assign new_P1_U4247 = ~new_P1_U3034 | ~new_P1_U3068;
  assign new_P1_U4248 = ~new_P1_R1150_U18 | ~new_P1_U4007;
  assign new_P1_U4249 = ~new_P1_R1117_U18 | ~new_P1_U4000;
  assign new_P1_U4250 = ~new_P1_R1138_U101 | ~new_P1_U3994;
  assign new_P1_U4251 = ~new_P1_R1192_U18 | ~new_P1_U4005;
  assign new_P1_U4252 = ~new_P1_R1207_U18 | ~new_P1_U4004;
  assign new_P1_U4253 = ~new_P1_R1171_U101 | ~new_P1_U4011;
  assign new_P1_U4254 = ~new_P1_R1240_U101 | ~new_P1_U3992;
  assign new_P1_U4255 = ~new_P1_U3380;
  assign new_P1_U4256 = ~new_P1_U3025 | ~new_P1_U3060;
  assign new_P1_U4257 = ~new_P1_R1222_U101 | ~new_P1_U3024;
  assign new_P1_U4258 = ~new_P1_R1282_U20 | ~new_P1_U4036;
  assign new_P1_U4259 = ~new_P1_U3467 | ~new_P1_U4185;
  assign new_P1_U4260 = ~new_P1_U3619 | ~new_P1_U4255;
  assign new_P1_U4261 = ~P1_REG2_REG_5_ | ~new_P1_U3018;
  assign new_P1_U4262 = ~P1_REG1_REG_5_ | ~new_P1_U3019;
  assign new_P1_U4263 = ~P1_REG0_REG_5_ | ~new_P1_U3020;
  assign new_P1_U4264 = ~new_P1_ADD_99_U58 | ~new_P1_U3017;
  assign new_P1_U4265 = ~new_P1_U3067;
  assign new_P1_U4266 = ~new_P1_U3034 | ~new_P1_U3064;
  assign new_P1_U4267 = ~new_P1_R1150_U107 | ~new_P1_U4007;
  assign new_P1_U4268 = ~new_P1_R1117_U107 | ~new_P1_U4000;
  assign new_P1_U4269 = ~new_P1_R1138_U100 | ~new_P1_U3994;
  assign new_P1_U4270 = ~new_P1_R1192_U107 | ~new_P1_U4005;
  assign new_P1_U4271 = ~new_P1_R1207_U107 | ~new_P1_U4004;
  assign new_P1_U4272 = ~new_P1_R1171_U100 | ~new_P1_U4011;
  assign new_P1_U4273 = ~new_P1_R1240_U100 | ~new_P1_U3992;
  assign new_P1_U4274 = ~new_P1_U3381;
  assign new_P1_U4275 = ~new_P1_U3025 | ~new_P1_U3067;
  assign new_P1_U4276 = ~new_P1_R1222_U100 | ~new_P1_U3024;
  assign new_P1_U4277 = ~new_P1_R1282_U21 | ~new_P1_U4036;
  assign new_P1_U4278 = ~new_P1_U3470 | ~new_P1_U4185;
  assign new_P1_U4279 = ~new_P1_U3623 | ~new_P1_U4274;
  assign new_P1_U4280 = ~P1_REG2_REG_6_ | ~new_P1_U3018;
  assign new_P1_U4281 = ~P1_REG1_REG_6_ | ~new_P1_U3019;
  assign new_P1_U4282 = ~P1_REG0_REG_6_ | ~new_P1_U3020;
  assign new_P1_U4283 = ~new_P1_ADD_99_U57 | ~new_P1_U3017;
  assign new_P1_U4284 = ~new_P1_U3071;
  assign new_P1_U4285 = ~new_P1_U3034 | ~new_P1_U3060;
  assign new_P1_U4286 = ~new_P1_R1150_U106 | ~new_P1_U4007;
  assign new_P1_U4287 = ~new_P1_R1117_U106 | ~new_P1_U4000;
  assign new_P1_U4288 = ~new_P1_R1138_U18 | ~new_P1_U3994;
  assign new_P1_U4289 = ~new_P1_R1192_U106 | ~new_P1_U4005;
  assign new_P1_U4290 = ~new_P1_R1207_U106 | ~new_P1_U4004;
  assign new_P1_U4291 = ~new_P1_R1171_U18 | ~new_P1_U4011;
  assign new_P1_U4292 = ~new_P1_R1240_U18 | ~new_P1_U3992;
  assign new_P1_U4293 = ~new_P1_U3382;
  assign new_P1_U4294 = ~new_P1_U3025 | ~new_P1_U3071;
  assign new_P1_U4295 = ~new_P1_R1222_U18 | ~new_P1_U3024;
  assign new_P1_U4296 = ~new_P1_R1282_U65 | ~new_P1_U4036;
  assign new_P1_U4297 = ~new_P1_U3473 | ~new_P1_U4185;
  assign new_P1_U4298 = ~new_P1_U3627 | ~new_P1_U4293;
  assign new_P1_U4299 = ~P1_REG2_REG_7_ | ~new_P1_U3018;
  assign new_P1_U4300 = ~P1_REG1_REG_7_ | ~new_P1_U3019;
  assign new_P1_U4301 = ~P1_REG0_REG_7_ | ~new_P1_U3020;
  assign new_P1_U4302 = ~new_P1_ADD_99_U56 | ~new_P1_U3017;
  assign new_P1_U4303 = ~new_P1_U3070;
  assign new_P1_U4304 = ~new_P1_U3034 | ~new_P1_U3067;
  assign new_P1_U4305 = ~new_P1_R1150_U19 | ~new_P1_U4007;
  assign new_P1_U4306 = ~new_P1_R1117_U19 | ~new_P1_U4000;
  assign new_P1_U4307 = ~new_P1_R1138_U99 | ~new_P1_U3994;
  assign new_P1_U4308 = ~new_P1_R1192_U19 | ~new_P1_U4005;
  assign new_P1_U4309 = ~new_P1_R1207_U19 | ~new_P1_U4004;
  assign new_P1_U4310 = ~new_P1_R1171_U99 | ~new_P1_U4011;
  assign new_P1_U4311 = ~new_P1_R1240_U99 | ~new_P1_U3992;
  assign new_P1_U4312 = ~new_P1_U3383;
  assign new_P1_U4313 = ~new_P1_U3025 | ~new_P1_U3070;
  assign new_P1_U4314 = ~new_P1_R1222_U99 | ~new_P1_U3024;
  assign new_P1_U4315 = ~new_P1_R1282_U22 | ~new_P1_U4036;
  assign new_P1_U4316 = ~new_P1_U3476 | ~new_P1_U4185;
  assign new_P1_U4317 = ~new_P1_U3631 | ~new_P1_U4312;
  assign new_P1_U4318 = ~P1_REG2_REG_8_ | ~new_P1_U3018;
  assign new_P1_U4319 = ~P1_REG1_REG_8_ | ~new_P1_U3019;
  assign new_P1_U4320 = ~P1_REG0_REG_8_ | ~new_P1_U3020;
  assign new_P1_U4321 = ~new_P1_ADD_99_U55 | ~new_P1_U3017;
  assign new_P1_U4322 = ~new_P1_U3084;
  assign new_P1_U4323 = ~new_P1_U3034 | ~new_P1_U3071;
  assign new_P1_U4324 = ~new_P1_R1150_U105 | ~new_P1_U4007;
  assign new_P1_U4325 = ~new_P1_R1117_U105 | ~new_P1_U4000;
  assign new_P1_U4326 = ~new_P1_R1138_U19 | ~new_P1_U3994;
  assign new_P1_U4327 = ~new_P1_R1192_U105 | ~new_P1_U4005;
  assign new_P1_U4328 = ~new_P1_R1207_U105 | ~new_P1_U4004;
  assign new_P1_U4329 = ~new_P1_R1171_U19 | ~new_P1_U4011;
  assign new_P1_U4330 = ~new_P1_R1240_U19 | ~new_P1_U3992;
  assign new_P1_U4331 = ~new_P1_U3384;
  assign new_P1_U4332 = ~new_P1_U3025 | ~new_P1_U3084;
  assign new_P1_U4333 = ~new_P1_R1222_U19 | ~new_P1_U3024;
  assign new_P1_U4334 = ~new_P1_R1282_U23 | ~new_P1_U4036;
  assign new_P1_U4335 = ~new_P1_U3479 | ~new_P1_U4185;
  assign new_P1_U4336 = ~new_P1_U3635 | ~new_P1_U4331;
  assign new_P1_U4337 = ~P1_REG2_REG_9_ | ~new_P1_U3018;
  assign new_P1_U4338 = ~P1_REG1_REG_9_ | ~new_P1_U3019;
  assign new_P1_U4339 = ~P1_REG0_REG_9_ | ~new_P1_U3020;
  assign new_P1_U4340 = ~new_P1_ADD_99_U54 | ~new_P1_U3017;
  assign new_P1_U4341 = ~new_P1_U3083;
  assign new_P1_U4342 = ~new_P1_U3034 | ~new_P1_U3070;
  assign new_P1_U4343 = ~new_P1_R1150_U20 | ~new_P1_U4007;
  assign new_P1_U4344 = ~new_P1_R1117_U20 | ~new_P1_U4000;
  assign new_P1_U4345 = ~new_P1_R1138_U98 | ~new_P1_U3994;
  assign new_P1_U4346 = ~new_P1_R1192_U20 | ~new_P1_U4005;
  assign new_P1_U4347 = ~new_P1_R1207_U20 | ~new_P1_U4004;
  assign new_P1_U4348 = ~new_P1_R1171_U98 | ~new_P1_U4011;
  assign new_P1_U4349 = ~new_P1_R1240_U98 | ~new_P1_U3992;
  assign new_P1_U4350 = ~new_P1_U3385;
  assign new_P1_U4351 = ~new_P1_U3025 | ~new_P1_U3083;
  assign new_P1_U4352 = ~new_P1_R1222_U98 | ~new_P1_U3024;
  assign new_P1_U4353 = ~new_P1_R1282_U24 | ~new_P1_U4036;
  assign new_P1_U4354 = ~new_P1_U3482 | ~new_P1_U4185;
  assign new_P1_U4355 = ~new_P1_U3639 | ~new_P1_U4350;
  assign new_P1_U4356 = ~P1_REG2_REG_10_ | ~new_P1_U3018;
  assign new_P1_U4357 = ~P1_REG1_REG_10_ | ~new_P1_U3019;
  assign new_P1_U4358 = ~P1_REG0_REG_10_ | ~new_P1_U3020;
  assign new_P1_U4359 = ~new_P1_ADD_99_U78 | ~new_P1_U3017;
  assign new_P1_U4360 = ~new_P1_U3062;
  assign new_P1_U4361 = ~new_P1_U3034 | ~new_P1_U3084;
  assign new_P1_U4362 = ~new_P1_R1150_U104 | ~new_P1_U4007;
  assign new_P1_U4363 = ~new_P1_R1117_U104 | ~new_P1_U4000;
  assign new_P1_U4364 = ~new_P1_R1138_U97 | ~new_P1_U3994;
  assign new_P1_U4365 = ~new_P1_R1192_U104 | ~new_P1_U4005;
  assign new_P1_U4366 = ~new_P1_R1207_U104 | ~new_P1_U4004;
  assign new_P1_U4367 = ~new_P1_R1171_U97 | ~new_P1_U4011;
  assign new_P1_U4368 = ~new_P1_R1240_U97 | ~new_P1_U3992;
  assign new_P1_U4369 = ~new_P1_U3386;
  assign new_P1_U4370 = ~new_P1_U3025 | ~new_P1_U3062;
  assign new_P1_U4371 = ~new_P1_R1222_U97 | ~new_P1_U3024;
  assign new_P1_U4372 = ~new_P1_R1282_U63 | ~new_P1_U4036;
  assign new_P1_U4373 = ~new_P1_U3485 | ~new_P1_U4185;
  assign new_P1_U4374 = ~new_P1_U3643 | ~new_P1_U4369;
  assign new_P1_U4375 = ~P1_REG2_REG_11_ | ~new_P1_U3018;
  assign new_P1_U4376 = ~P1_REG1_REG_11_ | ~new_P1_U3019;
  assign new_P1_U4377 = ~P1_REG0_REG_11_ | ~new_P1_U3020;
  assign new_P1_U4378 = ~new_P1_ADD_99_U77 | ~new_P1_U3017;
  assign new_P1_U4379 = ~new_P1_U3063;
  assign new_P1_U4380 = ~new_P1_U3034 | ~new_P1_U3083;
  assign new_P1_U4381 = ~new_P1_R1150_U114 | ~new_P1_U4007;
  assign new_P1_U4382 = ~new_P1_R1117_U114 | ~new_P1_U4000;
  assign new_P1_U4383 = ~new_P1_R1138_U11 | ~new_P1_U3994;
  assign new_P1_U4384 = ~new_P1_R1192_U114 | ~new_P1_U4005;
  assign new_P1_U4385 = ~new_P1_R1207_U114 | ~new_P1_U4004;
  assign new_P1_U4386 = ~new_P1_R1171_U11 | ~new_P1_U4011;
  assign new_P1_U4387 = ~new_P1_R1240_U11 | ~new_P1_U3992;
  assign new_P1_U4388 = ~new_P1_U3387;
  assign new_P1_U4389 = ~new_P1_U3025 | ~new_P1_U3063;
  assign new_P1_U4390 = ~new_P1_R1222_U11 | ~new_P1_U3024;
  assign new_P1_U4391 = ~new_P1_R1282_U6 | ~new_P1_U4036;
  assign new_P1_U4392 = ~new_P1_U3488 | ~new_P1_U4185;
  assign new_P1_U4393 = ~new_P1_U3647 | ~new_P1_U4388;
  assign new_P1_U4394 = ~P1_REG2_REG_12_ | ~new_P1_U3018;
  assign new_P1_U4395 = ~P1_REG1_REG_12_ | ~new_P1_U3019;
  assign new_P1_U4396 = ~P1_REG0_REG_12_ | ~new_P1_U3020;
  assign new_P1_U4397 = ~new_P1_ADD_99_U76 | ~new_P1_U3017;
  assign new_P1_U4398 = ~new_P1_U3072;
  assign new_P1_U4399 = ~new_P1_U3034 | ~new_P1_U3062;
  assign new_P1_U4400 = ~new_P1_R1150_U13 | ~new_P1_U4007;
  assign new_P1_U4401 = ~new_P1_R1117_U13 | ~new_P1_U4000;
  assign new_P1_U4402 = ~new_P1_R1138_U115 | ~new_P1_U3994;
  assign new_P1_U4403 = ~new_P1_R1192_U13 | ~new_P1_U4005;
  assign new_P1_U4404 = ~new_P1_R1207_U13 | ~new_P1_U4004;
  assign new_P1_U4405 = ~new_P1_R1171_U115 | ~new_P1_U4011;
  assign new_P1_U4406 = ~new_P1_R1240_U115 | ~new_P1_U3992;
  assign new_P1_U4407 = ~new_P1_U3388;
  assign new_P1_U4408 = ~new_P1_U3025 | ~new_P1_U3072;
  assign new_P1_U4409 = ~new_P1_R1222_U115 | ~new_P1_U3024;
  assign new_P1_U4410 = ~new_P1_R1282_U7 | ~new_P1_U4036;
  assign new_P1_U4411 = ~new_P1_U3491 | ~new_P1_U4185;
  assign new_P1_U4412 = ~new_P1_U3651 | ~new_P1_U4407;
  assign new_P1_U4413 = ~P1_REG2_REG_13_ | ~new_P1_U3018;
  assign new_P1_U4414 = ~P1_REG1_REG_13_ | ~new_P1_U3019;
  assign new_P1_U4415 = ~P1_REG0_REG_13_ | ~new_P1_U3020;
  assign new_P1_U4416 = ~new_P1_ADD_99_U75 | ~new_P1_U3017;
  assign new_P1_U4417 = ~new_P1_U3080;
  assign new_P1_U4418 = ~new_P1_U3034 | ~new_P1_U3063;
  assign new_P1_U4419 = ~new_P1_R1150_U103 | ~new_P1_U4007;
  assign new_P1_U4420 = ~new_P1_R1117_U103 | ~new_P1_U4000;
  assign new_P1_U4421 = ~new_P1_R1138_U114 | ~new_P1_U3994;
  assign new_P1_U4422 = ~new_P1_R1192_U103 | ~new_P1_U4005;
  assign new_P1_U4423 = ~new_P1_R1207_U103 | ~new_P1_U4004;
  assign new_P1_U4424 = ~new_P1_R1171_U114 | ~new_P1_U4011;
  assign new_P1_U4425 = ~new_P1_R1240_U114 | ~new_P1_U3992;
  assign new_P1_U4426 = ~new_P1_U3389;
  assign new_P1_U4427 = ~new_P1_U3025 | ~new_P1_U3080;
  assign new_P1_U4428 = ~new_P1_R1222_U114 | ~new_P1_U3024;
  assign new_P1_U4429 = ~new_P1_R1282_U8 | ~new_P1_U4036;
  assign new_P1_U4430 = ~new_P1_U3494 | ~new_P1_U4185;
  assign new_P1_U4431 = ~new_P1_U3655 | ~new_P1_U4426;
  assign new_P1_U4432 = ~P1_REG2_REG_14_ | ~new_P1_U3018;
  assign new_P1_U4433 = ~P1_REG1_REG_14_ | ~new_P1_U3019;
  assign new_P1_U4434 = ~P1_REG0_REG_14_ | ~new_P1_U3020;
  assign new_P1_U4435 = ~new_P1_ADD_99_U74 | ~new_P1_U3017;
  assign new_P1_U4436 = ~new_P1_U3079;
  assign new_P1_U4437 = ~new_P1_U3034 | ~new_P1_U3072;
  assign new_P1_U4438 = ~new_P1_R1150_U102 | ~new_P1_U4007;
  assign new_P1_U4439 = ~new_P1_R1117_U102 | ~new_P1_U4000;
  assign new_P1_U4440 = ~new_P1_R1138_U12 | ~new_P1_U3994;
  assign new_P1_U4441 = ~new_P1_R1192_U102 | ~new_P1_U4005;
  assign new_P1_U4442 = ~new_P1_R1207_U102 | ~new_P1_U4004;
  assign new_P1_U4443 = ~new_P1_R1171_U12 | ~new_P1_U4011;
  assign new_P1_U4444 = ~new_P1_R1240_U12 | ~new_P1_U3992;
  assign new_P1_U4445 = ~new_P1_U3390;
  assign new_P1_U4446 = ~new_P1_U3025 | ~new_P1_U3079;
  assign new_P1_U4447 = ~new_P1_R1222_U12 | ~new_P1_U3024;
  assign new_P1_U4448 = ~new_P1_R1282_U86 | ~new_P1_U4036;
  assign new_P1_U4449 = ~new_P1_U3497 | ~new_P1_U4185;
  assign new_P1_U4450 = ~new_P1_U3659 | ~new_P1_U4445;
  assign new_P1_U4451 = ~P1_REG2_REG_15_ | ~new_P1_U3018;
  assign new_P1_U4452 = ~P1_REG1_REG_15_ | ~new_P1_U3019;
  assign new_P1_U4453 = ~P1_REG0_REG_15_ | ~new_P1_U3020;
  assign new_P1_U4454 = ~new_P1_ADD_99_U73 | ~new_P1_U3017;
  assign new_P1_U4455 = ~new_P1_U3074;
  assign new_P1_U4456 = ~new_P1_U3034 | ~new_P1_U3080;
  assign new_P1_U4457 = ~new_P1_R1150_U113 | ~new_P1_U4007;
  assign new_P1_U4458 = ~new_P1_R1117_U113 | ~new_P1_U4000;
  assign new_P1_U4459 = ~new_P1_R1138_U113 | ~new_P1_U3994;
  assign new_P1_U4460 = ~new_P1_R1192_U113 | ~new_P1_U4005;
  assign new_P1_U4461 = ~new_P1_R1207_U113 | ~new_P1_U4004;
  assign new_P1_U4462 = ~new_P1_R1171_U113 | ~new_P1_U4011;
  assign new_P1_U4463 = ~new_P1_R1240_U113 | ~new_P1_U3992;
  assign new_P1_U4464 = ~new_P1_U3391;
  assign new_P1_U4465 = ~new_P1_U3025 | ~new_P1_U3074;
  assign new_P1_U4466 = ~new_P1_R1222_U113 | ~new_P1_U3024;
  assign new_P1_U4467 = ~new_P1_R1282_U9 | ~new_P1_U4036;
  assign new_P1_U4468 = ~new_P1_U3500 | ~new_P1_U4185;
  assign new_P1_U4469 = ~new_P1_U3663 | ~new_P1_U4464;
  assign new_P1_U4470 = ~P1_REG2_REG_16_ | ~new_P1_U3018;
  assign new_P1_U4471 = ~P1_REG1_REG_16_ | ~new_P1_U3019;
  assign new_P1_U4472 = ~P1_REG0_REG_16_ | ~new_P1_U3020;
  assign new_P1_U4473 = ~new_P1_ADD_99_U72 | ~new_P1_U3017;
  assign new_P1_U4474 = ~new_P1_U3073;
  assign new_P1_U4475 = ~new_P1_U3034 | ~new_P1_U3079;
  assign new_P1_U4476 = ~new_P1_R1150_U112 | ~new_P1_U4007;
  assign new_P1_U4477 = ~new_P1_R1117_U112 | ~new_P1_U4000;
  assign new_P1_U4478 = ~new_P1_R1138_U112 | ~new_P1_U3994;
  assign new_P1_U4479 = ~new_P1_R1192_U112 | ~new_P1_U4005;
  assign new_P1_U4480 = ~new_P1_R1207_U112 | ~new_P1_U4004;
  assign new_P1_U4481 = ~new_P1_R1171_U112 | ~new_P1_U4011;
  assign new_P1_U4482 = ~new_P1_R1240_U112 | ~new_P1_U3992;
  assign new_P1_U4483 = ~new_P1_U3392;
  assign new_P1_U4484 = ~new_P1_U3025 | ~new_P1_U3073;
  assign new_P1_U4485 = ~new_P1_R1222_U112 | ~new_P1_U3024;
  assign new_P1_U4486 = ~new_P1_R1282_U10 | ~new_P1_U4036;
  assign new_P1_U4487 = ~new_P1_U3503 | ~new_P1_U4185;
  assign new_P1_U4488 = ~new_P1_U3667 | ~new_P1_U4483;
  assign new_P1_U4489 = ~P1_REG2_REG_17_ | ~new_P1_U3018;
  assign new_P1_U4490 = ~P1_REG1_REG_17_ | ~new_P1_U3019;
  assign new_P1_U4491 = ~P1_REG0_REG_17_ | ~new_P1_U3020;
  assign new_P1_U4492 = ~new_P1_ADD_99_U71 | ~new_P1_U3017;
  assign new_P1_U4493 = ~new_P1_U3069;
  assign new_P1_U4494 = ~new_P1_U3034 | ~new_P1_U3074;
  assign new_P1_U4495 = ~new_P1_R1150_U14 | ~new_P1_U4007;
  assign new_P1_U4496 = ~new_P1_R1117_U14 | ~new_P1_U4000;
  assign new_P1_U4497 = ~new_P1_R1138_U111 | ~new_P1_U3994;
  assign new_P1_U4498 = ~new_P1_R1192_U14 | ~new_P1_U4005;
  assign new_P1_U4499 = ~new_P1_R1207_U14 | ~new_P1_U4004;
  assign new_P1_U4500 = ~new_P1_R1171_U111 | ~new_P1_U4011;
  assign new_P1_U4501 = ~new_P1_R1240_U111 | ~new_P1_U3992;
  assign new_P1_U4502 = ~new_P1_U3393;
  assign new_P1_U4503 = ~new_P1_U3025 | ~new_P1_U3069;
  assign new_P1_U4504 = ~new_P1_R1222_U111 | ~new_P1_U3024;
  assign new_P1_U4505 = ~new_P1_R1282_U11 | ~new_P1_U4036;
  assign new_P1_U4506 = ~new_P1_U3506 | ~new_P1_U4185;
  assign new_P1_U4507 = ~new_P1_U3671 | ~new_P1_U4502;
  assign new_P1_U4508 = ~P1_REG2_REG_18_ | ~new_P1_U3018;
  assign new_P1_U4509 = ~P1_REG1_REG_18_ | ~new_P1_U3019;
  assign new_P1_U4510 = ~P1_REG0_REG_18_ | ~new_P1_U3020;
  assign new_P1_U4511 = ~new_P1_ADD_99_U70 | ~new_P1_U3017;
  assign new_P1_U4512 = ~new_P1_U3082;
  assign new_P1_U4513 = ~new_P1_U3034 | ~new_P1_U3073;
  assign new_P1_U4514 = ~new_P1_R1150_U101 | ~new_P1_U4007;
  assign new_P1_U4515 = ~new_P1_R1117_U101 | ~new_P1_U4000;
  assign new_P1_U4516 = ~new_P1_R1138_U13 | ~new_P1_U3994;
  assign new_P1_U4517 = ~new_P1_R1192_U101 | ~new_P1_U4005;
  assign new_P1_U4518 = ~new_P1_R1207_U101 | ~new_P1_U4004;
  assign new_P1_U4519 = ~new_P1_R1171_U13 | ~new_P1_U4011;
  assign new_P1_U4520 = ~new_P1_R1240_U13 | ~new_P1_U3992;
  assign new_P1_U4521 = ~new_P1_U3394;
  assign new_P1_U4522 = ~new_P1_U3025 | ~new_P1_U3082;
  assign new_P1_U4523 = ~new_P1_R1222_U13 | ~new_P1_U3024;
  assign new_P1_U4524 = ~new_P1_R1282_U84 | ~new_P1_U4036;
  assign new_P1_U4525 = ~new_P1_U3509 | ~new_P1_U4185;
  assign new_P1_U4526 = ~new_P1_U3675 | ~new_P1_U4521;
  assign new_P1_U4527 = ~P1_REG2_REG_19_ | ~new_P1_U3018;
  assign new_P1_U4528 = ~P1_REG1_REG_19_ | ~new_P1_U3019;
  assign new_P1_U4529 = ~P1_REG0_REG_19_ | ~new_P1_U3020;
  assign new_P1_U4530 = ~new_P1_ADD_99_U69 | ~new_P1_U3017;
  assign new_P1_U4531 = ~new_P1_U3081;
  assign new_P1_U4532 = ~new_P1_U3034 | ~new_P1_U3069;
  assign new_P1_U4533 = ~new_P1_R1150_U100 | ~new_P1_U4007;
  assign new_P1_U4534 = ~new_P1_R1117_U100 | ~new_P1_U4000;
  assign new_P1_U4535 = ~new_P1_R1138_U110 | ~new_P1_U3994;
  assign new_P1_U4536 = ~new_P1_R1192_U100 | ~new_P1_U4005;
  assign new_P1_U4537 = ~new_P1_R1207_U100 | ~new_P1_U4004;
  assign new_P1_U4538 = ~new_P1_R1171_U110 | ~new_P1_U4011;
  assign new_P1_U4539 = ~new_P1_R1240_U110 | ~new_P1_U3992;
  assign new_P1_U4540 = ~new_P1_U3395;
  assign new_P1_U4541 = ~new_P1_U3025 | ~new_P1_U3081;
  assign new_P1_U4542 = ~new_P1_R1222_U110 | ~new_P1_U3024;
  assign new_P1_U4543 = ~new_P1_R1282_U12 | ~new_P1_U4036;
  assign new_P1_U4544 = ~new_P1_U3512 | ~new_P1_U4185;
  assign new_P1_U4545 = ~new_P1_U3679 | ~new_P1_U4540;
  assign new_P1_U4546 = ~P1_REG2_REG_20_ | ~new_P1_U3018;
  assign new_P1_U4547 = ~P1_REG1_REG_20_ | ~new_P1_U3019;
  assign new_P1_U4548 = ~P1_REG0_REG_20_ | ~new_P1_U3020;
  assign new_P1_U4549 = ~new_P1_ADD_99_U68 | ~new_P1_U3017;
  assign new_P1_U4550 = ~new_P1_U3076;
  assign new_P1_U4551 = ~new_P1_U3034 | ~new_P1_U3082;
  assign new_P1_U4552 = ~new_P1_R1150_U99 | ~new_P1_U4007;
  assign new_P1_U4553 = ~new_P1_R1117_U99 | ~new_P1_U4000;
  assign new_P1_U4554 = ~new_P1_R1138_U109 | ~new_P1_U3994;
  assign new_P1_U4555 = ~new_P1_R1192_U99 | ~new_P1_U4005;
  assign new_P1_U4556 = ~new_P1_R1207_U99 | ~new_P1_U4004;
  assign new_P1_U4557 = ~new_P1_R1171_U109 | ~new_P1_U4011;
  assign new_P1_U4558 = ~new_P1_R1240_U109 | ~new_P1_U3992;
  assign new_P1_U4559 = ~new_P1_U3396;
  assign new_P1_U4560 = ~new_P1_U3025 | ~new_P1_U3076;
  assign new_P1_U4561 = ~new_P1_R1222_U109 | ~new_P1_U3024;
  assign new_P1_U4562 = ~new_P1_R1282_U82 | ~new_P1_U4036;
  assign new_P1_U4563 = ~new_P1_U3514 | ~new_P1_U4185;
  assign new_P1_U4564 = ~new_P1_U3683 | ~new_P1_U4559;
  assign new_P1_U4565 = ~P1_REG2_REG_21_ | ~new_P1_U3018;
  assign new_P1_U4566 = ~P1_REG1_REG_21_ | ~new_P1_U3019;
  assign new_P1_U4567 = ~P1_REG0_REG_21_ | ~new_P1_U3020;
  assign new_P1_U4568 = ~new_P1_ADD_99_U67 | ~new_P1_U3017;
  assign new_P1_U4569 = ~new_P1_U3075;
  assign new_P1_U4570 = ~new_P1_U3034 | ~new_P1_U3081;
  assign new_P1_U4571 = ~new_P1_R1150_U97 | ~new_P1_U4007;
  assign new_P1_U4572 = ~new_P1_R1117_U97 | ~new_P1_U4000;
  assign new_P1_U4573 = ~new_P1_R1138_U14 | ~new_P1_U3994;
  assign new_P1_U4574 = ~new_P1_R1192_U97 | ~new_P1_U4005;
  assign new_P1_U4575 = ~new_P1_R1207_U97 | ~new_P1_U4004;
  assign new_P1_U4576 = ~new_P1_R1171_U14 | ~new_P1_U4011;
  assign new_P1_U4577 = ~new_P1_R1240_U14 | ~new_P1_U3992;
  assign new_P1_U4578 = ~new_P1_U3398;
  assign new_P1_U4579 = ~new_P1_U3025 | ~new_P1_U3075;
  assign new_P1_U4580 = ~new_P1_R1222_U14 | ~new_P1_U3024;
  assign new_P1_U4581 = ~new_P1_R1282_U13 | ~new_P1_U4036;
  assign new_P1_U4582 = ~new_P1_U4025 | ~new_P1_U4185;
  assign new_P1_U4583 = ~new_P1_U3687 | ~new_P1_U4578;
  assign new_P1_U4584 = ~P1_REG2_REG_22_ | ~new_P1_U3018;
  assign new_P1_U4585 = ~P1_REG1_REG_22_ | ~new_P1_U3019;
  assign new_P1_U4586 = ~P1_REG0_REG_22_ | ~new_P1_U3020;
  assign new_P1_U4587 = ~new_P1_ADD_99_U66 | ~new_P1_U3017;
  assign new_P1_U4588 = ~new_P1_U3061;
  assign new_P1_U4589 = ~new_P1_U3034 | ~new_P1_U3076;
  assign new_P1_U4590 = ~new_P1_R1150_U111 | ~new_P1_U4007;
  assign new_P1_U4591 = ~new_P1_R1117_U111 | ~new_P1_U4000;
  assign new_P1_U4592 = ~new_P1_R1138_U15 | ~new_P1_U3994;
  assign new_P1_U4593 = ~new_P1_R1192_U111 | ~new_P1_U4005;
  assign new_P1_U4594 = ~new_P1_R1207_U111 | ~new_P1_U4004;
  assign new_P1_U4595 = ~new_P1_R1171_U15 | ~new_P1_U4011;
  assign new_P1_U4596 = ~new_P1_R1240_U15 | ~new_P1_U3992;
  assign new_P1_U4597 = ~new_P1_U3400;
  assign new_P1_U4598 = ~new_P1_U3025 | ~new_P1_U3061;
  assign new_P1_U4599 = ~new_P1_R1222_U15 | ~new_P1_U3024;
  assign new_P1_U4600 = ~new_P1_R1282_U78 | ~new_P1_U4036;
  assign new_P1_U4601 = ~new_P1_U4024 | ~new_P1_U4185;
  assign new_P1_U4602 = ~new_P1_U3691 | ~new_P1_U4597;
  assign new_P1_U4603 = ~P1_REG2_REG_23_ | ~new_P1_U3018;
  assign new_P1_U4604 = ~P1_REG1_REG_23_ | ~new_P1_U3019;
  assign new_P1_U4605 = ~P1_REG0_REG_23_ | ~new_P1_U3020;
  assign new_P1_U4606 = ~new_P1_ADD_99_U65 | ~new_P1_U3017;
  assign new_P1_U4607 = ~new_P1_U3066;
  assign new_P1_U4608 = ~new_P1_U3034 | ~new_P1_U3075;
  assign new_P1_U4609 = ~new_P1_R1150_U110 | ~new_P1_U4007;
  assign new_P1_U4610 = ~new_P1_R1117_U110 | ~new_P1_U4000;
  assign new_P1_U4611 = ~new_P1_R1138_U108 | ~new_P1_U3994;
  assign new_P1_U4612 = ~new_P1_R1192_U110 | ~new_P1_U4005;
  assign new_P1_U4613 = ~new_P1_R1207_U110 | ~new_P1_U4004;
  assign new_P1_U4614 = ~new_P1_R1171_U108 | ~new_P1_U4011;
  assign new_P1_U4615 = ~new_P1_R1240_U108 | ~new_P1_U3992;
  assign new_P1_U4616 = ~new_P1_U3402;
  assign new_P1_U4617 = ~new_P1_U3025 | ~new_P1_U3066;
  assign new_P1_U4618 = ~new_P1_R1222_U108 | ~new_P1_U3024;
  assign new_P1_U4619 = ~new_P1_R1282_U14 | ~new_P1_U4036;
  assign new_P1_U4620 = ~new_P1_U4023 | ~new_P1_U4185;
  assign new_P1_U4621 = ~new_P1_U3695 | ~new_P1_U4616;
  assign new_P1_U4622 = ~P1_REG2_REG_24_ | ~new_P1_U3018;
  assign new_P1_U4623 = ~P1_REG1_REG_24_ | ~new_P1_U3019;
  assign new_P1_U4624 = ~P1_REG0_REG_24_ | ~new_P1_U3020;
  assign new_P1_U4625 = ~new_P1_ADD_99_U64 | ~new_P1_U3017;
  assign new_P1_U4626 = ~new_P1_U3065;
  assign new_P1_U4627 = ~new_P1_U3034 | ~new_P1_U3061;
  assign new_P1_U4628 = ~new_P1_R1150_U15 | ~new_P1_U4007;
  assign new_P1_U4629 = ~new_P1_R1117_U15 | ~new_P1_U4000;
  assign new_P1_U4630 = ~new_P1_R1138_U107 | ~new_P1_U3994;
  assign new_P1_U4631 = ~new_P1_R1192_U15 | ~new_P1_U4005;
  assign new_P1_U4632 = ~new_P1_R1207_U15 | ~new_P1_U4004;
  assign new_P1_U4633 = ~new_P1_R1171_U107 | ~new_P1_U4011;
  assign new_P1_U4634 = ~new_P1_R1240_U107 | ~new_P1_U3992;
  assign new_P1_U4635 = ~new_P1_U3404;
  assign new_P1_U4636 = ~new_P1_U3025 | ~new_P1_U3065;
  assign new_P1_U4637 = ~new_P1_R1222_U107 | ~new_P1_U3024;
  assign new_P1_U4638 = ~new_P1_R1282_U76 | ~new_P1_U4036;
  assign new_P1_U4639 = ~new_P1_U4022 | ~new_P1_U4185;
  assign new_P1_U4640 = ~new_P1_U3699 | ~new_P1_U4635;
  assign new_P1_U4641 = ~P1_REG2_REG_25_ | ~new_P1_U3018;
  assign new_P1_U4642 = ~P1_REG1_REG_25_ | ~new_P1_U3019;
  assign new_P1_U4643 = ~P1_REG0_REG_25_ | ~new_P1_U3020;
  assign new_P1_U4644 = ~new_P1_ADD_99_U63 | ~new_P1_U3017;
  assign new_P1_U4645 = ~new_P1_U3058;
  assign new_P1_U4646 = ~new_P1_U3034 | ~new_P1_U3066;
  assign new_P1_U4647 = ~new_P1_R1150_U96 | ~new_P1_U4007;
  assign new_P1_U4648 = ~new_P1_R1117_U96 | ~new_P1_U4000;
  assign new_P1_U4649 = ~new_P1_R1138_U106 | ~new_P1_U3994;
  assign new_P1_U4650 = ~new_P1_R1192_U96 | ~new_P1_U4005;
  assign new_P1_U4651 = ~new_P1_R1207_U96 | ~new_P1_U4004;
  assign new_P1_U4652 = ~new_P1_R1171_U106 | ~new_P1_U4011;
  assign new_P1_U4653 = ~new_P1_R1240_U106 | ~new_P1_U3992;
  assign new_P1_U4654 = ~new_P1_U3406;
  assign new_P1_U4655 = ~new_P1_U3025 | ~new_P1_U3058;
  assign new_P1_U4656 = ~new_P1_R1222_U106 | ~new_P1_U3024;
  assign new_P1_U4657 = ~new_P1_R1282_U15 | ~new_P1_U4036;
  assign new_P1_U4658 = ~new_P1_U4021 | ~new_P1_U4185;
  assign new_P1_U4659 = ~new_P1_U3703 | ~new_P1_U4654;
  assign new_P1_U4660 = ~P1_REG2_REG_26_ | ~new_P1_U3018;
  assign new_P1_U4661 = ~P1_REG1_REG_26_ | ~new_P1_U3019;
  assign new_P1_U4662 = ~P1_REG0_REG_26_ | ~new_P1_U3020;
  assign new_P1_U4663 = ~new_P1_ADD_99_U62 | ~new_P1_U3017;
  assign new_P1_U4664 = ~new_P1_U3057;
  assign new_P1_U4665 = ~new_P1_U3034 | ~new_P1_U3065;
  assign new_P1_U4666 = ~new_P1_R1150_U95 | ~new_P1_U4007;
  assign new_P1_U4667 = ~new_P1_R1117_U95 | ~new_P1_U4000;
  assign new_P1_U4668 = ~new_P1_R1138_U105 | ~new_P1_U3994;
  assign new_P1_U4669 = ~new_P1_R1192_U95 | ~new_P1_U4005;
  assign new_P1_U4670 = ~new_P1_R1207_U95 | ~new_P1_U4004;
  assign new_P1_U4671 = ~new_P1_R1171_U105 | ~new_P1_U4011;
  assign new_P1_U4672 = ~new_P1_R1240_U105 | ~new_P1_U3992;
  assign new_P1_U4673 = ~new_P1_U3408;
  assign new_P1_U4674 = ~new_P1_U3025 | ~new_P1_U3057;
  assign new_P1_U4675 = ~new_P1_R1222_U105 | ~new_P1_U3024;
  assign new_P1_U4676 = ~new_P1_R1282_U74 | ~new_P1_U4036;
  assign new_P1_U4677 = ~new_P1_U4020 | ~new_P1_U4185;
  assign new_P1_U4678 = ~new_P1_U3707 | ~new_P1_U4673;
  assign new_P1_U4679 = ~P1_REG2_REG_27_ | ~new_P1_U3018;
  assign new_P1_U4680 = ~P1_REG1_REG_27_ | ~new_P1_U3019;
  assign new_P1_U4681 = ~P1_REG0_REG_27_ | ~new_P1_U3020;
  assign new_P1_U4682 = ~new_P1_ADD_99_U61 | ~new_P1_U3017;
  assign new_P1_U4683 = ~new_P1_U3053;
  assign new_P1_U4684 = ~new_P1_U3034 | ~new_P1_U3058;
  assign new_P1_U4685 = ~new_P1_R1150_U109 | ~new_P1_U4007;
  assign new_P1_U4686 = ~new_P1_R1117_U109 | ~new_P1_U4000;
  assign new_P1_U4687 = ~new_P1_R1138_U16 | ~new_P1_U3994;
  assign new_P1_U4688 = ~new_P1_R1192_U109 | ~new_P1_U4005;
  assign new_P1_U4689 = ~new_P1_R1207_U109 | ~new_P1_U4004;
  assign new_P1_U4690 = ~new_P1_R1171_U16 | ~new_P1_U4011;
  assign new_P1_U4691 = ~new_P1_R1240_U16 | ~new_P1_U3992;
  assign new_P1_U4692 = ~new_P1_U3410;
  assign new_P1_U4693 = ~new_P1_U3025 | ~new_P1_U3053;
  assign new_P1_U4694 = ~new_P1_R1222_U16 | ~new_P1_U3024;
  assign new_P1_U4695 = ~new_P1_R1282_U16 | ~new_P1_U4036;
  assign new_P1_U4696 = ~new_P1_U4019 | ~new_P1_U4185;
  assign new_P1_U4697 = ~new_P1_U3711 | ~new_P1_U4692;
  assign new_P1_U4698 = ~P1_REG2_REG_28_ | ~new_P1_U3018;
  assign new_P1_U4699 = ~P1_REG1_REG_28_ | ~new_P1_U3019;
  assign new_P1_U4700 = ~P1_REG0_REG_28_ | ~new_P1_U3020;
  assign new_P1_U4701 = ~new_P1_ADD_99_U60 | ~new_P1_U3017;
  assign new_P1_U4702 = ~new_P1_U3054;
  assign new_P1_U4703 = ~new_P1_U3034 | ~new_P1_U3057;
  assign new_P1_U4704 = ~new_P1_R1150_U16 | ~new_P1_U4007;
  assign new_P1_U4705 = ~new_P1_R1117_U16 | ~new_P1_U4000;
  assign new_P1_U4706 = ~new_P1_R1138_U104 | ~new_P1_U3994;
  assign new_P1_U4707 = ~new_P1_R1192_U16 | ~new_P1_U4005;
  assign new_P1_U4708 = ~new_P1_R1207_U16 | ~new_P1_U4004;
  assign new_P1_U4709 = ~new_P1_R1171_U104 | ~new_P1_U4011;
  assign new_P1_U4710 = ~new_P1_R1240_U104 | ~new_P1_U3992;
  assign new_P1_U4711 = ~new_P1_U3412;
  assign new_P1_U4712 = ~new_P1_U3025 | ~new_P1_U3054;
  assign new_P1_U4713 = ~new_P1_R1222_U104 | ~new_P1_U3024;
  assign new_P1_U4714 = ~new_P1_R1282_U72 | ~new_P1_U4036;
  assign new_P1_U4715 = ~new_P1_U4018 | ~new_P1_U4185;
  assign new_P1_U4716 = ~new_P1_U3715 | ~new_P1_U4711;
  assign new_P1_U4717 = ~new_P1_ADD_99_U5 | ~new_P1_U3017;
  assign new_P1_U4718 = ~P1_REG2_REG_29_ | ~new_P1_U3018;
  assign new_P1_U4719 = ~P1_REG1_REG_29_ | ~new_P1_U3019;
  assign new_P1_U4720 = ~P1_REG0_REG_29_ | ~new_P1_U3020;
  assign new_P1_U4721 = ~new_P1_U3055;
  assign new_P1_U4722 = ~new_P1_U3034 | ~new_P1_U3053;
  assign new_P1_U4723 = ~new_P1_R1150_U94 | ~new_P1_U4007;
  assign new_P1_U4724 = ~new_P1_R1117_U94 | ~new_P1_U4000;
  assign new_P1_U4725 = ~new_P1_R1138_U103 | ~new_P1_U3994;
  assign new_P1_U4726 = ~new_P1_R1192_U94 | ~new_P1_U4005;
  assign new_P1_U4727 = ~new_P1_R1207_U94 | ~new_P1_U4004;
  assign new_P1_U4728 = ~new_P1_R1171_U103 | ~new_P1_U4011;
  assign new_P1_U4729 = ~new_P1_R1240_U103 | ~new_P1_U3992;
  assign new_P1_U4730 = ~new_P1_U3414;
  assign new_P1_U4731 = ~new_P1_U3025 | ~new_P1_U3055;
  assign new_P1_U4732 = ~new_P1_R1222_U103 | ~new_P1_U3024;
  assign new_P1_U4733 = ~new_P1_R1282_U17 | ~new_P1_U4036;
  assign new_P1_U4734 = ~new_P1_U4017 | ~new_P1_U4185;
  assign new_P1_U4735 = ~new_P1_U3719 | ~new_P1_U4730;
  assign new_P1_U4736 = ~P1_REG2_REG_30_ | ~new_P1_U3018;
  assign new_P1_U4737 = ~P1_REG1_REG_30_ | ~new_P1_U3019;
  assign new_P1_U4738 = ~P1_REG0_REG_30_ | ~new_P1_U3020;
  assign new_P1_U4739 = ~new_P1_U3059;
  assign new_P1_U4740 = ~new_P1_U5811 | ~new_P1_U3359;
  assign new_P1_U4741 = ~new_P1_U3954 | ~new_P1_U4740;
  assign new_P1_U4742 = ~new_P1_U3720 | ~new_P1_U3059;
  assign new_P1_U4743 = ~new_P1_U3034 | ~new_P1_U3054;
  assign new_P1_U4744 = ~new_P1_R1150_U17 | ~new_P1_U4007;
  assign new_P1_U4745 = ~new_P1_R1117_U17 | ~new_P1_U4000;
  assign new_P1_U4746 = ~new_P1_R1138_U102 | ~new_P1_U3994;
  assign new_P1_U4747 = ~new_P1_R1192_U17 | ~new_P1_U4005;
  assign new_P1_U4748 = ~new_P1_R1207_U17 | ~new_P1_U4004;
  assign new_P1_U4749 = ~new_P1_R1171_U102 | ~new_P1_U4011;
  assign new_P1_U4750 = ~new_P1_R1240_U102 | ~new_P1_U3992;
  assign new_P1_U4751 = ~new_P1_U3416;
  assign new_P1_U4752 = ~new_P1_R1222_U102 | ~new_P1_U3024;
  assign new_P1_U4753 = ~new_P1_R1282_U70 | ~new_P1_U4036;
  assign new_P1_U4754 = ~new_P1_U4028 | ~new_P1_U4185;
  assign new_P1_U4755 = ~new_P1_U3724 | ~new_P1_U4751;
  assign new_P1_U4756 = ~P1_REG2_REG_31_ | ~new_P1_U3018;
  assign new_P1_U4757 = ~P1_REG1_REG_31_ | ~new_P1_U3019;
  assign new_P1_U4758 = ~P1_REG0_REG_31_ | ~new_P1_U3020;
  assign new_P1_U4759 = ~new_P1_U3056;
  assign new_P1_U4760 = ~new_P1_R1282_U19 | ~new_P1_U4036;
  assign new_P1_U4761 = ~new_P1_U4027 | ~new_P1_U4185;
  assign new_P1_U4762 = ~new_P1_U4760 | ~new_P1_U4761 | ~new_P1_U3987;
  assign new_P1_U4763 = ~new_P1_R1282_U68 | ~new_P1_U4036;
  assign new_P1_U4764 = ~new_P1_U4026 | ~new_P1_U4185;
  assign new_P1_U4765 = ~new_P1_U4763 | ~new_P1_U4764 | ~new_P1_U3987;
  assign new_P1_U4766 = ~new_P1_U3727 | ~new_P1_U3016;
  assign new_P1_U4767 = ~new_P1_U3421 | ~new_P1_U4766;
  assign new_P1_U4768 = ~new_P1_U3995 | ~new_P1_U5802;
  assign new_P1_U4769 = ~new_P1_U3426;
  assign new_P1_U4770 = ~new_P1_U3036 | ~new_P1_U3078;
  assign new_P1_U4771 = ~new_P1_U3033 | ~P1_REG3_REG_0_;
  assign new_P1_U4772 = ~new_P1_U3032 | ~new_P1_R1222_U96;
  assign new_P1_U4773 = ~new_P1_U3031 | ~new_P1_U3456;
  assign new_P1_U4774 = ~new_P1_U3030 | ~new_P1_U3456;
  assign new_P1_U4775 = ~new_P1_U3036 | ~new_P1_U3068;
  assign new_P1_U4776 = ~new_P1_U3033 | ~P1_REG3_REG_1_;
  assign new_P1_U4777 = ~new_P1_U3032 | ~new_P1_R1222_U95;
  assign new_P1_U4778 = ~new_P1_U3031 | ~new_P1_U3461;
  assign new_P1_U4779 = ~new_P1_U3030 | ~new_P1_R1282_U56;
  assign new_P1_U4780 = ~new_P1_U3036 | ~new_P1_U3064;
  assign new_P1_U4781 = ~new_P1_U3033 | ~P1_REG3_REG_2_;
  assign new_P1_U4782 = ~new_P1_U3032 | ~new_P1_R1222_U17;
  assign new_P1_U4783 = ~new_P1_U3031 | ~new_P1_U3464;
  assign new_P1_U4784 = ~new_P1_U3030 | ~new_P1_R1282_U18;
  assign new_P1_U4785 = ~new_P1_U3036 | ~new_P1_U3060;
  assign new_P1_U4786 = ~new_P1_U3033 | ~new_P1_ADD_99_U4;
  assign new_P1_U4787 = ~new_P1_U3032 | ~new_P1_R1222_U101;
  assign new_P1_U4788 = ~new_P1_U3031 | ~new_P1_U3467;
  assign new_P1_U4789 = ~new_P1_U3030 | ~new_P1_R1282_U20;
  assign new_P1_U4790 = ~new_P1_U3036 | ~new_P1_U3067;
  assign new_P1_U4791 = ~new_P1_U3033 | ~new_P1_ADD_99_U59;
  assign new_P1_U4792 = ~new_P1_U3032 | ~new_P1_R1222_U100;
  assign new_P1_U4793 = ~new_P1_U3031 | ~new_P1_U3470;
  assign new_P1_U4794 = ~new_P1_U3030 | ~new_P1_R1282_U21;
  assign new_P1_U4795 = ~new_P1_U3036 | ~new_P1_U3071;
  assign new_P1_U4796 = ~new_P1_U3033 | ~new_P1_ADD_99_U58;
  assign new_P1_U4797 = ~new_P1_U3032 | ~new_P1_R1222_U18;
  assign new_P1_U4798 = ~new_P1_U3031 | ~new_P1_U3473;
  assign new_P1_U4799 = ~new_P1_U3030 | ~new_P1_R1282_U65;
  assign new_P1_U4800 = ~new_P1_U3036 | ~new_P1_U3070;
  assign new_P1_U4801 = ~new_P1_U3033 | ~new_P1_ADD_99_U57;
  assign new_P1_U4802 = ~new_P1_U3032 | ~new_P1_R1222_U99;
  assign new_P1_U4803 = ~new_P1_U3031 | ~new_P1_U3476;
  assign new_P1_U4804 = ~new_P1_U3030 | ~new_P1_R1282_U22;
  assign new_P1_U4805 = ~new_P1_U3036 | ~new_P1_U3084;
  assign new_P1_U4806 = ~new_P1_U3033 | ~new_P1_ADD_99_U56;
  assign new_P1_U4807 = ~new_P1_U3032 | ~new_P1_R1222_U19;
  assign new_P1_U4808 = ~new_P1_U3031 | ~new_P1_U3479;
  assign new_P1_U4809 = ~new_P1_U3030 | ~new_P1_R1282_U23;
  assign new_P1_U4810 = ~new_P1_U3036 | ~new_P1_U3083;
  assign new_P1_U4811 = ~new_P1_U3033 | ~new_P1_ADD_99_U55;
  assign new_P1_U4812 = ~new_P1_U3032 | ~new_P1_R1222_U98;
  assign new_P1_U4813 = ~new_P1_U3031 | ~new_P1_U3482;
  assign new_P1_U4814 = ~new_P1_U3030 | ~new_P1_R1282_U24;
  assign new_P1_U4815 = ~new_P1_U3036 | ~new_P1_U3062;
  assign new_P1_U4816 = ~new_P1_U3033 | ~new_P1_ADD_99_U54;
  assign new_P1_U4817 = ~new_P1_U3032 | ~new_P1_R1222_U97;
  assign new_P1_U4818 = ~new_P1_U3031 | ~new_P1_U3485;
  assign new_P1_U4819 = ~new_P1_U3030 | ~new_P1_R1282_U63;
  assign new_P1_U4820 = ~new_P1_U3036 | ~new_P1_U3063;
  assign new_P1_U4821 = ~new_P1_U3033 | ~new_P1_ADD_99_U78;
  assign new_P1_U4822 = ~new_P1_U3032 | ~new_P1_R1222_U11;
  assign new_P1_U4823 = ~new_P1_U3031 | ~new_P1_U3488;
  assign new_P1_U4824 = ~new_P1_U3030 | ~new_P1_R1282_U6;
  assign new_P1_U4825 = ~new_P1_U3036 | ~new_P1_U3072;
  assign new_P1_U4826 = ~new_P1_U3033 | ~new_P1_ADD_99_U77;
  assign new_P1_U4827 = ~new_P1_U3032 | ~new_P1_R1222_U115;
  assign new_P1_U4828 = ~new_P1_U3031 | ~new_P1_U3491;
  assign new_P1_U4829 = ~new_P1_U3030 | ~new_P1_R1282_U7;
  assign new_P1_U4830 = ~new_P1_U3036 | ~new_P1_U3080;
  assign new_P1_U4831 = ~new_P1_U3033 | ~new_P1_ADD_99_U76;
  assign new_P1_U4832 = ~new_P1_U3032 | ~new_P1_R1222_U114;
  assign new_P1_U4833 = ~new_P1_U3031 | ~new_P1_U3494;
  assign new_P1_U4834 = ~new_P1_U3030 | ~new_P1_R1282_U8;
  assign new_P1_U4835 = ~new_P1_U3036 | ~new_P1_U3079;
  assign new_P1_U4836 = ~new_P1_U3033 | ~new_P1_ADD_99_U75;
  assign new_P1_U4837 = ~new_P1_U3032 | ~new_P1_R1222_U12;
  assign new_P1_U4838 = ~new_P1_U3031 | ~new_P1_U3497;
  assign new_P1_U4839 = ~new_P1_U3030 | ~new_P1_R1282_U86;
  assign new_P1_U4840 = ~new_P1_U3036 | ~new_P1_U3074;
  assign new_P1_U4841 = ~new_P1_U3033 | ~new_P1_ADD_99_U74;
  assign new_P1_U4842 = ~new_P1_U3032 | ~new_P1_R1222_U113;
  assign new_P1_U4843 = ~new_P1_U3031 | ~new_P1_U3500;
  assign new_P1_U4844 = ~new_P1_U3030 | ~new_P1_R1282_U9;
  assign new_P1_U4845 = ~new_P1_U3036 | ~new_P1_U3073;
  assign new_P1_U4846 = ~new_P1_U3033 | ~new_P1_ADD_99_U73;
  assign new_P1_U4847 = ~new_P1_U3032 | ~new_P1_R1222_U112;
  assign new_P1_U4848 = ~new_P1_U3031 | ~new_P1_U3503;
  assign new_P1_U4849 = ~new_P1_U3030 | ~new_P1_R1282_U10;
  assign new_P1_U4850 = ~new_P1_U3036 | ~new_P1_U3069;
  assign new_P1_U4851 = ~new_P1_U3033 | ~new_P1_ADD_99_U72;
  assign new_P1_U4852 = ~new_P1_U3032 | ~new_P1_R1222_U111;
  assign new_P1_U4853 = ~new_P1_U3031 | ~new_P1_U3506;
  assign new_P1_U4854 = ~new_P1_U3030 | ~new_P1_R1282_U11;
  assign new_P1_U4855 = ~new_P1_U3036 | ~new_P1_U3082;
  assign new_P1_U4856 = ~new_P1_U3033 | ~new_P1_ADD_99_U71;
  assign new_P1_U4857 = ~new_P1_U3032 | ~new_P1_R1222_U13;
  assign new_P1_U4858 = ~new_P1_U3031 | ~new_P1_U3509;
  assign new_P1_U4859 = ~new_P1_U3030 | ~new_P1_R1282_U84;
  assign new_P1_U4860 = ~new_P1_U3036 | ~new_P1_U3081;
  assign new_P1_U4861 = ~new_P1_U3033 | ~new_P1_ADD_99_U70;
  assign new_P1_U4862 = ~new_P1_U3032 | ~new_P1_R1222_U110;
  assign new_P1_U4863 = ~new_P1_U3031 | ~new_P1_U3512;
  assign new_P1_U4864 = ~new_P1_U3030 | ~new_P1_R1282_U12;
  assign new_P1_U4865 = ~new_P1_U3036 | ~new_P1_U3076;
  assign new_P1_U4866 = ~new_P1_U3033 | ~new_P1_ADD_99_U69;
  assign new_P1_U4867 = ~new_P1_U3032 | ~new_P1_R1222_U109;
  assign new_P1_U4868 = ~new_P1_U3031 | ~new_P1_U3514;
  assign new_P1_U4869 = ~new_P1_U3030 | ~new_P1_R1282_U82;
  assign new_P1_U4870 = ~new_P1_U3036 | ~new_P1_U3075;
  assign new_P1_U4871 = ~new_P1_U3033 | ~new_P1_ADD_99_U68;
  assign new_P1_U4872 = ~new_P1_U3032 | ~new_P1_R1222_U14;
  assign new_P1_U4873 = ~new_P1_U3031 | ~new_P1_U4025;
  assign new_P1_U4874 = ~new_P1_U3030 | ~new_P1_R1282_U13;
  assign new_P1_U4875 = ~new_P1_U3036 | ~new_P1_U3061;
  assign new_P1_U4876 = ~new_P1_U3033 | ~new_P1_ADD_99_U67;
  assign new_P1_U4877 = ~new_P1_U3032 | ~new_P1_R1222_U15;
  assign new_P1_U4878 = ~new_P1_U3031 | ~new_P1_U4024;
  assign new_P1_U4879 = ~new_P1_U3030 | ~new_P1_R1282_U78;
  assign new_P1_U4880 = ~new_P1_U3036 | ~new_P1_U3066;
  assign new_P1_U4881 = ~new_P1_U3033 | ~new_P1_ADD_99_U66;
  assign new_P1_U4882 = ~new_P1_U3032 | ~new_P1_R1222_U108;
  assign new_P1_U4883 = ~new_P1_U3031 | ~new_P1_U4023;
  assign new_P1_U4884 = ~new_P1_U3030 | ~new_P1_R1282_U14;
  assign new_P1_U4885 = ~new_P1_U3036 | ~new_P1_U3065;
  assign new_P1_U4886 = ~new_P1_U3033 | ~new_P1_ADD_99_U65;
  assign new_P1_U4887 = ~new_P1_U3032 | ~new_P1_R1222_U107;
  assign new_P1_U4888 = ~new_P1_U3031 | ~new_P1_U4022;
  assign new_P1_U4889 = ~new_P1_U3030 | ~new_P1_R1282_U76;
  assign new_P1_U4890 = ~new_P1_U3036 | ~new_P1_U3058;
  assign new_P1_U4891 = ~new_P1_U3033 | ~new_P1_ADD_99_U64;
  assign new_P1_U4892 = ~new_P1_U3032 | ~new_P1_R1222_U106;
  assign new_P1_U4893 = ~new_P1_U3031 | ~new_P1_U4021;
  assign new_P1_U4894 = ~new_P1_U3030 | ~new_P1_R1282_U15;
  assign new_P1_U4895 = ~new_P1_U3036 | ~new_P1_U3057;
  assign new_P1_U4896 = ~new_P1_U3033 | ~new_P1_ADD_99_U63;
  assign new_P1_U4897 = ~new_P1_U3032 | ~new_P1_R1222_U105;
  assign new_P1_U4898 = ~new_P1_U3031 | ~new_P1_U4020;
  assign new_P1_U4899 = ~new_P1_U3030 | ~new_P1_R1282_U74;
  assign new_P1_U4900 = ~new_P1_U3036 | ~new_P1_U3053;
  assign new_P1_U4901 = ~new_P1_U3033 | ~new_P1_ADD_99_U62;
  assign new_P1_U4902 = ~new_P1_U3032 | ~new_P1_R1222_U16;
  assign new_P1_U4903 = ~new_P1_U3031 | ~new_P1_U4019;
  assign new_P1_U4904 = ~new_P1_U3030 | ~new_P1_R1282_U16;
  assign new_P1_U4905 = ~new_P1_U3036 | ~new_P1_U3054;
  assign new_P1_U4906 = ~new_P1_U3033 | ~new_P1_ADD_99_U61;
  assign new_P1_U4907 = ~new_P1_U3032 | ~new_P1_R1222_U104;
  assign new_P1_U4908 = ~new_P1_U3031 | ~new_P1_U4018;
  assign new_P1_U4909 = ~new_P1_U3030 | ~new_P1_R1282_U72;
  assign new_P1_U4910 = ~new_P1_U3036 | ~new_P1_U3055;
  assign new_P1_U4911 = ~new_P1_U3033 | ~new_P1_ADD_99_U60;
  assign new_P1_U4912 = ~new_P1_U3032 | ~new_P1_R1222_U103;
  assign new_P1_U4913 = ~new_P1_U3031 | ~new_P1_U4017;
  assign new_P1_U4914 = ~new_P1_U3030 | ~new_P1_R1282_U17;
  assign new_P1_U4915 = ~new_P1_U3033 | ~new_P1_ADD_99_U5;
  assign new_P1_U4916 = ~new_P1_U3032 | ~new_P1_R1222_U102;
  assign new_P1_U4917 = ~new_P1_U3031 | ~new_P1_U4028;
  assign new_P1_U4918 = ~new_P1_U3030 | ~new_P1_R1282_U70;
  assign new_P1_U4919 = ~new_P1_U3031 | ~new_P1_U4027;
  assign new_P1_U4920 = ~new_P1_U3030 | ~new_P1_R1282_U19;
  assign new_P1_U4921 = ~new_P1_U3031 | ~new_P1_U4026;
  assign new_P1_U4922 = ~new_P1_U3030 | ~new_P1_R1282_U68;
  assign new_P1_U4923 = ~new_P1_U3421 | ~new_P1_U4769 | ~new_P1_U3789 | ~new_P1_U3787 | ~new_P1_U3786;
  assign new_P1_U4924 = ~new_P1_R1105_U13 | ~new_P1_U3042;
  assign new_P1_U4925 = ~new_P1_U3040 | ~new_P1_U3452;
  assign new_P1_U4926 = ~new_P1_R1162_U13 | ~new_P1_U3038;
  assign new_P1_U4927 = ~new_P1_U4926 | ~new_P1_U4925 | ~new_P1_U4924;
  assign new_P1_U4928 = ~new_P1_U3425 | ~new_P1_U3372;
  assign new_P1_U4929 = ~new_P1_U5786 | ~new_P1_U4928;
  assign new_P1_U4930 = ~new_P1_U4929 | ~new_P1_U3954;
  assign new_P1_U4931 = ~n1389;
  assign new_P1_U4932 = ~new_P1_U3428;
  assign new_P1_U4933 = ~new_P1_U3044 | ~new_P1_U4927;
  assign new_P1_U4934 = ~new_P1_U3043 | ~new_P1_R1105_U13;
  assign new_P1_U4935 = ~P1_REG3_REG_19_ | ~n1384;
  assign new_P1_U4936 = ~new_P1_U3041 | ~new_P1_U3452;
  assign new_P1_U4937 = ~new_P1_U3039 | ~new_P1_R1162_U13;
  assign new_P1_U4938 = ~P1_ADDR_REG_19_ | ~new_P1_U4932;
  assign new_P1_U4939 = ~new_P1_R1105_U75 | ~new_P1_U3042;
  assign new_P1_U4940 = ~new_P1_U3040 | ~new_P1_U3511;
  assign new_P1_U4941 = ~new_P1_R1162_U75 | ~new_P1_U3038;
  assign new_P1_U4942 = ~new_P1_U4941 | ~new_P1_U4940 | ~new_P1_U4939;
  assign new_P1_U4943 = ~new_P1_U3044 | ~new_P1_U4942;
  assign new_P1_U4944 = ~new_P1_R1105_U75 | ~new_P1_U3043;
  assign new_P1_U4945 = ~P1_REG3_REG_18_ | ~n1384;
  assign new_P1_U4946 = ~new_P1_U3041 | ~new_P1_U3511;
  assign new_P1_U4947 = ~new_P1_R1162_U75 | ~new_P1_U3039;
  assign new_P1_U4948 = ~P1_ADDR_REG_18_ | ~new_P1_U4932;
  assign new_P1_U4949 = ~new_P1_R1105_U12 | ~new_P1_U3042;
  assign new_P1_U4950 = ~new_P1_U3040 | ~new_P1_U3508;
  assign new_P1_U4951 = ~new_P1_R1162_U12 | ~new_P1_U3038;
  assign new_P1_U4952 = ~new_P1_U4951 | ~new_P1_U4950 | ~new_P1_U4949;
  assign new_P1_U4953 = ~new_P1_U3044 | ~new_P1_U4952;
  assign new_P1_U4954 = ~new_P1_R1105_U12 | ~new_P1_U3043;
  assign new_P1_U4955 = ~P1_REG3_REG_17_ | ~n1384;
  assign new_P1_U4956 = ~new_P1_U3041 | ~new_P1_U3508;
  assign new_P1_U4957 = ~new_P1_R1162_U12 | ~new_P1_U3039;
  assign new_P1_U4958 = ~P1_ADDR_REG_17_ | ~new_P1_U4932;
  assign new_P1_U4959 = ~new_P1_R1105_U76 | ~new_P1_U3042;
  assign new_P1_U4960 = ~new_P1_U3040 | ~new_P1_U3505;
  assign new_P1_U4961 = ~new_P1_R1162_U76 | ~new_P1_U3038;
  assign new_P1_U4962 = ~new_P1_U4961 | ~new_P1_U4960 | ~new_P1_U4959;
  assign new_P1_U4963 = ~new_P1_U3044 | ~new_P1_U4962;
  assign new_P1_U4964 = ~new_P1_R1105_U76 | ~new_P1_U3043;
  assign new_P1_U4965 = ~P1_REG3_REG_16_ | ~n1384;
  assign new_P1_U4966 = ~new_P1_U3041 | ~new_P1_U3505;
  assign new_P1_U4967 = ~new_P1_R1162_U76 | ~new_P1_U3039;
  assign new_P1_U4968 = ~P1_ADDR_REG_16_ | ~new_P1_U4932;
  assign new_P1_U4969 = ~new_P1_R1105_U77 | ~new_P1_U3042;
  assign new_P1_U4970 = ~new_P1_U3040 | ~new_P1_U3502;
  assign new_P1_U4971 = ~new_P1_R1162_U77 | ~new_P1_U3038;
  assign new_P1_U4972 = ~new_P1_U4971 | ~new_P1_U4970 | ~new_P1_U4969;
  assign new_P1_U4973 = ~new_P1_U3044 | ~new_P1_U4972;
  assign new_P1_U4974 = ~new_P1_R1105_U77 | ~new_P1_U3043;
  assign new_P1_U4975 = ~P1_REG3_REG_15_ | ~n1384;
  assign new_P1_U4976 = ~new_P1_U3041 | ~new_P1_U3502;
  assign new_P1_U4977 = ~new_P1_R1162_U77 | ~new_P1_U3039;
  assign new_P1_U4978 = ~P1_ADDR_REG_15_ | ~new_P1_U4932;
  assign new_P1_U4979 = ~new_P1_R1105_U78 | ~new_P1_U3042;
  assign new_P1_U4980 = ~new_P1_U3040 | ~new_P1_U3499;
  assign new_P1_U4981 = ~new_P1_R1162_U78 | ~new_P1_U3038;
  assign new_P1_U4982 = ~new_P1_U4981 | ~new_P1_U4980 | ~new_P1_U4979;
  assign new_P1_U4983 = ~new_P1_U3044 | ~new_P1_U4982;
  assign new_P1_U4984 = ~new_P1_R1105_U78 | ~new_P1_U3043;
  assign new_P1_U4985 = ~P1_REG3_REG_14_ | ~n1384;
  assign new_P1_U4986 = ~new_P1_U3041 | ~new_P1_U3499;
  assign new_P1_U4987 = ~new_P1_R1162_U78 | ~new_P1_U3039;
  assign new_P1_U4988 = ~P1_ADDR_REG_14_ | ~new_P1_U4932;
  assign new_P1_U4989 = ~new_P1_R1105_U11 | ~new_P1_U3042;
  assign new_P1_U4990 = ~new_P1_U3040 | ~new_P1_U3496;
  assign new_P1_U4991 = ~new_P1_R1162_U11 | ~new_P1_U3038;
  assign new_P1_U4992 = ~new_P1_U4991 | ~new_P1_U4990 | ~new_P1_U4989;
  assign new_P1_U4993 = ~new_P1_U3044 | ~new_P1_U4992;
  assign new_P1_U4994 = ~new_P1_R1105_U11 | ~new_P1_U3043;
  assign new_P1_U4995 = ~P1_REG3_REG_13_ | ~n1384;
  assign new_P1_U4996 = ~new_P1_U3041 | ~new_P1_U3496;
  assign new_P1_U4997 = ~new_P1_R1162_U11 | ~new_P1_U3039;
  assign new_P1_U4998 = ~P1_ADDR_REG_13_ | ~new_P1_U4932;
  assign new_P1_U4999 = ~new_P1_R1105_U79 | ~new_P1_U3042;
  assign new_P1_U5000 = ~new_P1_U3040 | ~new_P1_U3493;
  assign new_P1_U5001 = ~new_P1_R1162_U79 | ~new_P1_U3038;
  assign new_P1_U5002 = ~new_P1_U5001 | ~new_P1_U5000 | ~new_P1_U4999;
  assign new_P1_U5003 = ~new_P1_U3044 | ~new_P1_U5002;
  assign new_P1_U5004 = ~new_P1_R1105_U79 | ~new_P1_U3043;
  assign new_P1_U5005 = ~P1_REG3_REG_12_ | ~n1384;
  assign new_P1_U5006 = ~new_P1_U3041 | ~new_P1_U3493;
  assign new_P1_U5007 = ~new_P1_R1162_U79 | ~new_P1_U3039;
  assign new_P1_U5008 = ~P1_ADDR_REG_12_ | ~new_P1_U4932;
  assign new_P1_U5009 = ~new_P1_R1105_U80 | ~new_P1_U3042;
  assign new_P1_U5010 = ~new_P1_U3040 | ~new_P1_U3490;
  assign new_P1_U5011 = ~new_P1_R1162_U80 | ~new_P1_U3038;
  assign new_P1_U5012 = ~new_P1_U5011 | ~new_P1_U5010 | ~new_P1_U5009;
  assign new_P1_U5013 = ~new_P1_U3044 | ~new_P1_U5012;
  assign new_P1_U5014 = ~new_P1_R1105_U80 | ~new_P1_U3043;
  assign new_P1_U5015 = ~P1_REG3_REG_11_ | ~n1384;
  assign new_P1_U5016 = ~new_P1_U3041 | ~new_P1_U3490;
  assign new_P1_U5017 = ~new_P1_R1162_U80 | ~new_P1_U3039;
  assign new_P1_U5018 = ~P1_ADDR_REG_11_ | ~new_P1_U4932;
  assign new_P1_U5019 = ~new_P1_R1105_U10 | ~new_P1_U3042;
  assign new_P1_U5020 = ~new_P1_U3040 | ~new_P1_U3487;
  assign new_P1_U5021 = ~new_P1_R1162_U10 | ~new_P1_U3038;
  assign new_P1_U5022 = ~new_P1_U5021 | ~new_P1_U5020 | ~new_P1_U5019;
  assign new_P1_U5023 = ~new_P1_U3044 | ~new_P1_U5022;
  assign new_P1_U5024 = ~new_P1_R1105_U10 | ~new_P1_U3043;
  assign new_P1_U5025 = ~P1_REG3_REG_10_ | ~n1384;
  assign new_P1_U5026 = ~new_P1_U3041 | ~new_P1_U3487;
  assign new_P1_U5027 = ~new_P1_R1162_U10 | ~new_P1_U3039;
  assign new_P1_U5028 = ~P1_ADDR_REG_10_ | ~new_P1_U4932;
  assign new_P1_U5029 = ~new_P1_R1105_U70 | ~new_P1_U3042;
  assign new_P1_U5030 = ~new_P1_U3040 | ~new_P1_U3484;
  assign new_P1_U5031 = ~new_P1_R1162_U70 | ~new_P1_U3038;
  assign new_P1_U5032 = ~new_P1_U5031 | ~new_P1_U5030 | ~new_P1_U5029;
  assign new_P1_U5033 = ~new_P1_U3044 | ~new_P1_U5032;
  assign new_P1_U5034 = ~new_P1_R1105_U70 | ~new_P1_U3043;
  assign new_P1_U5035 = ~P1_REG3_REG_9_ | ~n1384;
  assign new_P1_U5036 = ~new_P1_U3041 | ~new_P1_U3484;
  assign new_P1_U5037 = ~new_P1_R1162_U70 | ~new_P1_U3039;
  assign new_P1_U5038 = ~P1_ADDR_REG_9_ | ~new_P1_U4932;
  assign new_P1_U5039 = ~new_P1_R1105_U71 | ~new_P1_U3042;
  assign new_P1_U5040 = ~new_P1_U3040 | ~new_P1_U3481;
  assign new_P1_U5041 = ~new_P1_R1162_U71 | ~new_P1_U3038;
  assign new_P1_U5042 = ~new_P1_U5041 | ~new_P1_U5040 | ~new_P1_U5039;
  assign new_P1_U5043 = ~new_P1_U3044 | ~new_P1_U5042;
  assign new_P1_U5044 = ~new_P1_R1105_U71 | ~new_P1_U3043;
  assign new_P1_U5045 = ~P1_REG3_REG_8_ | ~n1384;
  assign new_P1_U5046 = ~new_P1_U3041 | ~new_P1_U3481;
  assign new_P1_U5047 = ~new_P1_R1162_U71 | ~new_P1_U3039;
  assign new_P1_U5048 = ~P1_ADDR_REG_8_ | ~new_P1_U4932;
  assign new_P1_U5049 = ~new_P1_R1105_U16 | ~new_P1_U3042;
  assign new_P1_U5050 = ~new_P1_U3040 | ~new_P1_U3478;
  assign new_P1_U5051 = ~new_P1_R1162_U16 | ~new_P1_U3038;
  assign new_P1_U5052 = ~new_P1_U5051 | ~new_P1_U5050 | ~new_P1_U5049;
  assign new_P1_U5053 = ~new_P1_U3044 | ~new_P1_U5052;
  assign new_P1_U5054 = ~new_P1_R1105_U16 | ~new_P1_U3043;
  assign new_P1_U5055 = ~P1_REG3_REG_7_ | ~n1384;
  assign new_P1_U5056 = ~new_P1_U3041 | ~new_P1_U3478;
  assign new_P1_U5057 = ~new_P1_R1162_U16 | ~new_P1_U3039;
  assign new_P1_U5058 = ~P1_ADDR_REG_7_ | ~new_P1_U4932;
  assign new_P1_U5059 = ~new_P1_R1105_U72 | ~new_P1_U3042;
  assign new_P1_U5060 = ~new_P1_U3040 | ~new_P1_U3475;
  assign new_P1_U5061 = ~new_P1_R1162_U72 | ~new_P1_U3038;
  assign new_P1_U5062 = ~new_P1_U5061 | ~new_P1_U5060 | ~new_P1_U5059;
  assign new_P1_U5063 = ~new_P1_U3044 | ~new_P1_U5062;
  assign new_P1_U5064 = ~new_P1_R1105_U72 | ~new_P1_U3043;
  assign new_P1_U5065 = ~P1_REG3_REG_6_ | ~n1384;
  assign new_P1_U5066 = ~new_P1_U3041 | ~new_P1_U3475;
  assign new_P1_U5067 = ~new_P1_R1162_U72 | ~new_P1_U3039;
  assign new_P1_U5068 = ~P1_ADDR_REG_6_ | ~new_P1_U4932;
  assign new_P1_U5069 = ~new_P1_R1105_U15 | ~new_P1_U3042;
  assign new_P1_U5070 = ~new_P1_U3040 | ~new_P1_U3472;
  assign new_P1_U5071 = ~new_P1_R1162_U15 | ~new_P1_U3038;
  assign new_P1_U5072 = ~new_P1_U5071 | ~new_P1_U5070 | ~new_P1_U5069;
  assign new_P1_U5073 = ~new_P1_U3044 | ~new_P1_U5072;
  assign new_P1_U5074 = ~new_P1_R1105_U15 | ~new_P1_U3043;
  assign new_P1_U5075 = ~P1_REG3_REG_5_ | ~n1384;
  assign new_P1_U5076 = ~new_P1_U3041 | ~new_P1_U3472;
  assign new_P1_U5077 = ~new_P1_R1162_U15 | ~new_P1_U3039;
  assign new_P1_U5078 = ~P1_ADDR_REG_5_ | ~new_P1_U4932;
  assign new_P1_U5079 = ~new_P1_R1105_U73 | ~new_P1_U3042;
  assign new_P1_U5080 = ~new_P1_U3040 | ~new_P1_U3469;
  assign new_P1_U5081 = ~new_P1_R1162_U73 | ~new_P1_U3038;
  assign new_P1_U5082 = ~new_P1_U5081 | ~new_P1_U5080 | ~new_P1_U5079;
  assign new_P1_U5083 = ~new_P1_U3044 | ~new_P1_U5082;
  assign new_P1_U5084 = ~new_P1_R1105_U73 | ~new_P1_U3043;
  assign new_P1_U5085 = ~P1_REG3_REG_4_ | ~n1384;
  assign new_P1_U5086 = ~new_P1_U3041 | ~new_P1_U3469;
  assign new_P1_U5087 = ~new_P1_R1162_U73 | ~new_P1_U3039;
  assign new_P1_U5088 = ~P1_ADDR_REG_4_ | ~new_P1_U4932;
  assign new_P1_U5089 = ~new_P1_R1105_U74 | ~new_P1_U3042;
  assign new_P1_U5090 = ~new_P1_U3040 | ~new_P1_U3466;
  assign new_P1_U5091 = ~new_P1_R1162_U74 | ~new_P1_U3038;
  assign new_P1_U5092 = ~new_P1_U5091 | ~new_P1_U5090 | ~new_P1_U5089;
  assign new_P1_U5093 = ~new_P1_U3044 | ~new_P1_U5092;
  assign new_P1_U5094 = ~new_P1_R1105_U74 | ~new_P1_U3043;
  assign new_P1_U5095 = ~P1_REG3_REG_3_ | ~n1384;
  assign new_P1_U5096 = ~new_P1_U3041 | ~new_P1_U3466;
  assign new_P1_U5097 = ~new_P1_R1162_U74 | ~new_P1_U3039;
  assign new_P1_U5098 = ~P1_ADDR_REG_3_ | ~new_P1_U4932;
  assign new_P1_U5099 = ~new_P1_R1105_U14 | ~new_P1_U3042;
  assign new_P1_U5100 = ~new_P1_U3040 | ~new_P1_U3463;
  assign new_P1_U5101 = ~new_P1_R1162_U14 | ~new_P1_U3038;
  assign new_P1_U5102 = ~new_P1_U5101 | ~new_P1_U5100 | ~new_P1_U5099;
  assign new_P1_U5103 = ~new_P1_U3044 | ~new_P1_U5102;
  assign new_P1_U5104 = ~new_P1_R1105_U14 | ~new_P1_U3043;
  assign new_P1_U5105 = ~P1_REG3_REG_2_ | ~n1384;
  assign new_P1_U5106 = ~new_P1_U3041 | ~new_P1_U3463;
  assign new_P1_U5107 = ~new_P1_R1162_U14 | ~new_P1_U3039;
  assign new_P1_U5108 = ~P1_ADDR_REG_2_ | ~new_P1_U4932;
  assign new_P1_U5109 = ~new_P1_R1105_U68 | ~new_P1_U3042;
  assign new_P1_U5110 = ~new_P1_U3040 | ~new_P1_U3460;
  assign new_P1_U5111 = ~new_P1_R1162_U68 | ~new_P1_U3038;
  assign new_P1_U5112 = ~new_P1_U5111 | ~new_P1_U5110 | ~new_P1_U5109;
  assign new_P1_U5113 = ~new_P1_U3044 | ~new_P1_U5112;
  assign new_P1_U5114 = ~new_P1_R1105_U68 | ~new_P1_U3043;
  assign new_P1_U5115 = ~P1_REG3_REG_1_ | ~n1384;
  assign new_P1_U5116 = ~new_P1_U3041 | ~new_P1_U3460;
  assign new_P1_U5117 = ~new_P1_R1162_U68 | ~new_P1_U3039;
  assign new_P1_U5118 = ~P1_ADDR_REG_1_ | ~new_P1_U4932;
  assign new_P1_U5119 = ~new_P1_R1105_U69 | ~new_P1_U3042;
  assign new_P1_U5120 = ~new_P1_U3040 | ~new_P1_U3454;
  assign new_P1_U5121 = ~new_P1_R1162_U69 | ~new_P1_U3038;
  assign new_P1_U5122 = ~new_P1_U5121 | ~new_P1_U5120 | ~new_P1_U5119;
  assign new_P1_U5123 = ~new_P1_U3044 | ~new_P1_U5122;
  assign new_P1_U5124 = ~new_P1_R1105_U69 | ~new_P1_U3043;
  assign new_P1_U5125 = ~P1_REG3_REG_0_ | ~n1384;
  assign new_P1_U5126 = ~new_P1_U3041 | ~new_P1_U3454;
  assign new_P1_U5127 = ~new_P1_R1162_U69 | ~new_P1_U3039;
  assign new_P1_U5128 = ~P1_ADDR_REG_0_ | ~new_P1_U4932;
  assign new_P1_U5129 = ~new_P1_U3991;
  assign new_P1_U5130 = ~new_P1_U3990 | ~new_P1_U6277 | ~new_P1_U6276;
  assign new_P1_U5131 = ~new_P1_U3370 | ~new_P1_U3373;
  assign new_P1_U5132 = ~new_P1_U5802 | ~new_P1_U3451;
  assign new_P1_U5133 = ~new_P1_U3422 | ~new_P1_U5132;
  assign new_P1_U5134 = ~new_P1_U5772 | ~new_P1_U6279 | ~new_P1_U6278;
  assign new_P1_U5135 = ~new_P1_U3845 | ~new_P1_U6281 | ~new_P1_U6280;
  assign new_P1_U5136 = ~new_P1_U3432 | ~new_P1_U3022 | ~new_P1_U4029;
  assign new_P1_U5137 = ~new_P1_U4043 | ~new_P1_U5134;
  assign new_P1_U5138 = ~P1_B_REG | ~new_P1_U5135;
  assign new_P1_U5139 = ~new_P1_U3037 | ~new_P1_U3079;
  assign new_P1_U5140 = ~new_P1_U3035 | ~new_P1_U3073;
  assign new_P1_U5141 = ~new_P1_ADD_99_U73 | ~new_P1_U3434;
  assign new_P1_U5142 = ~new_P1_U5140 | ~new_P1_U5141 | ~new_P1_U5139;
  assign new_P1_U5143 = ~new_P1_U3152;
  assign new_P1_U5144 = ~new_P1_U3423 | ~new_P1_U3999;
  assign new_P1_U5145 = ~new_P1_U3848 | ~new_P1_U3849 | ~new_P1_U6283 | ~new_P1_U6282;
  assign new_P1_U5146 = ~new_P1_U5145 | ~new_P1_U3434;
  assign new_P1_U5147 = ~new_P1_U4012 | ~new_P1_U5146;
  assign new_P1_U5148 = ~new_P1_U3022 | ~new_P1_U5147;
  assign new_P1_U5149 = ~new_P1_U3503 | ~new_P1_U5770;
  assign new_P1_U5150 = ~new_P1_ADD_99_U73 | ~new_P1_U5769;
  assign new_P1_U5151 = ~new_P1_R1165_U105 | ~new_P1_U3026;
  assign new_P1_U5152 = ~new_P1_U4037 | ~new_P1_U5142;
  assign new_P1_U5153 = ~P1_REG3_REG_15_ | ~n1384;
  assign new_P1_U5154 = ~new_P1_U3037 | ~new_P1_U3058;
  assign new_P1_U5155 = ~new_P1_U3035 | ~new_P1_U3053;
  assign new_P1_U5156 = ~new_P1_ADD_99_U62 | ~new_P1_U3434;
  assign new_P1_U5157 = ~new_P1_U5155 | ~new_P1_U5156 | ~new_P1_U5154;
  assign new_P1_U5158 = ~new_P1_U4015 | ~new_P1_U3426;
  assign new_P1_U5159 = ~new_P1_U3421 | ~new_P1_U5158;
  assign new_P1_U5160 = ~new_P1_U3045 | ~new_P1_U4019;
  assign new_P1_U5161 = ~new_P1_ADD_99_U62 | ~new_P1_U5769;
  assign new_P1_U5162 = ~new_P1_R1165_U12 | ~new_P1_U3026;
  assign new_P1_U5163 = ~new_P1_U4037 | ~new_P1_U5157;
  assign new_P1_U5164 = ~P1_REG3_REG_26_ | ~n1384;
  assign new_P1_U5165 = ~new_P1_U3037 | ~new_P1_U3067;
  assign new_P1_U5166 = ~new_P1_U3035 | ~new_P1_U3070;
  assign new_P1_U5167 = ~new_P1_ADD_99_U57 | ~new_P1_U3434;
  assign new_P1_U5168 = ~new_P1_U5167 | ~new_P1_U5166 | ~new_P1_U5165;
  assign new_P1_U5169 = ~new_P1_U3476 | ~new_P1_U5770;
  assign new_P1_U5170 = ~new_P1_ADD_99_U57 | ~new_P1_U5769;
  assign new_P1_U5171 = ~new_P1_R1165_U90 | ~new_P1_U3026;
  assign new_P1_U5172 = ~new_P1_U4037 | ~new_P1_U5168;
  assign new_P1_U5173 = ~P1_REG3_REG_6_ | ~n1384;
  assign new_P1_U5174 = ~new_P1_U3037 | ~new_P1_U3069;
  assign new_P1_U5175 = ~new_P1_U3035 | ~new_P1_U3081;
  assign new_P1_U5176 = ~new_P1_ADD_99_U70 | ~new_P1_U3434;
  assign new_P1_U5177 = ~new_P1_U5175 | ~new_P1_U5176 | ~new_P1_U5174;
  assign new_P1_U5178 = ~new_P1_U3512 | ~new_P1_U5770;
  assign new_P1_U5179 = ~new_P1_ADD_99_U70 | ~new_P1_U5769;
  assign new_P1_U5180 = ~new_P1_R1165_U103 | ~new_P1_U3026;
  assign new_P1_U5181 = ~new_P1_U4037 | ~new_P1_U5177;
  assign new_P1_U5182 = ~P1_REG3_REG_18_ | ~n1384;
  assign new_P1_U5183 = ~new_P1_U3037 | ~new_P1_U3078;
  assign new_P1_U5184 = ~new_P1_U3035 | ~new_P1_U3064;
  assign new_P1_U5185 = ~P1_REG3_REG_2_ | ~new_P1_U3434;
  assign new_P1_U5186 = ~new_P1_U5185 | ~new_P1_U5184 | ~new_P1_U5183;
  assign new_P1_U5187 = ~new_P1_U3464 | ~new_P1_U5770;
  assign new_P1_U5188 = ~P1_REG3_REG_2_ | ~new_P1_U5769;
  assign new_P1_U5189 = ~new_P1_R1165_U93 | ~new_P1_U3026;
  assign new_P1_U5190 = ~new_P1_U4037 | ~new_P1_U5186;
  assign new_P1_U5191 = ~P1_REG3_REG_2_ | ~n1384;
  assign new_P1_U5192 = ~new_P1_U3037 | ~new_P1_U3062;
  assign new_P1_U5193 = ~new_P1_U3035 | ~new_P1_U3072;
  assign new_P1_U5194 = ~new_P1_ADD_99_U77 | ~new_P1_U3434;
  assign new_P1_U5195 = ~new_P1_U5194 | ~new_P1_U5193 | ~new_P1_U5192;
  assign new_P1_U5196 = ~new_P1_U3491 | ~new_P1_U5770;
  assign new_P1_U5197 = ~new_P1_ADD_99_U77 | ~new_P1_U5769;
  assign new_P1_U5198 = ~new_P1_R1165_U108 | ~new_P1_U3026;
  assign new_P1_U5199 = ~new_P1_U4037 | ~new_P1_U5195;
  assign new_P1_U5200 = ~P1_REG3_REG_11_ | ~n1384;
  assign new_P1_U5201 = ~new_P1_U3037 | ~new_P1_U3075;
  assign new_P1_U5202 = ~new_P1_U3035 | ~new_P1_U3066;
  assign new_P1_U5203 = ~new_P1_ADD_99_U66 | ~new_P1_U3434;
  assign new_P1_U5204 = ~new_P1_U5202 | ~new_P1_U5203 | ~new_P1_U5201;
  assign new_P1_U5205 = ~new_P1_U3045 | ~new_P1_U4023;
  assign new_P1_U5206 = ~new_P1_ADD_99_U66 | ~new_P1_U5769;
  assign new_P1_U5207 = ~new_P1_R1165_U99 | ~new_P1_U3026;
  assign new_P1_U5208 = ~new_P1_U4037 | ~new_P1_U5204;
  assign new_P1_U5209 = ~P1_REG3_REG_22_ | ~n1384;
  assign new_P1_U5210 = ~new_P1_U3037 | ~new_P1_U3072;
  assign new_P1_U5211 = ~new_P1_U3035 | ~new_P1_U3079;
  assign new_P1_U5212 = ~new_P1_ADD_99_U75 | ~new_P1_U3434;
  assign new_P1_U5213 = ~new_P1_U5211 | ~new_P1_U5212 | ~new_P1_U5210;
  assign new_P1_U5214 = ~new_P1_U3497 | ~new_P1_U5770;
  assign new_P1_U5215 = ~new_P1_ADD_99_U75 | ~new_P1_U5769;
  assign new_P1_U5216 = ~new_P1_R1165_U9 | ~new_P1_U3026;
  assign new_P1_U5217 = ~new_P1_U4037 | ~new_P1_U5213;
  assign new_P1_U5218 = ~P1_REG3_REG_13_ | ~n1384;
  assign new_P1_U5219 = ~new_P1_U3037 | ~new_P1_U3081;
  assign new_P1_U5220 = ~new_P1_U3035 | ~new_P1_U3075;
  assign new_P1_U5221 = ~new_P1_ADD_99_U68 | ~new_P1_U3434;
  assign new_P1_U5222 = ~new_P1_U5220 | ~new_P1_U5221 | ~new_P1_U5219;
  assign new_P1_U5223 = ~new_P1_U3045 | ~new_P1_U4025;
  assign new_P1_U5224 = ~new_P1_ADD_99_U68 | ~new_P1_U5769;
  assign new_P1_U5225 = ~new_P1_R1165_U100 | ~new_P1_U3026;
  assign new_P1_U5226 = ~new_P1_U4037 | ~new_P1_U5222;
  assign new_P1_U5227 = ~P1_REG3_REG_20_ | ~n1384;
  assign new_P1_U5228 = ~new_P1_U3435 | ~new_P1_U3433;
  assign new_P1_U5229 = ~new_P1_U5228 | ~new_P1_U3434;
  assign new_P1_U5230 = ~new_P1_U3050 | ~new_P1_U5229;
  assign new_P1_U5231 = ~new_P1_U3858 | ~new_P1_U3035;
  assign new_P1_U5232 = ~new_P1_U3456 | ~new_P1_U5770;
  assign new_P1_U5233 = ~P1_REG3_REG_0_ | ~new_P1_U5230;
  assign new_P1_U5234 = ~new_P1_R1165_U87 | ~new_P1_U3026;
  assign new_P1_U5235 = ~P1_REG3_REG_0_ | ~n1384;
  assign new_P1_U5236 = ~new_P1_U3037 | ~new_P1_U3084;
  assign new_P1_U5237 = ~new_P1_U3035 | ~new_P1_U3062;
  assign new_P1_U5238 = ~new_P1_ADD_99_U54 | ~new_P1_U3434;
  assign new_P1_U5239 = ~new_P1_U5238 | ~new_P1_U5237 | ~new_P1_U5236;
  assign new_P1_U5240 = ~new_P1_U3485 | ~new_P1_U5770;
  assign new_P1_U5241 = ~new_P1_ADD_99_U54 | ~new_P1_U5769;
  assign new_P1_U5242 = ~new_P1_R1165_U88 | ~new_P1_U3026;
  assign new_P1_U5243 = ~new_P1_U4037 | ~new_P1_U5239;
  assign new_P1_U5244 = ~P1_REG3_REG_9_ | ~n1384;
  assign new_P1_U5245 = ~new_P1_U3037 | ~new_P1_U3064;
  assign new_P1_U5246 = ~new_P1_U3035 | ~new_P1_U3067;
  assign new_P1_U5247 = ~new_P1_ADD_99_U59 | ~new_P1_U3434;
  assign new_P1_U5248 = ~new_P1_U5247 | ~new_P1_U5246 | ~new_P1_U5245;
  assign new_P1_U5249 = ~new_P1_U3470 | ~new_P1_U5770;
  assign new_P1_U5250 = ~new_P1_ADD_99_U59 | ~new_P1_U5769;
  assign new_P1_U5251 = ~new_P1_R1165_U92 | ~new_P1_U3026;
  assign new_P1_U5252 = ~new_P1_U4037 | ~new_P1_U5248;
  assign new_P1_U5253 = ~P1_REG3_REG_4_ | ~n1384;
  assign new_P1_U5254 = ~new_P1_U3037 | ~new_P1_U3066;
  assign new_P1_U5255 = ~new_P1_U3035 | ~new_P1_U3058;
  assign new_P1_U5256 = ~new_P1_ADD_99_U64 | ~new_P1_U3434;
  assign new_P1_U5257 = ~new_P1_U5255 | ~new_P1_U5256 | ~new_P1_U5254;
  assign new_P1_U5258 = ~new_P1_U3045 | ~new_P1_U4021;
  assign new_P1_U5259 = ~new_P1_ADD_99_U64 | ~new_P1_U5769;
  assign new_P1_U5260 = ~new_P1_R1165_U97 | ~new_P1_U3026;
  assign new_P1_U5261 = ~new_P1_U4037 | ~new_P1_U5257;
  assign new_P1_U5262 = ~P1_REG3_REG_24_ | ~n1384;
  assign new_P1_U5263 = ~new_P1_U3037 | ~new_P1_U3073;
  assign new_P1_U5264 = ~new_P1_U3035 | ~new_P1_U3082;
  assign new_P1_U5265 = ~new_P1_ADD_99_U71 | ~new_P1_U3434;
  assign new_P1_U5266 = ~new_P1_U5264 | ~new_P1_U5265 | ~new_P1_U5263;
  assign new_P1_U5267 = ~new_P1_U3509 | ~new_P1_U5770;
  assign new_P1_U5268 = ~new_P1_ADD_99_U71 | ~new_P1_U5769;
  assign new_P1_U5269 = ~new_P1_R1165_U10 | ~new_P1_U3026;
  assign new_P1_U5270 = ~new_P1_U4037 | ~new_P1_U5266;
  assign new_P1_U5271 = ~P1_REG3_REG_17_ | ~n1384;
  assign new_P1_U5272 = ~new_P1_U3037 | ~new_P1_U3060;
  assign new_P1_U5273 = ~new_P1_U3035 | ~new_P1_U3071;
  assign new_P1_U5274 = ~new_P1_ADD_99_U58 | ~new_P1_U3434;
  assign new_P1_U5275 = ~new_P1_U5274 | ~new_P1_U5273 | ~new_P1_U5272;
  assign new_P1_U5276 = ~new_P1_U3473 | ~new_P1_U5770;
  assign new_P1_U5277 = ~new_P1_ADD_99_U58 | ~new_P1_U5769;
  assign new_P1_U5278 = ~new_P1_R1165_U91 | ~new_P1_U3026;
  assign new_P1_U5279 = ~new_P1_U4037 | ~new_P1_U5275;
  assign new_P1_U5280 = ~P1_REG3_REG_5_ | ~n1384;
  assign new_P1_U5281 = ~new_P1_U3037 | ~new_P1_U3074;
  assign new_P1_U5282 = ~new_P1_U3035 | ~new_P1_U3069;
  assign new_P1_U5283 = ~new_P1_ADD_99_U72 | ~new_P1_U3434;
  assign new_P1_U5284 = ~new_P1_U5282 | ~new_P1_U5283 | ~new_P1_U5281;
  assign new_P1_U5285 = ~new_P1_U3506 | ~new_P1_U5770;
  assign new_P1_U5286 = ~new_P1_ADD_99_U72 | ~new_P1_U5769;
  assign new_P1_U5287 = ~new_P1_R1165_U104 | ~new_P1_U3026;
  assign new_P1_U5288 = ~new_P1_U4037 | ~new_P1_U5284;
  assign new_P1_U5289 = ~P1_REG3_REG_16_ | ~n1384;
  assign new_P1_U5290 = ~new_P1_U3037 | ~new_P1_U3065;
  assign new_P1_U5291 = ~new_P1_U3035 | ~new_P1_U3057;
  assign new_P1_U5292 = ~new_P1_ADD_99_U63 | ~new_P1_U3434;
  assign new_P1_U5293 = ~new_P1_U5291 | ~new_P1_U5292 | ~new_P1_U5290;
  assign new_P1_U5294 = ~new_P1_U3045 | ~new_P1_U4020;
  assign new_P1_U5295 = ~new_P1_ADD_99_U63 | ~new_P1_U5769;
  assign new_P1_U5296 = ~new_P1_R1165_U96 | ~new_P1_U3026;
  assign new_P1_U5297 = ~new_P1_U4037 | ~new_P1_U5293;
  assign new_P1_U5298 = ~P1_REG3_REG_25_ | ~n1384;
  assign new_P1_U5299 = ~new_P1_U3037 | ~new_P1_U3063;
  assign new_P1_U5300 = ~new_P1_U3035 | ~new_P1_U3080;
  assign new_P1_U5301 = ~new_P1_ADD_99_U76 | ~new_P1_U3434;
  assign new_P1_U5302 = ~new_P1_U5300 | ~new_P1_U5301 | ~new_P1_U5299;
  assign new_P1_U5303 = ~new_P1_U3494 | ~new_P1_U5770;
  assign new_P1_U5304 = ~new_P1_ADD_99_U76 | ~new_P1_U5769;
  assign new_P1_U5305 = ~new_P1_R1165_U107 | ~new_P1_U3026;
  assign new_P1_U5306 = ~new_P1_U4037 | ~new_P1_U5302;
  assign new_P1_U5307 = ~P1_REG3_REG_12_ | ~n1384;
  assign new_P1_U5308 = ~new_P1_U3037 | ~new_P1_U3076;
  assign new_P1_U5309 = ~new_P1_U3035 | ~new_P1_U3061;
  assign new_P1_U5310 = ~new_P1_ADD_99_U67 | ~new_P1_U3434;
  assign new_P1_U5311 = ~new_P1_U5309 | ~new_P1_U5310 | ~new_P1_U5308;
  assign new_P1_U5312 = ~new_P1_U3045 | ~new_P1_U4024;
  assign new_P1_U5313 = ~new_P1_ADD_99_U67 | ~new_P1_U5769;
  assign new_P1_U5314 = ~new_P1_R1165_U11 | ~new_P1_U3026;
  assign new_P1_U5315 = ~new_P1_U4037 | ~new_P1_U5311;
  assign new_P1_U5316 = ~P1_REG3_REG_21_ | ~n1384;
  assign new_P1_U5317 = ~new_P1_U3037 | ~new_P1_U3077;
  assign new_P1_U5318 = ~new_P1_U3035 | ~new_P1_U3068;
  assign new_P1_U5319 = ~P1_REG3_REG_1_ | ~new_P1_U3434;
  assign new_P1_U5320 = ~new_P1_U5319 | ~new_P1_U5318 | ~new_P1_U5317;
  assign new_P1_U5321 = ~new_P1_U3461 | ~new_P1_U5770;
  assign new_P1_U5322 = ~P1_REG3_REG_1_ | ~new_P1_U5769;
  assign new_P1_U5323 = ~new_P1_R1165_U101 | ~new_P1_U3026;
  assign new_P1_U5324 = ~new_P1_U4037 | ~new_P1_U5320;
  assign new_P1_U5325 = ~P1_REG3_REG_1_ | ~n1384;
  assign new_P1_U5326 = ~new_P1_U3037 | ~new_P1_U3070;
  assign new_P1_U5327 = ~new_P1_U3035 | ~new_P1_U3083;
  assign new_P1_U5328 = ~new_P1_ADD_99_U55 | ~new_P1_U3434;
  assign new_P1_U5329 = ~new_P1_U5328 | ~new_P1_U5327 | ~new_P1_U5326;
  assign new_P1_U5330 = ~new_P1_U3482 | ~new_P1_U5770;
  assign new_P1_U5331 = ~new_P1_ADD_99_U55 | ~new_P1_U5769;
  assign new_P1_U5332 = ~new_P1_R1165_U89 | ~new_P1_U3026;
  assign new_P1_U5333 = ~new_P1_U4037 | ~new_P1_U5329;
  assign new_P1_U5334 = ~P1_REG3_REG_8_ | ~n1384;
  assign new_P1_U5335 = ~new_P1_U3037 | ~new_P1_U3053;
  assign new_P1_U5336 = ~new_P1_U3035 | ~new_P1_U3055;
  assign new_P1_U5337 = ~new_P1_ADD_99_U60 | ~new_P1_U3434;
  assign new_P1_U5338 = ~new_P1_U5337 | ~new_P1_U5336 | ~new_P1_U5335;
  assign new_P1_U5339 = ~new_P1_U3045 | ~new_P1_U4017;
  assign new_P1_U5340 = ~new_P1_ADD_99_U60 | ~new_P1_U5769;
  assign new_P1_U5341 = ~new_P1_R1165_U94 | ~new_P1_U3026;
  assign new_P1_U5342 = ~new_P1_U4037 | ~new_P1_U5338;
  assign new_P1_U5343 = ~P1_REG3_REG_28_ | ~n1384;
  assign new_P1_U5344 = ~new_P1_U3037 | ~new_P1_U3082;
  assign new_P1_U5345 = ~new_P1_U3035 | ~new_P1_U3076;
  assign new_P1_U5346 = ~new_P1_ADD_99_U69 | ~new_P1_U3434;
  assign new_P1_U5347 = ~new_P1_U5345 | ~new_P1_U5346 | ~new_P1_U5344;
  assign new_P1_U5348 = ~new_P1_U3514 | ~new_P1_U5770;
  assign new_P1_U5349 = ~new_P1_ADD_99_U69 | ~new_P1_U5769;
  assign new_P1_U5350 = ~new_P1_R1165_U102 | ~new_P1_U3026;
  assign new_P1_U5351 = ~new_P1_U4037 | ~new_P1_U5347;
  assign new_P1_U5352 = ~P1_REG3_REG_19_ | ~n1384;
  assign new_P1_U5353 = ~new_P1_U3037 | ~new_P1_U3068;
  assign new_P1_U5354 = ~new_P1_U3035 | ~new_P1_U3060;
  assign new_P1_U5355 = ~new_P1_ADD_99_U4 | ~new_P1_U3434;
  assign new_P1_U5356 = ~new_P1_U5355 | ~new_P1_U5354 | ~new_P1_U5353;
  assign new_P1_U5357 = ~new_P1_U3467 | ~new_P1_U5770;
  assign new_P1_U5358 = ~new_P1_ADD_99_U4 | ~new_P1_U5769;
  assign new_P1_U5359 = ~new_P1_R1165_U13 | ~new_P1_U3026;
  assign new_P1_U5360 = ~new_P1_U4037 | ~new_P1_U5356;
  assign new_P1_U5361 = ~P1_REG3_REG_3_ | ~n1384;
  assign new_P1_U5362 = ~new_P1_U3037 | ~new_P1_U3083;
  assign new_P1_U5363 = ~new_P1_U3035 | ~new_P1_U3063;
  assign new_P1_U5364 = ~new_P1_ADD_99_U78 | ~new_P1_U3434;
  assign new_P1_U5365 = ~new_P1_U5364 | ~new_P1_U5363 | ~new_P1_U5362;
  assign new_P1_U5366 = ~new_P1_U3488 | ~new_P1_U5770;
  assign new_P1_U5367 = ~new_P1_ADD_99_U78 | ~new_P1_U5769;
  assign new_P1_U5368 = ~new_P1_R1165_U109 | ~new_P1_U3026;
  assign new_P1_U5369 = ~new_P1_U4037 | ~new_P1_U5365;
  assign new_P1_U5370 = ~P1_REG3_REG_10_ | ~n1384;
  assign new_P1_U5371 = ~new_P1_U3037 | ~new_P1_U3061;
  assign new_P1_U5372 = ~new_P1_U3035 | ~new_P1_U3065;
  assign new_P1_U5373 = ~new_P1_ADD_99_U65 | ~new_P1_U3434;
  assign new_P1_U5374 = ~new_P1_U5372 | ~new_P1_U5373 | ~new_P1_U5371;
  assign new_P1_U5375 = ~new_P1_U3045 | ~new_P1_U4022;
  assign new_P1_U5376 = ~new_P1_ADD_99_U65 | ~new_P1_U5769;
  assign new_P1_U5377 = ~new_P1_R1165_U98 | ~new_P1_U3026;
  assign new_P1_U5378 = ~new_P1_U4037 | ~new_P1_U5374;
  assign new_P1_U5379 = ~P1_REG3_REG_23_ | ~n1384;
  assign new_P1_U5380 = ~new_P1_U3037 | ~new_P1_U3080;
  assign new_P1_U5381 = ~new_P1_U3035 | ~new_P1_U3074;
  assign new_P1_U5382 = ~new_P1_ADD_99_U74 | ~new_P1_U3434;
  assign new_P1_U5383 = ~new_P1_U5381 | ~new_P1_U5382 | ~new_P1_U5380;
  assign new_P1_U5384 = ~new_P1_U3500 | ~new_P1_U5770;
  assign new_P1_U5385 = ~new_P1_ADD_99_U74 | ~new_P1_U5769;
  assign new_P1_U5386 = ~new_P1_R1165_U106 | ~new_P1_U3026;
  assign new_P1_U5387 = ~new_P1_U4037 | ~new_P1_U5383;
  assign new_P1_U5388 = ~P1_REG3_REG_14_ | ~n1384;
  assign new_P1_U5389 = ~new_P1_U3037 | ~new_P1_U3057;
  assign new_P1_U5390 = ~new_P1_U3035 | ~new_P1_U3054;
  assign new_P1_U5391 = ~new_P1_ADD_99_U61 | ~new_P1_U3434;
  assign new_P1_U5392 = ~new_P1_U5390 | ~new_P1_U5391 | ~new_P1_U5389;
  assign new_P1_U5393 = ~new_P1_U3045 | ~new_P1_U4018;
  assign new_P1_U5394 = ~new_P1_ADD_99_U61 | ~new_P1_U5769;
  assign new_P1_U5395 = ~new_P1_R1165_U95 | ~new_P1_U3026;
  assign new_P1_U5396 = ~new_P1_U4037 | ~new_P1_U5392;
  assign new_P1_U5397 = ~P1_REG3_REG_27_ | ~n1384;
  assign new_P1_U5398 = ~new_P1_U3037 | ~new_P1_U3071;
  assign new_P1_U5399 = ~new_P1_U3035 | ~new_P1_U3084;
  assign new_P1_U5400 = ~new_P1_ADD_99_U56 | ~new_P1_U3434;
  assign new_P1_U5401 = ~new_P1_U5400 | ~new_P1_U5399 | ~new_P1_U5398;
  assign new_P1_U5402 = ~new_P1_U3479 | ~new_P1_U5770;
  assign new_P1_U5403 = ~new_P1_ADD_99_U56 | ~new_P1_U5769;
  assign new_P1_U5404 = ~new_P1_R1165_U14 | ~new_P1_U3026;
  assign new_P1_U5405 = ~new_P1_U4037 | ~new_P1_U5401;
  assign new_P1_U5406 = ~P1_REG3_REG_7_ | ~n1384;
  assign new_P1_U5407 = ~new_P1_U3455 | ~new_P1_U3377;
  assign new_P1_U5408 = ~new_P1_U3449 | ~new_P1_U5407;
  assign new_P1_U5409 = ~new_P1_R1165_U87 | ~new_P1_U5817 | ~new_P1_U3449;
  assign new_P1_U5410 = ~new_P1_U3450 | ~new_P1_U3453;
  assign new_P1_U5411 = ~new_P1_U3874 | ~new_P1_U4013;
  assign new_P1_U5412 = ~new_P1_U3370 | ~new_P1_U3422;
  assign new_P1_U5413 = ~new_P1_U3365 | ~new_P1_U4006 | ~new_P1_U3363;
  assign new_P1_U5414 = ~new_P1_U4041 | ~new_P1_U3425;
  assign new_P1_U5415 = ~new_P1_U5413 | ~new_P1_U3425;
  assign new_P1_U5416 = ~new_P1_U3436;
  assign new_P1_U5417 = ~new_P1_U5416 | ~new_P1_U4013;
  assign new_P1_U5418 = ~new_P1_U3485 | ~new_P1_U5417;
  assign new_P1_U5419 = ~new_P1_U3021 | ~new_P1_U3083;
  assign new_P1_U5420 = ~new_P1_U3482 | ~new_P1_U5417;
  assign new_P1_U5421 = ~new_P1_U3021 | ~new_P1_U3084;
  assign new_P1_U5422 = ~new_P1_U3479 | ~new_P1_U5417;
  assign new_P1_U5423 = ~new_P1_U3021 | ~new_P1_U3070;
  assign new_P1_U5424 = ~new_P1_U3476 | ~new_P1_U5417;
  assign new_P1_U5425 = ~new_P1_U3021 | ~new_P1_U3071;
  assign new_P1_U5426 = ~new_P1_U3473 | ~new_P1_U5417;
  assign new_P1_U5427 = ~new_P1_U3021 | ~new_P1_U3067;
  assign new_P1_U5428 = ~new_P1_U3470 | ~new_P1_U5417;
  assign new_P1_U5429 = ~new_P1_U3021 | ~new_P1_U3060;
  assign new_P1_U5430 = ~new_P1_U3467 | ~new_P1_U5417;
  assign new_P1_U5431 = ~new_P1_U3021 | ~new_P1_U3064;
  assign new_P1_U5432 = ~new_P1_U4017 | ~new_P1_U5417;
  assign new_P1_U5433 = ~new_P1_U3021 | ~new_P1_U3054;
  assign new_P1_U5434 = ~new_P1_U4018 | ~new_P1_U5417;
  assign new_P1_U5435 = ~new_P1_U3021 | ~new_P1_U3053;
  assign new_P1_U5436 = ~new_P1_U4019 | ~new_P1_U5417;
  assign new_P1_U5437 = ~new_P1_U3021 | ~new_P1_U3057;
  assign new_P1_U5438 = ~new_P1_U4020 | ~new_P1_U5417;
  assign new_P1_U5439 = ~new_P1_U3021 | ~new_P1_U3058;
  assign new_P1_U5440 = ~new_P1_U4021 | ~new_P1_U5417;
  assign new_P1_U5441 = ~new_P1_U3021 | ~new_P1_U3065;
  assign new_P1_U5442 = ~new_P1_U4022 | ~new_P1_U5417;
  assign new_P1_U5443 = ~new_P1_U3021 | ~new_P1_U3066;
  assign new_P1_U5444 = ~new_P1_U4023 | ~new_P1_U5417;
  assign new_P1_U5445 = ~new_P1_U3021 | ~new_P1_U3061;
  assign new_P1_U5446 = ~new_P1_U4024 | ~new_P1_U5417;
  assign new_P1_U5447 = ~new_P1_U3021 | ~new_P1_U3075;
  assign new_P1_U5448 = ~new_P1_U4025 | ~new_P1_U5417;
  assign new_P1_U5449 = ~new_P1_U3021 | ~new_P1_U3076;
  assign new_P1_U5450 = ~new_P1_U3464 | ~new_P1_U5417;
  assign new_P1_U5451 = ~new_P1_U3021 | ~new_P1_U3068;
  assign new_P1_U5452 = ~new_P1_U3514 | ~new_P1_U5417;
  assign new_P1_U5453 = ~new_P1_U3021 | ~new_P1_U3081;
  assign new_P1_U5454 = ~new_P1_U3512 | ~new_P1_U5417;
  assign new_P1_U5455 = ~new_P1_U3021 | ~new_P1_U3082;
  assign new_P1_U5456 = ~new_P1_U3509 | ~new_P1_U5417;
  assign new_P1_U5457 = ~new_P1_U3021 | ~new_P1_U3069;
  assign new_P1_U5458 = ~new_P1_U3506 | ~new_P1_U5417;
  assign new_P1_U5459 = ~new_P1_U3021 | ~new_P1_U3073;
  assign new_P1_U5460 = ~new_P1_U3503 | ~new_P1_U5417;
  assign new_P1_U5461 = ~new_P1_U3021 | ~new_P1_U3074;
  assign new_P1_U5462 = ~new_P1_U3500 | ~new_P1_U5417;
  assign new_P1_U5463 = ~new_P1_U3021 | ~new_P1_U3079;
  assign new_P1_U5464 = ~new_P1_U3497 | ~new_P1_U5417;
  assign new_P1_U5465 = ~new_P1_U3021 | ~new_P1_U3080;
  assign new_P1_U5466 = ~new_P1_U3494 | ~new_P1_U5417;
  assign new_P1_U5467 = ~new_P1_U3021 | ~new_P1_U3072;
  assign new_P1_U5468 = ~new_P1_U3491 | ~new_P1_U5417;
  assign new_P1_U5469 = ~new_P1_U3021 | ~new_P1_U3063;
  assign new_P1_U5470 = ~new_P1_U3488 | ~new_P1_U5417;
  assign new_P1_U5471 = ~new_P1_U3021 | ~new_P1_U3062;
  assign new_P1_U5472 = ~new_P1_U3461 | ~new_P1_U5417;
  assign new_P1_U5473 = ~new_P1_U3021 | ~new_P1_U3078;
  assign new_P1_U5474 = ~new_P1_U3456 | ~new_P1_U5417;
  assign new_P1_U5475 = ~new_P1_U3021 | ~new_P1_U3077;
  assign new_P1_U5476 = ~new_P1_U4145 | ~P1_REG1_REG_0_;
  assign new_P1_U5477 = ~new_P1_U3021 | ~new_P1_U3485;
  assign new_P1_U5478 = ~new_P1_U3436 | ~new_P1_U3083;
  assign new_P1_U5479 = ~new_P1_U3021 | ~new_P1_U3482;
  assign new_P1_U5480 = ~new_P1_U3436 | ~new_P1_U3084;
  assign new_P1_U5481 = ~new_P1_U3021 | ~new_P1_U3479;
  assign new_P1_U5482 = ~new_P1_U3436 | ~new_P1_U3070;
  assign new_P1_U5483 = ~new_P1_U3021 | ~new_P1_U3476;
  assign new_P1_U5484 = ~new_P1_U3436 | ~new_P1_U3071;
  assign new_P1_U5485 = ~new_P1_U3021 | ~new_P1_U3473;
  assign new_P1_U5486 = ~new_P1_U3436 | ~new_P1_U3067;
  assign new_P1_U5487 = ~new_P1_U3021 | ~new_P1_U3470;
  assign new_P1_U5488 = ~new_P1_U3436 | ~new_P1_U3060;
  assign new_P1_U5489 = ~new_P1_U3021 | ~new_P1_U3467;
  assign new_P1_U5490 = ~new_P1_U3436 | ~new_P1_U3064;
  assign new_P1_U5491 = ~new_P1_U3021 | ~new_P1_U4017;
  assign new_P1_U5492 = ~new_P1_U3436 | ~new_P1_U3054;
  assign new_P1_U5493 = ~new_P1_U3021 | ~new_P1_U4018;
  assign new_P1_U5494 = ~new_P1_U3436 | ~new_P1_U3053;
  assign new_P1_U5495 = ~new_P1_U3021 | ~new_P1_U4019;
  assign new_P1_U5496 = ~new_P1_U3436 | ~new_P1_U3057;
  assign new_P1_U5497 = ~new_P1_U3021 | ~new_P1_U4020;
  assign new_P1_U5498 = ~new_P1_U3436 | ~new_P1_U3058;
  assign new_P1_U5499 = ~new_P1_U3021 | ~new_P1_U4021;
  assign new_P1_U5500 = ~new_P1_U3436 | ~new_P1_U3065;
  assign new_P1_U5501 = ~new_P1_U3021 | ~new_P1_U4022;
  assign new_P1_U5502 = ~new_P1_U3436 | ~new_P1_U3066;
  assign new_P1_U5503 = ~new_P1_U3021 | ~new_P1_U4023;
  assign new_P1_U5504 = ~new_P1_U3436 | ~new_P1_U3061;
  assign new_P1_U5505 = ~new_P1_U3021 | ~new_P1_U4024;
  assign new_P1_U5506 = ~new_P1_U3436 | ~new_P1_U3075;
  assign new_P1_U5507 = ~new_P1_U3021 | ~new_P1_U4025;
  assign new_P1_U5508 = ~new_P1_U3436 | ~new_P1_U3076;
  assign new_P1_U5509 = ~new_P1_U3021 | ~new_P1_U3464;
  assign new_P1_U5510 = ~new_P1_U3436 | ~new_P1_U3068;
  assign new_P1_U5511 = ~new_P1_U3021 | ~new_P1_U3514;
  assign new_P1_U5512 = ~new_P1_U3436 | ~new_P1_U3081;
  assign new_P1_U5513 = ~new_P1_U3021 | ~new_P1_U3512;
  assign new_P1_U5514 = ~new_P1_U3436 | ~new_P1_U3082;
  assign new_P1_U5515 = ~new_P1_U3021 | ~new_P1_U3509;
  assign new_P1_U5516 = ~new_P1_U3436 | ~new_P1_U3069;
  assign new_P1_U5517 = ~new_P1_U3021 | ~new_P1_U3506;
  assign new_P1_U5518 = ~new_P1_U3436 | ~new_P1_U3073;
  assign new_P1_U5519 = ~new_P1_U3021 | ~new_P1_U3503;
  assign new_P1_U5520 = ~new_P1_U3436 | ~new_P1_U3074;
  assign new_P1_U5521 = ~new_P1_U3021 | ~new_P1_U3500;
  assign new_P1_U5522 = ~new_P1_U3436 | ~new_P1_U3079;
  assign new_P1_U5523 = ~new_P1_U3021 | ~new_P1_U3497;
  assign new_P1_U5524 = ~new_P1_U3436 | ~new_P1_U3080;
  assign new_P1_U5525 = ~new_P1_U3021 | ~new_P1_U3494;
  assign new_P1_U5526 = ~new_P1_U3436 | ~new_P1_U3072;
  assign new_P1_U5527 = ~new_P1_U3021 | ~new_P1_U3491;
  assign new_P1_U5528 = ~new_P1_U3436 | ~new_P1_U3063;
  assign new_P1_U5529 = ~new_P1_U3021 | ~new_P1_U3488;
  assign new_P1_U5530 = ~new_P1_U3436 | ~new_P1_U3062;
  assign new_P1_U5531 = ~new_P1_U3021 | ~new_P1_U3461;
  assign new_P1_U5532 = ~new_P1_U3436 | ~new_P1_U3078;
  assign new_P1_U5533 = ~new_P1_U3021 | ~new_P1_U3456;
  assign new_P1_U5534 = ~new_P1_U3436 | ~new_P1_U3077;
  assign new_P1_U5535 = ~new_P1_U4145 | ~new_P1_U3454;
  assign new_P1_U5536 = ~new_P1_U3437;
  assign new_P1_U5537 = ~new_P1_U3438;
  assign new_P1_U5538 = ~new_P1_U5799 | ~new_P1_U3450;
  assign new_P1_U5539 = ~new_P1_U3437 | ~new_P1_U3439;
  assign new_P1_U5540 = ~new_P1_U3051 | ~new_P1_U5539;
  assign new_P1_U5541 = ~new_P1_U3014 | ~new_P1_U3444;
  assign new_P1_U5542 = ~new_P1_U3440;
  assign new_P1_U5543 = ~new_P1_U3052 | ~new_P1_U5542;
  assign new_P1_U5544 = ~new_P1_U3083 | ~new_P1_U3027;
  assign new_P1_U5545 = ~new_P1_U3485 | ~new_P1_U5543;
  assign new_P1_U5546 = ~new_P1_U5540 | ~new_P1_U3083;
  assign new_P1_U5547 = ~new_P1_U3084 | ~new_P1_U3027;
  assign new_P1_U5548 = ~new_P1_U3482 | ~new_P1_U5543;
  assign new_P1_U5549 = ~new_P1_U5540 | ~new_P1_U3084;
  assign new_P1_U5550 = ~new_P1_U3070 | ~new_P1_U3027;
  assign new_P1_U5551 = ~new_P1_U3479 | ~new_P1_U5543;
  assign new_P1_U5552 = ~new_P1_U5540 | ~new_P1_U3070;
  assign new_P1_U5553 = ~new_P1_U3071 | ~new_P1_U3027;
  assign new_P1_U5554 = ~new_P1_U3476 | ~new_P1_U5543;
  assign new_P1_U5555 = ~new_P1_U5540 | ~new_P1_U3071;
  assign new_P1_U5556 = ~new_P1_U3067 | ~new_P1_U3027;
  assign new_P1_U5557 = ~new_P1_U3473 | ~new_P1_U5543;
  assign new_P1_U5558 = ~new_P1_U5540 | ~new_P1_U3067;
  assign new_P1_U5559 = ~new_P1_U3060 | ~new_P1_U3027;
  assign new_P1_U5560 = ~new_P1_U3470 | ~new_P1_U5543;
  assign new_P1_U5561 = ~new_P1_U5540 | ~new_P1_U3060;
  assign new_P1_U5562 = ~new_P1_R1309_U8 | ~new_P1_U3027;
  assign new_P1_U5563 = ~new_P1_U4026 | ~new_P1_U5543;
  assign new_P1_U5564 = ~new_P1_U5540 | ~new_P1_U3056;
  assign new_P1_U5565 = ~new_P1_R1309_U6 | ~new_P1_U3027;
  assign new_P1_U5566 = ~new_P1_U4027 | ~new_P1_U5543;
  assign new_P1_U5567 = ~new_P1_U5540 | ~new_P1_U3059;
  assign new_P1_U5568 = ~new_P1_U3064 | ~new_P1_U3027;
  assign new_P1_U5569 = ~new_P1_U3467 | ~new_P1_U5543;
  assign new_P1_U5570 = ~new_P1_U5540 | ~new_P1_U3064;
  assign new_P1_U5571 = ~new_P1_U3055 | ~new_P1_U3027;
  assign new_P1_U5572 = ~new_P1_U4028 | ~new_P1_U5543;
  assign new_P1_U5573 = ~new_P1_U5540 | ~new_P1_U3055;
  assign new_P1_U5574 = ~new_P1_U3054 | ~new_P1_U3027;
  assign new_P1_U5575 = ~new_P1_U4017 | ~new_P1_U5543;
  assign new_P1_U5576 = ~new_P1_U5540 | ~new_P1_U3054;
  assign new_P1_U5577 = ~new_P1_U3053 | ~new_P1_U3027;
  assign new_P1_U5578 = ~new_P1_U4018 | ~new_P1_U5543;
  assign new_P1_U5579 = ~new_P1_U5540 | ~new_P1_U3053;
  assign new_P1_U5580 = ~new_P1_U3057 | ~new_P1_U3027;
  assign new_P1_U5581 = ~new_P1_U4019 | ~new_P1_U5543;
  assign new_P1_U5582 = ~new_P1_U5540 | ~new_P1_U3057;
  assign new_P1_U5583 = ~new_P1_U3058 | ~new_P1_U3027;
  assign new_P1_U5584 = ~new_P1_U4020 | ~new_P1_U5543;
  assign new_P1_U5585 = ~new_P1_U5540 | ~new_P1_U3058;
  assign new_P1_U5586 = ~new_P1_U3065 | ~new_P1_U3027;
  assign new_P1_U5587 = ~new_P1_U4021 | ~new_P1_U5543;
  assign new_P1_U5588 = ~new_P1_U5540 | ~new_P1_U3065;
  assign new_P1_U5589 = ~new_P1_U3066 | ~new_P1_U3027;
  assign new_P1_U5590 = ~new_P1_U4022 | ~new_P1_U5543;
  assign new_P1_U5591 = ~new_P1_U5540 | ~new_P1_U3066;
  assign new_P1_U5592 = ~new_P1_U3061 | ~new_P1_U3027;
  assign new_P1_U5593 = ~new_P1_U4023 | ~new_P1_U5543;
  assign new_P1_U5594 = ~new_P1_U5540 | ~new_P1_U3061;
  assign new_P1_U5595 = ~new_P1_U3075 | ~new_P1_U3027;
  assign new_P1_U5596 = ~new_P1_U4024 | ~new_P1_U5543;
  assign new_P1_U5597 = ~new_P1_U5540 | ~new_P1_U3075;
  assign new_P1_U5598 = ~new_P1_U3076 | ~new_P1_U3027;
  assign new_P1_U5599 = ~new_P1_U4025 | ~new_P1_U5543;
  assign new_P1_U5600 = ~new_P1_U5540 | ~new_P1_U3076;
  assign new_P1_U5601 = ~new_P1_U3068 | ~new_P1_U3027;
  assign new_P1_U5602 = ~new_P1_U3464 | ~new_P1_U5543;
  assign new_P1_U5603 = ~new_P1_U5540 | ~new_P1_U3068;
  assign new_P1_U5604 = ~new_P1_U3081 | ~new_P1_U3027;
  assign new_P1_U5605 = ~new_P1_U3514 | ~new_P1_U5543;
  assign new_P1_U5606 = ~new_P1_U5540 | ~new_P1_U3081;
  assign new_P1_U5607 = ~new_P1_U3082 | ~new_P1_U3027;
  assign new_P1_U5608 = ~new_P1_U3512 | ~new_P1_U5543;
  assign new_P1_U5609 = ~new_P1_U5540 | ~new_P1_U3082;
  assign new_P1_U5610 = ~new_P1_U3069 | ~new_P1_U3027;
  assign new_P1_U5611 = ~new_P1_U3509 | ~new_P1_U5543;
  assign new_P1_U5612 = ~new_P1_U5540 | ~new_P1_U3069;
  assign new_P1_U5613 = ~new_P1_U3073 | ~new_P1_U3027;
  assign new_P1_U5614 = ~new_P1_U3506 | ~new_P1_U5543;
  assign new_P1_U5615 = ~new_P1_U5540 | ~new_P1_U3073;
  assign new_P1_U5616 = ~new_P1_U3074 | ~new_P1_U3027;
  assign new_P1_U5617 = ~new_P1_U3503 | ~new_P1_U5543;
  assign new_P1_U5618 = ~new_P1_U5540 | ~new_P1_U3074;
  assign new_P1_U5619 = ~new_P1_U3079 | ~new_P1_U3027;
  assign new_P1_U5620 = ~new_P1_U3500 | ~new_P1_U5543;
  assign new_P1_U5621 = ~new_P1_U5540 | ~new_P1_U3079;
  assign new_P1_U5622 = ~new_P1_U3080 | ~new_P1_U3027;
  assign new_P1_U5623 = ~new_P1_U3497 | ~new_P1_U5543;
  assign new_P1_U5624 = ~new_P1_U5540 | ~new_P1_U3080;
  assign new_P1_U5625 = ~new_P1_U3072 | ~new_P1_U3027;
  assign new_P1_U5626 = ~new_P1_U3494 | ~new_P1_U5543;
  assign new_P1_U5627 = ~new_P1_U5540 | ~new_P1_U3072;
  assign new_P1_U5628 = ~new_P1_U3063 | ~new_P1_U3027;
  assign new_P1_U5629 = ~new_P1_U3491 | ~new_P1_U5543;
  assign new_P1_U5630 = ~new_P1_U5540 | ~new_P1_U3063;
  assign new_P1_U5631 = ~new_P1_U3062 | ~new_P1_U3027;
  assign new_P1_U5632 = ~new_P1_U3488 | ~new_P1_U5543;
  assign new_P1_U5633 = ~new_P1_U5540 | ~new_P1_U3062;
  assign new_P1_U5634 = ~new_P1_U3078 | ~new_P1_U3027;
  assign new_P1_U5635 = ~new_P1_U3461 | ~new_P1_U5543;
  assign new_P1_U5636 = ~new_P1_U5540 | ~new_P1_U3078;
  assign new_P1_U5637 = ~new_P1_U3077 | ~new_P1_U3027;
  assign new_P1_U5638 = ~new_P1_U3456 | ~new_P1_U5543;
  assign new_P1_U5639 = ~new_P1_U5540 | ~new_P1_U3077;
  assign new_P1_U5640 = ~new_P1_U3440 | ~new_P1_U3439;
  assign new_P1_U5641 = ~new_P1_U3052 | ~new_P1_U5640;
  assign new_P1_U5642 = ~new_P1_U3028 | ~new_P1_U3083;
  assign new_P1_U5643 = ~new_P1_U3485 | ~new_P1_U3438;
  assign new_P1_U5644 = ~new_P1_U5641 | ~new_P1_U3083;
  assign new_P1_U5645 = ~new_P1_U5786 | ~new_P1_U3084;
  assign new_P1_U5646 = ~new_P1_U3028 | ~new_P1_U3084;
  assign new_P1_U5647 = ~new_P1_U3482 | ~new_P1_U3438;
  assign new_P1_U5648 = ~new_P1_U5641 | ~new_P1_U3084;
  assign new_P1_U5649 = ~new_P1_U5786 | ~new_P1_U3070;
  assign new_P1_U5650 = ~new_P1_U3028 | ~new_P1_U3070;
  assign new_P1_U5651 = ~new_P1_U3479 | ~new_P1_U3438;
  assign new_P1_U5652 = ~new_P1_U5641 | ~new_P1_U3070;
  assign new_P1_U5653 = ~new_P1_U5786 | ~new_P1_U3071;
  assign new_P1_U5654 = ~new_P1_U3028 | ~new_P1_U3071;
  assign new_P1_U5655 = ~new_P1_U3476 | ~new_P1_U3438;
  assign new_P1_U5656 = ~new_P1_U5641 | ~new_P1_U3071;
  assign new_P1_U5657 = ~new_P1_U5786 | ~new_P1_U3067;
  assign new_P1_U5658 = ~new_P1_U3028 | ~new_P1_U3067;
  assign new_P1_U5659 = ~new_P1_U3473 | ~new_P1_U3438;
  assign new_P1_U5660 = ~new_P1_U5641 | ~new_P1_U3067;
  assign new_P1_U5661 = ~new_P1_U5786 | ~new_P1_U3060;
  assign new_P1_U5662 = ~new_P1_U3028 | ~new_P1_U3060;
  assign new_P1_U5663 = ~new_P1_U3470 | ~new_P1_U3438;
  assign new_P1_U5664 = ~new_P1_U5641 | ~new_P1_U3060;
  assign new_P1_U5665 = ~new_P1_U5786 | ~new_P1_U3064;
  assign new_P1_U5666 = ~new_P1_U3028 | ~new_P1_R1309_U8;
  assign new_P1_U5667 = ~new_P1_U4026 | ~new_P1_U3438;
  assign new_P1_U5668 = ~new_P1_U5641 | ~new_P1_U3056;
  assign new_P1_U5669 = ~new_P1_U3028 | ~new_P1_R1309_U6;
  assign new_P1_U5670 = ~new_P1_U4027 | ~new_P1_U3438;
  assign new_P1_U5671 = ~new_P1_U5641 | ~new_P1_U3059;
  assign new_P1_U5672 = ~new_P1_U3028 | ~new_P1_U3064;
  assign new_P1_U5673 = ~new_P1_U3467 | ~new_P1_U3438;
  assign new_P1_U5674 = ~new_P1_U5641 | ~new_P1_U3064;
  assign new_P1_U5675 = ~new_P1_U5786 | ~new_P1_U3068;
  assign new_P1_U5676 = ~new_P1_U3028 | ~new_P1_U3055;
  assign new_P1_U5677 = ~new_P1_U4028 | ~new_P1_U3438;
  assign new_P1_U5678 = ~new_P1_U5641 | ~new_P1_U3055;
  assign new_P1_U5679 = ~new_P1_U5786 | ~new_P1_U3054;
  assign new_P1_U5680 = ~new_P1_U3028 | ~new_P1_U3054;
  assign new_P1_U5681 = ~new_P1_U4017 | ~new_P1_U3438;
  assign new_P1_U5682 = ~new_P1_U5641 | ~new_P1_U3054;
  assign new_P1_U5683 = ~new_P1_U5786 | ~new_P1_U3053;
  assign new_P1_U5684 = ~new_P1_U3028 | ~new_P1_U3053;
  assign new_P1_U5685 = ~new_P1_U4018 | ~new_P1_U3438;
  assign new_P1_U5686 = ~new_P1_U5641 | ~new_P1_U3053;
  assign new_P1_U5687 = ~new_P1_U5786 | ~new_P1_U3057;
  assign new_P1_U5688 = ~new_P1_U3028 | ~new_P1_U3057;
  assign new_P1_U5689 = ~new_P1_U4019 | ~new_P1_U3438;
  assign new_P1_U5690 = ~new_P1_U5641 | ~new_P1_U3057;
  assign new_P1_U5691 = ~new_P1_U5786 | ~new_P1_U3058;
  assign new_P1_U5692 = ~new_P1_U3028 | ~new_P1_U3058;
  assign new_P1_U5693 = ~new_P1_U4020 | ~new_P1_U3438;
  assign new_P1_U5694 = ~new_P1_U5641 | ~new_P1_U3058;
  assign new_P1_U5695 = ~new_P1_U5786 | ~new_P1_U3065;
  assign new_P1_U5696 = ~new_P1_U3028 | ~new_P1_U3065;
  assign new_P1_U5697 = ~new_P1_U4021 | ~new_P1_U3438;
  assign new_P1_U5698 = ~new_P1_U5641 | ~new_P1_U3065;
  assign new_P1_U5699 = ~new_P1_U5786 | ~new_P1_U3066;
  assign new_P1_U5700 = ~new_P1_U3028 | ~new_P1_U3066;
  assign new_P1_U5701 = ~new_P1_U4022 | ~new_P1_U3438;
  assign new_P1_U5702 = ~new_P1_U5641 | ~new_P1_U3066;
  assign new_P1_U5703 = ~new_P1_U5786 | ~new_P1_U3061;
  assign new_P1_U5704 = ~new_P1_U3028 | ~new_P1_U3061;
  assign new_P1_U5705 = ~new_P1_U4023 | ~new_P1_U3438;
  assign new_P1_U5706 = ~new_P1_U5641 | ~new_P1_U3061;
  assign new_P1_U5707 = ~new_P1_U5786 | ~new_P1_U3075;
  assign new_P1_U5708 = ~new_P1_U3028 | ~new_P1_U3075;
  assign new_P1_U5709 = ~new_P1_U4024 | ~new_P1_U3438;
  assign new_P1_U5710 = ~new_P1_U5641 | ~new_P1_U3075;
  assign new_P1_U5711 = ~new_P1_U5786 | ~new_P1_U3076;
  assign new_P1_U5712 = ~new_P1_U3028 | ~new_P1_U3076;
  assign new_P1_U5713 = ~new_P1_U4025 | ~new_P1_U3438;
  assign new_P1_U5714 = ~new_P1_U5641 | ~new_P1_U3076;
  assign new_P1_U5715 = ~new_P1_U5786 | ~new_P1_U3081;
  assign new_P1_U5716 = ~new_P1_U3028 | ~new_P1_U3068;
  assign new_P1_U5717 = ~new_P1_U3464 | ~new_P1_U3438;
  assign new_P1_U5718 = ~new_P1_U5641 | ~new_P1_U3068;
  assign new_P1_U5719 = ~new_P1_U5786 | ~new_P1_U3078;
  assign new_P1_U5720 = ~new_P1_U3028 | ~new_P1_U3081;
  assign new_P1_U5721 = ~new_P1_U3514 | ~new_P1_U3438;
  assign new_P1_U5722 = ~new_P1_U5641 | ~new_P1_U3081;
  assign new_P1_U5723 = ~new_P1_U5786 | ~new_P1_U3082;
  assign new_P1_U5724 = ~new_P1_U3028 | ~new_P1_U3082;
  assign new_P1_U5725 = ~new_P1_U3512 | ~new_P1_U3438;
  assign new_P1_U5726 = ~new_P1_U5641 | ~new_P1_U3082;
  assign new_P1_U5727 = ~new_P1_U5786 | ~new_P1_U3069;
  assign new_P1_U5728 = ~new_P1_U3028 | ~new_P1_U3069;
  assign new_P1_U5729 = ~new_P1_U3509 | ~new_P1_U3438;
  assign new_P1_U5730 = ~new_P1_U5641 | ~new_P1_U3069;
  assign new_P1_U5731 = ~new_P1_U5786 | ~new_P1_U3073;
  assign new_P1_U5732 = ~new_P1_U3028 | ~new_P1_U3073;
  assign new_P1_U5733 = ~new_P1_U3506 | ~new_P1_U3438;
  assign new_P1_U5734 = ~new_P1_U5641 | ~new_P1_U3073;
  assign new_P1_U5735 = ~new_P1_U5786 | ~new_P1_U3074;
  assign new_P1_U5736 = ~new_P1_U3028 | ~new_P1_U3074;
  assign new_P1_U5737 = ~new_P1_U3503 | ~new_P1_U3438;
  assign new_P1_U5738 = ~new_P1_U5641 | ~new_P1_U3074;
  assign new_P1_U5739 = ~new_P1_U5786 | ~new_P1_U3079;
  assign new_P1_U5740 = ~new_P1_U3028 | ~new_P1_U3079;
  assign new_P1_U5741 = ~new_P1_U3500 | ~new_P1_U3438;
  assign new_P1_U5742 = ~new_P1_U5641 | ~new_P1_U3079;
  assign new_P1_U5743 = ~new_P1_U5786 | ~new_P1_U3080;
  assign new_P1_U5744 = ~new_P1_U3028 | ~new_P1_U3080;
  assign new_P1_U5745 = ~new_P1_U3497 | ~new_P1_U3438;
  assign new_P1_U5746 = ~new_P1_U5641 | ~new_P1_U3080;
  assign new_P1_U5747 = ~new_P1_U5786 | ~new_P1_U3072;
  assign new_P1_U5748 = ~new_P1_U3028 | ~new_P1_U3072;
  assign new_P1_U5749 = ~new_P1_U3494 | ~new_P1_U3438;
  assign new_P1_U5750 = ~new_P1_U5641 | ~new_P1_U3072;
  assign new_P1_U5751 = ~new_P1_U5786 | ~new_P1_U3063;
  assign new_P1_U5752 = ~new_P1_U3028 | ~new_P1_U3063;
  assign new_P1_U5753 = ~new_P1_U3491 | ~new_P1_U3438;
  assign new_P1_U5754 = ~new_P1_U5641 | ~new_P1_U3063;
  assign new_P1_U5755 = ~new_P1_U5786 | ~new_P1_U3062;
  assign new_P1_U5756 = ~new_P1_U3028 | ~new_P1_U3062;
  assign new_P1_U5757 = ~new_P1_U3488 | ~new_P1_U3438;
  assign new_P1_U5758 = ~new_P1_U5641 | ~new_P1_U3062;
  assign new_P1_U5759 = ~new_P1_U5786 | ~new_P1_U3083;
  assign new_P1_U5760 = ~new_P1_U3028 | ~new_P1_U3078;
  assign new_P1_U5761 = ~new_P1_U3461 | ~new_P1_U3438;
  assign new_P1_U5762 = ~new_P1_U5641 | ~new_P1_U3078;
  assign new_P1_U5763 = ~new_P1_U5786 | ~new_P1_U3077;
  assign new_P1_U5764 = ~new_P1_U3028 | ~new_P1_U3077;
  assign new_P1_U5765 = ~new_P1_U3456 | ~new_P1_U3438;
  assign new_P1_U5766 = ~new_P1_U5641 | ~new_P1_U3077;
  assign new_P1_U5767 = ~new_P1_U4038 | ~new_P1_U3434;
  assign new_P1_U5768 = ~new_P1_U4015 | ~new_P1_U4038;
  assign new_P1_U5769 = ~new_P1_U3050 | ~new_P1_U5767;
  assign new_P1_U5770 = ~new_P1_U5768 | ~new_P1_U4039;
  assign new_P1_U5771 = ~new_P1_U5775 | ~new_P1_U5781;
  assign new_P1_U5772 = ~new_P1_R1375_U9 | ~new_P1_U5131;
  assign new_P1_U5773 = ~P1_IR_REG_24_ | ~new_P1_U3952;
  assign new_P1_U5774 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U17;
  assign new_P1_U5775 = ~new_P1_U3441;
  assign new_P1_U5776 = ~P1_IR_REG_25_ | ~new_P1_U3952;
  assign new_P1_U5777 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U170;
  assign new_P1_U5778 = ~new_P1_U3442;
  assign new_P1_U5779 = ~P1_IR_REG_26_ | ~new_P1_U3952;
  assign new_P1_U5780 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U18;
  assign new_P1_U5781 = ~new_P1_U3443;
  assign new_P1_U5782 = ~new_P1_U3441 | ~new_P1_U3359;
  assign new_P1_U5783 = ~P1_B_REG | ~new_P1_U4046 | ~new_P1_U5775;
  assign new_P1_U5784 = ~P1_IR_REG_23_ | ~new_P1_U3952;
  assign new_P1_U5785 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U16;
  assign new_P1_U5786 = ~new_P1_U3444;
  assign new_P1_U5787 = ~P1_D_REG_0_ | ~new_P1_U3953;
  assign new_P1_U5788 = ~new_P1_U4034 | ~new_P1_U4146;
  assign new_P1_U5789 = ~P1_D_REG_1_ | ~new_P1_U3953;
  assign new_P1_U5790 = ~new_P1_U4034 | ~new_P1_U4147;
  assign new_P1_U5791 = ~P1_IR_REG_22_ | ~new_P1_U3952;
  assign new_P1_U5792 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U15;
  assign new_P1_U5793 = ~new_P1_U3451;
  assign new_P1_U5794 = ~P1_IR_REG_19_ | ~new_P1_U3952;
  assign new_P1_U5795 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U13;
  assign new_P1_U5796 = ~new_P1_U3452;
  assign new_P1_U5797 = ~P1_IR_REG_20_ | ~new_P1_U3952;
  assign new_P1_U5798 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U14;
  assign new_P1_U5799 = ~new_P1_U3453;
  assign new_P1_U5800 = ~P1_IR_REG_21_ | ~new_P1_U3952;
  assign new_P1_U5801 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U173;
  assign new_P1_U5802 = ~new_P1_U3450;
  assign new_P1_U5803 = ~P1_IR_REG_30_ | ~new_P1_U3952;
  assign new_P1_U5804 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U165;
  assign new_P1_U5805 = ~new_P1_U3447;
  assign new_P1_U5806 = ~P1_IR_REG_29_ | ~new_P1_U3952;
  assign new_P1_U5807 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U20;
  assign new_P1_U5808 = ~new_P1_U3448;
  assign new_P1_U5809 = ~P1_IR_REG_28_ | ~new_P1_U3952;
  assign new_P1_U5810 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U19;
  assign new_P1_U5811 = ~new_P1_U3449;
  assign new_P1_U5812 = ~P1_IR_REG_0_ | ~new_P1_U3952;
  assign new_P1_U5813 = ~P1_IR_REG_31_ | ~P1_IR_REG_0_;
  assign new_P1_U5814 = ~new_P1_U3454;
  assign new_P1_U5815 = ~P1_IR_REG_27_ | ~new_P1_U3952;
  assign new_P1_U5816 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U42;
  assign new_P1_U5817 = ~new_P1_U3455;
  assign new_P1_U5818 = ~new_U125 | ~new_P1_U3954;
  assign new_P1_U5819 = ~new_P1_U4014 | ~new_P1_U3454;
  assign new_P1_U5820 = ~new_P1_U3456;
  assign new_P1_U5821 = ~new_P1_U3451 | ~new_P1_U5802;
  assign new_P1_U5822 = ~new_P1_U5793 | ~new_P1_U4178;
  assign new_P1_U5823 = ~P1_D_REG_1_ | ~new_P1_U4144;
  assign new_P1_U5824 = ~new_P1_U4147 | ~new_P1_U3360;
  assign new_P1_U5825 = ~new_P1_U3458;
  assign new_P1_U5826 = ~new_P1_U5771 | ~new_P1_U3360;
  assign new_P1_U5827 = ~P1_D_REG_0_ | ~new_P1_U4144;
  assign new_P1_U5828 = ~new_P1_U3457;
  assign new_P1_U5829 = ~P1_REG0_REG_0_ | ~new_P1_U3955;
  assign new_P1_U5830 = ~new_P1_U4033 | ~new_P1_U4198;
  assign new_P1_U5831 = ~P1_IR_REG_1_ | ~new_P1_U3952;
  assign new_P1_U5832 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U40;
  assign new_P1_U5833 = ~new_U114 | ~new_P1_U3954;
  assign new_P1_U5834 = ~new_P1_U3460 | ~new_P1_U4014;
  assign new_P1_U5835 = ~new_P1_U3461;
  assign new_P1_U5836 = ~P1_REG0_REG_1_ | ~new_P1_U3955;
  assign new_P1_U5837 = ~new_P1_U4033 | ~new_P1_U4222;
  assign new_P1_U5838 = ~P1_IR_REG_2_ | ~new_P1_U3952;
  assign new_P1_U5839 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U21;
  assign new_P1_U5840 = ~new_U103 | ~new_P1_U3954;
  assign new_P1_U5841 = ~new_P1_U3463 | ~new_P1_U4014;
  assign new_P1_U5842 = ~new_P1_U3464;
  assign new_P1_U5843 = ~P1_REG0_REG_2_ | ~new_P1_U3955;
  assign new_P1_U5844 = ~new_P1_U4033 | ~new_P1_U4241;
  assign new_P1_U5845 = ~P1_IR_REG_3_ | ~new_P1_U3952;
  assign new_P1_U5846 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U22;
  assign new_P1_U5847 = ~new_U100 | ~new_P1_U3954;
  assign new_P1_U5848 = ~new_P1_U3466 | ~new_P1_U4014;
  assign new_P1_U5849 = ~new_P1_U3467;
  assign new_P1_U5850 = ~P1_REG0_REG_3_ | ~new_P1_U3955;
  assign new_P1_U5851 = ~new_P1_U4033 | ~new_P1_U4260;
  assign new_P1_U5852 = ~P1_IR_REG_4_ | ~new_P1_U3952;
  assign new_P1_U5853 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U23;
  assign new_P1_U5854 = ~new_U99 | ~new_P1_U3954;
  assign new_P1_U5855 = ~new_P1_U3469 | ~new_P1_U4014;
  assign new_P1_U5856 = ~new_P1_U3470;
  assign new_P1_U5857 = ~P1_REG0_REG_4_ | ~new_P1_U3955;
  assign new_P1_U5858 = ~new_P1_U4033 | ~new_P1_U4279;
  assign new_P1_U5859 = ~P1_IR_REG_5_ | ~new_P1_U3952;
  assign new_P1_U5860 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U162;
  assign new_P1_U5861 = ~new_U98 | ~new_P1_U3954;
  assign new_P1_U5862 = ~new_P1_U3472 | ~new_P1_U4014;
  assign new_P1_U5863 = ~new_P1_U3473;
  assign new_P1_U5864 = ~P1_REG0_REG_5_ | ~new_P1_U3955;
  assign new_P1_U5865 = ~new_P1_U4033 | ~new_P1_U4298;
  assign new_P1_U5866 = ~P1_IR_REG_6_ | ~new_P1_U3952;
  assign new_P1_U5867 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U24;
  assign new_P1_U5868 = ~new_U97 | ~new_P1_U3954;
  assign new_P1_U5869 = ~new_P1_U3475 | ~new_P1_U4014;
  assign new_P1_U5870 = ~new_P1_U3476;
  assign new_P1_U5871 = ~P1_REG0_REG_6_ | ~new_P1_U3955;
  assign new_P1_U5872 = ~new_P1_U4033 | ~new_P1_U4317;
  assign new_P1_U5873 = ~P1_IR_REG_7_ | ~new_P1_U3952;
  assign new_P1_U5874 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U25;
  assign new_P1_U5875 = ~new_U96 | ~new_P1_U3954;
  assign new_P1_U5876 = ~new_P1_U3478 | ~new_P1_U4014;
  assign new_P1_U5877 = ~new_P1_U3479;
  assign new_P1_U5878 = ~P1_REG0_REG_7_ | ~new_P1_U3955;
  assign new_P1_U5879 = ~new_P1_U4033 | ~new_P1_U4336;
  assign new_P1_U5880 = ~P1_IR_REG_8_ | ~new_P1_U3952;
  assign new_P1_U5881 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U26;
  assign new_P1_U5882 = ~new_U95 | ~new_P1_U3954;
  assign new_P1_U5883 = ~new_P1_U3481 | ~new_P1_U4014;
  assign new_P1_U5884 = ~new_P1_U3482;
  assign new_P1_U5885 = ~P1_REG0_REG_8_ | ~new_P1_U3955;
  assign new_P1_U5886 = ~new_P1_U4033 | ~new_P1_U4355;
  assign new_P1_U5887 = ~P1_IR_REG_9_ | ~new_P1_U3952;
  assign new_P1_U5888 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U160;
  assign new_P1_U5889 = ~new_U94 | ~new_P1_U3954;
  assign new_P1_U5890 = ~new_P1_U3484 | ~new_P1_U4014;
  assign new_P1_U5891 = ~new_P1_U3485;
  assign new_P1_U5892 = ~P1_REG0_REG_9_ | ~new_P1_U3955;
  assign new_P1_U5893 = ~new_P1_U4033 | ~new_P1_U4374;
  assign new_P1_U5894 = ~P1_IR_REG_10_ | ~new_P1_U3952;
  assign new_P1_U5895 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U6;
  assign new_P1_U5896 = ~new_U124 | ~new_P1_U3954;
  assign new_P1_U5897 = ~new_P1_U3487 | ~new_P1_U4014;
  assign new_P1_U5898 = ~new_P1_U3488;
  assign new_P1_U5899 = ~P1_REG0_REG_10_ | ~new_P1_U3955;
  assign new_P1_U5900 = ~new_P1_U4033 | ~new_P1_U4393;
  assign new_P1_U5901 = ~P1_IR_REG_11_ | ~new_P1_U3952;
  assign new_P1_U5902 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U7;
  assign new_P1_U5903 = ~new_U123 | ~new_P1_U3954;
  assign new_P1_U5904 = ~new_P1_U3490 | ~new_P1_U4014;
  assign new_P1_U5905 = ~new_P1_U3491;
  assign new_P1_U5906 = ~P1_REG0_REG_11_ | ~new_P1_U3955;
  assign new_P1_U5907 = ~new_P1_U4033 | ~new_P1_U4412;
  assign new_P1_U5908 = ~P1_IR_REG_12_ | ~new_P1_U3952;
  assign new_P1_U5909 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U8;
  assign new_P1_U5910 = ~new_U122 | ~new_P1_U3954;
  assign new_P1_U5911 = ~new_P1_U3493 | ~new_P1_U4014;
  assign new_P1_U5912 = ~new_P1_U3494;
  assign new_P1_U5913 = ~P1_REG0_REG_12_ | ~new_P1_U3955;
  assign new_P1_U5914 = ~new_P1_U4033 | ~new_P1_U4431;
  assign new_P1_U5915 = ~P1_IR_REG_13_ | ~new_P1_U3952;
  assign new_P1_U5916 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U179;
  assign new_P1_U5917 = ~new_U121 | ~new_P1_U3954;
  assign new_P1_U5918 = ~new_P1_U3496 | ~new_P1_U4014;
  assign new_P1_U5919 = ~new_P1_U3497;
  assign new_P1_U5920 = ~P1_REG0_REG_13_ | ~new_P1_U3955;
  assign new_P1_U5921 = ~new_P1_U4033 | ~new_P1_U4450;
  assign new_P1_U5922 = ~P1_IR_REG_14_ | ~new_P1_U3952;
  assign new_P1_U5923 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U9;
  assign new_P1_U5924 = ~new_U120 | ~new_P1_U3954;
  assign new_P1_U5925 = ~new_P1_U3499 | ~new_P1_U4014;
  assign new_P1_U5926 = ~new_P1_U3500;
  assign new_P1_U5927 = ~P1_REG0_REG_14_ | ~new_P1_U3955;
  assign new_P1_U5928 = ~new_P1_U4033 | ~new_P1_U4469;
  assign new_P1_U5929 = ~P1_IR_REG_15_ | ~new_P1_U3952;
  assign new_P1_U5930 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U10;
  assign new_P1_U5931 = ~new_U119 | ~new_P1_U3954;
  assign new_P1_U5932 = ~new_P1_U3502 | ~new_P1_U4014;
  assign new_P1_U5933 = ~new_P1_U3503;
  assign new_P1_U5934 = ~P1_REG0_REG_15_ | ~new_P1_U3955;
  assign new_P1_U5935 = ~new_P1_U4033 | ~new_P1_U4488;
  assign new_P1_U5936 = ~P1_IR_REG_16_ | ~new_P1_U3952;
  assign new_P1_U5937 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U11;
  assign new_P1_U5938 = ~new_U118 | ~new_P1_U3954;
  assign new_P1_U5939 = ~new_P1_U3505 | ~new_P1_U4014;
  assign new_P1_U5940 = ~new_P1_U3506;
  assign new_P1_U5941 = ~P1_REG0_REG_16_ | ~new_P1_U3955;
  assign new_P1_U5942 = ~new_P1_U4033 | ~new_P1_U4507;
  assign new_P1_U5943 = ~P1_IR_REG_17_ | ~new_P1_U3952;
  assign new_P1_U5944 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U177;
  assign new_P1_U5945 = ~new_U117 | ~new_P1_U3954;
  assign new_P1_U5946 = ~new_P1_U3508 | ~new_P1_U4014;
  assign new_P1_U5947 = ~new_P1_U3509;
  assign new_P1_U5948 = ~P1_REG0_REG_17_ | ~new_P1_U3955;
  assign new_P1_U5949 = ~new_P1_U4033 | ~new_P1_U4526;
  assign new_P1_U5950 = ~P1_IR_REG_18_ | ~new_P1_U3952;
  assign new_P1_U5951 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U12;
  assign new_P1_U5952 = ~new_U116 | ~new_P1_U3954;
  assign new_P1_U5953 = ~new_P1_U3511 | ~new_P1_U4014;
  assign new_P1_U5954 = ~new_P1_U3512;
  assign new_P1_U5955 = ~P1_REG0_REG_18_ | ~new_P1_U3955;
  assign new_P1_U5956 = ~new_P1_U4033 | ~new_P1_U4545;
  assign new_P1_U5957 = ~new_U115 | ~new_P1_U3954;
  assign new_P1_U5958 = ~new_P1_U4014 | ~new_P1_U3452;
  assign new_P1_U5959 = ~new_P1_U3514;
  assign new_P1_U5960 = ~P1_REG0_REG_19_ | ~new_P1_U3955;
  assign new_P1_U5961 = ~new_P1_U4033 | ~new_P1_U4564;
  assign new_P1_U5962 = ~P1_REG0_REG_20_ | ~new_P1_U3955;
  assign new_P1_U5963 = ~new_P1_U4033 | ~new_P1_U4583;
  assign new_P1_U5964 = ~P1_REG0_REG_21_ | ~new_P1_U3955;
  assign new_P1_U5965 = ~new_P1_U4033 | ~new_P1_U4602;
  assign new_P1_U5966 = ~P1_REG0_REG_22_ | ~new_P1_U3955;
  assign new_P1_U5967 = ~new_P1_U4033 | ~new_P1_U4621;
  assign new_P1_U5968 = ~P1_REG0_REG_23_ | ~new_P1_U3955;
  assign new_P1_U5969 = ~new_P1_U4033 | ~new_P1_U4640;
  assign new_P1_U5970 = ~P1_REG0_REG_24_ | ~new_P1_U3955;
  assign new_P1_U5971 = ~new_P1_U4033 | ~new_P1_U4659;
  assign new_P1_U5972 = ~P1_REG0_REG_25_ | ~new_P1_U3955;
  assign new_P1_U5973 = ~new_P1_U4033 | ~new_P1_U4678;
  assign new_P1_U5974 = ~P1_REG0_REG_26_ | ~new_P1_U3955;
  assign new_P1_U5975 = ~new_P1_U4033 | ~new_P1_U4697;
  assign new_P1_U5976 = ~P1_REG0_REG_27_ | ~new_P1_U3955;
  assign new_P1_U5977 = ~new_P1_U4033 | ~new_P1_U4716;
  assign new_P1_U5978 = ~P1_REG0_REG_28_ | ~new_P1_U3955;
  assign new_P1_U5979 = ~new_P1_U4033 | ~new_P1_U4735;
  assign new_P1_U5980 = ~P1_REG0_REG_29_ | ~new_P1_U3955;
  assign new_P1_U5981 = ~new_P1_U4033 | ~new_P1_U4755;
  assign new_P1_U5982 = ~P1_REG0_REG_30_ | ~new_P1_U3955;
  assign new_P1_U5983 = ~new_P1_U4033 | ~new_P1_U4762;
  assign new_P1_U5984 = ~P1_REG0_REG_31_ | ~new_P1_U3955;
  assign new_P1_U5985 = ~new_P1_U4033 | ~new_P1_U4765;
  assign new_P1_U5986 = ~P1_REG1_REG_0_ | ~new_P1_U3956;
  assign new_P1_U5987 = ~new_P1_U4032 | ~new_P1_U4198;
  assign new_P1_U5988 = ~P1_REG1_REG_1_ | ~new_P1_U3956;
  assign new_P1_U5989 = ~new_P1_U4032 | ~new_P1_U4222;
  assign new_P1_U5990 = ~P1_REG1_REG_2_ | ~new_P1_U3956;
  assign new_P1_U5991 = ~new_P1_U4032 | ~new_P1_U4241;
  assign new_P1_U5992 = ~P1_REG1_REG_3_ | ~new_P1_U3956;
  assign new_P1_U5993 = ~new_P1_U4032 | ~new_P1_U4260;
  assign new_P1_U5994 = ~P1_REG1_REG_4_ | ~new_P1_U3956;
  assign new_P1_U5995 = ~new_P1_U4032 | ~new_P1_U4279;
  assign new_P1_U5996 = ~P1_REG1_REG_5_ | ~new_P1_U3956;
  assign new_P1_U5997 = ~new_P1_U4032 | ~new_P1_U4298;
  assign new_P1_U5998 = ~P1_REG1_REG_6_ | ~new_P1_U3956;
  assign new_P1_U5999 = ~new_P1_U4032 | ~new_P1_U4317;
  assign new_P1_U6000 = ~P1_REG1_REG_7_ | ~new_P1_U3956;
  assign new_P1_U6001 = ~new_P1_U4032 | ~new_P1_U4336;
  assign new_P1_U6002 = ~P1_REG1_REG_8_ | ~new_P1_U3956;
  assign new_P1_U6003 = ~new_P1_U4032 | ~new_P1_U4355;
  assign new_P1_U6004 = ~P1_REG1_REG_9_ | ~new_P1_U3956;
  assign new_P1_U6005 = ~new_P1_U4032 | ~new_P1_U4374;
  assign new_P1_U6006 = ~P1_REG1_REG_10_ | ~new_P1_U3956;
  assign new_P1_U6007 = ~new_P1_U4032 | ~new_P1_U4393;
  assign new_P1_U6008 = ~P1_REG1_REG_11_ | ~new_P1_U3956;
  assign new_P1_U6009 = ~new_P1_U4032 | ~new_P1_U4412;
  assign new_P1_U6010 = ~P1_REG1_REG_12_ | ~new_P1_U3956;
  assign new_P1_U6011 = ~new_P1_U4032 | ~new_P1_U4431;
  assign new_P1_U6012 = ~P1_REG1_REG_13_ | ~new_P1_U3956;
  assign new_P1_U6013 = ~new_P1_U4032 | ~new_P1_U4450;
  assign new_P1_U6014 = ~P1_REG1_REG_14_ | ~new_P1_U3956;
  assign new_P1_U6015 = ~new_P1_U4032 | ~new_P1_U4469;
  assign new_P1_U6016 = ~P1_REG1_REG_15_ | ~new_P1_U3956;
  assign new_P1_U6017 = ~new_P1_U4032 | ~new_P1_U4488;
  assign new_P1_U6018 = ~P1_REG1_REG_16_ | ~new_P1_U3956;
  assign new_P1_U6019 = ~new_P1_U4032 | ~new_P1_U4507;
  assign new_P1_U6020 = ~P1_REG1_REG_17_ | ~new_P1_U3956;
  assign new_P1_U6021 = ~new_P1_U4032 | ~new_P1_U4526;
  assign new_P1_U6022 = ~P1_REG1_REG_18_ | ~new_P1_U3956;
  assign new_P1_U6023 = ~new_P1_U4032 | ~new_P1_U4545;
  assign new_P1_U6024 = ~P1_REG1_REG_19_ | ~new_P1_U3956;
  assign new_P1_U6025 = ~new_P1_U4032 | ~new_P1_U4564;
  assign new_P1_U6026 = ~P1_REG1_REG_20_ | ~new_P1_U3956;
  assign new_P1_U6027 = ~new_P1_U4032 | ~new_P1_U4583;
  assign new_P1_U6028 = ~P1_REG1_REG_21_ | ~new_P1_U3956;
  assign new_P1_U6029 = ~new_P1_U4032 | ~new_P1_U4602;
  assign new_P1_U6030 = ~P1_REG1_REG_22_ | ~new_P1_U3956;
  assign new_P1_U6031 = ~new_P1_U4032 | ~new_P1_U4621;
  assign new_P1_U6032 = ~P1_REG1_REG_23_ | ~new_P1_U3956;
  assign new_P1_U6033 = ~new_P1_U4032 | ~new_P1_U4640;
  assign new_P1_U6034 = ~P1_REG1_REG_24_ | ~new_P1_U3956;
  assign new_P1_U6035 = ~new_P1_U4032 | ~new_P1_U4659;
  assign new_P1_U6036 = ~P1_REG1_REG_25_ | ~new_P1_U3956;
  assign new_P1_U6037 = ~new_P1_U4032 | ~new_P1_U4678;
  assign new_P1_U6038 = ~P1_REG1_REG_26_ | ~new_P1_U3956;
  assign new_P1_U6039 = ~new_P1_U4032 | ~new_P1_U4697;
  assign new_P1_U6040 = ~P1_REG1_REG_27_ | ~new_P1_U3956;
  assign new_P1_U6041 = ~new_P1_U4032 | ~new_P1_U4716;
  assign new_P1_U6042 = ~P1_REG1_REG_28_ | ~new_P1_U3956;
  assign new_P1_U6043 = ~new_P1_U4032 | ~new_P1_U4735;
  assign new_P1_U6044 = ~P1_REG1_REG_29_ | ~new_P1_U3956;
  assign new_P1_U6045 = ~new_P1_U4032 | ~new_P1_U4755;
  assign new_P1_U6046 = ~P1_REG1_REG_30_ | ~new_P1_U3956;
  assign new_P1_U6047 = ~new_P1_U4032 | ~new_P1_U4762;
  assign new_P1_U6048 = ~P1_REG1_REG_31_ | ~new_P1_U3956;
  assign new_P1_U6049 = ~new_P1_U4032 | ~new_P1_U4765;
  assign new_P1_U6050 = ~P1_REG2_REG_0_ | ~new_P1_U3420;
  assign new_P1_U6051 = ~new_P1_U4031 | ~new_P1_U3376;
  assign new_P1_U6052 = ~P1_REG2_REG_1_ | ~new_P1_U3420;
  assign new_P1_U6053 = ~new_P1_U4031 | ~new_P1_U3378;
  assign new_P1_U6054 = ~P1_REG2_REG_2_ | ~new_P1_U3420;
  assign new_P1_U6055 = ~new_P1_U4031 | ~new_P1_U3379;
  assign new_P1_U6056 = ~P1_REG2_REG_3_ | ~new_P1_U3420;
  assign new_P1_U6057 = ~new_P1_U4031 | ~new_P1_U3380;
  assign new_P1_U6058 = ~P1_REG2_REG_4_ | ~new_P1_U3420;
  assign new_P1_U6059 = ~new_P1_U4031 | ~new_P1_U3381;
  assign new_P1_U6060 = ~P1_REG2_REG_5_ | ~new_P1_U3420;
  assign new_P1_U6061 = ~new_P1_U4031 | ~new_P1_U3382;
  assign new_P1_U6062 = ~P1_REG2_REG_6_ | ~new_P1_U3420;
  assign new_P1_U6063 = ~new_P1_U4031 | ~new_P1_U3383;
  assign new_P1_U6064 = ~P1_REG2_REG_7_ | ~new_P1_U3420;
  assign new_P1_U6065 = ~new_P1_U4031 | ~new_P1_U3384;
  assign new_P1_U6066 = ~P1_REG2_REG_8_ | ~new_P1_U3420;
  assign new_P1_U6067 = ~new_P1_U4031 | ~new_P1_U3385;
  assign new_P1_U6068 = ~P1_REG2_REG_9_ | ~new_P1_U3420;
  assign new_P1_U6069 = ~new_P1_U4031 | ~new_P1_U3386;
  assign new_P1_U6070 = ~P1_REG2_REG_10_ | ~new_P1_U3420;
  assign new_P1_U6071 = ~new_P1_U4031 | ~new_P1_U3387;
  assign new_P1_U6072 = ~P1_REG2_REG_11_ | ~new_P1_U3420;
  assign new_P1_U6073 = ~new_P1_U4031 | ~new_P1_U3388;
  assign new_P1_U6074 = ~P1_REG2_REG_12_ | ~new_P1_U3420;
  assign new_P1_U6075 = ~new_P1_U4031 | ~new_P1_U3389;
  assign new_P1_U6076 = ~P1_REG2_REG_13_ | ~new_P1_U3420;
  assign new_P1_U6077 = ~new_P1_U4031 | ~new_P1_U3390;
  assign new_P1_U6078 = ~P1_REG2_REG_14_ | ~new_P1_U3420;
  assign new_P1_U6079 = ~new_P1_U4031 | ~new_P1_U3391;
  assign new_P1_U6080 = ~P1_REG2_REG_15_ | ~new_P1_U3420;
  assign new_P1_U6081 = ~new_P1_U4031 | ~new_P1_U3392;
  assign new_P1_U6082 = ~P1_REG2_REG_16_ | ~new_P1_U3420;
  assign new_P1_U6083 = ~new_P1_U4031 | ~new_P1_U3393;
  assign new_P1_U6084 = ~P1_REG2_REG_17_ | ~new_P1_U3420;
  assign new_P1_U6085 = ~new_P1_U4031 | ~new_P1_U3394;
  assign new_P1_U6086 = ~P1_REG2_REG_18_ | ~new_P1_U3420;
  assign new_P1_U6087 = ~new_P1_U4031 | ~new_P1_U3395;
  assign new_P1_U6088 = ~P1_REG2_REG_19_ | ~new_P1_U3420;
  assign new_P1_U6089 = ~new_P1_U4031 | ~new_P1_U3396;
  assign new_P1_U6090 = ~P1_REG2_REG_20_ | ~new_P1_U3420;
  assign new_P1_U6091 = ~new_P1_U4031 | ~new_P1_U3398;
  assign new_P1_U6092 = ~P1_REG2_REG_21_ | ~new_P1_U3420;
  assign new_P1_U6093 = ~new_P1_U4031 | ~new_P1_U3400;
  assign new_P1_U6094 = ~P1_REG2_REG_22_ | ~new_P1_U3420;
  assign new_P1_U6095 = ~new_P1_U4031 | ~new_P1_U3402;
  assign new_P1_U6096 = ~P1_REG2_REG_23_ | ~new_P1_U3420;
  assign new_P1_U6097 = ~new_P1_U4031 | ~new_P1_U3404;
  assign new_P1_U6098 = ~P1_REG2_REG_24_ | ~new_P1_U3420;
  assign new_P1_U6099 = ~new_P1_U4031 | ~new_P1_U3406;
  assign new_P1_U6100 = ~P1_REG2_REG_25_ | ~new_P1_U3420;
  assign new_P1_U6101 = ~new_P1_U4031 | ~new_P1_U3408;
  assign new_P1_U6102 = ~P1_REG2_REG_26_ | ~new_P1_U3420;
  assign new_P1_U6103 = ~new_P1_U4031 | ~new_P1_U3410;
  assign new_P1_U6104 = ~P1_REG2_REG_27_ | ~new_P1_U3420;
  assign new_P1_U6105 = ~new_P1_U4031 | ~new_P1_U3412;
  assign new_P1_U6106 = ~P1_REG2_REG_28_ | ~new_P1_U3420;
  assign new_P1_U6107 = ~new_P1_U4031 | ~new_P1_U3414;
  assign new_P1_U6108 = ~P1_REG2_REG_29_ | ~new_P1_U3420;
  assign new_P1_U6109 = ~new_P1_U4031 | ~new_P1_U3416;
  assign new_P1_U6110 = ~P1_REG2_REG_30_ | ~new_P1_U3420;
  assign new_P1_U6111 = ~new_P1_U4035 | ~new_P1_U4031;
  assign new_P1_U6112 = ~P1_REG2_REG_31_ | ~new_P1_U3420;
  assign new_P1_U6113 = ~new_P1_U4035 | ~new_P1_U4031;
  assign new_P1_U6114 = ~P1_DATAO_REG_0_ | ~new_P1_U3430;
  assign new_P1_U6115 = ~n1394 | ~new_P1_U3077;
  assign new_P1_U6116 = ~P1_DATAO_REG_1_ | ~new_P1_U3430;
  assign new_P1_U6117 = ~n1394 | ~new_P1_U3078;
  assign new_P1_U6118 = ~P1_DATAO_REG_2_ | ~new_P1_U3430;
  assign new_P1_U6119 = ~n1394 | ~new_P1_U3068;
  assign new_P1_U6120 = ~P1_DATAO_REG_3_ | ~new_P1_U3430;
  assign new_P1_U6121 = ~n1394 | ~new_P1_U3064;
  assign new_P1_U6122 = ~P1_DATAO_REG_4_ | ~new_P1_U3430;
  assign new_P1_U6123 = ~n1394 | ~new_P1_U3060;
  assign new_P1_U6124 = ~P1_DATAO_REG_5_ | ~new_P1_U3430;
  assign new_P1_U6125 = ~n1394 | ~new_P1_U3067;
  assign new_P1_U6126 = ~P1_DATAO_REG_6_ | ~new_P1_U3430;
  assign new_P1_U6127 = ~n1394 | ~new_P1_U3071;
  assign new_P1_U6128 = ~P1_DATAO_REG_7_ | ~new_P1_U3430;
  assign new_P1_U6129 = ~n1394 | ~new_P1_U3070;
  assign new_P1_U6130 = ~P1_DATAO_REG_8_ | ~new_P1_U3430;
  assign new_P1_U6131 = ~n1394 | ~new_P1_U3084;
  assign new_P1_U6132 = ~P1_DATAO_REG_9_ | ~new_P1_U3430;
  assign new_P1_U6133 = ~n1394 | ~new_P1_U3083;
  assign new_P1_U6134 = ~P1_DATAO_REG_10_ | ~new_P1_U3430;
  assign new_P1_U6135 = ~n1394 | ~new_P1_U3062;
  assign new_P1_U6136 = ~P1_DATAO_REG_11_ | ~new_P1_U3430;
  assign new_P1_U6137 = ~n1394 | ~new_P1_U3063;
  assign new_P1_U6138 = ~P1_DATAO_REG_12_ | ~new_P1_U3430;
  assign new_P1_U6139 = ~n1394 | ~new_P1_U3072;
  assign new_P1_U6140 = ~P1_DATAO_REG_13_ | ~new_P1_U3430;
  assign new_P1_U6141 = ~n1394 | ~new_P1_U3080;
  assign new_P1_U6142 = ~P1_DATAO_REG_14_ | ~new_P1_U3430;
  assign new_P1_U6143 = ~n1394 | ~new_P1_U3079;
  assign new_P1_U6144 = ~P1_DATAO_REG_15_ | ~new_P1_U3430;
  assign new_P1_U6145 = ~n1394 | ~new_P1_U3074;
  assign new_P1_U6146 = ~P1_DATAO_REG_16_ | ~new_P1_U3430;
  assign new_P1_U6147 = ~n1394 | ~new_P1_U3073;
  assign new_P1_U6148 = ~P1_DATAO_REG_17_ | ~new_P1_U3430;
  assign new_P1_U6149 = ~n1394 | ~new_P1_U3069;
  assign new_P1_U6150 = ~P1_DATAO_REG_18_ | ~new_P1_U3430;
  assign new_P1_U6151 = ~n1394 | ~new_P1_U3082;
  assign new_P1_U6152 = ~P1_DATAO_REG_19_ | ~new_P1_U3430;
  assign new_P1_U6153 = ~n1394 | ~new_P1_U3081;
  assign new_P1_U6154 = ~P1_DATAO_REG_20_ | ~new_P1_U3430;
  assign new_P1_U6155 = ~n1394 | ~new_P1_U3076;
  assign new_P1_U6156 = ~P1_DATAO_REG_21_ | ~new_P1_U3430;
  assign new_P1_U6157 = ~n1394 | ~new_P1_U3075;
  assign new_P1_U6158 = ~P1_DATAO_REG_22_ | ~new_P1_U3430;
  assign new_P1_U6159 = ~n1394 | ~new_P1_U3061;
  assign new_P1_U6160 = ~P1_DATAO_REG_23_ | ~new_P1_U3430;
  assign new_P1_U6161 = ~n1394 | ~new_P1_U3066;
  assign new_P1_U6162 = ~P1_DATAO_REG_24_ | ~new_P1_U3430;
  assign new_P1_U6163 = ~n1394 | ~new_P1_U3065;
  assign new_P1_U6164 = ~P1_DATAO_REG_25_ | ~new_P1_U3430;
  assign new_P1_U6165 = ~n1394 | ~new_P1_U3058;
  assign new_P1_U6166 = ~P1_DATAO_REG_26_ | ~new_P1_U3430;
  assign new_P1_U6167 = ~n1394 | ~new_P1_U3057;
  assign new_P1_U6168 = ~P1_DATAO_REG_27_ | ~new_P1_U3430;
  assign new_P1_U6169 = ~n1394 | ~new_P1_U3053;
  assign new_P1_U6170 = ~P1_DATAO_REG_28_ | ~new_P1_U3430;
  assign new_P1_U6171 = ~n1394 | ~new_P1_U3054;
  assign new_P1_U6172 = ~P1_DATAO_REG_29_ | ~new_P1_U3430;
  assign new_P1_U6173 = ~n1394 | ~new_P1_U3055;
  assign new_P1_U6174 = ~P1_DATAO_REG_30_ | ~new_P1_U3430;
  assign new_P1_U6175 = ~n1394 | ~new_P1_U3059;
  assign new_P1_U6176 = ~P1_DATAO_REG_31_ | ~new_P1_U3430;
  assign new_P1_U6177 = ~n1394 | ~new_P1_U3056;
  assign new_P1_U6178 = ~new_P1_U3432 | ~new_P1_U3450 | ~new_P1_U5793;
  assign new_P1_U6179 = ~new_P1_R1375_U9 | ~new_P1_U4030;
  assign new_P1_U6180 = ~new_P1_U4017 | ~new_P1_U3054;
  assign new_P1_U6181 = ~new_P1_U3413 | ~new_P1_U4702;
  assign new_P1_U6182 = ~new_P1_U6181 | ~new_P1_U6180;
  assign new_P1_U6183 = ~new_P1_U4026 | ~new_P1_U3056;
  assign new_P1_U6184 = ~new_P1_U3418 | ~new_P1_U4759;
  assign new_P1_U6185 = ~new_P1_U6184 | ~new_P1_U6183;
  assign new_P1_U6186 = ~new_P1_U4025 | ~new_P1_U3076;
  assign new_P1_U6187 = ~new_P1_U3397 | ~new_P1_U4550;
  assign new_P1_U6188 = ~new_P1_U6187 | ~new_P1_U6186;
  assign new_P1_U6189 = ~new_P1_U4027 | ~new_P1_U3059;
  assign new_P1_U6190 = ~new_P1_U3417 | ~new_P1_U4739;
  assign new_P1_U6191 = ~new_P1_U6190 | ~new_P1_U6189;
  assign new_P1_U6192 = ~new_P1_U5959 | ~new_P1_U4531;
  assign new_P1_U6193 = ~new_P1_U3514 | ~new_P1_U3081;
  assign new_P1_U6194 = ~new_P1_U6193 | ~new_P1_U6192;
  assign new_P1_U6195 = ~new_P1_U5905 | ~new_P1_U4379;
  assign new_P1_U6196 = ~new_P1_U3491 | ~new_P1_U3063;
  assign new_P1_U6197 = ~new_P1_U6196 | ~new_P1_U6195;
  assign new_P1_U6198 = ~new_P1_U5856 | ~new_P1_U4246;
  assign new_P1_U6199 = ~new_P1_U3470 | ~new_P1_U3060;
  assign new_P1_U6200 = ~new_P1_U6199 | ~new_P1_U6198;
  assign new_P1_U6201 = ~new_P1_U5898 | ~new_P1_U4360;
  assign new_P1_U6202 = ~new_P1_U3488 | ~new_P1_U3062;
  assign new_P1_U6203 = ~new_P1_U6202 | ~new_P1_U6201;
  assign new_P1_U6204 = ~new_P1_U4028 | ~new_P1_U3055;
  assign new_P1_U6205 = ~new_P1_U3415 | ~new_P1_U4721;
  assign new_P1_U6206 = ~new_P1_U6205 | ~new_P1_U6204;
  assign new_P1_U6207 = ~new_P1_U4018 | ~new_P1_U3053;
  assign new_P1_U6208 = ~new_P1_U3411 | ~new_P1_U4683;
  assign new_P1_U6209 = ~new_P1_U6208 | ~new_P1_U6207;
  assign new_P1_U6210 = ~new_P1_U5947 | ~new_P1_U4493;
  assign new_P1_U6211 = ~new_P1_U3509 | ~new_P1_U3069;
  assign new_P1_U6212 = ~new_P1_U6211 | ~new_P1_U6210;
  assign new_P1_U6213 = ~new_P1_U5884 | ~new_P1_U4322;
  assign new_P1_U6214 = ~new_P1_U3482 | ~new_P1_U3084;
  assign new_P1_U6215 = ~new_P1_U6214 | ~new_P1_U6213;
  assign new_P1_U6216 = ~new_P1_U5891 | ~new_P1_U4341;
  assign new_P1_U6217 = ~new_P1_U3485 | ~new_P1_U3083;
  assign new_P1_U6218 = ~new_P1_U6217 | ~new_P1_U6216;
  assign new_P1_U6219 = ~new_P1_U5919 | ~new_P1_U4417;
  assign new_P1_U6220 = ~new_P1_U3497 | ~new_P1_U3080;
  assign new_P1_U6221 = ~new_P1_U6220 | ~new_P1_U6219;
  assign new_P1_U6222 = ~new_P1_U5926 | ~new_P1_U4436;
  assign new_P1_U6223 = ~new_P1_U3500 | ~new_P1_U3079;
  assign new_P1_U6224 = ~new_P1_U6223 | ~new_P1_U6222;
  assign new_P1_U6225 = ~new_P1_U5820 | ~new_P1_U4208;
  assign new_P1_U6226 = ~new_P1_U3456 | ~new_P1_U3077;
  assign new_P1_U6227 = ~new_P1_U6226 | ~new_P1_U6225;
  assign new_P1_U6228 = ~new_P1_U5835 | ~new_P1_U4184;
  assign new_P1_U6229 = ~new_P1_U3461 | ~new_P1_U3078;
  assign new_P1_U6230 = ~new_P1_U6229 | ~new_P1_U6228;
  assign new_P1_U6231 = ~new_P1_U5933 | ~new_P1_U4455;
  assign new_P1_U6232 = ~new_P1_U3503 | ~new_P1_U3074;
  assign new_P1_U6233 = ~new_P1_U6232 | ~new_P1_U6231;
  assign new_P1_U6234 = ~new_P1_U5940 | ~new_P1_U4474;
  assign new_P1_U6235 = ~new_P1_U3506 | ~new_P1_U3073;
  assign new_P1_U6236 = ~new_P1_U6235 | ~new_P1_U6234;
  assign new_P1_U6237 = ~new_P1_U5870 | ~new_P1_U4284;
  assign new_P1_U6238 = ~new_P1_U3476 | ~new_P1_U3071;
  assign new_P1_U6239 = ~new_P1_U6238 | ~new_P1_U6237;
  assign new_P1_U6240 = ~new_P1_U5877 | ~new_P1_U4303;
  assign new_P1_U6241 = ~new_P1_U3479 | ~new_P1_U3070;
  assign new_P1_U6242 = ~new_P1_U6241 | ~new_P1_U6240;
  assign new_P1_U6243 = ~new_P1_U5912 | ~new_P1_U4398;
  assign new_P1_U6244 = ~new_P1_U3494 | ~new_P1_U3072;
  assign new_P1_U6245 = ~new_P1_U6244 | ~new_P1_U6243;
  assign new_P1_U6246 = ~new_P1_U5842 | ~new_P1_U4203;
  assign new_P1_U6247 = ~new_P1_U3464 | ~new_P1_U3068;
  assign new_P1_U6248 = ~new_P1_U6247 | ~new_P1_U6246;
  assign new_P1_U6249 = ~new_P1_U5849 | ~new_P1_U4227;
  assign new_P1_U6250 = ~new_P1_U3467 | ~new_P1_U3064;
  assign new_P1_U6251 = ~new_P1_U6250 | ~new_P1_U6249;
  assign new_P1_U6252 = ~new_P1_U5863 | ~new_P1_U4265;
  assign new_P1_U6253 = ~new_P1_U3473 | ~new_P1_U3067;
  assign new_P1_U6254 = ~new_P1_U6253 | ~new_P1_U6252;
  assign new_P1_U6255 = ~new_P1_U5954 | ~new_P1_U4512;
  assign new_P1_U6256 = ~new_P1_U3512 | ~new_P1_U3082;
  assign new_P1_U6257 = ~new_P1_U6256 | ~new_P1_U6255;
  assign new_P1_U6258 = ~new_P1_U4021 | ~new_P1_U3065;
  assign new_P1_U6259 = ~new_P1_U3405 | ~new_P1_U4626;
  assign new_P1_U6260 = ~new_P1_U6259 | ~new_P1_U6258;
  assign new_P1_U6261 = ~new_P1_U4022 | ~new_P1_U3066;
  assign new_P1_U6262 = ~new_P1_U3403 | ~new_P1_U4607;
  assign new_P1_U6263 = ~new_P1_U6262 | ~new_P1_U6261;
  assign new_P1_U6264 = ~new_P1_U4024 | ~new_P1_U3075;
  assign new_P1_U6265 = ~new_P1_U3399 | ~new_P1_U4569;
  assign new_P1_U6266 = ~new_P1_U6265 | ~new_P1_U6264;
  assign new_P1_U6267 = ~new_P1_U4023 | ~new_P1_U3061;
  assign new_P1_U6268 = ~new_P1_U3401 | ~new_P1_U4588;
  assign new_P1_U6269 = ~new_P1_U6268 | ~new_P1_U6267;
  assign new_P1_U6270 = ~new_P1_U4020 | ~new_P1_U3058;
  assign new_P1_U6271 = ~new_P1_U3407 | ~new_P1_U4645;
  assign new_P1_U6272 = ~new_P1_U6271 | ~new_P1_U6270;
  assign new_P1_U6273 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_U6274 = ~new_P1_U3409 | ~new_P1_U4664;
  assign new_P1_U6275 = ~new_P1_U6274 | ~new_P1_U6273;
  assign new_P1_U6276 = ~new_P1_U4041 | ~new_P1_U3991;
  assign new_P1_U6277 = ~new_P1_U5129 | ~new_P1_U3049;
  assign new_P1_U6278 = ~new_P1_U5799 | ~new_P1_U5133 | ~new_P1_U3432;
  assign new_P1_U6279 = ~new_P1_U3453 | ~new_P1_U5130;
  assign new_P1_U6280 = ~new_P1_U5786 | ~new_P1_U3431;
  assign new_P1_U6281 = ~new_P1_U3451 | ~new_P1_U3444;
  assign new_P1_U6282 = ~new_P1_U3450 | ~new_P1_U5144;
  assign new_P1_U6283 = ~new_P1_U5802 | ~new_P1_U3994;
  assign new_P1_U6284 = ~new_P1_U3454 | ~new_P1_U5408;
  assign new_P1_U6285 = ~new_P1_U5814 | ~new_P1_U3015 | ~P1_REG2_REG_0_;
  assign new_P3_R1161_U489 = ~new_P3_U3079 | ~new_P3_R1161_U69;
  assign new_P3_R1161_U488 = ~new_P3_R1161_U254 | ~new_P3_R1161_U486;
  assign new_P3_R1161_U487 = ~new_P3_R1161_U165 | ~new_P3_R1161_U166;
  assign new_P3_R1161_U486 = ~new_P3_R1161_U485 | ~new_P3_R1161_U484;
  assign new_P3_R1161_U485 = ~new_P3_U3431 | ~new_P3_R1161_U72;
  assign new_P3_R1161_U484 = ~new_P3_U3078 | ~new_P3_R1161_U71;
  assign new_P3_R1161_U483 = ~new_P3_U3431 | ~new_P3_R1161_U72;
  assign new_P3_R1161_U482 = ~new_P3_U3078 | ~new_P3_R1161_U71;
  assign new_P3_R1161_U481 = ~new_P3_R1161_U258 | ~new_P3_R1161_U479;
  assign new_P3_R1161_U480 = ~new_P3_R1161_U163 | ~new_P3_R1161_U164;
  assign new_P3_R1161_U479 = ~new_P3_R1161_U478 | ~new_P3_R1161_U477;
  assign new_P3_R1161_U478 = ~new_P3_U3434 | ~new_P3_R1161_U74;
  assign new_P3_R1161_U477 = ~new_P3_U3073 | ~new_P3_R1161_U73;
  assign new_P3_R1161_U476 = ~new_P3_U3434 | ~new_P3_R1161_U74;
  assign new_P3_R1161_U475 = ~new_P3_U3073 | ~new_P3_R1161_U73;
  assign new_P3_R1161_U474 = ~new_P3_R1161_U472 | ~new_P3_R1161_U262;
  assign new_P3_R1161_U473 = ~new_P3_R1161_U361 | ~new_P3_R1161_U92;
  assign new_P3_R1161_U472 = ~new_P3_R1161_U471 | ~new_P3_R1161_U470;
  assign new_P3_R1161_U471 = ~new_P3_U3437 | ~new_P3_R1161_U57;
  assign new_P3_R1161_U470 = ~new_P3_U3072 | ~new_P3_R1161_U56;
  assign new_P3_R1161_U469 = ~new_P3_U3440 | ~new_P3_R1161_U58;
  assign new_P2_U3014 = new_P2_U3924 & new_P2_U5671;
  assign new_P2_U3015 = new_P2_U3937 & new_P2_U3419;
  assign new_P2_U3016 = new_P2_U3575 & new_P2_U3570;
  assign new_P2_U3017 = new_P2_U5688 & new_P2_U3423;
  assign new_P2_U3018 = new_P2_U3426 & new_P2_U3423;
  assign new_P2_U3019 = new_P2_U3421 & new_P2_U3422;
  assign new_P2_U3020 = new_P2_U5680 & new_P2_U3421;
  assign new_P2_U3021 = new_P2_U5677 & new_P2_U3422;
  assign new_P2_U3022 = new_P2_U5677 & new_P2_U5680;
  assign new_P2_U3023 = new_P2_U3048 & P2_STATE_REG;
  assign new_P2_U3024 = new_P2_U3757 & new_P2_U3401;
  assign new_P2_U3025 = new_P2_U3976 & new_P2_U5671;
  assign new_P2_U3026 = new_P2_U3963 & new_P2_U5683;
  assign new_P2_U3027 = new_P2_U3944 & new_P2_U5671;
  assign new_P2_U3028 = new_P2_U3803 & new_P2_U3946;
  assign new_P2_U3029 = new_P2_R1299_U6 & new_P2_U3411;
  assign new_P2_U3030 = new_P2_U3329 & P2_STATE_REG;
  assign new_P2_U3031 = new_P2_U3932 & new_P2_U3964;
  assign new_P2_U3032 = new_P2_U3964 & new_P2_U3398;
  assign new_P2_U3033 = new_P2_U3933 & new_P2_U3964;
  assign new_P2_U3034 = new_P2_U3938 & new_P2_U3964;
  assign new_P2_U3035 = new_P2_U3963 & new_P2_U3423;
  assign new_P2_U3036 = new_P2_U3946 & new_P2_U5683;
  assign new_P2_U3037 = new_P2_U3964 & new_P2_U3026;
  assign new_P2_U3038 = new_P2_U3946 & new_P2_U3423;
  assign new_P2_U3039 = new_P2_U5688 & new_P2_U4854;
  assign new_P2_U3040 = new_P2_U3024 & new_P2_U5688;
  assign new_P2_U3041 = new_P2_U5683 & new_P2_U4854;
  assign new_P2_U3042 = new_P2_U3024 & new_P2_U5683;
  assign new_P2_U3043 = new_P2_U3018 & new_P2_U4854;
  assign new_P2_U3044 = new_P2_U3024 & new_P2_U3018;
  assign new_P2_U3045 = new_P2_U3023 & new_P2_U3401;
  assign new_P2_U3046 = new_P2_U5184 & P2_STATE_REG;
  assign new_P2_U3047 = new_P2_U3023 & new_P2_U5186;
  assign new_P2_U3048 = new_P2_U5658 & new_P2_U3396;
  assign new_P2_U3049 = new_P2_U3418 & new_P2_U5668;
  assign new_P2_U3050 = new_P2_U3576 & new_P2_U3016;
  assign new_P2_U3051 = new_P2_U3337 & new_P2_U3338 & new_P2_U3392 & new_P2_U3341 & new_P2_U3402;
  assign new_P2_U3052 = new_P2_U3399 & P2_STATE_REG;
  assign new_P2_U3053 = new_P2_U3819 & new_P2_U3820 & new_P2_U5439;
  assign new_P2_U3054 = new_P2_U5461 & new_P2_U5460;
  assign new_P2_U3055 = ~new_P2_U4613 | ~new_P2_U4610 | ~new_P2_U4611 | ~new_P2_U4612;
  assign new_P2_U3056 = ~new_P2_U4632 | ~new_P2_U4629 | ~new_P2_U4630 | ~new_P2_U4631;
  assign new_P2_U3057 = ~new_P2_U4648 | ~new_P2_U4649 | ~new_P2_U4651 | ~new_P2_U4650;
  assign new_P2_U3058 = ~new_P2_U4687 | ~new_P2_U4688 | ~new_P2_U4689;
  assign new_P2_U3059 = ~new_P2_U4594 | ~new_P2_U4591 | ~new_P2_U4592 | ~new_P2_U4593;
  assign new_P2_U3060 = ~new_P2_U4575 | ~new_P2_U4572 | ~new_P2_U4573 | ~new_P2_U4574;
  assign new_P2_U3061 = ~new_P2_U4667 | ~new_P2_U4668 | ~new_P2_U4669;
  assign new_P2_U3062 = ~new_P2_U4173 | ~new_P2_U4174 | ~new_P2_U4176 | ~new_P2_U4175;
  assign new_P2_U3063 = ~new_P2_U4518 | ~new_P2_U4515 | ~new_P2_U4516 | ~new_P2_U4517;
  assign new_P2_U3064 = ~new_P2_U4287 | ~new_P2_U4288 | ~new_P2_U4290 | ~new_P2_U4289;
  assign new_P2_U3065 = ~new_P2_U4306 | ~new_P2_U4307 | ~new_P2_U4309 | ~new_P2_U4308;
  assign new_P2_U3066 = ~new_P2_U4154 | ~new_P2_U4155 | ~new_P2_U4157 | ~new_P2_U4156;
  assign new_P2_U3067 = ~new_P2_U4556 | ~new_P2_U4553 | ~new_P2_U4554 | ~new_P2_U4555;
  assign new_P2_U3068 = ~new_P2_U4537 | ~new_P2_U4534 | ~new_P2_U4535 | ~new_P2_U4536;
  assign new_P2_U3069 = ~new_P2_U4192 | ~new_P2_U4193 | ~new_P2_U4195 | ~new_P2_U4194;
  assign new_P2_U3070 = ~new_P2_U4130 | ~new_P2_U4131 | ~new_P2_U4133 | ~new_P2_U4132;
  assign new_P2_U3071 = ~new_P2_U4423 | ~new_P2_U4420 | ~new_P2_U4421 | ~new_P2_U4422;
  assign new_P2_U3072 = ~new_P2_U4230 | ~new_P2_U4231 | ~new_P2_U4233 | ~new_P2_U4232;
  assign new_P2_U3073 = ~new_P2_U4211 | ~new_P2_U4212 | ~new_P2_U4214 | ~new_P2_U4213;
  assign new_P2_U3074 = ~new_P2_U4325 | ~new_P2_U4326 | ~new_P2_U4328 | ~new_P2_U4327;
  assign new_P2_U3075 = ~new_P2_U4401 | ~new_P2_U4402 | ~new_P2_U4404 | ~new_P2_U4403;
  assign new_P2_U3076 = ~new_P2_U4382 | ~new_P2_U4383 | ~new_P2_U4385 | ~new_P2_U4384;
  assign new_P2_U3077 = ~new_P2_U4499 | ~new_P2_U4496 | ~new_P2_U4497 | ~new_P2_U4498;
  assign new_P2_U3078 = ~new_P2_U4480 | ~new_P2_U4477 | ~new_P2_U4478 | ~new_P2_U4479;
  assign new_P2_U3079 = ~new_P2_U4135 | ~new_P2_U4136 | ~new_P2_U4138 | ~new_P2_U4137;
  assign new_P2_U3080 = ~new_P2_U4111 | ~new_P2_U4112 | ~new_P2_U4114 | ~new_P2_U4113;
  assign new_P2_U3081 = ~new_P2_U4363 | ~new_P2_U4364 | ~new_P2_U4366 | ~new_P2_U4365;
  assign new_P2_U3082 = ~new_P2_U4344 | ~new_P2_U4345 | ~new_P2_U4347 | ~new_P2_U4346;
  assign new_P2_U3083 = ~new_P2_U4461 | ~new_P2_U4458 | ~new_P2_U4459 | ~new_P2_U4460;
  assign new_P2_U3084 = ~new_P2_U4442 | ~new_P2_U4439 | ~new_P2_U4440 | ~new_P2_U4441;
  assign new_P2_U3085 = ~new_P2_U4268 | ~new_P2_U4269 | ~new_P2_U4271 | ~new_P2_U4270;
  assign new_P2_U3086 = ~new_P2_U4249 | ~new_P2_U4250 | ~new_P2_U4252 | ~new_P2_U4251;
  assign n2614 = ~new_P2_U3815 | ~new_P2_U5434;
  assign n2609 = ~P2_STATE_REG;
  assign new_P2_U3089 = ~new_P2_U5557 | ~new_P2_U5556;
  assign new_P2_U3090 = ~new_P2_U5559 | ~new_P2_U5558;
  assign new_P2_U3091 = ~new_P2_U3859 | ~new_P2_U5563;
  assign new_P2_U3092 = ~new_P2_U3860 | ~new_P2_U5566;
  assign new_P2_U3093 = ~new_P2_U3861 | ~new_P2_U5569;
  assign new_P2_U3094 = ~new_P2_U3862 | ~new_P2_U5572;
  assign new_P2_U3095 = ~new_P2_U3863 | ~new_P2_U5575;
  assign new_P2_U3096 = ~new_P2_U3864 | ~new_P2_U5578;
  assign new_P2_U3097 = ~new_P2_U3865 | ~new_P2_U5581;
  assign new_P2_U3098 = ~new_P2_U3866 | ~new_P2_U5584;
  assign new_P2_U3099 = ~new_P2_U3867 | ~new_P2_U5587;
  assign new_P2_U3100 = ~new_P2_U3868 | ~new_P2_U5590;
  assign new_P2_U3101 = ~new_P2_U3869 | ~new_P2_U5596;
  assign new_P2_U3102 = ~new_P2_U3870 | ~new_P2_U5599;
  assign new_P2_U3103 = ~new_P2_U3871 | ~new_P2_U5602;
  assign new_P2_U3104 = ~new_P2_U3872 | ~new_P2_U5605;
  assign new_P2_U3105 = ~new_P2_U3873 | ~new_P2_U5608;
  assign new_P2_U3106 = ~new_P2_U3874 | ~new_P2_U5611;
  assign new_P2_U3107 = ~new_P2_U3875 | ~new_P2_U5614;
  assign new_P2_U3108 = ~new_P2_U3876 | ~new_P2_U5617;
  assign new_P2_U3109 = ~new_P2_U3877 | ~new_P2_U5620;
  assign new_P2_U3110 = ~new_P2_U3878 | ~new_P2_U5623;
  assign new_P2_U3111 = ~new_P2_U3857 | ~new_P2_U5538;
  assign new_P2_U3112 = ~new_P2_U3858 | ~new_P2_U5541;
  assign new_P2_U3113 = ~new_P2_U5546 | ~new_P2_U5545 | ~new_P2_U5544;
  assign new_P2_U3114 = ~new_P2_U5549 | ~new_P2_U5548 | ~new_P2_U5547;
  assign new_P2_U3115 = ~new_P2_U5552 | ~new_P2_U5551 | ~new_P2_U5550;
  assign new_P2_U3116 = ~new_P2_U5555 | ~new_P2_U5554 | ~new_P2_U5553;
  assign new_P2_U3117 = ~new_P2_U5562 | ~new_P2_U5561 | ~new_P2_U5560;
  assign new_P2_U3118 = ~new_P2_U5595 | ~new_P2_U5594 | ~new_P2_U5593;
  assign new_P2_U3119 = ~new_P2_U5628 | ~new_P2_U5627 | ~new_P2_U5626;
  assign new_P2_U3120 = ~new_P2_U5630 | ~new_P2_U5629;
  assign new_P2_U3121 = new_P2_U5638 & new_P2_U5637 & new_P2_U5632;
  assign new_P2_U3122 = ~new_P2_U5464 | ~new_P2_U5463 | ~new_P2_U5462;
  assign new_P2_U3123 = ~new_P2_U5470 | ~new_P2_U5469 | ~new_P2_U3831;
  assign new_P2_U3124 = ~new_P2_U5473 | ~new_P2_U5472 | ~new_P2_U3832;
  assign new_P2_U3125 = ~new_P2_U5476 | ~new_P2_U5475 | ~new_P2_U3833;
  assign new_P2_U3126 = ~new_P2_U5479 | ~new_P2_U5478 | ~new_P2_U3834;
  assign new_P2_U3127 = ~new_P2_U5482 | ~new_P2_U5481 | ~new_P2_U3835;
  assign new_P2_U3128 = ~new_P2_U5485 | ~new_P2_U5484 | ~new_P2_U3836;
  assign new_P2_U3129 = ~new_P2_U5488 | ~new_P2_U5487 | ~new_P2_U3837;
  assign new_P2_U3130 = ~new_P2_U5491 | ~new_P2_U5490 | ~new_P2_U3838;
  assign new_P2_U3131 = ~new_P2_U5494 | ~new_P2_U5493 | ~new_P2_U3839;
  assign new_P2_U3132 = ~new_P2_U5497 | ~new_P2_U5496 | ~new_P2_U3840;
  assign new_P2_U3133 = ~new_P2_U5503 | ~new_P2_U5502 | ~new_P2_U3843;
  assign new_P2_U3134 = ~new_P2_U5506 | ~new_P2_U5505 | ~new_P2_U3844;
  assign new_P2_U3135 = ~new_P2_U5509 | ~new_P2_U5508 | ~new_P2_U3845;
  assign new_P2_U3136 = ~new_P2_U5512 | ~new_P2_U5511 | ~new_P2_U3846;
  assign new_P2_U3137 = ~new_P2_U5515 | ~new_P2_U5514 | ~new_P2_U3847;
  assign new_P2_U3138 = ~new_P2_U5518 | ~new_P2_U5517 | ~new_P2_U3848;
  assign new_P2_U3139 = ~new_P2_U5521 | ~new_P2_U5520 | ~new_P2_U3849;
  assign new_P2_U3140 = ~new_P2_U5524 | ~new_P2_U5523 | ~new_P2_U3850;
  assign new_P2_U3141 = ~new_P2_U3851 | ~new_P2_U5526 | ~new_P2_U5525;
  assign new_P2_U3142 = ~new_P2_U3852 | ~new_P2_U5529 | ~new_P2_U5528;
  assign new_P2_U3143 = ~new_P2_U3821 | ~new_P2_U5443 | ~new_P2_U5442;
  assign new_P2_U3144 = ~new_P2_U3822 | ~new_P2_U5446 | ~new_P2_U5445;
  assign new_P2_U3145 = ~new_P2_U3823 | ~new_P2_U5449 | ~new_P2_U5448;
  assign new_P2_U3146 = ~new_P2_U3824 | ~new_P2_U5452 | ~new_P2_U5451;
  assign new_P2_U3147 = ~new_P2_U3825 | ~new_P2_U5455 | ~new_P2_U5454;
  assign new_P2_U3148 = ~new_P2_U5458 | ~new_P2_U3826;
  assign new_P2_U3149 = ~new_P2_U5466 | ~new_P2_U3829;
  assign new_P2_U3150 = ~new_P2_U5499 | ~new_P2_U3841;
  assign new_P2_U3151 = ~new_P2_U5532 | ~new_P2_U3853;
  assign new_P2_U3152 = ~new_P2_U5535 | ~new_P2_U3855;
  assign new_P2_U3153 = ~new_P2_U3415 | ~new_P2_U3817 | ~new_P2_U3345;
  assign new_P2_U3154 = ~new_P2_U3015 | ~new_P2_U5658;
  assign new_P2_U3155 = new_P2_U5437 & new_P2_U3056;
  assign new_P2_U3156 = new_P2_U5437 & new_P2_U3055;
  assign new_P2_U3157 = new_P2_U5437 & new_P2_U3059;
  assign new_P2_U3158 = new_P2_U5437 & new_P2_U3060;
  assign new_P2_U3159 = new_P2_U5437 & new_P2_U3067;
  assign new_P2_U3160 = new_P2_U5437 & new_P2_U3068;
  assign new_P2_U3161 = new_P2_U5437 & new_P2_U3063;
  assign new_P2_U3162 = new_P2_U5437 & new_P2_U3077;
  assign new_P2_U3163 = new_P2_U5437 & new_P2_U3078;
  assign new_P2_U3164 = new_P2_U5437 & new_P2_U3083;
  assign new_P2_U3165 = new_P2_U5437 & new_P2_U3084;
  assign new_P2_U3166 = new_P2_U5437 & new_P2_U3071;
  assign new_P2_U3167 = new_P2_U5437 & new_P2_U3075;
  assign new_P2_U3168 = new_P2_U5437 & new_P2_U3076;
  assign new_P2_U3169 = new_P2_U5437 & new_P2_U3081;
  assign new_P2_U3170 = new_P2_U5437 & new_P2_U3082;
  assign new_P2_U3171 = new_P2_U5437 & new_P2_U3074;
  assign new_P2_U3172 = new_P2_U5437 & new_P2_U3065;
  assign new_P2_U3173 = new_P2_U5437 & new_P2_U3064;
  assign new_P2_U3174 = new_P2_U5437 & new_P2_U3085;
  assign new_P2_U3175 = new_P2_U5437 & new_P2_U3086;
  assign new_P2_U3176 = new_P2_U5437 & new_P2_U3072;
  assign new_P2_U3177 = new_P2_U5437 & new_P2_U3073;
  assign new_P2_U3178 = new_P2_U5437 & new_P2_U3069;
  assign new_P2_U3179 = new_P2_U5437 & new_P2_U3062;
  assign new_P2_U3180 = new_P2_U5437 & new_P2_U3066;
  assign new_P2_U3181 = new_P2_U5437 & new_P2_U3070;
  assign new_P2_U3182 = new_P2_U5437 & new_P2_U3080;
  assign new_P2_U3183 = new_P2_U5437 & new_P2_U3079;
  assign new_P2_U3184 = ~new_P2_U3343 | ~new_P2_U3404 | ~new_P2_U5436;
  assign n2604 = ~new_P2_U5430 | ~new_P2_U3814 | ~new_P2_U5433 | ~new_P2_U5432;
  assign n2599 = ~new_P2_U5422 | ~new_P2_U5420 | ~new_P2_U5421 | ~new_P2_U5424 | ~new_P2_U5423;
  assign n2594 = ~new_P2_U5413 | ~new_P2_U5414 | ~new_P2_U5415 | ~new_P2_U5412 | ~new_P2_U5411;
  assign n2589 = ~new_P2_U5404 | ~new_P2_U5402 | ~new_P2_U5403 | ~new_P2_U5406 | ~new_P2_U5405;
  assign n2584 = ~new_P2_U5396 | ~new_P2_U5397 | ~new_P2_U5395 | ~new_P2_U5394 | ~new_P2_U5393;
  assign n2579 = ~new_P2_U5385 | ~new_P2_U3813 | ~new_P2_U5388 | ~new_P2_U5387;
  assign n2574 = ~new_P2_U5377 | ~new_P2_U5378 | ~new_P2_U5379 | ~new_P2_U5376 | ~new_P2_U5375;
  assign n2569 = ~new_P2_U5368 | ~new_P2_U5366 | ~new_P2_U5367 | ~new_P2_U5370 | ~new_P2_U5369;
  assign n2564 = ~new_P2_U5358 | ~new_P2_U3812 | ~new_P2_U5361 | ~new_P2_U5360;
  assign n2559 = ~new_P2_U5349 | ~new_P2_U3811 | ~new_P2_U5352 | ~new_P2_U5351;
  assign n2554 = ~new_P2_U5341 | ~new_P2_U5342 | ~new_P2_U5343 | ~new_P2_U5340 | ~new_P2_U5339;
  assign n2549 = ~new_P2_U5332 | ~new_P2_U5333 | ~new_P2_U5334 | ~new_P2_U5331 | ~new_P2_U5330;
  assign n2544 = ~new_P2_U5323 | ~new_P2_U5321 | ~new_P2_U5322 | ~new_P2_U5325 | ~new_P2_U5324;
  assign n2539 = ~new_P2_U5314 | ~new_P2_U5315 | ~new_P2_U5316 | ~new_P2_U5313 | ~new_P2_U5312;
  assign n2534 = ~new_P2_U5304 | ~new_P2_U3810 | ~new_P2_U5307 | ~new_P2_U5306;
  assign n2529 = ~new_P2_U5296 | ~new_P2_U5297 | ~new_P2_U5298 | ~new_P2_U5295 | ~new_P2_U5294;
  assign n2524 = ~new_P2_U5287 | ~new_P2_U5285 | ~new_P2_U5286 | ~new_P2_U5289 | ~new_P2_U5288;
  assign n2519 = ~new_P2_U5277 | ~new_P2_U3809 | ~new_P2_U5280 | ~new_P2_U5279;
  assign n2514 = ~new_P2_U5270 | ~new_P2_U5271 | ~new_P2_U5269 | ~new_P2_U5268 | ~new_P2_U5267;
  assign n2509 = ~new_P2_U3807 | ~new_P2_U3808 | ~new_P2_U5260;
  assign n2504 = ~new_P2_U5252 | ~new_P2_U5253 | ~new_P2_U5254 | ~new_P2_U5251 | ~new_P2_U5250;
  assign n2499 = ~new_P2_U5243 | ~new_P2_U5244 | ~new_P2_U5245 | ~new_P2_U5242 | ~new_P2_U5241;
  assign n2494 = ~new_P2_U5234 | ~new_P2_U5232 | ~new_P2_U5233 | ~new_P2_U5236 | ~new_P2_U5235;
  assign n2489 = ~new_P2_U5226 | ~new_P2_U5227 | ~new_P2_U5225 | ~new_P2_U5224 | ~new_P2_U5223;
  assign n2484 = ~new_P2_U5215 | ~new_P2_U3805 | ~new_P2_U5218 | ~new_P2_U5217;
  assign n2479 = ~new_P2_U5207 | ~new_P2_U5208 | ~new_P2_U5209 | ~new_P2_U5206 | ~new_P2_U5205;
  assign n2474 = ~new_P2_U5197 | ~new_P2_U3804 | ~new_P2_U5200 | ~new_P2_U5199;
  assign n2469 = ~new_P2_U5189 | ~new_P2_U5187 | ~new_P2_U5188 | ~new_P2_U5191 | ~new_P2_U5190;
  assign n2464 = ~new_P2_U5176 | ~new_P2_U5177 | ~new_P2_U5178 | ~new_P2_U5175 | ~new_P2_U5174;
  assign n2294 = ~new_P2_U3786 | ~new_P2_U3785 | ~new_P2_U5150 | ~new_P2_U5149;
  assign n2289 = ~new_P2_U3784 | ~new_P2_U3783 | ~new_P2_U5135 | ~new_P2_U5134;
  assign n2284 = ~new_P2_U3782 | ~new_P2_U3781 | ~new_P2_U5120 | ~new_P2_U5119;
  assign n2279 = ~new_P2_U3780 | ~new_P2_U3779 | ~new_P2_U5105 | ~new_P2_U5104;
  assign n2274 = ~new_P2_U3778 | ~new_P2_U3777 | ~new_P2_U5090 | ~new_P2_U5089;
  assign n2269 = ~new_P2_U3776 | ~new_P2_U3775 | ~new_P2_U5075 | ~new_P2_U5074;
  assign n2264 = ~new_P2_U3774 | ~new_P2_U3773 | ~new_P2_U5060 | ~new_P2_U5059;
  assign n2259 = ~new_P2_U3772 | ~new_P2_U3771 | ~new_P2_U5045 | ~new_P2_U5044;
  assign n2254 = ~new_P2_U3770 | ~new_P2_U3769 | ~new_P2_U5030 | ~new_P2_U5029;
  assign n2249 = ~new_P2_U3768 | ~new_P2_U5015 | ~new_P2_U5014;
  assign n2244 = ~new_P2_U3767 | ~new_P2_U5000 | ~new_P2_U4999;
  assign n2239 = ~new_P2_U3766 | ~new_P2_U4985 | ~new_P2_U4984;
  assign n2234 = ~new_P2_U3765 | ~new_P2_U4970 | ~new_P2_U4969;
  assign n2229 = ~new_P2_U3764 | ~new_P2_U4955 | ~new_P2_U4954;
  assign n2224 = ~new_P2_U3763 | ~new_P2_U4940 | ~new_P2_U4939;
  assign n2219 = ~new_P2_U3762 | ~new_P2_U4925 | ~new_P2_U4924;
  assign n2214 = ~new_P2_U3761 | ~new_P2_U4910 | ~new_P2_U4909;
  assign n2209 = ~new_P2_U3760 | ~new_P2_U4895 | ~new_P2_U4894;
  assign n2204 = ~new_P2_U3759 | ~new_P2_U4880 | ~new_P2_U4879;
  assign n2199 = ~new_P2_U3758 | ~new_P2_U4865 | ~new_P2_U4864;
  assign n2194 = ~new_P2_U4853 | ~new_P2_U3915 | ~new_P2_U4852;
  assign n2189 = ~new_P2_U4851 | ~new_P2_U3914 | ~new_P2_U4850;
  assign n2184 = ~new_P2_U3912 | ~new_P2_U4846 | ~new_P2_U4849 | ~new_P2_U4847 | ~new_P2_U4848;
  assign n2179 = ~new_P2_U3911 | ~new_P2_U4842 | ~new_P2_U3753 | ~new_P2_U3754;
  assign n2174 = ~new_P2_U3910 | ~new_P2_U4837 | ~new_P2_U3751 | ~new_P2_U3752;
  assign n2169 = ~new_P2_U3909 | ~new_P2_U4832 | ~new_P2_U3749 | ~new_P2_U3750;
  assign n2164 = ~new_P2_U3908 | ~new_P2_U4827 | ~new_P2_U3747 | ~new_P2_U3748;
  assign n2159 = ~new_P2_U3907 | ~new_P2_U4822 | ~new_P2_U3745 | ~new_P2_U3746;
  assign n2154 = ~new_P2_U3906 | ~new_P2_U4817 | ~new_P2_U3743 | ~new_P2_U3744;
  assign n2149 = ~new_P2_U3905 | ~new_P2_U4812 | ~new_P2_U3741 | ~new_P2_U3742;
  assign n2144 = ~new_P2_U3904 | ~new_P2_U4807 | ~new_P2_U3739 | ~new_P2_U3740;
  assign n2139 = ~new_P2_U3903 | ~new_P2_U4802 | ~new_P2_U3737 | ~new_P2_U3738;
  assign n2134 = ~new_P2_U3902 | ~new_P2_U4797 | ~new_P2_U3735 | ~new_P2_U3736;
  assign n2129 = ~new_P2_U3901 | ~new_P2_U4792 | ~new_P2_U3733 | ~new_P2_U3734;
  assign n2124 = ~new_P2_U3900 | ~new_P2_U4787 | ~new_P2_U3731 | ~new_P2_U3732;
  assign n2119 = ~new_P2_U3899 | ~new_P2_U4782 | ~new_P2_U3729 | ~new_P2_U3730;
  assign n2114 = ~new_P2_U3898 | ~new_P2_U3728 | ~new_P2_U3727;
  assign n2109 = ~new_P2_U3897 | ~new_P2_U3726 | ~new_P2_U3725;
  assign n2104 = ~new_P2_U3896 | ~new_P2_U3724 | ~new_P2_U3723;
  assign n2099 = ~new_P2_U3895 | ~new_P2_U3722 | ~new_P2_U3721;
  assign n2094 = ~new_P2_U3894 | ~new_P2_U3720 | ~new_P2_U3719;
  assign n2089 = ~new_P2_U3893 | ~new_P2_U3718 | ~new_P2_U3717;
  assign n2084 = ~new_P2_U3716 | ~new_P2_U3715;
  assign n2079 = ~new_P2_U3714 | ~new_P2_U3713;
  assign n2074 = ~new_P2_U3712 | ~new_P2_U3711;
  assign n2069 = ~new_P2_U3710 | ~new_P2_U3709;
  assign n2064 = ~new_P2_U3708 | ~new_P2_U3707;
  assign n2059 = ~new_P2_U3706 | ~new_P2_U3705;
  assign n2054 = ~new_P2_U3704 | ~new_P2_U3703;
  assign n2049 = ~new_P2_U3702 | ~new_P2_U3701;
  assign n2044 = ~new_P2_U3700 | ~new_P2_U3699;
  assign n2039 = ~new_P2_U3698 | ~new_P2_U3697;
  assign n1714 = P2_D_REG_31_ & new_P2_U3880;
  assign n1709 = P2_D_REG_30_ & new_P2_U3880;
  assign n1704 = P2_D_REG_29_ & new_P2_U3880;
  assign n1699 = P2_D_REG_28_ & new_P2_U3880;
  assign n1694 = P2_D_REG_27_ & new_P2_U3880;
  assign n1689 = P2_D_REG_26_ & new_P2_U3880;
  assign n1684 = P2_D_REG_25_ & new_P2_U3880;
  assign n1679 = P2_D_REG_24_ & new_P2_U3880;
  assign n1674 = P2_D_REG_23_ & new_P2_U3880;
  assign n1669 = P2_D_REG_22_ & new_P2_U3880;
  assign n1664 = P2_D_REG_21_ & new_P2_U3880;
  assign n1659 = P2_D_REG_20_ & new_P2_U3880;
  assign n1654 = P2_D_REG_19_ & new_P2_U3880;
  assign n1649 = P2_D_REG_18_ & new_P2_U3880;
  assign n1644 = P2_D_REG_17_ & new_P2_U3880;
  assign n1639 = P2_D_REG_16_ & new_P2_U3880;
  assign n1634 = P2_D_REG_15_ & new_P2_U3880;
  assign n1629 = P2_D_REG_14_ & new_P2_U3880;
  assign n1624 = P2_D_REG_13_ & new_P2_U3880;
  assign n1619 = P2_D_REG_12_ & new_P2_U3880;
  assign n1614 = P2_D_REG_11_ & new_P2_U3880;
  assign n1609 = P2_D_REG_10_ & new_P2_U3880;
  assign n1604 = P2_D_REG_9_ & new_P2_U3880;
  assign n1599 = P2_D_REG_8_ & new_P2_U3880;
  assign n1594 = P2_D_REG_7_ & new_P2_U3880;
  assign n1589 = P2_D_REG_6_ & new_P2_U3880;
  assign n1584 = P2_D_REG_5_ & new_P2_U3880;
  assign n1579 = P2_D_REG_4_ & new_P2_U3880;
  assign n1574 = P2_D_REG_3_ & new_P2_U3880;
  assign n1569 = P2_D_REG_2_ & new_P2_U3880;
  assign n1554 = ~new_P2_U4072 | ~new_P2_U4073 | ~new_P2_U4074;
  assign n1549 = ~new_P2_U4069 | ~new_P2_U4070 | ~new_P2_U4071;
  assign n1544 = ~new_P2_U4066 | ~new_P2_U4067 | ~new_P2_U4068;
  assign n1539 = ~new_P2_U4063 | ~new_P2_U4064 | ~new_P2_U4065;
  assign n1534 = ~new_P2_U4060 | ~new_P2_U4061 | ~new_P2_U4062;
  assign n1529 = ~new_P2_U4057 | ~new_P2_U4058 | ~new_P2_U4059;
  assign n1524 = ~new_P2_U4054 | ~new_P2_U4055 | ~new_P2_U4056;
  assign n1519 = ~new_P2_U4051 | ~new_P2_U4052 | ~new_P2_U4053;
  assign n1514 = ~new_P2_U4048 | ~new_P2_U4049 | ~new_P2_U4050;
  assign n1509 = ~new_P2_U4045 | ~new_P2_U4046 | ~new_P2_U4047;
  assign n1504 = ~new_P2_U4042 | ~new_P2_U4043 | ~new_P2_U4044;
  assign n1499 = ~new_P2_U4039 | ~new_P2_U4040 | ~new_P2_U4041;
  assign n1494 = ~new_P2_U4036 | ~new_P2_U4037 | ~new_P2_U4038;
  assign n1489 = ~new_P2_U4033 | ~new_P2_U4034 | ~new_P2_U4035;
  assign n1484 = ~new_P2_U4030 | ~new_P2_U4031 | ~new_P2_U4032;
  assign n1479 = ~new_P2_U4027 | ~new_P2_U4028 | ~new_P2_U4029;
  assign n1474 = ~new_P2_U4024 | ~new_P2_U4025 | ~new_P2_U4026;
  assign n1469 = ~new_P2_U4021 | ~new_P2_U4022 | ~new_P2_U4023;
  assign n1464 = ~new_P2_U4018 | ~new_P2_U4019 | ~new_P2_U4020;
  assign n1459 = ~new_P2_U4015 | ~new_P2_U4016 | ~new_P2_U4017;
  assign n1454 = ~new_P2_U4012 | ~new_P2_U4013 | ~new_P2_U4014;
  assign n1449 = ~new_P2_U4009 | ~new_P2_U4010 | ~new_P2_U4011;
  assign n1444 = ~new_P2_U4006 | ~new_P2_U4007 | ~new_P2_U4008;
  assign n1439 = ~new_P2_U4003 | ~new_P2_U4004 | ~new_P2_U4005;
  assign n1434 = ~new_P2_U4000 | ~new_P2_U4001 | ~new_P2_U4002;
  assign n1429 = ~new_P2_U3997 | ~new_P2_U3998 | ~new_P2_U3999;
  assign n1424 = ~new_P2_U3994 | ~new_P2_U3995 | ~new_P2_U3996;
  assign n1419 = ~new_P2_U3991 | ~new_P2_U3992 | ~new_P2_U3993;
  assign n1414 = ~new_P2_U3988 | ~new_P2_U3989 | ~new_P2_U3990;
  assign n1409 = ~new_P2_U3985 | ~new_P2_U3986 | ~new_P2_U3987;
  assign n1404 = ~new_P2_U3982 | ~new_P2_U3983 | ~new_P2_U3984;
  assign n1399 = ~new_P2_U3979 | ~new_P2_U3980 | ~new_P2_U3981;
  assign n2459 = new_P2_U3797 & new_P2_U5641;
  assign new_P2_U3329 = ~P2_STATE_REG | ~new_P2_U3879;
  assign new_P2_U3330 = ~new_U69;
  assign new_P2_U3331 = ~P2_B_REG;
  assign new_P2_U3332 = ~new_P2_U3414 | ~new_P2_U5649;
  assign new_P2_U3333 = ~new_P2_U3414 | ~new_P2_U4075;
  assign new_P2_U3334 = ~new_P2_U3420 | ~new_P2_U5671 | ~new_P2_U3424;
  assign new_P2_U3335 = ~new_P2_U3420 | ~new_P2_U3418 | ~new_P2_U3424;
  assign new_P2_U3336 = ~new_P2_U3049 | ~new_P2_U3420;
  assign new_P2_U3337 = ~new_P2_U3419 | ~new_P2_U3418 | ~new_P2_U3424;
  assign new_P2_U3338 = ~new_P2_U3049 | ~new_P2_U3419;
  assign new_P2_U3339 = ~new_P2_U3420 | ~new_P2_U5668 | ~new_P2_U5674;
  assign new_P2_U3340 = ~new_P2_U5671 | ~new_P2_U5668;
  assign new_P2_U3341 = ~new_P2_U3974 | ~new_P2_U3419;
  assign new_P2_U3342 = ~new_P2_U3939 | ~new_P2_U5665;
  assign new_P2_U3343 = ~new_P2_U5665 | ~new_P2_U5674;
  assign new_P2_U3344 = ~new_P2_U3420 | ~new_P2_U3419;
  assign new_P2_U3345 = ~new_P2_U5665 | ~new_P2_U3424;
  assign new_P2_U3346 = ~new_P2_U3049 | ~new_P2_U5665;
  assign new_P2_U3347 = ~new_P2_U5688 | ~new_P2_U5683;
  assign new_P2_U3348 = ~new_P2_U3563 | ~new_P2_U3564 | ~new_P2_U4123;
  assign new_P2_U3349 = ~new_P2_U3580 | ~new_P2_U3578 | ~new_P2_U4141 | ~new_P2_U4140;
  assign new_P2_U3350 = ~new_P2_U3584 | ~new_P2_U3582 | ~new_P2_U4160 | ~new_P2_U4159;
  assign new_P2_U3351 = ~new_P2_U3588 | ~new_P2_U3586 | ~new_P2_U4179 | ~new_P2_U4178;
  assign new_P2_U3352 = ~new_P2_U3592 | ~new_P2_U3590 | ~new_P2_U4198 | ~new_P2_U4197;
  assign new_P2_U3353 = ~new_P2_U3596 | ~new_P2_U3594 | ~new_P2_U4217 | ~new_P2_U4216;
  assign new_P2_U3354 = ~new_P2_U3600 | ~new_P2_U3598 | ~new_P2_U4236 | ~new_P2_U4235;
  assign new_P2_U3355 = ~new_P2_U3604 | ~new_P2_U3602 | ~new_P2_U4255 | ~new_P2_U4254;
  assign new_P2_U3356 = ~new_P2_U3608 | ~new_P2_U3606 | ~new_P2_U4274 | ~new_P2_U4273;
  assign new_P2_U3357 = ~new_P2_U3612 | ~new_P2_U3610 | ~new_P2_U4293 | ~new_P2_U4292;
  assign new_P2_U3358 = ~new_P2_U3616 | ~new_P2_U3614 | ~new_P2_U4312 | ~new_P2_U4311;
  assign new_P2_U3359 = ~new_P2_U3620 | ~new_P2_U3618 | ~new_P2_U4331 | ~new_P2_U4330;
  assign new_P2_U3360 = ~new_P2_U3624 | ~new_P2_U3622 | ~new_P2_U4350 | ~new_P2_U4349;
  assign new_P2_U3361 = ~new_P2_U3628 | ~new_P2_U3626 | ~new_P2_U4369 | ~new_P2_U4368;
  assign new_P2_U3362 = ~new_P2_U3632 | ~new_P2_U3630 | ~new_P2_U4388 | ~new_P2_U4387;
  assign new_P2_U3363 = ~new_P2_U3636 | ~new_P2_U3634 | ~new_P2_U4407 | ~new_P2_U4406;
  assign new_P2_U3364 = ~new_P2_U3640 | ~new_P2_U3638 | ~new_P2_U4426 | ~new_P2_U4425;
  assign new_P2_U3365 = ~new_P2_U3644 | ~new_P2_U3642 | ~new_P2_U4445 | ~new_P2_U4444;
  assign new_P2_U3366 = ~new_P2_U3648 | ~new_P2_U3646 | ~new_P2_U4464 | ~new_P2_U4463;
  assign new_P2_U3367 = ~new_P2_U3652 | ~new_P2_U3650 | ~new_P2_U4483 | ~new_P2_U4482;
  assign new_P2_U3368 = ~new_U81 | ~new_P2_U3347;
  assign new_P2_U3369 = ~new_P2_U3656 | ~new_P2_U3654 | ~new_P2_U4502 | ~new_P2_U4501;
  assign new_P2_U3370 = ~new_U80 | ~new_P2_U3347;
  assign new_P2_U3371 = ~new_P2_U3660 | ~new_P2_U3658 | ~new_P2_U4521 | ~new_P2_U4520;
  assign new_P2_U3372 = ~new_U79 | ~new_P2_U3347;
  assign new_P2_U3373 = ~new_P2_U3664 | ~new_P2_U3662 | ~new_P2_U4540 | ~new_P2_U4539;
  assign new_P2_U3374 = ~new_U78 | ~new_P2_U3347;
  assign new_P2_U3375 = ~new_P2_U3668 | ~new_P2_U3666 | ~new_P2_U4559 | ~new_P2_U4558;
  assign new_P2_U3376 = ~new_U77 | ~new_P2_U3347;
  assign new_P2_U3377 = ~new_P2_U3672 | ~new_P2_U3670 | ~new_P2_U4578 | ~new_P2_U4577;
  assign new_P2_U3378 = ~new_U76 | ~new_P2_U3347;
  assign new_P2_U3379 = ~new_P2_U3676 | ~new_P2_U3674 | ~new_P2_U4597 | ~new_P2_U4596;
  assign new_P2_U3380 = ~new_U75 | ~new_P2_U3347;
  assign new_P2_U3381 = ~new_P2_U3680 | ~new_P2_U3678 | ~new_P2_U4616 | ~new_P2_U4615;
  assign new_P2_U3382 = ~new_U74 | ~new_P2_U3347;
  assign new_P2_U3383 = ~new_P2_U3684 | ~new_P2_U3682 | ~new_P2_U4635 | ~new_P2_U4634;
  assign new_P2_U3384 = ~new_U73 | ~new_P2_U3347;
  assign new_P2_U3385 = ~new_P2_U3687 | ~new_P2_U4656 | ~new_P2_U4655 | ~new_P2_U4654 | ~new_P2_U4653;
  assign new_P2_U3386 = ~new_U72 | ~new_P2_U3347;
  assign new_P2_U3387 = ~new_P2_U3692 | ~new_P2_U3690 | ~new_P2_U4675 | ~new_P2_U4674 | ~new_P2_U4673;
  assign new_P2_U3388 = ~new_U70 | ~new_P2_U3347;
  assign new_P2_U3389 = ~new_U69 | ~new_P2_U3347;
  assign new_P2_U3390 = ~new_P2_U3944 | ~new_P2_U3424;
  assign new_P2_U3391 = ~new_P2_U3023 | ~new_P2_U4698;
  assign new_P2_U3392 = ~new_P2_U3419 | ~new_P2_U5671 | ~new_P2_U3424;
  assign new_P2_U3393 = ~new_P2_U3921 | ~new_P2_U5671;
  assign new_P2_U3394 = ~new_P2_U3944 | ~new_P2_U5668;
  assign new_P2_U3395 = ~new_P2_U3927 | ~new_P2_U5671;
  assign new_P2_U3396 = ~new_P2_U3414 | ~new_P2_U3413 | ~new_P2_U3412;
  assign new_P2_U3397 = ~new_P2_U3344 | ~new_P2_U3347;
  assign new_P2_U3398 = ~new_P2_U3934 | ~new_P2_U4699;
  assign new_P2_U3399 = ~new_P2_U3962 | ~new_P2_U5658;
  assign new_P2_U3400 = ~new_P2_U3977 | ~P2_STATE_REG;
  assign new_P2_U3401 = ~new_P2_U3756 | ~new_P2_U3052;
  assign new_P2_U3402 = ~new_P2_U3974 | ~new_P2_U3420;
  assign new_P2_U3403 = ~new_P2_U3015 | ~new_P2_U3018;
  assign new_P2_U3404 = ~new_P2_U5674 | ~new_P2_U3424;
  assign new_P2_U3405 = ~new_P2_U3023 | ~new_P2_U3398;
  assign new_P2_U3406 = ~new_P2_U3798 | ~new_P2_U3016;
  assign new_P2_U3407 = ~new_P2_U3396 | ~new_P2_U5168 | ~P2_STATE_REG;
  assign new_P2_U3408 = ~new_P2_U3802 | ~new_P2_U5172;
  assign new_P2_U3409 = ~new_P2_R1299_U6;
  assign new_P2_U3410 = ~new_P2_U3938 | ~new_P2_U5665;
  assign new_P2_U3411 = ~new_P2_U3923 | ~new_P2_U3346 | ~new_P2_U3335 | ~new_P2_U3336;
  assign new_P2_U3412 = ~new_P2_U5645 | ~new_P2_U5644;
  assign new_P2_U3413 = ~new_P2_U5648 | ~new_P2_U5647;
  assign new_P2_U3414 = ~new_P2_U5651 | ~new_P2_U5650;
  assign new_P2_U3415 = ~new_P2_U5657 | ~new_P2_U5656;
  assign n1559 = ~new_P2_U5660 | ~new_P2_U5659;
  assign n1564 = ~new_P2_U5662 | ~new_P2_U5661;
  assign new_P2_U3418 = ~new_P2_U5670 | ~new_P2_U5669;
  assign new_P2_U3419 = ~new_P2_U5673 | ~new_P2_U5672;
  assign new_P2_U3420 = ~new_P2_U5664 | ~new_P2_U5663;
  assign new_P2_U3421 = ~new_P2_U5676 | ~new_P2_U5675;
  assign new_P2_U3422 = ~new_P2_U5679 | ~new_P2_U5678;
  assign new_P2_U3423 = ~new_P2_U5682 | ~new_P2_U5681;
  assign new_P2_U3424 = ~new_P2_U5667 | ~new_P2_U5666;
  assign new_P2_U3425 = ~new_P2_U5685 | ~new_P2_U5684;
  assign new_P2_U3426 = ~new_P2_U5687 | ~new_P2_U5686;
  assign new_P2_U3427 = ~new_P2_U5690 | ~new_P2_U5689;
  assign new_P2_U3428 = ~new_P2_U5698 | ~new_P2_U5697;
  assign new_P2_U3429 = ~new_P2_U5695 | ~new_P2_U5694;
  assign n1719 = ~new_P2_U5701 | ~new_P2_U5700;
  assign new_P2_U3431 = ~new_P2_U5703 | ~new_P2_U5702;
  assign new_P2_U3432 = ~new_P2_U5705 | ~new_P2_U5704;
  assign n1724 = ~new_P2_U5708 | ~new_P2_U5707;
  assign new_P2_U3434 = ~new_P2_U5710 | ~new_P2_U5709;
  assign new_P2_U3435 = ~new_P2_U5712 | ~new_P2_U5711;
  assign n1729 = ~new_P2_U5715 | ~new_P2_U5714;
  assign new_P2_U3437 = ~new_P2_U5717 | ~new_P2_U5716;
  assign new_P2_U3438 = ~new_P2_U5719 | ~new_P2_U5718;
  assign n1734 = ~new_P2_U5722 | ~new_P2_U5721;
  assign new_P2_U3440 = ~new_P2_U5724 | ~new_P2_U5723;
  assign new_P2_U3441 = ~new_P2_U5726 | ~new_P2_U5725;
  assign n1739 = ~new_P2_U5729 | ~new_P2_U5728;
  assign new_P2_U3443 = ~new_P2_U5731 | ~new_P2_U5730;
  assign new_P2_U3444 = ~new_P2_U5733 | ~new_P2_U5732;
  assign n1744 = ~new_P2_U5736 | ~new_P2_U5735;
  assign new_P2_U3446 = ~new_P2_U5738 | ~new_P2_U5737;
  assign new_P2_U3447 = ~new_P2_U5740 | ~new_P2_U5739;
  assign n1749 = ~new_P2_U5743 | ~new_P2_U5742;
  assign new_P2_U3449 = ~new_P2_U5745 | ~new_P2_U5744;
  assign new_P2_U3450 = ~new_P2_U5747 | ~new_P2_U5746;
  assign n1754 = ~new_P2_U5750 | ~new_P2_U5749;
  assign new_P2_U3452 = ~new_P2_U5752 | ~new_P2_U5751;
  assign new_P2_U3453 = ~new_P2_U5754 | ~new_P2_U5753;
  assign n1759 = ~new_P2_U5757 | ~new_P2_U5756;
  assign new_P2_U3455 = ~new_P2_U5759 | ~new_P2_U5758;
  assign new_P2_U3456 = ~new_P2_U5761 | ~new_P2_U5760;
  assign n1764 = ~new_P2_U5764 | ~new_P2_U5763;
  assign new_P2_U3458 = ~new_P2_U5766 | ~new_P2_U5765;
  assign new_P2_U3459 = ~new_P2_U5768 | ~new_P2_U5767;
  assign n1769 = ~new_P2_U5771 | ~new_P2_U5770;
  assign new_P2_U3461 = ~new_P2_U5773 | ~new_P2_U5772;
  assign new_P2_U3462 = ~new_P2_U5775 | ~new_P2_U5774;
  assign n1774 = ~new_P2_U5778 | ~new_P2_U5777;
  assign new_P2_U3464 = ~new_P2_U5780 | ~new_P2_U5779;
  assign new_P2_U3465 = ~new_P2_U5782 | ~new_P2_U5781;
  assign n1779 = ~new_P2_U5785 | ~new_P2_U5784;
  assign new_P2_U3467 = ~new_P2_U5787 | ~new_P2_U5786;
  assign new_P2_U3468 = ~new_P2_U5789 | ~new_P2_U5788;
  assign n1784 = ~new_P2_U5792 | ~new_P2_U5791;
  assign new_P2_U3470 = ~new_P2_U5794 | ~new_P2_U5793;
  assign new_P2_U3471 = ~new_P2_U5796 | ~new_P2_U5795;
  assign n1789 = ~new_P2_U5799 | ~new_P2_U5798;
  assign new_P2_U3473 = ~new_P2_U5801 | ~new_P2_U5800;
  assign new_P2_U3474 = ~new_P2_U5803 | ~new_P2_U5802;
  assign n1794 = ~new_P2_U5806 | ~new_P2_U5805;
  assign new_P2_U3476 = ~new_P2_U5808 | ~new_P2_U5807;
  assign new_P2_U3477 = ~new_P2_U5810 | ~new_P2_U5809;
  assign n1799 = ~new_P2_U5813 | ~new_P2_U5812;
  assign new_P2_U3479 = ~new_P2_U5815 | ~new_P2_U5814;
  assign new_P2_U3480 = ~new_P2_U5817 | ~new_P2_U5816;
  assign n1804 = ~new_P2_U5820 | ~new_P2_U5819;
  assign new_P2_U3482 = ~new_P2_U5822 | ~new_P2_U5821;
  assign new_P2_U3483 = ~new_P2_U5824 | ~new_P2_U5823;
  assign n1809 = ~new_P2_U5827 | ~new_P2_U5826;
  assign new_P2_U3485 = ~new_P2_U5829 | ~new_P2_U5828;
  assign n1814 = ~new_P2_U5832 | ~new_P2_U5831;
  assign n1819 = ~new_P2_U5834 | ~new_P2_U5833;
  assign n1824 = ~new_P2_U5836 | ~new_P2_U5835;
  assign n1829 = ~new_P2_U5838 | ~new_P2_U5837;
  assign n1834 = ~new_P2_U5840 | ~new_P2_U5839;
  assign n1839 = ~new_P2_U5842 | ~new_P2_U5841;
  assign n1844 = ~new_P2_U5844 | ~new_P2_U5843;
  assign n1849 = ~new_P2_U5846 | ~new_P2_U5845;
  assign n1854 = ~new_P2_U5848 | ~new_P2_U5847;
  assign n1859 = ~new_P2_U5850 | ~new_P2_U5849;
  assign n1864 = ~new_P2_U5852 | ~new_P2_U5851;
  assign n1869 = ~new_P2_U5854 | ~new_P2_U5853;
  assign n1874 = ~new_P2_U5856 | ~new_P2_U5855;
  assign n1879 = ~new_P2_U5858 | ~new_P2_U5857;
  assign n1884 = ~new_P2_U5860 | ~new_P2_U5859;
  assign n1889 = ~new_P2_U5862 | ~new_P2_U5861;
  assign n1894 = ~new_P2_U5864 | ~new_P2_U5863;
  assign n1899 = ~new_P2_U5866 | ~new_P2_U5865;
  assign n1904 = ~new_P2_U5868 | ~new_P2_U5867;
  assign n1909 = ~new_P2_U5870 | ~new_P2_U5869;
  assign n1914 = ~new_P2_U5872 | ~new_P2_U5871;
  assign n1919 = ~new_P2_U5874 | ~new_P2_U5873;
  assign n1924 = ~new_P2_U5876 | ~new_P2_U5875;
  assign n1929 = ~new_P2_U5878 | ~new_P2_U5877;
  assign n1934 = ~new_P2_U5880 | ~new_P2_U5879;
  assign n1939 = ~new_P2_U5882 | ~new_P2_U5881;
  assign n1944 = ~new_P2_U5884 | ~new_P2_U5883;
  assign n1949 = ~new_P2_U5886 | ~new_P2_U5885;
  assign n1954 = ~new_P2_U5888 | ~new_P2_U5887;
  assign n1959 = ~new_P2_U5890 | ~new_P2_U5889;
  assign n1964 = ~new_P2_U5892 | ~new_P2_U5891;
  assign n1969 = ~new_P2_U5894 | ~new_P2_U5893;
  assign n1974 = ~new_P2_U5896 | ~new_P2_U5895;
  assign n1979 = ~new_P2_U5898 | ~new_P2_U5897;
  assign n1984 = ~new_P2_U5900 | ~new_P2_U5899;
  assign n1989 = ~new_P2_U5902 | ~new_P2_U5901;
  assign n1994 = ~new_P2_U5904 | ~new_P2_U5903;
  assign n1999 = ~new_P2_U5906 | ~new_P2_U5905;
  assign n2004 = ~new_P2_U5908 | ~new_P2_U5907;
  assign n2009 = ~new_P2_U5910 | ~new_P2_U5909;
  assign n2014 = ~new_P2_U5912 | ~new_P2_U5911;
  assign n2019 = ~new_P2_U5914 | ~new_P2_U5913;
  assign n2024 = ~new_P2_U5916 | ~new_P2_U5915;
  assign n2029 = ~new_P2_U5918 | ~new_P2_U5917;
  assign n2034 = ~new_P2_U5920 | ~new_P2_U5919;
  assign n2299 = ~new_P2_U5986 | ~new_P2_U5985;
  assign n2304 = ~new_P2_U5988 | ~new_P2_U5987;
  assign n2309 = ~new_P2_U5990 | ~new_P2_U5989;
  assign n2314 = ~new_P2_U5992 | ~new_P2_U5991;
  assign n2319 = ~new_P2_U5994 | ~new_P2_U5993;
  assign n2324 = ~new_P2_U5996 | ~new_P2_U5995;
  assign n2329 = ~new_P2_U5998 | ~new_P2_U5997;
  assign n2334 = ~new_P2_U6000 | ~new_P2_U5999;
  assign n2339 = ~new_P2_U6002 | ~new_P2_U6001;
  assign n2344 = ~new_P2_U6004 | ~new_P2_U6003;
  assign n2349 = ~new_P2_U6006 | ~new_P2_U6005;
  assign n2354 = ~new_P2_U6008 | ~new_P2_U6007;
  assign n2359 = ~new_P2_U6010 | ~new_P2_U6009;
  assign n2364 = ~new_P2_U6012 | ~new_P2_U6011;
  assign n2369 = ~new_P2_U6014 | ~new_P2_U6013;
  assign n2374 = ~new_P2_U6016 | ~new_P2_U6015;
  assign n2379 = ~new_P2_U6018 | ~new_P2_U6017;
  assign n2384 = ~new_P2_U6020 | ~new_P2_U6019;
  assign n2389 = ~new_P2_U6022 | ~new_P2_U6021;
  assign n2394 = ~new_P2_U6024 | ~new_P2_U6023;
  assign n2399 = ~new_P2_U6026 | ~new_P2_U6025;
  assign n2404 = ~new_P2_U6028 | ~new_P2_U6027;
  assign n2409 = ~new_P2_U6030 | ~new_P2_U6029;
  assign n2414 = ~new_P2_U6032 | ~new_P2_U6031;
  assign n2419 = ~new_P2_U6034 | ~new_P2_U6033;
  assign n2424 = ~new_P2_U6036 | ~new_P2_U6035;
  assign n2429 = ~new_P2_U6038 | ~new_P2_U6037;
  assign n2434 = ~new_P2_U6040 | ~new_P2_U6039;
  assign n2439 = ~new_P2_U6042 | ~new_P2_U6041;
  assign n2444 = ~new_P2_U6044 | ~new_P2_U6043;
  assign n2449 = ~new_P2_U6046 | ~new_P2_U6045;
  assign n2454 = ~new_P2_U6048 | ~new_P2_U6047;
  assign new_P2_U3563 = new_P2_U4117 & new_P2_U4118 & new_P2_U4120 & new_P2_U4119;
  assign new_P2_U3564 = new_P2_U4122 & new_P2_U4121;
  assign new_P2_U3565 = new_P2_U4127 & new_P2_U4125;
  assign new_P2_U3566 = new_P2_U4079 & new_P2_U4080 & new_P2_U4082 & new_P2_U4081;
  assign new_P2_U3567 = new_P2_U4083 & new_P2_U4084 & new_P2_U4086 & new_P2_U4085;
  assign new_P2_U3568 = new_P2_U4087 & new_P2_U4088 & new_P2_U4090 & new_P2_U4089;
  assign new_P2_U3569 = new_P2_U4093 & new_P2_U4092 & new_P2_U4091;
  assign new_P2_U3570 = new_P2_U3566 & new_P2_U3567 & new_P2_U3569 & new_P2_U3568;
  assign new_P2_U3571 = new_P2_U4094 & new_P2_U4095 & new_P2_U4097 & new_P2_U4096;
  assign new_P2_U3572 = new_P2_U4098 & new_P2_U4099 & new_P2_U4101 & new_P2_U4100;
  assign new_P2_U3573 = new_P2_U4102 & new_P2_U4103 & new_P2_U4105 & new_P2_U4104;
  assign new_P2_U3574 = new_P2_U4108 & new_P2_U4107 & new_P2_U4106;
  assign new_P2_U3575 = new_P2_U3571 & new_P2_U3572 & new_P2_U3574 & new_P2_U3573;
  assign new_P2_U3576 = new_P2_U5696 & new_P2_U4110;
  assign new_P2_U3577 = new_P2_U5699 & new_P2_U3023;
  assign new_P2_U3578 = new_P2_U4143 & new_P2_U4142;
  assign new_P2_U3579 = new_P2_U4145 & new_P2_U4144;
  assign new_P2_U3580 = new_P2_U3579 & new_P2_U4147 & new_P2_U4146;
  assign new_P2_U3581 = new_P2_U4151 & new_P2_U4152 & new_P2_U4150 & new_P2_U4149;
  assign new_P2_U3582 = new_P2_U4162 & new_P2_U4161;
  assign new_P2_U3583 = new_P2_U4164 & new_P2_U4163;
  assign new_P2_U3584 = new_P2_U3583 & new_P2_U4166 & new_P2_U4165;
  assign new_P2_U3585 = new_P2_U4170 & new_P2_U4171 & new_P2_U4169 & new_P2_U4168;
  assign new_P2_U3586 = new_P2_U4181 & new_P2_U4180;
  assign new_P2_U3587 = new_P2_U4183 & new_P2_U4182;
  assign new_P2_U3588 = new_P2_U3587 & new_P2_U4185 & new_P2_U4184;
  assign new_P2_U3589 = new_P2_U4189 & new_P2_U4190 & new_P2_U4188 & new_P2_U4187;
  assign new_P2_U3590 = new_P2_U4200 & new_P2_U4199;
  assign new_P2_U3591 = new_P2_U4202 & new_P2_U4201;
  assign new_P2_U3592 = new_P2_U3591 & new_P2_U4204 & new_P2_U4203;
  assign new_P2_U3593 = new_P2_U4208 & new_P2_U4209 & new_P2_U4207 & new_P2_U4206;
  assign new_P2_U3594 = new_P2_U4219 & new_P2_U4218;
  assign new_P2_U3595 = new_P2_U4221 & new_P2_U4220;
  assign new_P2_U3596 = new_P2_U3595 & new_P2_U4223 & new_P2_U4222;
  assign new_P2_U3597 = new_P2_U4227 & new_P2_U4228 & new_P2_U4226 & new_P2_U4225;
  assign new_P2_U3598 = new_P2_U4238 & new_P2_U4237;
  assign new_P2_U3599 = new_P2_U4240 & new_P2_U4239;
  assign new_P2_U3600 = new_P2_U3599 & new_P2_U4242 & new_P2_U4241;
  assign new_P2_U3601 = new_P2_U4246 & new_P2_U4247 & new_P2_U4245 & new_P2_U4244;
  assign new_P2_U3602 = new_P2_U4257 & new_P2_U4256;
  assign new_P2_U3603 = new_P2_U4259 & new_P2_U4258;
  assign new_P2_U3604 = new_P2_U3603 & new_P2_U4261 & new_P2_U4260;
  assign new_P2_U3605 = new_P2_U4265 & new_P2_U4266 & new_P2_U4264 & new_P2_U4263;
  assign new_P2_U3606 = new_P2_U4276 & new_P2_U4275;
  assign new_P2_U3607 = new_P2_U4278 & new_P2_U4277;
  assign new_P2_U3608 = new_P2_U3607 & new_P2_U4280 & new_P2_U4279;
  assign new_P2_U3609 = new_P2_U4284 & new_P2_U4285 & new_P2_U4283 & new_P2_U4282;
  assign new_P2_U3610 = new_P2_U4295 & new_P2_U4294;
  assign new_P2_U3611 = new_P2_U4297 & new_P2_U4296;
  assign new_P2_U3612 = new_P2_U3611 & new_P2_U4299 & new_P2_U4298;
  assign new_P2_U3613 = new_P2_U4303 & new_P2_U4304 & new_P2_U4302 & new_P2_U4301;
  assign new_P2_U3614 = new_P2_U4314 & new_P2_U4313;
  assign new_P2_U3615 = new_P2_U4316 & new_P2_U4315;
  assign new_P2_U3616 = new_P2_U3615 & new_P2_U4318 & new_P2_U4317;
  assign new_P2_U3617 = new_P2_U4322 & new_P2_U4323 & new_P2_U4321 & new_P2_U4320;
  assign new_P2_U3618 = new_P2_U4333 & new_P2_U4332;
  assign new_P2_U3619 = new_P2_U4335 & new_P2_U4334;
  assign new_P2_U3620 = new_P2_U3619 & new_P2_U4337 & new_P2_U4336;
  assign new_P2_U3621 = new_P2_U4341 & new_P2_U4342 & new_P2_U4340 & new_P2_U4339;
  assign new_P2_U3622 = new_P2_U4352 & new_P2_U4351;
  assign new_P2_U3623 = new_P2_U4354 & new_P2_U4353;
  assign new_P2_U3624 = new_P2_U3623 & new_P2_U4356 & new_P2_U4355;
  assign new_P2_U3625 = new_P2_U4360 & new_P2_U4361 & new_P2_U4359 & new_P2_U4358;
  assign new_P2_U3626 = new_P2_U4371 & new_P2_U4370;
  assign new_P2_U3627 = new_P2_U4373 & new_P2_U4372;
  assign new_P2_U3628 = new_P2_U3627 & new_P2_U4375 & new_P2_U4374;
  assign new_P2_U3629 = new_P2_U4379 & new_P2_U4380 & new_P2_U4378 & new_P2_U4377;
  assign new_P2_U3630 = new_P2_U4390 & new_P2_U4389;
  assign new_P2_U3631 = new_P2_U4392 & new_P2_U4391;
  assign new_P2_U3632 = new_P2_U3631 & new_P2_U4394 & new_P2_U4393;
  assign new_P2_U3633 = new_P2_U4398 & new_P2_U4399 & new_P2_U4397 & new_P2_U4396;
  assign new_P2_U3634 = new_P2_U4409 & new_P2_U4408;
  assign new_P2_U3635 = new_P2_U4411 & new_P2_U4410;
  assign new_P2_U3636 = new_P2_U3635 & new_P2_U4413 & new_P2_U4412;
  assign new_P2_U3637 = new_P2_U4417 & new_P2_U4418 & new_P2_U4416 & new_P2_U4415;
  assign new_P2_U3638 = new_P2_U4428 & new_P2_U4427;
  assign new_P2_U3639 = new_P2_U4430 & new_P2_U4429;
  assign new_P2_U3640 = new_P2_U3639 & new_P2_U4432 & new_P2_U4431;
  assign new_P2_U3641 = new_P2_U4436 & new_P2_U4437 & new_P2_U4435 & new_P2_U4434;
  assign new_P2_U3642 = new_P2_U4447 & new_P2_U4446;
  assign new_P2_U3643 = new_P2_U4449 & new_P2_U4448;
  assign new_P2_U3644 = new_P2_U3643 & new_P2_U4451 & new_P2_U4450;
  assign new_P2_U3645 = new_P2_U4455 & new_P2_U4456 & new_P2_U4454 & new_P2_U4453;
  assign new_P2_U3646 = new_P2_U4466 & new_P2_U4465;
  assign new_P2_U3647 = new_P2_U4468 & new_P2_U4467;
  assign new_P2_U3648 = new_P2_U3647 & new_P2_U4470 & new_P2_U4469;
  assign new_P2_U3649 = new_P2_U4474 & new_P2_U4475 & new_P2_U4473 & new_P2_U4472;
  assign new_P2_U3650 = new_P2_U4485 & new_P2_U4484;
  assign new_P2_U3651 = new_P2_U4487 & new_P2_U4486;
  assign new_P2_U3652 = new_P2_U3651 & new_P2_U4489 & new_P2_U4488;
  assign new_P2_U3653 = new_P2_U4493 & new_P2_U4494 & new_P2_U4492 & new_P2_U4491;
  assign new_P2_U3654 = new_P2_U4504 & new_P2_U4503;
  assign new_P2_U3655 = new_P2_U4506 & new_P2_U4505;
  assign new_P2_U3656 = new_P2_U3655 & new_P2_U4508 & new_P2_U4507;
  assign new_P2_U3657 = new_P2_U4512 & new_P2_U4513 & new_P2_U4511 & new_P2_U4510;
  assign new_P2_U3658 = new_P2_U4523 & new_P2_U4522;
  assign new_P2_U3659 = new_P2_U4525 & new_P2_U4524;
  assign new_P2_U3660 = new_P2_U3659 & new_P2_U4527 & new_P2_U4526;
  assign new_P2_U3661 = new_P2_U4531 & new_P2_U4532 & new_P2_U4530 & new_P2_U4529;
  assign new_P2_U3662 = new_P2_U4542 & new_P2_U4541;
  assign new_P2_U3663 = new_P2_U4544 & new_P2_U4543;
  assign new_P2_U3664 = new_P2_U3663 & new_P2_U4546 & new_P2_U4545;
  assign new_P2_U3665 = new_P2_U4550 & new_P2_U4551 & new_P2_U4549 & new_P2_U4548;
  assign new_P2_U3666 = new_P2_U4561 & new_P2_U4560;
  assign new_P2_U3667 = new_P2_U4563 & new_P2_U4562;
  assign new_P2_U3668 = new_P2_U3667 & new_P2_U4565 & new_P2_U4564;
  assign new_P2_U3669 = new_P2_U4569 & new_P2_U4570 & new_P2_U4568 & new_P2_U4567;
  assign new_P2_U3670 = new_P2_U4580 & new_P2_U4579;
  assign new_P2_U3671 = new_P2_U4582 & new_P2_U4581;
  assign new_P2_U3672 = new_P2_U3671 & new_P2_U4584 & new_P2_U4583;
  assign new_P2_U3673 = new_P2_U4588 & new_P2_U4589 & new_P2_U4587 & new_P2_U4586;
  assign new_P2_U3674 = new_P2_U4599 & new_P2_U4598;
  assign new_P2_U3675 = new_P2_U4601 & new_P2_U4600;
  assign new_P2_U3676 = new_P2_U3675 & new_P2_U4603 & new_P2_U4602;
  assign new_P2_U3677 = new_P2_U4607 & new_P2_U4608 & new_P2_U4606 & new_P2_U4605;
  assign new_P2_U3678 = new_P2_U4618 & new_P2_U4617;
  assign new_P2_U3679 = new_P2_U4620 & new_P2_U4619;
  assign new_P2_U3680 = new_P2_U3679 & new_P2_U4622 & new_P2_U4621;
  assign new_P2_U3681 = new_P2_U4626 & new_P2_U4627 & new_P2_U4625 & new_P2_U4624;
  assign new_P2_U3682 = new_P2_U4637 & new_P2_U4636;
  assign new_P2_U3683 = new_P2_U4639 & new_P2_U4638;
  assign new_P2_U3684 = new_P2_U3683 & new_P2_U4641 & new_P2_U4640;
  assign new_P2_U3685 = new_P2_U4645 & new_P2_U4646 & new_P2_U4644 & new_P2_U4643;
  assign new_P2_U3686 = new_P2_U4658 & new_P2_U4657;
  assign new_P2_U3687 = new_P2_U3686 & new_P2_U4660 & new_P2_U4659;
  assign new_P2_U3688 = new_P2_U4664 & new_P2_U4665 & new_P2_U4663 & new_P2_U4662;
  assign new_P2_U3689 = new_P2_U4672 & new_P2_U3963;
  assign new_P2_U3690 = new_P2_U4677 & new_P2_U4676;
  assign new_P2_U3691 = new_P2_U4679 & new_P2_U4678;
  assign new_P2_U3692 = new_P2_U3691 & new_P2_U4681 & new_P2_U4680;
  assign new_P2_U3693 = new_P2_U4684 & new_P2_U4685 & new_P2_U4683;
  assign new_P2_U3694 = new_P2_U3963 & new_P2_U4672;
  assign new_P2_U3695 = new_P2_U3023 & new_P2_U3428;
  assign new_P2_U3696 = new_P2_U3429 & new_P2_U5699 & new_P2_U3935;
  assign new_P2_U3697 = new_P2_U4703 & new_P2_U4702 & new_P2_U4701;
  assign new_P2_U3698 = new_P2_U3883 & new_P2_U4705 & new_P2_U4704;
  assign new_P2_U3699 = new_P2_U4708 & new_P2_U4707 & new_P2_U4706;
  assign new_P2_U3700 = new_P2_U3884 & new_P2_U4710 & new_P2_U4709;
  assign new_P2_U3701 = new_P2_U4713 & new_P2_U4712 & new_P2_U4711;
  assign new_P2_U3702 = new_P2_U3885 & new_P2_U4715 & new_P2_U4714;
  assign new_P2_U3703 = new_P2_U4718 & new_P2_U4717 & new_P2_U4716;
  assign new_P2_U3704 = new_P2_U3886 & new_P2_U4720 & new_P2_U4719;
  assign new_P2_U3705 = new_P2_U4723 & new_P2_U4722 & new_P2_U4721;
  assign new_P2_U3706 = new_P2_U3887 & new_P2_U4725 & new_P2_U4724;
  assign new_P2_U3707 = new_P2_U4728 & new_P2_U4727 & new_P2_U4726;
  assign new_P2_U3708 = new_P2_U3888 & new_P2_U4730 & new_P2_U4729;
  assign new_P2_U3709 = new_P2_U4733 & new_P2_U4732 & new_P2_U4731;
  assign new_P2_U3710 = new_P2_U3889 & new_P2_U4735 & new_P2_U4734;
  assign new_P2_U3711 = new_P2_U4738 & new_P2_U4737 & new_P2_U4736;
  assign new_P2_U3712 = new_P2_U3890 & new_P2_U4740 & new_P2_U4739;
  assign new_P2_U3713 = new_P2_U4743 & new_P2_U4742 & new_P2_U4741;
  assign new_P2_U3714 = new_P2_U3891 & new_P2_U4745 & new_P2_U4744;
  assign new_P2_U3715 = new_P2_U4748 & new_P2_U4747 & new_P2_U4746;
  assign new_P2_U3716 = new_P2_U3892 & new_P2_U4750 & new_P2_U4749;
  assign new_P2_U3717 = new_P2_U4753 & new_P2_U4752 & new_P2_U4751;
  assign new_P2_U3718 = new_P2_U4755 & new_P2_U4754;
  assign new_P2_U3719 = new_P2_U4758 & new_P2_U4757 & new_P2_U4756;
  assign new_P2_U3720 = new_P2_U4760 & new_P2_U4759;
  assign new_P2_U3721 = new_P2_U4763 & new_P2_U4762 & new_P2_U4761;
  assign new_P2_U3722 = new_P2_U4765 & new_P2_U4764;
  assign new_P2_U3723 = new_P2_U4767 & new_P2_U4768 & new_P2_U4766;
  assign new_P2_U3724 = new_P2_U4770 & new_P2_U4769;
  assign new_P2_U3725 = new_P2_U4773 & new_P2_U4772 & new_P2_U4771;
  assign new_P2_U3726 = new_P2_U4775 & new_P2_U4774;
  assign new_P2_U3727 = new_P2_U4777 & new_P2_U4778 & new_P2_U4776;
  assign new_P2_U3728 = new_P2_U4780 & new_P2_U4779;
  assign new_P2_U3729 = new_P2_U4783 & new_P2_U4781;
  assign new_P2_U3730 = new_P2_U4785 & new_P2_U4784;
  assign new_P2_U3731 = new_P2_U4788 & new_P2_U4786;
  assign new_P2_U3732 = new_P2_U4790 & new_P2_U4789;
  assign new_P2_U3733 = new_P2_U4793 & new_P2_U4791;
  assign new_P2_U3734 = new_P2_U4795 & new_P2_U4794;
  assign new_P2_U3735 = new_P2_U4798 & new_P2_U4796;
  assign new_P2_U3736 = new_P2_U4800 & new_P2_U4799;
  assign new_P2_U3737 = new_P2_U4803 & new_P2_U4801;
  assign new_P2_U3738 = new_P2_U4805 & new_P2_U4804;
  assign new_P2_U3739 = new_P2_U4808 & new_P2_U4806;
  assign new_P2_U3740 = new_P2_U4810 & new_P2_U4809;
  assign new_P2_U3741 = new_P2_U4813 & new_P2_U4811;
  assign new_P2_U3742 = new_P2_U4815 & new_P2_U4814;
  assign new_P2_U3743 = new_P2_U4818 & new_P2_U4816;
  assign new_P2_U3744 = new_P2_U4820 & new_P2_U4819;
  assign new_P2_U3745 = new_P2_U4823 & new_P2_U4821;
  assign new_P2_U3746 = new_P2_U4825 & new_P2_U4824;
  assign new_P2_U3747 = new_P2_U4828 & new_P2_U4826;
  assign new_P2_U3748 = new_P2_U4830 & new_P2_U4829;
  assign new_P2_U3749 = new_P2_U4833 & new_P2_U4831;
  assign new_P2_U3750 = new_P2_U4835 & new_P2_U4834;
  assign new_P2_U3751 = new_P2_U4838 & new_P2_U4836;
  assign new_P2_U3752 = new_P2_U4840 & new_P2_U4839;
  assign new_P2_U3753 = new_P2_U4843 & new_P2_U4841;
  assign new_P2_U3754 = new_P2_U4845 & new_P2_U4844;
  assign new_P2_U3755 = new_P2_U3334 & new_P2_U3335 & new_P2_U3336;
  assign new_P2_U3756 = new_P2_U5643 & new_P2_U3397;
  assign new_P2_U3757 = new_P2_U3415 & P2_STATE_REG;
  assign new_P2_U3758 = new_P2_U4866 & new_P2_U4867 & new_P2_U4869 & new_P2_U4870 & new_P2_U4868;
  assign new_P2_U3759 = new_P2_U4881 & new_P2_U4882 & new_P2_U4884 & new_P2_U4885 & new_P2_U4883;
  assign new_P2_U3760 = new_P2_U4896 & new_P2_U4897 & new_P2_U4899 & new_P2_U4900 & new_P2_U4898;
  assign new_P2_U3761 = new_P2_U4911 & new_P2_U4912 & new_P2_U4914 & new_P2_U4915 & new_P2_U4913;
  assign new_P2_U3762 = new_P2_U4926 & new_P2_U4927 & new_P2_U4929 & new_P2_U4930 & new_P2_U4928;
  assign new_P2_U3763 = new_P2_U4941 & new_P2_U4942 & new_P2_U4944 & new_P2_U4945 & new_P2_U4943;
  assign new_P2_U3764 = new_P2_U4956 & new_P2_U4957 & new_P2_U4959 & new_P2_U4960 & new_P2_U4958;
  assign new_P2_U3765 = new_P2_U4971 & new_P2_U4972 & new_P2_U4974 & new_P2_U4975 & new_P2_U4973;
  assign new_P2_U3766 = new_P2_U4986 & new_P2_U4987 & new_P2_U4990 & new_P2_U4989 & new_P2_U4988;
  assign new_P2_U3767 = new_P2_U5001 & new_P2_U5002 & new_P2_U5004 & new_P2_U5005 & new_P2_U5003;
  assign new_P2_U3768 = new_P2_U5016 & new_P2_U5017 & new_P2_U5020 & new_P2_U5019 & new_P2_U5018;
  assign new_P2_U3769 = new_P2_U5032 & new_P2_U5031;
  assign new_P2_U3770 = new_P2_U5035 & new_P2_U5034 & new_P2_U5033;
  assign new_P2_U3771 = new_P2_U5047 & new_P2_U5046;
  assign new_P2_U3772 = new_P2_U5050 & new_P2_U5049 & new_P2_U5048;
  assign new_P2_U3773 = new_P2_U5062 & new_P2_U5061;
  assign new_P2_U3774 = new_P2_U5065 & new_P2_U5064 & new_P2_U5063;
  assign new_P2_U3775 = new_P2_U5077 & new_P2_U5076;
  assign new_P2_U3776 = new_P2_U5080 & new_P2_U5079 & new_P2_U5078;
  assign new_P2_U3777 = new_P2_U5092 & new_P2_U5091;
  assign new_P2_U3778 = new_P2_U5095 & new_P2_U5094 & new_P2_U5093;
  assign new_P2_U3779 = new_P2_U5107 & new_P2_U5106;
  assign new_P2_U3780 = new_P2_U5110 & new_P2_U5109 & new_P2_U5108;
  assign new_P2_U3781 = new_P2_U5122 & new_P2_U5121;
  assign new_P2_U3782 = new_P2_U5125 & new_P2_U5124 & new_P2_U5123;
  assign new_P2_U3783 = new_P2_U5137 & new_P2_U5136;
  assign new_P2_U3784 = new_P2_U5140 & new_P2_U5139 & new_P2_U5138;
  assign new_P2_U3785 = new_P2_U5152 & new_P2_U5151;
  assign new_P2_U3786 = new_P2_U5155 & new_P2_U5154 & new_P2_U5153;
  assign new_P2_U3787 = new_P2_U5639 & new_P2_U5658;
  assign new_P2_U3788 = new_P2_U6106 & new_P2_U6103 & new_P2_U6100;
  assign new_P2_U3789 = new_P2_U6088 & new_P2_U6091 & new_P2_U6097 & new_P2_U6094;
  assign new_P2_U3790 = new_P2_U6112 & new_P2_U6115 & new_P2_U6121 & new_P2_U6118;
  assign new_P2_U3791 = new_P2_U6133 & new_P2_U6130 & new_P2_U6127 & new_P2_U6124;
  assign new_P2_U3792 = new_P2_U3790 & new_P2_U3791 & new_P2_U6109 & new_P2_U3788 & new_P2_U3789;
  assign new_P2_U3793 = new_P2_U6055 & new_P2_U6058 & new_P2_U6061 & new_P2_U3796 & new_P2_U3795;
  assign new_P2_U3794 = new_P2_U6148 & new_P2_U6136 & new_P2_U6139 & new_P2_U6145 & new_P2_U6142;
  assign new_P2_U3795 = new_P2_U6064 & new_P2_U6067 & new_P2_U6073 & new_P2_U6070;
  assign new_P2_U3796 = new_P2_U6079 & new_P2_U6076;
  assign new_P2_U3797 = new_P2_U5640 & new_P2_U5631;
  assign new_P2_U3798 = new_P2_U3428 & new_P2_U3429;
  assign new_P2_U3799 = new_P2_U3339 & new_P2_U3928;
  assign new_P2_U3800 = new_P2_U3799 & new_P2_U3342;
  assign new_P2_U3801 = new_P2_U3395 & new_P2_U3410;
  assign new_P2_U3802 = new_P2_U3399 & new_P2_U5658 & new_P2_U3935;
  assign new_P2_U3803 = new_P2_U3023 & new_P2_U5171;
  assign new_P2_U3804 = new_P2_U5198 & new_P2_U5196;
  assign new_P2_U3805 = new_P2_U5216 & new_P2_U5214;
  assign new_P2_U3806 = new_P2_U3969 & new_P2_U3080;
  assign new_P2_U3807 = new_P2_U5259 & new_P2_U5258;
  assign new_P2_U3808 = new_P2_U5262 & new_P2_U5261;
  assign new_P2_U3809 = new_P2_U5278 & new_P2_U5276;
  assign new_P2_U3810 = new_P2_U5305 & new_P2_U5303;
  assign new_P2_U3811 = new_P2_U5350 & new_P2_U5348;
  assign new_P2_U3812 = new_P2_U5359 & new_P2_U5357;
  assign new_P2_U3813 = new_P2_U5386 & new_P2_U5384;
  assign new_P2_U3814 = new_P2_U5431 & new_P2_U5429;
  assign new_P2_U3815 = new_P2_U5435 & P2_STATE_REG;
  assign new_P2_U3816 = new_P2_U3920 & new_P2_U3919 & new_P2_U3936;
  assign new_P2_U3817 = new_P2_U5671 & new_P2_U3419;
  assign new_P2_U3818 = new_P2_U3394 & new_P2_U3339;
  assign new_P2_U3819 = new_P2_U3818 & new_P2_U3342 & new_P2_U3390;
  assign new_P2_U3820 = new_P2_U3334 & new_P2_U3928;
  assign new_P2_U3821 = new_P2_U3415 & new_P2_U5444;
  assign new_P2_U3822 = new_P2_U3415 & new_P2_U5447;
  assign new_P2_U3823 = new_P2_U3415 & new_P2_U5450;
  assign new_P2_U3824 = new_P2_U3415 & new_P2_U5453;
  assign new_P2_U3825 = new_P2_U3415 & new_P2_U5456;
  assign new_P2_U3826 = new_P2_U3827 & new_P2_U5457;
  assign new_P2_U3827 = new_P2_U3415 & new_P2_U5459;
  assign new_P2_U3828 = new_P2_U5460 & new_P2_U3410;
  assign new_P2_U3829 = new_P2_U3830 & new_P2_U5465;
  assign new_P2_U3830 = new_P2_U3415 & new_P2_U5467;
  assign new_P2_U3831 = new_P2_U3415 & new_P2_U5468;
  assign new_P2_U3832 = new_P2_U3415 & new_P2_U5471;
  assign new_P2_U3833 = new_P2_U3415 & new_P2_U5474;
  assign new_P2_U3834 = new_P2_U3415 & new_P2_U5477;
  assign new_P2_U3835 = new_P2_U3415 & new_P2_U5480;
  assign new_P2_U3836 = new_P2_U3415 & new_P2_U5483;
  assign new_P2_U3837 = new_P2_U3415 & new_P2_U5486;
  assign new_P2_U3838 = new_P2_U3415 & new_P2_U5489;
  assign new_P2_U3839 = new_P2_U3415 & new_P2_U5492;
  assign new_P2_U3840 = new_P2_U3415 & new_P2_U5495;
  assign new_P2_U3841 = new_P2_U3842 & new_P2_U5498;
  assign new_P2_U3842 = new_P2_U3415 & new_P2_U5500;
  assign new_P2_U3843 = new_P2_U3415 & new_P2_U5501;
  assign new_P2_U3844 = new_P2_U3415 & new_P2_U5504;
  assign new_P2_U3845 = new_P2_U3415 & new_P2_U5507;
  assign new_P2_U3846 = new_P2_U3415 & new_P2_U5510;
  assign new_P2_U3847 = new_P2_U3415 & new_P2_U5513;
  assign new_P2_U3848 = new_P2_U3415 & new_P2_U5516;
  assign new_P2_U3849 = new_P2_U3415 & new_P2_U5519;
  assign new_P2_U3850 = new_P2_U3415 & new_P2_U5522;
  assign new_P2_U3851 = new_P2_U3415 & new_P2_U5527;
  assign new_P2_U3852 = new_P2_U3415 & new_P2_U5530;
  assign new_P2_U3853 = new_P2_U3854 & new_P2_U5531;
  assign new_P2_U3854 = new_P2_U3415 & new_P2_U5533;
  assign new_P2_U3855 = new_P2_U3856 & new_P2_U5534;
  assign new_P2_U3856 = new_P2_U3415 & new_P2_U5536;
  assign new_P2_U3857 = new_P2_U5539 & new_P2_U5540;
  assign new_P2_U3858 = new_P2_U5542 & new_P2_U5543;
  assign new_P2_U3859 = new_P2_U5564 & new_P2_U5565;
  assign new_P2_U3860 = new_P2_U5567 & new_P2_U5568;
  assign new_P2_U3861 = new_P2_U5570 & new_P2_U5571;
  assign new_P2_U3862 = new_P2_U5573 & new_P2_U5574;
  assign new_P2_U3863 = new_P2_U5576 & new_P2_U5577;
  assign new_P2_U3864 = new_P2_U5579 & new_P2_U5580;
  assign new_P2_U3865 = new_P2_U5582 & new_P2_U5583;
  assign new_P2_U3866 = new_P2_U5585 & new_P2_U5586;
  assign new_P2_U3867 = new_P2_U5588 & new_P2_U5589;
  assign new_P2_U3868 = new_P2_U5591 & new_P2_U5592;
  assign new_P2_U3869 = new_P2_U5597 & new_P2_U5598;
  assign new_P2_U3870 = new_P2_U5600 & new_P2_U5601;
  assign new_P2_U3871 = new_P2_U5603 & new_P2_U5604;
  assign new_P2_U3872 = new_P2_U5606 & new_P2_U5607;
  assign new_P2_U3873 = new_P2_U5609 & new_P2_U5610;
  assign new_P2_U3874 = new_P2_U5612 & new_P2_U5613;
  assign new_P2_U3875 = new_P2_U5615 & new_P2_U5616;
  assign new_P2_U3876 = new_P2_U5618 & new_P2_U5619;
  assign new_P2_U3877 = new_P2_U5621 & new_P2_U5622;
  assign new_P2_U3878 = new_P2_U5624 & new_P2_U5625;
  assign new_P2_U3879 = ~P2_IR_REG_31_;
  assign new_P2_U3880 = ~new_P2_U3023 | ~new_P2_U3333;
  assign new_P2_U3881 = ~new_P2_U3577 | ~new_P2_U3050;
  assign new_P2_U3882 = ~new_P2_U3695 | ~new_P2_U3050;
  assign new_P2_U3883 = new_P2_U5922 & new_P2_U5921;
  assign new_P2_U3884 = new_P2_U5924 & new_P2_U5923;
  assign new_P2_U3885 = new_P2_U5926 & new_P2_U5925;
  assign new_P2_U3886 = new_P2_U5928 & new_P2_U5927;
  assign new_P2_U3887 = new_P2_U5930 & new_P2_U5929;
  assign new_P2_U3888 = new_P2_U5932 & new_P2_U5931;
  assign new_P2_U3889 = new_P2_U5934 & new_P2_U5933;
  assign new_P2_U3890 = new_P2_U5936 & new_P2_U5935;
  assign new_P2_U3891 = new_P2_U5938 & new_P2_U5937;
  assign new_P2_U3892 = new_P2_U5940 & new_P2_U5939;
  assign new_P2_U3893 = new_P2_U5942 & new_P2_U5941;
  assign new_P2_U3894 = new_P2_U5944 & new_P2_U5943;
  assign new_P2_U3895 = new_P2_U5946 & new_P2_U5945;
  assign new_P2_U3896 = new_P2_U5948 & new_P2_U5947;
  assign new_P2_U3897 = new_P2_U5950 & new_P2_U5949;
  assign new_P2_U3898 = new_P2_U5952 & new_P2_U5951;
  assign new_P2_U3899 = new_P2_U5954 & new_P2_U5953;
  assign new_P2_U3900 = new_P2_U5956 & new_P2_U5955;
  assign new_P2_U3901 = new_P2_U5958 & new_P2_U5957;
  assign new_P2_U3902 = new_P2_U5960 & new_P2_U5959;
  assign new_P2_U3903 = new_P2_U5962 & new_P2_U5961;
  assign new_P2_U3904 = new_P2_U5964 & new_P2_U5963;
  assign new_P2_U3905 = new_P2_U5966 & new_P2_U5965;
  assign new_P2_U3906 = new_P2_U5968 & new_P2_U5967;
  assign new_P2_U3907 = new_P2_U5970 & new_P2_U5969;
  assign new_P2_U3908 = new_P2_U5972 & new_P2_U5971;
  assign new_P2_U3909 = new_P2_U5974 & new_P2_U5973;
  assign new_P2_U3910 = new_P2_U5976 & new_P2_U5975;
  assign new_P2_U3911 = new_P2_U5978 & new_P2_U5977;
  assign new_P2_U3912 = new_P2_U5980 & new_P2_U5979;
  assign new_P2_U3913 = ~new_P2_U3694 | ~new_P2_U3058;
  assign new_P2_U3914 = new_P2_U5982 & new_P2_U5981;
  assign new_P2_U3915 = new_P2_U5984 & new_P2_U5983;
  assign new_P2_U3916 = ~new_P2_R1312_U18;
  assign new_P2_U3917 = new_P2_U6050 & new_P2_U6049;
  assign new_P2_U3918 = ~new_P2_U3793 | ~new_P2_U6082 | ~new_P2_U6085 | ~new_P2_U3794 | ~new_P2_U3792;
  assign new_P2_U3919 = ~new_P2_U3049 | ~new_P2_U5674;
  assign new_P2_U3920 = ~new_P2_U3973 | ~new_P2_U3418;
  assign new_P2_U3921 = ~new_P2_U3390;
  assign new_P2_U3922 = ~new_P2_U3342;
  assign new_P2_U3923 = ~new_P2_U3976 | ~new_P2_U3418;
  assign new_P2_U3924 = ~new_P2_U3339;
  assign new_P2_U3925 = ~new_P2_U3346;
  assign new_P2_U3926 = ~new_P2_U3336;
  assign new_P2_U3927 = ~new_P2_U3394;
  assign new_P2_U3928 = ~new_P2_U3973 | ~new_P2_U3420;
  assign new_P2_U3929 = ~new_P2_U3410;
  assign new_P2_U3930 = ~new_P2_U3335;
  assign new_P2_U3931 = ~new_P2_U3334;
  assign new_P2_U3932 = ~new_P2_U3395;
  assign new_P2_U3933 = ~new_P2_U3393;
  assign new_P2_U3934 = ~new_P2_U3925 | ~new_P2_U5674;
  assign new_P2_U3935 = ~new_P2_U3963 | ~new_P2_U3340;
  assign new_P2_U3936 = ~new_P2_U3973 | ~new_P2_U5671;
  assign new_P2_U3937 = ~new_P2_U3402;
  assign new_P2_U3938 = ~new_P2_U3392;
  assign new_P2_U3939 = ~new_P2_U3341;
  assign new_P2_U3940 = ~new_P2_U3919;
  assign new_P2_U3941 = ~new_P2_U3337;
  assign new_P2_U3942 = ~new_P2_U3920;
  assign new_P2_U3943 = ~new_P2_U3338;
  assign new_P2_U3944 = ~new_P2_U3343;
  assign new_P2_U3945 = ~new_P2_U3347;
  assign new_P2_U3946 = ~new_P2_U3406;
  assign n2619 = ~new_P2_U3400;
  assign new_P2_U3948 = ~new_P2_U3397;
  assign new_P2_U3949 = ~new_P2_U3384;
  assign new_P2_U3950 = ~new_P2_U3382;
  assign new_P2_U3951 = ~new_P2_U3380;
  assign new_P2_U3952 = ~new_P2_U3378;
  assign new_P2_U3953 = ~new_P2_U3376;
  assign new_P2_U3954 = ~new_P2_U3374;
  assign new_P2_U3955 = ~new_P2_U3372;
  assign new_P2_U3956 = ~new_P2_U3370;
  assign new_P2_U3957 = ~new_P2_U3368;
  assign new_P2_U3958 = ~new_P2_U3389;
  assign new_P2_U3959 = ~new_P2_U3388;
  assign new_P2_U3960 = ~new_P2_U3386;
  assign new_P2_U3961 = ~new_P2_U3403;
  assign new_P2_U3962 = ~new_P2_U3396;
  assign new_P2_U3963 = ~new_P2_U3344;
  assign new_P2_U3964 = ~new_P2_U3391;
  assign new_P2_U3965 = ~new_P2_U3882;
  assign new_P2_U3966 = ~new_P2_U3881;
  assign new_P2_U3967 = ~new_P2_U3880;
  assign new_P2_U3968 = ~new_P2_U3913;
  assign new_P2_U3969 = ~new_P2_U3407;
  assign new_P2_U3970 = ~new_P2_U3408 | ~P2_STATE_REG;
  assign new_P2_U3971 = ~new_P2_U3933 | ~new_P2_U3023;
  assign new_P2_U3972 = ~new_P2_U3405;
  assign new_P2_U3973 = ~new_P2_U3404;
  assign new_P2_U3974 = ~new_P2_U3340;
  assign new_P2_U3975 = ~new_P2_U3332;
  assign new_P2_U3976 = ~new_P2_U3345;
  assign new_P2_U3977 = ~new_P2_U3399;
  assign new_P2_U3978 = ~new_P2_U3329;
  assign new_P2_U3979 = ~new_U93 | ~n2609;
  assign new_P2_U3980 = ~P2_IR_REG_0_ | ~new_P2_U3030;
  assign new_P2_U3981 = ~P2_IR_REG_0_ | ~new_P2_U3978;
  assign new_P2_U3982 = ~new_U82 | ~n2609;
  assign new_P2_U3983 = ~new_P2_SUB_1108_U42 | ~new_P2_U3030;
  assign new_P2_U3984 = ~P2_IR_REG_1_ | ~new_P2_U3978;
  assign new_P2_U3985 = ~new_U71 | ~n2609;
  assign new_P2_U3986 = ~new_P2_SUB_1108_U17 | ~new_P2_U3030;
  assign new_P2_U3987 = ~P2_IR_REG_2_ | ~new_P2_U3978;
  assign new_P2_U3988 = ~new_U68 | ~n2609;
  assign new_P2_U3989 = ~new_P2_SUB_1108_U18 | ~new_P2_U3030;
  assign new_P2_U3990 = ~P2_IR_REG_3_ | ~new_P2_U3978;
  assign new_P2_U3991 = ~new_U67 | ~n2609;
  assign new_P2_U3992 = ~new_P2_SUB_1108_U19 | ~new_P2_U3030;
  assign new_P2_U3993 = ~P2_IR_REG_4_ | ~new_P2_U3978;
  assign new_P2_U3994 = ~new_U66 | ~n2609;
  assign new_P2_U3995 = ~new_P2_SUB_1108_U101 | ~new_P2_U3030;
  assign new_P2_U3996 = ~P2_IR_REG_5_ | ~new_P2_U3978;
  assign new_P2_U3997 = ~new_U65 | ~n2609;
  assign new_P2_U3998 = ~new_P2_SUB_1108_U20 | ~new_P2_U3030;
  assign new_P2_U3999 = ~P2_IR_REG_6_ | ~new_P2_U3978;
  assign new_P2_U4000 = ~new_U64 | ~n2609;
  assign new_P2_U4001 = ~new_P2_SUB_1108_U21 | ~new_P2_U3030;
  assign new_P2_U4002 = ~P2_IR_REG_7_ | ~new_P2_U3978;
  assign new_P2_U4003 = ~new_U63 | ~n2609;
  assign new_P2_U4004 = ~new_P2_SUB_1108_U22 | ~new_P2_U3030;
  assign new_P2_U4005 = ~P2_IR_REG_8_ | ~new_P2_U3978;
  assign new_P2_U4006 = ~new_U62 | ~n2609;
  assign new_P2_U4007 = ~new_P2_SUB_1108_U99 | ~new_P2_U3030;
  assign new_P2_U4008 = ~P2_IR_REG_9_ | ~new_P2_U3978;
  assign new_P2_U4009 = ~new_U92 | ~n2609;
  assign new_P2_U4010 = ~new_P2_SUB_1108_U6 | ~new_P2_U3030;
  assign new_P2_U4011 = ~P2_IR_REG_10_ | ~new_P2_U3978;
  assign new_P2_U4012 = ~new_U91 | ~n2609;
  assign new_P2_U4013 = ~new_P2_SUB_1108_U7 | ~new_P2_U3030;
  assign new_P2_U4014 = ~P2_IR_REG_11_ | ~new_P2_U3978;
  assign new_P2_U4015 = ~new_U90 | ~n2609;
  assign new_P2_U4016 = ~new_P2_SUB_1108_U8 | ~new_P2_U3030;
  assign new_P2_U4017 = ~P2_IR_REG_12_ | ~new_P2_U3978;
  assign new_P2_U4018 = ~new_U89 | ~n2609;
  assign new_P2_U4019 = ~new_P2_SUB_1108_U127 | ~new_P2_U3030;
  assign new_P2_U4020 = ~P2_IR_REG_13_ | ~new_P2_U3978;
  assign new_P2_U4021 = ~new_U88 | ~n2609;
  assign new_P2_U4022 = ~new_P2_SUB_1108_U9 | ~new_P2_U3030;
  assign new_P2_U4023 = ~P2_IR_REG_14_ | ~new_P2_U3978;
  assign new_P2_U4024 = ~new_U87 | ~n2609;
  assign new_P2_U4025 = ~new_P2_SUB_1108_U10 | ~new_P2_U3030;
  assign new_P2_U4026 = ~P2_IR_REG_15_ | ~new_P2_U3978;
  assign new_P2_U4027 = ~new_U86 | ~n2609;
  assign new_P2_U4028 = ~new_P2_SUB_1108_U11 | ~new_P2_U3030;
  assign new_P2_U4029 = ~P2_IR_REG_16_ | ~new_P2_U3978;
  assign new_P2_U4030 = ~new_U85 | ~n2609;
  assign new_P2_U4031 = ~new_P2_SUB_1108_U125 | ~new_P2_U3030;
  assign new_P2_U4032 = ~P2_IR_REG_17_ | ~new_P2_U3978;
  assign new_P2_U4033 = ~new_U84 | ~n2609;
  assign new_P2_U4034 = ~new_P2_SUB_1108_U12 | ~new_P2_U3030;
  assign new_P2_U4035 = ~P2_IR_REG_18_ | ~new_P2_U3978;
  assign new_P2_U4036 = ~new_U83 | ~n2609;
  assign new_P2_U4037 = ~new_P2_SUB_1108_U123 | ~new_P2_U3030;
  assign new_P2_U4038 = ~P2_IR_REG_19_ | ~new_P2_U3978;
  assign new_P2_U4039 = ~new_U81 | ~n2609;
  assign new_P2_U4040 = ~new_P2_SUB_1108_U119 | ~new_P2_U3030;
  assign new_P2_U4041 = ~P2_IR_REG_20_ | ~new_P2_U3978;
  assign new_P2_U4042 = ~new_U80 | ~n2609;
  assign new_P2_U4043 = ~new_P2_SUB_1108_U116 | ~new_P2_U3030;
  assign new_P2_U4044 = ~P2_IR_REG_21_ | ~new_P2_U3978;
  assign new_P2_U4045 = ~new_U79 | ~n2609;
  assign new_P2_U4046 = ~new_P2_SUB_1108_U114 | ~new_P2_U3030;
  assign new_P2_U4047 = ~P2_IR_REG_22_ | ~new_P2_U3978;
  assign new_P2_U4048 = ~new_U78 | ~n2609;
  assign new_P2_U4049 = ~new_P2_SUB_1108_U13 | ~new_P2_U3030;
  assign new_P2_U4050 = ~P2_IR_REG_23_ | ~new_P2_U3978;
  assign new_P2_U4051 = ~new_U77 | ~n2609;
  assign new_P2_U4052 = ~new_P2_SUB_1108_U14 | ~new_P2_U3030;
  assign new_P2_U4053 = ~P2_IR_REG_24_ | ~new_P2_U3978;
  assign new_P2_U4054 = ~new_U76 | ~n2609;
  assign new_P2_U4055 = ~new_P2_SUB_1108_U112 | ~new_P2_U3030;
  assign new_P2_U4056 = ~P2_IR_REG_25_ | ~new_P2_U3978;
  assign new_P2_U4057 = ~new_U75 | ~n2609;
  assign new_P2_U4058 = ~new_P2_SUB_1108_U15 | ~new_P2_U3030;
  assign new_P2_U4059 = ~P2_IR_REG_26_ | ~new_P2_U3978;
  assign new_P2_U4060 = ~new_U74 | ~n2609;
  assign new_P2_U4061 = ~new_P2_SUB_1108_U110 | ~new_P2_U3030;
  assign new_P2_U4062 = ~P2_IR_REG_27_ | ~new_P2_U3978;
  assign new_P2_U4063 = ~new_U73 | ~n2609;
  assign new_P2_U4064 = ~new_P2_SUB_1108_U107 | ~new_P2_U3030;
  assign new_P2_U4065 = ~P2_IR_REG_28_ | ~new_P2_U3978;
  assign new_P2_U4066 = ~new_U72 | ~n2609;
  assign new_P2_U4067 = ~new_P2_SUB_1108_U16 | ~new_P2_U3030;
  assign new_P2_U4068 = ~P2_IR_REG_29_ | ~new_P2_U3978;
  assign new_P2_U4069 = ~new_U70 | ~n2609;
  assign new_P2_U4070 = ~new_P2_SUB_1108_U104 | ~new_P2_U3030;
  assign new_P2_U4071 = ~P2_IR_REG_30_ | ~new_P2_U3978;
  assign new_P2_U4072 = ~new_U69 | ~n2609;
  assign new_P2_U4073 = ~new_P2_SUB_1108_U43 | ~new_P2_U3030;
  assign new_P2_U4074 = ~P2_IR_REG_31_ | ~new_P2_U3978;
  assign new_P2_U4075 = ~new_P2_U3975 | ~new_P2_U5655;
  assign new_P2_U4076 = ~new_P2_U3333;
  assign new_P2_U4077 = ~new_P2_U3332 | ~new_P2_U5646;
  assign new_P2_U4078 = ~new_P2_U3332 | ~new_P2_U5649;
  assign new_P2_U4079 = ~new_P2_U4076 | ~P2_D_REG_10_;
  assign new_P2_U4080 = ~new_P2_U4076 | ~P2_D_REG_11_;
  assign new_P2_U4081 = ~new_P2_U4076 | ~P2_D_REG_12_;
  assign new_P2_U4082 = ~new_P2_U4076 | ~P2_D_REG_13_;
  assign new_P2_U4083 = ~new_P2_U4076 | ~P2_D_REG_14_;
  assign new_P2_U4084 = ~new_P2_U4076 | ~P2_D_REG_15_;
  assign new_P2_U4085 = ~new_P2_U4076 | ~P2_D_REG_16_;
  assign new_P2_U4086 = ~new_P2_U4076 | ~P2_D_REG_17_;
  assign new_P2_U4087 = ~new_P2_U4076 | ~P2_D_REG_18_;
  assign new_P2_U4088 = ~new_P2_U4076 | ~P2_D_REG_19_;
  assign new_P2_U4089 = ~new_P2_U4076 | ~P2_D_REG_20_;
  assign new_P2_U4090 = ~new_P2_U4076 | ~P2_D_REG_21_;
  assign new_P2_U4091 = ~new_P2_U4076 | ~P2_D_REG_22_;
  assign new_P2_U4092 = ~new_P2_U4076 | ~P2_D_REG_23_;
  assign new_P2_U4093 = ~new_P2_U4076 | ~P2_D_REG_24_;
  assign new_P2_U4094 = ~new_P2_U4076 | ~P2_D_REG_25_;
  assign new_P2_U4095 = ~new_P2_U4076 | ~P2_D_REG_26_;
  assign new_P2_U4096 = ~new_P2_U4076 | ~P2_D_REG_27_;
  assign new_P2_U4097 = ~new_P2_U4076 | ~P2_D_REG_28_;
  assign new_P2_U4098 = ~new_P2_U4076 | ~P2_D_REG_29_;
  assign new_P2_U4099 = ~new_P2_U4076 | ~P2_D_REG_2_;
  assign new_P2_U4100 = ~new_P2_U4076 | ~P2_D_REG_30_;
  assign new_P2_U4101 = ~new_P2_U4076 | ~P2_D_REG_31_;
  assign new_P2_U4102 = ~new_P2_U4076 | ~P2_D_REG_3_;
  assign new_P2_U4103 = ~new_P2_U4076 | ~P2_D_REG_4_;
  assign new_P2_U4104 = ~new_P2_U4076 | ~P2_D_REG_5_;
  assign new_P2_U4105 = ~new_P2_U4076 | ~P2_D_REG_6_;
  assign new_P2_U4106 = ~new_P2_U4076 | ~P2_D_REG_7_;
  assign new_P2_U4107 = ~new_P2_U4076 | ~P2_D_REG_8_;
  assign new_P2_U4108 = ~new_P2_U4076 | ~P2_D_REG_9_;
  assign new_P2_U4109 = ~new_P2_U5674 | ~new_P2_U5671;
  assign new_P2_U4110 = ~new_P2_U3340 | ~new_P2_U5693 | ~new_P2_U5692;
  assign new_P2_U4111 = ~new_P2_U3020 | ~P2_REG2_REG_1_;
  assign new_P2_U4112 = ~new_P2_U3021 | ~P2_REG1_REG_1_;
  assign new_P2_U4113 = ~new_P2_U3022 | ~P2_REG0_REG_1_;
  assign new_P2_U4114 = ~P2_REG3_REG_1_ | ~new_P2_U3019;
  assign new_P2_U4115 = ~new_P2_U3080;
  assign new_P2_U4116 = ~new_P2_U3390 | ~new_P2_U3934;
  assign new_P2_U4117 = ~new_P2_U3931 | ~new_P2_R1146_U20;
  assign new_P2_U4118 = ~new_P2_U3930 | ~new_P2_R1113_U20;
  assign new_P2_U4119 = ~new_P2_U3926 | ~new_P2_R1131_U95;
  assign new_P2_U4120 = ~new_P2_U3941 | ~new_P2_R1179_U20;
  assign new_P2_U4121 = ~new_P2_U3943 | ~new_P2_R1203_U20;
  assign new_P2_U4122 = ~new_P2_U3014 | ~new_P2_R1164_U95;
  assign new_P2_U4123 = ~new_P2_U3922 | ~new_P2_R1233_U95;
  assign new_P2_U4124 = ~new_P2_U3348;
  assign new_P2_U4125 = ~new_P2_U3427 | ~new_P2_U3027;
  assign new_P2_U4126 = ~new_P2_U3026 | ~new_P2_U3080;
  assign new_P2_U4127 = ~new_P2_R1215_U96 | ~new_P2_U3025;
  assign new_P2_U4128 = ~new_P2_U3427 | ~new_P2_U4116;
  assign new_P2_U4129 = ~new_P2_U4124 | ~new_P2_U3565 | ~new_P2_U4128 | ~new_P2_U4126;
  assign new_P2_U4130 = ~P2_REG2_REG_2_ | ~new_P2_U3020;
  assign new_P2_U4131 = ~P2_REG1_REG_2_ | ~new_P2_U3021;
  assign new_P2_U4132 = ~P2_REG0_REG_2_ | ~new_P2_U3022;
  assign new_P2_U4133 = ~P2_REG3_REG_2_ | ~new_P2_U3019;
  assign new_P2_U4134 = ~new_P2_U3070;
  assign new_P2_U4135 = ~P2_REG2_REG_0_ | ~new_P2_U3020;
  assign new_P2_U4136 = ~P2_REG1_REG_0_ | ~new_P2_U3021;
  assign new_P2_U4137 = ~P2_REG0_REG_0_ | ~new_P2_U3022;
  assign new_P2_U4138 = ~P2_REG3_REG_0_ | ~new_P2_U3019;
  assign new_P2_U4139 = ~new_P2_U3079;
  assign new_P2_U4140 = ~new_P2_U3035 | ~new_P2_U3079;
  assign new_P2_U4141 = ~new_P2_R1146_U97 | ~new_P2_U3931;
  assign new_P2_U4142 = ~new_P2_R1113_U97 | ~new_P2_U3930;
  assign new_P2_U4143 = ~new_P2_R1131_U94 | ~new_P2_U3926;
  assign new_P2_U4144 = ~new_P2_R1179_U97 | ~new_P2_U3941;
  assign new_P2_U4145 = ~new_P2_R1203_U97 | ~new_P2_U3943;
  assign new_P2_U4146 = ~new_P2_R1164_U94 | ~new_P2_U3014;
  assign new_P2_U4147 = ~new_P2_R1233_U94 | ~new_P2_U3922;
  assign new_P2_U4148 = ~new_P2_U3349;
  assign new_P2_U4149 = ~new_P2_R1275_U55 | ~new_P2_U3027;
  assign new_P2_U4150 = ~new_P2_U3026 | ~new_P2_U3070;
  assign new_P2_U4151 = ~new_P2_R1215_U95 | ~new_P2_U3025;
  assign new_P2_U4152 = ~new_P2_U3432 | ~new_P2_U4116;
  assign new_P2_U4153 = ~new_P2_U3581 | ~new_P2_U4148;
  assign new_P2_U4154 = ~P2_REG2_REG_3_ | ~new_P2_U3020;
  assign new_P2_U4155 = ~P2_REG1_REG_3_ | ~new_P2_U3021;
  assign new_P2_U4156 = ~P2_REG0_REG_3_ | ~new_P2_U3022;
  assign new_P2_U4157 = ~new_P2_ADD_1119_U4 | ~new_P2_U3019;
  assign new_P2_U4158 = ~new_P2_U3066;
  assign new_P2_U4159 = ~new_P2_U3035 | ~new_P2_U3080;
  assign new_P2_U4160 = ~new_P2_R1146_U107 | ~new_P2_U3931;
  assign new_P2_U4161 = ~new_P2_R1113_U107 | ~new_P2_U3930;
  assign new_P2_U4162 = ~new_P2_R1131_U16 | ~new_P2_U3926;
  assign new_P2_U4163 = ~new_P2_R1179_U107 | ~new_P2_U3941;
  assign new_P2_U4164 = ~new_P2_R1203_U107 | ~new_P2_U3943;
  assign new_P2_U4165 = ~new_P2_R1164_U16 | ~new_P2_U3014;
  assign new_P2_U4166 = ~new_P2_R1233_U16 | ~new_P2_U3922;
  assign new_P2_U4167 = ~new_P2_U3350;
  assign new_P2_U4168 = ~new_P2_R1275_U18 | ~new_P2_U3027;
  assign new_P2_U4169 = ~new_P2_U3026 | ~new_P2_U3066;
  assign new_P2_U4170 = ~new_P2_R1215_U17 | ~new_P2_U3025;
  assign new_P2_U4171 = ~new_P2_U3435 | ~new_P2_U4116;
  assign new_P2_U4172 = ~new_P2_U3585 | ~new_P2_U4167;
  assign new_P2_U4173 = ~P2_REG2_REG_4_ | ~new_P2_U3020;
  assign new_P2_U4174 = ~P2_REG1_REG_4_ | ~new_P2_U3021;
  assign new_P2_U4175 = ~P2_REG0_REG_4_ | ~new_P2_U3022;
  assign new_P2_U4176 = ~new_P2_ADD_1119_U55 | ~new_P2_U3019;
  assign new_P2_U4177 = ~new_P2_U3062;
  assign new_P2_U4178 = ~new_P2_U3035 | ~new_P2_U3070;
  assign new_P2_U4179 = ~new_P2_R1146_U17 | ~new_P2_U3931;
  assign new_P2_U4180 = ~new_P2_R1113_U17 | ~new_P2_U3930;
  assign new_P2_U4181 = ~new_P2_R1131_U100 | ~new_P2_U3926;
  assign new_P2_U4182 = ~new_P2_R1179_U17 | ~new_P2_U3941;
  assign new_P2_U4183 = ~new_P2_R1203_U17 | ~new_P2_U3943;
  assign new_P2_U4184 = ~new_P2_R1164_U100 | ~new_P2_U3014;
  assign new_P2_U4185 = ~new_P2_R1233_U100 | ~new_P2_U3922;
  assign new_P2_U4186 = ~new_P2_U3351;
  assign new_P2_U4187 = ~new_P2_R1275_U20 | ~new_P2_U3027;
  assign new_P2_U4188 = ~new_P2_U3026 | ~new_P2_U3062;
  assign new_P2_U4189 = ~new_P2_R1215_U101 | ~new_P2_U3025;
  assign new_P2_U4190 = ~new_P2_U3438 | ~new_P2_U4116;
  assign new_P2_U4191 = ~new_P2_U3589 | ~new_P2_U4186;
  assign new_P2_U4192 = ~P2_REG2_REG_5_ | ~new_P2_U3020;
  assign new_P2_U4193 = ~P2_REG1_REG_5_ | ~new_P2_U3021;
  assign new_P2_U4194 = ~P2_REG0_REG_5_ | ~new_P2_U3022;
  assign new_P2_U4195 = ~new_P2_ADD_1119_U54 | ~new_P2_U3019;
  assign new_P2_U4196 = ~new_P2_U3069;
  assign new_P2_U4197 = ~new_P2_U3035 | ~new_P2_U3066;
  assign new_P2_U4198 = ~new_P2_R1146_U106 | ~new_P2_U3931;
  assign new_P2_U4199 = ~new_P2_R1113_U106 | ~new_P2_U3930;
  assign new_P2_U4200 = ~new_P2_R1131_U99 | ~new_P2_U3926;
  assign new_P2_U4201 = ~new_P2_R1179_U106 | ~new_P2_U3941;
  assign new_P2_U4202 = ~new_P2_R1203_U106 | ~new_P2_U3943;
  assign new_P2_U4203 = ~new_P2_R1164_U99 | ~new_P2_U3014;
  assign new_P2_U4204 = ~new_P2_R1233_U99 | ~new_P2_U3922;
  assign new_P2_U4205 = ~new_P2_U3352;
  assign new_P2_U4206 = ~new_P2_R1275_U21 | ~new_P2_U3027;
  assign new_P2_U4207 = ~new_P2_U3026 | ~new_P2_U3069;
  assign new_P2_U4208 = ~new_P2_R1215_U100 | ~new_P2_U3025;
  assign new_P2_U4209 = ~new_P2_U3441 | ~new_P2_U4116;
  assign new_P2_U4210 = ~new_P2_U3593 | ~new_P2_U4205;
  assign new_P2_U4211 = ~P2_REG2_REG_6_ | ~new_P2_U3020;
  assign new_P2_U4212 = ~P2_REG1_REG_6_ | ~new_P2_U3021;
  assign new_P2_U4213 = ~P2_REG0_REG_6_ | ~new_P2_U3022;
  assign new_P2_U4214 = ~new_P2_ADD_1119_U53 | ~new_P2_U3019;
  assign new_P2_U4215 = ~new_P2_U3073;
  assign new_P2_U4216 = ~new_P2_U3035 | ~new_P2_U3062;
  assign new_P2_U4217 = ~new_P2_R1146_U105 | ~new_P2_U3931;
  assign new_P2_U4218 = ~new_P2_R1113_U105 | ~new_P2_U3930;
  assign new_P2_U4219 = ~new_P2_R1131_U17 | ~new_P2_U3926;
  assign new_P2_U4220 = ~new_P2_R1179_U105 | ~new_P2_U3941;
  assign new_P2_U4221 = ~new_P2_R1203_U105 | ~new_P2_U3943;
  assign new_P2_U4222 = ~new_P2_R1164_U17 | ~new_P2_U3014;
  assign new_P2_U4223 = ~new_P2_R1233_U17 | ~new_P2_U3922;
  assign new_P2_U4224 = ~new_P2_U3353;
  assign new_P2_U4225 = ~new_P2_R1275_U65 | ~new_P2_U3027;
  assign new_P2_U4226 = ~new_P2_U3026 | ~new_P2_U3073;
  assign new_P2_U4227 = ~new_P2_R1215_U18 | ~new_P2_U3025;
  assign new_P2_U4228 = ~new_P2_U3444 | ~new_P2_U4116;
  assign new_P2_U4229 = ~new_P2_U3597 | ~new_P2_U4224;
  assign new_P2_U4230 = ~P2_REG2_REG_7_ | ~new_P2_U3020;
  assign new_P2_U4231 = ~P2_REG1_REG_7_ | ~new_P2_U3021;
  assign new_P2_U4232 = ~P2_REG0_REG_7_ | ~new_P2_U3022;
  assign new_P2_U4233 = ~new_P2_ADD_1119_U52 | ~new_P2_U3019;
  assign new_P2_U4234 = ~new_P2_U3072;
  assign new_P2_U4235 = ~new_P2_U3035 | ~new_P2_U3069;
  assign new_P2_U4236 = ~new_P2_R1146_U18 | ~new_P2_U3931;
  assign new_P2_U4237 = ~new_P2_R1113_U18 | ~new_P2_U3930;
  assign new_P2_U4238 = ~new_P2_R1131_U98 | ~new_P2_U3926;
  assign new_P2_U4239 = ~new_P2_R1179_U18 | ~new_P2_U3941;
  assign new_P2_U4240 = ~new_P2_R1203_U18 | ~new_P2_U3943;
  assign new_P2_U4241 = ~new_P2_R1164_U98 | ~new_P2_U3014;
  assign new_P2_U4242 = ~new_P2_R1233_U98 | ~new_P2_U3922;
  assign new_P2_U4243 = ~new_P2_U3354;
  assign new_P2_U4244 = ~new_P2_R1275_U22 | ~new_P2_U3027;
  assign new_P2_U4245 = ~new_P2_U3026 | ~new_P2_U3072;
  assign new_P2_U4246 = ~new_P2_R1215_U99 | ~new_P2_U3025;
  assign new_P2_U4247 = ~new_P2_U3447 | ~new_P2_U4116;
  assign new_P2_U4248 = ~new_P2_U3601 | ~new_P2_U4243;
  assign new_P2_U4249 = ~P2_REG2_REG_8_ | ~new_P2_U3020;
  assign new_P2_U4250 = ~P2_REG1_REG_8_ | ~new_P2_U3021;
  assign new_P2_U4251 = ~P2_REG0_REG_8_ | ~new_P2_U3022;
  assign new_P2_U4252 = ~new_P2_ADD_1119_U51 | ~new_P2_U3019;
  assign new_P2_U4253 = ~new_P2_U3086;
  assign new_P2_U4254 = ~new_P2_U3035 | ~new_P2_U3073;
  assign new_P2_U4255 = ~new_P2_R1146_U104 | ~new_P2_U3931;
  assign new_P2_U4256 = ~new_P2_R1113_U104 | ~new_P2_U3930;
  assign new_P2_U4257 = ~new_P2_R1131_U18 | ~new_P2_U3926;
  assign new_P2_U4258 = ~new_P2_R1179_U104 | ~new_P2_U3941;
  assign new_P2_U4259 = ~new_P2_R1203_U104 | ~new_P2_U3943;
  assign new_P2_U4260 = ~new_P2_R1164_U18 | ~new_P2_U3014;
  assign new_P2_U4261 = ~new_P2_R1233_U18 | ~new_P2_U3922;
  assign new_P2_U4262 = ~new_P2_U3355;
  assign new_P2_U4263 = ~new_P2_R1275_U23 | ~new_P2_U3027;
  assign new_P2_U4264 = ~new_P2_U3026 | ~new_P2_U3086;
  assign new_P2_U4265 = ~new_P2_R1215_U19 | ~new_P2_U3025;
  assign new_P2_U4266 = ~new_P2_U3450 | ~new_P2_U4116;
  assign new_P2_U4267 = ~new_P2_U3605 | ~new_P2_U4262;
  assign new_P2_U4268 = ~P2_REG2_REG_9_ | ~new_P2_U3020;
  assign new_P2_U4269 = ~P2_REG1_REG_9_ | ~new_P2_U3021;
  assign new_P2_U4270 = ~P2_REG0_REG_9_ | ~new_P2_U3022;
  assign new_P2_U4271 = ~new_P2_ADD_1119_U50 | ~new_P2_U3019;
  assign new_P2_U4272 = ~new_P2_U3085;
  assign new_P2_U4273 = ~new_P2_U3035 | ~new_P2_U3072;
  assign new_P2_U4274 = ~new_P2_R1146_U19 | ~new_P2_U3931;
  assign new_P2_U4275 = ~new_P2_R1113_U19 | ~new_P2_U3930;
  assign new_P2_U4276 = ~new_P2_R1131_U97 | ~new_P2_U3926;
  assign new_P2_U4277 = ~new_P2_R1179_U19 | ~new_P2_U3941;
  assign new_P2_U4278 = ~new_P2_R1203_U19 | ~new_P2_U3943;
  assign new_P2_U4279 = ~new_P2_R1164_U97 | ~new_P2_U3014;
  assign new_P2_U4280 = ~new_P2_R1233_U97 | ~new_P2_U3922;
  assign new_P2_U4281 = ~new_P2_U3356;
  assign new_P2_U4282 = ~new_P2_R1275_U24 | ~new_P2_U3027;
  assign new_P2_U4283 = ~new_P2_U3026 | ~new_P2_U3085;
  assign new_P2_U4284 = ~new_P2_R1215_U98 | ~new_P2_U3025;
  assign new_P2_U4285 = ~new_P2_U3453 | ~new_P2_U4116;
  assign new_P2_U4286 = ~new_P2_U3609 | ~new_P2_U4281;
  assign new_P2_U4287 = ~P2_REG2_REG_10_ | ~new_P2_U3020;
  assign new_P2_U4288 = ~P2_REG1_REG_10_ | ~new_P2_U3021;
  assign new_P2_U4289 = ~P2_REG0_REG_10_ | ~new_P2_U3022;
  assign new_P2_U4290 = ~new_P2_ADD_1119_U74 | ~new_P2_U3019;
  assign new_P2_U4291 = ~new_P2_U3064;
  assign new_P2_U4292 = ~new_P2_U3035 | ~new_P2_U3086;
  assign new_P2_U4293 = ~new_P2_R1146_U103 | ~new_P2_U3931;
  assign new_P2_U4294 = ~new_P2_R1113_U103 | ~new_P2_U3930;
  assign new_P2_U4295 = ~new_P2_R1131_U96 | ~new_P2_U3926;
  assign new_P2_U4296 = ~new_P2_R1179_U103 | ~new_P2_U3941;
  assign new_P2_U4297 = ~new_P2_R1203_U103 | ~new_P2_U3943;
  assign new_P2_U4298 = ~new_P2_R1164_U96 | ~new_P2_U3014;
  assign new_P2_U4299 = ~new_P2_R1233_U96 | ~new_P2_U3922;
  assign new_P2_U4300 = ~new_P2_U3357;
  assign new_P2_U4301 = ~new_P2_R1275_U63 | ~new_P2_U3027;
  assign new_P2_U4302 = ~new_P2_U3026 | ~new_P2_U3064;
  assign new_P2_U4303 = ~new_P2_R1215_U97 | ~new_P2_U3025;
  assign new_P2_U4304 = ~new_P2_U3456 | ~new_P2_U4116;
  assign new_P2_U4305 = ~new_P2_U3613 | ~new_P2_U4300;
  assign new_P2_U4306 = ~P2_REG2_REG_11_ | ~new_P2_U3020;
  assign new_P2_U4307 = ~P2_REG1_REG_11_ | ~new_P2_U3021;
  assign new_P2_U4308 = ~P2_REG0_REG_11_ | ~new_P2_U3022;
  assign new_P2_U4309 = ~new_P2_ADD_1119_U73 | ~new_P2_U3019;
  assign new_P2_U4310 = ~new_P2_U3065;
  assign new_P2_U4311 = ~new_P2_U3035 | ~new_P2_U3085;
  assign new_P2_U4312 = ~new_P2_R1146_U113 | ~new_P2_U3931;
  assign new_P2_U4313 = ~new_P2_R1113_U113 | ~new_P2_U3930;
  assign new_P2_U4314 = ~new_P2_R1131_U10 | ~new_P2_U3926;
  assign new_P2_U4315 = ~new_P2_R1179_U113 | ~new_P2_U3941;
  assign new_P2_U4316 = ~new_P2_R1203_U113 | ~new_P2_U3943;
  assign new_P2_U4317 = ~new_P2_R1164_U10 | ~new_P2_U3014;
  assign new_P2_U4318 = ~new_P2_R1233_U10 | ~new_P2_U3922;
  assign new_P2_U4319 = ~new_P2_U3358;
  assign new_P2_U4320 = ~new_P2_R1275_U6 | ~new_P2_U3027;
  assign new_P2_U4321 = ~new_P2_U3026 | ~new_P2_U3065;
  assign new_P2_U4322 = ~new_P2_R1215_U11 | ~new_P2_U3025;
  assign new_P2_U4323 = ~new_P2_U3459 | ~new_P2_U4116;
  assign new_P2_U4324 = ~new_P2_U3617 | ~new_P2_U4319;
  assign new_P2_U4325 = ~P2_REG2_REG_12_ | ~new_P2_U3020;
  assign new_P2_U4326 = ~P2_REG1_REG_12_ | ~new_P2_U3021;
  assign new_P2_U4327 = ~P2_REG0_REG_12_ | ~new_P2_U3022;
  assign new_P2_U4328 = ~new_P2_ADD_1119_U72 | ~new_P2_U3019;
  assign new_P2_U4329 = ~new_P2_U3074;
  assign new_P2_U4330 = ~new_P2_U3035 | ~new_P2_U3064;
  assign new_P2_U4331 = ~new_P2_R1146_U12 | ~new_P2_U3931;
  assign new_P2_U4332 = ~new_P2_R1113_U12 | ~new_P2_U3930;
  assign new_P2_U4333 = ~new_P2_R1131_U114 | ~new_P2_U3926;
  assign new_P2_U4334 = ~new_P2_R1179_U12 | ~new_P2_U3941;
  assign new_P2_U4335 = ~new_P2_R1203_U12 | ~new_P2_U3943;
  assign new_P2_U4336 = ~new_P2_R1164_U114 | ~new_P2_U3014;
  assign new_P2_U4337 = ~new_P2_R1233_U114 | ~new_P2_U3922;
  assign new_P2_U4338 = ~new_P2_U3359;
  assign new_P2_U4339 = ~new_P2_R1275_U7 | ~new_P2_U3027;
  assign new_P2_U4340 = ~new_P2_U3026 | ~new_P2_U3074;
  assign new_P2_U4341 = ~new_P2_R1215_U115 | ~new_P2_U3025;
  assign new_P2_U4342 = ~new_P2_U3462 | ~new_P2_U4116;
  assign new_P2_U4343 = ~new_P2_U3621 | ~new_P2_U4338;
  assign new_P2_U4344 = ~P2_REG2_REG_13_ | ~new_P2_U3020;
  assign new_P2_U4345 = ~P2_REG1_REG_13_ | ~new_P2_U3021;
  assign new_P2_U4346 = ~P2_REG0_REG_13_ | ~new_P2_U3022;
  assign new_P2_U4347 = ~new_P2_ADD_1119_U71 | ~new_P2_U3019;
  assign new_P2_U4348 = ~new_P2_U3082;
  assign new_P2_U4349 = ~new_P2_U3035 | ~new_P2_U3065;
  assign new_P2_U4350 = ~new_P2_R1146_U102 | ~new_P2_U3931;
  assign new_P2_U4351 = ~new_P2_R1113_U102 | ~new_P2_U3930;
  assign new_P2_U4352 = ~new_P2_R1131_U113 | ~new_P2_U3926;
  assign new_P2_U4353 = ~new_P2_R1179_U102 | ~new_P2_U3941;
  assign new_P2_U4354 = ~new_P2_R1203_U102 | ~new_P2_U3943;
  assign new_P2_U4355 = ~new_P2_R1164_U113 | ~new_P2_U3014;
  assign new_P2_U4356 = ~new_P2_R1233_U113 | ~new_P2_U3922;
  assign new_P2_U4357 = ~new_P2_U3360;
  assign new_P2_U4358 = ~new_P2_R1275_U8 | ~new_P2_U3027;
  assign new_P2_U4359 = ~new_P2_U3026 | ~new_P2_U3082;
  assign new_P2_U4360 = ~new_P2_R1215_U114 | ~new_P2_U3025;
  assign new_P2_U4361 = ~new_P2_U3465 | ~new_P2_U4116;
  assign new_P2_U4362 = ~new_P2_U3625 | ~new_P2_U4357;
  assign new_P2_U4363 = ~P2_REG2_REG_14_ | ~new_P2_U3020;
  assign new_P2_U4364 = ~P2_REG1_REG_14_ | ~new_P2_U3021;
  assign new_P2_U4365 = ~P2_REG0_REG_14_ | ~new_P2_U3022;
  assign new_P2_U4366 = ~new_P2_ADD_1119_U70 | ~new_P2_U3019;
  assign new_P2_U4367 = ~new_P2_U3081;
  assign new_P2_U4368 = ~new_P2_U3035 | ~new_P2_U3074;
  assign new_P2_U4369 = ~new_P2_R1146_U101 | ~new_P2_U3931;
  assign new_P2_U4370 = ~new_P2_R1113_U101 | ~new_P2_U3930;
  assign new_P2_U4371 = ~new_P2_R1131_U11 | ~new_P2_U3926;
  assign new_P2_U4372 = ~new_P2_R1179_U101 | ~new_P2_U3941;
  assign new_P2_U4373 = ~new_P2_R1203_U101 | ~new_P2_U3943;
  assign new_P2_U4374 = ~new_P2_R1164_U11 | ~new_P2_U3014;
  assign new_P2_U4375 = ~new_P2_R1233_U11 | ~new_P2_U3922;
  assign new_P2_U4376 = ~new_P2_U3361;
  assign new_P2_U4377 = ~new_P2_R1275_U86 | ~new_P2_U3027;
  assign new_P2_U4378 = ~new_P2_U3026 | ~new_P2_U3081;
  assign new_P2_U4379 = ~new_P2_R1215_U12 | ~new_P2_U3025;
  assign new_P2_U4380 = ~new_P2_U3468 | ~new_P2_U4116;
  assign new_P2_U4381 = ~new_P2_U3629 | ~new_P2_U4376;
  assign new_P2_U4382 = ~P2_REG2_REG_15_ | ~new_P2_U3020;
  assign new_P2_U4383 = ~P2_REG1_REG_15_ | ~new_P2_U3021;
  assign new_P2_U4384 = ~P2_REG0_REG_15_ | ~new_P2_U3022;
  assign new_P2_U4385 = ~new_P2_ADD_1119_U69 | ~new_P2_U3019;
  assign new_P2_U4386 = ~new_P2_U3076;
  assign new_P2_U4387 = ~new_P2_U3035 | ~new_P2_U3082;
  assign new_P2_U4388 = ~new_P2_R1146_U112 | ~new_P2_U3931;
  assign new_P2_U4389 = ~new_P2_R1113_U112 | ~new_P2_U3930;
  assign new_P2_U4390 = ~new_P2_R1131_U112 | ~new_P2_U3926;
  assign new_P2_U4391 = ~new_P2_R1179_U112 | ~new_P2_U3941;
  assign new_P2_U4392 = ~new_P2_R1203_U112 | ~new_P2_U3943;
  assign new_P2_U4393 = ~new_P2_R1164_U112 | ~new_P2_U3014;
  assign new_P2_U4394 = ~new_P2_R1233_U112 | ~new_P2_U3922;
  assign new_P2_U4395 = ~new_P2_U3362;
  assign new_P2_U4396 = ~new_P2_R1275_U9 | ~new_P2_U3027;
  assign new_P2_U4397 = ~new_P2_U3026 | ~new_P2_U3076;
  assign new_P2_U4398 = ~new_P2_R1215_U113 | ~new_P2_U3025;
  assign new_P2_U4399 = ~new_P2_U3471 | ~new_P2_U4116;
  assign new_P2_U4400 = ~new_P2_U3633 | ~new_P2_U4395;
  assign new_P2_U4401 = ~P2_REG2_REG_16_ | ~new_P2_U3020;
  assign new_P2_U4402 = ~P2_REG1_REG_16_ | ~new_P2_U3021;
  assign new_P2_U4403 = ~P2_REG0_REG_16_ | ~new_P2_U3022;
  assign new_P2_U4404 = ~new_P2_ADD_1119_U68 | ~new_P2_U3019;
  assign new_P2_U4405 = ~new_P2_U3075;
  assign new_P2_U4406 = ~new_P2_U3035 | ~new_P2_U3081;
  assign new_P2_U4407 = ~new_P2_R1146_U111 | ~new_P2_U3931;
  assign new_P2_U4408 = ~new_P2_R1113_U111 | ~new_P2_U3930;
  assign new_P2_U4409 = ~new_P2_R1131_U111 | ~new_P2_U3926;
  assign new_P2_U4410 = ~new_P2_R1179_U111 | ~new_P2_U3941;
  assign new_P2_U4411 = ~new_P2_R1203_U111 | ~new_P2_U3943;
  assign new_P2_U4412 = ~new_P2_R1164_U111 | ~new_P2_U3014;
  assign new_P2_U4413 = ~new_P2_R1233_U111 | ~new_P2_U3922;
  assign new_P2_U4414 = ~new_P2_U3363;
  assign new_P2_U4415 = ~new_P2_R1275_U10 | ~new_P2_U3027;
  assign new_P2_U4416 = ~new_P2_U3026 | ~new_P2_U3075;
  assign new_P2_U4417 = ~new_P2_R1215_U112 | ~new_P2_U3025;
  assign new_P2_U4418 = ~new_P2_U3474 | ~new_P2_U4116;
  assign new_P2_U4419 = ~new_P2_U3637 | ~new_P2_U4414;
  assign new_P2_U4420 = ~P2_REG2_REG_17_ | ~new_P2_U3020;
  assign new_P2_U4421 = ~P2_REG1_REG_17_ | ~new_P2_U3021;
  assign new_P2_U4422 = ~P2_REG0_REG_17_ | ~new_P2_U3022;
  assign new_P2_U4423 = ~new_P2_ADD_1119_U67 | ~new_P2_U3019;
  assign new_P2_U4424 = ~new_P2_U3071;
  assign new_P2_U4425 = ~new_P2_U3035 | ~new_P2_U3076;
  assign new_P2_U4426 = ~new_P2_R1146_U13 | ~new_P2_U3931;
  assign new_P2_U4427 = ~new_P2_R1113_U13 | ~new_P2_U3930;
  assign new_P2_U4428 = ~new_P2_R1131_U110 | ~new_P2_U3926;
  assign new_P2_U4429 = ~new_P2_R1179_U13 | ~new_P2_U3941;
  assign new_P2_U4430 = ~new_P2_R1203_U13 | ~new_P2_U3943;
  assign new_P2_U4431 = ~new_P2_R1164_U110 | ~new_P2_U3014;
  assign new_P2_U4432 = ~new_P2_R1233_U110 | ~new_P2_U3922;
  assign new_P2_U4433 = ~new_P2_U3364;
  assign new_P2_U4434 = ~new_P2_R1275_U11 | ~new_P2_U3027;
  assign new_P2_U4435 = ~new_P2_U3026 | ~new_P2_U3071;
  assign new_P2_U4436 = ~new_P2_R1215_U111 | ~new_P2_U3025;
  assign new_P2_U4437 = ~new_P2_U3477 | ~new_P2_U4116;
  assign new_P2_U4438 = ~new_P2_U3641 | ~new_P2_U4433;
  assign new_P2_U4439 = ~P2_REG2_REG_18_ | ~new_P2_U3020;
  assign new_P2_U4440 = ~P2_REG1_REG_18_ | ~new_P2_U3021;
  assign new_P2_U4441 = ~P2_REG0_REG_18_ | ~new_P2_U3022;
  assign new_P2_U4442 = ~new_P2_ADD_1119_U66 | ~new_P2_U3019;
  assign new_P2_U4443 = ~new_P2_U3084;
  assign new_P2_U4444 = ~new_P2_U3035 | ~new_P2_U3075;
  assign new_P2_U4445 = ~new_P2_R1146_U100 | ~new_P2_U3931;
  assign new_P2_U4446 = ~new_P2_R1113_U100 | ~new_P2_U3930;
  assign new_P2_U4447 = ~new_P2_R1131_U12 | ~new_P2_U3926;
  assign new_P2_U4448 = ~new_P2_R1179_U100 | ~new_P2_U3941;
  assign new_P2_U4449 = ~new_P2_R1203_U100 | ~new_P2_U3943;
  assign new_P2_U4450 = ~new_P2_R1164_U12 | ~new_P2_U3014;
  assign new_P2_U4451 = ~new_P2_R1233_U12 | ~new_P2_U3922;
  assign new_P2_U4452 = ~new_P2_U3365;
  assign new_P2_U4453 = ~new_P2_R1275_U84 | ~new_P2_U3027;
  assign new_P2_U4454 = ~new_P2_U3026 | ~new_P2_U3084;
  assign new_P2_U4455 = ~new_P2_R1215_U13 | ~new_P2_U3025;
  assign new_P2_U4456 = ~new_P2_U3480 | ~new_P2_U4116;
  assign new_P2_U4457 = ~new_P2_U3645 | ~new_P2_U4452;
  assign new_P2_U4458 = ~P2_REG2_REG_19_ | ~new_P2_U3020;
  assign new_P2_U4459 = ~P2_REG1_REG_19_ | ~new_P2_U3021;
  assign new_P2_U4460 = ~P2_REG0_REG_19_ | ~new_P2_U3022;
  assign new_P2_U4461 = ~new_P2_ADD_1119_U65 | ~new_P2_U3019;
  assign new_P2_U4462 = ~new_P2_U3083;
  assign new_P2_U4463 = ~new_P2_U3035 | ~new_P2_U3071;
  assign new_P2_U4464 = ~new_P2_R1146_U99 | ~new_P2_U3931;
  assign new_P2_U4465 = ~new_P2_R1113_U99 | ~new_P2_U3930;
  assign new_P2_U4466 = ~new_P2_R1131_U109 | ~new_P2_U3926;
  assign new_P2_U4467 = ~new_P2_R1179_U99 | ~new_P2_U3941;
  assign new_P2_U4468 = ~new_P2_R1203_U99 | ~new_P2_U3943;
  assign new_P2_U4469 = ~new_P2_R1164_U109 | ~new_P2_U3014;
  assign new_P2_U4470 = ~new_P2_R1233_U109 | ~new_P2_U3922;
  assign new_P2_U4471 = ~new_P2_U3366;
  assign new_P2_U4472 = ~new_P2_R1275_U12 | ~new_P2_U3027;
  assign new_P2_U4473 = ~new_P2_U3026 | ~new_P2_U3083;
  assign new_P2_U4474 = ~new_P2_R1215_U110 | ~new_P2_U3025;
  assign new_P2_U4475 = ~new_P2_U3483 | ~new_P2_U4116;
  assign new_P2_U4476 = ~new_P2_U3649 | ~new_P2_U4471;
  assign new_P2_U4477 = ~P2_REG2_REG_20_ | ~new_P2_U3020;
  assign new_P2_U4478 = ~P2_REG1_REG_20_ | ~new_P2_U3021;
  assign new_P2_U4479 = ~P2_REG0_REG_20_ | ~new_P2_U3022;
  assign new_P2_U4480 = ~new_P2_ADD_1119_U64 | ~new_P2_U3019;
  assign new_P2_U4481 = ~new_P2_U3078;
  assign new_P2_U4482 = ~new_P2_U3035 | ~new_P2_U3084;
  assign new_P2_U4483 = ~new_P2_R1146_U98 | ~new_P2_U3931;
  assign new_P2_U4484 = ~new_P2_R1113_U98 | ~new_P2_U3930;
  assign new_P2_U4485 = ~new_P2_R1131_U108 | ~new_P2_U3926;
  assign new_P2_U4486 = ~new_P2_R1179_U98 | ~new_P2_U3941;
  assign new_P2_U4487 = ~new_P2_R1203_U98 | ~new_P2_U3943;
  assign new_P2_U4488 = ~new_P2_R1164_U108 | ~new_P2_U3014;
  assign new_P2_U4489 = ~new_P2_R1233_U108 | ~new_P2_U3922;
  assign new_P2_U4490 = ~new_P2_U3367;
  assign new_P2_U4491 = ~new_P2_R1275_U82 | ~new_P2_U3027;
  assign new_P2_U4492 = ~new_P2_U3026 | ~new_P2_U3078;
  assign new_P2_U4493 = ~new_P2_R1215_U109 | ~new_P2_U3025;
  assign new_P2_U4494 = ~new_P2_U3485 | ~new_P2_U4116;
  assign new_P2_U4495 = ~new_P2_U3653 | ~new_P2_U4490;
  assign new_P2_U4496 = ~P2_REG2_REG_21_ | ~new_P2_U3020;
  assign new_P2_U4497 = ~P2_REG1_REG_21_ | ~new_P2_U3021;
  assign new_P2_U4498 = ~P2_REG0_REG_21_ | ~new_P2_U3022;
  assign new_P2_U4499 = ~new_P2_ADD_1119_U63 | ~new_P2_U3019;
  assign new_P2_U4500 = ~new_P2_U3077;
  assign new_P2_U4501 = ~new_P2_U3035 | ~new_P2_U3083;
  assign new_P2_U4502 = ~new_P2_R1146_U96 | ~new_P2_U3931;
  assign new_P2_U4503 = ~new_P2_R1113_U96 | ~new_P2_U3930;
  assign new_P2_U4504 = ~new_P2_R1131_U13 | ~new_P2_U3926;
  assign new_P2_U4505 = ~new_P2_R1179_U96 | ~new_P2_U3941;
  assign new_P2_U4506 = ~new_P2_R1203_U96 | ~new_P2_U3943;
  assign new_P2_U4507 = ~new_P2_R1164_U13 | ~new_P2_U3014;
  assign new_P2_U4508 = ~new_P2_R1233_U13 | ~new_P2_U3922;
  assign new_P2_U4509 = ~new_P2_U3369;
  assign new_P2_U4510 = ~new_P2_R1275_U13 | ~new_P2_U3027;
  assign new_P2_U4511 = ~new_P2_U3026 | ~new_P2_U3077;
  assign new_P2_U4512 = ~new_P2_R1215_U14 | ~new_P2_U3025;
  assign new_P2_U4513 = ~new_P2_U3957 | ~new_P2_U4116;
  assign new_P2_U4514 = ~new_P2_U3657 | ~new_P2_U4509;
  assign new_P2_U4515 = ~P2_REG2_REG_22_ | ~new_P2_U3020;
  assign new_P2_U4516 = ~P2_REG1_REG_22_ | ~new_P2_U3021;
  assign new_P2_U4517 = ~P2_REG0_REG_22_ | ~new_P2_U3022;
  assign new_P2_U4518 = ~new_P2_ADD_1119_U62 | ~new_P2_U3019;
  assign new_P2_U4519 = ~new_P2_U3063;
  assign new_P2_U4520 = ~new_P2_U3035 | ~new_P2_U3078;
  assign new_P2_U4521 = ~new_P2_R1146_U110 | ~new_P2_U3931;
  assign new_P2_U4522 = ~new_P2_R1113_U110 | ~new_P2_U3930;
  assign new_P2_U4523 = ~new_P2_R1131_U14 | ~new_P2_U3926;
  assign new_P2_U4524 = ~new_P2_R1179_U110 | ~new_P2_U3941;
  assign new_P2_U4525 = ~new_P2_R1203_U110 | ~new_P2_U3943;
  assign new_P2_U4526 = ~new_P2_R1164_U14 | ~new_P2_U3014;
  assign new_P2_U4527 = ~new_P2_R1233_U14 | ~new_P2_U3922;
  assign new_P2_U4528 = ~new_P2_U3371;
  assign new_P2_U4529 = ~new_P2_R1275_U78 | ~new_P2_U3027;
  assign new_P2_U4530 = ~new_P2_U3026 | ~new_P2_U3063;
  assign new_P2_U4531 = ~new_P2_R1215_U15 | ~new_P2_U3025;
  assign new_P2_U4532 = ~new_P2_U3956 | ~new_P2_U4116;
  assign new_P2_U4533 = ~new_P2_U3661 | ~new_P2_U4528;
  assign new_P2_U4534 = ~P2_REG2_REG_23_ | ~new_P2_U3020;
  assign new_P2_U4535 = ~P2_REG1_REG_23_ | ~new_P2_U3021;
  assign new_P2_U4536 = ~P2_REG0_REG_23_ | ~new_P2_U3022;
  assign new_P2_U4537 = ~new_P2_ADD_1119_U61 | ~new_P2_U3019;
  assign new_P2_U4538 = ~new_P2_U3068;
  assign new_P2_U4539 = ~new_P2_U3035 | ~new_P2_U3077;
  assign new_P2_U4540 = ~new_P2_R1146_U109 | ~new_P2_U3931;
  assign new_P2_U4541 = ~new_P2_R1113_U109 | ~new_P2_U3930;
  assign new_P2_U4542 = ~new_P2_R1131_U107 | ~new_P2_U3926;
  assign new_P2_U4543 = ~new_P2_R1179_U109 | ~new_P2_U3941;
  assign new_P2_U4544 = ~new_P2_R1203_U109 | ~new_P2_U3943;
  assign new_P2_U4545 = ~new_P2_R1164_U107 | ~new_P2_U3014;
  assign new_P2_U4546 = ~new_P2_R1233_U107 | ~new_P2_U3922;
  assign new_P2_U4547 = ~new_P2_U3373;
  assign new_P2_U4548 = ~new_P2_R1275_U14 | ~new_P2_U3027;
  assign new_P2_U4549 = ~new_P2_U3026 | ~new_P2_U3068;
  assign new_P2_U4550 = ~new_P2_R1215_U108 | ~new_P2_U3025;
  assign new_P2_U4551 = ~new_P2_U3955 | ~new_P2_U4116;
  assign new_P2_U4552 = ~new_P2_U3665 | ~new_P2_U4547;
  assign new_P2_U4553 = ~P2_REG2_REG_24_ | ~new_P2_U3020;
  assign new_P2_U4554 = ~P2_REG1_REG_24_ | ~new_P2_U3021;
  assign new_P2_U4555 = ~P2_REG0_REG_24_ | ~new_P2_U3022;
  assign new_P2_U4556 = ~new_P2_ADD_1119_U60 | ~new_P2_U3019;
  assign new_P2_U4557 = ~new_P2_U3067;
  assign new_P2_U4558 = ~new_P2_U3035 | ~new_P2_U3063;
  assign new_P2_U4559 = ~new_P2_R1146_U14 | ~new_P2_U3931;
  assign new_P2_U4560 = ~new_P2_R1113_U14 | ~new_P2_U3930;
  assign new_P2_U4561 = ~new_P2_R1131_U106 | ~new_P2_U3926;
  assign new_P2_U4562 = ~new_P2_R1179_U14 | ~new_P2_U3941;
  assign new_P2_U4563 = ~new_P2_R1203_U14 | ~new_P2_U3943;
  assign new_P2_U4564 = ~new_P2_R1164_U106 | ~new_P2_U3014;
  assign new_P2_U4565 = ~new_P2_R1233_U106 | ~new_P2_U3922;
  assign new_P2_U4566 = ~new_P2_U3375;
  assign new_P2_U4567 = ~new_P2_R1275_U76 | ~new_P2_U3027;
  assign new_P2_U4568 = ~new_P2_U3026 | ~new_P2_U3067;
  assign new_P2_U4569 = ~new_P2_R1215_U107 | ~new_P2_U3025;
  assign new_P2_U4570 = ~new_P2_U3954 | ~new_P2_U4116;
  assign new_P2_U4571 = ~new_P2_U3669 | ~new_P2_U4566;
  assign new_P2_U4572 = ~P2_REG2_REG_25_ | ~new_P2_U3020;
  assign new_P2_U4573 = ~P2_REG1_REG_25_ | ~new_P2_U3021;
  assign new_P2_U4574 = ~P2_REG0_REG_25_ | ~new_P2_U3022;
  assign new_P2_U4575 = ~new_P2_ADD_1119_U59 | ~new_P2_U3019;
  assign new_P2_U4576 = ~new_P2_U3060;
  assign new_P2_U4577 = ~new_P2_U3035 | ~new_P2_U3068;
  assign new_P2_U4578 = ~new_P2_R1146_U95 | ~new_P2_U3931;
  assign new_P2_U4579 = ~new_P2_R1113_U95 | ~new_P2_U3930;
  assign new_P2_U4580 = ~new_P2_R1131_U105 | ~new_P2_U3926;
  assign new_P2_U4581 = ~new_P2_R1179_U95 | ~new_P2_U3941;
  assign new_P2_U4582 = ~new_P2_R1203_U95 | ~new_P2_U3943;
  assign new_P2_U4583 = ~new_P2_R1164_U105 | ~new_P2_U3014;
  assign new_P2_U4584 = ~new_P2_R1233_U105 | ~new_P2_U3922;
  assign new_P2_U4585 = ~new_P2_U3377;
  assign new_P2_U4586 = ~new_P2_R1275_U15 | ~new_P2_U3027;
  assign new_P2_U4587 = ~new_P2_U3026 | ~new_P2_U3060;
  assign new_P2_U4588 = ~new_P2_R1215_U106 | ~new_P2_U3025;
  assign new_P2_U4589 = ~new_P2_U3953 | ~new_P2_U4116;
  assign new_P2_U4590 = ~new_P2_U3673 | ~new_P2_U4585;
  assign new_P2_U4591 = ~P2_REG2_REG_26_ | ~new_P2_U3020;
  assign new_P2_U4592 = ~P2_REG1_REG_26_ | ~new_P2_U3021;
  assign new_P2_U4593 = ~P2_REG0_REG_26_ | ~new_P2_U3022;
  assign new_P2_U4594 = ~new_P2_ADD_1119_U58 | ~new_P2_U3019;
  assign new_P2_U4595 = ~new_P2_U3059;
  assign new_P2_U4596 = ~new_P2_U3035 | ~new_P2_U3067;
  assign new_P2_U4597 = ~new_P2_R1146_U94 | ~new_P2_U3931;
  assign new_P2_U4598 = ~new_P2_R1113_U94 | ~new_P2_U3930;
  assign new_P2_U4599 = ~new_P2_R1131_U104 | ~new_P2_U3926;
  assign new_P2_U4600 = ~new_P2_R1179_U94 | ~new_P2_U3941;
  assign new_P2_U4601 = ~new_P2_R1203_U94 | ~new_P2_U3943;
  assign new_P2_U4602 = ~new_P2_R1164_U104 | ~new_P2_U3014;
  assign new_P2_U4603 = ~new_P2_R1233_U104 | ~new_P2_U3922;
  assign new_P2_U4604 = ~new_P2_U3379;
  assign new_P2_U4605 = ~new_P2_R1275_U74 | ~new_P2_U3027;
  assign new_P2_U4606 = ~new_P2_U3026 | ~new_P2_U3059;
  assign new_P2_U4607 = ~new_P2_R1215_U105 | ~new_P2_U3025;
  assign new_P2_U4608 = ~new_P2_U3952 | ~new_P2_U4116;
  assign new_P2_U4609 = ~new_P2_U3677 | ~new_P2_U4604;
  assign new_P2_U4610 = ~P2_REG2_REG_27_ | ~new_P2_U3020;
  assign new_P2_U4611 = ~P2_REG1_REG_27_ | ~new_P2_U3021;
  assign new_P2_U4612 = ~P2_REG0_REG_27_ | ~new_P2_U3022;
  assign new_P2_U4613 = ~new_P2_ADD_1119_U57 | ~new_P2_U3019;
  assign new_P2_U4614 = ~new_P2_U3055;
  assign new_P2_U4615 = ~new_P2_U3035 | ~new_P2_U3060;
  assign new_P2_U4616 = ~new_P2_R1146_U108 | ~new_P2_U3931;
  assign new_P2_U4617 = ~new_P2_R1113_U108 | ~new_P2_U3930;
  assign new_P2_U4618 = ~new_P2_R1131_U15 | ~new_P2_U3926;
  assign new_P2_U4619 = ~new_P2_R1179_U108 | ~new_P2_U3941;
  assign new_P2_U4620 = ~new_P2_R1203_U108 | ~new_P2_U3943;
  assign new_P2_U4621 = ~new_P2_R1164_U15 | ~new_P2_U3014;
  assign new_P2_U4622 = ~new_P2_R1233_U15 | ~new_P2_U3922;
  assign new_P2_U4623 = ~new_P2_U3381;
  assign new_P2_U4624 = ~new_P2_R1275_U16 | ~new_P2_U3027;
  assign new_P2_U4625 = ~new_P2_U3026 | ~new_P2_U3055;
  assign new_P2_U4626 = ~new_P2_R1215_U16 | ~new_P2_U3025;
  assign new_P2_U4627 = ~new_P2_U3951 | ~new_P2_U4116;
  assign new_P2_U4628 = ~new_P2_U3681 | ~new_P2_U4623;
  assign new_P2_U4629 = ~P2_REG2_REG_28_ | ~new_P2_U3020;
  assign new_P2_U4630 = ~P2_REG1_REG_28_ | ~new_P2_U3021;
  assign new_P2_U4631 = ~P2_REG0_REG_28_ | ~new_P2_U3022;
  assign new_P2_U4632 = ~new_P2_ADD_1119_U56 | ~new_P2_U3019;
  assign new_P2_U4633 = ~new_P2_U3056;
  assign new_P2_U4634 = ~new_P2_U3035 | ~new_P2_U3059;
  assign new_P2_U4635 = ~new_P2_R1146_U15 | ~new_P2_U3931;
  assign new_P2_U4636 = ~new_P2_R1113_U15 | ~new_P2_U3930;
  assign new_P2_U4637 = ~new_P2_R1131_U103 | ~new_P2_U3926;
  assign new_P2_U4638 = ~new_P2_R1179_U15 | ~new_P2_U3941;
  assign new_P2_U4639 = ~new_P2_R1203_U15 | ~new_P2_U3943;
  assign new_P2_U4640 = ~new_P2_R1164_U103 | ~new_P2_U3014;
  assign new_P2_U4641 = ~new_P2_R1233_U103 | ~new_P2_U3922;
  assign new_P2_U4642 = ~new_P2_U3383;
  assign new_P2_U4643 = ~new_P2_R1275_U72 | ~new_P2_U3027;
  assign new_P2_U4644 = ~new_P2_U3026 | ~new_P2_U3056;
  assign new_P2_U4645 = ~new_P2_R1215_U104 | ~new_P2_U3025;
  assign new_P2_U4646 = ~new_P2_U3950 | ~new_P2_U4116;
  assign new_P2_U4647 = ~new_P2_U3685 | ~new_P2_U4642;
  assign new_P2_U4648 = ~new_P2_ADD_1119_U5 | ~new_P2_U3019;
  assign new_P2_U4649 = ~P2_REG2_REG_29_ | ~new_P2_U3020;
  assign new_P2_U4650 = ~P2_REG1_REG_29_ | ~new_P2_U3021;
  assign new_P2_U4651 = ~P2_REG0_REG_29_ | ~new_P2_U3022;
  assign new_P2_U4652 = ~new_P2_U3057;
  assign new_P2_U4653 = ~new_P2_U3035 | ~new_P2_U3055;
  assign new_P2_U4654 = ~new_P2_R1146_U93 | ~new_P2_U3931;
  assign new_P2_U4655 = ~new_P2_R1113_U93 | ~new_P2_U3930;
  assign new_P2_U4656 = ~new_P2_R1131_U102 | ~new_P2_U3926;
  assign new_P2_U4657 = ~new_P2_R1179_U93 | ~new_P2_U3941;
  assign new_P2_U4658 = ~new_P2_R1203_U93 | ~new_P2_U3943;
  assign new_P2_U4659 = ~new_P2_R1164_U102 | ~new_P2_U3014;
  assign new_P2_U4660 = ~new_P2_R1233_U102 | ~new_P2_U3922;
  assign new_P2_U4661 = ~new_P2_U3385;
  assign new_P2_U4662 = ~new_P2_R1275_U17 | ~new_P2_U3027;
  assign new_P2_U4663 = ~new_P2_U3026 | ~new_P2_U3057;
  assign new_P2_U4664 = ~new_P2_R1215_U103 | ~new_P2_U3025;
  assign new_P2_U4665 = ~new_P2_U3949 | ~new_P2_U4116;
  assign new_P2_U4666 = ~new_P2_U3688 | ~new_P2_U4661;
  assign new_P2_U4667 = ~P2_REG2_REG_30_ | ~new_P2_U3020;
  assign new_P2_U4668 = ~P2_REG1_REG_30_ | ~new_P2_U3021;
  assign new_P2_U4669 = ~P2_REG0_REG_30_ | ~new_P2_U3022;
  assign new_P2_U4670 = ~new_P2_U3061;
  assign new_P2_U4671 = ~new_P2_U5683 | ~new_P2_U3331;
  assign new_P2_U4672 = ~new_P2_U3347 | ~new_P2_U4671;
  assign new_P2_U4673 = ~new_P2_U3689 | ~new_P2_U3061;
  assign new_P2_U4674 = ~new_P2_U3035 | ~new_P2_U3056;
  assign new_P2_U4675 = ~new_P2_R1146_U16 | ~new_P2_U3931;
  assign new_P2_U4676 = ~new_P2_R1113_U16 | ~new_P2_U3930;
  assign new_P2_U4677 = ~new_P2_R1131_U101 | ~new_P2_U3926;
  assign new_P2_U4678 = ~new_P2_R1179_U16 | ~new_P2_U3941;
  assign new_P2_U4679 = ~new_P2_R1203_U16 | ~new_P2_U3943;
  assign new_P2_U4680 = ~new_P2_R1164_U101 | ~new_P2_U3014;
  assign new_P2_U4681 = ~new_P2_R1233_U101 | ~new_P2_U3922;
  assign new_P2_U4682 = ~new_P2_U3387;
  assign new_P2_U4683 = ~new_P2_R1275_U70 | ~new_P2_U3027;
  assign new_P2_U4684 = ~new_P2_R1215_U102 | ~new_P2_U3025;
  assign new_P2_U4685 = ~new_P2_U3960 | ~new_P2_U4116;
  assign new_P2_U4686 = ~new_P2_U3693 | ~new_P2_U4682;
  assign new_P2_U4687 = ~P2_REG2_REG_31_ | ~new_P2_U3020;
  assign new_P2_U4688 = ~P2_REG1_REG_31_ | ~new_P2_U3021;
  assign new_P2_U4689 = ~P2_REG0_REG_31_ | ~new_P2_U3022;
  assign new_P2_U4690 = ~new_P2_U3058;
  assign new_P2_U4691 = ~new_P2_R1275_U19 | ~new_P2_U3027;
  assign new_P2_U4692 = ~new_P2_U3959 | ~new_P2_U4116;
  assign new_P2_U4693 = ~new_P2_U4691 | ~new_P2_U4692 | ~new_P2_U3913;
  assign new_P2_U4694 = ~new_P2_R1275_U68 | ~new_P2_U3027;
  assign new_P2_U4695 = ~new_P2_U3958 | ~new_P2_U4116;
  assign new_P2_U4696 = ~new_P2_U4694 | ~new_P2_U4695 | ~new_P2_U3913;
  assign new_P2_U4697 = ~new_P2_U3696 | ~new_P2_U3016;
  assign new_P2_U4698 = ~new_P2_U3393 | ~new_P2_U4697;
  assign new_P2_U4699 = ~new_P2_U3921 | ~new_P2_U3418;
  assign new_P2_U4700 = ~new_P2_U3398;
  assign new_P2_U4701 = ~new_P2_U3037 | ~new_P2_U3080;
  assign new_P2_U4702 = ~new_P2_U3034 | ~new_P2_R1215_U96;
  assign new_P2_U4703 = ~new_P2_U3033 | ~P2_REG3_REG_0_;
  assign new_P2_U4704 = ~new_P2_U3032 | ~new_P2_U3427;
  assign new_P2_U4705 = ~new_P2_U3031 | ~new_P2_U3427;
  assign new_P2_U4706 = ~new_P2_U3037 | ~new_P2_U3070;
  assign new_P2_U4707 = ~new_P2_U3034 | ~new_P2_R1215_U95;
  assign new_P2_U4708 = ~new_P2_U3033 | ~P2_REG3_REG_1_;
  assign new_P2_U4709 = ~new_P2_U3032 | ~new_P2_U3432;
  assign new_P2_U4710 = ~new_P2_U3031 | ~new_P2_R1275_U55;
  assign new_P2_U4711 = ~new_P2_U3037 | ~new_P2_U3066;
  assign new_P2_U4712 = ~new_P2_U3034 | ~new_P2_R1215_U17;
  assign new_P2_U4713 = ~new_P2_U3033 | ~P2_REG3_REG_2_;
  assign new_P2_U4714 = ~new_P2_U3032 | ~new_P2_U3435;
  assign new_P2_U4715 = ~new_P2_U3031 | ~new_P2_R1275_U18;
  assign new_P2_U4716 = ~new_P2_U3037 | ~new_P2_U3062;
  assign new_P2_U4717 = ~new_P2_U3034 | ~new_P2_R1215_U101;
  assign new_P2_U4718 = ~new_P2_U3033 | ~new_P2_ADD_1119_U4;
  assign new_P2_U4719 = ~new_P2_U3032 | ~new_P2_U3438;
  assign new_P2_U4720 = ~new_P2_U3031 | ~new_P2_R1275_U20;
  assign new_P2_U4721 = ~new_P2_U3037 | ~new_P2_U3069;
  assign new_P2_U4722 = ~new_P2_U3034 | ~new_P2_R1215_U100;
  assign new_P2_U4723 = ~new_P2_U3033 | ~new_P2_ADD_1119_U55;
  assign new_P2_U4724 = ~new_P2_U3032 | ~new_P2_U3441;
  assign new_P2_U4725 = ~new_P2_U3031 | ~new_P2_R1275_U21;
  assign new_P2_U4726 = ~new_P2_U3037 | ~new_P2_U3073;
  assign new_P2_U4727 = ~new_P2_U3034 | ~new_P2_R1215_U18;
  assign new_P2_U4728 = ~new_P2_U3033 | ~new_P2_ADD_1119_U54;
  assign new_P2_U4729 = ~new_P2_U3032 | ~new_P2_U3444;
  assign new_P2_U4730 = ~new_P2_U3031 | ~new_P2_R1275_U65;
  assign new_P2_U4731 = ~new_P2_U3037 | ~new_P2_U3072;
  assign new_P2_U4732 = ~new_P2_U3034 | ~new_P2_R1215_U99;
  assign new_P2_U4733 = ~new_P2_U3033 | ~new_P2_ADD_1119_U53;
  assign new_P2_U4734 = ~new_P2_U3032 | ~new_P2_U3447;
  assign new_P2_U4735 = ~new_P2_U3031 | ~new_P2_R1275_U22;
  assign new_P2_U4736 = ~new_P2_U3037 | ~new_P2_U3086;
  assign new_P2_U4737 = ~new_P2_U3034 | ~new_P2_R1215_U19;
  assign new_P2_U4738 = ~new_P2_U3033 | ~new_P2_ADD_1119_U52;
  assign new_P2_U4739 = ~new_P2_U3032 | ~new_P2_U3450;
  assign new_P2_U4740 = ~new_P2_U3031 | ~new_P2_R1275_U23;
  assign new_P2_U4741 = ~new_P2_U3037 | ~new_P2_U3085;
  assign new_P2_U4742 = ~new_P2_U3034 | ~new_P2_R1215_U98;
  assign new_P2_U4743 = ~new_P2_U3033 | ~new_P2_ADD_1119_U51;
  assign new_P2_U4744 = ~new_P2_U3032 | ~new_P2_U3453;
  assign new_P2_U4745 = ~new_P2_U3031 | ~new_P2_R1275_U24;
  assign new_P2_U4746 = ~new_P2_U3037 | ~new_P2_U3064;
  assign new_P2_U4747 = ~new_P2_U3034 | ~new_P2_R1215_U97;
  assign new_P2_U4748 = ~new_P2_U3033 | ~new_P2_ADD_1119_U50;
  assign new_P2_U4749 = ~new_P2_U3032 | ~new_P2_U3456;
  assign new_P2_U4750 = ~new_P2_U3031 | ~new_P2_R1275_U63;
  assign new_P2_U4751 = ~new_P2_U3037 | ~new_P2_U3065;
  assign new_P2_U4752 = ~new_P2_U3034 | ~new_P2_R1215_U11;
  assign new_P2_U4753 = ~new_P2_U3033 | ~new_P2_ADD_1119_U74;
  assign new_P2_U4754 = ~new_P2_U3032 | ~new_P2_U3459;
  assign new_P2_U4755 = ~new_P2_U3031 | ~new_P2_R1275_U6;
  assign new_P2_U4756 = ~new_P2_U3037 | ~new_P2_U3074;
  assign new_P2_U4757 = ~new_P2_U3034 | ~new_P2_R1215_U115;
  assign new_P2_U4758 = ~new_P2_U3033 | ~new_P2_ADD_1119_U73;
  assign new_P2_U4759 = ~new_P2_U3032 | ~new_P2_U3462;
  assign new_P2_U4760 = ~new_P2_U3031 | ~new_P2_R1275_U7;
  assign new_P2_U4761 = ~new_P2_U3037 | ~new_P2_U3082;
  assign new_P2_U4762 = ~new_P2_U3034 | ~new_P2_R1215_U114;
  assign new_P2_U4763 = ~new_P2_U3033 | ~new_P2_ADD_1119_U72;
  assign new_P2_U4764 = ~new_P2_U3032 | ~new_P2_U3465;
  assign new_P2_U4765 = ~new_P2_U3031 | ~new_P2_R1275_U8;
  assign new_P2_U4766 = ~new_P2_U3037 | ~new_P2_U3081;
  assign new_P2_U4767 = ~new_P2_U3034 | ~new_P2_R1215_U12;
  assign new_P2_U4768 = ~new_P2_U3033 | ~new_P2_ADD_1119_U71;
  assign new_P2_U4769 = ~new_P2_U3032 | ~new_P2_U3468;
  assign new_P2_U4770 = ~new_P2_U3031 | ~new_P2_R1275_U86;
  assign new_P2_U4771 = ~new_P2_U3037 | ~new_P2_U3076;
  assign new_P2_U4772 = ~new_P2_U3034 | ~new_P2_R1215_U113;
  assign new_P2_U4773 = ~new_P2_U3033 | ~new_P2_ADD_1119_U70;
  assign new_P2_U4774 = ~new_P2_U3032 | ~new_P2_U3471;
  assign new_P2_U4775 = ~new_P2_U3031 | ~new_P2_R1275_U9;
  assign new_P2_U4776 = ~new_P2_U3037 | ~new_P2_U3075;
  assign new_P2_U4777 = ~new_P2_U3034 | ~new_P2_R1215_U112;
  assign new_P2_U4778 = ~new_P2_U3033 | ~new_P2_ADD_1119_U69;
  assign new_P2_U4779 = ~new_P2_U3032 | ~new_P2_U3474;
  assign new_P2_U4780 = ~new_P2_U3031 | ~new_P2_R1275_U10;
  assign new_P2_U4781 = ~new_P2_U3037 | ~new_P2_U3071;
  assign new_P2_U4782 = ~new_P2_U3034 | ~new_P2_R1215_U111;
  assign new_P2_U4783 = ~new_P2_U3033 | ~new_P2_ADD_1119_U68;
  assign new_P2_U4784 = ~new_P2_U3032 | ~new_P2_U3477;
  assign new_P2_U4785 = ~new_P2_U3031 | ~new_P2_R1275_U11;
  assign new_P2_U4786 = ~new_P2_U3037 | ~new_P2_U3084;
  assign new_P2_U4787 = ~new_P2_U3034 | ~new_P2_R1215_U13;
  assign new_P2_U4788 = ~new_P2_U3033 | ~new_P2_ADD_1119_U67;
  assign new_P2_U4789 = ~new_P2_U3032 | ~new_P2_U3480;
  assign new_P2_U4790 = ~new_P2_U3031 | ~new_P2_R1275_U84;
  assign new_P2_U4791 = ~new_P2_U3037 | ~new_P2_U3083;
  assign new_P2_U4792 = ~new_P2_U3034 | ~new_P2_R1215_U110;
  assign new_P2_U4793 = ~new_P2_U3033 | ~new_P2_ADD_1119_U66;
  assign new_P2_U4794 = ~new_P2_U3032 | ~new_P2_U3483;
  assign new_P2_U4795 = ~new_P2_U3031 | ~new_P2_R1275_U12;
  assign new_P2_U4796 = ~new_P2_U3037 | ~new_P2_U3078;
  assign new_P2_U4797 = ~new_P2_U3034 | ~new_P2_R1215_U109;
  assign new_P2_U4798 = ~new_P2_U3033 | ~new_P2_ADD_1119_U65;
  assign new_P2_U4799 = ~new_P2_U3032 | ~new_P2_U3485;
  assign new_P2_U4800 = ~new_P2_U3031 | ~new_P2_R1275_U82;
  assign new_P2_U4801 = ~new_P2_U3037 | ~new_P2_U3077;
  assign new_P2_U4802 = ~new_P2_U3034 | ~new_P2_R1215_U14;
  assign new_P2_U4803 = ~new_P2_U3033 | ~new_P2_ADD_1119_U64;
  assign new_P2_U4804 = ~new_P2_U3032 | ~new_P2_U3957;
  assign new_P2_U4805 = ~new_P2_U3031 | ~new_P2_R1275_U13;
  assign new_P2_U4806 = ~new_P2_U3037 | ~new_P2_U3063;
  assign new_P2_U4807 = ~new_P2_U3034 | ~new_P2_R1215_U15;
  assign new_P2_U4808 = ~new_P2_U3033 | ~new_P2_ADD_1119_U63;
  assign new_P2_U4809 = ~new_P2_U3032 | ~new_P2_U3956;
  assign new_P2_U4810 = ~new_P2_U3031 | ~new_P2_R1275_U78;
  assign new_P2_U4811 = ~new_P2_U3037 | ~new_P2_U3068;
  assign new_P2_U4812 = ~new_P2_U3034 | ~new_P2_R1215_U108;
  assign new_P2_U4813 = ~new_P2_U3033 | ~new_P2_ADD_1119_U62;
  assign new_P2_U4814 = ~new_P2_U3032 | ~new_P2_U3955;
  assign new_P2_U4815 = ~new_P2_U3031 | ~new_P2_R1275_U14;
  assign new_P2_U4816 = ~new_P2_U3037 | ~new_P2_U3067;
  assign new_P2_U4817 = ~new_P2_U3034 | ~new_P2_R1215_U107;
  assign new_P2_U4818 = ~new_P2_U3033 | ~new_P2_ADD_1119_U61;
  assign new_P2_U4819 = ~new_P2_U3032 | ~new_P2_U3954;
  assign new_P2_U4820 = ~new_P2_U3031 | ~new_P2_R1275_U76;
  assign new_P2_U4821 = ~new_P2_U3037 | ~new_P2_U3060;
  assign new_P2_U4822 = ~new_P2_U3034 | ~new_P2_R1215_U106;
  assign new_P2_U4823 = ~new_P2_U3033 | ~new_P2_ADD_1119_U60;
  assign new_P2_U4824 = ~new_P2_U3032 | ~new_P2_U3953;
  assign new_P2_U4825 = ~new_P2_U3031 | ~new_P2_R1275_U15;
  assign new_P2_U4826 = ~new_P2_U3037 | ~new_P2_U3059;
  assign new_P2_U4827 = ~new_P2_U3034 | ~new_P2_R1215_U105;
  assign new_P2_U4828 = ~new_P2_U3033 | ~new_P2_ADD_1119_U59;
  assign new_P2_U4829 = ~new_P2_U3032 | ~new_P2_U3952;
  assign new_P2_U4830 = ~new_P2_U3031 | ~new_P2_R1275_U74;
  assign new_P2_U4831 = ~new_P2_U3037 | ~new_P2_U3055;
  assign new_P2_U4832 = ~new_P2_U3034 | ~new_P2_R1215_U16;
  assign new_P2_U4833 = ~new_P2_U3033 | ~new_P2_ADD_1119_U58;
  assign new_P2_U4834 = ~new_P2_U3032 | ~new_P2_U3951;
  assign new_P2_U4835 = ~new_P2_U3031 | ~new_P2_R1275_U16;
  assign new_P2_U4836 = ~new_P2_U3037 | ~new_P2_U3056;
  assign new_P2_U4837 = ~new_P2_U3034 | ~new_P2_R1215_U104;
  assign new_P2_U4838 = ~new_P2_U3033 | ~new_P2_ADD_1119_U57;
  assign new_P2_U4839 = ~new_P2_U3032 | ~new_P2_U3950;
  assign new_P2_U4840 = ~new_P2_U3031 | ~new_P2_R1275_U72;
  assign new_P2_U4841 = ~new_P2_U3037 | ~new_P2_U3057;
  assign new_P2_U4842 = ~new_P2_U3034 | ~new_P2_R1215_U103;
  assign new_P2_U4843 = ~new_P2_U3033 | ~new_P2_ADD_1119_U56;
  assign new_P2_U4844 = ~new_P2_U3032 | ~new_P2_U3949;
  assign new_P2_U4845 = ~new_P2_U3031 | ~new_P2_R1275_U17;
  assign new_P2_U4846 = ~new_P2_U3034 | ~new_P2_R1215_U102;
  assign new_P2_U4847 = ~new_P2_U3033 | ~new_P2_ADD_1119_U5;
  assign new_P2_U4848 = ~new_P2_U3032 | ~new_P2_U3960;
  assign new_P2_U4849 = ~new_P2_U3031 | ~new_P2_R1275_U70;
  assign new_P2_U4850 = ~new_P2_U3032 | ~new_P2_U3959;
  assign new_P2_U4851 = ~new_P2_U3031 | ~new_P2_R1275_U19;
  assign new_P2_U4852 = ~new_P2_U3032 | ~new_P2_U3958;
  assign new_P2_U4853 = ~new_P2_U3031 | ~new_P2_R1275_U68;
  assign new_P2_U4854 = ~new_P2_U3393 | ~new_P2_U4700 | ~new_P2_U3051 | ~new_P2_U3755 | ~new_P2_U3395;
  assign new_P2_U4855 = ~new_P2_R1170_U13 | ~new_P2_U3043;
  assign new_P2_U4856 = ~new_P2_U3041 | ~new_P2_U3424;
  assign new_P2_U4857 = ~new_P2_R1209_U13 | ~new_P2_U3039;
  assign new_P2_U4858 = ~new_P2_U4857 | ~new_P2_U4856 | ~new_P2_U4855;
  assign new_P2_U4859 = ~new_P2_R1170_U13 | ~new_P2_U3018;
  assign new_P2_U4860 = ~new_P2_U3017 | ~new_P2_R1209_U13;
  assign new_P2_U4861 = ~new_P2_U5683 | ~new_P2_U3424;
  assign new_P2_U4862 = ~new_P2_U4861 | ~new_P2_U4860 | ~new_P2_U4859;
  assign new_P2_U4863 = ~new_P2_U3401;
  assign new_P2_U4864 = ~new_P2_U3045 | ~new_P2_U4858;
  assign new_P2_U4865 = ~n2619 | ~new_P2_U4862;
  assign new_P2_U4866 = ~new_P2_U3044 | ~new_P2_R1170_U13;
  assign new_P2_U4867 = ~P2_REG3_REG_19_ | ~n2609;
  assign new_P2_U4868 = ~new_P2_U3042 | ~new_P2_U3424;
  assign new_P2_U4869 = ~new_P2_U3040 | ~new_P2_R1209_U13;
  assign new_P2_U4870 = ~P2_ADDR_REG_19_ | ~new_P2_U4863;
  assign new_P2_U4871 = ~new_P2_R1170_U75 | ~new_P2_U3043;
  assign new_P2_U4872 = ~new_P2_U3041 | ~new_P2_U3482;
  assign new_P2_U4873 = ~new_P2_R1209_U75 | ~new_P2_U3039;
  assign new_P2_U4874 = ~new_P2_U4873 | ~new_P2_U4872 | ~new_P2_U4871;
  assign new_P2_U4875 = ~new_P2_R1170_U75 | ~new_P2_U3018;
  assign new_P2_U4876 = ~new_P2_R1209_U75 | ~new_P2_U3017;
  assign new_P2_U4877 = ~new_P2_U5683 | ~new_P2_U3482;
  assign new_P2_U4878 = ~new_P2_U4877 | ~new_P2_U4876 | ~new_P2_U4875;
  assign new_P2_U4879 = ~new_P2_U3045 | ~new_P2_U4874;
  assign new_P2_U4880 = ~n2619 | ~new_P2_U4878;
  assign new_P2_U4881 = ~new_P2_R1170_U75 | ~new_P2_U3044;
  assign new_P2_U4882 = ~P2_REG3_REG_18_ | ~n2609;
  assign new_P2_U4883 = ~new_P2_U3042 | ~new_P2_U3482;
  assign new_P2_U4884 = ~new_P2_R1209_U75 | ~new_P2_U3040;
  assign new_P2_U4885 = ~P2_ADDR_REG_18_ | ~new_P2_U4863;
  assign new_P2_U4886 = ~new_P2_R1170_U12 | ~new_P2_U3043;
  assign new_P2_U4887 = ~new_P2_U3041 | ~new_P2_U3479;
  assign new_P2_U4888 = ~new_P2_R1209_U12 | ~new_P2_U3039;
  assign new_P2_U4889 = ~new_P2_U4888 | ~new_P2_U4887 | ~new_P2_U4886;
  assign new_P2_U4890 = ~new_P2_R1170_U12 | ~new_P2_U3018;
  assign new_P2_U4891 = ~new_P2_R1209_U12 | ~new_P2_U3017;
  assign new_P2_U4892 = ~new_P2_U5683 | ~new_P2_U3479;
  assign new_P2_U4893 = ~new_P2_U4892 | ~new_P2_U4891 | ~new_P2_U4890;
  assign new_P2_U4894 = ~new_P2_U3045 | ~new_P2_U4889;
  assign new_P2_U4895 = ~n2619 | ~new_P2_U4893;
  assign new_P2_U4896 = ~new_P2_R1170_U12 | ~new_P2_U3044;
  assign new_P2_U4897 = ~P2_REG3_REG_17_ | ~n2609;
  assign new_P2_U4898 = ~new_P2_U3042 | ~new_P2_U3479;
  assign new_P2_U4899 = ~new_P2_R1209_U12 | ~new_P2_U3040;
  assign new_P2_U4900 = ~P2_ADDR_REG_17_ | ~new_P2_U4863;
  assign new_P2_U4901 = ~new_P2_R1170_U76 | ~new_P2_U3043;
  assign new_P2_U4902 = ~new_P2_U3041 | ~new_P2_U3476;
  assign new_P2_U4903 = ~new_P2_R1209_U76 | ~new_P2_U3039;
  assign new_P2_U4904 = ~new_P2_U4903 | ~new_P2_U4902 | ~new_P2_U4901;
  assign new_P2_U4905 = ~new_P2_R1170_U76 | ~new_P2_U3018;
  assign new_P2_U4906 = ~new_P2_R1209_U76 | ~new_P2_U3017;
  assign new_P2_U4907 = ~new_P2_U5683 | ~new_P2_U3476;
  assign new_P2_U4908 = ~new_P2_U4907 | ~new_P2_U4906 | ~new_P2_U4905;
  assign new_P2_U4909 = ~new_P2_U3045 | ~new_P2_U4904;
  assign new_P2_U4910 = ~n2619 | ~new_P2_U4908;
  assign new_P2_U4911 = ~new_P2_R1170_U76 | ~new_P2_U3044;
  assign new_P2_U4912 = ~P2_REG3_REG_16_ | ~n2609;
  assign new_P2_U4913 = ~new_P2_U3042 | ~new_P2_U3476;
  assign new_P2_U4914 = ~new_P2_R1209_U76 | ~new_P2_U3040;
  assign new_P2_U4915 = ~P2_ADDR_REG_16_ | ~new_P2_U4863;
  assign new_P2_U4916 = ~new_P2_R1170_U77 | ~new_P2_U3043;
  assign new_P2_U4917 = ~new_P2_U3041 | ~new_P2_U3473;
  assign new_P2_U4918 = ~new_P2_R1209_U77 | ~new_P2_U3039;
  assign new_P2_U4919 = ~new_P2_U4918 | ~new_P2_U4917 | ~new_P2_U4916;
  assign new_P2_U4920 = ~new_P2_R1170_U77 | ~new_P2_U3018;
  assign new_P2_U4921 = ~new_P2_R1209_U77 | ~new_P2_U3017;
  assign new_P2_U4922 = ~new_P2_U5683 | ~new_P2_U3473;
  assign new_P2_U4923 = ~new_P2_U4922 | ~new_P2_U4921 | ~new_P2_U4920;
  assign new_P2_U4924 = ~new_P2_U3045 | ~new_P2_U4919;
  assign new_P2_U4925 = ~n2619 | ~new_P2_U4923;
  assign new_P2_U4926 = ~new_P2_R1170_U77 | ~new_P2_U3044;
  assign new_P2_U4927 = ~P2_REG3_REG_15_ | ~n2609;
  assign new_P2_U4928 = ~new_P2_U3042 | ~new_P2_U3473;
  assign new_P2_U4929 = ~new_P2_R1209_U77 | ~new_P2_U3040;
  assign new_P2_U4930 = ~P2_ADDR_REG_15_ | ~new_P2_U4863;
  assign new_P2_U4931 = ~new_P2_R1170_U78 | ~new_P2_U3043;
  assign new_P2_U4932 = ~new_P2_U3041 | ~new_P2_U3470;
  assign new_P2_U4933 = ~new_P2_R1209_U78 | ~new_P2_U3039;
  assign new_P2_U4934 = ~new_P2_U4933 | ~new_P2_U4932 | ~new_P2_U4931;
  assign new_P2_U4935 = ~new_P2_R1170_U78 | ~new_P2_U3018;
  assign new_P2_U4936 = ~new_P2_R1209_U78 | ~new_P2_U3017;
  assign new_P2_U4937 = ~new_P2_U5683 | ~new_P2_U3470;
  assign new_P2_U4938 = ~new_P2_U4937 | ~new_P2_U4936 | ~new_P2_U4935;
  assign new_P2_U4939 = ~new_P2_U3045 | ~new_P2_U4934;
  assign new_P2_U4940 = ~n2619 | ~new_P2_U4938;
  assign new_P2_U4941 = ~new_P2_R1170_U78 | ~new_P2_U3044;
  assign new_P2_U4942 = ~P2_REG3_REG_14_ | ~n2609;
  assign new_P2_U4943 = ~new_P2_U3042 | ~new_P2_U3470;
  assign new_P2_U4944 = ~new_P2_R1209_U78 | ~new_P2_U3040;
  assign new_P2_U4945 = ~P2_ADDR_REG_14_ | ~new_P2_U4863;
  assign new_P2_U4946 = ~new_P2_R1170_U11 | ~new_P2_U3043;
  assign new_P2_U4947 = ~new_P2_U3041 | ~new_P2_U3467;
  assign new_P2_U4948 = ~new_P2_R1209_U11 | ~new_P2_U3039;
  assign new_P2_U4949 = ~new_P2_U4948 | ~new_P2_U4947 | ~new_P2_U4946;
  assign new_P2_U4950 = ~new_P2_R1170_U11 | ~new_P2_U3018;
  assign new_P2_U4951 = ~new_P2_R1209_U11 | ~new_P2_U3017;
  assign new_P2_U4952 = ~new_P2_U5683 | ~new_P2_U3467;
  assign new_P2_U4953 = ~new_P2_U4952 | ~new_P2_U4951 | ~new_P2_U4950;
  assign new_P2_U4954 = ~new_P2_U3045 | ~new_P2_U4949;
  assign new_P2_U4955 = ~n2619 | ~new_P2_U4953;
  assign new_P2_U4956 = ~new_P2_R1170_U11 | ~new_P2_U3044;
  assign new_P2_U4957 = ~P2_REG3_REG_13_ | ~n2609;
  assign new_P2_U4958 = ~new_P2_U3042 | ~new_P2_U3467;
  assign new_P2_U4959 = ~new_P2_R1209_U11 | ~new_P2_U3040;
  assign new_P2_U4960 = ~P2_ADDR_REG_13_ | ~new_P2_U4863;
  assign new_P2_U4961 = ~new_P2_R1170_U79 | ~new_P2_U3043;
  assign new_P2_U4962 = ~new_P2_U3041 | ~new_P2_U3464;
  assign new_P2_U4963 = ~new_P2_R1209_U79 | ~new_P2_U3039;
  assign new_P2_U4964 = ~new_P2_U4963 | ~new_P2_U4962 | ~new_P2_U4961;
  assign new_P2_U4965 = ~new_P2_R1170_U79 | ~new_P2_U3018;
  assign new_P2_U4966 = ~new_P2_R1209_U79 | ~new_P2_U3017;
  assign new_P2_U4967 = ~new_P2_U5683 | ~new_P2_U3464;
  assign new_P2_U4968 = ~new_P2_U4967 | ~new_P2_U4966 | ~new_P2_U4965;
  assign new_P2_U4969 = ~new_P2_U3045 | ~new_P2_U4964;
  assign new_P2_U4970 = ~n2619 | ~new_P2_U4968;
  assign new_P2_U4971 = ~new_P2_R1170_U79 | ~new_P2_U3044;
  assign new_P2_U4972 = ~P2_REG3_REG_12_ | ~n2609;
  assign new_P2_U4973 = ~new_P2_U3042 | ~new_P2_U3464;
  assign new_P2_U4974 = ~new_P2_R1209_U79 | ~new_P2_U3040;
  assign new_P2_U4975 = ~P2_ADDR_REG_12_ | ~new_P2_U4863;
  assign new_P2_U4976 = ~new_P2_R1170_U80 | ~new_P2_U3043;
  assign new_P2_U4977 = ~new_P2_U3041 | ~new_P2_U3461;
  assign new_P2_U4978 = ~new_P2_R1209_U80 | ~new_P2_U3039;
  assign new_P2_U4979 = ~new_P2_U4978 | ~new_P2_U4977 | ~new_P2_U4976;
  assign new_P2_U4980 = ~new_P2_R1170_U80 | ~new_P2_U3018;
  assign new_P2_U4981 = ~new_P2_R1209_U80 | ~new_P2_U3017;
  assign new_P2_U4982 = ~new_P2_U5683 | ~new_P2_U3461;
  assign new_P2_U4983 = ~new_P2_U4982 | ~new_P2_U4981 | ~new_P2_U4980;
  assign new_P2_U4984 = ~new_P2_U3045 | ~new_P2_U4979;
  assign new_P2_U4985 = ~n2619 | ~new_P2_U4983;
  assign new_P2_U4986 = ~new_P2_R1170_U80 | ~new_P2_U3044;
  assign new_P2_U4987 = ~P2_REG3_REG_11_ | ~n2609;
  assign new_P2_U4988 = ~new_P2_U3042 | ~new_P2_U3461;
  assign new_P2_U4989 = ~new_P2_R1209_U80 | ~new_P2_U3040;
  assign new_P2_U4990 = ~P2_ADDR_REG_11_ | ~new_P2_U4863;
  assign new_P2_U4991 = ~new_P2_R1170_U10 | ~new_P2_U3043;
  assign new_P2_U4992 = ~new_P2_U3041 | ~new_P2_U3458;
  assign new_P2_U4993 = ~new_P2_R1209_U10 | ~new_P2_U3039;
  assign new_P2_U4994 = ~new_P2_U4993 | ~new_P2_U4992 | ~new_P2_U4991;
  assign new_P2_U4995 = ~new_P2_R1170_U10 | ~new_P2_U3018;
  assign new_P2_U4996 = ~new_P2_R1209_U10 | ~new_P2_U3017;
  assign new_P2_U4997 = ~new_P2_U5683 | ~new_P2_U3458;
  assign new_P2_U4998 = ~new_P2_U4997 | ~new_P2_U4996 | ~new_P2_U4995;
  assign new_P2_U4999 = ~new_P2_U3045 | ~new_P2_U4994;
  assign new_P2_U5000 = ~n2619 | ~new_P2_U4998;
  assign new_P2_U5001 = ~new_P2_R1170_U10 | ~new_P2_U3044;
  assign new_P2_U5002 = ~P2_REG3_REG_10_ | ~n2609;
  assign new_P2_U5003 = ~new_P2_U3042 | ~new_P2_U3458;
  assign new_P2_U5004 = ~new_P2_R1209_U10 | ~new_P2_U3040;
  assign new_P2_U5005 = ~P2_ADDR_REG_10_ | ~new_P2_U4863;
  assign new_P2_U5006 = ~new_P2_R1170_U70 | ~new_P2_U3043;
  assign new_P2_U5007 = ~new_P2_U3041 | ~new_P2_U3455;
  assign new_P2_U5008 = ~new_P2_R1209_U70 | ~new_P2_U3039;
  assign new_P2_U5009 = ~new_P2_U5008 | ~new_P2_U5007 | ~new_P2_U5006;
  assign new_P2_U5010 = ~new_P2_R1170_U70 | ~new_P2_U3018;
  assign new_P2_U5011 = ~new_P2_R1209_U70 | ~new_P2_U3017;
  assign new_P2_U5012 = ~new_P2_U5683 | ~new_P2_U3455;
  assign new_P2_U5013 = ~new_P2_U5012 | ~new_P2_U5011 | ~new_P2_U5010;
  assign new_P2_U5014 = ~new_P2_U3045 | ~new_P2_U5009;
  assign new_P2_U5015 = ~n2619 | ~new_P2_U5013;
  assign new_P2_U5016 = ~new_P2_R1170_U70 | ~new_P2_U3044;
  assign new_P2_U5017 = ~P2_REG3_REG_9_ | ~n2609;
  assign new_P2_U5018 = ~new_P2_U3042 | ~new_P2_U3455;
  assign new_P2_U5019 = ~new_P2_R1209_U70 | ~new_P2_U3040;
  assign new_P2_U5020 = ~P2_ADDR_REG_9_ | ~new_P2_U4863;
  assign new_P2_U5021 = ~new_P2_R1170_U71 | ~new_P2_U3043;
  assign new_P2_U5022 = ~new_P2_U3041 | ~new_P2_U3452;
  assign new_P2_U5023 = ~new_P2_R1209_U71 | ~new_P2_U3039;
  assign new_P2_U5024 = ~new_P2_U5023 | ~new_P2_U5022 | ~new_P2_U5021;
  assign new_P2_U5025 = ~new_P2_R1170_U71 | ~new_P2_U3018;
  assign new_P2_U5026 = ~new_P2_R1209_U71 | ~new_P2_U3017;
  assign new_P2_U5027 = ~new_P2_U5683 | ~new_P2_U3452;
  assign new_P2_U5028 = ~new_P2_U5027 | ~new_P2_U5026 | ~new_P2_U5025;
  assign new_P2_U5029 = ~new_P2_U3045 | ~new_P2_U5024;
  assign new_P2_U5030 = ~n2619 | ~new_P2_U5028;
  assign new_P2_U5031 = ~new_P2_R1170_U71 | ~new_P2_U3044;
  assign new_P2_U5032 = ~P2_REG3_REG_8_ | ~n2609;
  assign new_P2_U5033 = ~new_P2_U3042 | ~new_P2_U3452;
  assign new_P2_U5034 = ~new_P2_R1209_U71 | ~new_P2_U3040;
  assign new_P2_U5035 = ~P2_ADDR_REG_8_ | ~new_P2_U4863;
  assign new_P2_U5036 = ~new_P2_R1170_U16 | ~new_P2_U3043;
  assign new_P2_U5037 = ~new_P2_U3041 | ~new_P2_U3449;
  assign new_P2_U5038 = ~new_P2_R1209_U16 | ~new_P2_U3039;
  assign new_P2_U5039 = ~new_P2_U5038 | ~new_P2_U5037 | ~new_P2_U5036;
  assign new_P2_U5040 = ~new_P2_R1170_U16 | ~new_P2_U3018;
  assign new_P2_U5041 = ~new_P2_R1209_U16 | ~new_P2_U3017;
  assign new_P2_U5042 = ~new_P2_U5683 | ~new_P2_U3449;
  assign new_P2_U5043 = ~new_P2_U5042 | ~new_P2_U5041 | ~new_P2_U5040;
  assign new_P2_U5044 = ~new_P2_U3045 | ~new_P2_U5039;
  assign new_P2_U5045 = ~n2619 | ~new_P2_U5043;
  assign new_P2_U5046 = ~new_P2_R1170_U16 | ~new_P2_U3044;
  assign new_P2_U5047 = ~P2_REG3_REG_7_ | ~n2609;
  assign new_P2_U5048 = ~new_P2_U3042 | ~new_P2_U3449;
  assign new_P2_U5049 = ~new_P2_R1209_U16 | ~new_P2_U3040;
  assign new_P2_U5050 = ~P2_ADDR_REG_7_ | ~new_P2_U4863;
  assign new_P2_U5051 = ~new_P2_R1170_U72 | ~new_P2_U3043;
  assign new_P2_U5052 = ~new_P2_U3041 | ~new_P2_U3446;
  assign new_P2_U5053 = ~new_P2_R1209_U72 | ~new_P2_U3039;
  assign new_P2_U5054 = ~new_P2_U5053 | ~new_P2_U5052 | ~new_P2_U5051;
  assign new_P2_U5055 = ~new_P2_R1170_U72 | ~new_P2_U3018;
  assign new_P2_U5056 = ~new_P2_R1209_U72 | ~new_P2_U3017;
  assign new_P2_U5057 = ~new_P2_U5683 | ~new_P2_U3446;
  assign new_P2_U5058 = ~new_P2_U5057 | ~new_P2_U5056 | ~new_P2_U5055;
  assign new_P2_U5059 = ~new_P2_U3045 | ~new_P2_U5054;
  assign new_P2_U5060 = ~n2619 | ~new_P2_U5058;
  assign new_P2_U5061 = ~new_P2_R1170_U72 | ~new_P2_U3044;
  assign new_P2_U5062 = ~P2_REG3_REG_6_ | ~n2609;
  assign new_P2_U5063 = ~new_P2_U3042 | ~new_P2_U3446;
  assign new_P2_U5064 = ~new_P2_R1209_U72 | ~new_P2_U3040;
  assign new_P2_U5065 = ~P2_ADDR_REG_6_ | ~new_P2_U4863;
  assign new_P2_U5066 = ~new_P2_R1170_U15 | ~new_P2_U3043;
  assign new_P2_U5067 = ~new_P2_U3041 | ~new_P2_U3443;
  assign new_P2_U5068 = ~new_P2_R1209_U15 | ~new_P2_U3039;
  assign new_P2_U5069 = ~new_P2_U5068 | ~new_P2_U5067 | ~new_P2_U5066;
  assign new_P2_U5070 = ~new_P2_R1170_U15 | ~new_P2_U3018;
  assign new_P2_U5071 = ~new_P2_R1209_U15 | ~new_P2_U3017;
  assign new_P2_U5072 = ~new_P2_U5683 | ~new_P2_U3443;
  assign new_P2_U5073 = ~new_P2_U5072 | ~new_P2_U5071 | ~new_P2_U5070;
  assign new_P2_U5074 = ~new_P2_U3045 | ~new_P2_U5069;
  assign new_P2_U5075 = ~n2619 | ~new_P2_U5073;
  assign new_P2_U5076 = ~new_P2_R1170_U15 | ~new_P2_U3044;
  assign new_P2_U5077 = ~P2_REG3_REG_5_ | ~n2609;
  assign new_P2_U5078 = ~new_P2_U3042 | ~new_P2_U3443;
  assign new_P2_U5079 = ~new_P2_R1209_U15 | ~new_P2_U3040;
  assign new_P2_U5080 = ~P2_ADDR_REG_5_ | ~new_P2_U4863;
  assign new_P2_U5081 = ~new_P2_R1170_U73 | ~new_P2_U3043;
  assign new_P2_U5082 = ~new_P2_U3041 | ~new_P2_U3440;
  assign new_P2_U5083 = ~new_P2_R1209_U73 | ~new_P2_U3039;
  assign new_P2_U5084 = ~new_P2_U5083 | ~new_P2_U5082 | ~new_P2_U5081;
  assign new_P2_U5085 = ~new_P2_R1170_U73 | ~new_P2_U3018;
  assign new_P2_U5086 = ~new_P2_R1209_U73 | ~new_P2_U3017;
  assign new_P2_U5087 = ~new_P2_U5683 | ~new_P2_U3440;
  assign new_P2_U5088 = ~new_P2_U5087 | ~new_P2_U5086 | ~new_P2_U5085;
  assign new_P2_U5089 = ~new_P2_U3045 | ~new_P2_U5084;
  assign new_P2_U5090 = ~n2619 | ~new_P2_U5088;
  assign new_P2_U5091 = ~new_P2_R1170_U73 | ~new_P2_U3044;
  assign new_P2_U5092 = ~P2_REG3_REG_4_ | ~n2609;
  assign new_P2_U5093 = ~new_P2_U3042 | ~new_P2_U3440;
  assign new_P2_U5094 = ~new_P2_R1209_U73 | ~new_P2_U3040;
  assign new_P2_U5095 = ~P2_ADDR_REG_4_ | ~new_P2_U4863;
  assign new_P2_U5096 = ~new_P2_R1170_U74 | ~new_P2_U3043;
  assign new_P2_U5097 = ~new_P2_U3041 | ~new_P2_U3437;
  assign new_P2_U5098 = ~new_P2_R1209_U74 | ~new_P2_U3039;
  assign new_P2_U5099 = ~new_P2_U5098 | ~new_P2_U5097 | ~new_P2_U5096;
  assign new_P2_U5100 = ~new_P2_R1170_U74 | ~new_P2_U3018;
  assign new_P2_U5101 = ~new_P2_R1209_U74 | ~new_P2_U3017;
  assign new_P2_U5102 = ~new_P2_U5683 | ~new_P2_U3437;
  assign new_P2_U5103 = ~new_P2_U5102 | ~new_P2_U5101 | ~new_P2_U5100;
  assign new_P2_U5104 = ~new_P2_U3045 | ~new_P2_U5099;
  assign new_P2_U5105 = ~n2619 | ~new_P2_U5103;
  assign new_P2_U5106 = ~new_P2_R1170_U74 | ~new_P2_U3044;
  assign new_P2_U5107 = ~P2_REG3_REG_3_ | ~n2609;
  assign new_P2_U5108 = ~new_P2_U3042 | ~new_P2_U3437;
  assign new_P2_U5109 = ~new_P2_R1209_U74 | ~new_P2_U3040;
  assign new_P2_U5110 = ~P2_ADDR_REG_3_ | ~new_P2_U4863;
  assign new_P2_U5111 = ~new_P2_R1170_U14 | ~new_P2_U3043;
  assign new_P2_U5112 = ~new_P2_U3041 | ~new_P2_U3434;
  assign new_P2_U5113 = ~new_P2_R1209_U14 | ~new_P2_U3039;
  assign new_P2_U5114 = ~new_P2_U5113 | ~new_P2_U5112 | ~new_P2_U5111;
  assign new_P2_U5115 = ~new_P2_R1170_U14 | ~new_P2_U3018;
  assign new_P2_U5116 = ~new_P2_R1209_U14 | ~new_P2_U3017;
  assign new_P2_U5117 = ~new_P2_U5683 | ~new_P2_U3434;
  assign new_P2_U5118 = ~new_P2_U5117 | ~new_P2_U5116 | ~new_P2_U5115;
  assign new_P2_U5119 = ~new_P2_U3045 | ~new_P2_U5114;
  assign new_P2_U5120 = ~n2619 | ~new_P2_U5118;
  assign new_P2_U5121 = ~new_P2_R1170_U14 | ~new_P2_U3044;
  assign new_P2_U5122 = ~P2_REG3_REG_2_ | ~n2609;
  assign new_P2_U5123 = ~new_P2_U3042 | ~new_P2_U3434;
  assign new_P2_U5124 = ~new_P2_R1209_U14 | ~new_P2_U3040;
  assign new_P2_U5125 = ~P2_ADDR_REG_2_ | ~new_P2_U4863;
  assign new_P2_U5126 = ~new_P2_R1170_U68 | ~new_P2_U3043;
  assign new_P2_U5127 = ~new_P2_U3041 | ~new_P2_U3431;
  assign new_P2_U5128 = ~new_P2_R1209_U68 | ~new_P2_U3039;
  assign new_P2_U5129 = ~new_P2_U5128 | ~new_P2_U5127 | ~new_P2_U5126;
  assign new_P2_U5130 = ~new_P2_R1170_U68 | ~new_P2_U3018;
  assign new_P2_U5131 = ~new_P2_R1209_U68 | ~new_P2_U3017;
  assign new_P2_U5132 = ~new_P2_U5683 | ~new_P2_U3431;
  assign new_P2_U5133 = ~new_P2_U5132 | ~new_P2_U5131 | ~new_P2_U5130;
  assign new_P2_U5134 = ~new_P2_U3045 | ~new_P2_U5129;
  assign new_P2_U5135 = ~n2619 | ~new_P2_U5133;
  assign new_P2_U5136 = ~new_P2_R1170_U68 | ~new_P2_U3044;
  assign new_P2_U5137 = ~P2_REG3_REG_1_ | ~n2609;
  assign new_P2_U5138 = ~new_P2_U3042 | ~new_P2_U3431;
  assign new_P2_U5139 = ~new_P2_R1209_U68 | ~new_P2_U3040;
  assign new_P2_U5140 = ~P2_ADDR_REG_1_ | ~new_P2_U4863;
  assign new_P2_U5141 = ~new_P2_R1170_U69 | ~new_P2_U3043;
  assign new_P2_U5142 = ~new_P2_U3041 | ~new_P2_U3425;
  assign new_P2_U5143 = ~new_P2_R1209_U69 | ~new_P2_U3039;
  assign new_P2_U5144 = ~new_P2_U5143 | ~new_P2_U5142 | ~new_P2_U5141;
  assign new_P2_U5145 = ~new_P2_R1170_U69 | ~new_P2_U3018;
  assign new_P2_U5146 = ~new_P2_R1209_U69 | ~new_P2_U3017;
  assign new_P2_U5147 = ~new_P2_U5683 | ~new_P2_U3425;
  assign new_P2_U5148 = ~new_P2_U5147 | ~new_P2_U5146 | ~new_P2_U5145;
  assign new_P2_U5149 = ~new_P2_U3045 | ~new_P2_U5144;
  assign new_P2_U5150 = ~n2619 | ~new_P2_U5148;
  assign new_P2_U5151 = ~new_P2_R1170_U69 | ~new_P2_U3044;
  assign new_P2_U5152 = ~P2_REG3_REG_0_ | ~n2609;
  assign new_P2_U5153 = ~new_P2_U3042 | ~new_P2_U3425;
  assign new_P2_U5154 = ~new_P2_R1209_U69 | ~new_P2_U3040;
  assign new_P2_U5155 = ~P2_ADDR_REG_0_ | ~new_P2_U4863;
  assign new_P2_U5156 = ~new_P2_U3918;
  assign new_P2_U5157 = ~new_P2_U3337 | ~new_P2_U3936 | ~new_P2_U3334;
  assign new_P2_U5158 = ~new_P2_U5665 | ~new_P2_U5671;
  assign new_P2_U5159 = ~new_P2_U3424 | ~new_P2_U5158;
  assign new_P2_U5160 = ~new_P2_U3419 | ~new_P2_U5159;
  assign new_P2_U5161 = ~new_P2_U3340 | ~new_P2_U5160;
  assign new_P2_U5162 = ~new_P2_U3052 | ~new_P2_U6052 | ~new_P2_U6051;
  assign new_P2_U5163 = ~P2_B_REG | ~new_P2_U5162;
  assign new_P2_U5164 = ~new_P2_U3038 | ~new_P2_U3081;
  assign new_P2_U5165 = ~new_P2_U3036 | ~new_P2_U3075;
  assign new_P2_U5166 = ~new_P2_ADD_1119_U69 | ~new_P2_U3406;
  assign new_P2_U5167 = ~new_P2_U5166 | ~new_P2_U5165 | ~new_P2_U5164;
  assign new_P2_U5168 = ~new_P2_U3154;
  assign new_P2_U5169 = ~new_P2_U3923 | ~new_P2_U3346;
  assign new_P2_U5170 = ~new_P2_U3419 | ~new_P2_U5169;
  assign new_P2_U5171 = ~new_P2_U3801 | ~new_P2_U3800 | ~new_P2_U5170;
  assign new_P2_U5172 = ~new_P2_U5171 | ~new_P2_U3406;
  assign new_P2_U5173 = ~new_P2_U3408;
  assign new_P2_U5174 = ~new_P2_U3474 | ~new_P2_U5636;
  assign new_P2_U5175 = ~new_P2_ADD_1119_U69 | ~new_P2_U5635;
  assign new_P2_U5176 = ~new_P2_R1176_U111 | ~new_P2_U3028;
  assign new_P2_U5177 = ~new_P2_U3969 | ~new_P2_U5167;
  assign new_P2_U5178 = ~P2_REG3_REG_15_ | ~n2609;
  assign new_P2_U5179 = ~new_P2_U3038 | ~new_P2_U3060;
  assign new_P2_U5180 = ~new_P2_U3036 | ~new_P2_U3055;
  assign new_P2_U5181 = ~new_P2_ADD_1119_U58 | ~new_P2_U3406;
  assign new_P2_U5182 = ~new_P2_U5180 | ~new_P2_U5181 | ~new_P2_U5179;
  assign new_P2_U5183 = ~new_P2_U3398 | ~new_P2_U3406;
  assign new_P2_U5184 = ~new_P2_U5173 | ~new_P2_U5183;
  assign new_P2_U5185 = ~new_P2_U3946 | ~new_P2_U3398;
  assign new_P2_U5186 = ~new_P2_U3393 | ~new_P2_U5185;
  assign new_P2_U5187 = ~new_P2_U3047 | ~new_P2_U3951;
  assign new_P2_U5188 = ~new_P2_U3046 | ~new_P2_ADD_1119_U58;
  assign new_P2_U5189 = ~new_P2_R1176_U16 | ~new_P2_U3028;
  assign new_P2_U5190 = ~new_P2_U3969 | ~new_P2_U5182;
  assign new_P2_U5191 = ~P2_REG3_REG_26_ | ~n2609;
  assign new_P2_U5192 = ~new_P2_U3038 | ~new_P2_U3069;
  assign new_P2_U5193 = ~new_P2_U3036 | ~new_P2_U3072;
  assign new_P2_U5194 = ~new_P2_ADD_1119_U53 | ~new_P2_U3406;
  assign new_P2_U5195 = ~new_P2_U5194 | ~new_P2_U5193 | ~new_P2_U5192;
  assign new_P2_U5196 = ~new_P2_U3447 | ~new_P2_U5636;
  assign new_P2_U5197 = ~new_P2_ADD_1119_U53 | ~new_P2_U5635;
  assign new_P2_U5198 = ~new_P2_R1176_U96 | ~new_P2_U3028;
  assign new_P2_U5199 = ~new_P2_U3969 | ~new_P2_U5195;
  assign new_P2_U5200 = ~P2_REG3_REG_6_ | ~n2609;
  assign new_P2_U5201 = ~new_P2_U3038 | ~new_P2_U3071;
  assign new_P2_U5202 = ~new_P2_U3036 | ~new_P2_U3083;
  assign new_P2_U5203 = ~new_P2_ADD_1119_U66 | ~new_P2_U3406;
  assign new_P2_U5204 = ~new_P2_U5203 | ~new_P2_U5202 | ~new_P2_U5201;
  assign new_P2_U5205 = ~new_P2_U3483 | ~new_P2_U5636;
  assign new_P2_U5206 = ~new_P2_ADD_1119_U66 | ~new_P2_U5635;
  assign new_P2_U5207 = ~new_P2_R1176_U109 | ~new_P2_U3028;
  assign new_P2_U5208 = ~new_P2_U3969 | ~new_P2_U5204;
  assign new_P2_U5209 = ~P2_REG3_REG_18_ | ~n2609;
  assign new_P2_U5210 = ~new_P2_U3038 | ~new_P2_U3080;
  assign new_P2_U5211 = ~new_P2_U3036 | ~new_P2_U3066;
  assign new_P2_U5212 = ~P2_REG3_REG_2_ | ~new_P2_U3406;
  assign new_P2_U5213 = ~new_P2_U5212 | ~new_P2_U5211 | ~new_P2_U5210;
  assign new_P2_U5214 = ~new_P2_U3435 | ~new_P2_U5636;
  assign new_P2_U5215 = ~P2_REG3_REG_2_ | ~new_P2_U5635;
  assign new_P2_U5216 = ~new_P2_R1176_U99 | ~new_P2_U3028;
  assign new_P2_U5217 = ~new_P2_U3969 | ~new_P2_U5213;
  assign new_P2_U5218 = ~P2_REG3_REG_2_ | ~n2609;
  assign new_P2_U5219 = ~new_P2_U3038 | ~new_P2_U3064;
  assign new_P2_U5220 = ~new_P2_U3036 | ~new_P2_U3074;
  assign new_P2_U5221 = ~new_P2_ADD_1119_U73 | ~new_P2_U3406;
  assign new_P2_U5222 = ~new_P2_U5221 | ~new_P2_U5220 | ~new_P2_U5219;
  assign new_P2_U5223 = ~new_P2_U3462 | ~new_P2_U5636;
  assign new_P2_U5224 = ~new_P2_ADD_1119_U73 | ~new_P2_U5635;
  assign new_P2_U5225 = ~new_P2_R1176_U114 | ~new_P2_U3028;
  assign new_P2_U5226 = ~new_P2_U3969 | ~new_P2_U5222;
  assign new_P2_U5227 = ~P2_REG3_REG_11_ | ~n2609;
  assign new_P2_U5228 = ~new_P2_U3038 | ~new_P2_U3077;
  assign new_P2_U5229 = ~new_P2_U3036 | ~new_P2_U3068;
  assign new_P2_U5230 = ~new_P2_ADD_1119_U62 | ~new_P2_U3406;
  assign new_P2_U5231 = ~new_P2_U5230 | ~new_P2_U5229 | ~new_P2_U5228;
  assign new_P2_U5232 = ~new_P2_U3047 | ~new_P2_U3955;
  assign new_P2_U5233 = ~new_P2_U3046 | ~new_P2_ADD_1119_U62;
  assign new_P2_U5234 = ~new_P2_R1176_U105 | ~new_P2_U3028;
  assign new_P2_U5235 = ~new_P2_U3969 | ~new_P2_U5231;
  assign new_P2_U5236 = ~P2_REG3_REG_22_ | ~n2609;
  assign new_P2_U5237 = ~new_P2_U3038 | ~new_P2_U3074;
  assign new_P2_U5238 = ~new_P2_U3036 | ~new_P2_U3081;
  assign new_P2_U5239 = ~new_P2_ADD_1119_U71 | ~new_P2_U3406;
  assign new_P2_U5240 = ~new_P2_U5239 | ~new_P2_U5238 | ~new_P2_U5237;
  assign new_P2_U5241 = ~new_P2_U3468 | ~new_P2_U5636;
  assign new_P2_U5242 = ~new_P2_ADD_1119_U71 | ~new_P2_U5635;
  assign new_P2_U5243 = ~new_P2_R1176_U13 | ~new_P2_U3028;
  assign new_P2_U5244 = ~new_P2_U3969 | ~new_P2_U5240;
  assign new_P2_U5245 = ~P2_REG3_REG_13_ | ~n2609;
  assign new_P2_U5246 = ~new_P2_U3038 | ~new_P2_U3083;
  assign new_P2_U5247 = ~new_P2_U3036 | ~new_P2_U3077;
  assign new_P2_U5248 = ~new_P2_ADD_1119_U64 | ~new_P2_U3406;
  assign new_P2_U5249 = ~new_P2_U5248 | ~new_P2_U5247 | ~new_P2_U5246;
  assign new_P2_U5250 = ~new_P2_U3047 | ~new_P2_U3957;
  assign new_P2_U5251 = ~new_P2_U3046 | ~new_P2_ADD_1119_U64;
  assign new_P2_U5252 = ~new_P2_R1176_U106 | ~new_P2_U3028;
  assign new_P2_U5253 = ~new_P2_U3969 | ~new_P2_U5249;
  assign new_P2_U5254 = ~P2_REG3_REG_20_ | ~n2609;
  assign new_P2_U5255 = ~new_P2_U3407 | ~new_P2_U3405;
  assign new_P2_U5256 = ~new_P2_U5255 | ~new_P2_U3406;
  assign new_P2_U5257 = ~new_P2_U3970 | ~new_P2_U5256;
  assign new_P2_U5258 = ~new_P2_U3806 | ~new_P2_U3036;
  assign new_P2_U5259 = ~new_P2_U3427 | ~new_P2_U5636;
  assign new_P2_U5260 = ~P2_REG3_REG_0_ | ~new_P2_U5257;
  assign new_P2_U5261 = ~new_P2_R1176_U93 | ~new_P2_U3028;
  assign new_P2_U5262 = ~P2_REG3_REG_0_ | ~n2609;
  assign new_P2_U5263 = ~new_P2_U3038 | ~new_P2_U3086;
  assign new_P2_U5264 = ~new_P2_U3036 | ~new_P2_U3064;
  assign new_P2_U5265 = ~new_P2_ADD_1119_U50 | ~new_P2_U3406;
  assign new_P2_U5266 = ~new_P2_U5265 | ~new_P2_U5264 | ~new_P2_U5263;
  assign new_P2_U5267 = ~new_P2_U3456 | ~new_P2_U5636;
  assign new_P2_U5268 = ~new_P2_ADD_1119_U50 | ~new_P2_U5635;
  assign new_P2_U5269 = ~new_P2_R1176_U94 | ~new_P2_U3028;
  assign new_P2_U5270 = ~new_P2_U3969 | ~new_P2_U5266;
  assign new_P2_U5271 = ~P2_REG3_REG_9_ | ~n2609;
  assign new_P2_U5272 = ~new_P2_U3038 | ~new_P2_U3066;
  assign new_P2_U5273 = ~new_P2_U3036 | ~new_P2_U3069;
  assign new_P2_U5274 = ~new_P2_ADD_1119_U55 | ~new_P2_U3406;
  assign new_P2_U5275 = ~new_P2_U5274 | ~new_P2_U5273 | ~new_P2_U5272;
  assign new_P2_U5276 = ~new_P2_U3441 | ~new_P2_U5636;
  assign new_P2_U5277 = ~new_P2_ADD_1119_U55 | ~new_P2_U5635;
  assign new_P2_U5278 = ~new_P2_R1176_U98 | ~new_P2_U3028;
  assign new_P2_U5279 = ~new_P2_U3969 | ~new_P2_U5275;
  assign new_P2_U5280 = ~P2_REG3_REG_4_ | ~n2609;
  assign new_P2_U5281 = ~new_P2_U3038 | ~new_P2_U3068;
  assign new_P2_U5282 = ~new_P2_U3036 | ~new_P2_U3060;
  assign new_P2_U5283 = ~new_P2_ADD_1119_U60 | ~new_P2_U3406;
  assign new_P2_U5284 = ~new_P2_U5283 | ~new_P2_U5282 | ~new_P2_U5281;
  assign new_P2_U5285 = ~new_P2_U3047 | ~new_P2_U3953;
  assign new_P2_U5286 = ~new_P2_U3046 | ~new_P2_ADD_1119_U60;
  assign new_P2_U5287 = ~new_P2_R1176_U103 | ~new_P2_U3028;
  assign new_P2_U5288 = ~new_P2_U3969 | ~new_P2_U5284;
  assign new_P2_U5289 = ~P2_REG3_REG_24_ | ~n2609;
  assign new_P2_U5290 = ~new_P2_U3038 | ~new_P2_U3075;
  assign new_P2_U5291 = ~new_P2_U3036 | ~new_P2_U3084;
  assign new_P2_U5292 = ~new_P2_ADD_1119_U67 | ~new_P2_U3406;
  assign new_P2_U5293 = ~new_P2_U5292 | ~new_P2_U5291 | ~new_P2_U5290;
  assign new_P2_U5294 = ~new_P2_U3480 | ~new_P2_U5636;
  assign new_P2_U5295 = ~new_P2_ADD_1119_U67 | ~new_P2_U5635;
  assign new_P2_U5296 = ~new_P2_R1176_U14 | ~new_P2_U3028;
  assign new_P2_U5297 = ~new_P2_U3969 | ~new_P2_U5293;
  assign new_P2_U5298 = ~P2_REG3_REG_17_ | ~n2609;
  assign new_P2_U5299 = ~new_P2_U3038 | ~new_P2_U3062;
  assign new_P2_U5300 = ~new_P2_U3036 | ~new_P2_U3073;
  assign new_P2_U5301 = ~new_P2_ADD_1119_U54 | ~new_P2_U3406;
  assign new_P2_U5302 = ~new_P2_U5301 | ~new_P2_U5300 | ~new_P2_U5299;
  assign new_P2_U5303 = ~new_P2_U3444 | ~new_P2_U5636;
  assign new_P2_U5304 = ~new_P2_ADD_1119_U54 | ~new_P2_U5635;
  assign new_P2_U5305 = ~new_P2_R1176_U97 | ~new_P2_U3028;
  assign new_P2_U5306 = ~new_P2_U3969 | ~new_P2_U5302;
  assign new_P2_U5307 = ~P2_REG3_REG_5_ | ~n2609;
  assign new_P2_U5308 = ~new_P2_U3038 | ~new_P2_U3076;
  assign new_P2_U5309 = ~new_P2_U3036 | ~new_P2_U3071;
  assign new_P2_U5310 = ~new_P2_ADD_1119_U68 | ~new_P2_U3406;
  assign new_P2_U5311 = ~new_P2_U5310 | ~new_P2_U5309 | ~new_P2_U5308;
  assign new_P2_U5312 = ~new_P2_U3477 | ~new_P2_U5636;
  assign new_P2_U5313 = ~new_P2_ADD_1119_U68 | ~new_P2_U5635;
  assign new_P2_U5314 = ~new_P2_R1176_U110 | ~new_P2_U3028;
  assign new_P2_U5315 = ~new_P2_U3969 | ~new_P2_U5311;
  assign new_P2_U5316 = ~P2_REG3_REG_16_ | ~n2609;
  assign new_P2_U5317 = ~new_P2_U3038 | ~new_P2_U3067;
  assign new_P2_U5318 = ~new_P2_U3036 | ~new_P2_U3059;
  assign new_P2_U5319 = ~new_P2_ADD_1119_U59 | ~new_P2_U3406;
  assign new_P2_U5320 = ~new_P2_U5319 | ~new_P2_U5318 | ~new_P2_U5317;
  assign new_P2_U5321 = ~new_P2_U3047 | ~new_P2_U3952;
  assign new_P2_U5322 = ~new_P2_U3046 | ~new_P2_ADD_1119_U59;
  assign new_P2_U5323 = ~new_P2_R1176_U102 | ~new_P2_U3028;
  assign new_P2_U5324 = ~new_P2_U3969 | ~new_P2_U5320;
  assign new_P2_U5325 = ~P2_REG3_REG_25_ | ~n2609;
  assign new_P2_U5326 = ~new_P2_U3038 | ~new_P2_U3065;
  assign new_P2_U5327 = ~new_P2_U3036 | ~new_P2_U3082;
  assign new_P2_U5328 = ~new_P2_ADD_1119_U72 | ~new_P2_U3406;
  assign new_P2_U5329 = ~new_P2_U5328 | ~new_P2_U5327 | ~new_P2_U5326;
  assign new_P2_U5330 = ~new_P2_U3465 | ~new_P2_U5636;
  assign new_P2_U5331 = ~new_P2_ADD_1119_U72 | ~new_P2_U5635;
  assign new_P2_U5332 = ~new_P2_R1176_U113 | ~new_P2_U3028;
  assign new_P2_U5333 = ~new_P2_U3969 | ~new_P2_U5329;
  assign new_P2_U5334 = ~P2_REG3_REG_12_ | ~n2609;
  assign new_P2_U5335 = ~new_P2_U3038 | ~new_P2_U3078;
  assign new_P2_U5336 = ~new_P2_U3036 | ~new_P2_U3063;
  assign new_P2_U5337 = ~new_P2_ADD_1119_U63 | ~new_P2_U3406;
  assign new_P2_U5338 = ~new_P2_U5337 | ~new_P2_U5336 | ~new_P2_U5335;
  assign new_P2_U5339 = ~new_P2_U3047 | ~new_P2_U3956;
  assign new_P2_U5340 = ~new_P2_U3046 | ~new_P2_ADD_1119_U63;
  assign new_P2_U5341 = ~new_P2_R1176_U15 | ~new_P2_U3028;
  assign new_P2_U5342 = ~new_P2_U3969 | ~new_P2_U5338;
  assign new_P2_U5343 = ~P2_REG3_REG_21_ | ~n2609;
  assign new_P2_U5344 = ~new_P2_U3038 | ~new_P2_U3079;
  assign new_P2_U5345 = ~new_P2_U3036 | ~new_P2_U3070;
  assign new_P2_U5346 = ~P2_REG3_REG_1_ | ~new_P2_U3406;
  assign new_P2_U5347 = ~new_P2_U5346 | ~new_P2_U5345 | ~new_P2_U5344;
  assign new_P2_U5348 = ~new_P2_U3432 | ~new_P2_U5636;
  assign new_P2_U5349 = ~P2_REG3_REG_1_ | ~new_P2_U5635;
  assign new_P2_U5350 = ~new_P2_R1176_U107 | ~new_P2_U3028;
  assign new_P2_U5351 = ~new_P2_U3969 | ~new_P2_U5347;
  assign new_P2_U5352 = ~P2_REG3_REG_1_ | ~n2609;
  assign new_P2_U5353 = ~new_P2_U3038 | ~new_P2_U3072;
  assign new_P2_U5354 = ~new_P2_U3036 | ~new_P2_U3085;
  assign new_P2_U5355 = ~new_P2_ADD_1119_U51 | ~new_P2_U3406;
  assign new_P2_U5356 = ~new_P2_U5355 | ~new_P2_U5354 | ~new_P2_U5353;
  assign new_P2_U5357 = ~new_P2_U3453 | ~new_P2_U5636;
  assign new_P2_U5358 = ~new_P2_ADD_1119_U51 | ~new_P2_U5635;
  assign new_P2_U5359 = ~new_P2_R1176_U95 | ~new_P2_U3028;
  assign new_P2_U5360 = ~new_P2_U3969 | ~new_P2_U5356;
  assign new_P2_U5361 = ~P2_REG3_REG_8_ | ~n2609;
  assign new_P2_U5362 = ~new_P2_U3038 | ~new_P2_U3055;
  assign new_P2_U5363 = ~new_P2_U3036 | ~new_P2_U3057;
  assign new_P2_U5364 = ~new_P2_ADD_1119_U56 | ~new_P2_U3406;
  assign new_P2_U5365 = ~new_P2_U5362 | ~new_P2_U5363 | ~new_P2_U5364;
  assign new_P2_U5366 = ~new_P2_U3047 | ~new_P2_U3949;
  assign new_P2_U5367 = ~new_P2_U3046 | ~new_P2_ADD_1119_U56;
  assign new_P2_U5368 = ~new_P2_R1176_U100 | ~new_P2_U3028;
  assign new_P2_U5369 = ~new_P2_U3969 | ~new_P2_U5365;
  assign new_P2_U5370 = ~P2_REG3_REG_28_ | ~n2609;
  assign new_P2_U5371 = ~new_P2_U3038 | ~new_P2_U3084;
  assign new_P2_U5372 = ~new_P2_U3036 | ~new_P2_U3078;
  assign new_P2_U5373 = ~new_P2_ADD_1119_U65 | ~new_P2_U3406;
  assign new_P2_U5374 = ~new_P2_U5373 | ~new_P2_U5372 | ~new_P2_U5371;
  assign new_P2_U5375 = ~new_P2_U3485 | ~new_P2_U5636;
  assign new_P2_U5376 = ~new_P2_ADD_1119_U65 | ~new_P2_U5635;
  assign new_P2_U5377 = ~new_P2_R1176_U108 | ~new_P2_U3028;
  assign new_P2_U5378 = ~new_P2_U3969 | ~new_P2_U5374;
  assign new_P2_U5379 = ~P2_REG3_REG_19_ | ~n2609;
  assign new_P2_U5380 = ~new_P2_U3038 | ~new_P2_U3070;
  assign new_P2_U5381 = ~new_P2_U3036 | ~new_P2_U3062;
  assign new_P2_U5382 = ~new_P2_ADD_1119_U4 | ~new_P2_U3406;
  assign new_P2_U5383 = ~new_P2_U5382 | ~new_P2_U5381 | ~new_P2_U5380;
  assign new_P2_U5384 = ~new_P2_U3438 | ~new_P2_U5636;
  assign new_P2_U5385 = ~new_P2_ADD_1119_U4 | ~new_P2_U5635;
  assign new_P2_U5386 = ~new_P2_R1176_U17 | ~new_P2_U3028;
  assign new_P2_U5387 = ~new_P2_U3969 | ~new_P2_U5383;
  assign new_P2_U5388 = ~P2_REG3_REG_3_ | ~n2609;
  assign new_P2_U5389 = ~new_P2_U3038 | ~new_P2_U3085;
  assign new_P2_U5390 = ~new_P2_U3036 | ~new_P2_U3065;
  assign new_P2_U5391 = ~new_P2_ADD_1119_U74 | ~new_P2_U3406;
  assign new_P2_U5392 = ~new_P2_U5391 | ~new_P2_U5390 | ~new_P2_U5389;
  assign new_P2_U5393 = ~new_P2_U3459 | ~new_P2_U5636;
  assign new_P2_U5394 = ~new_P2_ADD_1119_U74 | ~new_P2_U5635;
  assign new_P2_U5395 = ~new_P2_R1176_U115 | ~new_P2_U3028;
  assign new_P2_U5396 = ~new_P2_U3969 | ~new_P2_U5392;
  assign new_P2_U5397 = ~P2_REG3_REG_10_ | ~n2609;
  assign new_P2_U5398 = ~new_P2_U3038 | ~new_P2_U3063;
  assign new_P2_U5399 = ~new_P2_U3036 | ~new_P2_U3067;
  assign new_P2_U5400 = ~new_P2_ADD_1119_U61 | ~new_P2_U3406;
  assign new_P2_U5401 = ~new_P2_U5400 | ~new_P2_U5399 | ~new_P2_U5398;
  assign new_P2_U5402 = ~new_P2_U3047 | ~new_P2_U3954;
  assign new_P2_U5403 = ~new_P2_U3046 | ~new_P2_ADD_1119_U61;
  assign new_P2_U5404 = ~new_P2_R1176_U104 | ~new_P2_U3028;
  assign new_P2_U5405 = ~new_P2_U3969 | ~new_P2_U5401;
  assign new_P2_U5406 = ~P2_REG3_REG_23_ | ~n2609;
  assign new_P2_U5407 = ~new_P2_U3038 | ~new_P2_U3082;
  assign new_P2_U5408 = ~new_P2_U3036 | ~new_P2_U3076;
  assign new_P2_U5409 = ~new_P2_ADD_1119_U70 | ~new_P2_U3406;
  assign new_P2_U5410 = ~new_P2_U5409 | ~new_P2_U5408 | ~new_P2_U5407;
  assign new_P2_U5411 = ~new_P2_U3471 | ~new_P2_U5636;
  assign new_P2_U5412 = ~new_P2_ADD_1119_U70 | ~new_P2_U5635;
  assign new_P2_U5413 = ~new_P2_R1176_U112 | ~new_P2_U3028;
  assign new_P2_U5414 = ~new_P2_U3969 | ~new_P2_U5410;
  assign new_P2_U5415 = ~P2_REG3_REG_14_ | ~n2609;
  assign new_P2_U5416 = ~new_P2_U3038 | ~new_P2_U3059;
  assign new_P2_U5417 = ~new_P2_U3036 | ~new_P2_U3056;
  assign new_P2_U5418 = ~new_P2_ADD_1119_U57 | ~new_P2_U3406;
  assign new_P2_U5419 = ~new_P2_U5417 | ~new_P2_U5418 | ~new_P2_U5416;
  assign new_P2_U5420 = ~new_P2_U3047 | ~new_P2_U3950;
  assign new_P2_U5421 = ~new_P2_U3046 | ~new_P2_ADD_1119_U57;
  assign new_P2_U5422 = ~new_P2_R1176_U101 | ~new_P2_U3028;
  assign new_P2_U5423 = ~new_P2_U3969 | ~new_P2_U5419;
  assign new_P2_U5424 = ~P2_REG3_REG_27_ | ~n2609;
  assign new_P2_U5425 = ~new_P2_U3038 | ~new_P2_U3073;
  assign new_P2_U5426 = ~new_P2_U3036 | ~new_P2_U3086;
  assign new_P2_U5427 = ~new_P2_ADD_1119_U52 | ~new_P2_U3406;
  assign new_P2_U5428 = ~new_P2_U5427 | ~new_P2_U5426 | ~new_P2_U5425;
  assign new_P2_U5429 = ~new_P2_U3450 | ~new_P2_U5636;
  assign new_P2_U5430 = ~new_P2_ADD_1119_U52 | ~new_P2_U5635;
  assign new_P2_U5431 = ~new_P2_R1176_U18 | ~new_P2_U3028;
  assign new_P2_U5432 = ~new_P2_U3969 | ~new_P2_U5428;
  assign new_P2_U5433 = ~P2_REG3_REG_7_ | ~n2609;
  assign new_P2_U5434 = ~new_P2_U3948 | ~new_P2_U3048;
  assign new_P2_U5435 = ~new_P2_U3415 | ~new_P2_U3347;
  assign new_P2_U5436 = ~new_P2_U3419 | ~new_P2_U3418;
  assign new_P2_U5437 = ~new_P2_U3816 | ~new_P2_U3051;
  assign new_P2_U5438 = ~new_P2_U3411;
  assign new_P2_U5439 = ~new_P2_U3015 | ~new_P2_U3415;
  assign new_P2_U5440 = ~new_P2_U3411 | ~new_P2_U3409;
  assign new_P2_U5441 = ~new_P2_U3053 | ~new_P2_U5440;
  assign new_P2_U5442 = ~new_P2_U3085 | ~new_P2_U3029;
  assign new_P2_U5443 = ~new_P2_U5441 | ~new_P2_U3085;
  assign new_P2_U5444 = ~new_P2_U3929 | ~new_P2_U3456;
  assign new_P2_U5445 = ~new_P2_U3086 | ~new_P2_U3029;
  assign new_P2_U5446 = ~new_P2_U5441 | ~new_P2_U3086;
  assign new_P2_U5447 = ~new_P2_U3929 | ~new_P2_U3453;
  assign new_P2_U5448 = ~new_P2_U3072 | ~new_P2_U3029;
  assign new_P2_U5449 = ~new_P2_U5441 | ~new_P2_U3072;
  assign new_P2_U5450 = ~new_P2_U3929 | ~new_P2_U3450;
  assign new_P2_U5451 = ~new_P2_U3073 | ~new_P2_U3029;
  assign new_P2_U5452 = ~new_P2_U5441 | ~new_P2_U3073;
  assign new_P2_U5453 = ~new_P2_U3929 | ~new_P2_U3447;
  assign new_P2_U5454 = ~new_P2_U3069 | ~new_P2_U3029;
  assign new_P2_U5455 = ~new_P2_U5441 | ~new_P2_U3069;
  assign new_P2_U5456 = ~new_P2_U3929 | ~new_P2_U3444;
  assign new_P2_U5457 = ~new_P2_U3062 | ~new_P2_U3029;
  assign new_P2_U5458 = ~new_P2_U5441 | ~new_P2_U3062;
  assign new_P2_U5459 = ~new_P2_U3929 | ~new_P2_U3441;
  assign new_P2_U5460 = ~new_P2_R1335_U8 | ~new_P2_U3029;
  assign new_P2_U5461 = ~new_P2_U5441 | ~new_P2_U3058;
  assign new_P2_U5462 = ~new_P2_R1335_U6 | ~new_P2_U3029;
  assign new_P2_U5463 = ~new_P2_U5441 | ~new_P2_U3061;
  assign new_P2_U5464 = ~new_U70 | ~new_P2_U3929 | ~new_P2_U3347;
  assign new_P2_U5465 = ~new_P2_U3066 | ~new_P2_U3029;
  assign new_P2_U5466 = ~new_P2_U5441 | ~new_P2_U3066;
  assign new_P2_U5467 = ~new_P2_U3929 | ~new_P2_U3438;
  assign new_P2_U5468 = ~new_P2_U3057 | ~new_P2_U3029;
  assign new_P2_U5469 = ~new_P2_U5441 | ~new_P2_U3057;
  assign new_P2_U5470 = ~new_P2_U3929 | ~new_P2_U3960;
  assign new_P2_U5471 = ~new_P2_U3056 | ~new_P2_U3029;
  assign new_P2_U5472 = ~new_P2_U5441 | ~new_P2_U3056;
  assign new_P2_U5473 = ~new_P2_U3929 | ~new_P2_U3949;
  assign new_P2_U5474 = ~new_P2_U3055 | ~new_P2_U3029;
  assign new_P2_U5475 = ~new_P2_U5441 | ~new_P2_U3055;
  assign new_P2_U5476 = ~new_P2_U3929 | ~new_P2_U3950;
  assign new_P2_U5477 = ~new_P2_U3059 | ~new_P2_U3029;
  assign new_P2_U5478 = ~new_P2_U5441 | ~new_P2_U3059;
  assign new_P2_U5479 = ~new_P2_U3929 | ~new_P2_U3951;
  assign new_P2_U5480 = ~new_P2_U3060 | ~new_P2_U3029;
  assign new_P2_U5481 = ~new_P2_U5441 | ~new_P2_U3060;
  assign new_P2_U5482 = ~new_P2_U3929 | ~new_P2_U3952;
  assign new_P2_U5483 = ~new_P2_U3067 | ~new_P2_U3029;
  assign new_P2_U5484 = ~new_P2_U5441 | ~new_P2_U3067;
  assign new_P2_U5485 = ~new_P2_U3929 | ~new_P2_U3953;
  assign new_P2_U5486 = ~new_P2_U3068 | ~new_P2_U3029;
  assign new_P2_U5487 = ~new_P2_U5441 | ~new_P2_U3068;
  assign new_P2_U5488 = ~new_P2_U3929 | ~new_P2_U3954;
  assign new_P2_U5489 = ~new_P2_U3063 | ~new_P2_U3029;
  assign new_P2_U5490 = ~new_P2_U5441 | ~new_P2_U3063;
  assign new_P2_U5491 = ~new_P2_U3929 | ~new_P2_U3955;
  assign new_P2_U5492 = ~new_P2_U3077 | ~new_P2_U3029;
  assign new_P2_U5493 = ~new_P2_U5441 | ~new_P2_U3077;
  assign new_P2_U5494 = ~new_P2_U3929 | ~new_P2_U3956;
  assign new_P2_U5495 = ~new_P2_U3078 | ~new_P2_U3029;
  assign new_P2_U5496 = ~new_P2_U5441 | ~new_P2_U3078;
  assign new_P2_U5497 = ~new_P2_U3929 | ~new_P2_U3957;
  assign new_P2_U5498 = ~new_P2_U3070 | ~new_P2_U3029;
  assign new_P2_U5499 = ~new_P2_U5441 | ~new_P2_U3070;
  assign new_P2_U5500 = ~new_P2_U3929 | ~new_P2_U3435;
  assign new_P2_U5501 = ~new_P2_U3083 | ~new_P2_U3029;
  assign new_P2_U5502 = ~new_P2_U5441 | ~new_P2_U3083;
  assign new_P2_U5503 = ~new_P2_U3929 | ~new_P2_U3485;
  assign new_P2_U5504 = ~new_P2_U3084 | ~new_P2_U3029;
  assign new_P2_U5505 = ~new_P2_U5441 | ~new_P2_U3084;
  assign new_P2_U5506 = ~new_P2_U3929 | ~new_P2_U3483;
  assign new_P2_U5507 = ~new_P2_U3071 | ~new_P2_U3029;
  assign new_P2_U5508 = ~new_P2_U5441 | ~new_P2_U3071;
  assign new_P2_U5509 = ~new_P2_U3929 | ~new_P2_U3480;
  assign new_P2_U5510 = ~new_P2_U3075 | ~new_P2_U3029;
  assign new_P2_U5511 = ~new_P2_U5441 | ~new_P2_U3075;
  assign new_P2_U5512 = ~new_P2_U3929 | ~new_P2_U3477;
  assign new_P2_U5513 = ~new_P2_U3076 | ~new_P2_U3029;
  assign new_P2_U5514 = ~new_P2_U5441 | ~new_P2_U3076;
  assign new_P2_U5515 = ~new_P2_U3929 | ~new_P2_U3474;
  assign new_P2_U5516 = ~new_P2_U3081 | ~new_P2_U3029;
  assign new_P2_U5517 = ~new_P2_U5441 | ~new_P2_U3081;
  assign new_P2_U5518 = ~new_P2_U3929 | ~new_P2_U3471;
  assign new_P2_U5519 = ~new_P2_U3082 | ~new_P2_U3029;
  assign new_P2_U5520 = ~new_P2_U5441 | ~new_P2_U3082;
  assign new_P2_U5521 = ~new_P2_U3929 | ~new_P2_U3468;
  assign new_P2_U5522 = ~new_P2_U3074 | ~new_P2_U3029;
  assign new_P2_U5523 = ~new_P2_U5441 | ~new_P2_U3074;
  assign new_P2_U5524 = ~new_P2_U3929 | ~new_P2_U3465;
  assign new_P2_U5525 = ~new_P2_U3065 | ~new_P2_U3029;
  assign new_P2_U5526 = ~new_P2_U5441 | ~new_P2_U3065;
  assign new_P2_U5527 = ~new_P2_U3929 | ~new_P2_U3462;
  assign new_P2_U5528 = ~new_P2_U3064 | ~new_P2_U3029;
  assign new_P2_U5529 = ~new_P2_U5441 | ~new_P2_U3064;
  assign new_P2_U5530 = ~new_P2_U3929 | ~new_P2_U3459;
  assign new_P2_U5531 = ~new_P2_U3080 | ~new_P2_U3029;
  assign new_P2_U5532 = ~new_P2_U5441 | ~new_P2_U3080;
  assign new_P2_U5533 = ~new_P2_U3929 | ~new_P2_U3432;
  assign new_P2_U5534 = ~new_P2_U3079 | ~new_P2_U3029;
  assign new_P2_U5535 = ~new_P2_U5441 | ~new_P2_U3079;
  assign new_P2_U5536 = ~new_P2_U3929 | ~new_P2_U3427;
  assign new_P2_U5537 = ~new_P2_U5438 | ~new_P2_U3053;
  assign new_P2_U5538 = ~new_P2_U3456 | ~new_P2_U5537;
  assign new_P2_U5539 = ~new_P2_U3929 | ~new_P2_U3085;
  assign new_P2_U5540 = ~new_P2_U5658 | ~new_P2_U3086;
  assign new_P2_U5541 = ~new_P2_U3453 | ~new_P2_U5537;
  assign new_P2_U5542 = ~new_P2_U3929 | ~new_P2_U3086;
  assign new_P2_U5543 = ~new_P2_U5658 | ~new_P2_U3072;
  assign new_P2_U5544 = ~new_P2_U3450 | ~new_P2_U5537;
  assign new_P2_U5545 = ~new_P2_U3929 | ~new_P2_U3072;
  assign new_P2_U5546 = ~new_P2_U5658 | ~new_P2_U3073;
  assign new_P2_U5547 = ~new_P2_U3447 | ~new_P2_U5537;
  assign new_P2_U5548 = ~new_P2_U3929 | ~new_P2_U3073;
  assign new_P2_U5549 = ~new_P2_U5658 | ~new_P2_U3069;
  assign new_P2_U5550 = ~new_P2_U3444 | ~new_P2_U5537;
  assign new_P2_U5551 = ~new_P2_U3929 | ~new_P2_U3069;
  assign new_P2_U5552 = ~new_P2_U5658 | ~new_P2_U3062;
  assign new_P2_U5553 = ~new_P2_U3441 | ~new_P2_U5537;
  assign new_P2_U5554 = ~new_P2_U3929 | ~new_P2_U3062;
  assign new_P2_U5555 = ~new_P2_U5658 | ~new_P2_U3066;
  assign new_P2_U5556 = ~new_U69 | ~new_P2_U5537 | ~new_P2_U3347;
  assign new_P2_U5557 = ~new_P2_U3929 | ~new_P2_U3058;
  assign new_P2_U5558 = ~new_P2_U3959 | ~new_P2_U5537;
  assign new_P2_U5559 = ~new_P2_U3929 | ~new_P2_U3061;
  assign new_P2_U5560 = ~new_P2_U3438 | ~new_P2_U5537;
  assign new_P2_U5561 = ~new_P2_U3929 | ~new_P2_U3066;
  assign new_P2_U5562 = ~new_P2_U5658 | ~new_P2_U3070;
  assign new_P2_U5563 = ~new_P2_U3960 | ~new_P2_U5537;
  assign new_P2_U5564 = ~new_P2_U3929 | ~new_P2_U3057;
  assign new_P2_U5565 = ~new_P2_U5658 | ~new_P2_U3056;
  assign new_P2_U5566 = ~new_P2_U3949 | ~new_P2_U5537;
  assign new_P2_U5567 = ~new_P2_U3929 | ~new_P2_U3056;
  assign new_P2_U5568 = ~new_P2_U5658 | ~new_P2_U3055;
  assign new_P2_U5569 = ~new_P2_U3950 | ~new_P2_U5537;
  assign new_P2_U5570 = ~new_P2_U3929 | ~new_P2_U3055;
  assign new_P2_U5571 = ~new_P2_U5658 | ~new_P2_U3059;
  assign new_P2_U5572 = ~new_P2_U3951 | ~new_P2_U5537;
  assign new_P2_U5573 = ~new_P2_U3929 | ~new_P2_U3059;
  assign new_P2_U5574 = ~new_P2_U5658 | ~new_P2_U3060;
  assign new_P2_U5575 = ~new_P2_U3952 | ~new_P2_U5537;
  assign new_P2_U5576 = ~new_P2_U3929 | ~new_P2_U3060;
  assign new_P2_U5577 = ~new_P2_U5658 | ~new_P2_U3067;
  assign new_P2_U5578 = ~new_P2_U3953 | ~new_P2_U5537;
  assign new_P2_U5579 = ~new_P2_U3929 | ~new_P2_U3067;
  assign new_P2_U5580 = ~new_P2_U5658 | ~new_P2_U3068;
  assign new_P2_U5581 = ~new_P2_U3954 | ~new_P2_U5537;
  assign new_P2_U5582 = ~new_P2_U3929 | ~new_P2_U3068;
  assign new_P2_U5583 = ~new_P2_U5658 | ~new_P2_U3063;
  assign new_P2_U5584 = ~new_P2_U3955 | ~new_P2_U5537;
  assign new_P2_U5585 = ~new_P2_U3929 | ~new_P2_U3063;
  assign new_P2_U5586 = ~new_P2_U5658 | ~new_P2_U3077;
  assign new_P2_U5587 = ~new_P2_U3956 | ~new_P2_U5537;
  assign new_P2_U5588 = ~new_P2_U3929 | ~new_P2_U3077;
  assign new_P2_U5589 = ~new_P2_U5658 | ~new_P2_U3078;
  assign new_P2_U5590 = ~new_P2_U3957 | ~new_P2_U5537;
  assign new_P2_U5591 = ~new_P2_U3929 | ~new_P2_U3078;
  assign new_P2_U5592 = ~new_P2_U5658 | ~new_P2_U3083;
  assign new_P2_U5593 = ~new_P2_U3435 | ~new_P2_U5537;
  assign new_P2_U5594 = ~new_P2_U3929 | ~new_P2_U3070;
  assign new_P2_U5595 = ~new_P2_U5658 | ~new_P2_U3080;
  assign new_P2_U5596 = ~new_P2_U3485 | ~new_P2_U5537;
  assign new_P2_U5597 = ~new_P2_U3929 | ~new_P2_U3083;
  assign new_P2_U5598 = ~new_P2_U5658 | ~new_P2_U3084;
  assign new_P2_U5599 = ~new_P2_U3483 | ~new_P2_U5537;
  assign new_P2_U5600 = ~new_P2_U3929 | ~new_P2_U3084;
  assign new_P2_U5601 = ~new_P2_U5658 | ~new_P2_U3071;
  assign new_P2_U5602 = ~new_P2_U3480 | ~new_P2_U5537;
  assign new_P2_U5603 = ~new_P2_U3929 | ~new_P2_U3071;
  assign new_P2_U5604 = ~new_P2_U5658 | ~new_P2_U3075;
  assign new_P2_U5605 = ~new_P2_U3477 | ~new_P2_U5537;
  assign new_P2_U5606 = ~new_P2_U3929 | ~new_P2_U3075;
  assign new_P2_U5607 = ~new_P2_U5658 | ~new_P2_U3076;
  assign new_P2_U5608 = ~new_P2_U3474 | ~new_P2_U5537;
  assign new_P2_U5609 = ~new_P2_U3929 | ~new_P2_U3076;
  assign new_P2_U5610 = ~new_P2_U5658 | ~new_P2_U3081;
  assign new_P2_U5611 = ~new_P2_U3471 | ~new_P2_U5537;
  assign new_P2_U5612 = ~new_P2_U3929 | ~new_P2_U3081;
  assign new_P2_U5613 = ~new_P2_U5658 | ~new_P2_U3082;
  assign new_P2_U5614 = ~new_P2_U3468 | ~new_P2_U5537;
  assign new_P2_U5615 = ~new_P2_U3929 | ~new_P2_U3082;
  assign new_P2_U5616 = ~new_P2_U5658 | ~new_P2_U3074;
  assign new_P2_U5617 = ~new_P2_U3465 | ~new_P2_U5537;
  assign new_P2_U5618 = ~new_P2_U3929 | ~new_P2_U3074;
  assign new_P2_U5619 = ~new_P2_U5658 | ~new_P2_U3065;
  assign new_P2_U5620 = ~new_P2_U3462 | ~new_P2_U5537;
  assign new_P2_U5621 = ~new_P2_U3929 | ~new_P2_U3065;
  assign new_P2_U5622 = ~new_P2_U5658 | ~new_P2_U3064;
  assign new_P2_U5623 = ~new_P2_U3459 | ~new_P2_U5537;
  assign new_P2_U5624 = ~new_P2_U3929 | ~new_P2_U3064;
  assign new_P2_U5625 = ~new_P2_U5658 | ~new_P2_U3085;
  assign new_P2_U5626 = ~new_P2_U3432 | ~new_P2_U5537;
  assign new_P2_U5627 = ~new_P2_U3929 | ~new_P2_U3080;
  assign new_P2_U5628 = ~new_P2_U5658 | ~new_P2_U3079;
  assign new_P2_U5629 = ~new_P2_U3427 | ~new_P2_U5537;
  assign new_P2_U5630 = ~new_P2_U3929 | ~new_P2_U3079;
  assign new_P2_U5631 = ~new_P2_U5163 | ~n2609;
  assign new_P2_U5632 = ~new_P2_U3828 | ~new_P2_U5461;
  assign new_P2_U5633 = ~new_P2_U3972 | ~new_P2_U3406;
  assign new_P2_U5634 = ~new_P2_U3946 | ~new_P2_U3972;
  assign new_P2_U5635 = ~new_P2_U5633 | ~new_P2_U3970;
  assign new_P2_U5636 = ~new_P2_U5634 | ~new_P2_U3971;
  assign new_P2_U5637 = ~new_P2_U3054 | ~new_P2_U3945;
  assign new_P2_U5638 = ~new_P2_U3054 | ~new_P2_U3330;
  assign new_P2_U5639 = ~new_P2_U3961 | ~new_P2_U3023;
  assign new_P2_U5640 = ~new_P2_U3787 | ~new_P2_U5163;
  assign new_P2_U5641 = ~new_P2_U3917 | ~new_P2_U5163 | ~new_P2_U6150 | ~new_P2_U6149;
  assign new_P2_U5642 = ~new_P2_U5652 | ~new_P2_U5646;
  assign new_P2_U5643 = ~new_P2_U3415 | ~new_P2_U3347;
  assign new_P2_U5644 = ~P2_IR_REG_24_ | ~new_P2_U3879;
  assign new_P2_U5645 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U14;
  assign new_P2_U5646 = ~new_P2_U3412;
  assign new_P2_U5647 = ~P2_IR_REG_25_ | ~new_P2_U3879;
  assign new_P2_U5648 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U112;
  assign new_P2_U5649 = ~new_P2_U3413;
  assign new_P2_U5650 = ~P2_IR_REG_26_ | ~new_P2_U3879;
  assign new_P2_U5651 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U15;
  assign new_P2_U5652 = ~new_P2_U3414;
  assign new_P2_U5653 = ~new_P2_U5646 | ~P2_B_REG;
  assign new_P2_U5654 = ~new_P2_U3412 | ~new_P2_U3331;
  assign new_P2_U5655 = ~new_P2_U5654 | ~new_P2_U5653;
  assign new_P2_U5656 = ~P2_IR_REG_23_ | ~new_P2_U3879;
  assign new_P2_U5657 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U13;
  assign new_P2_U5658 = ~new_P2_U3415;
  assign new_P2_U5659 = ~P2_D_REG_0_ | ~new_P2_U3880;
  assign new_P2_U5660 = ~new_P2_U3967 | ~new_P2_U4077;
  assign new_P2_U5661 = ~P2_D_REG_1_ | ~new_P2_U3880;
  assign new_P2_U5662 = ~new_P2_U3967 | ~new_P2_U4078;
  assign new_P2_U5663 = ~P2_IR_REG_22_ | ~new_P2_U3879;
  assign new_P2_U5664 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U114;
  assign new_P2_U5665 = ~new_P2_U3420;
  assign new_P2_U5666 = ~P2_IR_REG_19_ | ~new_P2_U3879;
  assign new_P2_U5667 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U123;
  assign new_P2_U5668 = ~new_P2_U3424;
  assign new_P2_U5669 = ~P2_IR_REG_20_ | ~new_P2_U3879;
  assign new_P2_U5670 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U119;
  assign new_P2_U5671 = ~new_P2_U3418;
  assign new_P2_U5672 = ~P2_IR_REG_21_ | ~new_P2_U3879;
  assign new_P2_U5673 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U116;
  assign new_P2_U5674 = ~new_P2_U3419;
  assign new_P2_U5675 = ~P2_IR_REG_30_ | ~new_P2_U3879;
  assign new_P2_U5676 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U104;
  assign new_P2_U5677 = ~new_P2_U3421;
  assign new_P2_U5678 = ~P2_IR_REG_29_ | ~new_P2_U3879;
  assign new_P2_U5679 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U16;
  assign new_P2_U5680 = ~new_P2_U3422;
  assign new_P2_U5681 = ~P2_IR_REG_28_ | ~new_P2_U3879;
  assign new_P2_U5682 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U107;
  assign new_P2_U5683 = ~new_P2_U3423;
  assign new_P2_U5684 = ~P2_IR_REG_0_ | ~new_P2_U3879;
  assign new_P2_U5685 = ~P2_IR_REG_31_ | ~P2_IR_REG_0_;
  assign new_P2_U5686 = ~P2_IR_REG_27_ | ~new_P2_U3879;
  assign new_P2_U5687 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U110;
  assign new_P2_U5688 = ~new_P2_U3426;
  assign new_P2_U5689 = ~new_U93 | ~new_P2_U3347;
  assign new_P2_U5690 = ~new_P2_U3425 | ~new_P2_U3945;
  assign new_P2_U5691 = ~new_P2_U3427;
  assign new_P2_U5692 = ~new_P2_U3420 | ~new_P2_U5674;
  assign new_P2_U5693 = ~new_P2_U5665 | ~new_P2_U4109;
  assign new_P2_U5694 = ~P2_D_REG_1_ | ~new_P2_U4076;
  assign new_P2_U5695 = ~new_P2_U4078 | ~new_P2_U3333;
  assign new_P2_U5696 = ~new_P2_U3429;
  assign new_P2_U5697 = ~new_P2_U5642 | ~new_P2_U3333;
  assign new_P2_U5698 = ~P2_D_REG_0_ | ~new_P2_U4076;
  assign new_P2_U5699 = ~new_P2_U3428;
  assign new_P2_U5700 = ~P2_REG0_REG_0_ | ~new_P2_U3881;
  assign new_P2_U5701 = ~new_P2_U3966 | ~new_P2_U4129;
  assign new_P2_U5702 = ~P2_IR_REG_1_ | ~new_P2_U3879;
  assign new_P2_U5703 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U42;
  assign new_P2_U5704 = ~new_U82 | ~new_P2_U3347;
  assign new_P2_U5705 = ~new_P2_U3431 | ~new_P2_U3945;
  assign new_P2_U5706 = ~new_P2_U3432;
  assign new_P2_U5707 = ~P2_REG0_REG_1_ | ~new_P2_U3881;
  assign new_P2_U5708 = ~new_P2_U3966 | ~new_P2_U4153;
  assign new_P2_U5709 = ~P2_IR_REG_2_ | ~new_P2_U3879;
  assign new_P2_U5710 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U17;
  assign new_P2_U5711 = ~new_U71 | ~new_P2_U3347;
  assign new_P2_U5712 = ~new_P2_U3434 | ~new_P2_U3945;
  assign new_P2_U5713 = ~new_P2_U3435;
  assign new_P2_U5714 = ~P2_REG0_REG_2_ | ~new_P2_U3881;
  assign new_P2_U5715 = ~new_P2_U3966 | ~new_P2_U4172;
  assign new_P2_U5716 = ~P2_IR_REG_3_ | ~new_P2_U3879;
  assign new_P2_U5717 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U18;
  assign new_P2_U5718 = ~new_U68 | ~new_P2_U3347;
  assign new_P2_U5719 = ~new_P2_U3437 | ~new_P2_U3945;
  assign new_P2_U5720 = ~new_P2_U3438;
  assign new_P2_U5721 = ~P2_REG0_REG_3_ | ~new_P2_U3881;
  assign new_P2_U5722 = ~new_P2_U3966 | ~new_P2_U4191;
  assign new_P2_U5723 = ~P2_IR_REG_4_ | ~new_P2_U3879;
  assign new_P2_U5724 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U19;
  assign new_P2_U5725 = ~new_U67 | ~new_P2_U3347;
  assign new_P2_U5726 = ~new_P2_U3440 | ~new_P2_U3945;
  assign new_P2_U5727 = ~new_P2_U3441;
  assign new_P2_U5728 = ~P2_REG0_REG_4_ | ~new_P2_U3881;
  assign new_P2_U5729 = ~new_P2_U3966 | ~new_P2_U4210;
  assign new_P2_U5730 = ~P2_IR_REG_5_ | ~new_P2_U3879;
  assign new_P2_U5731 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U101;
  assign new_P2_U5732 = ~new_U66 | ~new_P2_U3347;
  assign new_P2_U5733 = ~new_P2_U3443 | ~new_P2_U3945;
  assign new_P2_U5734 = ~new_P2_U3444;
  assign new_P2_U5735 = ~P2_REG0_REG_5_ | ~new_P2_U3881;
  assign new_P2_U5736 = ~new_P2_U3966 | ~new_P2_U4229;
  assign new_P2_U5737 = ~P2_IR_REG_6_ | ~new_P2_U3879;
  assign new_P2_U5738 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U20;
  assign new_P2_U5739 = ~new_U65 | ~new_P2_U3347;
  assign new_P2_U5740 = ~new_P2_U3446 | ~new_P2_U3945;
  assign new_P2_U5741 = ~new_P2_U3447;
  assign new_P2_U5742 = ~P2_REG0_REG_6_ | ~new_P2_U3881;
  assign new_P2_U5743 = ~new_P2_U3966 | ~new_P2_U4248;
  assign new_P2_U5744 = ~P2_IR_REG_7_ | ~new_P2_U3879;
  assign new_P2_U5745 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U21;
  assign new_P2_U5746 = ~new_U64 | ~new_P2_U3347;
  assign new_P2_U5747 = ~new_P2_U3449 | ~new_P2_U3945;
  assign new_P2_U5748 = ~new_P2_U3450;
  assign new_P2_U5749 = ~P2_REG0_REG_7_ | ~new_P2_U3881;
  assign new_P2_U5750 = ~new_P2_U3966 | ~new_P2_U4267;
  assign new_P2_U5751 = ~P2_IR_REG_8_ | ~new_P2_U3879;
  assign new_P2_U5752 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U22;
  assign new_P2_U5753 = ~new_U63 | ~new_P2_U3347;
  assign new_P2_U5754 = ~new_P2_U3452 | ~new_P2_U3945;
  assign new_P2_U5755 = ~new_P2_U3453;
  assign new_P2_U5756 = ~P2_REG0_REG_8_ | ~new_P2_U3881;
  assign new_P2_U5757 = ~new_P2_U3966 | ~new_P2_U4286;
  assign new_P2_U5758 = ~P2_IR_REG_9_ | ~new_P2_U3879;
  assign new_P2_U5759 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U99;
  assign new_P2_U5760 = ~new_U62 | ~new_P2_U3347;
  assign new_P2_U5761 = ~new_P2_U3455 | ~new_P2_U3945;
  assign new_P2_U5762 = ~new_P2_U3456;
  assign new_P2_U5763 = ~P2_REG0_REG_9_ | ~new_P2_U3881;
  assign new_P2_U5764 = ~new_P2_U3966 | ~new_P2_U4305;
  assign new_P2_U5765 = ~P2_IR_REG_10_ | ~new_P2_U3879;
  assign new_P2_U5766 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U6;
  assign new_P2_U5767 = ~new_U92 | ~new_P2_U3347;
  assign new_P2_U5768 = ~new_P2_U3458 | ~new_P2_U3945;
  assign new_P2_U5769 = ~new_P2_U3459;
  assign new_P2_U5770 = ~P2_REG0_REG_10_ | ~new_P2_U3881;
  assign new_P2_U5771 = ~new_P2_U3966 | ~new_P2_U4324;
  assign new_P2_U5772 = ~P2_IR_REG_11_ | ~new_P2_U3879;
  assign new_P2_U5773 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U7;
  assign new_P2_U5774 = ~new_U91 | ~new_P2_U3347;
  assign new_P2_U5775 = ~new_P2_U3461 | ~new_P2_U3945;
  assign new_P2_U5776 = ~new_P2_U3462;
  assign new_P2_U5777 = ~P2_REG0_REG_11_ | ~new_P2_U3881;
  assign new_P2_U5778 = ~new_P2_U3966 | ~new_P2_U4343;
  assign new_P2_U5779 = ~P2_IR_REG_12_ | ~new_P2_U3879;
  assign new_P2_U5780 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U8;
  assign new_P2_U5781 = ~new_U90 | ~new_P2_U3347;
  assign new_P2_U5782 = ~new_P2_U3464 | ~new_P2_U3945;
  assign new_P2_U5783 = ~new_P2_U3465;
  assign new_P2_U5784 = ~P2_REG0_REG_12_ | ~new_P2_U3881;
  assign new_P2_U5785 = ~new_P2_U3966 | ~new_P2_U4362;
  assign new_P2_U5786 = ~P2_IR_REG_13_ | ~new_P2_U3879;
  assign new_P2_U5787 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U127;
  assign new_P2_U5788 = ~new_U89 | ~new_P2_U3347;
  assign new_P2_U5789 = ~new_P2_U3467 | ~new_P2_U3945;
  assign new_P2_U5790 = ~new_P2_U3468;
  assign new_P2_U5791 = ~P2_REG0_REG_13_ | ~new_P2_U3881;
  assign new_P2_U5792 = ~new_P2_U3966 | ~new_P2_U4381;
  assign new_P2_U5793 = ~P2_IR_REG_14_ | ~new_P2_U3879;
  assign new_P2_U5794 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U9;
  assign new_P2_U5795 = ~new_U88 | ~new_P2_U3347;
  assign new_P2_U5796 = ~new_P2_U3470 | ~new_P2_U3945;
  assign new_P2_U5797 = ~new_P2_U3471;
  assign new_P2_U5798 = ~P2_REG0_REG_14_ | ~new_P2_U3881;
  assign new_P2_U5799 = ~new_P2_U3966 | ~new_P2_U4400;
  assign new_P2_U5800 = ~P2_IR_REG_15_ | ~new_P2_U3879;
  assign new_P2_U5801 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U10;
  assign new_P2_U5802 = ~new_U87 | ~new_P2_U3347;
  assign new_P2_U5803 = ~new_P2_U3473 | ~new_P2_U3945;
  assign new_P2_U5804 = ~new_P2_U3474;
  assign new_P2_U5805 = ~P2_REG0_REG_15_ | ~new_P2_U3881;
  assign new_P2_U5806 = ~new_P2_U3966 | ~new_P2_U4419;
  assign new_P2_U5807 = ~P2_IR_REG_16_ | ~new_P2_U3879;
  assign new_P2_U5808 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U11;
  assign new_P2_U5809 = ~new_U86 | ~new_P2_U3347;
  assign new_P2_U5810 = ~new_P2_U3476 | ~new_P2_U3945;
  assign new_P2_U5811 = ~new_P2_U3477;
  assign new_P2_U5812 = ~P2_REG0_REG_16_ | ~new_P2_U3881;
  assign new_P2_U5813 = ~new_P2_U3966 | ~new_P2_U4438;
  assign new_P2_U5814 = ~P2_IR_REG_17_ | ~new_P2_U3879;
  assign new_P2_U5815 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U125;
  assign new_P2_U5816 = ~new_U85 | ~new_P2_U3347;
  assign new_P2_U5817 = ~new_P2_U3479 | ~new_P2_U3945;
  assign new_P2_U5818 = ~new_P2_U3480;
  assign new_P2_U5819 = ~P2_REG0_REG_17_ | ~new_P2_U3881;
  assign new_P2_U5820 = ~new_P2_U3966 | ~new_P2_U4457;
  assign new_P2_U5821 = ~P2_IR_REG_18_ | ~new_P2_U3879;
  assign new_P2_U5822 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U12;
  assign new_P2_U5823 = ~new_U84 | ~new_P2_U3347;
  assign new_P2_U5824 = ~new_P2_U3482 | ~new_P2_U3945;
  assign new_P2_U5825 = ~new_P2_U3483;
  assign new_P2_U5826 = ~P2_REG0_REG_18_ | ~new_P2_U3881;
  assign new_P2_U5827 = ~new_P2_U3966 | ~new_P2_U4476;
  assign new_P2_U5828 = ~new_U83 | ~new_P2_U3347;
  assign new_P2_U5829 = ~new_P2_U3424 | ~new_P2_U3945;
  assign new_P2_U5830 = ~new_P2_U3485;
  assign new_P2_U5831 = ~P2_REG0_REG_19_ | ~new_P2_U3881;
  assign new_P2_U5832 = ~new_P2_U3966 | ~new_P2_U4495;
  assign new_P2_U5833 = ~P2_REG0_REG_20_ | ~new_P2_U3881;
  assign new_P2_U5834 = ~new_P2_U3966 | ~new_P2_U4514;
  assign new_P2_U5835 = ~P2_REG0_REG_21_ | ~new_P2_U3881;
  assign new_P2_U5836 = ~new_P2_U3966 | ~new_P2_U4533;
  assign new_P2_U5837 = ~P2_REG0_REG_22_ | ~new_P2_U3881;
  assign new_P2_U5838 = ~new_P2_U3966 | ~new_P2_U4552;
  assign new_P2_U5839 = ~P2_REG0_REG_23_ | ~new_P2_U3881;
  assign new_P2_U5840 = ~new_P2_U3966 | ~new_P2_U4571;
  assign new_P2_U5841 = ~P2_REG0_REG_24_ | ~new_P2_U3881;
  assign new_P2_U5842 = ~new_P2_U3966 | ~new_P2_U4590;
  assign new_P2_U5843 = ~P2_REG0_REG_25_ | ~new_P2_U3881;
  assign new_P2_U5844 = ~new_P2_U3966 | ~new_P2_U4609;
  assign new_P2_U5845 = ~P2_REG0_REG_26_ | ~new_P2_U3881;
  assign new_P2_U5846 = ~new_P2_U3966 | ~new_P2_U4628;
  assign new_P2_U5847 = ~P2_REG0_REG_27_ | ~new_P2_U3881;
  assign new_P2_U5848 = ~new_P2_U3966 | ~new_P2_U4647;
  assign new_P2_U5849 = ~P2_REG0_REG_28_ | ~new_P2_U3881;
  assign new_P2_U5850 = ~new_P2_U3966 | ~new_P2_U4666;
  assign new_P2_U5851 = ~P2_REG0_REG_29_ | ~new_P2_U3881;
  assign new_P2_U5852 = ~new_P2_U3966 | ~new_P2_U4686;
  assign new_P2_U5853 = ~P2_REG0_REG_30_ | ~new_P2_U3881;
  assign new_P2_U5854 = ~new_P2_U3966 | ~new_P2_U4693;
  assign new_P2_U5855 = ~P2_REG0_REG_31_ | ~new_P2_U3881;
  assign new_P2_U5856 = ~new_P2_U3966 | ~new_P2_U4696;
  assign new_P2_U5857 = ~P2_REG1_REG_0_ | ~new_P2_U3882;
  assign new_P2_U5858 = ~new_P2_U3965 | ~new_P2_U4129;
  assign new_P2_U5859 = ~P2_REG1_REG_1_ | ~new_P2_U3882;
  assign new_P2_U5860 = ~new_P2_U3965 | ~new_P2_U4153;
  assign new_P2_U5861 = ~P2_REG1_REG_2_ | ~new_P2_U3882;
  assign new_P2_U5862 = ~new_P2_U3965 | ~new_P2_U4172;
  assign new_P2_U5863 = ~P2_REG1_REG_3_ | ~new_P2_U3882;
  assign new_P2_U5864 = ~new_P2_U3965 | ~new_P2_U4191;
  assign new_P2_U5865 = ~P2_REG1_REG_4_ | ~new_P2_U3882;
  assign new_P2_U5866 = ~new_P2_U3965 | ~new_P2_U4210;
  assign new_P2_U5867 = ~P2_REG1_REG_5_ | ~new_P2_U3882;
  assign new_P2_U5868 = ~new_P2_U3965 | ~new_P2_U4229;
  assign new_P2_U5869 = ~P2_REG1_REG_6_ | ~new_P2_U3882;
  assign new_P2_U5870 = ~new_P2_U3965 | ~new_P2_U4248;
  assign new_P2_U5871 = ~P2_REG1_REG_7_ | ~new_P2_U3882;
  assign new_P2_U5872 = ~new_P2_U3965 | ~new_P2_U4267;
  assign new_P2_U5873 = ~P2_REG1_REG_8_ | ~new_P2_U3882;
  assign new_P2_U5874 = ~new_P2_U3965 | ~new_P2_U4286;
  assign new_P2_U5875 = ~P2_REG1_REG_9_ | ~new_P2_U3882;
  assign new_P2_U5876 = ~new_P2_U3965 | ~new_P2_U4305;
  assign new_P2_U5877 = ~P2_REG1_REG_10_ | ~new_P2_U3882;
  assign new_P2_U5878 = ~new_P2_U3965 | ~new_P2_U4324;
  assign new_P2_U5879 = ~P2_REG1_REG_11_ | ~new_P2_U3882;
  assign new_P2_U5880 = ~new_P2_U3965 | ~new_P2_U4343;
  assign new_P2_U5881 = ~P2_REG1_REG_12_ | ~new_P2_U3882;
  assign new_P2_U5882 = ~new_P2_U3965 | ~new_P2_U4362;
  assign new_P2_U5883 = ~P2_REG1_REG_13_ | ~new_P2_U3882;
  assign new_P2_U5884 = ~new_P2_U3965 | ~new_P2_U4381;
  assign new_P2_U5885 = ~P2_REG1_REG_14_ | ~new_P2_U3882;
  assign new_P2_U5886 = ~new_P2_U3965 | ~new_P2_U4400;
  assign new_P2_U5887 = ~P2_REG1_REG_15_ | ~new_P2_U3882;
  assign new_P2_U5888 = ~new_P2_U3965 | ~new_P2_U4419;
  assign new_P2_U5889 = ~P2_REG1_REG_16_ | ~new_P2_U3882;
  assign new_P2_U5890 = ~new_P2_U3965 | ~new_P2_U4438;
  assign new_P2_U5891 = ~P2_REG1_REG_17_ | ~new_P2_U3882;
  assign new_P2_U5892 = ~new_P2_U3965 | ~new_P2_U4457;
  assign new_P2_U5893 = ~P2_REG1_REG_18_ | ~new_P2_U3882;
  assign new_P2_U5894 = ~new_P2_U3965 | ~new_P2_U4476;
  assign new_P2_U5895 = ~P2_REG1_REG_19_ | ~new_P2_U3882;
  assign new_P2_U5896 = ~new_P2_U3965 | ~new_P2_U4495;
  assign new_P2_U5897 = ~P2_REG1_REG_20_ | ~new_P2_U3882;
  assign new_P2_U5898 = ~new_P2_U3965 | ~new_P2_U4514;
  assign new_P2_U5899 = ~P2_REG1_REG_21_ | ~new_P2_U3882;
  assign new_P2_U5900 = ~new_P2_U3965 | ~new_P2_U4533;
  assign new_P2_U5901 = ~P2_REG1_REG_22_ | ~new_P2_U3882;
  assign new_P2_U5902 = ~new_P2_U3965 | ~new_P2_U4552;
  assign new_P2_U5903 = ~P2_REG1_REG_23_ | ~new_P2_U3882;
  assign new_P2_U5904 = ~new_P2_U3965 | ~new_P2_U4571;
  assign new_P2_U5905 = ~P2_REG1_REG_24_ | ~new_P2_U3882;
  assign new_P2_U5906 = ~new_P2_U3965 | ~new_P2_U4590;
  assign new_P2_U5907 = ~P2_REG1_REG_25_ | ~new_P2_U3882;
  assign new_P2_U5908 = ~new_P2_U3965 | ~new_P2_U4609;
  assign new_P2_U5909 = ~P2_REG1_REG_26_ | ~new_P2_U3882;
  assign new_P2_U5910 = ~new_P2_U3965 | ~new_P2_U4628;
  assign new_P2_U5911 = ~P2_REG1_REG_27_ | ~new_P2_U3882;
  assign new_P2_U5912 = ~new_P2_U3965 | ~new_P2_U4647;
  assign new_P2_U5913 = ~P2_REG1_REG_28_ | ~new_P2_U3882;
  assign new_P2_U5914 = ~new_P2_U3965 | ~new_P2_U4666;
  assign new_P2_U5915 = ~P2_REG1_REG_29_ | ~new_P2_U3882;
  assign new_P2_U5916 = ~new_P2_U3965 | ~new_P2_U4686;
  assign new_P2_U5917 = ~P2_REG1_REG_30_ | ~new_P2_U3882;
  assign new_P2_U5918 = ~new_P2_U3965 | ~new_P2_U4693;
  assign new_P2_U5919 = ~P2_REG1_REG_31_ | ~new_P2_U3882;
  assign new_P2_U5920 = ~new_P2_U3965 | ~new_P2_U4696;
  assign new_P2_U5921 = ~P2_REG2_REG_0_ | ~new_P2_U3391;
  assign new_P2_U5922 = ~new_P2_U3964 | ~new_P2_U3348;
  assign new_P2_U5923 = ~P2_REG2_REG_1_ | ~new_P2_U3391;
  assign new_P2_U5924 = ~new_P2_U3964 | ~new_P2_U3349;
  assign new_P2_U5925 = ~P2_REG2_REG_2_ | ~new_P2_U3391;
  assign new_P2_U5926 = ~new_P2_U3964 | ~new_P2_U3350;
  assign new_P2_U5927 = ~P2_REG2_REG_3_ | ~new_P2_U3391;
  assign new_P2_U5928 = ~new_P2_U3964 | ~new_P2_U3351;
  assign new_P2_U5929 = ~P2_REG2_REG_4_ | ~new_P2_U3391;
  assign new_P2_U5930 = ~new_P2_U3964 | ~new_P2_U3352;
  assign new_P2_U5931 = ~P2_REG2_REG_5_ | ~new_P2_U3391;
  assign new_P2_U5932 = ~new_P2_U3964 | ~new_P2_U3353;
  assign new_P2_U5933 = ~P2_REG2_REG_6_ | ~new_P2_U3391;
  assign new_P2_U5934 = ~new_P2_U3964 | ~new_P2_U3354;
  assign new_P2_U5935 = ~P2_REG2_REG_7_ | ~new_P2_U3391;
  assign new_P2_U5936 = ~new_P2_U3964 | ~new_P2_U3355;
  assign new_P2_U5937 = ~P2_REG2_REG_8_ | ~new_P2_U3391;
  assign new_P2_U5938 = ~new_P2_U3964 | ~new_P2_U3356;
  assign new_P2_U5939 = ~P2_REG2_REG_9_ | ~new_P2_U3391;
  assign new_P2_U5940 = ~new_P2_U3964 | ~new_P2_U3357;
  assign new_P2_U5941 = ~P2_REG2_REG_10_ | ~new_P2_U3391;
  assign new_P2_U5942 = ~new_P2_U3964 | ~new_P2_U3358;
  assign new_P2_U5943 = ~P2_REG2_REG_11_ | ~new_P2_U3391;
  assign new_P2_U5944 = ~new_P2_U3964 | ~new_P2_U3359;
  assign new_P2_U5945 = ~P2_REG2_REG_12_ | ~new_P2_U3391;
  assign new_P2_U5946 = ~new_P2_U3964 | ~new_P2_U3360;
  assign new_P2_U5947 = ~P2_REG2_REG_13_ | ~new_P2_U3391;
  assign new_P2_U5948 = ~new_P2_U3964 | ~new_P2_U3361;
  assign new_P2_U5949 = ~P2_REG2_REG_14_ | ~new_P2_U3391;
  assign new_P2_U5950 = ~new_P2_U3964 | ~new_P2_U3362;
  assign new_P2_U5951 = ~P2_REG2_REG_15_ | ~new_P2_U3391;
  assign new_P2_U5952 = ~new_P2_U3964 | ~new_P2_U3363;
  assign new_P2_U5953 = ~P2_REG2_REG_16_ | ~new_P2_U3391;
  assign new_P2_U5954 = ~new_P2_U3964 | ~new_P2_U3364;
  assign new_P2_U5955 = ~P2_REG2_REG_17_ | ~new_P2_U3391;
  assign new_P2_U5956 = ~new_P2_U3964 | ~new_P2_U3365;
  assign new_P2_U5957 = ~P2_REG2_REG_18_ | ~new_P2_U3391;
  assign new_P2_U5958 = ~new_P2_U3964 | ~new_P2_U3366;
  assign new_P2_U5959 = ~P2_REG2_REG_19_ | ~new_P2_U3391;
  assign new_P2_U5960 = ~new_P2_U3964 | ~new_P2_U3367;
  assign new_P2_U5961 = ~P2_REG2_REG_20_ | ~new_P2_U3391;
  assign new_P2_U5962 = ~new_P2_U3964 | ~new_P2_U3369;
  assign new_P2_U5963 = ~P2_REG2_REG_21_ | ~new_P2_U3391;
  assign new_P2_U5964 = ~new_P2_U3964 | ~new_P2_U3371;
  assign new_P2_U5965 = ~P2_REG2_REG_22_ | ~new_P2_U3391;
  assign new_P2_U5966 = ~new_P2_U3964 | ~new_P2_U3373;
  assign new_P2_U5967 = ~P2_REG2_REG_23_ | ~new_P2_U3391;
  assign new_P2_U5968 = ~new_P2_U3964 | ~new_P2_U3375;
  assign new_P2_U5969 = ~P2_REG2_REG_24_ | ~new_P2_U3391;
  assign new_P2_U5970 = ~new_P2_U3964 | ~new_P2_U3377;
  assign new_P2_U5971 = ~P2_REG2_REG_25_ | ~new_P2_U3391;
  assign new_P2_U5972 = ~new_P2_U3964 | ~new_P2_U3379;
  assign new_P2_U5973 = ~P2_REG2_REG_26_ | ~new_P2_U3391;
  assign new_P2_U5974 = ~new_P2_U3964 | ~new_P2_U3381;
  assign new_P2_U5975 = ~P2_REG2_REG_27_ | ~new_P2_U3391;
  assign new_P2_U5976 = ~new_P2_U3964 | ~new_P2_U3383;
  assign new_P2_U5977 = ~P2_REG2_REG_28_ | ~new_P2_U3391;
  assign new_P2_U5978 = ~new_P2_U3964 | ~new_P2_U3385;
  assign new_P2_U5979 = ~P2_REG2_REG_29_ | ~new_P2_U3391;
  assign new_P2_U5980 = ~new_P2_U3964 | ~new_P2_U3387;
  assign new_P2_U5981 = ~P2_REG2_REG_30_ | ~new_P2_U3391;
  assign new_P2_U5982 = ~new_P2_U3968 | ~new_P2_U3964;
  assign new_P2_U5983 = ~P2_REG2_REG_31_ | ~new_P2_U3391;
  assign new_P2_U5984 = ~new_P2_U3968 | ~new_P2_U3964;
  assign new_P2_U5985 = ~P2_DATAO_REG_0_ | ~new_P2_U3400;
  assign new_P2_U5986 = ~n2619 | ~new_P2_U3079;
  assign new_P2_U5987 = ~P2_DATAO_REG_1_ | ~new_P2_U3400;
  assign new_P2_U5988 = ~n2619 | ~new_P2_U3080;
  assign new_P2_U5989 = ~P2_DATAO_REG_2_ | ~new_P2_U3400;
  assign new_P2_U5990 = ~n2619 | ~new_P2_U3070;
  assign new_P2_U5991 = ~P2_DATAO_REG_3_ | ~new_P2_U3400;
  assign new_P2_U5992 = ~n2619 | ~new_P2_U3066;
  assign new_P2_U5993 = ~P2_DATAO_REG_4_ | ~new_P2_U3400;
  assign new_P2_U5994 = ~n2619 | ~new_P2_U3062;
  assign new_P2_U5995 = ~P2_DATAO_REG_5_ | ~new_P2_U3400;
  assign new_P2_U5996 = ~n2619 | ~new_P2_U3069;
  assign new_P2_U5997 = ~P2_DATAO_REG_6_ | ~new_P2_U3400;
  assign new_P2_U5998 = ~n2619 | ~new_P2_U3073;
  assign new_P2_U5999 = ~P2_DATAO_REG_7_ | ~new_P2_U3400;
  assign new_P2_U6000 = ~n2619 | ~new_P2_U3072;
  assign new_P2_U6001 = ~P2_DATAO_REG_8_ | ~new_P2_U3400;
  assign new_P2_U6002 = ~n2619 | ~new_P2_U3086;
  assign new_P2_U6003 = ~P2_DATAO_REG_9_ | ~new_P2_U3400;
  assign new_P2_U6004 = ~n2619 | ~new_P2_U3085;
  assign new_P2_U6005 = ~P2_DATAO_REG_10_ | ~new_P2_U3400;
  assign new_P2_U6006 = ~n2619 | ~new_P2_U3064;
  assign new_P2_U6007 = ~P2_DATAO_REG_11_ | ~new_P2_U3400;
  assign new_P2_U6008 = ~n2619 | ~new_P2_U3065;
  assign new_P2_U6009 = ~P2_DATAO_REG_12_ | ~new_P2_U3400;
  assign new_P2_U6010 = ~n2619 | ~new_P2_U3074;
  assign new_P2_U6011 = ~P2_DATAO_REG_13_ | ~new_P2_U3400;
  assign new_P2_U6012 = ~n2619 | ~new_P2_U3082;
  assign new_P2_U6013 = ~P2_DATAO_REG_14_ | ~new_P2_U3400;
  assign new_P2_U6014 = ~n2619 | ~new_P2_U3081;
  assign new_P2_U6015 = ~P2_DATAO_REG_15_ | ~new_P2_U3400;
  assign new_P2_U6016 = ~n2619 | ~new_P2_U3076;
  assign new_P2_U6017 = ~P2_DATAO_REG_16_ | ~new_P2_U3400;
  assign new_P2_U6018 = ~n2619 | ~new_P2_U3075;
  assign new_P2_U6019 = ~P2_DATAO_REG_17_ | ~new_P2_U3400;
  assign new_P2_U6020 = ~n2619 | ~new_P2_U3071;
  assign new_P2_U6021 = ~P2_DATAO_REG_18_ | ~new_P2_U3400;
  assign new_P2_U6022 = ~n2619 | ~new_P2_U3084;
  assign new_P2_U6023 = ~P2_DATAO_REG_19_ | ~new_P2_U3400;
  assign new_P2_U6024 = ~n2619 | ~new_P2_U3083;
  assign new_P2_U6025 = ~P2_DATAO_REG_20_ | ~new_P2_U3400;
  assign new_P2_U6026 = ~n2619 | ~new_P2_U3078;
  assign new_P2_U6027 = ~P2_DATAO_REG_21_ | ~new_P2_U3400;
  assign new_P2_U6028 = ~n2619 | ~new_P2_U3077;
  assign new_P2_U6029 = ~P2_DATAO_REG_22_ | ~new_P2_U3400;
  assign new_P2_U6030 = ~n2619 | ~new_P2_U3063;
  assign new_P2_U6031 = ~P2_DATAO_REG_23_ | ~new_P2_U3400;
  assign new_P2_U6032 = ~n2619 | ~new_P2_U3068;
  assign new_P2_U6033 = ~P2_DATAO_REG_24_ | ~new_P2_U3400;
  assign new_P2_U6034 = ~n2619 | ~new_P2_U3067;
  assign new_P2_U6035 = ~P2_DATAO_REG_25_ | ~new_P2_U3400;
  assign new_P2_U6036 = ~n2619 | ~new_P2_U3060;
  assign new_P2_U6037 = ~P2_DATAO_REG_26_ | ~new_P2_U3400;
  assign new_P2_U6038 = ~n2619 | ~new_P2_U3059;
  assign new_P2_U6039 = ~P2_DATAO_REG_27_ | ~new_P2_U3400;
  assign new_P2_U6040 = ~n2619 | ~new_P2_U3055;
  assign new_P2_U6041 = ~P2_DATAO_REG_28_ | ~new_P2_U3400;
  assign new_P2_U6042 = ~n2619 | ~new_P2_U3056;
  assign new_P2_U6043 = ~P2_DATAO_REG_29_ | ~new_P2_U3400;
  assign new_P2_U6044 = ~n2619 | ~new_P2_U3057;
  assign new_P2_U6045 = ~P2_DATAO_REG_30_ | ~new_P2_U3400;
  assign new_P2_U6046 = ~n2619 | ~new_P2_U3061;
  assign new_P2_U6047 = ~P2_DATAO_REG_31_ | ~new_P2_U3400;
  assign new_P2_U6048 = ~n2619 | ~new_P2_U3058;
  assign new_P2_U6049 = ~new_P2_R1312_U18 | ~new_P2_U5157;
  assign new_P2_U6050 = ~new_P2_U5161 | ~new_P2_U3916;
  assign new_P2_U6051 = ~new_P2_U5658 | ~new_P2_U3403;
  assign new_P2_U6052 = ~new_P2_U3420 | ~new_P2_U3415;
  assign new_P2_U6053 = ~new_P2_U3960 | ~new_P2_U3057;
  assign new_P2_U6054 = ~new_P2_U3386 | ~new_P2_U4652;
  assign new_P2_U6055 = ~new_P2_U6054 | ~new_P2_U6053;
  assign new_P2_U6056 = ~new_P2_U3949 | ~new_P2_U3056;
  assign new_P2_U6057 = ~new_P2_U3384 | ~new_P2_U4633;
  assign new_P2_U6058 = ~new_P2_U6057 | ~new_P2_U6056;
  assign new_P2_U6059 = ~new_P2_U3950 | ~new_P2_U3055;
  assign new_P2_U6060 = ~new_P2_U3382 | ~new_P2_U4614;
  assign new_P2_U6061 = ~new_P2_U6060 | ~new_P2_U6059;
  assign new_P2_U6062 = ~new_P2_U3953 | ~new_P2_U3067;
  assign new_P2_U6063 = ~new_P2_U3376 | ~new_P2_U4557;
  assign new_P2_U6064 = ~new_P2_U6063 | ~new_P2_U6062;
  assign new_P2_U6065 = ~new_P2_U3954 | ~new_P2_U3068;
  assign new_P2_U6066 = ~new_P2_U3374 | ~new_P2_U4538;
  assign new_P2_U6067 = ~new_P2_U6066 | ~new_P2_U6065;
  assign new_P2_U6068 = ~new_P2_U3956 | ~new_P2_U3077;
  assign new_P2_U6069 = ~new_P2_U3370 | ~new_P2_U4500;
  assign new_P2_U6070 = ~new_P2_U6069 | ~new_P2_U6068;
  assign new_P2_U6071 = ~new_P2_U3955 | ~new_P2_U3063;
  assign new_P2_U6072 = ~new_P2_U3372 | ~new_P2_U4519;
  assign new_P2_U6073 = ~new_P2_U6072 | ~new_P2_U6071;
  assign new_P2_U6074 = ~new_P2_U3952 | ~new_P2_U3060;
  assign new_P2_U6075 = ~new_P2_U3378 | ~new_P2_U4576;
  assign new_P2_U6076 = ~new_P2_U6075 | ~new_P2_U6074;
  assign new_P2_U6077 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_U6078 = ~new_P2_U3380 | ~new_P2_U4595;
  assign new_P2_U6079 = ~new_P2_U6078 | ~new_P2_U6077;
  assign new_P2_U6080 = ~new_P2_U3959 | ~new_P2_U3061;
  assign new_P2_U6081 = ~new_P2_U3388 | ~new_P2_U4670;
  assign new_P2_U6082 = ~new_P2_U6081 | ~new_P2_U6080;
  assign new_P2_U6083 = ~new_P2_U3958 | ~new_P2_U3058;
  assign new_P2_U6084 = ~new_P2_U3389 | ~new_P2_U4690;
  assign new_P2_U6085 = ~new_P2_U6084 | ~new_P2_U6083;
  assign new_P2_U6086 = ~new_P2_U5797 | ~new_P2_U4367;
  assign new_P2_U6087 = ~new_P2_U3471 | ~new_P2_U3081;
  assign new_P2_U6088 = ~new_P2_U6087 | ~new_P2_U6086;
  assign new_P2_U6089 = ~new_P2_U5706 | ~new_P2_U4115;
  assign new_P2_U6090 = ~new_P2_U3432 | ~new_P2_U3080;
  assign new_P2_U6091 = ~new_P2_U6090 | ~new_P2_U6089;
  assign new_P2_U6092 = ~new_P2_U5691 | ~new_P2_U4139;
  assign new_P2_U6093 = ~new_P2_U3427 | ~new_P2_U3079;
  assign new_P2_U6094 = ~new_P2_U6093 | ~new_P2_U6092;
  assign new_P2_U6095 = ~new_P2_U5804 | ~new_P2_U4386;
  assign new_P2_U6096 = ~new_P2_U3474 | ~new_P2_U3076;
  assign new_P2_U6097 = ~new_P2_U6096 | ~new_P2_U6095;
  assign new_P2_U6098 = ~new_P2_U5755 | ~new_P2_U4253;
  assign new_P2_U6099 = ~new_P2_U3453 | ~new_P2_U3086;
  assign new_P2_U6100 = ~new_P2_U6099 | ~new_P2_U6098;
  assign new_P2_U6101 = ~new_P2_U5762 | ~new_P2_U4272;
  assign new_P2_U6102 = ~new_P2_U3456 | ~new_P2_U3085;
  assign new_P2_U6103 = ~new_P2_U6102 | ~new_P2_U6101;
  assign new_P2_U6104 = ~new_P2_U5790 | ~new_P2_U4348;
  assign new_P2_U6105 = ~new_P2_U3468 | ~new_P2_U3082;
  assign new_P2_U6106 = ~new_P2_U6105 | ~new_P2_U6104;
  assign new_P2_U6107 = ~new_P2_U5825 | ~new_P2_U4443;
  assign new_P2_U6108 = ~new_P2_U3483 | ~new_P2_U3084;
  assign new_P2_U6109 = ~new_P2_U6108 | ~new_P2_U6107;
  assign new_P2_U6110 = ~new_P2_U5811 | ~new_P2_U4405;
  assign new_P2_U6111 = ~new_P2_U3477 | ~new_P2_U3075;
  assign new_P2_U6112 = ~new_P2_U6111 | ~new_P2_U6110;
  assign new_P2_U6113 = ~new_P2_U5783 | ~new_P2_U4329;
  assign new_P2_U6114 = ~new_P2_U3465 | ~new_P2_U3074;
  assign new_P2_U6115 = ~new_P2_U6114 | ~new_P2_U6113;
  assign new_P2_U6116 = ~new_P2_U5741 | ~new_P2_U4215;
  assign new_P2_U6117 = ~new_P2_U3447 | ~new_P2_U3073;
  assign new_P2_U6118 = ~new_P2_U6117 | ~new_P2_U6116;
  assign new_P2_U6119 = ~new_P2_U5748 | ~new_P2_U4234;
  assign new_P2_U6120 = ~new_P2_U3450 | ~new_P2_U3072;
  assign new_P2_U6121 = ~new_P2_U6120 | ~new_P2_U6119;
  assign new_P2_U6122 = ~new_P2_U5734 | ~new_P2_U4196;
  assign new_P2_U6123 = ~new_P2_U3444 | ~new_P2_U3069;
  assign new_P2_U6124 = ~new_P2_U6123 | ~new_P2_U6122;
  assign new_P2_U6125 = ~new_P2_U5720 | ~new_P2_U4158;
  assign new_P2_U6126 = ~new_P2_U3438 | ~new_P2_U3066;
  assign new_P2_U6127 = ~new_P2_U6126 | ~new_P2_U6125;
  assign new_P2_U6128 = ~new_P2_U5713 | ~new_P2_U4134;
  assign new_P2_U6129 = ~new_P2_U3435 | ~new_P2_U3070;
  assign new_P2_U6130 = ~new_P2_U6129 | ~new_P2_U6128;
  assign new_P2_U6131 = ~new_P2_U5818 | ~new_P2_U4424;
  assign new_P2_U6132 = ~new_P2_U3480 | ~new_P2_U3071;
  assign new_P2_U6133 = ~new_P2_U6132 | ~new_P2_U6131;
  assign new_P2_U6134 = ~new_P2_U5830 | ~new_P2_U4462;
  assign new_P2_U6135 = ~new_P2_U3485 | ~new_P2_U3083;
  assign new_P2_U6136 = ~new_P2_U6135 | ~new_P2_U6134;
  assign new_P2_U6137 = ~new_P2_U5727 | ~new_P2_U4177;
  assign new_P2_U6138 = ~new_P2_U3441 | ~new_P2_U3062;
  assign new_P2_U6139 = ~new_P2_U6138 | ~new_P2_U6137;
  assign new_P2_U6140 = ~new_P2_U5776 | ~new_P2_U4310;
  assign new_P2_U6141 = ~new_P2_U3462 | ~new_P2_U3065;
  assign new_P2_U6142 = ~new_P2_U6141 | ~new_P2_U6140;
  assign new_P2_U6143 = ~new_P2_U5769 | ~new_P2_U4291;
  assign new_P2_U6144 = ~new_P2_U3459 | ~new_P2_U3064;
  assign new_P2_U6145 = ~new_P2_U6144 | ~new_P2_U6143;
  assign new_P2_U6146 = ~new_P2_U3957 | ~new_P2_U3078;
  assign new_P2_U6147 = ~new_P2_U3368 | ~new_P2_U4481;
  assign new_P2_U6148 = ~new_P2_U6147 | ~new_P2_U6146;
  assign new_P2_U6149 = ~new_P2_U3940 | ~new_P2_U5156;
  assign new_P2_U6150 = ~new_P2_U3942 | ~new_P2_U3918;
  assign new_P3_R1161_U468 = ~new_P3_U3068 | ~new_P3_R1161_U60;
  assign new_P3_R1161_U467 = ~new_P3_R1161_U270 | ~new_P3_R1161_U465;
  assign new_P3_R1161_U466 = ~new_P3_R1161_U360 | ~new_P3_R1161_U162;
  assign new_P3_R1161_U465 = ~new_P3_R1161_U464 | ~new_P3_R1161_U463;
  assign new_P3_R1161_U464 = ~new_P3_U3443 | ~new_P3_R1161_U76;
  assign new_P3_R1161_U463 = ~new_P3_U3081 | ~new_P3_R1161_U75;
  assign new_P3_R1161_U462 = ~new_P3_R1161_U460 | ~new_P3_R1161_U316;
  assign new_P3_R1161_U461 = ~new_P3_R1161_U359 | ~new_P3_R1161_U91;
  assign new_P3_R1161_U460 = ~new_P3_R1161_U459 | ~new_P3_R1161_U458;
  assign new_P3_R1161_U459 = ~new_P3_U3445 | ~new_P3_R1161_U79;
  assign new_P3_R1161_U458 = ~new_P3_U3080 | ~new_P3_R1161_U78;
  assign new_P3_R1161_U457 = ~new_P3_R1161_U328 | ~new_P3_R1161_U31;
  assign new_P3_R1161_U456 = ~new_P3_R1161_U182 | ~new_P3_R1161_U161;
  assign new_P3_R1161_U455 = ~new_P3_U3907 | ~new_P3_R1161_U90;
  assign new_P3_R1161_U454 = ~new_P3_U3075 | ~new_P3_R1161_U81;
  assign new_P3_R1161_U453 = ~new_P3_R1161_U452 | ~new_P3_R1161_U451;
  assign new_P3_R1161_U452 = ~new_P3_U3906 | ~new_P3_R1161_U55;
  assign new_P3_R1161_U451 = ~new_P3_U3074 | ~new_P3_R1161_U54;
  assign new_P3_R1161_U450 = ~new_P3_U3906 | ~new_P3_R1161_U55;
  assign new_P3_R1161_U449 = ~new_P3_U3074 | ~new_P3_R1161_U54;
  assign new_P3_U3013 = new_P3_U3380 & new_P3_U5450;
  assign new_P3_U3014 = new_P3_U3380 & new_P3_U3379;
  assign new_P3_U3015 = new_P3_U5453 & new_P3_U3379;
  assign new_P3_U3016 = new_P3_U5453 & new_P3_U5450;
  assign new_P3_U3017 = new_P3_U3874 & new_P3_U5447;
  assign new_P3_U3018 = new_P3_U3587 & new_P3_U3582;
  assign new_P3_U3019 = new_P3_U3381 & new_P3_U3382;
  assign new_P3_U3020 = new_P3_U5462 & new_P3_U3381;
  assign new_P3_U3021 = new_P3_U5459 & new_P3_U3382;
  assign new_P3_U3022 = new_P3_U5462 & new_P3_U5459;
  assign new_P3_U3023 = new_P3_U3046 & P3_STATE_REG;
  assign new_P3_U3024 = new_P3_U3696 & new_P3_U3366;
  assign new_P3_U3025 = new_P3_U3911 & new_P3_U4073;
  assign new_P3_U3026 = new_P3_U3015 & new_P3_U5447;
  assign new_P3_U3027 = new_P3_U3297 & P3_STATE_REG;
  assign new_P3_U3028 = new_P3_U3886 & new_P3_U3912;
  assign new_P3_U3029 = new_P3_U3912 & new_P3_U3365;
  assign new_P3_U3030 = new_P3_U3693 & new_P3_U3912;
  assign new_P3_U3031 = new_P3_U3890 & new_P3_U3023;
  assign new_P3_U3032 = new_P3_U3895 & new_P3_U4073;
  assign new_P3_U3033 = new_P3_U3911 & new_P3_U4089;
  assign new_P3_U3034 = new_P3_U3912 & new_P3_U3025;
  assign new_P3_U3035 = new_P3_U3023 & new_P3_U4989;
  assign new_P3_U3036 = new_P3_U3895 & new_P3_U4089;
  assign new_P3_U3037 = new_P3_U5468 & new_P3_U4754;
  assign new_P3_U3038 = new_P3_U3024 & new_P3_U5468;
  assign new_P3_U3039 = new_P3_U5465 & new_P3_U4754;
  assign new_P3_U3040 = new_P3_U3892 & new_P3_U4754;
  assign new_P3_U3041 = new_P3_U3024 & new_P3_U3892;
  assign new_P3_U3042 = new_P3_U3023 & new_P3_U3366;
  assign new_P3_U3043 = new_P3_U3023 & new_P3_U3365;
  assign new_P3_U3044 = new_P3_U5004 & P3_STATE_REG;
  assign new_P3_U3045 = new_P3_U3023 & new_P3_U5006;
  assign new_P3_U3046 = new_P3_U5440 & new_P3_U3362;
  assign new_P3_U3047 = new_P3_U3692 & new_P3_U3018;
  assign new_P3_U3048 = new_P3_U3691 & new_P3_U3018;
  assign new_P3_U3049 = new_P3_U4749 & new_P3_U4748;
  assign new_P3_U3050 = new_P3_U4759 & P3_STATE_REG;
  assign new_P3_U3051 = n3844 & new_P3_U4761;
  assign new_P3_U3052 = ~new_P3_U4538 | ~new_P3_U4535 | ~new_P3_U4536 | ~new_P3_U4537;
  assign new_P3_U3053 = ~new_P3_U4553 | ~new_P3_U4554 | ~new_P3_U4556 | ~new_P3_U4555;
  assign new_P3_U3054 = ~new_P3_U4571 | ~new_P3_U4572 | ~new_P3_U4574 | ~new_P3_U4573;
  assign new_P3_U3055 = ~new_P3_U4609 | ~new_P3_U4610 | ~new_P3_U4612 | ~new_P3_U4611;
  assign new_P3_U3056 = ~new_P3_U4517 | ~new_P3_U4518 | ~new_P3_U4520 | ~new_P3_U4519;
  assign new_P3_U3057 = ~new_P3_U4499 | ~new_P3_U4500 | ~new_P3_U4502 | ~new_P3_U4501;
  assign new_P3_U3058 = ~new_P3_U4589 | ~new_P3_U4590 | ~new_P3_U4592 | ~new_P3_U4591;
  assign new_P3_U3059 = ~new_P3_U4121 | ~new_P3_U4122 | ~new_P3_U4124 | ~new_P3_U4123;
  assign new_P3_U3060 = ~new_P3_U4445 | ~new_P3_U4446 | ~new_P3_U4448 | ~new_P3_U4447;
  assign new_P3_U3061 = ~new_P3_U4229 | ~new_P3_U4230 | ~new_P3_U4232 | ~new_P3_U4231;
  assign new_P3_U3062 = ~new_P3_U4247 | ~new_P3_U4248 | ~new_P3_U4250 | ~new_P3_U4249;
  assign new_P3_U3063 = ~new_P3_U4103 | ~new_P3_U4104 | ~new_P3_U4106 | ~new_P3_U4105;
  assign new_P3_U3064 = ~new_P3_U4481 | ~new_P3_U4482 | ~new_P3_U4484 | ~new_P3_U4483;
  assign new_P3_U3065 = ~new_P3_U4463 | ~new_P3_U4464 | ~new_P3_U4466 | ~new_P3_U4465;
  assign new_P3_U3066 = ~new_P3_U4139 | ~new_P3_U4140 | ~new_P3_U4142 | ~new_P3_U4141;
  assign new_P3_U3067 = ~new_P3_U4078 | ~new_P3_U4079 | ~new_P3_U4081 | ~new_P3_U4080;
  assign new_P3_U3068 = ~new_P3_U4355 | ~new_P3_U4356 | ~new_P3_U4358 | ~new_P3_U4357;
  assign new_P3_U3069 = ~new_P3_U4175 | ~new_P3_U4176 | ~new_P3_U4178 | ~new_P3_U4177;
  assign new_P3_U3070 = ~new_P3_U4157 | ~new_P3_U4158 | ~new_P3_U4160 | ~new_P3_U4159;
  assign new_P3_U3071 = ~new_P3_U4265 | ~new_P3_U4266 | ~new_P3_U4268 | ~new_P3_U4267;
  assign new_P3_U3072 = ~new_P3_U4337 | ~new_P3_U4338 | ~new_P3_U4340 | ~new_P3_U4339;
  assign new_P3_U3073 = ~new_P3_U4319 | ~new_P3_U4320 | ~new_P3_U4322 | ~new_P3_U4321;
  assign new_P3_U3074 = ~new_P3_U4427 | ~new_P3_U4428 | ~new_P3_U4430 | ~new_P3_U4429;
  assign new_P3_U3075 = ~new_P3_U4409 | ~new_P3_U4410 | ~new_P3_U4412 | ~new_P3_U4411;
  assign new_P3_U3076 = ~new_P3_U4083 | ~new_P3_U4084 | ~new_P3_U4086 | ~new_P3_U4085;
  assign new_P3_U3077 = ~new_P3_U4059 | ~new_P3_U4060 | ~new_P3_U4062 | ~new_P3_U4061;
  assign new_P3_U3078 = ~new_P3_U4301 | ~new_P3_U4302 | ~new_P3_U4304 | ~new_P3_U4303;
  assign new_P3_U3079 = ~new_P3_U4283 | ~new_P3_U4284 | ~new_P3_U4286 | ~new_P3_U4285;
  assign new_P3_U3080 = ~new_P3_U4391 | ~new_P3_U4392 | ~new_P3_U4394 | ~new_P3_U4393;
  assign new_P3_U3081 = ~new_P3_U4373 | ~new_P3_U4374 | ~new_P3_U4376 | ~new_P3_U4375;
  assign new_P3_U3082 = ~new_P3_U4211 | ~new_P3_U4212 | ~new_P3_U4214 | ~new_P3_U4213;
  assign new_P3_U3083 = ~new_P3_U4193 | ~new_P3_U4194 | ~new_P3_U4196 | ~new_P3_U4195;
  assign new_P3_U3084 = ~new_P3_U5341 | ~new_P3_U5340;
  assign new_P3_U3085 = ~new_P3_U5343 | ~new_P3_U5342;
  assign new_P3_U3086 = ~new_P3_U5348 | ~new_P3_U5349 | ~new_P3_U5347;
  assign new_P3_U3087 = ~new_P3_U5351 | ~new_P3_U5352 | ~new_P3_U5350;
  assign new_P3_U3088 = ~new_P3_U5354 | ~new_P3_U5355 | ~new_P3_U5353;
  assign new_P3_U3089 = ~new_P3_U5357 | ~new_P3_U5358 | ~new_P3_U5356;
  assign new_P3_U3090 = ~new_P3_U5360 | ~new_P3_U5361 | ~new_P3_U5359;
  assign new_P3_U3091 = ~new_P3_U5363 | ~new_P3_U5364 | ~new_P3_U5362;
  assign new_P3_U3092 = ~new_P3_U5366 | ~new_P3_U5367 | ~new_P3_U5365;
  assign new_P3_U3093 = ~new_P3_U5369 | ~new_P3_U5370 | ~new_P3_U5368;
  assign new_P3_U3094 = ~new_P3_U5372 | ~new_P3_U5373 | ~new_P3_U5371;
  assign new_P3_U3095 = ~new_P3_U5375 | ~new_P3_U5376 | ~new_P3_U5374;
  assign new_P3_U3096 = ~new_P3_U5380 | ~new_P3_U5381 | ~new_P3_U5382;
  assign new_P3_U3097 = ~new_P3_U5383 | ~new_P3_U5384 | ~new_P3_U5385;
  assign new_P3_U3098 = ~new_P3_U5386 | ~new_P3_U5387 | ~new_P3_U5388;
  assign new_P3_U3099 = ~new_P3_U5389 | ~new_P3_U5390 | ~new_P3_U5391;
  assign new_P3_U3100 = ~new_P3_U5392 | ~new_P3_U5393 | ~new_P3_U5394;
  assign new_P3_U3101 = ~new_P3_U5395 | ~new_P3_U5396 | ~new_P3_U5397;
  assign new_P3_U3102 = ~new_P3_U5400 | ~new_P3_U5399 | ~new_P3_U5398;
  assign new_P3_U3103 = ~new_P3_U5403 | ~new_P3_U5402 | ~new_P3_U5401;
  assign new_P3_U3104 = ~new_P3_U5406 | ~new_P3_U5405 | ~new_P3_U5404;
  assign new_P3_U3105 = ~new_P3_U5409 | ~new_P3_U5408 | ~new_P3_U5407;
  assign new_P3_U3106 = ~new_P3_U5324 | ~new_P3_U5323 | ~new_P3_U5322;
  assign new_P3_U3107 = ~new_P3_U5327 | ~new_P3_U5326 | ~new_P3_U5325;
  assign new_P3_U3108 = ~new_P3_U5330 | ~new_P3_U5329 | ~new_P3_U5328;
  assign new_P3_U3109 = ~new_P3_U5333 | ~new_P3_U5332 | ~new_P3_U5331;
  assign new_P3_U3110 = ~new_P3_U5336 | ~new_P3_U5335 | ~new_P3_U5334;
  assign new_P3_U3111 = ~new_P3_U5339 | ~new_P3_U5338 | ~new_P3_U5337;
  assign new_P3_U3112 = ~new_P3_U5346 | ~new_P3_U5345 | ~new_P3_U5344;
  assign new_P3_U3113 = ~new_P3_U5379 | ~new_P3_U5378 | ~new_P3_U5377;
  assign new_P3_U3114 = ~new_P3_U5412 | ~new_P3_U5411 | ~new_P3_U5410;
  assign new_P3_U3115 = ~new_P3_U5414 | ~new_P3_U5413;
  assign new_P3_U3116 = ~new_P3_U5271 | ~new_P3_U5270;
  assign new_P3_U3117 = ~new_P3_U5273 | ~new_P3_U5272;
  assign new_P3_U3118 = ~new_P3_U5276 | ~new_P3_U5277 | ~new_P3_U3375;
  assign new_P3_U3119 = ~new_P3_U5278 | ~new_P3_U5279 | ~new_P3_U3375;
  assign new_P3_U3120 = ~new_P3_U5280 | ~new_P3_U5281 | ~new_P3_U3375;
  assign new_P3_U3121 = ~new_P3_U5282 | ~new_P3_U5283 | ~new_P3_U3375;
  assign new_P3_U3122 = ~new_P3_U5284 | ~new_P3_U5285 | ~new_P3_U3375;
  assign new_P3_U3123 = ~new_P3_U5286 | ~new_P3_U5287 | ~new_P3_U3375;
  assign new_P3_U3124 = ~new_P3_U5288 | ~new_P3_U5289 | ~new_P3_U3375;
  assign new_P3_U3125 = ~new_P3_U5290 | ~new_P3_U5291 | ~new_P3_U3375;
  assign new_P3_U3126 = ~new_P3_U5292 | ~new_P3_U5293 | ~new_P3_U3375;
  assign new_P3_U3127 = ~new_P3_U5294 | ~new_P3_U5295 | ~new_P3_U3375;
  assign new_P3_U3128 = ~new_P3_U5298 | ~new_P3_U5299 | ~new_P3_U3375;
  assign new_P3_U3129 = ~new_P3_U5300 | ~new_P3_U5301 | ~new_P3_U3375;
  assign new_P3_U3130 = ~new_P3_U5302 | ~new_P3_U5303 | ~new_P3_U3375;
  assign new_P3_U3131 = ~new_P3_U5304 | ~new_P3_U5305 | ~new_P3_U3375;
  assign new_P3_U3132 = ~new_P3_U5306 | ~new_P3_U5307 | ~new_P3_U3375;
  assign new_P3_U3133 = ~new_P3_U5308 | ~new_P3_U5309 | ~new_P3_U3375;
  assign new_P3_U3134 = ~new_P3_U3825 | ~new_P3_U5311;
  assign new_P3_U3135 = ~new_P3_U3826 | ~new_P3_U5313;
  assign new_P3_U3136 = ~new_P3_U3827 | ~new_P3_U5315;
  assign new_P3_U3137 = ~new_P3_U3828 | ~new_P3_U5317;
  assign new_P3_U3138 = ~new_P3_U3817 | ~new_P3_U5259;
  assign new_P3_U3139 = ~new_P3_U3818 | ~new_P3_U5261;
  assign new_P3_U3140 = ~new_P3_U3819 | ~new_P3_U5263;
  assign new_P3_U3141 = ~new_P3_U3820 | ~new_P3_U5265;
  assign new_P3_U3142 = ~new_P3_U3821 | ~new_P3_U5267;
  assign new_P3_U3143 = ~new_P3_U3822 | ~new_P3_U5269;
  assign new_P3_U3144 = ~new_P3_U3823 | ~new_P3_U5275;
  assign new_P3_U3145 = ~new_P3_U3824 | ~new_P3_U5297;
  assign new_P3_U3146 = ~new_P3_U3829 | ~new_P3_U5319;
  assign new_P3_U3147 = ~new_P3_U3830 | ~new_P3_U5321;
  assign new_P3_U3148 = ~new_P3_U3375 | ~new_P3_U3385 | ~new_P3_U5453;
  assign new_P3_U3149 = ~new_P3_U3813 | ~new_P3_U3013;
  assign n3839 = ~new_P3_U3812 | ~new_P3_U5253;
  assign n3834 = ~P3_STATE_REG;
  assign new_P3_U3152 = ~new_P3_U3359 | ~new_P3_U5944 | ~new_P3_U5943;
  assign n3829 = ~new_P3_U5250 | ~new_P3_U3811 | ~new_P3_U5249 | ~new_P3_U5248;
  assign n3824 = ~new_P3_U5241 | ~new_P3_U5239 | ~new_P3_U5240 | ~new_P3_U3810;
  assign n3819 = ~new_P3_U5232 | ~new_P3_U3809 | ~new_P3_U5231 | ~new_P3_U5230;
  assign n3814 = ~new_P3_U5223 | ~new_P3_U5221 | ~new_P3_U5222 | ~new_P3_U3808;
  assign n3809 = ~new_P3_U5214 | ~new_P3_U3807 | ~new_P3_U5213 | ~new_P3_U5212;
  assign n3804 = ~new_P3_U3806 | ~new_P3_U3805 | ~new_P3_U5204;
  assign n3799 = ~new_P3_U5196 | ~new_P3_U5194 | ~new_P3_U5195 | ~new_P3_U3804;
  assign n3794 = ~new_P3_U5187 | ~new_P3_U5185 | ~new_P3_U5186 | ~new_P3_U3803;
  assign n3789 = ~new_P3_U5178 | ~new_P3_U3802 | ~new_P3_U5177 | ~new_P3_U5176;
  assign n3784 = ~new_P3_U3801 | ~new_P3_U3800 | ~new_P3_U5168;
  assign n3779 = ~new_P3_U5160 | ~new_P3_U5158 | ~new_P3_U5159 | ~new_P3_U3799;
  assign n3774 = ~new_P3_U5151 | ~new_P3_U3798 | ~new_P3_U5150 | ~new_P3_U5149;
  assign n3769 = ~new_P3_U5142 | ~new_P3_U5140 | ~new_P3_U5141 | ~new_P3_U3797;
  assign n3764 = ~new_P3_U5133 | ~new_P3_U3796 | ~new_P3_U5132 | ~new_P3_U5131;
  assign n3759 = ~new_P3_U5124 | ~new_P3_U3795 | ~new_P3_U5123 | ~new_P3_U5122;
  assign n3754 = ~new_P3_U5115 | ~new_P3_U3794 | ~new_P3_U5114 | ~new_P3_U5113;
  assign n3749 = ~new_P3_U5106 | ~new_P3_U5104 | ~new_P3_U5105 | ~new_P3_U3793;
  assign n3744 = ~new_P3_U3792 | ~new_P3_U3791 | ~new_P3_U5096;
  assign n3739 = ~new_P3_U5088 | ~new_P3_U3790 | ~new_P3_U5087 | ~new_P3_U5086;
  assign n3734 = ~new_P3_U5079 | ~new_P3_U3789;
  assign n3729 = ~new_P3_U5072 | ~new_P3_U5070 | ~new_P3_U5071 | ~new_P3_U3786;
  assign n3724 = ~new_P3_U5063 | ~new_P3_U3785 | ~new_P3_U5062 | ~new_P3_U5061;
  assign n3719 = ~new_P3_U5054 | ~new_P3_U5052 | ~new_P3_U5053 | ~new_P3_U3784;
  assign n3714 = ~new_P3_U5045 | ~new_P3_U3783 | ~new_P3_U5044 | ~new_P3_U5043;
  assign n3709 = ~new_P3_U3782 | ~new_P3_U3781 | ~new_P3_U5035;
  assign n3704 = ~new_P3_U5027 | ~new_P3_U3780 | ~new_P3_U5026 | ~new_P3_U5025;
  assign n3699 = ~new_P3_U5018 | ~new_P3_U3779 | ~new_P3_U5017 | ~new_P3_U5016;
  assign n3694 = ~new_P3_U5009 | ~new_P3_U5007 | ~new_P3_U5008 | ~new_P3_U3778;
  assign n3689 = ~new_P3_U4996 | ~new_P3_U3777 | ~new_P3_U4995 | ~new_P3_U4994;
  assign n3519 = ~new_P3_U4973 | ~new_P3_U3756;
  assign n3514 = ~new_P3_U4962 | ~new_P3_U3753;
  assign n3509 = ~new_P3_U4951 | ~new_P3_U3750;
  assign n3504 = ~new_P3_U3747 | ~new_P3_U4941 | ~new_P3_U4940;
  assign n3499 = ~new_P3_U3744 | ~new_P3_U4930 | ~new_P3_U4929;
  assign n3494 = ~new_P3_U4916 | ~new_P3_U3743 | ~new_P3_U4918 | ~new_P3_U3741;
  assign n3489 = ~new_P3_U4905 | ~new_P3_U4907 | ~new_P3_U3738;
  assign n3484 = ~new_P3_U4896 | ~new_P3_U3735;
  assign n3479 = ~new_P3_U4885 | ~new_P3_U3732;
  assign n3474 = ~new_P3_U4874 | ~new_P3_U3729;
  assign n3469 = ~new_P3_U4863 | ~new_P3_U3726;
  assign n3464 = ~new_P3_U4852 | ~new_P3_U3723;
  assign n3459 = ~new_P3_U4841 | ~new_P3_U3720;
  assign n3454 = ~new_P3_U4830 | ~new_P3_U3717;
  assign n3449 = ~new_P3_U4819 | ~new_P3_U3714;
  assign n3444 = ~new_P3_U4808 | ~new_P3_U3711;
  assign n3439 = ~new_P3_U4797 | ~new_P3_U3708;
  assign n3434 = ~new_P3_U4786 | ~new_P3_U3705;
  assign n3429 = ~new_P3_U4775 | ~new_P3_U3702;
  assign n3424 = ~new_P3_U4764 | ~new_P3_U3699;
  assign n3419 = ~new_P3_U4752 | ~new_P3_U4753 | ~new_P3_U3049;
  assign n3414 = ~new_P3_U4750 | ~new_P3_U4751 | ~new_P3_U3049;
  assign n3409 = ~new_P3_U3866 | ~new_P3_U4745 | ~new_P3_U4746 | ~new_P3_U4747;
  assign n3404 = ~new_P3_U3865 | ~new_P3_U4742 | ~new_P3_U4744 | ~new_P3_U4743 | ~new_P3_U4741;
  assign n3399 = ~new_P3_U3864 | ~new_P3_U4738 | ~new_P3_U4740 | ~new_P3_U4739 | ~new_P3_U4737;
  assign n3394 = ~new_P3_U3863 | ~new_P3_U4734 | ~new_P3_U4736 | ~new_P3_U4735 | ~new_P3_U4733;
  assign n3389 = ~new_P3_U3862 | ~new_P3_U4730 | ~new_P3_U4732 | ~new_P3_U4731 | ~new_P3_U4729;
  assign n3384 = ~new_P3_U3861 | ~new_P3_U4726 | ~new_P3_U4728 | ~new_P3_U4727 | ~new_P3_U4725;
  assign n3379 = ~new_P3_U3860 | ~new_P3_U4722 | ~new_P3_U4724 | ~new_P3_U4723 | ~new_P3_U4721;
  assign n3374 = ~new_P3_U3859 | ~new_P3_U4718 | ~new_P3_U4720 | ~new_P3_U4719 | ~new_P3_U4717;
  assign n3369 = ~new_P3_U3858 | ~new_P3_U4714 | ~new_P3_U4716 | ~new_P3_U4715 | ~new_P3_U4713;
  assign n3364 = ~new_P3_U3857 | ~new_P3_U4710 | ~new_P3_U4712 | ~new_P3_U4711 | ~new_P3_U4709;
  assign n3359 = ~new_P3_U3856 | ~new_P3_U4706 | ~new_P3_U4708 | ~new_P3_U4707 | ~new_P3_U4705;
  assign n3354 = ~new_P3_U3855 | ~new_P3_U4702 | ~new_P3_U4704 | ~new_P3_U4703 | ~new_P3_U4701;
  assign n3349 = ~new_P3_U3854 | ~new_P3_U4698 | ~new_P3_U4700 | ~new_P3_U4699 | ~new_P3_U4697;
  assign n3344 = ~new_P3_U3853 | ~new_P3_U4694 | ~new_P3_U4696 | ~new_P3_U4695 | ~new_P3_U4693;
  assign n3339 = ~new_P3_U3852 | ~new_P3_U4690 | ~new_P3_U4692 | ~new_P3_U4691 | ~new_P3_U4689;
  assign n3334 = ~new_P3_U3851 | ~new_P3_U4686 | ~new_P3_U4688 | ~new_P3_U4687 | ~new_P3_U4685;
  assign n3329 = ~new_P3_U3850 | ~new_P3_U4681 | ~new_P3_U4683 | ~new_P3_U4684 | ~new_P3_U4682;
  assign n3324 = ~new_P3_U3849 | ~new_P3_U4677 | ~new_P3_U4678 | ~new_P3_U4680 | ~new_P3_U4679;
  assign n3319 = ~new_P3_U3848 | ~new_P3_U4673 | ~new_P3_U4675 | ~new_P3_U4676 | ~new_P3_U4674;
  assign n3314 = ~new_P3_U3847 | ~new_P3_U4669 | ~new_P3_U4670 | ~new_P3_U4672 | ~new_P3_U4671;
  assign n3309 = ~new_P3_U4668 | ~new_P3_U3846 | ~new_P3_U4667 | ~new_P3_U4666 | ~new_P3_U4665;
  assign n3304 = ~new_P3_U4664 | ~new_P3_U3845 | ~new_P3_U4663 | ~new_P3_U4662 | ~new_P3_U4661;
  assign n3299 = ~new_P3_U4660 | ~new_P3_U3844 | ~new_P3_U4659 | ~new_P3_U4658 | ~new_P3_U4657;
  assign n3294 = ~new_P3_U4656 | ~new_P3_U3843 | ~new_P3_U4655 | ~new_P3_U4654 | ~new_P3_U4653;
  assign n3289 = ~new_P3_U4652 | ~new_P3_U3842 | ~new_P3_U4651 | ~new_P3_U4650 | ~new_P3_U4649;
  assign n3284 = ~new_P3_U4648 | ~new_P3_U3841 | ~new_P3_U4647 | ~new_P3_U4646 | ~new_P3_U4645;
  assign n3279 = ~new_P3_U4644 | ~new_P3_U3840 | ~new_P3_U4643 | ~new_P3_U4642 | ~new_P3_U4641;
  assign n3274 = ~new_P3_U4640 | ~new_P3_U3839 | ~new_P3_U4639 | ~new_P3_U4638 | ~new_P3_U4637;
  assign n3269 = ~new_P3_U4636 | ~new_P3_U3838 | ~new_P3_U4635 | ~new_P3_U4634 | ~new_P3_U4633;
  assign n3264 = ~new_P3_U4632 | ~new_P3_U3837 | ~new_P3_U4631 | ~new_P3_U4630 | ~new_P3_U4629;
  assign n2939 = P3_D_REG_31_ & new_P3_U3832;
  assign n2934 = P3_D_REG_30_ & new_P3_U3832;
  assign n2929 = P3_D_REG_29_ & new_P3_U3832;
  assign n2924 = P3_D_REG_28_ & new_P3_U3832;
  assign n2919 = P3_D_REG_27_ & new_P3_U3832;
  assign n2914 = P3_D_REG_26_ & new_P3_U3832;
  assign n2909 = P3_D_REG_25_ & new_P3_U3832;
  assign n2904 = P3_D_REG_24_ & new_P3_U3832;
  assign n2899 = P3_D_REG_23_ & new_P3_U3832;
  assign n2894 = P3_D_REG_22_ & new_P3_U3832;
  assign n2889 = P3_D_REG_21_ & new_P3_U3832;
  assign n2884 = P3_D_REG_20_ & new_P3_U3832;
  assign n2879 = P3_D_REG_19_ & new_P3_U3832;
  assign n2874 = P3_D_REG_18_ & new_P3_U3832;
  assign n2869 = P3_D_REG_17_ & new_P3_U3832;
  assign n2864 = P3_D_REG_16_ & new_P3_U3832;
  assign n2859 = P3_D_REG_15_ & new_P3_U3832;
  assign n2854 = P3_D_REG_14_ & new_P3_U3832;
  assign n2849 = P3_D_REG_13_ & new_P3_U3832;
  assign n2844 = P3_D_REG_12_ & new_P3_U3832;
  assign n2839 = P3_D_REG_11_ & new_P3_U3832;
  assign n2834 = P3_D_REG_10_ & new_P3_U3832;
  assign n2829 = P3_D_REG_9_ & new_P3_U3832;
  assign n2824 = P3_D_REG_8_ & new_P3_U3832;
  assign n2819 = P3_D_REG_7_ & new_P3_U3832;
  assign n2814 = P3_D_REG_6_ & new_P3_U3832;
  assign n2809 = P3_D_REG_5_ & new_P3_U3832;
  assign n2804 = P3_D_REG_4_ & new_P3_U3832;
  assign n2799 = P3_D_REG_3_ & new_P3_U3832;
  assign n2794 = P3_D_REG_2_ & new_P3_U3832;
  assign n2779 = ~new_P3_U4015 | ~new_P3_U4016 | ~new_P3_U4017;
  assign n2774 = ~new_P3_U4012 | ~new_P3_U4013 | ~new_P3_U4014;
  assign n2769 = ~new_P3_U4009 | ~new_P3_U4010 | ~new_P3_U4011;
  assign n2764 = ~new_P3_U4006 | ~new_P3_U4007 | ~new_P3_U4008;
  assign n2759 = ~new_P3_U4003 | ~new_P3_U4004 | ~new_P3_U4005;
  assign n2754 = ~new_P3_U4000 | ~new_P3_U4001 | ~new_P3_U4002;
  assign n2749 = ~new_P3_U3997 | ~new_P3_U3998 | ~new_P3_U3999;
  assign n2744 = ~new_P3_U3994 | ~new_P3_U3995 | ~new_P3_U3996;
  assign n2739 = ~new_P3_U3991 | ~new_P3_U3992 | ~new_P3_U3993;
  assign n2734 = ~new_P3_U3988 | ~new_P3_U3989 | ~new_P3_U3990;
  assign n2729 = ~new_P3_U3985 | ~new_P3_U3986 | ~new_P3_U3987;
  assign n2724 = ~new_P3_U3982 | ~new_P3_U3983 | ~new_P3_U3984;
  assign n2719 = ~new_P3_U3979 | ~new_P3_U3980 | ~new_P3_U3981;
  assign n2714 = ~new_P3_U3976 | ~new_P3_U3977 | ~new_P3_U3978;
  assign n2709 = ~new_P3_U3973 | ~new_P3_U3974 | ~new_P3_U3975;
  assign n2704 = ~new_P3_U3970 | ~new_P3_U3971 | ~new_P3_U3972;
  assign n2699 = ~new_P3_U3967 | ~new_P3_U3968 | ~new_P3_U3969;
  assign n2694 = ~new_P3_U3964 | ~new_P3_U3965 | ~new_P3_U3966;
  assign n2689 = ~new_P3_U3961 | ~new_P3_U3962 | ~new_P3_U3963;
  assign n2684 = ~new_P3_U3958 | ~new_P3_U3959 | ~new_P3_U3960;
  assign n2679 = ~new_P3_U3955 | ~new_P3_U3956 | ~new_P3_U3957;
  assign n2674 = ~new_P3_U3952 | ~new_P3_U3953 | ~new_P3_U3954;
  assign n2669 = ~new_P3_U3949 | ~new_P3_U3950 | ~new_P3_U3951;
  assign n2664 = ~new_P3_U3946 | ~new_P3_U3947 | ~new_P3_U3948;
  assign n2659 = ~new_P3_U3943 | ~new_P3_U3944 | ~new_P3_U3945;
  assign n2654 = ~new_P3_U3940 | ~new_P3_U3941 | ~new_P3_U3942;
  assign n2649 = ~new_P3_U3937 | ~new_P3_U3938 | ~new_P3_U3939;
  assign n2644 = ~new_P3_U3934 | ~new_P3_U3935 | ~new_P3_U3936;
  assign n2639 = ~new_P3_U3931 | ~new_P3_U3932 | ~new_P3_U3933;
  assign n2634 = ~new_P3_U3928 | ~new_P3_U3929 | ~new_P3_U3930;
  assign n2629 = ~new_P3_U3925 | ~new_P3_U3926 | ~new_P3_U3927;
  assign n2624 = ~new_P3_U3922 | ~new_P3_U3923 | ~new_P3_U3924;
  assign n3684 = new_P3_U3775 & new_P3_U5421;
  assign new_P3_U3297 = ~P3_STATE_REG | ~new_P3_U3831;
  assign new_P3_U3298 = ~P3_B_REG;
  assign new_P3_U3299 = ~new_P3_U3374 | ~new_P3_U5431;
  assign new_P3_U3300 = ~new_P3_U3374 | ~new_P3_U4018;
  assign new_P3_U3301 = ~new_P3_U3013 | ~new_P3_U5447;
  assign new_P3_U3302 = ~new_P3_U3014 | ~new_P3_U5456;
  assign new_P3_U3303 = ~new_P3_U3588 | ~new_P3_U3018;
  assign new_P3_U3304 = ~new_P3_U3589 | ~new_P3_U3018;
  assign new_P3_U3305 = ~new_P3_U3014 | ~new_P3_U5447;
  assign new_P3_U3306 = ~new_P3_U3014 | ~new_P3_U3378;
  assign new_P3_U3307 = ~new_P3_U3013 | ~new_P3_U3378;
  assign new_P3_U3308 = ~new_P3_U3378 | ~new_P3_U3385 | ~new_P3_U3379;
  assign new_P3_U3309 = ~new_P3_U3378 | ~new_P3_U5450 | ~new_P3_U3385;
  assign new_P3_U3310 = ~new_P3_U5456 | ~new_P3_U3013;
  assign new_P3_U3311 = ~new_P3_U3878 | ~new_P3_U5447;
  assign new_P3_U3312 = ~new_P3_U3016 | ~new_P3_U3385;
  assign new_P3_U3313 = ~new_P3_U3385 | ~new_P3_U3380;
  assign new_P3_U3314 = ~new_P3_U3575 | ~new_P3_U3576 | ~new_P3_U4071 | ~new_P3_U4070 | ~new_P3_U4069;
  assign new_P3_U3315 = ~new_P3_U3592 | ~new_P3_U3590 | ~new_P3_U4091 | ~new_P3_U4090;
  assign new_P3_U3316 = ~new_P3_U3596 | ~new_P3_U3594 | ~new_P3_U4109 | ~new_P3_U4108;
  assign new_P3_U3317 = ~new_P3_U3600 | ~new_P3_U3598 | ~new_P3_U4127 | ~new_P3_U4126;
  assign new_P3_U3318 = ~new_P3_U3603 | ~new_P3_U4147 | ~new_P3_U4146 | ~new_P3_U4145 | ~new_P3_U4144;
  assign new_P3_U3319 = ~new_P3_U3606 | ~new_P3_U4165 | ~new_P3_U4164 | ~new_P3_U4163 | ~new_P3_U4162;
  assign new_P3_U3320 = ~new_P3_U3609 | ~new_P3_U4183 | ~new_P3_U4182 | ~new_P3_U4181 | ~new_P3_U4180;
  assign new_P3_U3321 = ~new_P3_U3612 | ~new_P3_U4201 | ~new_P3_U4200 | ~new_P3_U4199 | ~new_P3_U4198;
  assign new_P3_U3322 = ~new_P3_U3615 | ~new_P3_U4219 | ~new_P3_U4218 | ~new_P3_U4217 | ~new_P3_U4216;
  assign new_P3_U3323 = ~new_P3_U3619 | ~new_P3_U3617 | ~new_P3_U4235 | ~new_P3_U4234;
  assign new_P3_U3324 = ~new_P3_U3623 | ~new_P3_U3621 | ~new_P3_U4253 | ~new_P3_U4252;
  assign new_P3_U3325 = ~new_P3_U3626 | ~new_P3_U4273 | ~new_P3_U4272 | ~new_P3_U4271 | ~new_P3_U4270;
  assign new_P3_U3326 = ~new_P3_U3630 | ~new_P3_U3628 | ~new_P3_U4289 | ~new_P3_U4288;
  assign new_P3_U3327 = ~new_P3_U3634 | ~new_P3_U3632 | ~new_P3_U4307 | ~new_P3_U4306;
  assign new_P3_U3328 = ~new_P3_U3637 | ~new_P3_U4327 | ~new_P3_U4326 | ~new_P3_U4325 | ~new_P3_U4324;
  assign new_P3_U3329 = ~new_P3_U3640 | ~new_P3_U4345 | ~new_P3_U4344 | ~new_P3_U4343 | ~new_P3_U4342;
  assign new_P3_U3330 = ~new_P3_U3643 | ~new_P3_U4363 | ~new_P3_U4362 | ~new_P3_U4361 | ~new_P3_U4360;
  assign new_P3_U3331 = ~new_P3_U3647 | ~new_P3_U3645 | ~new_P3_U4379 | ~new_P3_U4378;
  assign new_P3_U3332 = ~new_P3_U3650 | ~new_P3_U4399 | ~new_P3_U4398 | ~new_P3_U4397 | ~new_P3_U4396;
  assign new_P3_U3333 = ~new_P3_U3653 | ~new_P3_U4417 | ~new_P3_U4416 | ~new_P3_U4415 | ~new_P3_U4414;
  assign new_P3_U3334 = ~new_U49 | ~new_P3_U3833;
  assign new_P3_U3335 = ~new_P3_U3656 | ~new_P3_U4435 | ~new_P3_U4434 | ~new_P3_U4433 | ~new_P3_U4432;
  assign new_P3_U3336 = ~new_U48 | ~new_P3_U3833;
  assign new_P3_U3337 = ~new_P3_U3659 | ~new_P3_U4453 | ~new_P3_U4452 | ~new_P3_U4451 | ~new_P3_U4450;
  assign new_P3_U3338 = ~new_U47 | ~new_P3_U3833;
  assign new_P3_U3339 = ~new_P3_U3662 | ~new_P3_U4471 | ~new_P3_U4470 | ~new_P3_U4469 | ~new_P3_U4468;
  assign new_P3_U3340 = ~new_U46 | ~new_P3_U3833;
  assign new_P3_U3341 = ~new_P3_U3665 | ~new_P3_U4489 | ~new_P3_U4488 | ~new_P3_U4487 | ~new_P3_U4486;
  assign new_P3_U3342 = ~new_U45 | ~new_P3_U3833;
  assign new_P3_U3343 = ~new_P3_U3669 | ~new_P3_U3667 | ~new_P3_U4505 | ~new_P3_U4504;
  assign new_P3_U3344 = ~new_U44 | ~new_P3_U3833;
  assign new_P3_U3345 = ~new_P3_U3673 | ~new_P3_U3671 | ~new_P3_U4523 | ~new_P3_U4522;
  assign new_P3_U3346 = ~new_U43 | ~new_P3_U3833;
  assign new_P3_U3347 = ~new_P3_U3677 | ~new_P3_U3675 | ~new_P3_U4541 | ~new_P3_U4540;
  assign new_P3_U3348 = ~new_U42 | ~new_P3_U3833;
  assign new_P3_U3349 = ~new_P3_U3681 | ~new_P3_U3679 | ~new_P3_U4559 | ~new_P3_U4558;
  assign new_P3_U3350 = ~new_U41 | ~new_P3_U3833;
  assign new_P3_U3351 = ~new_P3_U3685 | ~new_P3_U3683 | ~new_P3_U4577 | ~new_P3_U4576;
  assign new_P3_U3352 = ~new_P3_U3383 | ~new_P3_U3384;
  assign new_P3_U3353 = ~new_U40 | ~new_P3_U3833;
  assign new_P3_U3354 = ~new_P3_U3689 | ~new_P3_U3687 | ~new_P3_U4598 | ~new_P3_U4597 | ~new_P3_U4596;
  assign new_P3_U3355 = ~new_U38 | ~new_P3_U3833;
  assign new_P3_U3356 = ~new_U37 | ~new_P3_U3833;
  assign new_P3_U3357 = ~new_P3_U3015 | ~new_P3_U5456;
  assign new_P3_U3358 = ~new_P3_U3023 | ~new_P3_U4627;
  assign new_P3_U3359 = ~new_P3_U5447 | ~new_P3_U3385;
  assign new_P3_U3360 = ~new_P3_U3879 | ~new_P3_U5447;
  assign new_P3_U3361 = ~new_P3_U3055 | ~new_P3_U3911 | ~new_P3_U4595;
  assign new_P3_U3362 = ~new_P3_U3372 | ~new_P3_U3373 | ~new_P3_U3374;
  assign new_P3_U3363 = ~new_P3_U3694 | ~new_P3_U3910;
  assign new_P3_U3364 = ~new_P3_U3313 | ~new_P3_U3833;
  assign new_P3_U3365 = ~new_P3_U3877 | ~new_P3_U5423;
  assign new_P3_U3366 = ~new_P3_U3695 | ~new_P3_U3050;
  assign new_P3_U3367 = ~new_P3_U3882 | ~new_P3_U3385;
  assign new_P3_U3368 = ~new_P3_U3759 | ~new_P3_U3890;
  assign new_P3_U3369 = ~new_P3_U3876 | ~new_P3_U3378;
  assign new_P3_U3370 = ~new_P3_U3776 | ~new_P3_U4992 | ~new_P3_U4991;
  assign new_P3_U3371 = ~new_P3_U5417 | ~new_P3_U3917;
  assign new_P3_U3372 = ~new_P3_U5427 | ~new_P3_U5426;
  assign new_P3_U3373 = ~new_P3_U5430 | ~new_P3_U5429;
  assign new_P3_U3374 = ~new_P3_U5433 | ~new_P3_U5432;
  assign new_P3_U3375 = ~new_P3_U5439 | ~new_P3_U5438;
  assign n2784 = ~new_P3_U5442 | ~new_P3_U5441;
  assign n2789 = ~new_P3_U5444 | ~new_P3_U5443;
  assign new_P3_U3378 = ~new_P3_U5446 | ~new_P3_U5445;
  assign new_P3_U3379 = ~new_P3_U5449 | ~new_P3_U5448;
  assign new_P3_U3380 = ~new_P3_U5452 | ~new_P3_U5451;
  assign new_P3_U3381 = ~new_P3_U5458 | ~new_P3_U5457;
  assign new_P3_U3382 = ~new_P3_U5461 | ~new_P3_U5460;
  assign new_P3_U3383 = ~new_P3_U5464 | ~new_P3_U5463;
  assign new_P3_U3384 = ~new_P3_U5467 | ~new_P3_U5466;
  assign new_P3_U3385 = ~new_P3_U5455 | ~new_P3_U5454;
  assign new_P3_U3386 = ~new_P3_U5470 | ~new_P3_U5469;
  assign new_P3_U3387 = ~new_P3_U5472 | ~new_P3_U5471;
  assign new_P3_U3388 = ~new_P3_U5475 | ~new_P3_U5474;
  assign new_P3_U3389 = ~new_P3_U5478 | ~new_P3_U5477;
  assign n2944 = ~new_P3_U5484 | ~new_P3_U5483;
  assign new_P3_U3391 = ~new_P3_U5486 | ~new_P3_U5485;
  assign new_P3_U3392 = ~new_P3_U5488 | ~new_P3_U5487;
  assign n2949 = ~new_P3_U5491 | ~new_P3_U5490;
  assign new_P3_U3394 = ~new_P3_U5493 | ~new_P3_U5492;
  assign new_P3_U3395 = ~new_P3_U5495 | ~new_P3_U5494;
  assign n2954 = ~new_P3_U5498 | ~new_P3_U5497;
  assign new_P3_U3397 = ~new_P3_U5500 | ~new_P3_U5499;
  assign new_P3_U3398 = ~new_P3_U5502 | ~new_P3_U5501;
  assign n2959 = ~new_P3_U5505 | ~new_P3_U5504;
  assign new_P3_U3400 = ~new_P3_U5507 | ~new_P3_U5506;
  assign new_P3_U3401 = ~new_P3_U5509 | ~new_P3_U5508;
  assign n2964 = ~new_P3_U5512 | ~new_P3_U5511;
  assign new_P3_U3403 = ~new_P3_U5514 | ~new_P3_U5513;
  assign new_P3_U3404 = ~new_P3_U5516 | ~new_P3_U5515;
  assign n2969 = ~new_P3_U5519 | ~new_P3_U5518;
  assign new_P3_U3406 = ~new_P3_U5521 | ~new_P3_U5520;
  assign new_P3_U3407 = ~new_P3_U5523 | ~new_P3_U5522;
  assign n2974 = ~new_P3_U5526 | ~new_P3_U5525;
  assign new_P3_U3409 = ~new_P3_U5528 | ~new_P3_U5527;
  assign new_P3_U3410 = ~new_P3_U5530 | ~new_P3_U5529;
  assign n2979 = ~new_P3_U5533 | ~new_P3_U5532;
  assign new_P3_U3412 = ~new_P3_U5535 | ~new_P3_U5534;
  assign new_P3_U3413 = ~new_P3_U5537 | ~new_P3_U5536;
  assign n2984 = ~new_P3_U5540 | ~new_P3_U5539;
  assign new_P3_U3415 = ~new_P3_U5542 | ~new_P3_U5541;
  assign new_P3_U3416 = ~new_P3_U5544 | ~new_P3_U5543;
  assign n2989 = ~new_P3_U5547 | ~new_P3_U5546;
  assign new_P3_U3418 = ~new_P3_U5549 | ~new_P3_U5548;
  assign new_P3_U3419 = ~new_P3_U5551 | ~new_P3_U5550;
  assign n2994 = ~new_P3_U5554 | ~new_P3_U5553;
  assign new_P3_U3421 = ~new_P3_U5556 | ~new_P3_U5555;
  assign new_P3_U3422 = ~new_P3_U5558 | ~new_P3_U5557;
  assign n2999 = ~new_P3_U5561 | ~new_P3_U5560;
  assign new_P3_U3424 = ~new_P3_U5563 | ~new_P3_U5562;
  assign new_P3_U3425 = ~new_P3_U5565 | ~new_P3_U5564;
  assign n3004 = ~new_P3_U5568 | ~new_P3_U5567;
  assign new_P3_U3427 = ~new_P3_U5570 | ~new_P3_U5569;
  assign new_P3_U3428 = ~new_P3_U5572 | ~new_P3_U5571;
  assign n3009 = ~new_P3_U5575 | ~new_P3_U5574;
  assign new_P3_U3430 = ~new_P3_U5577 | ~new_P3_U5576;
  assign new_P3_U3431 = ~new_P3_U5579 | ~new_P3_U5578;
  assign n3014 = ~new_P3_U5582 | ~new_P3_U5581;
  assign new_P3_U3433 = ~new_P3_U5584 | ~new_P3_U5583;
  assign new_P3_U3434 = ~new_P3_U5586 | ~new_P3_U5585;
  assign n3019 = ~new_P3_U5589 | ~new_P3_U5588;
  assign new_P3_U3436 = ~new_P3_U5591 | ~new_P3_U5590;
  assign new_P3_U3437 = ~new_P3_U5593 | ~new_P3_U5592;
  assign n3024 = ~new_P3_U5596 | ~new_P3_U5595;
  assign new_P3_U3439 = ~new_P3_U5598 | ~new_P3_U5597;
  assign new_P3_U3440 = ~new_P3_U5600 | ~new_P3_U5599;
  assign n3029 = ~new_P3_U5603 | ~new_P3_U5602;
  assign new_P3_U3442 = ~new_P3_U5605 | ~new_P3_U5604;
  assign new_P3_U3443 = ~new_P3_U5607 | ~new_P3_U5606;
  assign n3034 = ~new_P3_U5610 | ~new_P3_U5609;
  assign new_P3_U3445 = ~new_P3_U5612 | ~new_P3_U5611;
  assign n3039 = ~new_P3_U5615 | ~new_P3_U5614;
  assign n3044 = ~new_P3_U5617 | ~new_P3_U5616;
  assign n3049 = ~new_P3_U5619 | ~new_P3_U5618;
  assign n3054 = ~new_P3_U5621 | ~new_P3_U5620;
  assign n3059 = ~new_P3_U5623 | ~new_P3_U5622;
  assign n3064 = ~new_P3_U5625 | ~new_P3_U5624;
  assign n3069 = ~new_P3_U5627 | ~new_P3_U5626;
  assign n3074 = ~new_P3_U5629 | ~new_P3_U5628;
  assign n3079 = ~new_P3_U5631 | ~new_P3_U5630;
  assign n3084 = ~new_P3_U5633 | ~new_P3_U5632;
  assign n3089 = ~new_P3_U5635 | ~new_P3_U5634;
  assign n3094 = ~new_P3_U5637 | ~new_P3_U5636;
  assign n3099 = ~new_P3_U5639 | ~new_P3_U5638;
  assign n3104 = ~new_P3_U5643 | ~new_P3_U5642;
  assign n3109 = ~new_P3_U5645 | ~new_P3_U5644;
  assign n3114 = ~new_P3_U5647 | ~new_P3_U5646;
  assign n3119 = ~new_P3_U5649 | ~new_P3_U5648;
  assign n3124 = ~new_P3_U5651 | ~new_P3_U5650;
  assign n3129 = ~new_P3_U5653 | ~new_P3_U5652;
  assign n3134 = ~new_P3_U5655 | ~new_P3_U5654;
  assign n3139 = ~new_P3_U5657 | ~new_P3_U5656;
  assign n3144 = ~new_P3_U5659 | ~new_P3_U5658;
  assign n3149 = ~new_P3_U5661 | ~new_P3_U5660;
  assign n3154 = ~new_P3_U5663 | ~new_P3_U5662;
  assign n3159 = ~new_P3_U5665 | ~new_P3_U5664;
  assign n3164 = ~new_P3_U5667 | ~new_P3_U5666;
  assign n3169 = ~new_P3_U5669 | ~new_P3_U5668;
  assign n3174 = ~new_P3_U5671 | ~new_P3_U5670;
  assign n3179 = ~new_P3_U5673 | ~new_P3_U5672;
  assign n3184 = ~new_P3_U5675 | ~new_P3_U5674;
  assign n3189 = ~new_P3_U5677 | ~new_P3_U5676;
  assign n3194 = ~new_P3_U5679 | ~new_P3_U5678;
  assign n3199 = ~new_P3_U5681 | ~new_P3_U5680;
  assign n3204 = ~new_P3_U5683 | ~new_P3_U5682;
  assign n3209 = ~new_P3_U5685 | ~new_P3_U5684;
  assign n3214 = ~new_P3_U5687 | ~new_P3_U5686;
  assign n3219 = ~new_P3_U5689 | ~new_P3_U5688;
  assign n3224 = ~new_P3_U5691 | ~new_P3_U5690;
  assign n3229 = ~new_P3_U5693 | ~new_P3_U5692;
  assign n3234 = ~new_P3_U5695 | ~new_P3_U5694;
  assign n3239 = ~new_P3_U5697 | ~new_P3_U5696;
  assign n3244 = ~new_P3_U5699 | ~new_P3_U5698;
  assign n3249 = ~new_P3_U5701 | ~new_P3_U5700;
  assign n3254 = ~new_P3_U5703 | ~new_P3_U5702;
  assign n3259 = ~new_P3_U5705 | ~new_P3_U5704;
  assign n3524 = ~new_P3_U5770 | ~new_P3_U5769;
  assign n3529 = ~new_P3_U5772 | ~new_P3_U5771;
  assign n3534 = ~new_P3_U5774 | ~new_P3_U5773;
  assign n3539 = ~new_P3_U5776 | ~new_P3_U5775;
  assign n3544 = ~new_P3_U5778 | ~new_P3_U5777;
  assign n3549 = ~new_P3_U5780 | ~new_P3_U5779;
  assign n3554 = ~new_P3_U5782 | ~new_P3_U5781;
  assign n3559 = ~new_P3_U5784 | ~new_P3_U5783;
  assign n3564 = ~new_P3_U5786 | ~new_P3_U5785;
  assign n3569 = ~new_P3_U5788 | ~new_P3_U5787;
  assign n3574 = ~new_P3_U5790 | ~new_P3_U5789;
  assign n3579 = ~new_P3_U5792 | ~new_P3_U5791;
  assign n3584 = ~new_P3_U5794 | ~new_P3_U5793;
  assign n3589 = ~new_P3_U5796 | ~new_P3_U5795;
  assign n3594 = ~new_P3_U5798 | ~new_P3_U5797;
  assign n3599 = ~new_P3_U5800 | ~new_P3_U5799;
  assign n3604 = ~new_P3_U5802 | ~new_P3_U5801;
  assign n3609 = ~new_P3_U5804 | ~new_P3_U5803;
  assign n3614 = ~new_P3_U5806 | ~new_P3_U5805;
  assign n3619 = ~new_P3_U5808 | ~new_P3_U5807;
  assign n3624 = ~new_P3_U5810 | ~new_P3_U5809;
  assign n3629 = ~new_P3_U5812 | ~new_P3_U5811;
  assign n3634 = ~new_P3_U5814 | ~new_P3_U5813;
  assign n3639 = ~new_P3_U5816 | ~new_P3_U5815;
  assign n3644 = ~new_P3_U5818 | ~new_P3_U5817;
  assign n3649 = ~new_P3_U5820 | ~new_P3_U5819;
  assign n3654 = ~new_P3_U5822 | ~new_P3_U5821;
  assign n3659 = ~new_P3_U5824 | ~new_P3_U5823;
  assign n3664 = ~new_P3_U5826 | ~new_P3_U5825;
  assign n3669 = ~new_P3_U5828 | ~new_P3_U5827;
  assign n3674 = ~new_P3_U5830 | ~new_P3_U5829;
  assign n3679 = ~new_P3_U5832 | ~new_P3_U5831;
  assign new_P3_U3523 = ~new_P3_U5946 | ~new_P3_U5945;
  assign new_P3_U3524 = ~new_P3_U5948 | ~new_P3_U5947;
  assign new_P3_U3525 = ~new_P3_U5950 | ~new_P3_U5949;
  assign new_P3_U3526 = ~new_P3_U5952 | ~new_P3_U5951;
  assign new_P3_U3527 = ~new_P3_U5954 | ~new_P3_U5953;
  assign new_P3_U3528 = ~new_P3_U5956 | ~new_P3_U5955;
  assign new_P3_U3529 = ~new_P3_U5958 | ~new_P3_U5957;
  assign new_P3_U3530 = ~new_P3_U5960 | ~new_P3_U5959;
  assign new_P3_U3531 = ~new_P3_U5962 | ~new_P3_U5961;
  assign new_P3_U3532 = ~new_P3_U5964 | ~new_P3_U5963;
  assign new_P3_U3533 = ~new_P3_U5966 | ~new_P3_U5965;
  assign new_P3_U3534 = ~new_P3_U5968 | ~new_P3_U5967;
  assign new_P3_U3535 = ~new_P3_U5970 | ~new_P3_U5969;
  assign new_P3_U3536 = ~new_P3_U5972 | ~new_P3_U5971;
  assign new_P3_U3537 = ~new_P3_U5974 | ~new_P3_U5973;
  assign new_P3_U3538 = ~new_P3_U5976 | ~new_P3_U5975;
  assign new_P3_U3539 = ~new_P3_U5978 | ~new_P3_U5977;
  assign new_P3_U3540 = ~new_P3_U5980 | ~new_P3_U5979;
  assign new_P3_U3541 = ~new_P3_U5982 | ~new_P3_U5981;
  assign new_P3_U3542 = ~new_P3_U5984 | ~new_P3_U5983;
  assign new_P3_U3543 = ~new_P3_U5986 | ~new_P3_U5985;
  assign new_P3_U3544 = ~new_P3_U5988 | ~new_P3_U5987;
  assign new_P3_U3545 = ~new_P3_U5990 | ~new_P3_U5989;
  assign new_P3_U3546 = ~new_P3_U5992 | ~new_P3_U5991;
  assign new_P3_U3547 = ~new_P3_U5994 | ~new_P3_U5993;
  assign new_P3_U3548 = ~new_P3_U5996 | ~new_P3_U5995;
  assign new_P3_U3549 = ~new_P3_U5998 | ~new_P3_U5997;
  assign new_P3_U3550 = ~new_P3_U6000 | ~new_P3_U5999;
  assign new_P3_U3551 = ~new_P3_U6002 | ~new_P3_U6001;
  assign new_P3_U3552 = ~new_P3_U6004 | ~new_P3_U6003;
  assign new_P3_U3553 = ~new_P3_U6006 | ~new_P3_U6005;
  assign new_P3_U3554 = ~new_P3_U6008 | ~new_P3_U6007;
  assign new_P3_U3555 = ~new_P3_U6010 | ~new_P3_U6009;
  assign new_P3_U3556 = ~new_P3_U6012 | ~new_P3_U6011;
  assign new_P3_U3557 = ~new_P3_U6014 | ~new_P3_U6013;
  assign new_P3_U3558 = ~new_P3_U6016 | ~new_P3_U6015;
  assign new_P3_U3559 = ~new_P3_U6018 | ~new_P3_U6017;
  assign new_P3_U3560 = ~new_P3_U6020 | ~new_P3_U6019;
  assign new_P3_U3561 = ~new_P3_U6022 | ~new_P3_U6021;
  assign new_P3_U3562 = ~new_P3_U6024 | ~new_P3_U6023;
  assign new_P3_U3563 = ~new_P3_U6026 | ~new_P3_U6025;
  assign new_P3_U3564 = ~new_P3_U6028 | ~new_P3_U6027;
  assign new_P3_U3565 = ~new_P3_U6030 | ~new_P3_U6029;
  assign new_P3_U3566 = ~new_P3_U6032 | ~new_P3_U6031;
  assign new_P3_U3567 = ~new_P3_U6034 | ~new_P3_U6033;
  assign new_P3_U3568 = ~new_P3_U6036 | ~new_P3_U6035;
  assign new_P3_U3569 = ~new_P3_U6038 | ~new_P3_U6037;
  assign new_P3_U3570 = ~new_P3_U6040 | ~new_P3_U6039;
  assign new_P3_U3571 = ~new_P3_U6042 | ~new_P3_U6041;
  assign new_P3_U3572 = ~new_P3_U6044 | ~new_P3_U6043;
  assign new_P3_U3573 = ~new_P3_U6046 | ~new_P3_U6045;
  assign new_P3_U3574 = ~new_P3_U6048 | ~new_P3_U6047;
  assign new_P3_U3575 = new_P3_U4066 & new_P3_U4065;
  assign new_P3_U3576 = new_P3_U4068 & new_P3_U4067;
  assign new_P3_U3577 = new_P3_U4075 & new_P3_U4076 & new_P3_U4074;
  assign new_P3_U3578 = new_P3_U4022 & new_P3_U4023 & new_P3_U4025 & new_P3_U4024;
  assign new_P3_U3579 = new_P3_U4026 & new_P3_U4027 & new_P3_U4029 & new_P3_U4028;
  assign new_P3_U3580 = new_P3_U4030 & new_P3_U4031 & new_P3_U4033 & new_P3_U4032;
  assign new_P3_U3581 = new_P3_U4036 & new_P3_U4035 & new_P3_U4034;
  assign new_P3_U3582 = new_P3_U3578 & new_P3_U3579 & new_P3_U3581 & new_P3_U3580;
  assign new_P3_U3583 = new_P3_U4037 & new_P3_U4038 & new_P3_U4040 & new_P3_U4039;
  assign new_P3_U3584 = new_P3_U4041 & new_P3_U4042 & new_P3_U4044 & new_P3_U4043;
  assign new_P3_U3585 = new_P3_U4045 & new_P3_U4046 & new_P3_U4048 & new_P3_U4047;
  assign new_P3_U3586 = new_P3_U4051 & new_P3_U4050 & new_P3_U4049;
  assign new_P3_U3587 = new_P3_U3583 & new_P3_U3584 & new_P3_U3586 & new_P3_U3585;
  assign new_P3_U3588 = new_P3_U3389 & new_P3_U3388;
  assign new_P3_U3589 = new_P3_U5479 & new_P3_U5476;
  assign new_P3_U3590 = new_P3_U4093 & new_P3_U4092;
  assign new_P3_U3591 = new_P3_U4095 & new_P3_U4094;
  assign new_P3_U3592 = new_P3_U3591 & new_P3_U4097 & new_P3_U4096;
  assign new_P3_U3593 = new_P3_U4099 & new_P3_U4100 & new_P3_U4101;
  assign new_P3_U3594 = new_P3_U4111 & new_P3_U4110;
  assign new_P3_U3595 = new_P3_U4113 & new_P3_U4112;
  assign new_P3_U3596 = new_P3_U3595 & new_P3_U4115 & new_P3_U4114;
  assign new_P3_U3597 = new_P3_U4117 & new_P3_U4118 & new_P3_U4119;
  assign new_P3_U3598 = new_P3_U4129 & new_P3_U4128;
  assign new_P3_U3599 = new_P3_U4131 & new_P3_U4130;
  assign new_P3_U3600 = new_P3_U3599 & new_P3_U4133 & new_P3_U4132;
  assign new_P3_U3601 = new_P3_U4135 & new_P3_U4136 & new_P3_U4137;
  assign new_P3_U3602 = new_P3_U4149 & new_P3_U4148;
  assign new_P3_U3603 = new_P3_U3602 & new_P3_U4151 & new_P3_U4150;
  assign new_P3_U3604 = new_P3_U4153 & new_P3_U4154 & new_P3_U4155;
  assign new_P3_U3605 = new_P3_U4167 & new_P3_U4166;
  assign new_P3_U3606 = new_P3_U3605 & new_P3_U4169 & new_P3_U4168;
  assign new_P3_U3607 = new_P3_U4171 & new_P3_U4172 & new_P3_U4173;
  assign new_P3_U3608 = new_P3_U4185 & new_P3_U4184;
  assign new_P3_U3609 = new_P3_U3608 & new_P3_U4187 & new_P3_U4186;
  assign new_P3_U3610 = new_P3_U4189 & new_P3_U4190 & new_P3_U4191;
  assign new_P3_U3611 = new_P3_U4203 & new_P3_U4202;
  assign new_P3_U3612 = new_P3_U3611 & new_P3_U4205 & new_P3_U4204;
  assign new_P3_U3613 = new_P3_U4207 & new_P3_U4208 & new_P3_U4209;
  assign new_P3_U3614 = new_P3_U4221 & new_P3_U4220;
  assign new_P3_U3615 = new_P3_U3614 & new_P3_U4223 & new_P3_U4222;
  assign new_P3_U3616 = new_P3_U4225 & new_P3_U4226 & new_P3_U4227;
  assign new_P3_U3617 = new_P3_U4237 & new_P3_U4236;
  assign new_P3_U3618 = new_P3_U4239 & new_P3_U4238;
  assign new_P3_U3619 = new_P3_U3618 & new_P3_U4241 & new_P3_U4240;
  assign new_P3_U3620 = new_P3_U4243 & new_P3_U4244 & new_P3_U4245;
  assign new_P3_U3621 = new_P3_U4255 & new_P3_U4254;
  assign new_P3_U3622 = new_P3_U4257 & new_P3_U4256;
  assign new_P3_U3623 = new_P3_U3622 & new_P3_U4259 & new_P3_U4258;
  assign new_P3_U3624 = new_P3_U4261 & new_P3_U4262 & new_P3_U4263;
  assign new_P3_U3625 = new_P3_U4275 & new_P3_U4274;
  assign new_P3_U3626 = new_P3_U3625 & new_P3_U4277 & new_P3_U4276;
  assign new_P3_U3627 = new_P3_U4279 & new_P3_U4280 & new_P3_U4281;
  assign new_P3_U3628 = new_P3_U4291 & new_P3_U4290;
  assign new_P3_U3629 = new_P3_U4293 & new_P3_U4292;
  assign new_P3_U3630 = new_P3_U3629 & new_P3_U4295 & new_P3_U4294;
  assign new_P3_U3631 = new_P3_U4297 & new_P3_U4298 & new_P3_U4299;
  assign new_P3_U3632 = new_P3_U4309 & new_P3_U4308;
  assign new_P3_U3633 = new_P3_U4311 & new_P3_U4310;
  assign new_P3_U3634 = new_P3_U3633 & new_P3_U4313 & new_P3_U4312;
  assign new_P3_U3635 = new_P3_U4315 & new_P3_U4316 & new_P3_U4317;
  assign new_P3_U3636 = new_P3_U4329 & new_P3_U4328;
  assign new_P3_U3637 = new_P3_U3636 & new_P3_U4331 & new_P3_U4330;
  assign new_P3_U3638 = new_P3_U4333 & new_P3_U4334 & new_P3_U4335;
  assign new_P3_U3639 = new_P3_U4347 & new_P3_U4346;
  assign new_P3_U3640 = new_P3_U3639 & new_P3_U4349 & new_P3_U4348;
  assign new_P3_U3641 = new_P3_U4351 & new_P3_U4352 & new_P3_U4353;
  assign new_P3_U3642 = new_P3_U4365 & new_P3_U4364;
  assign new_P3_U3643 = new_P3_U3642 & new_P3_U4367 & new_P3_U4366;
  assign new_P3_U3644 = new_P3_U4369 & new_P3_U4370 & new_P3_U4371;
  assign new_P3_U3645 = new_P3_U4381 & new_P3_U4380;
  assign new_P3_U3646 = new_P3_U4383 & new_P3_U4382;
  assign new_P3_U3647 = new_P3_U3646 & new_P3_U4385 & new_P3_U4384;
  assign new_P3_U3648 = new_P3_U4387 & new_P3_U4388 & new_P3_U4389;
  assign new_P3_U3649 = new_P3_U4401 & new_P3_U4400;
  assign new_P3_U3650 = new_P3_U3649 & new_P3_U4403 & new_P3_U4402;
  assign new_P3_U3651 = new_P3_U4405 & new_P3_U4406 & new_P3_U4407;
  assign new_P3_U3652 = new_P3_U4419 & new_P3_U4418;
  assign new_P3_U3653 = new_P3_U3652 & new_P3_U4421 & new_P3_U4420;
  assign new_P3_U3654 = new_P3_U4423 & new_P3_U4424 & new_P3_U4425;
  assign new_P3_U3655 = new_P3_U4437 & new_P3_U4436;
  assign new_P3_U3656 = new_P3_U3655 & new_P3_U4439 & new_P3_U4438;
  assign new_P3_U3657 = new_P3_U4441 & new_P3_U4442 & new_P3_U4443;
  assign new_P3_U3658 = new_P3_U4455 & new_P3_U4454;
  assign new_P3_U3659 = new_P3_U3658 & new_P3_U4457 & new_P3_U4456;
  assign new_P3_U3660 = new_P3_U4459 & new_P3_U4460 & new_P3_U4461;
  assign new_P3_U3661 = new_P3_U4473 & new_P3_U4472;
  assign new_P3_U3662 = new_P3_U3661 & new_P3_U4475 & new_P3_U4474;
  assign new_P3_U3663 = new_P3_U4477 & new_P3_U4478 & new_P3_U4479;
  assign new_P3_U3664 = new_P3_U4491 & new_P3_U4490;
  assign new_P3_U3665 = new_P3_U3664 & new_P3_U4493 & new_P3_U4492;
  assign new_P3_U3666 = new_P3_U4495 & new_P3_U4496 & new_P3_U4497;
  assign new_P3_U3667 = new_P3_U4507 & new_P3_U4506;
  assign new_P3_U3668 = new_P3_U4509 & new_P3_U4508;
  assign new_P3_U3669 = new_P3_U3668 & new_P3_U4511 & new_P3_U4510;
  assign new_P3_U3670 = new_P3_U4513 & new_P3_U4514 & new_P3_U4515;
  assign new_P3_U3671 = new_P3_U4525 & new_P3_U4524;
  assign new_P3_U3672 = new_P3_U4527 & new_P3_U4526;
  assign new_P3_U3673 = new_P3_U3672 & new_P3_U4529 & new_P3_U4528;
  assign new_P3_U3674 = new_P3_U4531 & new_P3_U4532 & new_P3_U4533;
  assign new_P3_U3675 = new_P3_U4543 & new_P3_U4542;
  assign new_P3_U3676 = new_P3_U4545 & new_P3_U4544;
  assign new_P3_U3677 = new_P3_U3676 & new_P3_U4547 & new_P3_U4546;
  assign new_P3_U3678 = new_P3_U4549 & new_P3_U4550 & new_P3_U4551;
  assign new_P3_U3679 = new_P3_U4561 & new_P3_U4560;
  assign new_P3_U3680 = new_P3_U4563 & new_P3_U4562;
  assign new_P3_U3681 = new_P3_U3680 & new_P3_U4565 & new_P3_U4564;
  assign new_P3_U3682 = new_P3_U4567 & new_P3_U4568 & new_P3_U4569;
  assign new_P3_U3683 = new_P3_U4579 & new_P3_U4578;
  assign new_P3_U3684 = new_P3_U4581 & new_P3_U4580;
  assign new_P3_U3685 = new_P3_U3684 & new_P3_U4583 & new_P3_U4582;
  assign new_P3_U3686 = new_P3_U4585 & new_P3_U4586 & new_P3_U4587;
  assign new_P3_U3687 = new_P3_U4600 & new_P3_U4599;
  assign new_P3_U3688 = new_P3_U4602 & new_P3_U4601;
  assign new_P3_U3689 = new_P3_U3688 & new_P3_U4604 & new_P3_U4603;
  assign new_P3_U3690 = new_P3_U4607 & new_P3_U4606;
  assign new_P3_U3691 = new_P3_U5476 & new_P3_U3389;
  assign new_P3_U3692 = new_P3_U5479 & new_P3_U3388;
  assign new_P3_U3693 = new_P3_U3920 & new_P3_U3379;
  assign new_P3_U3694 = new_P3_U5440 & P3_STATE_REG;
  assign new_P3_U3695 = new_P3_U5424 & new_P3_U3364;
  assign new_P3_U3696 = new_P3_U3375 & P3_STATE_REG;
  assign new_P3_U3697 = new_P3_U3307 & new_P3_U3306 & new_P3_U3305 & new_P3_U3301 & new_P3_U3308;
  assign new_P3_U3698 = new_P3_U3309 & new_P3_U3360;
  assign new_P3_U3699 = new_P3_U3701 & new_P3_U4765 & new_P3_U4763 & new_P3_U4762;
  assign new_P3_U3700 = new_P3_U4768 & new_P3_U4766;
  assign new_P3_U3701 = new_P3_U3700 & new_P3_U4767;
  assign new_P3_U3702 = new_P3_U3704 & new_P3_U4776 & new_P3_U4774 & new_P3_U4773;
  assign new_P3_U3703 = new_P3_U4779 & new_P3_U4777;
  assign new_P3_U3704 = new_P3_U3703 & new_P3_U4778;
  assign new_P3_U3705 = new_P3_U3707 & new_P3_U4787 & new_P3_U4785 & new_P3_U4784;
  assign new_P3_U3706 = new_P3_U4790 & new_P3_U4788;
  assign new_P3_U3707 = new_P3_U3706 & new_P3_U4789;
  assign new_P3_U3708 = new_P3_U3710 & new_P3_U4798 & new_P3_U4796 & new_P3_U4795;
  assign new_P3_U3709 = new_P3_U4801 & new_P3_U4799;
  assign new_P3_U3710 = new_P3_U3709 & new_P3_U4800;
  assign new_P3_U3711 = new_P3_U3713 & new_P3_U4809 & new_P3_U4807 & new_P3_U4806;
  assign new_P3_U3712 = new_P3_U4812 & new_P3_U4810;
  assign new_P3_U3713 = new_P3_U3712 & new_P3_U4811;
  assign new_P3_U3714 = new_P3_U3716 & new_P3_U4820 & new_P3_U4818 & new_P3_U4817;
  assign new_P3_U3715 = new_P3_U4823 & new_P3_U4821;
  assign new_P3_U3716 = new_P3_U3715 & new_P3_U4822;
  assign new_P3_U3717 = new_P3_U3719 & new_P3_U4831 & new_P3_U4829 & new_P3_U4828;
  assign new_P3_U3718 = new_P3_U4834 & new_P3_U4832;
  assign new_P3_U3719 = new_P3_U3718 & new_P3_U4833;
  assign new_P3_U3720 = new_P3_U3722 & new_P3_U4842 & new_P3_U4840 & new_P3_U4839;
  assign new_P3_U3721 = new_P3_U4845 & new_P3_U4843;
  assign new_P3_U3722 = new_P3_U3721 & new_P3_U4844;
  assign new_P3_U3723 = new_P3_U3725 & new_P3_U4853 & new_P3_U4851 & new_P3_U4850;
  assign new_P3_U3724 = new_P3_U4856 & new_P3_U4854;
  assign new_P3_U3725 = new_P3_U3724 & new_P3_U4855;
  assign new_P3_U3726 = new_P3_U3728 & new_P3_U4864 & new_P3_U4862 & new_P3_U4861;
  assign new_P3_U3727 = new_P3_U4867 & new_P3_U4865;
  assign new_P3_U3728 = new_P3_U3727 & new_P3_U4866;
  assign new_P3_U3729 = new_P3_U3731 & new_P3_U4875 & new_P3_U4873 & new_P3_U4872;
  assign new_P3_U3730 = new_P3_U4878 & new_P3_U4876;
  assign new_P3_U3731 = new_P3_U3730 & new_P3_U4877;
  assign new_P3_U3732 = new_P3_U3734 & new_P3_U4883 & new_P3_U4884 & new_P3_U4886;
  assign new_P3_U3733 = new_P3_U4889 & new_P3_U4887;
  assign new_P3_U3734 = new_P3_U3733 & new_P3_U4888;
  assign new_P3_U3735 = new_P3_U3737 & new_P3_U4894 & new_P3_U4895 & new_P3_U4897;
  assign new_P3_U3736 = new_P3_U4900 & new_P3_U4898;
  assign new_P3_U3737 = new_P3_U3736 & new_P3_U4899;
  assign new_P3_U3738 = new_P3_U3740 & new_P3_U4908 & new_P3_U4906;
  assign new_P3_U3739 = new_P3_U4911 & new_P3_U4909;
  assign new_P3_U3740 = new_P3_U3739 & new_P3_U4910;
  assign new_P3_U3741 = new_P3_U4919 & new_P3_U4917;
  assign new_P3_U3742 = new_P3_U4922 & new_P3_U4920;
  assign new_P3_U3743 = new_P3_U3742 & new_P3_U4921;
  assign new_P3_U3744 = new_P3_U4927 & new_P3_U4928 & new_P3_U3746;
  assign new_P3_U3745 = new_P3_U4933 & new_P3_U4931;
  assign new_P3_U3746 = new_P3_U3745 & new_P3_U4932;
  assign new_P3_U3747 = new_P3_U4938 & new_P3_U4939 & new_P3_U3749;
  assign new_P3_U3748 = new_P3_U4944 & new_P3_U4942;
  assign new_P3_U3749 = new_P3_U3748 & new_P3_U4943;
  assign new_P3_U3750 = new_P3_U3752 & new_P3_U4949 & new_P3_U4950 & new_P3_U4952;
  assign new_P3_U3751 = new_P3_U4955 & new_P3_U4953;
  assign new_P3_U3752 = new_P3_U3751 & new_P3_U4954;
  assign new_P3_U3753 = new_P3_U3755 & new_P3_U4963 & new_P3_U4961 & new_P3_U4960;
  assign new_P3_U3754 = new_P3_U4966 & new_P3_U4964;
  assign new_P3_U3755 = new_P3_U3754 & new_P3_U4965;
  assign new_P3_U3756 = new_P3_U3758 & new_P3_U4974 & new_P3_U4972 & new_P3_U4971;
  assign new_P3_U3757 = new_P3_U4977 & new_P3_U4975;
  assign new_P3_U3758 = new_P3_U3757 & new_P3_U4976;
  assign new_P3_U3759 = new_P3_U5468 & new_P3_U3383;
  assign new_P3_U3760 = ~new_P3_U5834 | ~new_P3_U5833;
  assign new_P3_U3761 = new_P3_U5915 & new_P3_U5912;
  assign new_P3_U3762 = new_P3_U5897 & new_P3_U3761 & new_P3_U3764 & new_P3_U3763;
  assign new_P3_U3763 = new_P3_U5903 & new_P3_U5900;
  assign new_P3_U3764 = new_P3_U5909 & new_P3_U5906;
  assign new_P3_U3765 = new_P3_U5879 & new_P3_U5885 & new_P3_U5882;
  assign new_P3_U3766 = new_P3_U5888 & new_P3_U5894 & new_P3_U5891;
  assign new_P3_U3767 = new_P3_U5873 & new_P3_U5876 & new_P3_U3766 & new_P3_U3765;
  assign new_P3_U3768 = new_P3_U5858 & new_P3_U5861 & new_P3_U5867 & new_P3_U5864;
  assign new_P3_U3769 = new_P3_U5855 & new_P3_U5852;
  assign new_P3_U3770 = new_P3_U5921 & new_P3_U5924 & new_P3_U5930 & new_P3_U5927;
  assign new_P3_U3771 = new_P3_U5846 & new_P3_U5843 & new_P3_U5840;
  assign new_P3_U3772 = new_P3_U3771 & new_P3_U5849 & new_P3_U5870 & new_P3_U3768 & new_P3_U3769;
  assign new_P3_U3773 = new_P3_U5933 & new_P3_U3770 & new_P3_U5918 & new_P3_U3762 & new_P3_U3767;
  assign new_P3_U3774 = new_P3_U4980 & new_P3_U4981 & new_P3_U3870;
  assign new_P3_U3775 = new_P3_U5416 & new_P3_U5415;
  assign new_P3_U3776 = new_P3_U3880 & new_P3_U4990 & new_P3_U5440 & new_P3_U3362;
  assign new_P3_U3777 = new_P3_U4998 & new_P3_U4997;
  assign new_P3_U3778 = new_P3_U5011 & new_P3_U5010;
  assign new_P3_U3779 = new_P3_U5020 & new_P3_U5019;
  assign new_P3_U3780 = new_P3_U5029 & new_P3_U5028;
  assign new_P3_U3781 = new_P3_U5036 & new_P3_U5034;
  assign new_P3_U3782 = new_P3_U5038 & new_P3_U5037;
  assign new_P3_U3783 = new_P3_U5047 & new_P3_U5046;
  assign new_P3_U3784 = new_P3_U5056 & new_P3_U5055;
  assign new_P3_U3785 = new_P3_U5065 & new_P3_U5064;
  assign new_P3_U3786 = new_P3_U5074 & new_P3_U5073;
  assign new_P3_U3787 = new_P3_U3031 & new_P3_U3077;
  assign new_P3_U3788 = new_P3_U5078 & new_P3_U5077;
  assign new_P3_U3789 = new_P3_U3788 & new_P3_U5081 & new_P3_U5080;
  assign new_P3_U3790 = new_P3_U5090 & new_P3_U5089;
  assign new_P3_U3791 = new_P3_U5097 & new_P3_U5095;
  assign new_P3_U3792 = new_P3_U5099 & new_P3_U5098;
  assign new_P3_U3793 = new_P3_U5108 & new_P3_U5107;
  assign new_P3_U3794 = new_P3_U5117 & new_P3_U5116;
  assign new_P3_U3795 = new_P3_U5126 & new_P3_U5125;
  assign new_P3_U3796 = new_P3_U5135 & new_P3_U5134;
  assign new_P3_U3797 = new_P3_U5144 & new_P3_U5143;
  assign new_P3_U3798 = new_P3_U5153 & new_P3_U5152;
  assign new_P3_U3799 = new_P3_U5162 & new_P3_U5161;
  assign new_P3_U3800 = new_P3_U5169 & new_P3_U5167;
  assign new_P3_U3801 = new_P3_U5171 & new_P3_U5170;
  assign new_P3_U3802 = new_P3_U5180 & new_P3_U5179;
  assign new_P3_U3803 = new_P3_U5189 & new_P3_U5188;
  assign new_P3_U3804 = new_P3_U5198 & new_P3_U5197;
  assign new_P3_U3805 = new_P3_U5205 & new_P3_U5203;
  assign new_P3_U3806 = new_P3_U5207 & new_P3_U5206;
  assign new_P3_U3807 = new_P3_U5216 & new_P3_U5215;
  assign new_P3_U3808 = new_P3_U5225 & new_P3_U5224;
  assign new_P3_U3809 = new_P3_U5234 & new_P3_U5233;
  assign new_P3_U3810 = new_P3_U5243 & new_P3_U5242;
  assign new_P3_U3811 = new_P3_U5252 & new_P3_U5251;
  assign new_P3_U3812 = new_P3_U5254 & P3_STATE_REG;
  assign new_P3_U3813 = new_P3_U5440 & new_P3_U3385;
  assign new_P3_U3814 = new_P3_U3385 & new_P3_U3375;
  assign new_P3_U3815 = new_P3_U3302 & new_P3_U3875 & new_P3_U3312;
  assign new_P3_U3816 = new_P3_U3310 & new_P3_U3357 & new_P3_U3877;
  assign new_P3_U3817 = new_P3_U3375 & new_P3_U5258;
  assign new_P3_U3818 = new_P3_U3375 & new_P3_U5260;
  assign new_P3_U3819 = new_P3_U3375 & new_P3_U5262;
  assign new_P3_U3820 = new_P3_U3375 & new_P3_U5264;
  assign new_P3_U3821 = new_P3_U3375 & new_P3_U5266;
  assign new_P3_U3822 = new_P3_U3375 & new_P3_U5268;
  assign new_P3_U3823 = new_P3_U3375 & new_P3_U5274;
  assign new_P3_U3824 = new_P3_U3375 & new_P3_U5296;
  assign new_P3_U3825 = new_P3_U3375 & new_P3_U5310;
  assign new_P3_U3826 = new_P3_U3375 & new_P3_U5312;
  assign new_P3_U3827 = new_P3_U3375 & new_P3_U5314;
  assign new_P3_U3828 = new_P3_U3375 & new_P3_U5316;
  assign new_P3_U3829 = new_P3_U3375 & new_P3_U5318;
  assign new_P3_U3830 = new_P3_U3375 & new_P3_U5320;
  assign new_P3_U3831 = ~P3_IR_REG_31_;
  assign new_P3_U3832 = ~new_P3_U3023 | ~new_P3_U3300;
  assign new_P3_U3833 = ~new_P3_U5468 | ~new_P3_U5465;
  assign new_P3_U3834 = ~new_P3_U5456 | ~new_P3_U5447;
  assign new_P3_U3835 = ~new_P3_U3023 | ~new_P3_U4058;
  assign new_P3_U3836 = ~new_P3_U3023 | ~new_P3_U4622;
  assign new_P3_U3837 = new_P3_U5707 & new_P3_U5706;
  assign new_P3_U3838 = new_P3_U5709 & new_P3_U5708;
  assign new_P3_U3839 = new_P3_U5711 & new_P3_U5710;
  assign new_P3_U3840 = new_P3_U5713 & new_P3_U5712;
  assign new_P3_U3841 = new_P3_U5715 & new_P3_U5714;
  assign new_P3_U3842 = new_P3_U5717 & new_P3_U5716;
  assign new_P3_U3843 = new_P3_U5719 & new_P3_U5718;
  assign new_P3_U3844 = new_P3_U5721 & new_P3_U5720;
  assign new_P3_U3845 = new_P3_U5723 & new_P3_U5722;
  assign new_P3_U3846 = new_P3_U5725 & new_P3_U5724;
  assign new_P3_U3847 = new_P3_U5727 & new_P3_U5726;
  assign new_P3_U3848 = new_P3_U5729 & new_P3_U5728;
  assign new_P3_U3849 = new_P3_U5731 & new_P3_U5730;
  assign new_P3_U3850 = new_P3_U5733 & new_P3_U5732;
  assign new_P3_U3851 = new_P3_U5735 & new_P3_U5734;
  assign new_P3_U3852 = new_P3_U5737 & new_P3_U5736;
  assign new_P3_U3853 = new_P3_U5739 & new_P3_U5738;
  assign new_P3_U3854 = new_P3_U5741 & new_P3_U5740;
  assign new_P3_U3855 = new_P3_U5743 & new_P3_U5742;
  assign new_P3_U3856 = new_P3_U5745 & new_P3_U5744;
  assign new_P3_U3857 = new_P3_U5747 & new_P3_U5746;
  assign new_P3_U3858 = new_P3_U5749 & new_P3_U5748;
  assign new_P3_U3859 = new_P3_U5751 & new_P3_U5750;
  assign new_P3_U3860 = new_P3_U5753 & new_P3_U5752;
  assign new_P3_U3861 = new_P3_U5755 & new_P3_U5754;
  assign new_P3_U3862 = new_P3_U5757 & new_P3_U5756;
  assign new_P3_U3863 = new_P3_U5759 & new_P3_U5758;
  assign new_P3_U3864 = new_P3_U5761 & new_P3_U5760;
  assign new_P3_U3865 = new_P3_U5763 & new_P3_U5762;
  assign new_P3_U3866 = new_P3_U5765 & new_P3_U5764;
  assign new_P3_U3867 = ~new_P3_R1269_U11;
  assign new_P3_U3868 = ~new_P3_U3773 | ~new_P3_U3772;
  assign new_P3_U3869 = ~new_P3_R693_U14;
  assign new_P3_U3870 = new_P3_U5940 & new_P3_U5939;
  assign new_P3_U3871 = ~new_P3_R1297_U6;
  assign new_P3_U3872 = ~new_P3_U3356;
  assign new_P3_U3873 = ~new_P3_U3355;
  assign new_P3_U3874 = ~new_P3_U3312;
  assign new_P3_U3875 = ~new_P3_U3015 | ~new_P3_U3385;
  assign new_P3_U3876 = ~new_P3_U3302;
  assign new_P3_U3877 = ~new_P3_U3016 | ~new_P3_U5456;
  assign new_P3_U3878 = ~new_P3_U3310;
  assign new_P3_U3879 = ~new_P3_U3357;
  assign new_P3_U3880 = ~new_P3_U3014 | ~new_P3_U3385;
  assign new_P3_U3881 = ~new_P3_U3308;
  assign new_P3_U3882 = ~new_P3_U3301;
  assign new_P3_U3883 = ~new_P3_U3305;
  assign new_P3_U3884 = ~new_P3_U3307;
  assign new_P3_U3885 = ~new_P3_U3306;
  assign new_P3_U3886 = ~new_P3_U3360;
  assign new_P3_U3887 = ~new_P3_U3311;
  assign new_P3_U3888 = ~new_P3_U3878 | ~new_P3_U3378;
  assign new_P3_U3889 = ~new_P3_U3369;
  assign new_P3_U3890 = ~new_P3_U3367;
  assign new_P3_U3891 = ~new_P3_U3309;
  assign new_P3_U3892 = ~new_P3_U3352;
  assign new_P3_U3893 = ~new_P3_U3833;
  assign new_P3_U3894 = ~new_P3_U3303;
  assign new_P3_U3895 = ~new_P3_U3304;
  assign new_P3_U3896 = ~new_P3_U5465 | ~new_P3_U3384;
  assign n3844 = ~new_P3_U3363;
  assign new_P3_U3898 = ~new_P3_U3364;
  assign new_P3_U3899 = ~new_P3_U3350;
  assign new_P3_U3900 = ~new_P3_U3348;
  assign new_P3_U3901 = ~new_P3_U3346;
  assign new_P3_U3902 = ~new_P3_U3344;
  assign new_P3_U3903 = ~new_P3_U3342;
  assign new_P3_U3904 = ~new_P3_U3340;
  assign new_P3_U3905 = ~new_P3_U3338;
  assign new_P3_U3906 = ~new_P3_U3336;
  assign new_P3_U3907 = ~new_P3_U3334;
  assign new_P3_U3908 = ~new_P3_U3353;
  assign new_P3_U3909 = ~new_P3_U3368;
  assign new_P3_U3910 = ~new_P3_U3362;
  assign new_P3_U3911 = ~new_P3_U3313;
  assign new_P3_U3912 = ~new_P3_U3358;
  assign new_P3_U3913 = ~new_P3_U3836;
  assign new_P3_U3914 = ~new_P3_U3835;
  assign new_P3_U3915 = ~new_P3_U3832;
  assign new_P3_U3916 = ~new_P3_U3361;
  assign new_P3_U3917 = ~new_P3_U3370 | ~P3_STATE_REG;
  assign new_P3_U3918 = ~new_P3_U3886 | ~new_P3_U3023;
  assign new_P3_U3919 = ~new_P3_U3299;
  assign new_P3_U3920 = ~new_P3_U3359;
  assign new_P3_U3921 = ~new_P3_U3297;
  assign new_P3_U3922 = ~new_U61 | ~n3834;
  assign new_P3_U3923 = ~P3_IR_REG_0_ | ~new_P3_U3027;
  assign new_P3_U3924 = ~P3_IR_REG_0_ | ~new_P3_U3921;
  assign new_P3_U3925 = ~new_U50 | ~n3834;
  assign new_P3_U3926 = ~new_P3_SUB_598_U51 | ~new_P3_U3027;
  assign new_P3_U3927 = ~P3_IR_REG_1_ | ~new_P3_U3921;
  assign new_P3_U3928 = ~new_U39 | ~n3834;
  assign new_P3_U3929 = ~new_P3_SUB_598_U22 | ~new_P3_U3027;
  assign new_P3_U3930 = ~P3_IR_REG_2_ | ~new_P3_U3921;
  assign new_P3_U3931 = ~new_U36 | ~n3834;
  assign new_P3_U3932 = ~new_P3_SUB_598_U23 | ~new_P3_U3027;
  assign new_P3_U3933 = ~P3_IR_REG_3_ | ~new_P3_U3921;
  assign new_P3_U3934 = ~new_U35 | ~n3834;
  assign new_P3_U3935 = ~new_P3_SUB_598_U24 | ~new_P3_U3027;
  assign new_P3_U3936 = ~P3_IR_REG_4_ | ~new_P3_U3921;
  assign new_P3_U3937 = ~new_U34 | ~n3834;
  assign new_P3_U3938 = ~new_P3_SUB_598_U74 | ~new_P3_U3027;
  assign new_P3_U3939 = ~P3_IR_REG_5_ | ~new_P3_U3921;
  assign new_P3_U3940 = ~new_U33 | ~n3834;
  assign new_P3_U3941 = ~new_P3_SUB_598_U25 | ~new_P3_U3027;
  assign new_P3_U3942 = ~P3_IR_REG_6_ | ~new_P3_U3921;
  assign new_P3_U3943 = ~new_U32 | ~n3834;
  assign new_P3_U3944 = ~new_P3_SUB_598_U26 | ~new_P3_U3027;
  assign new_P3_U3945 = ~P3_IR_REG_7_ | ~new_P3_U3921;
  assign new_P3_U3946 = ~new_U31 | ~n3834;
  assign new_P3_U3947 = ~new_P3_SUB_598_U27 | ~new_P3_U3027;
  assign new_P3_U3948 = ~P3_IR_REG_8_ | ~new_P3_U3921;
  assign new_P3_U3949 = ~new_U30 | ~n3834;
  assign new_P3_U3950 = ~new_P3_SUB_598_U72 | ~new_P3_U3027;
  assign new_P3_U3951 = ~P3_IR_REG_9_ | ~new_P3_U3921;
  assign new_P3_U3952 = ~new_U60 | ~n3834;
  assign new_P3_U3953 = ~new_P3_SUB_598_U7 | ~new_P3_U3027;
  assign new_P3_U3954 = ~P3_IR_REG_10_ | ~new_P3_U3921;
  assign new_P3_U3955 = ~new_U59 | ~n3834;
  assign new_P3_U3956 = ~new_P3_SUB_598_U8 | ~new_P3_U3027;
  assign new_P3_U3957 = ~P3_IR_REG_11_ | ~new_P3_U3921;
  assign new_P3_U3958 = ~new_U58 | ~n3834;
  assign new_P3_U3959 = ~new_P3_SUB_598_U9 | ~new_P3_U3027;
  assign new_P3_U3960 = ~P3_IR_REG_12_ | ~new_P3_U3921;
  assign new_P3_U3961 = ~new_U57 | ~n3834;
  assign new_P3_U3962 = ~new_P3_SUB_598_U89 | ~new_P3_U3027;
  assign new_P3_U3963 = ~P3_IR_REG_13_ | ~new_P3_U3921;
  assign new_P3_U3964 = ~new_U56 | ~n3834;
  assign new_P3_U3965 = ~new_P3_SUB_598_U10 | ~new_P3_U3027;
  assign new_P3_U3966 = ~P3_IR_REG_14_ | ~new_P3_U3921;
  assign new_P3_U3967 = ~new_U55 | ~n3834;
  assign new_P3_U3968 = ~new_P3_SUB_598_U11 | ~new_P3_U3027;
  assign new_P3_U3969 = ~P3_IR_REG_15_ | ~new_P3_U3921;
  assign new_P3_U3970 = ~new_U54 | ~n3834;
  assign new_P3_U3971 = ~new_P3_SUB_598_U12 | ~new_P3_U3027;
  assign new_P3_U3972 = ~P3_IR_REG_16_ | ~new_P3_U3921;
  assign new_P3_U3973 = ~new_U53 | ~n3834;
  assign new_P3_U3974 = ~new_P3_SUB_598_U87 | ~new_P3_U3027;
  assign new_P3_U3975 = ~P3_IR_REG_17_ | ~new_P3_U3921;
  assign new_P3_U3976 = ~new_U52 | ~n3834;
  assign new_P3_U3977 = ~new_P3_SUB_598_U13 | ~new_P3_U3027;
  assign new_P3_U3978 = ~P3_IR_REG_18_ | ~new_P3_U3921;
  assign new_P3_U3979 = ~new_U51 | ~n3834;
  assign new_P3_U3980 = ~new_P3_SUB_598_U14 | ~new_P3_U3027;
  assign new_P3_U3981 = ~P3_IR_REG_19_ | ~new_P3_U3921;
  assign new_P3_U3982 = ~new_U49 | ~n3834;
  assign new_P3_U3983 = ~new_P3_SUB_598_U15 | ~new_P3_U3027;
  assign new_P3_U3984 = ~P3_IR_REG_20_ | ~new_P3_U3921;
  assign new_P3_U3985 = ~new_U48 | ~n3834;
  assign new_P3_U3986 = ~new_P3_SUB_598_U83 | ~new_P3_U3027;
  assign new_P3_U3987 = ~P3_IR_REG_21_ | ~new_P3_U3921;
  assign new_P3_U3988 = ~new_U47 | ~n3834;
  assign new_P3_U3989 = ~new_P3_SUB_598_U16 | ~new_P3_U3027;
  assign new_P3_U3990 = ~P3_IR_REG_22_ | ~new_P3_U3921;
  assign new_P3_U3991 = ~new_U46 | ~n3834;
  assign new_P3_U3992 = ~new_P3_SUB_598_U17 | ~new_P3_U3027;
  assign new_P3_U3993 = ~P3_IR_REG_23_ | ~new_P3_U3921;
  assign new_P3_U3994 = ~new_U45 | ~n3834;
  assign new_P3_U3995 = ~new_P3_SUB_598_U18 | ~new_P3_U3027;
  assign new_P3_U3996 = ~P3_IR_REG_24_ | ~new_P3_U3921;
  assign new_P3_U3997 = ~new_U44 | ~n3834;
  assign new_P3_U3998 = ~new_P3_SUB_598_U81 | ~new_P3_U3027;
  assign new_P3_U3999 = ~P3_IR_REG_25_ | ~new_P3_U3921;
  assign new_P3_U4000 = ~new_U43 | ~n3834;
  assign new_P3_U4001 = ~new_P3_SUB_598_U19 | ~new_P3_U3027;
  assign new_P3_U4002 = ~P3_IR_REG_26_ | ~new_P3_U3921;
  assign new_P3_U4003 = ~new_U42 | ~n3834;
  assign new_P3_U4004 = ~new_P3_SUB_598_U79 | ~new_P3_U3027;
  assign new_P3_U4005 = ~P3_IR_REG_27_ | ~new_P3_U3921;
  assign new_P3_U4006 = ~new_U41 | ~n3834;
  assign new_P3_U4007 = ~new_P3_SUB_598_U20 | ~new_P3_U3027;
  assign new_P3_U4008 = ~P3_IR_REG_28_ | ~new_P3_U3921;
  assign new_P3_U4009 = ~new_U40 | ~n3834;
  assign new_P3_U4010 = ~new_P3_SUB_598_U21 | ~new_P3_U3027;
  assign new_P3_U4011 = ~P3_IR_REG_29_ | ~new_P3_U3921;
  assign new_P3_U4012 = ~new_U38 | ~n3834;
  assign new_P3_U4013 = ~new_P3_SUB_598_U77 | ~new_P3_U3027;
  assign new_P3_U4014 = ~P3_IR_REG_30_ | ~new_P3_U3921;
  assign new_P3_U4015 = ~new_U37 | ~n3834;
  assign new_P3_U4016 = ~new_P3_SUB_598_U52 | ~new_P3_U3027;
  assign new_P3_U4017 = ~P3_IR_REG_31_ | ~new_P3_U3921;
  assign new_P3_U4018 = ~new_P3_U3919 | ~new_P3_U5437;
  assign new_P3_U4019 = ~new_P3_U3300;
  assign new_P3_U4020 = ~new_P3_U3299 | ~new_P3_U5428;
  assign new_P3_U4021 = ~new_P3_U3299 | ~new_P3_U5431;
  assign new_P3_U4022 = ~new_P3_U4019 | ~P3_D_REG_10_;
  assign new_P3_U4023 = ~new_P3_U4019 | ~P3_D_REG_11_;
  assign new_P3_U4024 = ~new_P3_U4019 | ~P3_D_REG_12_;
  assign new_P3_U4025 = ~new_P3_U4019 | ~P3_D_REG_13_;
  assign new_P3_U4026 = ~new_P3_U4019 | ~P3_D_REG_14_;
  assign new_P3_U4027 = ~new_P3_U4019 | ~P3_D_REG_15_;
  assign new_P3_U4028 = ~new_P3_U4019 | ~P3_D_REG_16_;
  assign new_P3_U4029 = ~new_P3_U4019 | ~P3_D_REG_17_;
  assign new_P3_U4030 = ~new_P3_U4019 | ~P3_D_REG_18_;
  assign new_P3_U4031 = ~new_P3_U4019 | ~P3_D_REG_19_;
  assign new_P3_U4032 = ~new_P3_U4019 | ~P3_D_REG_20_;
  assign new_P3_U4033 = ~new_P3_U4019 | ~P3_D_REG_21_;
  assign new_P3_U4034 = ~new_P3_U4019 | ~P3_D_REG_22_;
  assign new_P3_U4035 = ~new_P3_U4019 | ~P3_D_REG_23_;
  assign new_P3_U4036 = ~new_P3_U4019 | ~P3_D_REG_24_;
  assign new_P3_U4037 = ~new_P3_U4019 | ~P3_D_REG_25_;
  assign new_P3_U4038 = ~new_P3_U4019 | ~P3_D_REG_26_;
  assign new_P3_U4039 = ~new_P3_U4019 | ~P3_D_REG_27_;
  assign new_P3_U4040 = ~new_P3_U4019 | ~P3_D_REG_28_;
  assign new_P3_U4041 = ~new_P3_U4019 | ~P3_D_REG_29_;
  assign new_P3_U4042 = ~new_P3_U4019 | ~P3_D_REG_2_;
  assign new_P3_U4043 = ~new_P3_U4019 | ~P3_D_REG_30_;
  assign new_P3_U4044 = ~new_P3_U4019 | ~P3_D_REG_31_;
  assign new_P3_U4045 = ~new_P3_U4019 | ~P3_D_REG_3_;
  assign new_P3_U4046 = ~new_P3_U4019 | ~P3_D_REG_4_;
  assign new_P3_U4047 = ~new_P3_U4019 | ~P3_D_REG_5_;
  assign new_P3_U4048 = ~new_P3_U4019 | ~P3_D_REG_6_;
  assign new_P3_U4049 = ~new_P3_U4019 | ~P3_D_REG_7_;
  assign new_P3_U4050 = ~new_P3_U4019 | ~P3_D_REG_8_;
  assign new_P3_U4051 = ~new_P3_U4019 | ~P3_D_REG_9_;
  assign new_P3_U4052 = ~new_P3_U3834;
  assign new_P3_U4053 = ~new_P3_U5456 | ~new_P3_U5450;
  assign new_P3_U4054 = ~new_P3_U5482 | ~new_P3_U4053;
  assign new_P3_U4055 = ~new_P3_U3369 | ~new_P3_U3367;
  assign new_P3_U4056 = ~new_P3_U3894 | ~new_P3_U4055;
  assign new_P3_U4057 = ~new_P3_U3895 | ~new_P3_U4054;
  assign new_P3_U4058 = ~new_P3_U4057 | ~new_P3_U4056;
  assign new_P3_U4059 = ~new_P3_U3022 | ~P3_REG0_REG_1_;
  assign new_P3_U4060 = ~P3_REG1_REG_1_ | ~new_P3_U3021;
  assign new_P3_U4061 = ~P3_REG2_REG_1_ | ~new_P3_U3020;
  assign new_P3_U4062 = ~P3_REG3_REG_1_ | ~new_P3_U3019;
  assign new_P3_U4063 = ~new_P3_U3077;
  assign new_P3_U4064 = ~new_P3_U3877 | ~new_P3_U3357;
  assign new_P3_U4065 = ~new_P3_U3883 | ~new_P3_R1110_U95;
  assign new_P3_U4066 = ~new_P3_U3885 | ~new_P3_R1077_U95;
  assign new_P3_U4067 = ~new_P3_U3884 | ~new_P3_R1095_U24;
  assign new_P3_U4068 = ~new_P3_U3881 | ~new_P3_R1143_U95;
  assign new_P3_U4069 = ~new_P3_U3891 | ~new_P3_R1161_U95;
  assign new_P3_U4070 = ~new_P3_U3887 | ~new_P3_R1131_U24;
  assign new_P3_U4071 = ~new_P3_U3017 | ~new_P3_R1200_U24;
  assign new_P3_U4072 = ~new_P3_U3314;
  assign new_P3_U4073 = ~new_P3_U3352 | ~new_P3_U3833;
  assign new_P3_U4074 = ~new_P3_R1179_U24 | ~new_P3_U3026;
  assign new_P3_U4075 = ~new_P3_U3025 | ~new_P3_U3077;
  assign new_P3_U4076 = ~new_P3_U3387 | ~new_P3_U4064;
  assign new_P3_U4077 = ~new_P3_U3577 | ~new_P3_U4072;
  assign new_P3_U4078 = ~P3_REG0_REG_2_ | ~new_P3_U3022;
  assign new_P3_U4079 = ~P3_REG1_REG_2_ | ~new_P3_U3021;
  assign new_P3_U4080 = ~P3_REG2_REG_2_ | ~new_P3_U3020;
  assign new_P3_U4081 = ~P3_REG3_REG_2_ | ~new_P3_U3019;
  assign new_P3_U4082 = ~new_P3_U3067;
  assign new_P3_U4083 = ~P3_REG0_REG_0_ | ~new_P3_U3022;
  assign new_P3_U4084 = ~P3_REG1_REG_0_ | ~new_P3_U3021;
  assign new_P3_U4085 = ~P3_REG2_REG_0_ | ~new_P3_U3020;
  assign new_P3_U4086 = ~P3_REG3_REG_0_ | ~new_P3_U3019;
  assign new_P3_U4087 = ~new_P3_U3076;
  assign new_P3_U4088 = ~new_P3_U5468 | ~new_P3_U3383;
  assign new_P3_U4089 = ~new_P3_U3896 | ~new_P3_U4088;
  assign new_P3_U4090 = ~new_P3_U3033 | ~new_P3_U3076;
  assign new_P3_U4091 = ~new_P3_R1110_U94 | ~new_P3_U3883;
  assign new_P3_U4092 = ~new_P3_R1077_U94 | ~new_P3_U3885;
  assign new_P3_U4093 = ~new_P3_R1095_U100 | ~new_P3_U3884;
  assign new_P3_U4094 = ~new_P3_R1143_U94 | ~new_P3_U3881;
  assign new_P3_U4095 = ~new_P3_R1161_U94 | ~new_P3_U3891;
  assign new_P3_U4096 = ~new_P3_R1131_U100 | ~new_P3_U3887;
  assign new_P3_U4097 = ~new_P3_R1200_U100 | ~new_P3_U3017;
  assign new_P3_U4098 = ~new_P3_U3315;
  assign new_P3_U4099 = ~new_P3_R1179_U100 | ~new_P3_U3026;
  assign new_P3_U4100 = ~new_P3_U3025 | ~new_P3_U3067;
  assign new_P3_U4101 = ~new_P3_U3392 | ~new_P3_U4064;
  assign new_P3_U4102 = ~new_P3_U3593 | ~new_P3_U4098;
  assign new_P3_U4103 = ~P3_REG0_REG_3_ | ~new_P3_U3022;
  assign new_P3_U4104 = ~P3_REG1_REG_3_ | ~new_P3_U3021;
  assign new_P3_U4105 = ~P3_REG2_REG_3_ | ~new_P3_U3020;
  assign new_P3_U4106 = ~new_P3_SUB_609_U25 | ~new_P3_U3019;
  assign new_P3_U4107 = ~new_P3_U3063;
  assign new_P3_U4108 = ~new_P3_U3033 | ~new_P3_U3077;
  assign new_P3_U4109 = ~new_P3_R1110_U16 | ~new_P3_U3883;
  assign new_P3_U4110 = ~new_P3_R1077_U16 | ~new_P3_U3885;
  assign new_P3_U4111 = ~new_P3_R1095_U110 | ~new_P3_U3884;
  assign new_P3_U4112 = ~new_P3_R1143_U16 | ~new_P3_U3881;
  assign new_P3_U4113 = ~new_P3_R1161_U16 | ~new_P3_U3891;
  assign new_P3_U4114 = ~new_P3_R1131_U110 | ~new_P3_U3887;
  assign new_P3_U4115 = ~new_P3_R1200_U110 | ~new_P3_U3017;
  assign new_P3_U4116 = ~new_P3_U3316;
  assign new_P3_U4117 = ~new_P3_R1179_U110 | ~new_P3_U3026;
  assign new_P3_U4118 = ~new_P3_U3025 | ~new_P3_U3063;
  assign new_P3_U4119 = ~new_P3_U3395 | ~new_P3_U4064;
  assign new_P3_U4120 = ~new_P3_U3597 | ~new_P3_U4116;
  assign new_P3_U4121 = ~P3_REG0_REG_4_ | ~new_P3_U3022;
  assign new_P3_U4122 = ~P3_REG1_REG_4_ | ~new_P3_U3021;
  assign new_P3_U4123 = ~P3_REG2_REG_4_ | ~new_P3_U3020;
  assign new_P3_U4124 = ~new_P3_SUB_609_U29 | ~new_P3_U3019;
  assign new_P3_U4125 = ~new_P3_U3059;
  assign new_P3_U4126 = ~new_P3_U3033 | ~new_P3_U3067;
  assign new_P3_U4127 = ~new_P3_R1110_U100 | ~new_P3_U3883;
  assign new_P3_U4128 = ~new_P3_R1077_U100 | ~new_P3_U3885;
  assign new_P3_U4129 = ~new_P3_R1095_U21 | ~new_P3_U3884;
  assign new_P3_U4130 = ~new_P3_R1143_U100 | ~new_P3_U3881;
  assign new_P3_U4131 = ~new_P3_R1161_U100 | ~new_P3_U3891;
  assign new_P3_U4132 = ~new_P3_R1131_U21 | ~new_P3_U3887;
  assign new_P3_U4133 = ~new_P3_R1200_U21 | ~new_P3_U3017;
  assign new_P3_U4134 = ~new_P3_U3317;
  assign new_P3_U4135 = ~new_P3_R1179_U21 | ~new_P3_U3026;
  assign new_P3_U4136 = ~new_P3_U3025 | ~new_P3_U3059;
  assign new_P3_U4137 = ~new_P3_U3398 | ~new_P3_U4064;
  assign new_P3_U4138 = ~new_P3_U3601 | ~new_P3_U4134;
  assign new_P3_U4139 = ~P3_REG0_REG_5_ | ~new_P3_U3022;
  assign new_P3_U4140 = ~P3_REG1_REG_5_ | ~new_P3_U3021;
  assign new_P3_U4141 = ~P3_REG2_REG_5_ | ~new_P3_U3020;
  assign new_P3_U4142 = ~new_P3_SUB_609_U53 | ~new_P3_U3019;
  assign new_P3_U4143 = ~new_P3_U3066;
  assign new_P3_U4144 = ~new_P3_U3033 | ~new_P3_U3063;
  assign new_P3_U4145 = ~new_P3_R1110_U99 | ~new_P3_U3883;
  assign new_P3_U4146 = ~new_P3_R1077_U99 | ~new_P3_U3885;
  assign new_P3_U4147 = ~new_P3_R1095_U109 | ~new_P3_U3884;
  assign new_P3_U4148 = ~new_P3_R1143_U99 | ~new_P3_U3881;
  assign new_P3_U4149 = ~new_P3_R1161_U99 | ~new_P3_U3891;
  assign new_P3_U4150 = ~new_P3_R1131_U109 | ~new_P3_U3887;
  assign new_P3_U4151 = ~new_P3_R1200_U109 | ~new_P3_U3017;
  assign new_P3_U4152 = ~new_P3_U3318;
  assign new_P3_U4153 = ~new_P3_R1179_U109 | ~new_P3_U3026;
  assign new_P3_U4154 = ~new_P3_U3025 | ~new_P3_U3066;
  assign new_P3_U4155 = ~new_P3_U3401 | ~new_P3_U4064;
  assign new_P3_U4156 = ~new_P3_U3604 | ~new_P3_U4152;
  assign new_P3_U4157 = ~P3_REG0_REG_6_ | ~new_P3_U3022;
  assign new_P3_U4158 = ~P3_REG1_REG_6_ | ~new_P3_U3021;
  assign new_P3_U4159 = ~P3_REG2_REG_6_ | ~new_P3_U3020;
  assign new_P3_U4160 = ~new_P3_SUB_609_U8 | ~new_P3_U3019;
  assign new_P3_U4161 = ~new_P3_U3070;
  assign new_P3_U4162 = ~new_P3_U3033 | ~new_P3_U3059;
  assign new_P3_U4163 = ~new_P3_R1110_U17 | ~new_P3_U3883;
  assign new_P3_U4164 = ~new_P3_R1077_U17 | ~new_P3_U3885;
  assign new_P3_U4165 = ~new_P3_R1095_U108 | ~new_P3_U3884;
  assign new_P3_U4166 = ~new_P3_R1143_U17 | ~new_P3_U3881;
  assign new_P3_U4167 = ~new_P3_R1161_U17 | ~new_P3_U3891;
  assign new_P3_U4168 = ~new_P3_R1131_U108 | ~new_P3_U3887;
  assign new_P3_U4169 = ~new_P3_R1200_U108 | ~new_P3_U3017;
  assign new_P3_U4170 = ~new_P3_U3319;
  assign new_P3_U4171 = ~new_P3_R1179_U108 | ~new_P3_U3026;
  assign new_P3_U4172 = ~new_P3_U3025 | ~new_P3_U3070;
  assign new_P3_U4173 = ~new_P3_U3404 | ~new_P3_U4064;
  assign new_P3_U4174 = ~new_P3_U3607 | ~new_P3_U4170;
  assign new_P3_U4175 = ~P3_REG0_REG_7_ | ~new_P3_U3022;
  assign new_P3_U4176 = ~P3_REG1_REG_7_ | ~new_P3_U3021;
  assign new_P3_U4177 = ~P3_REG2_REG_7_ | ~new_P3_U3020;
  assign new_P3_U4178 = ~new_P3_SUB_609_U18 | ~new_P3_U3019;
  assign new_P3_U4179 = ~new_P3_U3069;
  assign new_P3_U4180 = ~new_P3_U3033 | ~new_P3_U3066;
  assign new_P3_U4181 = ~new_P3_R1110_U98 | ~new_P3_U3883;
  assign new_P3_U4182 = ~new_P3_R1077_U98 | ~new_P3_U3885;
  assign new_P3_U4183 = ~new_P3_R1095_U22 | ~new_P3_U3884;
  assign new_P3_U4184 = ~new_P3_R1143_U98 | ~new_P3_U3881;
  assign new_P3_U4185 = ~new_P3_R1161_U98 | ~new_P3_U3891;
  assign new_P3_U4186 = ~new_P3_R1131_U22 | ~new_P3_U3887;
  assign new_P3_U4187 = ~new_P3_R1200_U22 | ~new_P3_U3017;
  assign new_P3_U4188 = ~new_P3_U3320;
  assign new_P3_U4189 = ~new_P3_R1179_U22 | ~new_P3_U3026;
  assign new_P3_U4190 = ~new_P3_U3025 | ~new_P3_U3069;
  assign new_P3_U4191 = ~new_P3_U3407 | ~new_P3_U4064;
  assign new_P3_U4192 = ~new_P3_U3610 | ~new_P3_U4188;
  assign new_P3_U4193 = ~P3_REG0_REG_8_ | ~new_P3_U3022;
  assign new_P3_U4194 = ~P3_REG1_REG_8_ | ~new_P3_U3021;
  assign new_P3_U4195 = ~P3_REG2_REG_8_ | ~new_P3_U3020;
  assign new_P3_U4196 = ~new_P3_SUB_609_U12 | ~new_P3_U3019;
  assign new_P3_U4197 = ~new_P3_U3083;
  assign new_P3_U4198 = ~new_P3_U3033 | ~new_P3_U3070;
  assign new_P3_U4199 = ~new_P3_R1110_U18 | ~new_P3_U3883;
  assign new_P3_U4200 = ~new_P3_R1077_U18 | ~new_P3_U3885;
  assign new_P3_U4201 = ~new_P3_R1095_U107 | ~new_P3_U3884;
  assign new_P3_U4202 = ~new_P3_R1143_U18 | ~new_P3_U3881;
  assign new_P3_U4203 = ~new_P3_R1161_U18 | ~new_P3_U3891;
  assign new_P3_U4204 = ~new_P3_R1131_U107 | ~new_P3_U3887;
  assign new_P3_U4205 = ~new_P3_R1200_U107 | ~new_P3_U3017;
  assign new_P3_U4206 = ~new_P3_U3321;
  assign new_P3_U4207 = ~new_P3_R1179_U107 | ~new_P3_U3026;
  assign new_P3_U4208 = ~new_P3_U3025 | ~new_P3_U3083;
  assign new_P3_U4209 = ~new_P3_U3410 | ~new_P3_U4064;
  assign new_P3_U4210 = ~new_P3_U3613 | ~new_P3_U4206;
  assign new_P3_U4211 = ~P3_REG0_REG_9_ | ~new_P3_U3022;
  assign new_P3_U4212 = ~P3_REG1_REG_9_ | ~new_P3_U3021;
  assign new_P3_U4213 = ~P3_REG2_REG_9_ | ~new_P3_U3020;
  assign new_P3_U4214 = ~new_P3_SUB_609_U14 | ~new_P3_U3019;
  assign new_P3_U4215 = ~new_P3_U3082;
  assign new_P3_U4216 = ~new_P3_U3033 | ~new_P3_U3069;
  assign new_P3_U4217 = ~new_P3_R1110_U97 | ~new_P3_U3883;
  assign new_P3_U4218 = ~new_P3_R1077_U97 | ~new_P3_U3885;
  assign new_P3_U4219 = ~new_P3_R1095_U23 | ~new_P3_U3884;
  assign new_P3_U4220 = ~new_P3_R1143_U97 | ~new_P3_U3881;
  assign new_P3_U4221 = ~new_P3_R1161_U97 | ~new_P3_U3891;
  assign new_P3_U4222 = ~new_P3_R1131_U23 | ~new_P3_U3887;
  assign new_P3_U4223 = ~new_P3_R1200_U23 | ~new_P3_U3017;
  assign new_P3_U4224 = ~new_P3_U3322;
  assign new_P3_U4225 = ~new_P3_R1179_U23 | ~new_P3_U3026;
  assign new_P3_U4226 = ~new_P3_U3025 | ~new_P3_U3082;
  assign new_P3_U4227 = ~new_P3_U3413 | ~new_P3_U4064;
  assign new_P3_U4228 = ~new_P3_U3616 | ~new_P3_U4224;
  assign new_P3_U4229 = ~P3_REG0_REG_10_ | ~new_P3_U3022;
  assign new_P3_U4230 = ~P3_REG1_REG_10_ | ~new_P3_U3021;
  assign new_P3_U4231 = ~P3_REG2_REG_10_ | ~new_P3_U3020;
  assign new_P3_U4232 = ~new_P3_SUB_609_U13 | ~new_P3_U3019;
  assign new_P3_U4233 = ~new_P3_U3061;
  assign new_P3_U4234 = ~new_P3_U3033 | ~new_P3_U3083;
  assign new_P3_U4235 = ~new_P3_R1110_U96 | ~new_P3_U3883;
  assign new_P3_U4236 = ~new_P3_R1077_U96 | ~new_P3_U3885;
  assign new_P3_U4237 = ~new_P3_R1095_U106 | ~new_P3_U3884;
  assign new_P3_U4238 = ~new_P3_R1143_U96 | ~new_P3_U3881;
  assign new_P3_U4239 = ~new_P3_R1161_U96 | ~new_P3_U3891;
  assign new_P3_U4240 = ~new_P3_R1131_U106 | ~new_P3_U3887;
  assign new_P3_U4241 = ~new_P3_R1200_U106 | ~new_P3_U3017;
  assign new_P3_U4242 = ~new_P3_U3323;
  assign new_P3_U4243 = ~new_P3_R1179_U106 | ~new_P3_U3026;
  assign new_P3_U4244 = ~new_P3_U3025 | ~new_P3_U3061;
  assign new_P3_U4245 = ~new_P3_U3416 | ~new_P3_U4064;
  assign new_P3_U4246 = ~new_P3_U3620 | ~new_P3_U4242;
  assign new_P3_U4247 = ~P3_REG0_REG_11_ | ~new_P3_U3022;
  assign new_P3_U4248 = ~P3_REG1_REG_11_ | ~new_P3_U3021;
  assign new_P3_U4249 = ~P3_REG2_REG_11_ | ~new_P3_U3020;
  assign new_P3_U4250 = ~new_P3_SUB_609_U9 | ~new_P3_U3019;
  assign new_P3_U4251 = ~new_P3_U3062;
  assign new_P3_U4252 = ~new_P3_U3033 | ~new_P3_U3082;
  assign new_P3_U4253 = ~new_P3_R1110_U10 | ~new_P3_U3883;
  assign new_P3_U4254 = ~new_P3_R1077_U10 | ~new_P3_U3885;
  assign new_P3_U4255 = ~new_P3_R1095_U116 | ~new_P3_U3884;
  assign new_P3_U4256 = ~new_P3_R1143_U10 | ~new_P3_U3881;
  assign new_P3_U4257 = ~new_P3_R1161_U10 | ~new_P3_U3891;
  assign new_P3_U4258 = ~new_P3_R1131_U116 | ~new_P3_U3887;
  assign new_P3_U4259 = ~new_P3_R1200_U116 | ~new_P3_U3017;
  assign new_P3_U4260 = ~new_P3_U3324;
  assign new_P3_U4261 = ~new_P3_R1179_U116 | ~new_P3_U3026;
  assign new_P3_U4262 = ~new_P3_U3025 | ~new_P3_U3062;
  assign new_P3_U4263 = ~new_P3_U3419 | ~new_P3_U4064;
  assign new_P3_U4264 = ~new_P3_U3624 | ~new_P3_U4260;
  assign new_P3_U4265 = ~P3_REG0_REG_12_ | ~new_P3_U3022;
  assign new_P3_U4266 = ~P3_REG1_REG_12_ | ~new_P3_U3021;
  assign new_P3_U4267 = ~P3_REG2_REG_12_ | ~new_P3_U3020;
  assign new_P3_U4268 = ~new_P3_SUB_609_U23 | ~new_P3_U3019;
  assign new_P3_U4269 = ~new_P3_U3071;
  assign new_P3_U4270 = ~new_P3_U3033 | ~new_P3_U3061;
  assign new_P3_U4271 = ~new_P3_R1110_U114 | ~new_P3_U3883;
  assign new_P3_U4272 = ~new_P3_R1077_U114 | ~new_P3_U3885;
  assign new_P3_U4273 = ~new_P3_R1095_U16 | ~new_P3_U3884;
  assign new_P3_U4274 = ~new_P3_R1143_U114 | ~new_P3_U3881;
  assign new_P3_U4275 = ~new_P3_R1161_U114 | ~new_P3_U3891;
  assign new_P3_U4276 = ~new_P3_R1131_U16 | ~new_P3_U3887;
  assign new_P3_U4277 = ~new_P3_R1200_U16 | ~new_P3_U3017;
  assign new_P3_U4278 = ~new_P3_U3325;
  assign new_P3_U4279 = ~new_P3_R1179_U16 | ~new_P3_U3026;
  assign new_P3_U4280 = ~new_P3_U3025 | ~new_P3_U3071;
  assign new_P3_U4281 = ~new_P3_U3422 | ~new_P3_U4064;
  assign new_P3_U4282 = ~new_P3_U3627 | ~new_P3_U4278;
  assign new_P3_U4283 = ~P3_REG0_REG_13_ | ~new_P3_U3022;
  assign new_P3_U4284 = ~P3_REG1_REG_13_ | ~new_P3_U3021;
  assign new_P3_U4285 = ~P3_REG2_REG_13_ | ~new_P3_U3020;
  assign new_P3_U4286 = ~new_P3_SUB_609_U24 | ~new_P3_U3019;
  assign new_P3_U4287 = ~new_P3_U3079;
  assign new_P3_U4288 = ~new_P3_U3033 | ~new_P3_U3062;
  assign new_P3_U4289 = ~new_P3_R1110_U113 | ~new_P3_U3883;
  assign new_P3_U4290 = ~new_P3_R1077_U113 | ~new_P3_U3885;
  assign new_P3_U4291 = ~new_P3_R1095_U105 | ~new_P3_U3884;
  assign new_P3_U4292 = ~new_P3_R1143_U113 | ~new_P3_U3881;
  assign new_P3_U4293 = ~new_P3_R1161_U113 | ~new_P3_U3891;
  assign new_P3_U4294 = ~new_P3_R1131_U105 | ~new_P3_U3887;
  assign new_P3_U4295 = ~new_P3_R1200_U105 | ~new_P3_U3017;
  assign new_P3_U4296 = ~new_P3_U3326;
  assign new_P3_U4297 = ~new_P3_R1179_U105 | ~new_P3_U3026;
  assign new_P3_U4298 = ~new_P3_U3025 | ~new_P3_U3079;
  assign new_P3_U4299 = ~new_P3_U3425 | ~new_P3_U4064;
  assign new_P3_U4300 = ~new_P3_U3631 | ~new_P3_U4296;
  assign new_P3_U4301 = ~P3_REG0_REG_14_ | ~new_P3_U3022;
  assign new_P3_U4302 = ~P3_REG1_REG_14_ | ~new_P3_U3021;
  assign new_P3_U4303 = ~P3_REG2_REG_14_ | ~new_P3_U3020;
  assign new_P3_U4304 = ~new_P3_SUB_609_U30 | ~new_P3_U3019;
  assign new_P3_U4305 = ~new_P3_U3078;
  assign new_P3_U4306 = ~new_P3_U3033 | ~new_P3_U3071;
  assign new_P3_U4307 = ~new_P3_R1110_U11 | ~new_P3_U3883;
  assign new_P3_U4308 = ~new_P3_R1077_U11 | ~new_P3_U3885;
  assign new_P3_U4309 = ~new_P3_R1095_U104 | ~new_P3_U3884;
  assign new_P3_U4310 = ~new_P3_R1143_U11 | ~new_P3_U3881;
  assign new_P3_U4311 = ~new_P3_R1161_U11 | ~new_P3_U3891;
  assign new_P3_U4312 = ~new_P3_R1131_U104 | ~new_P3_U3887;
  assign new_P3_U4313 = ~new_P3_R1200_U104 | ~new_P3_U3017;
  assign new_P3_U4314 = ~new_P3_U3327;
  assign new_P3_U4315 = ~new_P3_R1179_U104 | ~new_P3_U3026;
  assign new_P3_U4316 = ~new_P3_U3025 | ~new_P3_U3078;
  assign new_P3_U4317 = ~new_P3_U3428 | ~new_P3_U4064;
  assign new_P3_U4318 = ~new_P3_U3635 | ~new_P3_U4314;
  assign new_P3_U4319 = ~P3_REG0_REG_15_ | ~new_P3_U3022;
  assign new_P3_U4320 = ~P3_REG1_REG_15_ | ~new_P3_U3021;
  assign new_P3_U4321 = ~P3_REG2_REG_15_ | ~new_P3_U3020;
  assign new_P3_U4322 = ~new_P3_SUB_609_U21 | ~new_P3_U3019;
  assign new_P3_U4323 = ~new_P3_U3073;
  assign new_P3_U4324 = ~new_P3_U3033 | ~new_P3_U3079;
  assign new_P3_U4325 = ~new_P3_R1110_U112 | ~new_P3_U3883;
  assign new_P3_U4326 = ~new_P3_R1077_U112 | ~new_P3_U3885;
  assign new_P3_U4327 = ~new_P3_R1095_U115 | ~new_P3_U3884;
  assign new_P3_U4328 = ~new_P3_R1143_U112 | ~new_P3_U3881;
  assign new_P3_U4329 = ~new_P3_R1161_U112 | ~new_P3_U3891;
  assign new_P3_U4330 = ~new_P3_R1131_U115 | ~new_P3_U3887;
  assign new_P3_U4331 = ~new_P3_R1200_U115 | ~new_P3_U3017;
  assign new_P3_U4332 = ~new_P3_U3328;
  assign new_P3_U4333 = ~new_P3_R1179_U115 | ~new_P3_U3026;
  assign new_P3_U4334 = ~new_P3_U3025 | ~new_P3_U3073;
  assign new_P3_U4335 = ~new_P3_U3431 | ~new_P3_U4064;
  assign new_P3_U4336 = ~new_P3_U3638 | ~new_P3_U4332;
  assign new_P3_U4337 = ~P3_REG0_REG_16_ | ~new_P3_U3022;
  assign new_P3_U4338 = ~P3_REG1_REG_16_ | ~new_P3_U3021;
  assign new_P3_U4339 = ~P3_REG2_REG_16_ | ~new_P3_U3020;
  assign new_P3_U4340 = ~new_P3_SUB_609_U7 | ~new_P3_U3019;
  assign new_P3_U4341 = ~new_P3_U3072;
  assign new_P3_U4342 = ~new_P3_U3033 | ~new_P3_U3078;
  assign new_P3_U4343 = ~new_P3_R1110_U111 | ~new_P3_U3883;
  assign new_P3_U4344 = ~new_P3_R1077_U111 | ~new_P3_U3885;
  assign new_P3_U4345 = ~new_P3_R1095_U114 | ~new_P3_U3884;
  assign new_P3_U4346 = ~new_P3_R1143_U111 | ~new_P3_U3881;
  assign new_P3_U4347 = ~new_P3_R1161_U111 | ~new_P3_U3891;
  assign new_P3_U4348 = ~new_P3_R1131_U114 | ~new_P3_U3887;
  assign new_P3_U4349 = ~new_P3_R1200_U114 | ~new_P3_U3017;
  assign new_P3_U4350 = ~new_P3_U3329;
  assign new_P3_U4351 = ~new_P3_R1179_U114 | ~new_P3_U3026;
  assign new_P3_U4352 = ~new_P3_U3025 | ~new_P3_U3072;
  assign new_P3_U4353 = ~new_P3_U3434 | ~new_P3_U4064;
  assign new_P3_U4354 = ~new_P3_U3641 | ~new_P3_U4350;
  assign new_P3_U4355 = ~P3_REG0_REG_17_ | ~new_P3_U3022;
  assign new_P3_U4356 = ~P3_REG1_REG_17_ | ~new_P3_U3021;
  assign new_P3_U4357 = ~P3_REG2_REG_17_ | ~new_P3_U3020;
  assign new_P3_U4358 = ~new_P3_SUB_609_U19 | ~new_P3_U3019;
  assign new_P3_U4359 = ~new_P3_U3068;
  assign new_P3_U4360 = ~new_P3_U3033 | ~new_P3_U3073;
  assign new_P3_U4361 = ~new_P3_R1110_U110 | ~new_P3_U3883;
  assign new_P3_U4362 = ~new_P3_R1077_U110 | ~new_P3_U3885;
  assign new_P3_U4363 = ~new_P3_R1095_U17 | ~new_P3_U3884;
  assign new_P3_U4364 = ~new_P3_R1143_U110 | ~new_P3_U3881;
  assign new_P3_U4365 = ~new_P3_R1161_U110 | ~new_P3_U3891;
  assign new_P3_U4366 = ~new_P3_R1131_U17 | ~new_P3_U3887;
  assign new_P3_U4367 = ~new_P3_R1200_U17 | ~new_P3_U3017;
  assign new_P3_U4368 = ~new_P3_U3330;
  assign new_P3_U4369 = ~new_P3_R1179_U17 | ~new_P3_U3026;
  assign new_P3_U4370 = ~new_P3_U3025 | ~new_P3_U3068;
  assign new_P3_U4371 = ~new_P3_U3437 | ~new_P3_U4064;
  assign new_P3_U4372 = ~new_P3_U3644 | ~new_P3_U4368;
  assign new_P3_U4373 = ~P3_REG0_REG_18_ | ~new_P3_U3022;
  assign new_P3_U4374 = ~P3_REG1_REG_18_ | ~new_P3_U3021;
  assign new_P3_U4375 = ~P3_REG2_REG_18_ | ~new_P3_U3020;
  assign new_P3_U4376 = ~new_P3_SUB_609_U11 | ~new_P3_U3019;
  assign new_P3_U4377 = ~new_P3_U3081;
  assign new_P3_U4378 = ~new_P3_U3033 | ~new_P3_U3072;
  assign new_P3_U4379 = ~new_P3_R1110_U12 | ~new_P3_U3883;
  assign new_P3_U4380 = ~new_P3_R1077_U12 | ~new_P3_U3885;
  assign new_P3_U4381 = ~new_P3_R1095_U103 | ~new_P3_U3884;
  assign new_P3_U4382 = ~new_P3_R1143_U12 | ~new_P3_U3881;
  assign new_P3_U4383 = ~new_P3_R1161_U12 | ~new_P3_U3891;
  assign new_P3_U4384 = ~new_P3_R1131_U103 | ~new_P3_U3887;
  assign new_P3_U4385 = ~new_P3_R1200_U103 | ~new_P3_U3017;
  assign new_P3_U4386 = ~new_P3_U3331;
  assign new_P3_U4387 = ~new_P3_R1179_U103 | ~new_P3_U3026;
  assign new_P3_U4388 = ~new_P3_U3025 | ~new_P3_U3081;
  assign new_P3_U4389 = ~new_P3_U3440 | ~new_P3_U4064;
  assign new_P3_U4390 = ~new_P3_U3648 | ~new_P3_U4386;
  assign new_P3_U4391 = ~P3_REG0_REG_19_ | ~new_P3_U3022;
  assign new_P3_U4392 = ~P3_REG1_REG_19_ | ~new_P3_U3021;
  assign new_P3_U4393 = ~P3_REG2_REG_19_ | ~new_P3_U3020;
  assign new_P3_U4394 = ~new_P3_SUB_609_U15 | ~new_P3_U3019;
  assign new_P3_U4395 = ~new_P3_U3080;
  assign new_P3_U4396 = ~new_P3_U3033 | ~new_P3_U3068;
  assign new_P3_U4397 = ~new_P3_R1110_U109 | ~new_P3_U3883;
  assign new_P3_U4398 = ~new_P3_R1077_U109 | ~new_P3_U3885;
  assign new_P3_U4399 = ~new_P3_R1095_U102 | ~new_P3_U3884;
  assign new_P3_U4400 = ~new_P3_R1143_U109 | ~new_P3_U3881;
  assign new_P3_U4401 = ~new_P3_R1161_U109 | ~new_P3_U3891;
  assign new_P3_U4402 = ~new_P3_R1131_U102 | ~new_P3_U3887;
  assign new_P3_U4403 = ~new_P3_R1200_U102 | ~new_P3_U3017;
  assign new_P3_U4404 = ~new_P3_U3332;
  assign new_P3_U4405 = ~new_P3_R1179_U102 | ~new_P3_U3026;
  assign new_P3_U4406 = ~new_P3_U3025 | ~new_P3_U3080;
  assign new_P3_U4407 = ~new_P3_U3443 | ~new_P3_U4064;
  assign new_P3_U4408 = ~new_P3_U3651 | ~new_P3_U4404;
  assign new_P3_U4409 = ~P3_REG2_REG_20_ | ~new_P3_U3020;
  assign new_P3_U4410 = ~P3_REG1_REG_20_ | ~new_P3_U3021;
  assign new_P3_U4411 = ~P3_REG0_REG_20_ | ~new_P3_U3022;
  assign new_P3_U4412 = ~new_P3_SUB_609_U20 | ~new_P3_U3019;
  assign new_P3_U4413 = ~new_P3_U3075;
  assign new_P3_U4414 = ~new_P3_U3033 | ~new_P3_U3081;
  assign new_P3_U4415 = ~new_P3_R1110_U108 | ~new_P3_U3883;
  assign new_P3_U4416 = ~new_P3_R1077_U108 | ~new_P3_U3885;
  assign new_P3_U4417 = ~new_P3_R1095_U101 | ~new_P3_U3884;
  assign new_P3_U4418 = ~new_P3_R1143_U108 | ~new_P3_U3881;
  assign new_P3_U4419 = ~new_P3_R1161_U108 | ~new_P3_U3891;
  assign new_P3_U4420 = ~new_P3_R1131_U101 | ~new_P3_U3887;
  assign new_P3_U4421 = ~new_P3_R1200_U101 | ~new_P3_U3017;
  assign new_P3_U4422 = ~new_P3_U3333;
  assign new_P3_U4423 = ~new_P3_R1179_U101 | ~new_P3_U3026;
  assign new_P3_U4424 = ~new_P3_U3025 | ~new_P3_U3075;
  assign new_P3_U4425 = ~new_P3_U3445 | ~new_P3_U4064;
  assign new_P3_U4426 = ~new_P3_U3654 | ~new_P3_U4422;
  assign new_P3_U4427 = ~P3_REG2_REG_21_ | ~new_P3_U3020;
  assign new_P3_U4428 = ~P3_REG1_REG_21_ | ~new_P3_U3021;
  assign new_P3_U4429 = ~P3_REG0_REG_21_ | ~new_P3_U3022;
  assign new_P3_U4430 = ~new_P3_SUB_609_U27 | ~new_P3_U3019;
  assign new_P3_U4431 = ~new_P3_U3074;
  assign new_P3_U4432 = ~new_P3_U3033 | ~new_P3_U3080;
  assign new_P3_U4433 = ~new_P3_R1110_U13 | ~new_P3_U3883;
  assign new_P3_U4434 = ~new_P3_R1077_U13 | ~new_P3_U3885;
  assign new_P3_U4435 = ~new_P3_R1095_U99 | ~new_P3_U3884;
  assign new_P3_U4436 = ~new_P3_R1143_U13 | ~new_P3_U3881;
  assign new_P3_U4437 = ~new_P3_R1161_U13 | ~new_P3_U3891;
  assign new_P3_U4438 = ~new_P3_R1131_U99 | ~new_P3_U3887;
  assign new_P3_U4439 = ~new_P3_R1200_U99 | ~new_P3_U3017;
  assign new_P3_U4440 = ~new_P3_U3335;
  assign new_P3_U4441 = ~new_P3_R1179_U99 | ~new_P3_U3026;
  assign new_P3_U4442 = ~new_P3_U3025 | ~new_P3_U3074;
  assign new_P3_U4443 = ~new_P3_U3907 | ~new_P3_U4064;
  assign new_P3_U4444 = ~new_P3_U3657 | ~new_P3_U4440;
  assign new_P3_U4445 = ~P3_REG2_REG_22_ | ~new_P3_U3020;
  assign new_P3_U4446 = ~P3_REG1_REG_22_ | ~new_P3_U3021;
  assign new_P3_U4447 = ~P3_REG0_REG_22_ | ~new_P3_U3022;
  assign new_P3_U4448 = ~new_P3_SUB_609_U17 | ~new_P3_U3019;
  assign new_P3_U4449 = ~new_P3_U3060;
  assign new_P3_U4450 = ~new_P3_U3033 | ~new_P3_U3075;
  assign new_P3_U4451 = ~new_P3_R1110_U14 | ~new_P3_U3883;
  assign new_P3_U4452 = ~new_P3_R1077_U14 | ~new_P3_U3885;
  assign new_P3_U4453 = ~new_P3_R1095_U113 | ~new_P3_U3884;
  assign new_P3_U4454 = ~new_P3_R1143_U14 | ~new_P3_U3881;
  assign new_P3_U4455 = ~new_P3_R1161_U14 | ~new_P3_U3891;
  assign new_P3_U4456 = ~new_P3_R1131_U113 | ~new_P3_U3887;
  assign new_P3_U4457 = ~new_P3_R1200_U113 | ~new_P3_U3017;
  assign new_P3_U4458 = ~new_P3_U3337;
  assign new_P3_U4459 = ~new_P3_R1179_U113 | ~new_P3_U3026;
  assign new_P3_U4460 = ~new_P3_U3025 | ~new_P3_U3060;
  assign new_P3_U4461 = ~new_P3_U3906 | ~new_P3_U4064;
  assign new_P3_U4462 = ~new_P3_U3660 | ~new_P3_U4458;
  assign new_P3_U4463 = ~P3_REG2_REG_23_ | ~new_P3_U3020;
  assign new_P3_U4464 = ~P3_REG1_REG_23_ | ~new_P3_U3021;
  assign new_P3_U4465 = ~P3_REG0_REG_23_ | ~new_P3_U3022;
  assign new_P3_U4466 = ~new_P3_SUB_609_U6 | ~new_P3_U3019;
  assign new_P3_U4467 = ~new_P3_U3065;
  assign new_P3_U4468 = ~new_P3_U3033 | ~new_P3_U3074;
  assign new_P3_U4469 = ~new_P3_R1110_U107 | ~new_P3_U3883;
  assign new_P3_U4470 = ~new_P3_R1077_U107 | ~new_P3_U3885;
  assign new_P3_U4471 = ~new_P3_R1095_U112 | ~new_P3_U3884;
  assign new_P3_U4472 = ~new_P3_R1143_U107 | ~new_P3_U3881;
  assign new_P3_U4473 = ~new_P3_R1161_U107 | ~new_P3_U3891;
  assign new_P3_U4474 = ~new_P3_R1131_U112 | ~new_P3_U3887;
  assign new_P3_U4475 = ~new_P3_R1200_U112 | ~new_P3_U3017;
  assign new_P3_U4476 = ~new_P3_U3339;
  assign new_P3_U4477 = ~new_P3_R1179_U112 | ~new_P3_U3026;
  assign new_P3_U4478 = ~new_P3_U3025 | ~new_P3_U3065;
  assign new_P3_U4479 = ~new_P3_U3905 | ~new_P3_U4064;
  assign new_P3_U4480 = ~new_P3_U3663 | ~new_P3_U4476;
  assign new_P3_U4481 = ~P3_REG2_REG_24_ | ~new_P3_U3020;
  assign new_P3_U4482 = ~P3_REG1_REG_24_ | ~new_P3_U3021;
  assign new_P3_U4483 = ~P3_REG0_REG_24_ | ~new_P3_U3022;
  assign new_P3_U4484 = ~new_P3_SUB_609_U10 | ~new_P3_U3019;
  assign new_P3_U4485 = ~new_P3_U3064;
  assign new_P3_U4486 = ~new_P3_U3033 | ~new_P3_U3060;
  assign new_P3_U4487 = ~new_P3_R1110_U106 | ~new_P3_U3883;
  assign new_P3_U4488 = ~new_P3_R1077_U106 | ~new_P3_U3885;
  assign new_P3_U4489 = ~new_P3_R1095_U18 | ~new_P3_U3884;
  assign new_P3_U4490 = ~new_P3_R1143_U106 | ~new_P3_U3881;
  assign new_P3_U4491 = ~new_P3_R1161_U106 | ~new_P3_U3891;
  assign new_P3_U4492 = ~new_P3_R1131_U18 | ~new_P3_U3887;
  assign new_P3_U4493 = ~new_P3_R1200_U18 | ~new_P3_U3017;
  assign new_P3_U4494 = ~new_P3_U3341;
  assign new_P3_U4495 = ~new_P3_R1179_U18 | ~new_P3_U3026;
  assign new_P3_U4496 = ~new_P3_U3025 | ~new_P3_U3064;
  assign new_P3_U4497 = ~new_P3_U3904 | ~new_P3_U4064;
  assign new_P3_U4498 = ~new_P3_U3666 | ~new_P3_U4494;
  assign new_P3_U4499 = ~P3_REG2_REG_25_ | ~new_P3_U3020;
  assign new_P3_U4500 = ~P3_REG1_REG_25_ | ~new_P3_U3021;
  assign new_P3_U4501 = ~P3_REG0_REG_25_ | ~new_P3_U3022;
  assign new_P3_U4502 = ~new_P3_SUB_609_U16 | ~new_P3_U3019;
  assign new_P3_U4503 = ~new_P3_U3057;
  assign new_P3_U4504 = ~new_P3_U3033 | ~new_P3_U3065;
  assign new_P3_U4505 = ~new_P3_R1110_U105 | ~new_P3_U3883;
  assign new_P3_U4506 = ~new_P3_R1077_U105 | ~new_P3_U3885;
  assign new_P3_U4507 = ~new_P3_R1095_U98 | ~new_P3_U3884;
  assign new_P3_U4508 = ~new_P3_R1143_U105 | ~new_P3_U3881;
  assign new_P3_U4509 = ~new_P3_R1161_U105 | ~new_P3_U3891;
  assign new_P3_U4510 = ~new_P3_R1131_U98 | ~new_P3_U3887;
  assign new_P3_U4511 = ~new_P3_R1200_U98 | ~new_P3_U3017;
  assign new_P3_U4512 = ~new_P3_U3343;
  assign new_P3_U4513 = ~new_P3_R1179_U98 | ~new_P3_U3026;
  assign new_P3_U4514 = ~new_P3_U3025 | ~new_P3_U3057;
  assign new_P3_U4515 = ~new_P3_U3903 | ~new_P3_U4064;
  assign new_P3_U4516 = ~new_P3_U3670 | ~new_P3_U4512;
  assign new_P3_U4517 = ~P3_REG2_REG_26_ | ~new_P3_U3020;
  assign new_P3_U4518 = ~P3_REG1_REG_26_ | ~new_P3_U3021;
  assign new_P3_U4519 = ~P3_REG0_REG_26_ | ~new_P3_U3022;
  assign new_P3_U4520 = ~new_P3_SUB_609_U26 | ~new_P3_U3019;
  assign new_P3_U4521 = ~new_P3_U3056;
  assign new_P3_U4522 = ~new_P3_U3033 | ~new_P3_U3064;
  assign new_P3_U4523 = ~new_P3_R1110_U104 | ~new_P3_U3883;
  assign new_P3_U4524 = ~new_P3_R1077_U104 | ~new_P3_U3885;
  assign new_P3_U4525 = ~new_P3_R1095_U97 | ~new_P3_U3884;
  assign new_P3_U4526 = ~new_P3_R1143_U104 | ~new_P3_U3881;
  assign new_P3_U4527 = ~new_P3_R1161_U104 | ~new_P3_U3891;
  assign new_P3_U4528 = ~new_P3_R1131_U97 | ~new_P3_U3887;
  assign new_P3_U4529 = ~new_P3_R1200_U97 | ~new_P3_U3017;
  assign new_P3_U4530 = ~new_P3_U3345;
  assign new_P3_U4531 = ~new_P3_R1179_U97 | ~new_P3_U3026;
  assign new_P3_U4532 = ~new_P3_U3025 | ~new_P3_U3056;
  assign new_P3_U4533 = ~new_P3_U3902 | ~new_P3_U4064;
  assign new_P3_U4534 = ~new_P3_U3674 | ~new_P3_U4530;
  assign new_P3_U4535 = ~P3_REG2_REG_27_ | ~new_P3_U3020;
  assign new_P3_U4536 = ~P3_REG1_REG_27_ | ~new_P3_U3021;
  assign new_P3_U4537 = ~P3_REG0_REG_27_ | ~new_P3_U3022;
  assign new_P3_U4538 = ~new_P3_SUB_609_U22 | ~new_P3_U3019;
  assign new_P3_U4539 = ~new_P3_U3052;
  assign new_P3_U4540 = ~new_P3_U3033 | ~new_P3_U3057;
  assign new_P3_U4541 = ~new_P3_R1110_U15 | ~new_P3_U3883;
  assign new_P3_U4542 = ~new_P3_R1077_U15 | ~new_P3_U3885;
  assign new_P3_U4543 = ~new_P3_R1095_U111 | ~new_P3_U3884;
  assign new_P3_U4544 = ~new_P3_R1143_U15 | ~new_P3_U3881;
  assign new_P3_U4545 = ~new_P3_R1161_U15 | ~new_P3_U3891;
  assign new_P3_U4546 = ~new_P3_R1131_U111 | ~new_P3_U3887;
  assign new_P3_U4547 = ~new_P3_R1200_U111 | ~new_P3_U3017;
  assign new_P3_U4548 = ~new_P3_U3347;
  assign new_P3_U4549 = ~new_P3_R1179_U111 | ~new_P3_U3026;
  assign new_P3_U4550 = ~new_P3_U3025 | ~new_P3_U3052;
  assign new_P3_U4551 = ~new_P3_U3901 | ~new_P3_U4064;
  assign new_P3_U4552 = ~new_P3_U3678 | ~new_P3_U4548;
  assign new_P3_U4553 = ~P3_REG2_REG_28_ | ~new_P3_U3020;
  assign new_P3_U4554 = ~P3_REG1_REG_28_ | ~new_P3_U3021;
  assign new_P3_U4555 = ~P3_REG0_REG_28_ | ~new_P3_U3022;
  assign new_P3_U4556 = ~new_P3_SUB_609_U28 | ~new_P3_U3019;
  assign new_P3_U4557 = ~new_P3_U3053;
  assign new_P3_U4558 = ~new_P3_U3033 | ~new_P3_U3056;
  assign new_P3_U4559 = ~new_P3_R1110_U103 | ~new_P3_U3883;
  assign new_P3_U4560 = ~new_P3_R1077_U103 | ~new_P3_U3885;
  assign new_P3_U4561 = ~new_P3_R1095_U19 | ~new_P3_U3884;
  assign new_P3_U4562 = ~new_P3_R1143_U103 | ~new_P3_U3881;
  assign new_P3_U4563 = ~new_P3_R1161_U103 | ~new_P3_U3891;
  assign new_P3_U4564 = ~new_P3_R1131_U19 | ~new_P3_U3887;
  assign new_P3_U4565 = ~new_P3_R1200_U19 | ~new_P3_U3017;
  assign new_P3_U4566 = ~new_P3_U3349;
  assign new_P3_U4567 = ~new_P3_R1179_U19 | ~new_P3_U3026;
  assign new_P3_U4568 = ~new_P3_U3025 | ~new_P3_U3053;
  assign new_P3_U4569 = ~new_P3_U3900 | ~new_P3_U4064;
  assign new_P3_U4570 = ~new_P3_U3682 | ~new_P3_U4566;
  assign new_P3_U4571 = ~new_P3_SUB_609_U92 | ~new_P3_U3019;
  assign new_P3_U4572 = ~P3_REG2_REG_29_ | ~new_P3_U3020;
  assign new_P3_U4573 = ~P3_REG1_REG_29_ | ~new_P3_U3021;
  assign new_P3_U4574 = ~P3_REG0_REG_29_ | ~new_P3_U3022;
  assign new_P3_U4575 = ~new_P3_U3054;
  assign new_P3_U4576 = ~new_P3_U3033 | ~new_P3_U3052;
  assign new_P3_U4577 = ~new_P3_R1110_U102 | ~new_P3_U3883;
  assign new_P3_U4578 = ~new_P3_R1077_U102 | ~new_P3_U3885;
  assign new_P3_U4579 = ~new_P3_R1095_U96 | ~new_P3_U3884;
  assign new_P3_U4580 = ~new_P3_R1143_U102 | ~new_P3_U3881;
  assign new_P3_U4581 = ~new_P3_R1161_U102 | ~new_P3_U3891;
  assign new_P3_U4582 = ~new_P3_R1131_U96 | ~new_P3_U3887;
  assign new_P3_U4583 = ~new_P3_R1200_U96 | ~new_P3_U3017;
  assign new_P3_U4584 = ~new_P3_U3351;
  assign new_P3_U4585 = ~new_P3_R1179_U96 | ~new_P3_U3026;
  assign new_P3_U4586 = ~new_P3_U3025 | ~new_P3_U3054;
  assign new_P3_U4587 = ~new_P3_U3899 | ~new_P3_U4064;
  assign new_P3_U4588 = ~new_P3_U3686 | ~new_P3_U4584;
  assign new_P3_U4589 = ~P3_REG2_REG_30_ | ~new_P3_U3020;
  assign new_P3_U4590 = ~P3_REG1_REG_30_ | ~new_P3_U3021;
  assign new_P3_U4591 = ~P3_REG0_REG_30_ | ~new_P3_U3022;
  assign new_P3_U4592 = ~new_P3_SUB_609_U92 | ~new_P3_U3019;
  assign new_P3_U4593 = ~new_P3_U3058;
  assign new_P3_U4594 = ~new_P3_U3892 | ~new_P3_U3298;
  assign new_P3_U4595 = ~new_P3_U3833 | ~new_P3_U4594;
  assign new_P3_U4596 = ~new_P3_U3058 | ~new_P3_U4595 | ~new_P3_U3911;
  assign new_P3_U4597 = ~new_P3_U3033 | ~new_P3_U3053;
  assign new_P3_U4598 = ~new_P3_R1110_U101 | ~new_P3_U3883;
  assign new_P3_U4599 = ~new_P3_R1077_U101 | ~new_P3_U3885;
  assign new_P3_U4600 = ~new_P3_R1095_U20 | ~new_P3_U3884;
  assign new_P3_U4601 = ~new_P3_R1143_U101 | ~new_P3_U3881;
  assign new_P3_U4602 = ~new_P3_R1161_U101 | ~new_P3_U3891;
  assign new_P3_U4603 = ~new_P3_R1131_U20 | ~new_P3_U3887;
  assign new_P3_U4604 = ~new_P3_R1200_U20 | ~new_P3_U3017;
  assign new_P3_U4605 = ~new_P3_U3354;
  assign new_P3_U4606 = ~new_P3_R1179_U20 | ~new_P3_U3026;
  assign new_P3_U4607 = ~new_P3_U3908 | ~new_P3_U4064;
  assign new_P3_U4608 = ~new_P3_U3690 | ~new_P3_U4605;
  assign new_P3_U4609 = ~new_P3_SUB_609_U92 | ~new_P3_U3019;
  assign new_P3_U4610 = ~P3_REG2_REG_31_ | ~new_P3_U3020;
  assign new_P3_U4611 = ~P3_REG1_REG_31_ | ~new_P3_U3021;
  assign new_P3_U4612 = ~P3_REG0_REG_31_ | ~new_P3_U3022;
  assign new_P3_U4613 = ~new_P3_U3055;
  assign new_P3_U4614 = ~new_P3_U3873 | ~new_P3_U4064;
  assign new_P3_U4615 = ~new_P3_U3361 | ~new_P3_U4614;
  assign new_P3_U4616 = ~new_P3_U3872 | ~new_P3_U4064;
  assign new_P3_U4617 = ~new_P3_U3361 | ~new_P3_U4616;
  assign new_P3_U4618 = ~new_P3_U3302 | ~new_P3_U5641 | ~new_P3_U5640;
  assign new_P3_U4619 = ~new_P3_U3888 | ~new_P3_U3367;
  assign new_P3_U4620 = ~new_P3_U3048 | ~new_P3_U4619;
  assign new_P3_U4621 = ~new_P3_U3047 | ~new_P3_U4618;
  assign new_P3_U4622 = ~new_P3_U4621 | ~new_P3_U4620;
  assign new_P3_U4623 = ~new_P3_U5456 | ~new_P3_U3379;
  assign new_P3_U4624 = ~new_P3_U3834 | ~new_P3_U4623 | ~new_P3_U3380;
  assign new_P3_U4625 = ~new_P3_U3048 | ~new_P3_U4624;
  assign new_P3_U4626 = ~new_P3_U3047 | ~new_P3_U4619;
  assign new_P3_U4627 = ~new_P3_U4626 | ~new_P3_U4625 | ~new_P3_U3360;
  assign new_P3_U4628 = ~new_P3_U3365;
  assign new_P3_U4629 = ~new_P3_U3034 | ~new_P3_U3077;
  assign new_P3_U4630 = ~new_P3_U3030 | ~new_P3_R1179_U24;
  assign new_P3_U4631 = ~new_P3_U3029 | ~new_P3_U3387;
  assign new_P3_U4632 = ~new_P3_U3028 | ~P3_REG3_REG_0_;
  assign new_P3_U4633 = ~new_P3_U3034 | ~new_P3_U3067;
  assign new_P3_U4634 = ~new_P3_U3030 | ~new_P3_R1179_U100;
  assign new_P3_U4635 = ~new_P3_U3029 | ~new_P3_U3392;
  assign new_P3_U4636 = ~new_P3_U3028 | ~P3_REG3_REG_1_;
  assign new_P3_U4637 = ~new_P3_U3034 | ~new_P3_U3063;
  assign new_P3_U4638 = ~new_P3_U3030 | ~new_P3_R1179_U110;
  assign new_P3_U4639 = ~new_P3_U3029 | ~new_P3_U3395;
  assign new_P3_U4640 = ~new_P3_U3028 | ~P3_REG3_REG_2_;
  assign new_P3_U4641 = ~new_P3_U3034 | ~new_P3_U3059;
  assign new_P3_U4642 = ~new_P3_U3030 | ~new_P3_R1179_U21;
  assign new_P3_U4643 = ~new_P3_U3029 | ~new_P3_U3398;
  assign new_P3_U4644 = ~new_P3_U3028 | ~new_P3_SUB_609_U25;
  assign new_P3_U4645 = ~new_P3_U3034 | ~new_P3_U3066;
  assign new_P3_U4646 = ~new_P3_U3030 | ~new_P3_R1179_U109;
  assign new_P3_U4647 = ~new_P3_U3029 | ~new_P3_U3401;
  assign new_P3_U4648 = ~new_P3_U3028 | ~new_P3_SUB_609_U29;
  assign new_P3_U4649 = ~new_P3_U3034 | ~new_P3_U3070;
  assign new_P3_U4650 = ~new_P3_U3030 | ~new_P3_R1179_U108;
  assign new_P3_U4651 = ~new_P3_U3029 | ~new_P3_U3404;
  assign new_P3_U4652 = ~new_P3_U3028 | ~new_P3_SUB_609_U53;
  assign new_P3_U4653 = ~new_P3_U3034 | ~new_P3_U3069;
  assign new_P3_U4654 = ~new_P3_U3030 | ~new_P3_R1179_U22;
  assign new_P3_U4655 = ~new_P3_U3029 | ~new_P3_U3407;
  assign new_P3_U4656 = ~new_P3_U3028 | ~new_P3_SUB_609_U8;
  assign new_P3_U4657 = ~new_P3_U3034 | ~new_P3_U3083;
  assign new_P3_U4658 = ~new_P3_U3030 | ~new_P3_R1179_U107;
  assign new_P3_U4659 = ~new_P3_U3029 | ~new_P3_U3410;
  assign new_P3_U4660 = ~new_P3_U3028 | ~new_P3_SUB_609_U18;
  assign new_P3_U4661 = ~new_P3_U3034 | ~new_P3_U3082;
  assign new_P3_U4662 = ~new_P3_U3030 | ~new_P3_R1179_U23;
  assign new_P3_U4663 = ~new_P3_U3029 | ~new_P3_U3413;
  assign new_P3_U4664 = ~new_P3_U3028 | ~new_P3_SUB_609_U12;
  assign new_P3_U4665 = ~new_P3_U3034 | ~new_P3_U3061;
  assign new_P3_U4666 = ~new_P3_U3030 | ~new_P3_R1179_U106;
  assign new_P3_U4667 = ~new_P3_U3029 | ~new_P3_U3416;
  assign new_P3_U4668 = ~new_P3_U3028 | ~new_P3_SUB_609_U14;
  assign new_P3_U4669 = ~new_P3_U3034 | ~new_P3_U3062;
  assign new_P3_U4670 = ~new_P3_U3030 | ~new_P3_R1179_U116;
  assign new_P3_U4671 = ~new_P3_U3029 | ~new_P3_U3419;
  assign new_P3_U4672 = ~new_P3_U3028 | ~new_P3_SUB_609_U13;
  assign new_P3_U4673 = ~new_P3_U3034 | ~new_P3_U3071;
  assign new_P3_U4674 = ~new_P3_U3030 | ~new_P3_R1179_U16;
  assign new_P3_U4675 = ~new_P3_U3029 | ~new_P3_U3422;
  assign new_P3_U4676 = ~new_P3_U3028 | ~new_P3_SUB_609_U9;
  assign new_P3_U4677 = ~new_P3_U3034 | ~new_P3_U3079;
  assign new_P3_U4678 = ~new_P3_U3030 | ~new_P3_R1179_U105;
  assign new_P3_U4679 = ~new_P3_U3029 | ~new_P3_U3425;
  assign new_P3_U4680 = ~new_P3_U3028 | ~new_P3_SUB_609_U23;
  assign new_P3_U4681 = ~new_P3_U3034 | ~new_P3_U3078;
  assign new_P3_U4682 = ~new_P3_U3030 | ~new_P3_R1179_U104;
  assign new_P3_U4683 = ~new_P3_U3029 | ~new_P3_U3428;
  assign new_P3_U4684 = ~new_P3_U3028 | ~new_P3_SUB_609_U24;
  assign new_P3_U4685 = ~new_P3_U3034 | ~new_P3_U3073;
  assign new_P3_U4686 = ~new_P3_U3030 | ~new_P3_R1179_U115;
  assign new_P3_U4687 = ~new_P3_U3029 | ~new_P3_U3431;
  assign new_P3_U4688 = ~new_P3_U3028 | ~new_P3_SUB_609_U30;
  assign new_P3_U4689 = ~new_P3_U3034 | ~new_P3_U3072;
  assign new_P3_U4690 = ~new_P3_U3030 | ~new_P3_R1179_U114;
  assign new_P3_U4691 = ~new_P3_U3029 | ~new_P3_U3434;
  assign new_P3_U4692 = ~new_P3_U3028 | ~new_P3_SUB_609_U21;
  assign new_P3_U4693 = ~new_P3_U3034 | ~new_P3_U3068;
  assign new_P3_U4694 = ~new_P3_U3030 | ~new_P3_R1179_U17;
  assign new_P3_U4695 = ~new_P3_U3029 | ~new_P3_U3437;
  assign new_P3_U4696 = ~new_P3_U3028 | ~new_P3_SUB_609_U7;
  assign new_P3_U4697 = ~new_P3_U3034 | ~new_P3_U3081;
  assign new_P3_U4698 = ~new_P3_U3030 | ~new_P3_R1179_U103;
  assign new_P3_U4699 = ~new_P3_U3029 | ~new_P3_U3440;
  assign new_P3_U4700 = ~new_P3_U3028 | ~new_P3_SUB_609_U19;
  assign new_P3_U4701 = ~new_P3_U3034 | ~new_P3_U3080;
  assign new_P3_U4702 = ~new_P3_U3030 | ~new_P3_R1179_U102;
  assign new_P3_U4703 = ~new_P3_U3029 | ~new_P3_U3443;
  assign new_P3_U4704 = ~new_P3_U3028 | ~new_P3_SUB_609_U11;
  assign new_P3_U4705 = ~new_P3_U3034 | ~new_P3_U3075;
  assign new_P3_U4706 = ~new_P3_U3030 | ~new_P3_R1179_U101;
  assign new_P3_U4707 = ~new_P3_U3029 | ~new_P3_U3445;
  assign new_P3_U4708 = ~new_P3_U3028 | ~new_P3_SUB_609_U15;
  assign new_P3_U4709 = ~new_P3_U3034 | ~new_P3_U3074;
  assign new_P3_U4710 = ~new_P3_U3030 | ~new_P3_R1179_U99;
  assign new_P3_U4711 = ~new_P3_U3029 | ~new_P3_U3907;
  assign new_P3_U4712 = ~new_P3_U3028 | ~new_P3_SUB_609_U20;
  assign new_P3_U4713 = ~new_P3_U3034 | ~new_P3_U3060;
  assign new_P3_U4714 = ~new_P3_U3030 | ~new_P3_R1179_U113;
  assign new_P3_U4715 = ~new_P3_U3029 | ~new_P3_U3906;
  assign new_P3_U4716 = ~new_P3_U3028 | ~new_P3_SUB_609_U27;
  assign new_P3_U4717 = ~new_P3_U3034 | ~new_P3_U3065;
  assign new_P3_U4718 = ~new_P3_U3030 | ~new_P3_R1179_U112;
  assign new_P3_U4719 = ~new_P3_U3029 | ~new_P3_U3905;
  assign new_P3_U4720 = ~new_P3_U3028 | ~new_P3_SUB_609_U17;
  assign new_P3_U4721 = ~new_P3_U3034 | ~new_P3_U3064;
  assign new_P3_U4722 = ~new_P3_U3030 | ~new_P3_R1179_U18;
  assign new_P3_U4723 = ~new_P3_U3029 | ~new_P3_U3904;
  assign new_P3_U4724 = ~new_P3_U3028 | ~new_P3_SUB_609_U6;
  assign new_P3_U4725 = ~new_P3_U3034 | ~new_P3_U3057;
  assign new_P3_U4726 = ~new_P3_U3030 | ~new_P3_R1179_U98;
  assign new_P3_U4727 = ~new_P3_U3029 | ~new_P3_U3903;
  assign new_P3_U4728 = ~new_P3_U3028 | ~new_P3_SUB_609_U10;
  assign new_P3_U4729 = ~new_P3_U3034 | ~new_P3_U3056;
  assign new_P3_U4730 = ~new_P3_U3030 | ~new_P3_R1179_U97;
  assign new_P3_U4731 = ~new_P3_U3029 | ~new_P3_U3902;
  assign new_P3_U4732 = ~new_P3_U3028 | ~new_P3_SUB_609_U16;
  assign new_P3_U4733 = ~new_P3_U3034 | ~new_P3_U3052;
  assign new_P3_U4734 = ~new_P3_U3030 | ~new_P3_R1179_U111;
  assign new_P3_U4735 = ~new_P3_U3029 | ~new_P3_U3901;
  assign new_P3_U4736 = ~new_P3_U3028 | ~new_P3_SUB_609_U26;
  assign new_P3_U4737 = ~new_P3_U3034 | ~new_P3_U3053;
  assign new_P3_U4738 = ~new_P3_U3030 | ~new_P3_R1179_U19;
  assign new_P3_U4739 = ~new_P3_U3029 | ~new_P3_U3900;
  assign new_P3_U4740 = ~new_P3_U3028 | ~new_P3_SUB_609_U22;
  assign new_P3_U4741 = ~new_P3_U3034 | ~new_P3_U3054;
  assign new_P3_U4742 = ~new_P3_U3030 | ~new_P3_R1179_U96;
  assign new_P3_U4743 = ~new_P3_U3029 | ~new_P3_U3899;
  assign new_P3_U4744 = ~new_P3_U3028 | ~new_P3_SUB_609_U28;
  assign new_P3_U4745 = ~new_P3_U3030 | ~new_P3_R1179_U20;
  assign new_P3_U4746 = ~new_P3_U3029 | ~new_P3_U3908;
  assign new_P3_U4747 = ~new_P3_U3028 | ~new_P3_SUB_609_U92;
  assign new_P3_U4748 = ~new_P3_U3028 | ~new_P3_SUB_609_U92;
  assign new_P3_U4749 = ~new_P3_U3916 | ~new_P3_U3912;
  assign new_P3_U4750 = ~new_P3_U3029 | ~new_P3_U3873;
  assign new_P3_U4751 = ~P3_REG2_REG_30_ | ~new_P3_U3358;
  assign new_P3_U4752 = ~new_P3_U3029 | ~new_P3_U3872;
  assign new_P3_U4753 = ~P3_REG2_REG_31_ | ~new_P3_U3358;
  assign new_P3_U4754 = ~new_P3_U3697 | ~new_P3_U3698 | ~new_P3_U4628 | ~new_P3_U3359;
  assign new_P3_U4755 = ~new_P3_R1212_U6 | ~new_P3_U3040;
  assign new_P3_U4756 = ~new_P3_U3039 | ~new_P3_U3379;
  assign new_P3_U4757 = ~new_P3_R1209_U6 | ~new_P3_U3037;
  assign new_P3_U4758 = ~new_P3_U4757 | ~new_P3_U4756 | ~new_P3_U4755;
  assign new_P3_U4759 = ~new_P3_U3910 | ~new_P3_U5440;
  assign new_P3_U4760 = ~new_P3_U3366;
  assign new_P3_U4761 = ~new_P3_U3833 | ~new_P3_U3896;
  assign new_P3_U4762 = ~new_P3_R1054_U67 | ~new_P3_U3051;
  assign new_P3_U4763 = ~new_P3_U5768 | ~new_P3_U3379;
  assign new_P3_U4764 = ~new_P3_U3042 | ~new_P3_U4758;
  assign new_P3_U4765 = ~new_P3_U3041 | ~new_P3_R1212_U6;
  assign new_P3_U4766 = ~P3_REG3_REG_19_ | ~n3834;
  assign new_P3_U4767 = ~new_P3_U3038 | ~new_P3_R1209_U6;
  assign new_P3_U4768 = ~P3_ADDR_REG_19_ | ~new_P3_U4760;
  assign new_P3_U4769 = ~new_P3_R1212_U58 | ~new_P3_U3040;
  assign new_P3_U4770 = ~new_P3_U3039 | ~new_P3_U3442;
  assign new_P3_U4771 = ~new_P3_R1209_U58 | ~new_P3_U3037;
  assign new_P3_U4772 = ~new_P3_U4771 | ~new_P3_U4770 | ~new_P3_U4769;
  assign new_P3_U4773 = ~new_P3_R1054_U68 | ~new_P3_U3051;
  assign new_P3_U4774 = ~new_P3_U5768 | ~new_P3_U3442;
  assign new_P3_U4775 = ~new_P3_U3042 | ~new_P3_U4772;
  assign new_P3_U4776 = ~new_P3_R1212_U58 | ~new_P3_U3041;
  assign new_P3_U4777 = ~P3_REG3_REG_18_ | ~n3834;
  assign new_P3_U4778 = ~new_P3_R1209_U58 | ~new_P3_U3038;
  assign new_P3_U4779 = ~P3_ADDR_REG_18_ | ~new_P3_U4760;
  assign new_P3_U4780 = ~new_P3_R1212_U59 | ~new_P3_U3040;
  assign new_P3_U4781 = ~new_P3_U3039 | ~new_P3_U3439;
  assign new_P3_U4782 = ~new_P3_R1209_U59 | ~new_P3_U3037;
  assign new_P3_U4783 = ~new_P3_U4782 | ~new_P3_U4781 | ~new_P3_U4780;
  assign new_P3_U4784 = ~new_P3_R1054_U69 | ~new_P3_U3051;
  assign new_P3_U4785 = ~new_P3_U5768 | ~new_P3_U3439;
  assign new_P3_U4786 = ~new_P3_U3042 | ~new_P3_U4783;
  assign new_P3_U4787 = ~new_P3_R1212_U59 | ~new_P3_U3041;
  assign new_P3_U4788 = ~P3_REG3_REG_17_ | ~n3834;
  assign new_P3_U4789 = ~new_P3_R1209_U59 | ~new_P3_U3038;
  assign new_P3_U4790 = ~P3_ADDR_REG_17_ | ~new_P3_U4760;
  assign new_P3_U4791 = ~new_P3_R1212_U60 | ~new_P3_U3040;
  assign new_P3_U4792 = ~new_P3_U3039 | ~new_P3_U3436;
  assign new_P3_U4793 = ~new_P3_R1209_U60 | ~new_P3_U3037;
  assign new_P3_U4794 = ~new_P3_U4793 | ~new_P3_U4792 | ~new_P3_U4791;
  assign new_P3_U4795 = ~new_P3_R1054_U13 | ~new_P3_U3051;
  assign new_P3_U4796 = ~new_P3_U5768 | ~new_P3_U3436;
  assign new_P3_U4797 = ~new_P3_U3042 | ~new_P3_U4794;
  assign new_P3_U4798 = ~new_P3_R1212_U60 | ~new_P3_U3041;
  assign new_P3_U4799 = ~P3_REG3_REG_16_ | ~n3834;
  assign new_P3_U4800 = ~new_P3_R1209_U60 | ~new_P3_U3038;
  assign new_P3_U4801 = ~P3_ADDR_REG_16_ | ~new_P3_U4760;
  assign new_P3_U4802 = ~new_P3_R1212_U61 | ~new_P3_U3040;
  assign new_P3_U4803 = ~new_P3_U3039 | ~new_P3_U3433;
  assign new_P3_U4804 = ~new_P3_R1209_U61 | ~new_P3_U3037;
  assign new_P3_U4805 = ~new_P3_U4804 | ~new_P3_U4803 | ~new_P3_U4802;
  assign new_P3_U4806 = ~new_P3_R1054_U77 | ~new_P3_U3051;
  assign new_P3_U4807 = ~new_P3_U5768 | ~new_P3_U3433;
  assign new_P3_U4808 = ~new_P3_U3042 | ~new_P3_U4805;
  assign new_P3_U4809 = ~new_P3_R1212_U61 | ~new_P3_U3041;
  assign new_P3_U4810 = ~P3_REG3_REG_15_ | ~n3834;
  assign new_P3_U4811 = ~new_P3_R1209_U61 | ~new_P3_U3038;
  assign new_P3_U4812 = ~P3_ADDR_REG_15_ | ~new_P3_U4760;
  assign new_P3_U4813 = ~new_P3_R1212_U62 | ~new_P3_U3040;
  assign new_P3_U4814 = ~new_P3_U3039 | ~new_P3_U3430;
  assign new_P3_U4815 = ~new_P3_R1209_U62 | ~new_P3_U3037;
  assign new_P3_U4816 = ~new_P3_U4815 | ~new_P3_U4814 | ~new_P3_U4813;
  assign new_P3_U4817 = ~new_P3_R1054_U78 | ~new_P3_U3051;
  assign new_P3_U4818 = ~new_P3_U5768 | ~new_P3_U3430;
  assign new_P3_U4819 = ~new_P3_U3042 | ~new_P3_U4816;
  assign new_P3_U4820 = ~new_P3_R1212_U62 | ~new_P3_U3041;
  assign new_P3_U4821 = ~P3_REG3_REG_14_ | ~n3834;
  assign new_P3_U4822 = ~new_P3_R1209_U62 | ~new_P3_U3038;
  assign new_P3_U4823 = ~P3_ADDR_REG_14_ | ~new_P3_U4760;
  assign new_P3_U4824 = ~new_P3_R1212_U63 | ~new_P3_U3040;
  assign new_P3_U4825 = ~new_P3_U3039 | ~new_P3_U3427;
  assign new_P3_U4826 = ~new_P3_R1209_U63 | ~new_P3_U3037;
  assign new_P3_U4827 = ~new_P3_U4826 | ~new_P3_U4825 | ~new_P3_U4824;
  assign new_P3_U4828 = ~new_P3_R1054_U70 | ~new_P3_U3051;
  assign new_P3_U4829 = ~new_P3_U5768 | ~new_P3_U3427;
  assign new_P3_U4830 = ~new_P3_U3042 | ~new_P3_U4827;
  assign new_P3_U4831 = ~new_P3_R1212_U63 | ~new_P3_U3041;
  assign new_P3_U4832 = ~P3_REG3_REG_13_ | ~n3834;
  assign new_P3_U4833 = ~new_P3_R1209_U63 | ~new_P3_U3038;
  assign new_P3_U4834 = ~P3_ADDR_REG_13_ | ~new_P3_U4760;
  assign new_P3_U4835 = ~new_P3_R1212_U64 | ~new_P3_U3040;
  assign new_P3_U4836 = ~new_P3_U3039 | ~new_P3_U3424;
  assign new_P3_U4837 = ~new_P3_R1209_U64 | ~new_P3_U3037;
  assign new_P3_U4838 = ~new_P3_U4837 | ~new_P3_U4836 | ~new_P3_U4835;
  assign new_P3_U4839 = ~new_P3_R1054_U71 | ~new_P3_U3051;
  assign new_P3_U4840 = ~new_P3_U5768 | ~new_P3_U3424;
  assign new_P3_U4841 = ~new_P3_U3042 | ~new_P3_U4838;
  assign new_P3_U4842 = ~new_P3_R1212_U64 | ~new_P3_U3041;
  assign new_P3_U4843 = ~P3_REG3_REG_12_ | ~n3834;
  assign new_P3_U4844 = ~new_P3_R1209_U64 | ~new_P3_U3038;
  assign new_P3_U4845 = ~P3_ADDR_REG_12_ | ~new_P3_U4760;
  assign new_P3_U4846 = ~new_P3_R1212_U65 | ~new_P3_U3040;
  assign new_P3_U4847 = ~new_P3_U3039 | ~new_P3_U3421;
  assign new_P3_U4848 = ~new_P3_R1209_U65 | ~new_P3_U3037;
  assign new_P3_U4849 = ~new_P3_U4848 | ~new_P3_U4847 | ~new_P3_U4846;
  assign new_P3_U4850 = ~new_P3_R1054_U12 | ~new_P3_U3051;
  assign new_P3_U4851 = ~new_P3_U5768 | ~new_P3_U3421;
  assign new_P3_U4852 = ~new_P3_U3042 | ~new_P3_U4849;
  assign new_P3_U4853 = ~new_P3_R1212_U65 | ~new_P3_U3041;
  assign new_P3_U4854 = ~P3_REG3_REG_11_ | ~n3834;
  assign new_P3_U4855 = ~new_P3_R1209_U65 | ~new_P3_U3038;
  assign new_P3_U4856 = ~P3_ADDR_REG_11_ | ~new_P3_U4760;
  assign new_P3_U4857 = ~new_P3_R1212_U66 | ~new_P3_U3040;
  assign new_P3_U4858 = ~new_P3_U3039 | ~new_P3_U3418;
  assign new_P3_U4859 = ~new_P3_R1209_U66 | ~new_P3_U3037;
  assign new_P3_U4860 = ~new_P3_U4859 | ~new_P3_U4858 | ~new_P3_U4857;
  assign new_P3_U4861 = ~new_P3_R1054_U79 | ~new_P3_U3051;
  assign new_P3_U4862 = ~new_P3_U5768 | ~new_P3_U3418;
  assign new_P3_U4863 = ~new_P3_U3042 | ~new_P3_U4860;
  assign new_P3_U4864 = ~new_P3_R1212_U66 | ~new_P3_U3041;
  assign new_P3_U4865 = ~P3_REG3_REG_10_ | ~n3834;
  assign new_P3_U4866 = ~new_P3_R1209_U66 | ~new_P3_U3038;
  assign new_P3_U4867 = ~P3_ADDR_REG_10_ | ~new_P3_U4760;
  assign new_P3_U4868 = ~new_P3_R1212_U49 | ~new_P3_U3040;
  assign new_P3_U4869 = ~new_P3_U3039 | ~new_P3_U3415;
  assign new_P3_U4870 = ~new_P3_R1209_U49 | ~new_P3_U3037;
  assign new_P3_U4871 = ~new_P3_U4870 | ~new_P3_U4869 | ~new_P3_U4868;
  assign new_P3_U4872 = ~new_P3_R1054_U72 | ~new_P3_U3051;
  assign new_P3_U4873 = ~new_P3_U5768 | ~new_P3_U3415;
  assign new_P3_U4874 = ~new_P3_U3042 | ~new_P3_U4871;
  assign new_P3_U4875 = ~new_P3_R1212_U49 | ~new_P3_U3041;
  assign new_P3_U4876 = ~P3_REG3_REG_9_ | ~n3834;
  assign new_P3_U4877 = ~new_P3_R1209_U49 | ~new_P3_U3038;
  assign new_P3_U4878 = ~P3_ADDR_REG_9_ | ~new_P3_U4760;
  assign new_P3_U4879 = ~new_P3_R1212_U50 | ~new_P3_U3040;
  assign new_P3_U4880 = ~new_P3_U3039 | ~new_P3_U3412;
  assign new_P3_U4881 = ~new_P3_R1209_U50 | ~new_P3_U3037;
  assign new_P3_U4882 = ~new_P3_U4881 | ~new_P3_U4880 | ~new_P3_U4879;
  assign new_P3_U4883 = ~new_P3_R1054_U16 | ~new_P3_U3051;
  assign new_P3_U4884 = ~new_P3_U5768 | ~new_P3_U3412;
  assign new_P3_U4885 = ~new_P3_U3042 | ~new_P3_U4882;
  assign new_P3_U4886 = ~new_P3_R1212_U50 | ~new_P3_U3041;
  assign new_P3_U4887 = ~P3_REG3_REG_8_ | ~n3834;
  assign new_P3_U4888 = ~new_P3_R1209_U50 | ~new_P3_U3038;
  assign new_P3_U4889 = ~P3_ADDR_REG_8_ | ~new_P3_U4760;
  assign new_P3_U4890 = ~new_P3_R1212_U51 | ~new_P3_U3040;
  assign new_P3_U4891 = ~new_P3_U3039 | ~new_P3_U3409;
  assign new_P3_U4892 = ~new_P3_R1209_U51 | ~new_P3_U3037;
  assign new_P3_U4893 = ~new_P3_U4892 | ~new_P3_U4891 | ~new_P3_U4890;
  assign new_P3_U4894 = ~new_P3_R1054_U73 | ~new_P3_U3051;
  assign new_P3_U4895 = ~new_P3_U5768 | ~new_P3_U3409;
  assign new_P3_U4896 = ~new_P3_U3042 | ~new_P3_U4893;
  assign new_P3_U4897 = ~new_P3_R1212_U51 | ~new_P3_U3041;
  assign new_P3_U4898 = ~P3_REG3_REG_7_ | ~n3834;
  assign new_P3_U4899 = ~new_P3_R1209_U51 | ~new_P3_U3038;
  assign new_P3_U4900 = ~P3_ADDR_REG_7_ | ~new_P3_U4760;
  assign new_P3_U4901 = ~new_P3_R1212_U52 | ~new_P3_U3040;
  assign new_P3_U4902 = ~new_P3_U3039 | ~new_P3_U3406;
  assign new_P3_U4903 = ~new_P3_R1209_U52 | ~new_P3_U3037;
  assign new_P3_U4904 = ~new_P3_U4903 | ~new_P3_U4902 | ~new_P3_U4901;
  assign new_P3_U4905 = ~new_P3_R1054_U15 | ~new_P3_U3051;
  assign new_P3_U4906 = ~new_P3_U5768 | ~new_P3_U3406;
  assign new_P3_U4907 = ~new_P3_U3042 | ~new_P3_U4904;
  assign new_P3_U4908 = ~new_P3_R1212_U52 | ~new_P3_U3041;
  assign new_P3_U4909 = ~P3_REG3_REG_6_ | ~n3834;
  assign new_P3_U4910 = ~new_P3_R1209_U52 | ~new_P3_U3038;
  assign new_P3_U4911 = ~P3_ADDR_REG_6_ | ~new_P3_U4760;
  assign new_P3_U4912 = ~new_P3_R1212_U53 | ~new_P3_U3040;
  assign new_P3_U4913 = ~new_P3_U3039 | ~new_P3_U3403;
  assign new_P3_U4914 = ~new_P3_R1209_U53 | ~new_P3_U3037;
  assign new_P3_U4915 = ~new_P3_U4914 | ~new_P3_U4913 | ~new_P3_U4912;
  assign new_P3_U4916 = ~new_P3_R1054_U74 | ~new_P3_U3051;
  assign new_P3_U4917 = ~new_P3_U5768 | ~new_P3_U3403;
  assign new_P3_U4918 = ~new_P3_U3042 | ~new_P3_U4915;
  assign new_P3_U4919 = ~new_P3_R1212_U53 | ~new_P3_U3041;
  assign new_P3_U4920 = ~P3_REG3_REG_5_ | ~n3834;
  assign new_P3_U4921 = ~new_P3_R1209_U53 | ~new_P3_U3038;
  assign new_P3_U4922 = ~P3_ADDR_REG_5_ | ~new_P3_U4760;
  assign new_P3_U4923 = ~new_P3_R1212_U54 | ~new_P3_U3040;
  assign new_P3_U4924 = ~new_P3_U3039 | ~new_P3_U3400;
  assign new_P3_U4925 = ~new_P3_R1209_U54 | ~new_P3_U3037;
  assign new_P3_U4926 = ~new_P3_U4925 | ~new_P3_U4924 | ~new_P3_U4923;
  assign new_P3_U4927 = ~new_P3_R1054_U75 | ~new_P3_U3051;
  assign new_P3_U4928 = ~new_P3_U5768 | ~new_P3_U3400;
  assign new_P3_U4929 = ~new_P3_U3042 | ~new_P3_U4926;
  assign new_P3_U4930 = ~new_P3_R1212_U54 | ~new_P3_U3041;
  assign new_P3_U4931 = ~P3_REG3_REG_4_ | ~n3834;
  assign new_P3_U4932 = ~new_P3_R1209_U54 | ~new_P3_U3038;
  assign new_P3_U4933 = ~P3_ADDR_REG_4_ | ~new_P3_U4760;
  assign new_P3_U4934 = ~new_P3_R1212_U55 | ~new_P3_U3040;
  assign new_P3_U4935 = ~new_P3_U3039 | ~new_P3_U3397;
  assign new_P3_U4936 = ~new_P3_R1209_U55 | ~new_P3_U3037;
  assign new_P3_U4937 = ~new_P3_U4936 | ~new_P3_U4935 | ~new_P3_U4934;
  assign new_P3_U4938 = ~new_P3_R1054_U14 | ~new_P3_U3051;
  assign new_P3_U4939 = ~new_P3_U5768 | ~new_P3_U3397;
  assign new_P3_U4940 = ~new_P3_U3042 | ~new_P3_U4937;
  assign new_P3_U4941 = ~new_P3_R1212_U55 | ~new_P3_U3041;
  assign new_P3_U4942 = ~P3_REG3_REG_3_ | ~n3834;
  assign new_P3_U4943 = ~new_P3_R1209_U55 | ~new_P3_U3038;
  assign new_P3_U4944 = ~P3_ADDR_REG_3_ | ~new_P3_U4760;
  assign new_P3_U4945 = ~new_P3_R1212_U56 | ~new_P3_U3040;
  assign new_P3_U4946 = ~new_P3_U3039 | ~new_P3_U3394;
  assign new_P3_U4947 = ~new_P3_R1209_U56 | ~new_P3_U3037;
  assign new_P3_U4948 = ~new_P3_U4947 | ~new_P3_U4946 | ~new_P3_U4945;
  assign new_P3_U4949 = ~new_P3_R1054_U76 | ~new_P3_U3051;
  assign new_P3_U4950 = ~new_P3_U5768 | ~new_P3_U3394;
  assign new_P3_U4951 = ~new_P3_U3042 | ~new_P3_U4948;
  assign new_P3_U4952 = ~new_P3_R1212_U56 | ~new_P3_U3041;
  assign new_P3_U4953 = ~P3_REG3_REG_2_ | ~n3834;
  assign new_P3_U4954 = ~new_P3_R1209_U56 | ~new_P3_U3038;
  assign new_P3_U4955 = ~P3_ADDR_REG_2_ | ~new_P3_U4760;
  assign new_P3_U4956 = ~new_P3_R1212_U57 | ~new_P3_U3040;
  assign new_P3_U4957 = ~new_P3_U3039 | ~new_P3_U3391;
  assign new_P3_U4958 = ~new_P3_R1209_U57 | ~new_P3_U3037;
  assign new_P3_U4959 = ~new_P3_U4958 | ~new_P3_U4957 | ~new_P3_U4956;
  assign new_P3_U4960 = ~new_P3_R1054_U66 | ~new_P3_U3051;
  assign new_P3_U4961 = ~new_P3_U5768 | ~new_P3_U3391;
  assign new_P3_U4962 = ~new_P3_U3042 | ~new_P3_U4959;
  assign new_P3_U4963 = ~new_P3_R1212_U57 | ~new_P3_U3041;
  assign new_P3_U4964 = ~P3_REG3_REG_1_ | ~n3834;
  assign new_P3_U4965 = ~new_P3_R1209_U57 | ~new_P3_U3038;
  assign new_P3_U4966 = ~P3_ADDR_REG_1_ | ~new_P3_U4760;
  assign new_P3_U4967 = ~new_P3_R1212_U7 | ~new_P3_U3040;
  assign new_P3_U4968 = ~new_P3_U3039 | ~new_P3_U3386;
  assign new_P3_U4969 = ~new_P3_R1209_U7 | ~new_P3_U3037;
  assign new_P3_U4970 = ~new_P3_U4969 | ~new_P3_U4968 | ~new_P3_U4967;
  assign new_P3_U4971 = ~new_P3_R1054_U17 | ~new_P3_U3051;
  assign new_P3_U4972 = ~new_P3_U5768 | ~new_P3_U3386;
  assign new_P3_U4973 = ~new_P3_U3042 | ~new_P3_U4970;
  assign new_P3_U4974 = ~new_P3_R1212_U7 | ~new_P3_U3041;
  assign new_P3_U4975 = ~P3_REG3_REG_0_ | ~n3834;
  assign new_P3_U4976 = ~new_P3_R1209_U7 | ~new_P3_U3038;
  assign new_P3_U4977 = ~P3_ADDR_REG_0_ | ~new_P3_U4760;
  assign new_P3_U4978 = ~new_P3_U3868;
  assign new_P3_U4979 = ~new_P3_U3050 | ~new_P3_U5942 | ~new_P3_U5941;
  assign new_P3_U4980 = ~new_P3_U3867 | ~new_P3_U3023 | ~new_P3_U3909;
  assign new_P3_U4981 = ~P3_B_REG | ~new_P3_U4979;
  assign new_P3_U4982 = ~new_P3_U3036 | ~new_P3_U3078;
  assign new_P3_U4983 = ~new_P3_U3032 | ~new_P3_U3072;
  assign new_P3_U4984 = ~new_P3_SUB_609_U21 | ~new_P3_U3304;
  assign new_P3_U4985 = ~new_P3_U4984 | ~new_P3_U4983 | ~new_P3_U4982;
  assign new_P3_U4986 = ~new_P3_U3312 | ~new_P3_U5425 | ~new_P3_U3888 | ~new_P3_U3311 | ~new_P3_U3875;
  assign new_P3_U4987 = ~new_P3_U3894 | ~new_P3_U4986;
  assign new_P3_U4988 = ~new_P3_U3889 | ~new_P3_U3895;
  assign new_P3_U4989 = ~new_P3_U4988 | ~new_P3_U4987;
  assign new_P3_U4990 = ~new_P3_U3911 | ~new_P3_U3378;
  assign new_P3_U4991 = ~new_P3_U3889 | ~new_P3_U3304;
  assign new_P3_U4992 = ~new_P3_U4986 | ~new_P3_U3303;
  assign new_P3_U4993 = ~new_P3_U3370;
  assign new_P3_U4994 = ~new_P3_U3434 | ~new_P3_U5420;
  assign new_P3_U4995 = ~new_P3_SUB_609_U21 | ~new_P3_U3371;
  assign new_P3_U4996 = ~new_P3_R1158_U114 | ~new_P3_U3035;
  assign new_P3_U4997 = ~new_P3_U3031 | ~new_P3_U4985;
  assign new_P3_U4998 = ~P3_REG3_REG_15_ | ~n3834;
  assign new_P3_U4999 = ~new_P3_U3036 | ~new_P3_U3057;
  assign new_P3_U5000 = ~new_P3_U3032 | ~new_P3_U3052;
  assign new_P3_U5001 = ~new_P3_SUB_609_U26 | ~new_P3_U3304;
  assign new_P3_U5002 = ~new_P3_U5001 | ~new_P3_U5000 | ~new_P3_U4999;
  assign new_P3_U5003 = ~new_P3_U3365 | ~new_P3_U3303;
  assign new_P3_U5004 = ~new_P3_U4993 | ~new_P3_U5003;
  assign new_P3_U5005 = ~new_P3_U3894 | ~new_P3_U3365;
  assign new_P3_U5006 = ~new_P3_U3360 | ~new_P3_U5005;
  assign new_P3_U5007 = ~new_P3_U3045 | ~new_P3_U3901;
  assign new_P3_U5008 = ~new_P3_U3044 | ~new_P3_SUB_609_U26;
  assign new_P3_U5009 = ~new_P3_R1158_U16 | ~new_P3_U3035;
  assign new_P3_U5010 = ~new_P3_U3031 | ~new_P3_U5002;
  assign new_P3_U5011 = ~P3_REG3_REG_26_ | ~n3834;
  assign new_P3_U5012 = ~new_P3_U3036 | ~new_P3_U3066;
  assign new_P3_U5013 = ~new_P3_U3032 | ~new_P3_U3069;
  assign new_P3_U5014 = ~new_P3_SUB_609_U8 | ~new_P3_U3304;
  assign new_P3_U5015 = ~new_P3_U5014 | ~new_P3_U5013 | ~new_P3_U5012;
  assign new_P3_U5016 = ~new_P3_U3407 | ~new_P3_U5420;
  assign new_P3_U5017 = ~new_P3_SUB_609_U8 | ~new_P3_U3371;
  assign new_P3_U5018 = ~new_P3_R1158_U97 | ~new_P3_U3035;
  assign new_P3_U5019 = ~new_P3_U3031 | ~new_P3_U5015;
  assign new_P3_U5020 = ~P3_REG3_REG_6_ | ~n3834;
  assign new_P3_U5021 = ~new_P3_U3036 | ~new_P3_U3068;
  assign new_P3_U5022 = ~new_P3_U3032 | ~new_P3_U3080;
  assign new_P3_U5023 = ~new_P3_SUB_609_U11 | ~new_P3_U3304;
  assign new_P3_U5024 = ~new_P3_U5023 | ~new_P3_U5022 | ~new_P3_U5021;
  assign new_P3_U5025 = ~new_P3_U3443 | ~new_P3_U5420;
  assign new_P3_U5026 = ~new_P3_SUB_609_U11 | ~new_P3_U3371;
  assign new_P3_U5027 = ~new_P3_R1158_U112 | ~new_P3_U3035;
  assign new_P3_U5028 = ~new_P3_U3031 | ~new_P3_U5024;
  assign new_P3_U5029 = ~P3_REG3_REG_18_ | ~n3834;
  assign new_P3_U5030 = ~new_P3_U3036 | ~new_P3_U3077;
  assign new_P3_U5031 = ~new_P3_U3032 | ~new_P3_U3063;
  assign new_P3_U5032 = ~P3_REG3_REG_2_ | ~new_P3_U3304;
  assign new_P3_U5033 = ~new_P3_U5032 | ~new_P3_U5031 | ~new_P3_U5030;
  assign new_P3_U5034 = ~new_P3_U3395 | ~new_P3_U5420;
  assign new_P3_U5035 = ~P3_REG3_REG_2_ | ~new_P3_U3371;
  assign new_P3_U5036 = ~new_P3_R1158_U100 | ~new_P3_U3035;
  assign new_P3_U5037 = ~new_P3_U3031 | ~new_P3_U5033;
  assign new_P3_U5038 = ~P3_REG3_REG_2_ | ~n3834;
  assign new_P3_U5039 = ~new_P3_U3036 | ~new_P3_U3061;
  assign new_P3_U5040 = ~new_P3_U3032 | ~new_P3_U3071;
  assign new_P3_U5041 = ~new_P3_SUB_609_U9 | ~new_P3_U3304;
  assign new_P3_U5042 = ~new_P3_U5041 | ~new_P3_U5040 | ~new_P3_U5039;
  assign new_P3_U5043 = ~new_P3_U3422 | ~new_P3_U5420;
  assign new_P3_U5044 = ~new_P3_SUB_609_U9 | ~new_P3_U3371;
  assign new_P3_U5045 = ~new_P3_R1158_U117 | ~new_P3_U3035;
  assign new_P3_U5046 = ~new_P3_U3031 | ~new_P3_U5042;
  assign new_P3_U5047 = ~P3_REG3_REG_11_ | ~n3834;
  assign new_P3_U5048 = ~new_P3_U3036 | ~new_P3_U3074;
  assign new_P3_U5049 = ~new_P3_U3032 | ~new_P3_U3065;
  assign new_P3_U5050 = ~new_P3_SUB_609_U17 | ~new_P3_U3304;
  assign new_P3_U5051 = ~new_P3_U5050 | ~new_P3_U5049 | ~new_P3_U5048;
  assign new_P3_U5052 = ~new_P3_U3045 | ~new_P3_U3905;
  assign new_P3_U5053 = ~new_P3_U3044 | ~new_P3_SUB_609_U17;
  assign new_P3_U5054 = ~new_P3_R1158_U108 | ~new_P3_U3035;
  assign new_P3_U5055 = ~new_P3_U3031 | ~new_P3_U5051;
  assign new_P3_U5056 = ~P3_REG3_REG_22_ | ~n3834;
  assign new_P3_U5057 = ~new_P3_U3036 | ~new_P3_U3071;
  assign new_P3_U5058 = ~new_P3_U3032 | ~new_P3_U3078;
  assign new_P3_U5059 = ~new_P3_SUB_609_U24 | ~new_P3_U3304;
  assign new_P3_U5060 = ~new_P3_U5059 | ~new_P3_U5058 | ~new_P3_U5057;
  assign new_P3_U5061 = ~new_P3_U3428 | ~new_P3_U5420;
  assign new_P3_U5062 = ~new_P3_SUB_609_U24 | ~new_P3_U3371;
  assign new_P3_U5063 = ~new_P3_R1158_U13 | ~new_P3_U3035;
  assign new_P3_U5064 = ~new_P3_U3031 | ~new_P3_U5060;
  assign new_P3_U5065 = ~P3_REG3_REG_13_ | ~n3834;
  assign new_P3_U5066 = ~new_P3_U3036 | ~new_P3_U3080;
  assign new_P3_U5067 = ~new_P3_U3032 | ~new_P3_U3074;
  assign new_P3_U5068 = ~new_P3_SUB_609_U20 | ~new_P3_U3304;
  assign new_P3_U5069 = ~new_P3_U5068 | ~new_P3_U5067 | ~new_P3_U5066;
  assign new_P3_U5070 = ~new_P3_U3045 | ~new_P3_U3907;
  assign new_P3_U5071 = ~new_P3_U3044 | ~new_P3_SUB_609_U20;
  assign new_P3_U5072 = ~new_P3_R1158_U109 | ~new_P3_U3035;
  assign new_P3_U5073 = ~new_P3_U3031 | ~new_P3_U5069;
  assign new_P3_U5074 = ~P3_REG3_REG_20_ | ~n3834;
  assign new_P3_U5075 = ~new_P3_U3031 | ~new_P3_U3304;
  assign new_P3_U5076 = ~new_P3_U5419 | ~new_P3_U5075;
  assign new_P3_U5077 = ~new_P3_U3787 | ~new_P3_U3032;
  assign new_P3_U5078 = ~new_P3_U3387 | ~new_P3_U5420;
  assign new_P3_U5079 = ~P3_REG3_REG_0_ | ~new_P3_U5076;
  assign new_P3_U5080 = ~new_P3_R1158_U94 | ~new_P3_U3035;
  assign new_P3_U5081 = ~P3_REG3_REG_0_ | ~n3834;
  assign new_P3_U5082 = ~new_P3_U3036 | ~new_P3_U3083;
  assign new_P3_U5083 = ~new_P3_U3032 | ~new_P3_U3061;
  assign new_P3_U5084 = ~new_P3_SUB_609_U14 | ~new_P3_U3304;
  assign new_P3_U5085 = ~new_P3_U5084 | ~new_P3_U5083 | ~new_P3_U5082;
  assign new_P3_U5086 = ~new_P3_U3416 | ~new_P3_U5420;
  assign new_P3_U5087 = ~new_P3_SUB_609_U14 | ~new_P3_U3371;
  assign new_P3_U5088 = ~new_P3_R1158_U95 | ~new_P3_U3035;
  assign new_P3_U5089 = ~new_P3_U3031 | ~new_P3_U5085;
  assign new_P3_U5090 = ~P3_REG3_REG_9_ | ~n3834;
  assign new_P3_U5091 = ~new_P3_U3036 | ~new_P3_U3063;
  assign new_P3_U5092 = ~new_P3_U3032 | ~new_P3_U3066;
  assign new_P3_U5093 = ~new_P3_SUB_609_U29 | ~new_P3_U3304;
  assign new_P3_U5094 = ~new_P3_U5093 | ~new_P3_U5092 | ~new_P3_U5091;
  assign new_P3_U5095 = ~new_P3_U3401 | ~new_P3_U5420;
  assign new_P3_U5096 = ~new_P3_SUB_609_U29 | ~new_P3_U3371;
  assign new_P3_U5097 = ~new_P3_R1158_U99 | ~new_P3_U3035;
  assign new_P3_U5098 = ~new_P3_U3031 | ~new_P3_U5094;
  assign new_P3_U5099 = ~P3_REG3_REG_4_ | ~n3834;
  assign new_P3_U5100 = ~new_P3_U3036 | ~new_P3_U3065;
  assign new_P3_U5101 = ~new_P3_U3032 | ~new_P3_U3057;
  assign new_P3_U5102 = ~new_P3_SUB_609_U10 | ~new_P3_U3304;
  assign new_P3_U5103 = ~new_P3_U5102 | ~new_P3_U5101 | ~new_P3_U5100;
  assign new_P3_U5104 = ~new_P3_U3045 | ~new_P3_U3903;
  assign new_P3_U5105 = ~new_P3_U3044 | ~new_P3_SUB_609_U10;
  assign new_P3_U5106 = ~new_P3_R1158_U106 | ~new_P3_U3035;
  assign new_P3_U5107 = ~new_P3_U3031 | ~new_P3_U5103;
  assign new_P3_U5108 = ~P3_REG3_REG_24_ | ~n3834;
  assign new_P3_U5109 = ~new_P3_U3036 | ~new_P3_U3072;
  assign new_P3_U5110 = ~new_P3_U3032 | ~new_P3_U3081;
  assign new_P3_U5111 = ~new_P3_SUB_609_U19 | ~new_P3_U3304;
  assign new_P3_U5112 = ~new_P3_U5111 | ~new_P3_U5110 | ~new_P3_U5109;
  assign new_P3_U5113 = ~new_P3_U3440 | ~new_P3_U5420;
  assign new_P3_U5114 = ~new_P3_SUB_609_U19 | ~new_P3_U3371;
  assign new_P3_U5115 = ~new_P3_R1158_U14 | ~new_P3_U3035;
  assign new_P3_U5116 = ~new_P3_U3031 | ~new_P3_U5112;
  assign new_P3_U5117 = ~P3_REG3_REG_17_ | ~n3834;
  assign new_P3_U5118 = ~new_P3_U3036 | ~new_P3_U3059;
  assign new_P3_U5119 = ~new_P3_U3032 | ~new_P3_U3070;
  assign new_P3_U5120 = ~new_P3_SUB_609_U53 | ~new_P3_U3304;
  assign new_P3_U5121 = ~new_P3_U5120 | ~new_P3_U5119 | ~new_P3_U5118;
  assign new_P3_U5122 = ~new_P3_U3404 | ~new_P3_U5420;
  assign new_P3_U5123 = ~new_P3_SUB_609_U53 | ~new_P3_U3371;
  assign new_P3_U5124 = ~new_P3_R1158_U98 | ~new_P3_U3035;
  assign new_P3_U5125 = ~new_P3_U3031 | ~new_P3_U5121;
  assign new_P3_U5126 = ~P3_REG3_REG_5_ | ~n3834;
  assign new_P3_U5127 = ~new_P3_U3036 | ~new_P3_U3073;
  assign new_P3_U5128 = ~new_P3_U3032 | ~new_P3_U3068;
  assign new_P3_U5129 = ~new_P3_SUB_609_U7 | ~new_P3_U3304;
  assign new_P3_U5130 = ~new_P3_U5129 | ~new_P3_U5128 | ~new_P3_U5127;
  assign new_P3_U5131 = ~new_P3_U3437 | ~new_P3_U5420;
  assign new_P3_U5132 = ~new_P3_SUB_609_U7 | ~new_P3_U3371;
  assign new_P3_U5133 = ~new_P3_R1158_U113 | ~new_P3_U3035;
  assign new_P3_U5134 = ~new_P3_U3031 | ~new_P3_U5130;
  assign new_P3_U5135 = ~P3_REG3_REG_16_ | ~n3834;
  assign new_P3_U5136 = ~new_P3_U3036 | ~new_P3_U3064;
  assign new_P3_U5137 = ~new_P3_U3032 | ~new_P3_U3056;
  assign new_P3_U5138 = ~new_P3_SUB_609_U16 | ~new_P3_U3304;
  assign new_P3_U5139 = ~new_P3_U5138 | ~new_P3_U5137 | ~new_P3_U5136;
  assign new_P3_U5140 = ~new_P3_U3045 | ~new_P3_U3902;
  assign new_P3_U5141 = ~new_P3_U3044 | ~new_P3_SUB_609_U16;
  assign new_P3_U5142 = ~new_P3_R1158_U105 | ~new_P3_U3035;
  assign new_P3_U5143 = ~new_P3_U3031 | ~new_P3_U5139;
  assign new_P3_U5144 = ~P3_REG3_REG_25_ | ~n3834;
  assign new_P3_U5145 = ~new_P3_U3036 | ~new_P3_U3062;
  assign new_P3_U5146 = ~new_P3_U3032 | ~new_P3_U3079;
  assign new_P3_U5147 = ~new_P3_SUB_609_U23 | ~new_P3_U3304;
  assign new_P3_U5148 = ~new_P3_U5147 | ~new_P3_U5146 | ~new_P3_U5145;
  assign new_P3_U5149 = ~new_P3_U3425 | ~new_P3_U5420;
  assign new_P3_U5150 = ~new_P3_SUB_609_U23 | ~new_P3_U3371;
  assign new_P3_U5151 = ~new_P3_R1158_U116 | ~new_P3_U3035;
  assign new_P3_U5152 = ~new_P3_U3031 | ~new_P3_U5148;
  assign new_P3_U5153 = ~P3_REG3_REG_12_ | ~n3834;
  assign new_P3_U5154 = ~new_P3_U3036 | ~new_P3_U3075;
  assign new_P3_U5155 = ~new_P3_U3032 | ~new_P3_U3060;
  assign new_P3_U5156 = ~new_P3_SUB_609_U27 | ~new_P3_U3304;
  assign new_P3_U5157 = ~new_P3_U5156 | ~new_P3_U5155 | ~new_P3_U5154;
  assign new_P3_U5158 = ~new_P3_U3045 | ~new_P3_U3906;
  assign new_P3_U5159 = ~new_P3_U3044 | ~new_P3_SUB_609_U27;
  assign new_P3_U5160 = ~new_P3_R1158_U15 | ~new_P3_U3035;
  assign new_P3_U5161 = ~new_P3_U3031 | ~new_P3_U5157;
  assign new_P3_U5162 = ~P3_REG3_REG_21_ | ~n3834;
  assign new_P3_U5163 = ~new_P3_U3036 | ~new_P3_U3076;
  assign new_P3_U5164 = ~new_P3_U3032 | ~new_P3_U3067;
  assign new_P3_U5165 = ~P3_REG3_REG_1_ | ~new_P3_U3304;
  assign new_P3_U5166 = ~new_P3_U5165 | ~new_P3_U5164 | ~new_P3_U5163;
  assign new_P3_U5167 = ~new_P3_U3392 | ~new_P3_U5420;
  assign new_P3_U5168 = ~P3_REG3_REG_1_ | ~new_P3_U3371;
  assign new_P3_U5169 = ~new_P3_R1158_U110 | ~new_P3_U3035;
  assign new_P3_U5170 = ~new_P3_U3031 | ~new_P3_U5166;
  assign new_P3_U5171 = ~P3_REG3_REG_1_ | ~n3834;
  assign new_P3_U5172 = ~new_P3_U3036 | ~new_P3_U3069;
  assign new_P3_U5173 = ~new_P3_U3032 | ~new_P3_U3082;
  assign new_P3_U5174 = ~new_P3_SUB_609_U12 | ~new_P3_U3304;
  assign new_P3_U5175 = ~new_P3_U5174 | ~new_P3_U5173 | ~new_P3_U5172;
  assign new_P3_U5176 = ~new_P3_U3413 | ~new_P3_U5420;
  assign new_P3_U5177 = ~new_P3_SUB_609_U12 | ~new_P3_U3371;
  assign new_P3_U5178 = ~new_P3_R1158_U96 | ~new_P3_U3035;
  assign new_P3_U5179 = ~new_P3_U3031 | ~new_P3_U5175;
  assign new_P3_U5180 = ~P3_REG3_REG_8_ | ~n3834;
  assign new_P3_U5181 = ~new_P3_U3036 | ~new_P3_U3052;
  assign new_P3_U5182 = ~new_P3_U3032 | ~new_P3_U3054;
  assign new_P3_U5183 = ~new_P3_SUB_609_U28 | ~new_P3_U3304;
  assign new_P3_U5184 = ~new_P3_U5183 | ~new_P3_U5182 | ~new_P3_U5181;
  assign new_P3_U5185 = ~new_P3_U3045 | ~new_P3_U3899;
  assign new_P3_U5186 = ~new_P3_U3044 | ~new_P3_SUB_609_U28;
  assign new_P3_U5187 = ~new_P3_R1158_U101 | ~new_P3_U3035;
  assign new_P3_U5188 = ~new_P3_U3031 | ~new_P3_U5184;
  assign new_P3_U5189 = ~P3_REG3_REG_28_ | ~n3834;
  assign new_P3_U5190 = ~new_P3_U3036 | ~new_P3_U3081;
  assign new_P3_U5191 = ~new_P3_U3032 | ~new_P3_U3075;
  assign new_P3_U5192 = ~new_P3_SUB_609_U15 | ~new_P3_U3304;
  assign new_P3_U5193 = ~new_P3_U5192 | ~new_P3_U5191 | ~new_P3_U5190;
  assign new_P3_U5194 = ~new_P3_U3445 | ~new_P3_U5420;
  assign new_P3_U5195 = ~new_P3_SUB_609_U15 | ~new_P3_U3371;
  assign new_P3_U5196 = ~new_P3_R1158_U111 | ~new_P3_U3035;
  assign new_P3_U5197 = ~new_P3_U3031 | ~new_P3_U5193;
  assign new_P3_U5198 = ~P3_REG3_REG_19_ | ~n3834;
  assign new_P3_U5199 = ~new_P3_U3036 | ~new_P3_U3067;
  assign new_P3_U5200 = ~new_P3_U3032 | ~new_P3_U3059;
  assign new_P3_U5201 = ~new_P3_SUB_609_U25 | ~new_P3_U3304;
  assign new_P3_U5202 = ~new_P3_U5201 | ~new_P3_U5200 | ~new_P3_U5199;
  assign new_P3_U5203 = ~new_P3_U3398 | ~new_P3_U5420;
  assign new_P3_U5204 = ~new_P3_SUB_609_U25 | ~new_P3_U3371;
  assign new_P3_U5205 = ~new_P3_R1158_U17 | ~new_P3_U3035;
  assign new_P3_U5206 = ~new_P3_U3031 | ~new_P3_U5202;
  assign new_P3_U5207 = ~P3_REG3_REG_3_ | ~n3834;
  assign new_P3_U5208 = ~new_P3_U3036 | ~new_P3_U3082;
  assign new_P3_U5209 = ~new_P3_U3032 | ~new_P3_U3062;
  assign new_P3_U5210 = ~new_P3_SUB_609_U13 | ~new_P3_U3304;
  assign new_P3_U5211 = ~new_P3_U5210 | ~new_P3_U5209 | ~new_P3_U5208;
  assign new_P3_U5212 = ~new_P3_U3419 | ~new_P3_U5420;
  assign new_P3_U5213 = ~new_P3_SUB_609_U13 | ~new_P3_U3371;
  assign new_P3_U5214 = ~new_P3_R1158_U118 | ~new_P3_U3035;
  assign new_P3_U5215 = ~new_P3_U3031 | ~new_P3_U5211;
  assign new_P3_U5216 = ~P3_REG3_REG_10_ | ~n3834;
  assign new_P3_U5217 = ~new_P3_U3036 | ~new_P3_U3060;
  assign new_P3_U5218 = ~new_P3_U3032 | ~new_P3_U3064;
  assign new_P3_U5219 = ~new_P3_SUB_609_U6 | ~new_P3_U3304;
  assign new_P3_U5220 = ~new_P3_U5219 | ~new_P3_U5218 | ~new_P3_U5217;
  assign new_P3_U5221 = ~new_P3_U3045 | ~new_P3_U3904;
  assign new_P3_U5222 = ~new_P3_U3044 | ~new_P3_SUB_609_U6;
  assign new_P3_U5223 = ~new_P3_R1158_U107 | ~new_P3_U3035;
  assign new_P3_U5224 = ~new_P3_U3031 | ~new_P3_U5220;
  assign new_P3_U5225 = ~P3_REG3_REG_23_ | ~n3834;
  assign new_P3_U5226 = ~new_P3_U3036 | ~new_P3_U3079;
  assign new_P3_U5227 = ~new_P3_U3032 | ~new_P3_U3073;
  assign new_P3_U5228 = ~new_P3_SUB_609_U30 | ~new_P3_U3304;
  assign new_P3_U5229 = ~new_P3_U5228 | ~new_P3_U5227 | ~new_P3_U5226;
  assign new_P3_U5230 = ~new_P3_U3431 | ~new_P3_U5420;
  assign new_P3_U5231 = ~new_P3_SUB_609_U30 | ~new_P3_U3371;
  assign new_P3_U5232 = ~new_P3_R1158_U115 | ~new_P3_U3035;
  assign new_P3_U5233 = ~new_P3_U3031 | ~new_P3_U5229;
  assign new_P3_U5234 = ~P3_REG3_REG_14_ | ~n3834;
  assign new_P3_U5235 = ~new_P3_U3036 | ~new_P3_U3056;
  assign new_P3_U5236 = ~new_P3_U3032 | ~new_P3_U3053;
  assign new_P3_U5237 = ~new_P3_SUB_609_U22 | ~new_P3_U3304;
  assign new_P3_U5238 = ~new_P3_U5237 | ~new_P3_U5236 | ~new_P3_U5235;
  assign new_P3_U5239 = ~new_P3_U3045 | ~new_P3_U3900;
  assign new_P3_U5240 = ~new_P3_U3044 | ~new_P3_SUB_609_U22;
  assign new_P3_U5241 = ~new_P3_R1158_U102 | ~new_P3_U3035;
  assign new_P3_U5242 = ~new_P3_U3031 | ~new_P3_U5238;
  assign new_P3_U5243 = ~P3_REG3_REG_27_ | ~n3834;
  assign new_P3_U5244 = ~new_P3_U3036 | ~new_P3_U3070;
  assign new_P3_U5245 = ~new_P3_U3032 | ~new_P3_U3083;
  assign new_P3_U5246 = ~new_P3_SUB_609_U18 | ~new_P3_U3304;
  assign new_P3_U5247 = ~new_P3_U5246 | ~new_P3_U5245 | ~new_P3_U5244;
  assign new_P3_U5248 = ~new_P3_U3410 | ~new_P3_U5420;
  assign new_P3_U5249 = ~new_P3_SUB_609_U18 | ~new_P3_U3371;
  assign new_P3_U5250 = ~new_P3_R1158_U18 | ~new_P3_U3035;
  assign new_P3_U5251 = ~new_P3_U3031 | ~new_P3_U5247;
  assign new_P3_U5252 = ~P3_REG3_REG_7_ | ~n3834;
  assign new_P3_U5253 = ~new_P3_U3898 | ~new_P3_U3046;
  assign new_P3_U5254 = ~new_P3_U3375 | ~new_P3_U3833;
  assign new_P3_U5255 = ~new_P3_U3816 | ~new_P3_U3815;
  assign new_P3_U5256 = ~new_P3_U3814 | ~new_P3_U3013;
  assign new_P3_U5257 = ~new_P3_U3880 | ~new_P3_U5256;
  assign new_P3_U5258 = ~new_P3_U3416 | ~new_P3_U5257;
  assign new_P3_U5259 = ~new_P3_U5255 | ~new_P3_U3082;
  assign new_P3_U5260 = ~new_P3_U3413 | ~new_P3_U5257;
  assign new_P3_U5261 = ~new_P3_U5255 | ~new_P3_U3083;
  assign new_P3_U5262 = ~new_P3_U3410 | ~new_P3_U5257;
  assign new_P3_U5263 = ~new_P3_U5255 | ~new_P3_U3069;
  assign new_P3_U5264 = ~new_P3_U3407 | ~new_P3_U5257;
  assign new_P3_U5265 = ~new_P3_U5255 | ~new_P3_U3070;
  assign new_P3_U5266 = ~new_P3_U3404 | ~new_P3_U5257;
  assign new_P3_U5267 = ~new_P3_U5255 | ~new_P3_U3066;
  assign new_P3_U5268 = ~new_P3_U3401 | ~new_P3_U5257;
  assign new_P3_U5269 = ~new_P3_U5255 | ~new_P3_U3059;
  assign new_P3_U5270 = ~new_P3_U3872 | ~new_P3_U5257;
  assign new_P3_U5271 = ~new_P3_U5255 | ~new_P3_U3055;
  assign new_P3_U5272 = ~new_P3_U3873 | ~new_P3_U5257;
  assign new_P3_U5273 = ~new_P3_U5255 | ~new_P3_U3058;
  assign new_P3_U5274 = ~new_P3_U3398 | ~new_P3_U5257;
  assign new_P3_U5275 = ~new_P3_U5255 | ~new_P3_U3063;
  assign new_P3_U5276 = ~new_P3_U3908 | ~new_P3_U5257;
  assign new_P3_U5277 = ~new_P3_U5255 | ~new_P3_U3054;
  assign new_P3_U5278 = ~new_P3_U3899 | ~new_P3_U5257;
  assign new_P3_U5279 = ~new_P3_U5255 | ~new_P3_U3053;
  assign new_P3_U5280 = ~new_P3_U3900 | ~new_P3_U5257;
  assign new_P3_U5281 = ~new_P3_U5255 | ~new_P3_U3052;
  assign new_P3_U5282 = ~new_P3_U3901 | ~new_P3_U5257;
  assign new_P3_U5283 = ~new_P3_U5255 | ~new_P3_U3056;
  assign new_P3_U5284 = ~new_P3_U3902 | ~new_P3_U5257;
  assign new_P3_U5285 = ~new_P3_U5255 | ~new_P3_U3057;
  assign new_P3_U5286 = ~new_P3_U3903 | ~new_P3_U5257;
  assign new_P3_U5287 = ~new_P3_U5255 | ~new_P3_U3064;
  assign new_P3_U5288 = ~new_P3_U3904 | ~new_P3_U5257;
  assign new_P3_U5289 = ~new_P3_U5255 | ~new_P3_U3065;
  assign new_P3_U5290 = ~new_P3_U3905 | ~new_P3_U5257;
  assign new_P3_U5291 = ~new_P3_U5255 | ~new_P3_U3060;
  assign new_P3_U5292 = ~new_P3_U3906 | ~new_P3_U5257;
  assign new_P3_U5293 = ~new_P3_U5255 | ~new_P3_U3074;
  assign new_P3_U5294 = ~new_P3_U3907 | ~new_P3_U5257;
  assign new_P3_U5295 = ~new_P3_U5255 | ~new_P3_U3075;
  assign new_P3_U5296 = ~new_P3_U3395 | ~new_P3_U5257;
  assign new_P3_U5297 = ~new_P3_U5255 | ~new_P3_U3067;
  assign new_P3_U5298 = ~new_P3_U3445 | ~new_P3_U5257;
  assign new_P3_U5299 = ~new_P3_U5255 | ~new_P3_U3080;
  assign new_P3_U5300 = ~new_P3_U3443 | ~new_P3_U5257;
  assign new_P3_U5301 = ~new_P3_U5255 | ~new_P3_U3081;
  assign new_P3_U5302 = ~new_P3_U3440 | ~new_P3_U5257;
  assign new_P3_U5303 = ~new_P3_U5255 | ~new_P3_U3068;
  assign new_P3_U5304 = ~new_P3_U3437 | ~new_P3_U5257;
  assign new_P3_U5305 = ~new_P3_U5255 | ~new_P3_U3072;
  assign new_P3_U5306 = ~new_P3_U3434 | ~new_P3_U5257;
  assign new_P3_U5307 = ~new_P3_U5255 | ~new_P3_U3073;
  assign new_P3_U5308 = ~new_P3_U3431 | ~new_P3_U5257;
  assign new_P3_U5309 = ~new_P3_U5255 | ~new_P3_U3078;
  assign new_P3_U5310 = ~new_P3_U3428 | ~new_P3_U5257;
  assign new_P3_U5311 = ~new_P3_U5255 | ~new_P3_U3079;
  assign new_P3_U5312 = ~new_P3_U3425 | ~new_P3_U5257;
  assign new_P3_U5313 = ~new_P3_U5255 | ~new_P3_U3071;
  assign new_P3_U5314 = ~new_P3_U3422 | ~new_P3_U5257;
  assign new_P3_U5315 = ~new_P3_U5255 | ~new_P3_U3062;
  assign new_P3_U5316 = ~new_P3_U3419 | ~new_P3_U5257;
  assign new_P3_U5317 = ~new_P3_U5255 | ~new_P3_U3061;
  assign new_P3_U5318 = ~new_P3_U3392 | ~new_P3_U5257;
  assign new_P3_U5319 = ~new_P3_U5255 | ~new_P3_U3077;
  assign new_P3_U5320 = ~new_P3_U3387 | ~new_P3_U5257;
  assign new_P3_U5321 = ~new_P3_U5255 | ~new_P3_U3076;
  assign new_P3_U5322 = ~new_P3_U3416 | ~new_P3_U5255;
  assign new_P3_U5323 = ~new_P3_U5257 | ~new_P3_U3082;
  assign new_P3_U5324 = ~new_P3_U5440 | ~new_P3_U3083;
  assign new_P3_U5325 = ~new_P3_U3413 | ~new_P3_U5255;
  assign new_P3_U5326 = ~new_P3_U5257 | ~new_P3_U3083;
  assign new_P3_U5327 = ~new_P3_U5440 | ~new_P3_U3069;
  assign new_P3_U5328 = ~new_P3_U3410 | ~new_P3_U5255;
  assign new_P3_U5329 = ~new_P3_U5257 | ~new_P3_U3069;
  assign new_P3_U5330 = ~new_P3_U5440 | ~new_P3_U3070;
  assign new_P3_U5331 = ~new_P3_U3407 | ~new_P3_U5255;
  assign new_P3_U5332 = ~new_P3_U5257 | ~new_P3_U3070;
  assign new_P3_U5333 = ~new_P3_U5440 | ~new_P3_U3066;
  assign new_P3_U5334 = ~new_P3_U3404 | ~new_P3_U5255;
  assign new_P3_U5335 = ~new_P3_U5257 | ~new_P3_U3066;
  assign new_P3_U5336 = ~new_P3_U5440 | ~new_P3_U3059;
  assign new_P3_U5337 = ~new_P3_U3401 | ~new_P3_U5255;
  assign new_P3_U5338 = ~new_P3_U5257 | ~new_P3_U3059;
  assign new_P3_U5339 = ~new_P3_U5440 | ~new_P3_U3063;
  assign new_P3_U5340 = ~new_P3_U5257 | ~new_P3_U3055;
  assign new_P3_U5341 = ~new_P3_U3872 | ~new_P3_U5255;
  assign new_P3_U5342 = ~new_P3_U5257 | ~new_P3_U3058;
  assign new_P3_U5343 = ~new_P3_U3873 | ~new_P3_U5255;
  assign new_P3_U5344 = ~new_P3_U3398 | ~new_P3_U5255;
  assign new_P3_U5345 = ~new_P3_U5257 | ~new_P3_U3063;
  assign new_P3_U5346 = ~new_P3_U5440 | ~new_P3_U3067;
  assign new_P3_U5347 = ~new_P3_U5257 | ~new_P3_U3054;
  assign new_P3_U5348 = ~new_P3_U3908 | ~new_P3_U5255;
  assign new_P3_U5349 = ~new_P3_U5440 | ~new_P3_U3053;
  assign new_P3_U5350 = ~new_P3_U5257 | ~new_P3_U3053;
  assign new_P3_U5351 = ~new_P3_U3899 | ~new_P3_U5255;
  assign new_P3_U5352 = ~new_P3_U5440 | ~new_P3_U3052;
  assign new_P3_U5353 = ~new_P3_U5257 | ~new_P3_U3052;
  assign new_P3_U5354 = ~new_P3_U3900 | ~new_P3_U5255;
  assign new_P3_U5355 = ~new_P3_U5440 | ~new_P3_U3056;
  assign new_P3_U5356 = ~new_P3_U5257 | ~new_P3_U3056;
  assign new_P3_U5357 = ~new_P3_U3901 | ~new_P3_U5255;
  assign new_P3_U5358 = ~new_P3_U5440 | ~new_P3_U3057;
  assign new_P3_U5359 = ~new_P3_U5257 | ~new_P3_U3057;
  assign new_P3_U5360 = ~new_P3_U3902 | ~new_P3_U5255;
  assign new_P3_U5361 = ~new_P3_U5440 | ~new_P3_U3064;
  assign new_P3_U5362 = ~new_P3_U5257 | ~new_P3_U3064;
  assign new_P3_U5363 = ~new_P3_U3903 | ~new_P3_U5255;
  assign new_P3_U5364 = ~new_P3_U5440 | ~new_P3_U3065;
  assign new_P3_U5365 = ~new_P3_U5257 | ~new_P3_U3065;
  assign new_P3_U5366 = ~new_P3_U3904 | ~new_P3_U5255;
  assign new_P3_U5367 = ~new_P3_U5440 | ~new_P3_U3060;
  assign new_P3_U5368 = ~new_P3_U5257 | ~new_P3_U3060;
  assign new_P3_U5369 = ~new_P3_U3905 | ~new_P3_U5255;
  assign new_P3_U5370 = ~new_P3_U5440 | ~new_P3_U3074;
  assign new_P3_U5371 = ~new_P3_U5257 | ~new_P3_U3074;
  assign new_P3_U5372 = ~new_P3_U3906 | ~new_P3_U5255;
  assign new_P3_U5373 = ~new_P3_U5440 | ~new_P3_U3075;
  assign new_P3_U5374 = ~new_P3_U5257 | ~new_P3_U3075;
  assign new_P3_U5375 = ~new_P3_U3907 | ~new_P3_U5255;
  assign new_P3_U5376 = ~new_P3_U5440 | ~new_P3_U3080;
  assign new_P3_U5377 = ~new_P3_U3395 | ~new_P3_U5255;
  assign new_P3_U5378 = ~new_P3_U5257 | ~new_P3_U3067;
  assign new_P3_U5379 = ~new_P3_U5440 | ~new_P3_U3077;
  assign new_P3_U5380 = ~new_P3_U3445 | ~new_P3_U5255;
  assign new_P3_U5381 = ~new_P3_U5257 | ~new_P3_U3080;
  assign new_P3_U5382 = ~new_P3_U5440 | ~new_P3_U3081;
  assign new_P3_U5383 = ~new_P3_U3443 | ~new_P3_U5255;
  assign new_P3_U5384 = ~new_P3_U5257 | ~new_P3_U3081;
  assign new_P3_U5385 = ~new_P3_U5440 | ~new_P3_U3068;
  assign new_P3_U5386 = ~new_P3_U3440 | ~new_P3_U5255;
  assign new_P3_U5387 = ~new_P3_U5257 | ~new_P3_U3068;
  assign new_P3_U5388 = ~new_P3_U5440 | ~new_P3_U3072;
  assign new_P3_U5389 = ~new_P3_U3437 | ~new_P3_U5255;
  assign new_P3_U5390 = ~new_P3_U5257 | ~new_P3_U3072;
  assign new_P3_U5391 = ~new_P3_U5440 | ~new_P3_U3073;
  assign new_P3_U5392 = ~new_P3_U3434 | ~new_P3_U5255;
  assign new_P3_U5393 = ~new_P3_U5257 | ~new_P3_U3073;
  assign new_P3_U5394 = ~new_P3_U5440 | ~new_P3_U3078;
  assign new_P3_U5395 = ~new_P3_U3431 | ~new_P3_U5255;
  assign new_P3_U5396 = ~new_P3_U5257 | ~new_P3_U3078;
  assign new_P3_U5397 = ~new_P3_U5440 | ~new_P3_U3079;
  assign new_P3_U5398 = ~new_P3_U3428 | ~new_P3_U5255;
  assign new_P3_U5399 = ~new_P3_U5257 | ~new_P3_U3079;
  assign new_P3_U5400 = ~new_P3_U5440 | ~new_P3_U3071;
  assign new_P3_U5401 = ~new_P3_U3425 | ~new_P3_U5255;
  assign new_P3_U5402 = ~new_P3_U5257 | ~new_P3_U3071;
  assign new_P3_U5403 = ~new_P3_U5440 | ~new_P3_U3062;
  assign new_P3_U5404 = ~new_P3_U3422 | ~new_P3_U5255;
  assign new_P3_U5405 = ~new_P3_U5257 | ~new_P3_U3062;
  assign new_P3_U5406 = ~new_P3_U5440 | ~new_P3_U3061;
  assign new_P3_U5407 = ~new_P3_U3419 | ~new_P3_U5255;
  assign new_P3_U5408 = ~new_P3_U5257 | ~new_P3_U3061;
  assign new_P3_U5409 = ~new_P3_U5440 | ~new_P3_U3082;
  assign new_P3_U5410 = ~new_P3_U3392 | ~new_P3_U5255;
  assign new_P3_U5411 = ~new_P3_U5257 | ~new_P3_U3077;
  assign new_P3_U5412 = ~new_P3_U5440 | ~new_P3_U3076;
  assign new_P3_U5413 = ~new_P3_U3387 | ~new_P3_U5255;
  assign new_P3_U5414 = ~new_P3_U5257 | ~new_P3_U3076;
  assign new_P3_U5415 = ~new_P3_U4981 | ~n3834;
  assign new_P3_U5416 = ~new_P3_U4980 | ~new_P3_U4981 | ~new_P3_U5440;
  assign new_P3_U5417 = ~new_P3_U3043 | ~new_P3_U3303;
  assign new_P3_U5418 = ~new_P3_U3043 | ~new_P3_U3894;
  assign new_P3_U5419 = ~new_P3_U3371;
  assign new_P3_U5420 = ~new_P3_U5418 | ~new_P3_U3918;
  assign new_P3_U5421 = ~new_P3_U3774 | ~new_P3_U5938 | ~new_P3_U5937;
  assign new_P3_U5422 = ~new_P3_U5434 | ~new_P3_U5428;
  assign new_P3_U5423 = ~new_P3_U3879 | ~new_P3_U3378;
  assign new_P3_U5424 = ~new_P3_U3375 | ~new_P3_U3833;
  assign new_P3_U5425 = ~new_P3_U3876 | ~new_P3_U5447;
  assign new_P3_U5426 = ~P3_IR_REG_24_ | ~new_P3_U3831;
  assign new_P3_U5427 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U18;
  assign new_P3_U5428 = ~new_P3_U3372;
  assign new_P3_U5429 = ~P3_IR_REG_25_ | ~new_P3_U3831;
  assign new_P3_U5430 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U81;
  assign new_P3_U5431 = ~new_P3_U3373;
  assign new_P3_U5432 = ~P3_IR_REG_26_ | ~new_P3_U3831;
  assign new_P3_U5433 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U19;
  assign new_P3_U5434 = ~new_P3_U3374;
  assign new_P3_U5435 = ~new_P3_U5428 | ~P3_B_REG;
  assign new_P3_U5436 = ~new_P3_U3372 | ~new_P3_U3298;
  assign new_P3_U5437 = ~new_P3_U5436 | ~new_P3_U5435;
  assign new_P3_U5438 = ~P3_IR_REG_23_ | ~new_P3_U3831;
  assign new_P3_U5439 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U17;
  assign new_P3_U5440 = ~new_P3_U3375;
  assign new_P3_U5441 = ~P3_D_REG_0_ | ~new_P3_U3832;
  assign new_P3_U5442 = ~new_P3_U3915 | ~new_P3_U4020;
  assign new_P3_U5443 = ~P3_D_REG_1_ | ~new_P3_U3832;
  assign new_P3_U5444 = ~new_P3_U3915 | ~new_P3_U4021;
  assign new_P3_U5445 = ~P3_IR_REG_20_ | ~new_P3_U3831;
  assign new_P3_U5446 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U15;
  assign new_P3_U5447 = ~new_P3_U3378;
  assign new_P3_U5448 = ~P3_IR_REG_19_ | ~new_P3_U3831;
  assign new_P3_U5449 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U14;
  assign new_P3_U5450 = ~new_P3_U3379;
  assign new_P3_U5451 = ~P3_IR_REG_22_ | ~new_P3_U3831;
  assign new_P3_U5452 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U16;
  assign new_P3_U5453 = ~new_P3_U3380;
  assign new_P3_U5454 = ~P3_IR_REG_21_ | ~new_P3_U3831;
  assign new_P3_U5455 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U83;
  assign new_P3_U5456 = ~new_P3_U3385;
  assign new_P3_U5457 = ~P3_IR_REG_30_ | ~new_P3_U3831;
  assign new_P3_U5458 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U77;
  assign new_P3_U5459 = ~new_P3_U3381;
  assign new_P3_U5460 = ~P3_IR_REG_29_ | ~new_P3_U3831;
  assign new_P3_U5461 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U21;
  assign new_P3_U5462 = ~new_P3_U3382;
  assign new_P3_U5463 = ~P3_IR_REG_28_ | ~new_P3_U3831;
  assign new_P3_U5464 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U20;
  assign new_P3_U5465 = ~new_P3_U3383;
  assign new_P3_U5466 = ~P3_IR_REG_27_ | ~new_P3_U3831;
  assign new_P3_U5467 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U79;
  assign new_P3_U5468 = ~new_P3_U3384;
  assign new_P3_U5469 = ~P3_IR_REG_0_ | ~new_P3_U3831;
  assign new_P3_U5470 = ~P3_IR_REG_31_ | ~P3_IR_REG_0_;
  assign new_P3_U5471 = ~new_U61 | ~new_P3_U3833;
  assign new_P3_U5472 = ~new_P3_U3893 | ~new_P3_U3386;
  assign new_P3_U5473 = ~new_P3_U3387;
  assign new_P3_U5474 = ~new_P3_U5422 | ~new_P3_U3300;
  assign new_P3_U5475 = ~P3_D_REG_0_ | ~new_P3_U4019;
  assign new_P3_U5476 = ~new_P3_U3388;
  assign new_P3_U5477 = ~P3_D_REG_1_ | ~new_P3_U4019;
  assign new_P3_U5478 = ~new_P3_U4021 | ~new_P3_U3300;
  assign new_P3_U5479 = ~new_P3_U3389;
  assign new_P3_U5480 = ~new_P3_U4052 | ~new_P3_U5453;
  assign new_P3_U5481 = ~new_P3_U3380 | ~new_P3_U3834;
  assign new_P3_U5482 = ~new_P3_U5481 | ~new_P3_U5480;
  assign new_P3_U5483 = ~P3_REG0_REG_0_ | ~new_P3_U3835;
  assign new_P3_U5484 = ~new_P3_U3914 | ~new_P3_U4077;
  assign new_P3_U5485 = ~P3_IR_REG_1_ | ~new_P3_U3831;
  assign new_P3_U5486 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U51;
  assign new_P3_U5487 = ~new_U50 | ~new_P3_U3833;
  assign new_P3_U5488 = ~new_P3_U3391 | ~new_P3_U3893;
  assign new_P3_U5489 = ~new_P3_U3392;
  assign new_P3_U5490 = ~P3_REG0_REG_1_ | ~new_P3_U3835;
  assign new_P3_U5491 = ~new_P3_U3914 | ~new_P3_U4102;
  assign new_P3_U5492 = ~P3_IR_REG_2_ | ~new_P3_U3831;
  assign new_P3_U5493 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U22;
  assign new_P3_U5494 = ~new_U39 | ~new_P3_U3833;
  assign new_P3_U5495 = ~new_P3_U3394 | ~new_P3_U3893;
  assign new_P3_U5496 = ~new_P3_U3395;
  assign new_P3_U5497 = ~P3_REG0_REG_2_ | ~new_P3_U3835;
  assign new_P3_U5498 = ~new_P3_U3914 | ~new_P3_U4120;
  assign new_P3_U5499 = ~P3_IR_REG_3_ | ~new_P3_U3831;
  assign new_P3_U5500 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U23;
  assign new_P3_U5501 = ~new_U36 | ~new_P3_U3833;
  assign new_P3_U5502 = ~new_P3_U3397 | ~new_P3_U3893;
  assign new_P3_U5503 = ~new_P3_U3398;
  assign new_P3_U5504 = ~P3_REG0_REG_3_ | ~new_P3_U3835;
  assign new_P3_U5505 = ~new_P3_U3914 | ~new_P3_U4138;
  assign new_P3_U5506 = ~P3_IR_REG_4_ | ~new_P3_U3831;
  assign new_P3_U5507 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U24;
  assign new_P3_U5508 = ~new_U35 | ~new_P3_U3833;
  assign new_P3_U5509 = ~new_P3_U3400 | ~new_P3_U3893;
  assign new_P3_U5510 = ~new_P3_U3401;
  assign new_P3_U5511 = ~P3_REG0_REG_4_ | ~new_P3_U3835;
  assign new_P3_U5512 = ~new_P3_U3914 | ~new_P3_U4156;
  assign new_P3_U5513 = ~P3_IR_REG_5_ | ~new_P3_U3831;
  assign new_P3_U5514 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U74;
  assign new_P3_U5515 = ~new_U34 | ~new_P3_U3833;
  assign new_P3_U5516 = ~new_P3_U3403 | ~new_P3_U3893;
  assign new_P3_U5517 = ~new_P3_U3404;
  assign new_P3_U5518 = ~P3_REG0_REG_5_ | ~new_P3_U3835;
  assign new_P3_U5519 = ~new_P3_U3914 | ~new_P3_U4174;
  assign new_P3_U5520 = ~P3_IR_REG_6_ | ~new_P3_U3831;
  assign new_P3_U5521 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U25;
  assign new_P3_U5522 = ~new_U33 | ~new_P3_U3833;
  assign new_P3_U5523 = ~new_P3_U3406 | ~new_P3_U3893;
  assign new_P3_U5524 = ~new_P3_U3407;
  assign new_P3_U5525 = ~P3_REG0_REG_6_ | ~new_P3_U3835;
  assign new_P3_U5526 = ~new_P3_U3914 | ~new_P3_U4192;
  assign new_P3_U5527 = ~P3_IR_REG_7_ | ~new_P3_U3831;
  assign new_P3_U5528 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U26;
  assign new_P3_U5529 = ~new_U32 | ~new_P3_U3833;
  assign new_P3_U5530 = ~new_P3_U3409 | ~new_P3_U3893;
  assign new_P3_U5531 = ~new_P3_U3410;
  assign new_P3_U5532 = ~P3_REG0_REG_7_ | ~new_P3_U3835;
  assign new_P3_U5533 = ~new_P3_U3914 | ~new_P3_U4210;
  assign new_P3_U5534 = ~P3_IR_REG_8_ | ~new_P3_U3831;
  assign new_P3_U5535 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U27;
  assign new_P3_U5536 = ~new_U31 | ~new_P3_U3833;
  assign new_P3_U5537 = ~new_P3_U3412 | ~new_P3_U3893;
  assign new_P3_U5538 = ~new_P3_U3413;
  assign new_P3_U5539 = ~P3_REG0_REG_8_ | ~new_P3_U3835;
  assign new_P3_U5540 = ~new_P3_U3914 | ~new_P3_U4228;
  assign new_P3_U5541 = ~P3_IR_REG_9_ | ~new_P3_U3831;
  assign new_P3_U5542 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U72;
  assign new_P3_U5543 = ~new_U30 | ~new_P3_U3833;
  assign new_P3_U5544 = ~new_P3_U3415 | ~new_P3_U3893;
  assign new_P3_U5545 = ~new_P3_U3416;
  assign new_P3_U5546 = ~P3_REG0_REG_9_ | ~new_P3_U3835;
  assign new_P3_U5547 = ~new_P3_U3914 | ~new_P3_U4246;
  assign new_P3_U5548 = ~P3_IR_REG_10_ | ~new_P3_U3831;
  assign new_P3_U5549 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U7;
  assign new_P3_U5550 = ~new_U60 | ~new_P3_U3833;
  assign new_P3_U5551 = ~new_P3_U3418 | ~new_P3_U3893;
  assign new_P3_U5552 = ~new_P3_U3419;
  assign new_P3_U5553 = ~P3_REG0_REG_10_ | ~new_P3_U3835;
  assign new_P3_U5554 = ~new_P3_U3914 | ~new_P3_U4264;
  assign new_P3_U5555 = ~P3_IR_REG_11_ | ~new_P3_U3831;
  assign new_P3_U5556 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U8;
  assign new_P3_U5557 = ~new_U59 | ~new_P3_U3833;
  assign new_P3_U5558 = ~new_P3_U3421 | ~new_P3_U3893;
  assign new_P3_U5559 = ~new_P3_U3422;
  assign new_P3_U5560 = ~P3_REG0_REG_11_ | ~new_P3_U3835;
  assign new_P3_U5561 = ~new_P3_U3914 | ~new_P3_U4282;
  assign new_P3_U5562 = ~P3_IR_REG_12_ | ~new_P3_U3831;
  assign new_P3_U5563 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U9;
  assign new_P3_U5564 = ~new_U58 | ~new_P3_U3833;
  assign new_P3_U5565 = ~new_P3_U3424 | ~new_P3_U3893;
  assign new_P3_U5566 = ~new_P3_U3425;
  assign new_P3_U5567 = ~P3_REG0_REG_12_ | ~new_P3_U3835;
  assign new_P3_U5568 = ~new_P3_U3914 | ~new_P3_U4300;
  assign new_P3_U5569 = ~P3_IR_REG_13_ | ~new_P3_U3831;
  assign new_P3_U5570 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U89;
  assign new_P3_U5571 = ~new_U57 | ~new_P3_U3833;
  assign new_P3_U5572 = ~new_P3_U3427 | ~new_P3_U3893;
  assign new_P3_U5573 = ~new_P3_U3428;
  assign new_P3_U5574 = ~P3_REG0_REG_13_ | ~new_P3_U3835;
  assign new_P3_U5575 = ~new_P3_U3914 | ~new_P3_U4318;
  assign new_P3_U5576 = ~P3_IR_REG_14_ | ~new_P3_U3831;
  assign new_P3_U5577 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U10;
  assign new_P3_U5578 = ~new_U56 | ~new_P3_U3833;
  assign new_P3_U5579 = ~new_P3_U3430 | ~new_P3_U3893;
  assign new_P3_U5580 = ~new_P3_U3431;
  assign new_P3_U5581 = ~P3_REG0_REG_14_ | ~new_P3_U3835;
  assign new_P3_U5582 = ~new_P3_U3914 | ~new_P3_U4336;
  assign new_P3_U5583 = ~P3_IR_REG_15_ | ~new_P3_U3831;
  assign new_P3_U5584 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U11;
  assign new_P3_U5585 = ~new_U55 | ~new_P3_U3833;
  assign new_P3_U5586 = ~new_P3_U3433 | ~new_P3_U3893;
  assign new_P3_U5587 = ~new_P3_U3434;
  assign new_P3_U5588 = ~P3_REG0_REG_15_ | ~new_P3_U3835;
  assign new_P3_U5589 = ~new_P3_U3914 | ~new_P3_U4354;
  assign new_P3_U5590 = ~P3_IR_REG_16_ | ~new_P3_U3831;
  assign new_P3_U5591 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U12;
  assign new_P3_U5592 = ~new_U54 | ~new_P3_U3833;
  assign new_P3_U5593 = ~new_P3_U3436 | ~new_P3_U3893;
  assign new_P3_U5594 = ~new_P3_U3437;
  assign new_P3_U5595 = ~P3_REG0_REG_16_ | ~new_P3_U3835;
  assign new_P3_U5596 = ~new_P3_U3914 | ~new_P3_U4372;
  assign new_P3_U5597 = ~P3_IR_REG_17_ | ~new_P3_U3831;
  assign new_P3_U5598 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U87;
  assign new_P3_U5599 = ~new_U53 | ~new_P3_U3833;
  assign new_P3_U5600 = ~new_P3_U3439 | ~new_P3_U3893;
  assign new_P3_U5601 = ~new_P3_U3440;
  assign new_P3_U5602 = ~P3_REG0_REG_17_ | ~new_P3_U3835;
  assign new_P3_U5603 = ~new_P3_U3914 | ~new_P3_U4390;
  assign new_P3_U5604 = ~P3_IR_REG_18_ | ~new_P3_U3831;
  assign new_P3_U5605 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U13;
  assign new_P3_U5606 = ~new_U52 | ~new_P3_U3833;
  assign new_P3_U5607 = ~new_P3_U3442 | ~new_P3_U3893;
  assign new_P3_U5608 = ~new_P3_U3443;
  assign new_P3_U5609 = ~P3_REG0_REG_18_ | ~new_P3_U3835;
  assign new_P3_U5610 = ~new_P3_U3914 | ~new_P3_U4408;
  assign new_P3_U5611 = ~new_U51 | ~new_P3_U3833;
  assign new_P3_U5612 = ~new_P3_U3893 | ~new_P3_U3379;
  assign new_P3_U5613 = ~new_P3_U3445;
  assign new_P3_U5614 = ~P3_REG0_REG_19_ | ~new_P3_U3835;
  assign new_P3_U5615 = ~new_P3_U3914 | ~new_P3_U4426;
  assign new_P3_U5616 = ~P3_REG0_REG_20_ | ~new_P3_U3835;
  assign new_P3_U5617 = ~new_P3_U3914 | ~new_P3_U4444;
  assign new_P3_U5618 = ~P3_REG0_REG_21_ | ~new_P3_U3835;
  assign new_P3_U5619 = ~new_P3_U3914 | ~new_P3_U4462;
  assign new_P3_U5620 = ~P3_REG0_REG_22_ | ~new_P3_U3835;
  assign new_P3_U5621 = ~new_P3_U3914 | ~new_P3_U4480;
  assign new_P3_U5622 = ~P3_REG0_REG_23_ | ~new_P3_U3835;
  assign new_P3_U5623 = ~new_P3_U3914 | ~new_P3_U4498;
  assign new_P3_U5624 = ~P3_REG0_REG_24_ | ~new_P3_U3835;
  assign new_P3_U5625 = ~new_P3_U3914 | ~new_P3_U4516;
  assign new_P3_U5626 = ~P3_REG0_REG_25_ | ~new_P3_U3835;
  assign new_P3_U5627 = ~new_P3_U3914 | ~new_P3_U4534;
  assign new_P3_U5628 = ~P3_REG0_REG_26_ | ~new_P3_U3835;
  assign new_P3_U5629 = ~new_P3_U3914 | ~new_P3_U4552;
  assign new_P3_U5630 = ~P3_REG0_REG_27_ | ~new_P3_U3835;
  assign new_P3_U5631 = ~new_P3_U3914 | ~new_P3_U4570;
  assign new_P3_U5632 = ~P3_REG0_REG_28_ | ~new_P3_U3835;
  assign new_P3_U5633 = ~new_P3_U3914 | ~new_P3_U4588;
  assign new_P3_U5634 = ~P3_REG0_REG_29_ | ~new_P3_U3835;
  assign new_P3_U5635 = ~new_P3_U3914 | ~new_P3_U4608;
  assign new_P3_U5636 = ~P3_REG0_REG_30_ | ~new_P3_U3835;
  assign new_P3_U5637 = ~new_P3_U3914 | ~new_P3_U4615;
  assign new_P3_U5638 = ~P3_REG0_REG_31_ | ~new_P3_U3835;
  assign new_P3_U5639 = ~new_P3_U3914 | ~new_P3_U4617;
  assign new_P3_U5640 = ~new_P3_U5453 | ~new_P3_U3834;
  assign new_P3_U5641 = ~new_P3_U4052 | ~new_P3_U5450;
  assign new_P3_U5642 = ~P3_REG1_REG_0_ | ~new_P3_U3836;
  assign new_P3_U5643 = ~new_P3_U3913 | ~new_P3_U4077;
  assign new_P3_U5644 = ~P3_REG1_REG_1_ | ~new_P3_U3836;
  assign new_P3_U5645 = ~new_P3_U3913 | ~new_P3_U4102;
  assign new_P3_U5646 = ~P3_REG1_REG_2_ | ~new_P3_U3836;
  assign new_P3_U5647 = ~new_P3_U3913 | ~new_P3_U4120;
  assign new_P3_U5648 = ~P3_REG1_REG_3_ | ~new_P3_U3836;
  assign new_P3_U5649 = ~new_P3_U3913 | ~new_P3_U4138;
  assign new_P3_U5650 = ~P3_REG1_REG_4_ | ~new_P3_U3836;
  assign new_P3_U5651 = ~new_P3_U3913 | ~new_P3_U4156;
  assign new_P3_U5652 = ~P3_REG1_REG_5_ | ~new_P3_U3836;
  assign new_P3_U5653 = ~new_P3_U3913 | ~new_P3_U4174;
  assign new_P3_U5654 = ~P3_REG1_REG_6_ | ~new_P3_U3836;
  assign new_P3_U5655 = ~new_P3_U3913 | ~new_P3_U4192;
  assign new_P3_U5656 = ~P3_REG1_REG_7_ | ~new_P3_U3836;
  assign new_P3_U5657 = ~new_P3_U3913 | ~new_P3_U4210;
  assign new_P3_U5658 = ~P3_REG1_REG_8_ | ~new_P3_U3836;
  assign new_P3_U5659 = ~new_P3_U3913 | ~new_P3_U4228;
  assign new_P3_U5660 = ~P3_REG1_REG_9_ | ~new_P3_U3836;
  assign new_P3_U5661 = ~new_P3_U3913 | ~new_P3_U4246;
  assign new_P3_U5662 = ~P3_REG1_REG_10_ | ~new_P3_U3836;
  assign new_P3_U5663 = ~new_P3_U3913 | ~new_P3_U4264;
  assign new_P3_U5664 = ~P3_REG1_REG_11_ | ~new_P3_U3836;
  assign new_P3_U5665 = ~new_P3_U3913 | ~new_P3_U4282;
  assign new_P3_U5666 = ~P3_REG1_REG_12_ | ~new_P3_U3836;
  assign new_P3_U5667 = ~new_P3_U3913 | ~new_P3_U4300;
  assign new_P3_U5668 = ~P3_REG1_REG_13_ | ~new_P3_U3836;
  assign new_P3_U5669 = ~new_P3_U3913 | ~new_P3_U4318;
  assign new_P3_U5670 = ~P3_REG1_REG_14_ | ~new_P3_U3836;
  assign new_P3_U5671 = ~new_P3_U3913 | ~new_P3_U4336;
  assign new_P3_U5672 = ~P3_REG1_REG_15_ | ~new_P3_U3836;
  assign new_P3_U5673 = ~new_P3_U3913 | ~new_P3_U4354;
  assign new_P3_U5674 = ~P3_REG1_REG_16_ | ~new_P3_U3836;
  assign new_P3_U5675 = ~new_P3_U3913 | ~new_P3_U4372;
  assign new_P3_U5676 = ~P3_REG1_REG_17_ | ~new_P3_U3836;
  assign new_P3_U5677 = ~new_P3_U3913 | ~new_P3_U4390;
  assign new_P3_U5678 = ~P3_REG1_REG_18_ | ~new_P3_U3836;
  assign new_P3_U5679 = ~new_P3_U3913 | ~new_P3_U4408;
  assign new_P3_U5680 = ~P3_REG1_REG_19_ | ~new_P3_U3836;
  assign new_P3_U5681 = ~new_P3_U3913 | ~new_P3_U4426;
  assign new_P3_U5682 = ~P3_REG1_REG_20_ | ~new_P3_U3836;
  assign new_P3_U5683 = ~new_P3_U3913 | ~new_P3_U4444;
  assign new_P3_U5684 = ~P3_REG1_REG_21_ | ~new_P3_U3836;
  assign new_P3_U5685 = ~new_P3_U3913 | ~new_P3_U4462;
  assign new_P3_U5686 = ~P3_REG1_REG_22_ | ~new_P3_U3836;
  assign new_P3_U5687 = ~new_P3_U3913 | ~new_P3_U4480;
  assign new_P3_U5688 = ~P3_REG1_REG_23_ | ~new_P3_U3836;
  assign new_P3_U5689 = ~new_P3_U3913 | ~new_P3_U4498;
  assign new_P3_U5690 = ~P3_REG1_REG_24_ | ~new_P3_U3836;
  assign new_P3_U5691 = ~new_P3_U3913 | ~new_P3_U4516;
  assign new_P3_U5692 = ~P3_REG1_REG_25_ | ~new_P3_U3836;
  assign new_P3_U5693 = ~new_P3_U3913 | ~new_P3_U4534;
  assign new_P3_U5694 = ~P3_REG1_REG_26_ | ~new_P3_U3836;
  assign new_P3_U5695 = ~new_P3_U3913 | ~new_P3_U4552;
  assign new_P3_U5696 = ~P3_REG1_REG_27_ | ~new_P3_U3836;
  assign new_P3_U5697 = ~new_P3_U3913 | ~new_P3_U4570;
  assign new_P3_U5698 = ~P3_REG1_REG_28_ | ~new_P3_U3836;
  assign new_P3_U5699 = ~new_P3_U3913 | ~new_P3_U4588;
  assign new_P3_U5700 = ~P3_REG1_REG_29_ | ~new_P3_U3836;
  assign new_P3_U5701 = ~new_P3_U3913 | ~new_P3_U4608;
  assign new_P3_U5702 = ~P3_REG1_REG_30_ | ~new_P3_U3836;
  assign new_P3_U5703 = ~new_P3_U3913 | ~new_P3_U4615;
  assign new_P3_U5704 = ~P3_REG1_REG_31_ | ~new_P3_U3836;
  assign new_P3_U5705 = ~new_P3_U3913 | ~new_P3_U4617;
  assign new_P3_U5706 = ~P3_REG2_REG_0_ | ~new_P3_U3358;
  assign new_P3_U5707 = ~new_P3_U3912 | ~new_P3_U3314;
  assign new_P3_U5708 = ~P3_REG2_REG_1_ | ~new_P3_U3358;
  assign new_P3_U5709 = ~new_P3_U3912 | ~new_P3_U3315;
  assign new_P3_U5710 = ~P3_REG2_REG_2_ | ~new_P3_U3358;
  assign new_P3_U5711 = ~new_P3_U3912 | ~new_P3_U3316;
  assign new_P3_U5712 = ~P3_REG2_REG_3_ | ~new_P3_U3358;
  assign new_P3_U5713 = ~new_P3_U3912 | ~new_P3_U3317;
  assign new_P3_U5714 = ~P3_REG2_REG_4_ | ~new_P3_U3358;
  assign new_P3_U5715 = ~new_P3_U3912 | ~new_P3_U3318;
  assign new_P3_U5716 = ~P3_REG2_REG_5_ | ~new_P3_U3358;
  assign new_P3_U5717 = ~new_P3_U3912 | ~new_P3_U3319;
  assign new_P3_U5718 = ~P3_REG2_REG_6_ | ~new_P3_U3358;
  assign new_P3_U5719 = ~new_P3_U3912 | ~new_P3_U3320;
  assign new_P3_U5720 = ~P3_REG2_REG_7_ | ~new_P3_U3358;
  assign new_P3_U5721 = ~new_P3_U3912 | ~new_P3_U3321;
  assign new_P3_U5722 = ~P3_REG2_REG_8_ | ~new_P3_U3358;
  assign new_P3_U5723 = ~new_P3_U3912 | ~new_P3_U3322;
  assign new_P3_U5724 = ~P3_REG2_REG_9_ | ~new_P3_U3358;
  assign new_P3_U5725 = ~new_P3_U3912 | ~new_P3_U3323;
  assign new_P3_U5726 = ~P3_REG2_REG_10_ | ~new_P3_U3358;
  assign new_P3_U5727 = ~new_P3_U3912 | ~new_P3_U3324;
  assign new_P3_U5728 = ~P3_REG2_REG_11_ | ~new_P3_U3358;
  assign new_P3_U5729 = ~new_P3_U3912 | ~new_P3_U3325;
  assign new_P3_U5730 = ~P3_REG2_REG_12_ | ~new_P3_U3358;
  assign new_P3_U5731 = ~new_P3_U3912 | ~new_P3_U3326;
  assign new_P3_U5732 = ~P3_REG2_REG_13_ | ~new_P3_U3358;
  assign new_P3_U5733 = ~new_P3_U3912 | ~new_P3_U3327;
  assign new_P3_U5734 = ~P3_REG2_REG_14_ | ~new_P3_U3358;
  assign new_P3_U5735 = ~new_P3_U3912 | ~new_P3_U3328;
  assign new_P3_U5736 = ~P3_REG2_REG_15_ | ~new_P3_U3358;
  assign new_P3_U5737 = ~new_P3_U3912 | ~new_P3_U3329;
  assign new_P3_U5738 = ~P3_REG2_REG_16_ | ~new_P3_U3358;
  assign new_P3_U5739 = ~new_P3_U3912 | ~new_P3_U3330;
  assign new_P3_U5740 = ~P3_REG2_REG_17_ | ~new_P3_U3358;
  assign new_P3_U5741 = ~new_P3_U3912 | ~new_P3_U3331;
  assign new_P3_U5742 = ~P3_REG2_REG_18_ | ~new_P3_U3358;
  assign new_P3_U5743 = ~new_P3_U3912 | ~new_P3_U3332;
  assign new_P3_U5744 = ~P3_REG2_REG_19_ | ~new_P3_U3358;
  assign new_P3_U5745 = ~new_P3_U3912 | ~new_P3_U3333;
  assign new_P3_U5746 = ~P3_REG2_REG_20_ | ~new_P3_U3358;
  assign new_P3_U5747 = ~new_P3_U3912 | ~new_P3_U3335;
  assign new_P3_U5748 = ~P3_REG2_REG_21_ | ~new_P3_U3358;
  assign new_P3_U5749 = ~new_P3_U3912 | ~new_P3_U3337;
  assign new_P3_U5750 = ~P3_REG2_REG_22_ | ~new_P3_U3358;
  assign new_P3_U5751 = ~new_P3_U3912 | ~new_P3_U3339;
  assign new_P3_U5752 = ~P3_REG2_REG_23_ | ~new_P3_U3358;
  assign new_P3_U5753 = ~new_P3_U3912 | ~new_P3_U3341;
  assign new_P3_U5754 = ~P3_REG2_REG_24_ | ~new_P3_U3358;
  assign new_P3_U5755 = ~new_P3_U3912 | ~new_P3_U3343;
  assign new_P3_U5756 = ~P3_REG2_REG_25_ | ~new_P3_U3358;
  assign new_P3_U5757 = ~new_P3_U3912 | ~new_P3_U3345;
  assign new_P3_U5758 = ~P3_REG2_REG_26_ | ~new_P3_U3358;
  assign new_P3_U5759 = ~new_P3_U3912 | ~new_P3_U3347;
  assign new_P3_U5760 = ~P3_REG2_REG_27_ | ~new_P3_U3358;
  assign new_P3_U5761 = ~new_P3_U3912 | ~new_P3_U3349;
  assign new_P3_U5762 = ~P3_REG2_REG_28_ | ~new_P3_U3358;
  assign new_P3_U5763 = ~new_P3_U3912 | ~new_P3_U3351;
  assign new_P3_U5764 = ~P3_REG2_REG_29_ | ~new_P3_U3358;
  assign new_P3_U5765 = ~new_P3_U3912 | ~new_P3_U3354;
  assign new_P3_U5766 = ~new_P3_U5465 | ~new_P3_U3024;
  assign new_P3_U5767 = ~new_P3_U3383 | ~n3844;
  assign new_P3_U5768 = ~new_P3_U5767 | ~new_P3_U5766;
  assign new_P3_U5769 = ~P3_DATAO_REG_0_ | ~new_P3_U3363;
  assign new_P3_U5770 = ~n3844 | ~new_P3_U3076;
  assign new_P3_U5771 = ~P3_DATAO_REG_1_ | ~new_P3_U3363;
  assign new_P3_U5772 = ~n3844 | ~new_P3_U3077;
  assign new_P3_U5773 = ~P3_DATAO_REG_2_ | ~new_P3_U3363;
  assign new_P3_U5774 = ~n3844 | ~new_P3_U3067;
  assign new_P3_U5775 = ~P3_DATAO_REG_3_ | ~new_P3_U3363;
  assign new_P3_U5776 = ~n3844 | ~new_P3_U3063;
  assign new_P3_U5777 = ~P3_DATAO_REG_4_ | ~new_P3_U3363;
  assign new_P3_U5778 = ~n3844 | ~new_P3_U3059;
  assign new_P3_U5779 = ~P3_DATAO_REG_5_ | ~new_P3_U3363;
  assign new_P3_U5780 = ~n3844 | ~new_P3_U3066;
  assign new_P3_U5781 = ~P3_DATAO_REG_6_ | ~new_P3_U3363;
  assign new_P3_U5782 = ~n3844 | ~new_P3_U3070;
  assign new_P3_U5783 = ~P3_DATAO_REG_7_ | ~new_P3_U3363;
  assign new_P3_U5784 = ~n3844 | ~new_P3_U3069;
  assign new_P3_U5785 = ~P3_DATAO_REG_8_ | ~new_P3_U3363;
  assign new_P3_U5786 = ~n3844 | ~new_P3_U3083;
  assign new_P3_U5787 = ~P3_DATAO_REG_9_ | ~new_P3_U3363;
  assign new_P3_U5788 = ~n3844 | ~new_P3_U3082;
  assign new_P3_U5789 = ~P3_DATAO_REG_10_ | ~new_P3_U3363;
  assign new_P3_U5790 = ~n3844 | ~new_P3_U3061;
  assign new_P3_U5791 = ~P3_DATAO_REG_11_ | ~new_P3_U3363;
  assign new_P3_U5792 = ~n3844 | ~new_P3_U3062;
  assign new_P3_U5793 = ~P3_DATAO_REG_12_ | ~new_P3_U3363;
  assign new_P3_U5794 = ~n3844 | ~new_P3_U3071;
  assign new_P3_U5795 = ~P3_DATAO_REG_13_ | ~new_P3_U3363;
  assign new_P3_U5796 = ~n3844 | ~new_P3_U3079;
  assign new_P3_U5797 = ~P3_DATAO_REG_14_ | ~new_P3_U3363;
  assign new_P3_U5798 = ~n3844 | ~new_P3_U3078;
  assign new_P3_U5799 = ~P3_DATAO_REG_15_ | ~new_P3_U3363;
  assign new_P3_U5800 = ~n3844 | ~new_P3_U3073;
  assign new_P3_U5801 = ~P3_DATAO_REG_16_ | ~new_P3_U3363;
  assign new_P3_U5802 = ~n3844 | ~new_P3_U3072;
  assign new_P3_U5803 = ~P3_DATAO_REG_17_ | ~new_P3_U3363;
  assign new_P3_U5804 = ~n3844 | ~new_P3_U3068;
  assign new_P3_U5805 = ~P3_DATAO_REG_18_ | ~new_P3_U3363;
  assign new_P3_U5806 = ~n3844 | ~new_P3_U3081;
  assign new_P3_U5807 = ~P3_DATAO_REG_19_ | ~new_P3_U3363;
  assign new_P3_U5808 = ~n3844 | ~new_P3_U3080;
  assign new_P3_U5809 = ~P3_DATAO_REG_20_ | ~new_P3_U3363;
  assign new_P3_U5810 = ~n3844 | ~new_P3_U3075;
  assign new_P3_U5811 = ~P3_DATAO_REG_21_ | ~new_P3_U3363;
  assign new_P3_U5812 = ~n3844 | ~new_P3_U3074;
  assign new_P3_U5813 = ~P3_DATAO_REG_22_ | ~new_P3_U3363;
  assign new_P3_U5814 = ~n3844 | ~new_P3_U3060;
  assign new_P3_U5815 = ~P3_DATAO_REG_23_ | ~new_P3_U3363;
  assign new_P3_U5816 = ~n3844 | ~new_P3_U3065;
  assign new_P3_U5817 = ~P3_DATAO_REG_24_ | ~new_P3_U3363;
  assign new_P3_U5818 = ~n3844 | ~new_P3_U3064;
  assign new_P3_U5819 = ~P3_DATAO_REG_25_ | ~new_P3_U3363;
  assign new_P3_U5820 = ~n3844 | ~new_P3_U3057;
  assign new_P3_U5821 = ~P3_DATAO_REG_26_ | ~new_P3_U3363;
  assign new_P3_U5822 = ~n3844 | ~new_P3_U3056;
  assign new_P3_U5823 = ~P3_DATAO_REG_27_ | ~new_P3_U3363;
  assign new_P3_U5824 = ~n3844 | ~new_P3_U3052;
  assign new_P3_U5825 = ~P3_DATAO_REG_28_ | ~new_P3_U3363;
  assign new_P3_U5826 = ~n3844 | ~new_P3_U3053;
  assign new_P3_U5827 = ~P3_DATAO_REG_29_ | ~new_P3_U3363;
  assign new_P3_U5828 = ~n3844 | ~new_P3_U3054;
  assign new_P3_U5829 = ~P3_DATAO_REG_30_ | ~new_P3_U3363;
  assign new_P3_U5830 = ~n3844 | ~new_P3_U3058;
  assign new_P3_U5831 = ~P3_DATAO_REG_31_ | ~new_P3_U3363;
  assign new_P3_U5832 = ~n3844 | ~new_P3_U3055;
  assign new_P3_U5833 = ~new_P3_U3379 | ~new_P3_U3313;
  assign new_P3_U5834 = ~new_P3_U5450 | ~new_P3_U3911;
  assign new_P3_U5835 = ~new_P3_U3760;
  assign new_P3_U5836 = ~new_P3_R1269_U11 | ~new_P3_U5835;
  assign new_P3_U5837 = ~new_P3_U3760 | ~new_P3_U3867;
  assign new_P3_U5838 = ~new_P3_U3900 | ~new_P3_U3052;
  assign new_P3_U5839 = ~new_P3_U3348 | ~new_P3_U4539;
  assign new_P3_U5840 = ~new_P3_U5839 | ~new_P3_U5838;
  assign new_P3_U5841 = ~new_P3_U3899 | ~new_P3_U3053;
  assign new_P3_U5842 = ~new_P3_U3350 | ~new_P3_U4557;
  assign new_P3_U5843 = ~new_P3_U5842 | ~new_P3_U5841;
  assign new_P3_U5844 = ~new_P3_U3872 | ~new_P3_U3055;
  assign new_P3_U5845 = ~new_P3_U3356 | ~new_P3_U4613;
  assign new_P3_U5846 = ~new_P3_U5845 | ~new_P3_U5844;
  assign new_P3_U5847 = ~new_P3_U3908 | ~new_P3_U3054;
  assign new_P3_U5848 = ~new_P3_U3353 | ~new_P3_U4575;
  assign new_P3_U5849 = ~new_P3_U5848 | ~new_P3_U5847;
  assign new_P3_U5850 = ~new_P3_U3906 | ~new_P3_U3074;
  assign new_P3_U5851 = ~new_P3_U3336 | ~new_P3_U4431;
  assign new_P3_U5852 = ~new_P3_U5851 | ~new_P3_U5850;
  assign new_P3_U5853 = ~new_P3_U3907 | ~new_P3_U3075;
  assign new_P3_U5854 = ~new_P3_U3334 | ~new_P3_U4413;
  assign new_P3_U5855 = ~new_P3_U5854 | ~new_P3_U5853;
  assign new_P3_U5856 = ~new_P3_U5503 | ~new_P3_U4107;
  assign new_P3_U5857 = ~new_P3_U3398 | ~new_P3_U3063;
  assign new_P3_U5858 = ~new_P3_U5857 | ~new_P3_U5856;
  assign new_P3_U5859 = ~new_P3_U5559 | ~new_P3_U4251;
  assign new_P3_U5860 = ~new_P3_U3422 | ~new_P3_U3062;
  assign new_P3_U5861 = ~new_P3_U5860 | ~new_P3_U5859;
  assign new_P3_U5862 = ~new_P3_U5552 | ~new_P3_U4233;
  assign new_P3_U5863 = ~new_P3_U3419 | ~new_P3_U3061;
  assign new_P3_U5864 = ~new_P3_U5863 | ~new_P3_U5862;
  assign new_P3_U5865 = ~new_P3_U5510 | ~new_P3_U4125;
  assign new_P3_U5866 = ~new_P3_U3401 | ~new_P3_U3059;
  assign new_P3_U5867 = ~new_P3_U5866 | ~new_P3_U5865;
  assign new_P3_U5868 = ~new_P3_U3905 | ~new_P3_U3060;
  assign new_P3_U5869 = ~new_P3_U3338 | ~new_P3_U4449;
  assign new_P3_U5870 = ~new_P3_U5869 | ~new_P3_U5868;
  assign new_P3_U5871 = ~new_P3_U5601 | ~new_P3_U4359;
  assign new_P3_U5872 = ~new_P3_U3440 | ~new_P3_U3068;
  assign new_P3_U5873 = ~new_P3_U5872 | ~new_P3_U5871;
  assign new_P3_U5874 = ~new_P3_U5594 | ~new_P3_U4341;
  assign new_P3_U5875 = ~new_P3_U3437 | ~new_P3_U3072;
  assign new_P3_U5876 = ~new_P3_U5875 | ~new_P3_U5874;
  assign new_P3_U5877 = ~new_P3_U5587 | ~new_P3_U4323;
  assign new_P3_U5878 = ~new_P3_U3434 | ~new_P3_U3073;
  assign new_P3_U5879 = ~new_P3_U5878 | ~new_P3_U5877;
  assign new_P3_U5880 = ~new_P3_U5566 | ~new_P3_U4269;
  assign new_P3_U5881 = ~new_P3_U3425 | ~new_P3_U3071;
  assign new_P3_U5882 = ~new_P3_U5881 | ~new_P3_U5880;
  assign new_P3_U5883 = ~new_P3_U5524 | ~new_P3_U4161;
  assign new_P3_U5884 = ~new_P3_U3407 | ~new_P3_U3070;
  assign new_P3_U5885 = ~new_P3_U5884 | ~new_P3_U5883;
  assign new_P3_U5886 = ~new_P3_U5531 | ~new_P3_U4179;
  assign new_P3_U5887 = ~new_P3_U3410 | ~new_P3_U3069;
  assign new_P3_U5888 = ~new_P3_U5887 | ~new_P3_U5886;
  assign new_P3_U5889 = ~new_P3_U5496 | ~new_P3_U4082;
  assign new_P3_U5890 = ~new_P3_U3395 | ~new_P3_U3067;
  assign new_P3_U5891 = ~new_P3_U5890 | ~new_P3_U5889;
  assign new_P3_U5892 = ~new_P3_U5517 | ~new_P3_U4143;
  assign new_P3_U5893 = ~new_P3_U3404 | ~new_P3_U3066;
  assign new_P3_U5894 = ~new_P3_U5893 | ~new_P3_U5892;
  assign new_P3_U5895 = ~new_P3_U5608 | ~new_P3_U4377;
  assign new_P3_U5896 = ~new_P3_U3443 | ~new_P3_U3081;
  assign new_P3_U5897 = ~new_P3_U5896 | ~new_P3_U5895;
  assign new_P3_U5898 = ~new_P3_U5573 | ~new_P3_U4287;
  assign new_P3_U5899 = ~new_P3_U3428 | ~new_P3_U3079;
  assign new_P3_U5900 = ~new_P3_U5899 | ~new_P3_U5898;
  assign new_P3_U5901 = ~new_P3_U5580 | ~new_P3_U4305;
  assign new_P3_U5902 = ~new_P3_U3431 | ~new_P3_U3078;
  assign new_P3_U5903 = ~new_P3_U5902 | ~new_P3_U5901;
  assign new_P3_U5904 = ~new_P3_U5489 | ~new_P3_U4063;
  assign new_P3_U5905 = ~new_P3_U3392 | ~new_P3_U3077;
  assign new_P3_U5906 = ~new_P3_U5905 | ~new_P3_U5904;
  assign new_P3_U5907 = ~new_P3_U5473 | ~new_P3_U4087;
  assign new_P3_U5908 = ~new_P3_U3387 | ~new_P3_U3076;
  assign new_P3_U5909 = ~new_P3_U5908 | ~new_P3_U5907;
  assign new_P3_U5910 = ~new_P3_U5538 | ~new_P3_U4197;
  assign new_P3_U5911 = ~new_P3_U3413 | ~new_P3_U3083;
  assign new_P3_U5912 = ~new_P3_U5911 | ~new_P3_U5910;
  assign new_P3_U5913 = ~new_P3_U5545 | ~new_P3_U4215;
  assign new_P3_U5914 = ~new_P3_U3416 | ~new_P3_U3082;
  assign new_P3_U5915 = ~new_P3_U5914 | ~new_P3_U5913;
  assign new_P3_U5916 = ~new_P3_U5613 | ~new_P3_U4395;
  assign new_P3_U5917 = ~new_P3_U3445 | ~new_P3_U3080;
  assign new_P3_U5918 = ~new_P3_U5917 | ~new_P3_U5916;
  assign new_P3_U5919 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_U5920 = ~new_P3_U3346 | ~new_P3_U4521;
  assign new_P3_U5921 = ~new_P3_U5920 | ~new_P3_U5919;
  assign new_P3_U5922 = ~new_P3_U3902 | ~new_P3_U3057;
  assign new_P3_U5923 = ~new_P3_U3344 | ~new_P3_U4503;
  assign new_P3_U5924 = ~new_P3_U5923 | ~new_P3_U5922;
  assign new_P3_U5925 = ~new_P3_U3904 | ~new_P3_U3065;
  assign new_P3_U5926 = ~new_P3_U3340 | ~new_P3_U4467;
  assign new_P3_U5927 = ~new_P3_U5926 | ~new_P3_U5925;
  assign new_P3_U5928 = ~new_P3_U3903 | ~new_P3_U3064;
  assign new_P3_U5929 = ~new_P3_U3342 | ~new_P3_U4485;
  assign new_P3_U5930 = ~new_P3_U5929 | ~new_P3_U5928;
  assign new_P3_U5931 = ~new_P3_U3873 | ~new_P3_U3058;
  assign new_P3_U5932 = ~new_P3_U3355 | ~new_P3_U4593;
  assign new_P3_U5933 = ~new_P3_U5932 | ~new_P3_U5931;
  assign new_P3_U5934 = ~new_P3_U4978 | ~new_P3_U5450;
  assign new_P3_U5935 = ~new_P3_U3379 | ~new_P3_U3868;
  assign new_P3_U5936 = ~new_P3_U5935 | ~new_P3_U5934;
  assign new_P3_U5937 = ~new_P3_U5447 | ~new_P3_U5837 | ~new_P3_U5836;
  assign new_P3_U5938 = ~new_P3_U3378 | ~new_P3_U5456 | ~new_P3_U5936;
  assign new_P3_U5939 = ~new_P3_U3881 | ~new_P3_U3869;
  assign new_P3_U5940 = ~new_P3_R693_U14 | ~new_P3_U3891;
  assign new_P3_U5941 = ~new_P3_U5440 | ~new_P3_U3368;
  assign new_P3_U5942 = ~new_P3_U3380 | ~new_P3_U3375;
  assign new_P3_U5943 = ~new_P3_U5450 | ~new_P3_U5447;
  assign new_P3_U5944 = ~new_P3_U3378 | ~new_P3_U3388 | ~new_P3_U5456;
  assign new_P3_U5945 = ~new_P3_U3082 | ~new_P3_R1297_U6;
  assign new_P3_U5946 = ~new_P3_U3082 | ~new_P3_U3871;
  assign new_P3_U5947 = ~new_P3_U3083 | ~new_P3_R1297_U6;
  assign new_P3_U5948 = ~new_P3_U3083 | ~new_P3_U3871;
  assign new_P3_U5949 = ~new_P3_U3069 | ~new_P3_R1297_U6;
  assign new_P3_U5950 = ~new_P3_U3069 | ~new_P3_U3871;
  assign new_P3_U5951 = ~new_P3_U3070 | ~new_P3_R1297_U6;
  assign new_P3_U5952 = ~new_P3_U3070 | ~new_P3_U3871;
  assign new_P3_U5953 = ~new_P3_U3066 | ~new_P3_R1297_U6;
  assign new_P3_U5954 = ~new_P3_U3066 | ~new_P3_U3871;
  assign new_P3_U5955 = ~new_P3_U3059 | ~new_P3_R1297_U6;
  assign new_P3_U5956 = ~new_P3_U3059 | ~new_P3_U3871;
  assign new_P3_U5957 = ~new_P3_R1300_U8 | ~new_P3_R1297_U6;
  assign new_P3_U5958 = ~new_P3_U3055 | ~new_P3_U3871;
  assign new_P3_U5959 = ~new_P3_R1300_U6 | ~new_P3_R1297_U6;
  assign new_P3_U5960 = ~new_P3_U3058 | ~new_P3_U3871;
  assign new_P3_U5961 = ~new_P3_U3063 | ~new_P3_R1297_U6;
  assign new_P3_U5962 = ~new_P3_U3063 | ~new_P3_U3871;
  assign new_P3_U5963 = ~new_P3_U3054 | ~new_P3_R1297_U6;
  assign new_P3_U5964 = ~new_P3_U3054 | ~new_P3_U3871;
  assign new_P3_U5965 = ~new_P3_U3053 | ~new_P3_R1297_U6;
  assign new_P3_U5966 = ~new_P3_U3053 | ~new_P3_U3871;
  assign new_P3_U5967 = ~new_P3_U3052 | ~new_P3_R1297_U6;
  assign new_P3_U5968 = ~new_P3_U3052 | ~new_P3_U3871;
  assign new_P3_U5969 = ~new_P3_U3056 | ~new_P3_R1297_U6;
  assign new_P3_U5970 = ~new_P3_U3056 | ~new_P3_U3871;
  assign new_P3_U5971 = ~new_P3_U3057 | ~new_P3_R1297_U6;
  assign new_P3_U5972 = ~new_P3_U3057 | ~new_P3_U3871;
  assign new_P3_U5973 = ~new_P3_U3064 | ~new_P3_R1297_U6;
  assign new_P3_U5974 = ~new_P3_U3064 | ~new_P3_U3871;
  assign new_P3_U5975 = ~new_P3_U3065 | ~new_P3_R1297_U6;
  assign new_P3_U5976 = ~new_P3_U3065 | ~new_P3_U3871;
  assign new_P3_U5977 = ~new_P3_U3060 | ~new_P3_R1297_U6;
  assign new_P3_U5978 = ~new_P3_U3060 | ~new_P3_U3871;
  assign new_P3_U5979 = ~new_P3_U3074 | ~new_P3_R1297_U6;
  assign new_P3_U5980 = ~new_P3_U3074 | ~new_P3_U3871;
  assign new_P3_U5981 = ~new_P3_U3075 | ~new_P3_R1297_U6;
  assign new_P3_U5982 = ~new_P3_U3075 | ~new_P3_U3871;
  assign new_P3_U5983 = ~new_P3_U3067 | ~new_P3_R1297_U6;
  assign new_P3_U5984 = ~new_P3_U3067 | ~new_P3_U3871;
  assign new_P3_U5985 = ~new_P3_U3080 | ~new_P3_R1297_U6;
  assign new_P3_U5986 = ~new_P3_U3080 | ~new_P3_U3871;
  assign new_P3_U5987 = ~new_P3_U3081 | ~new_P3_R1297_U6;
  assign new_P3_U5988 = ~new_P3_U3081 | ~new_P3_U3871;
  assign new_P3_U5989 = ~new_P3_U3068 | ~new_P3_R1297_U6;
  assign new_P3_U5990 = ~new_P3_U3068 | ~new_P3_U3871;
  assign new_P3_U5991 = ~new_P3_U3072 | ~new_P3_R1297_U6;
  assign new_P3_U5992 = ~new_P3_U3072 | ~new_P3_U3871;
  assign new_P3_U5993 = ~new_P3_U3073 | ~new_P3_R1297_U6;
  assign new_P3_U5994 = ~new_P3_U3073 | ~new_P3_U3871;
  assign new_P3_U5995 = ~new_P3_U3078 | ~new_P3_R1297_U6;
  assign new_P3_U5996 = ~new_P3_U3078 | ~new_P3_U3871;
  assign new_P3_U5997 = ~new_P3_U3079 | ~new_P3_R1297_U6;
  assign new_P3_U5998 = ~new_P3_U3079 | ~new_P3_U3871;
  assign new_P3_U5999 = ~new_P3_U3071 | ~new_P3_R1297_U6;
  assign new_P3_U6000 = ~new_P3_U3071 | ~new_P3_U3871;
  assign new_P3_U6001 = ~new_P3_U3062 | ~new_P3_R1297_U6;
  assign new_P3_U6002 = ~new_P3_U3062 | ~new_P3_U3871;
  assign new_P3_U6003 = ~new_P3_U3061 | ~new_P3_R1297_U6;
  assign new_P3_U6004 = ~new_P3_U3061 | ~new_P3_U3871;
  assign new_P3_U6005 = ~new_P3_U3077 | ~new_P3_R1297_U6;
  assign new_P3_U6006 = ~new_P3_U3077 | ~new_P3_U3871;
  assign new_P3_U6007 = ~new_P3_U3076 | ~new_P3_R1297_U6;
  assign new_P3_U6008 = ~new_P3_U3076 | ~new_P3_U3871;
  assign new_P3_U6009 = ~new_P3_U5468 | ~P3_REG1_REG_9_;
  assign new_P3_U6010 = ~new_P3_U3384 | ~P3_REG2_REG_9_;
  assign new_P3_U6011 = ~new_P3_U5468 | ~P3_REG1_REG_8_;
  assign new_P3_U6012 = ~new_P3_U3384 | ~P3_REG2_REG_8_;
  assign new_P3_U6013 = ~new_P3_U5468 | ~P3_REG1_REG_7_;
  assign new_P3_U6014 = ~new_P3_U3384 | ~P3_REG2_REG_7_;
  assign new_P3_U6015 = ~new_P3_U5468 | ~P3_REG1_REG_6_;
  assign new_P3_U6016 = ~new_P3_U3384 | ~P3_REG2_REG_6_;
  assign new_P3_U6017 = ~new_P3_U5468 | ~P3_REG1_REG_5_;
  assign new_P3_U6018 = ~new_P3_U3384 | ~P3_REG2_REG_5_;
  assign new_P3_U6019 = ~new_P3_U5468 | ~P3_REG1_REG_4_;
  assign new_P3_U6020 = ~new_P3_U3384 | ~P3_REG2_REG_4_;
  assign new_P3_U6021 = ~new_P3_U5468 | ~P3_REG1_REG_3_;
  assign new_P3_U6022 = ~new_P3_U3384 | ~P3_REG2_REG_3_;
  assign new_P3_U6023 = ~new_P3_U5468 | ~P3_REG1_REG_2_;
  assign new_P3_U6024 = ~new_P3_U3384 | ~P3_REG2_REG_2_;
  assign new_P3_U6025 = ~new_P3_U5468 | ~P3_REG1_REG_19_;
  assign new_P3_U6026 = ~new_P3_U3384 | ~P3_REG2_REG_19_;
  assign new_P3_U6027 = ~new_P3_U5468 | ~P3_REG1_REG_18_;
  assign new_P3_U6028 = ~new_P3_U3384 | ~P3_REG2_REG_18_;
  assign new_P3_U6029 = ~new_P3_U5468 | ~P3_REG1_REG_17_;
  assign new_P3_U6030 = ~new_P3_U3384 | ~P3_REG2_REG_17_;
  assign new_P3_U6031 = ~new_P3_U5468 | ~P3_REG1_REG_16_;
  assign new_P3_U6032 = ~new_P3_U3384 | ~P3_REG2_REG_16_;
  assign new_P3_U6033 = ~new_P3_U5468 | ~P3_REG1_REG_15_;
  assign new_P3_U6034 = ~new_P3_U3384 | ~P3_REG2_REG_15_;
  assign new_P3_U6035 = ~new_P3_U5468 | ~P3_REG1_REG_14_;
  assign new_P3_U6036 = ~new_P3_U3384 | ~P3_REG2_REG_14_;
  assign new_P3_U6037 = ~new_P3_U5468 | ~P3_REG1_REG_13_;
  assign new_P3_U6038 = ~new_P3_U3384 | ~P3_REG2_REG_13_;
  assign new_P3_U6039 = ~new_P3_U5468 | ~P3_REG1_REG_12_;
  assign new_P3_U6040 = ~new_P3_U3384 | ~P3_REG2_REG_12_;
  assign new_P3_U6041 = ~new_P3_U5468 | ~P3_REG1_REG_11_;
  assign new_P3_U6042 = ~new_P3_U3384 | ~P3_REG2_REG_11_;
  assign new_P3_U6043 = ~new_P3_U5468 | ~P3_REG1_REG_10_;
  assign new_P3_U6044 = ~new_P3_U3384 | ~P3_REG2_REG_10_;
  assign new_P3_U6045 = ~new_P3_U5468 | ~P3_REG1_REG_1_;
  assign new_P3_U6046 = ~new_P3_U3384 | ~P3_REG2_REG_1_;
  assign new_P3_U6047 = ~new_P3_U5468 | ~P3_REG1_REG_0_;
  assign new_P3_U6048 = ~new_P3_U3384 | ~P3_REG2_REG_0_;
  assign new_P3_R1161_U448 = ~new_P3_R1161_U286 | ~new_P3_R1161_U446;
  assign new_P3_R1161_U447 = ~new_P3_R1161_U158 | ~new_P3_R1161_U159;
  assign new_P3_R1161_U446 = ~new_P3_R1161_U445 | ~new_P3_R1161_U444;
  assign new_P3_R1161_U445 = ~new_P3_U3905 | ~new_P3_R1161_U83;
  assign new_P3_R1161_U444 = ~new_P3_U3060 | ~new_P3_R1161_U82;
  assign new_P3_R1161_U443 = ~new_P3_U3905 | ~new_P3_R1161_U83;
  assign new_P3_R1161_U442 = ~new_P3_U3060 | ~new_P3_R1161_U82;
  assign new_P3_R1161_U441 = ~new_P3_R1161_U290 | ~new_P3_R1161_U439;
  assign new_P3_R1161_U440 = ~new_P3_R1161_U156 | ~new_P3_R1161_U157;
  assign new_P3_R1161_U439 = ~new_P3_R1161_U438 | ~new_P3_R1161_U437;
  assign new_P3_R1161_U438 = ~new_P3_U3904 | ~new_P3_R1161_U85;
  assign new_P3_R1161_U437 = ~new_P3_U3065 | ~new_P3_R1161_U84;
  assign new_P3_R1161_U436 = ~new_P3_U3904 | ~new_P3_R1161_U85;
  assign new_P3_R1161_U435 = ~new_P3_U3065 | ~new_P3_R1161_U84;
  assign new_P3_R1161_U434 = ~new_P3_R1161_U294 | ~new_P3_R1161_U432;
  assign new_P3_R1161_U433 = ~new_P3_R1161_U358 | ~new_P3_R1161_U155;
  assign new_P3_R1161_U432 = ~new_P3_R1161_U431 | ~new_P3_R1161_U430;
  assign new_P3_R1161_U431 = ~new_P3_U3903 | ~new_P3_R1161_U53;
  assign new_P3_R1161_U430 = ~new_P3_U3064 | ~new_P3_R1161_U52;
  assign new_SUB_1605_U6 = new_SUB_1605_U194 & new_SUB_1605_U190;
  assign new_SUB_1605_U7 = new_SUB_1605_U202 & new_SUB_1605_U200;
  assign new_SUB_1605_U8 = new_SUB_1605_U7 & new_SUB_1605_U204;
  assign new_SUB_1605_U9 = new_SUB_1605_U212 & new_SUB_1605_U208;
  assign new_SUB_1605_U10 = new_SUB_1605_U9 & new_SUB_1605_U215;
  assign new_SUB_1605_U11 = new_SUB_1605_U363 & new_SUB_1605_U362;
  assign new_SUB_1605_U12 = ~new_SUB_1605_U128 | ~new_SUB_1605_U323;
  assign new_SUB_1605_U13 = ~new_SUB_1605_U175 | ~new_SUB_1605_U291;
  assign new_SUB_1605_U14 = ~P1_DATAO_REG_8_;
  assign new_SUB_1605_U15 = ~P2_DATAO_REG_8_;
  assign new_SUB_1605_U16 = ~P2_DATAO_REG_7_;
  assign new_SUB_1605_U17 = ~P1_DATAO_REG_6_;
  assign new_SUB_1605_U18 = ~P1_DATAO_REG_7_;
  assign new_SUB_1605_U19 = ~P2_DATAO_REG_6_;
  assign new_SUB_1605_U20 = ~P1_DATAO_REG_5_;
  assign new_SUB_1605_U21 = ~new_SUB_1605_U303 | ~new_SUB_1605_U204;
  assign new_SUB_1605_U22 = ~P1_DATAO_REG_4_;
  assign new_SUB_1605_U23 = ~P2_DATAO_REG_0_;
  assign new_SUB_1605_U24 = ~P1_DATAO_REG_1_;
  assign new_SUB_1605_U25 = ~P2_DATAO_REG_4_;
  assign new_SUB_1605_U26 = ~P2_DATAO_REG_2_;
  assign new_SUB_1605_U27 = ~P2_DATAO_REG_3_;
  assign new_SUB_1605_U28 = ~P1_DATAO_REG_2_;
  assign new_SUB_1605_U29 = ~P1_DATAO_REG_3_;
  assign new_SUB_1605_U30 = ~P2_DATAO_REG_5_;
  assign new_SUB_1605_U31 = ~P2_DATAO_REG_9_;
  assign new_SUB_1605_U32 = ~P1_DATAO_REG_9_;
  assign new_SUB_1605_U33 = ~P1_DATAO_REG_12_;
  assign new_SUB_1605_U34 = ~P2_DATAO_REG_12_;
  assign new_SUB_1605_U35 = ~P2_DATAO_REG_11_;
  assign new_SUB_1605_U36 = ~P2_DATAO_REG_10_;
  assign new_SUB_1605_U37 = ~P1_DATAO_REG_11_;
  assign new_SUB_1605_U38 = ~P1_DATAO_REG_10_;
  assign new_SUB_1605_U39 = ~P1_DATAO_REG_9_ | ~new_SUB_1605_U31;
  assign new_SUB_1605_U40 = ~P2_DATAO_REG_13_;
  assign new_SUB_1605_U41 = ~P1_DATAO_REG_13_;
  assign new_SUB_1605_U42 = ~P2_DATAO_REG_14_;
  assign new_SUB_1605_U43 = ~P1_DATAO_REG_14_;
  assign new_SUB_1605_U44 = ~P2_DATAO_REG_15_;
  assign new_SUB_1605_U45 = ~P1_DATAO_REG_15_;
  assign new_SUB_1605_U46 = ~P2_DATAO_REG_16_;
  assign new_SUB_1605_U47 = ~P1_DATAO_REG_16_;
  assign new_SUB_1605_U48 = ~P2_DATAO_REG_17_;
  assign new_SUB_1605_U49 = ~P1_DATAO_REG_17_;
  assign new_SUB_1605_U50 = ~P2_DATAO_REG_18_;
  assign new_SUB_1605_U51 = ~P1_DATAO_REG_18_;
  assign new_SUB_1605_U52 = ~P2_DATAO_REG_19_;
  assign new_SUB_1605_U53 = ~P1_DATAO_REG_19_;
  assign new_SUB_1605_U54 = ~P2_DATAO_REG_20_;
  assign new_SUB_1605_U55 = ~P1_DATAO_REG_20_;
  assign new_SUB_1605_U56 = ~P2_DATAO_REG_21_;
  assign new_SUB_1605_U57 = ~P1_DATAO_REG_21_;
  assign new_SUB_1605_U58 = ~P2_DATAO_REG_22_;
  assign new_SUB_1605_U59 = ~P1_DATAO_REG_22_;
  assign new_SUB_1605_U60 = ~P2_DATAO_REG_23_;
  assign new_SUB_1605_U61 = ~P1_DATAO_REG_23_;
  assign new_SUB_1605_U62 = ~P2_DATAO_REG_24_;
  assign new_SUB_1605_U63 = ~P1_DATAO_REG_24_;
  assign new_SUB_1605_U64 = ~P2_DATAO_REG_25_;
  assign new_SUB_1605_U65 = ~P1_DATAO_REG_25_;
  assign new_SUB_1605_U66 = ~P2_DATAO_REG_26_;
  assign new_SUB_1605_U67 = ~P1_DATAO_REG_26_;
  assign new_SUB_1605_U68 = ~P2_DATAO_REG_27_;
  assign new_SUB_1605_U69 = ~P1_DATAO_REG_27_;
  assign new_SUB_1605_U70 = ~P2_DATAO_REG_28_;
  assign new_SUB_1605_U71 = ~P1_DATAO_REG_28_;
  assign new_SUB_1605_U72 = ~P2_DATAO_REG_29_;
  assign new_SUB_1605_U73 = ~P1_DATAO_REG_29_;
  assign new_SUB_1605_U74 = ~P1_DATAO_REG_30_;
  assign new_SUB_1605_U75 = ~P2_DATAO_REG_30_;
  assign new_SUB_1605_U76 = ~new_SUB_1605_U308 | ~new_SUB_1605_U216;
  assign new_SUB_1605_U77 = ~new_SUB_1605_U305 | ~new_SUB_1605_U213;
  assign new_SUB_1605_U78 = ~P1_DATAO_REG_0_;
  assign new_SUB_1605_U79 = ~new_SUB_1605_U328 | ~new_SUB_1605_U327;
  assign new_SUB_1605_U80 = ~new_SUB_1605_U333 | ~new_SUB_1605_U332;
  assign new_SUB_1605_U81 = ~new_SUB_1605_U338 | ~new_SUB_1605_U337;
  assign new_SUB_1605_U82 = ~new_SUB_1605_U343 | ~new_SUB_1605_U342;
  assign new_SUB_1605_U83 = ~new_SUB_1605_U348 | ~new_SUB_1605_U347;
  assign new_SUB_1605_U84 = ~new_SUB_1605_U353 | ~new_SUB_1605_U352;
  assign new_SUB_1605_U85 = ~new_SUB_1605_U358 | ~new_SUB_1605_U357;
  assign new_SUB_1605_U86 = ~new_SUB_1605_U370 | ~new_SUB_1605_U369;
  assign new_SUB_1605_U87 = ~new_SUB_1605_U375 | ~new_SUB_1605_U374;
  assign new_SUB_1605_U88 = ~new_SUB_1605_U380 | ~new_SUB_1605_U379;
  assign new_SUB_1605_U89 = ~new_SUB_1605_U385 | ~new_SUB_1605_U384;
  assign new_SUB_1605_U90 = ~new_SUB_1605_U390 | ~new_SUB_1605_U389;
  assign new_SUB_1605_U91 = ~new_SUB_1605_U395 | ~new_SUB_1605_U394;
  assign new_SUB_1605_U92 = ~new_SUB_1605_U400 | ~new_SUB_1605_U399;
  assign new_SUB_1605_U93 = ~new_SUB_1605_U405 | ~new_SUB_1605_U404;
  assign new_SUB_1605_U94 = ~new_SUB_1605_U410 | ~new_SUB_1605_U409;
  assign new_SUB_1605_U95 = ~new_SUB_1605_U415 | ~new_SUB_1605_U414;
  assign new_SUB_1605_U96 = ~new_SUB_1605_U420 | ~new_SUB_1605_U419;
  assign new_SUB_1605_U97 = ~new_SUB_1605_U425 | ~new_SUB_1605_U424;
  assign new_SUB_1605_U98 = ~new_SUB_1605_U430 | ~new_SUB_1605_U429;
  assign new_SUB_1605_U99 = ~new_SUB_1605_U435 | ~new_SUB_1605_U434;
  assign new_SUB_1605_U100 = ~new_SUB_1605_U440 | ~new_SUB_1605_U439;
  assign new_SUB_1605_U101 = ~new_SUB_1605_U445 | ~new_SUB_1605_U444;
  assign new_SUB_1605_U102 = ~new_SUB_1605_U450 | ~new_SUB_1605_U449;
  assign new_SUB_1605_U103 = ~new_SUB_1605_U455 | ~new_SUB_1605_U454;
  assign new_SUB_1605_U104 = ~new_SUB_1605_U460 | ~new_SUB_1605_U459;
  assign new_SUB_1605_U105 = ~new_SUB_1605_U465 | ~new_SUB_1605_U464;
  assign new_SUB_1605_U106 = ~new_SUB_1605_U470 | ~new_SUB_1605_U469;
  assign new_SUB_1605_U107 = ~new_SUB_1605_U475 | ~new_SUB_1605_U474;
  assign new_SUB_1605_U108 = ~new_SUB_1605_U480 | ~new_SUB_1605_U479;
  assign new_SUB_1605_U109 = P1_DATAO_REG_5_ & new_SUB_1605_U30;
  assign new_SUB_1605_U110 = new_SUB_1605_U205 & new_SUB_1605_U203;
  assign new_SUB_1605_U111 = new_SUB_1605_U197 & new_SUB_1605_U6;
  assign new_SUB_1605_U112 = new_SUB_1605_U299 & new_SUB_1605_U197;
  assign new_SUB_1605_U113 = new_SUB_1605_U298 & new_SUB_1605_U198;
  assign new_SUB_1605_U114 = new_SUB_1605_U206 & new_SUB_1605_U8;
  assign new_SUB_1605_U115 = new_SUB_1605_U302 & new_SUB_1605_U207;
  assign new_SUB_1605_U116 = ~new_SUB_1605_U325 | ~new_SUB_1605_U324;
  assign new_SUB_1605_U117 = ~new_SUB_1605_U330 | ~new_SUB_1605_U329;
  assign new_SUB_1605_U118 = new_SUB_1605_U300 & new_SUB_1605_U203;
  assign new_SUB_1605_U119 = ~new_SUB_1605_U335 | ~new_SUB_1605_U334;
  assign new_SUB_1605_U120 = ~new_SUB_1605_U340 | ~new_SUB_1605_U339;
  assign new_SUB_1605_U121 = ~new_SUB_1605_U345 | ~new_SUB_1605_U344;
  assign new_SUB_1605_U122 = ~new_SUB_1605_U350 | ~new_SUB_1605_U349;
  assign new_SUB_1605_U123 = ~new_SUB_1605_U355 | ~new_SUB_1605_U354;
  assign new_SUB_1605_U124 = new_SUB_1605_U10 & new_SUB_1605_U218;
  assign new_SUB_1605_U125 = new_SUB_1605_U311 & new_SUB_1605_U219;
  assign new_SUB_1605_U126 = new_SUB_1605_U287 & new_SUB_1605_U11 & new_SUB_1605_U290;
  assign new_SUB_1605_U127 = new_SUB_1605_U289 & new_SUB_1605_U361;
  assign new_SUB_1605_U128 = new_SUB_1605_U161 & new_SUB_1605_U293;
  assign new_SUB_1605_U129 = ~new_SUB_1605_U367 | ~new_SUB_1605_U366;
  assign new_SUB_1605_U130 = ~new_SUB_1605_U372 | ~new_SUB_1605_U371;
  assign new_SUB_1605_U131 = ~new_SUB_1605_U377 | ~new_SUB_1605_U376;
  assign new_SUB_1605_U132 = ~new_SUB_1605_U382 | ~new_SUB_1605_U381;
  assign new_SUB_1605_U133 = ~new_SUB_1605_U387 | ~new_SUB_1605_U386;
  assign new_SUB_1605_U134 = ~new_SUB_1605_U392 | ~new_SUB_1605_U391;
  assign new_SUB_1605_U135 = ~new_SUB_1605_U397 | ~new_SUB_1605_U396;
  assign new_SUB_1605_U136 = ~new_SUB_1605_U402 | ~new_SUB_1605_U401;
  assign new_SUB_1605_U137 = ~new_SUB_1605_U407 | ~new_SUB_1605_U406;
  assign new_SUB_1605_U138 = ~new_SUB_1605_U412 | ~new_SUB_1605_U411;
  assign new_SUB_1605_U139 = ~new_SUB_1605_U417 | ~new_SUB_1605_U416;
  assign new_SUB_1605_U140 = ~new_SUB_1605_U422 | ~new_SUB_1605_U421;
  assign new_SUB_1605_U141 = ~new_SUB_1605_U427 | ~new_SUB_1605_U426;
  assign new_SUB_1605_U142 = ~new_SUB_1605_U432 | ~new_SUB_1605_U431;
  assign new_SUB_1605_U143 = ~new_SUB_1605_U437 | ~new_SUB_1605_U436;
  assign new_SUB_1605_U144 = ~new_SUB_1605_U442 | ~new_SUB_1605_U441;
  assign new_SUB_1605_U145 = ~new_SUB_1605_U447 | ~new_SUB_1605_U446;
  assign new_SUB_1605_U146 = ~new_SUB_1605_U452 | ~new_SUB_1605_U451;
  assign new_SUB_1605_U147 = ~new_SUB_1605_U457 | ~new_SUB_1605_U456;
  assign new_SUB_1605_U148 = ~new_SUB_1605_U462 | ~new_SUB_1605_U461;
  assign new_SUB_1605_U149 = ~new_SUB_1605_U467 | ~new_SUB_1605_U466;
  assign new_SUB_1605_U150 = ~new_SUB_1605_U472 | ~new_SUB_1605_U471;
  assign new_SUB_1605_U151 = ~new_SUB_1605_U477 | ~new_SUB_1605_U476;
  assign new_SUB_1605_U152 = ~new_SUB_1605_U115 | ~new_SUB_1605_U321;
  assign new_SUB_1605_U153 = ~new_SUB_1605_U319 | ~new_SUB_1605_U21;
  assign new_SUB_1605_U154 = ~new_SUB_1605_U118 | ~new_SUB_1605_U317;
  assign new_SUB_1605_U155 = ~new_SUB_1605_U315 | ~new_SUB_1605_U201;
  assign new_SUB_1605_U156 = ~new_SUB_1605_U113 | ~new_SUB_1605_U297;
  assign new_SUB_1605_U157 = ~new_SUB_1605_U296 | ~new_SUB_1605_U294;
  assign new_SUB_1605_U158 = ~new_SUB_1605_U192 | ~new_SUB_1605_U191;
  assign new_SUB_1605_U159 = ~P2_DATAO_REG_31_;
  assign new_SUB_1605_U160 = ~P1_DATAO_REG_31_;
  assign new_SUB_1605_U161 = new_SUB_1605_U365 & new_SUB_1605_U364;
  assign new_SUB_1605_U162 = ~new_SUB_1605_U287 | ~new_SUB_1605_U286;
  assign new_SUB_1605_U163 = ~new_SUB_1605_U292 | ~new_SUB_1605_U188 | ~new_SUB_1605_U186;
  assign new_SUB_1605_U164 = ~new_SUB_1605_U283 | ~new_SUB_1605_U282;
  assign new_SUB_1605_U165 = ~new_SUB_1605_U279 | ~new_SUB_1605_U278;
  assign new_SUB_1605_U166 = ~new_SUB_1605_U275 | ~new_SUB_1605_U274;
  assign new_SUB_1605_U167 = ~new_SUB_1605_U271 | ~new_SUB_1605_U270;
  assign new_SUB_1605_U168 = ~new_SUB_1605_U267 | ~new_SUB_1605_U266;
  assign new_SUB_1605_U169 = ~new_SUB_1605_U263 | ~new_SUB_1605_U262;
  assign new_SUB_1605_U170 = ~new_SUB_1605_U259 | ~new_SUB_1605_U258;
  assign new_SUB_1605_U171 = ~new_SUB_1605_U255 | ~new_SUB_1605_U254;
  assign new_SUB_1605_U172 = ~new_SUB_1605_U251 | ~new_SUB_1605_U250;
  assign new_SUB_1605_U173 = ~new_SUB_1605_U247 | ~new_SUB_1605_U246;
  assign new_SUB_1605_U174 = ~P2_DATAO_REG_1_;
  assign new_SUB_1605_U175 = ~P2_DATAO_REG_0_ | ~new_SUB_1605_U78;
  assign new_SUB_1605_U176 = ~new_SUB_1605_U243 | ~new_SUB_1605_U242;
  assign new_SUB_1605_U177 = ~new_SUB_1605_U239 | ~new_SUB_1605_U238;
  assign new_SUB_1605_U178 = ~new_SUB_1605_U235 | ~new_SUB_1605_U234;
  assign new_SUB_1605_U179 = ~new_SUB_1605_U231 | ~new_SUB_1605_U230;
  assign new_SUB_1605_U180 = ~new_SUB_1605_U227 | ~new_SUB_1605_U226;
  assign new_SUB_1605_U181 = ~new_SUB_1605_U223 | ~new_SUB_1605_U222;
  assign new_SUB_1605_U182 = ~new_SUB_1605_U125 | ~new_SUB_1605_U310;
  assign new_SUB_1605_U183 = ~new_SUB_1605_U309 | ~new_SUB_1605_U307;
  assign new_SUB_1605_U184 = ~new_SUB_1605_U306 | ~new_SUB_1605_U304;
  assign new_SUB_1605_U185 = ~new_SUB_1605_U39 | ~new_SUB_1605_U209;
  assign new_SUB_1605_U186 = ~new_SUB_1605_U175 | ~new_SUB_1605_U174;
  assign new_SUB_1605_U187 = ~new_SUB_1605_U175;
  assign new_SUB_1605_U188 = ~P1_DATAO_REG_1_ | ~new_SUB_1605_U175;
  assign new_SUB_1605_U189 = ~new_SUB_1605_U163;
  assign new_SUB_1605_U190 = ~P2_DATAO_REG_2_ | ~new_SUB_1605_U28;
  assign new_SUB_1605_U191 = ~new_SUB_1605_U190 | ~new_SUB_1605_U312;
  assign new_SUB_1605_U192 = ~P1_DATAO_REG_2_ | ~new_SUB_1605_U26;
  assign new_SUB_1605_U193 = ~new_SUB_1605_U158;
  assign new_SUB_1605_U194 = ~P2_DATAO_REG_3_ | ~new_SUB_1605_U29;
  assign new_SUB_1605_U195 = ~P1_DATAO_REG_3_ | ~new_SUB_1605_U27;
  assign new_SUB_1605_U196 = ~new_SUB_1605_U157;
  assign new_SUB_1605_U197 = ~P2_DATAO_REG_4_ | ~new_SUB_1605_U22;
  assign new_SUB_1605_U198 = ~P1_DATAO_REG_4_ | ~new_SUB_1605_U25;
  assign new_SUB_1605_U199 = ~new_SUB_1605_U156;
  assign new_SUB_1605_U200 = ~P2_DATAO_REG_5_ | ~new_SUB_1605_U20;
  assign new_SUB_1605_U201 = ~P1_DATAO_REG_5_ | ~new_SUB_1605_U30;
  assign new_SUB_1605_U202 = ~P2_DATAO_REG_6_ | ~new_SUB_1605_U17;
  assign new_SUB_1605_U203 = ~P1_DATAO_REG_6_ | ~new_SUB_1605_U19;
  assign new_SUB_1605_U204 = ~P2_DATAO_REG_7_ | ~new_SUB_1605_U18;
  assign new_SUB_1605_U205 = ~P1_DATAO_REG_7_ | ~new_SUB_1605_U16;
  assign new_SUB_1605_U206 = ~P2_DATAO_REG_8_ | ~new_SUB_1605_U14;
  assign new_SUB_1605_U207 = ~P1_DATAO_REG_8_ | ~new_SUB_1605_U15;
  assign new_SUB_1605_U208 = ~P2_DATAO_REG_9_ | ~new_SUB_1605_U32;
  assign new_SUB_1605_U209 = ~new_SUB_1605_U208 | ~new_SUB_1605_U152;
  assign new_SUB_1605_U210 = ~new_SUB_1605_U39;
  assign new_SUB_1605_U211 = ~new_SUB_1605_U185;
  assign new_SUB_1605_U212 = ~P2_DATAO_REG_10_ | ~new_SUB_1605_U38;
  assign new_SUB_1605_U213 = ~P1_DATAO_REG_10_ | ~new_SUB_1605_U36;
  assign new_SUB_1605_U214 = ~new_SUB_1605_U184;
  assign new_SUB_1605_U215 = ~P2_DATAO_REG_11_ | ~new_SUB_1605_U37;
  assign new_SUB_1605_U216 = ~P1_DATAO_REG_11_ | ~new_SUB_1605_U35;
  assign new_SUB_1605_U217 = ~new_SUB_1605_U183;
  assign new_SUB_1605_U218 = ~P2_DATAO_REG_12_ | ~new_SUB_1605_U33;
  assign new_SUB_1605_U219 = ~P1_DATAO_REG_12_ | ~new_SUB_1605_U34;
  assign new_SUB_1605_U220 = ~new_SUB_1605_U182;
  assign new_SUB_1605_U221 = ~P2_DATAO_REG_13_ | ~new_SUB_1605_U41;
  assign new_SUB_1605_U222 = ~new_SUB_1605_U221 | ~new_SUB_1605_U182;
  assign new_SUB_1605_U223 = ~P1_DATAO_REG_13_ | ~new_SUB_1605_U40;
  assign new_SUB_1605_U224 = ~new_SUB_1605_U181;
  assign new_SUB_1605_U225 = ~P2_DATAO_REG_14_ | ~new_SUB_1605_U43;
  assign new_SUB_1605_U226 = ~new_SUB_1605_U225 | ~new_SUB_1605_U181;
  assign new_SUB_1605_U227 = ~P1_DATAO_REG_14_ | ~new_SUB_1605_U42;
  assign new_SUB_1605_U228 = ~new_SUB_1605_U180;
  assign new_SUB_1605_U229 = ~P2_DATAO_REG_15_ | ~new_SUB_1605_U45;
  assign new_SUB_1605_U230 = ~new_SUB_1605_U229 | ~new_SUB_1605_U180;
  assign new_SUB_1605_U231 = ~P1_DATAO_REG_15_ | ~new_SUB_1605_U44;
  assign new_SUB_1605_U232 = ~new_SUB_1605_U179;
  assign new_SUB_1605_U233 = ~P2_DATAO_REG_16_ | ~new_SUB_1605_U47;
  assign new_SUB_1605_U234 = ~new_SUB_1605_U233 | ~new_SUB_1605_U179;
  assign new_SUB_1605_U235 = ~P1_DATAO_REG_16_ | ~new_SUB_1605_U46;
  assign new_SUB_1605_U236 = ~new_SUB_1605_U178;
  assign new_SUB_1605_U237 = ~P2_DATAO_REG_17_ | ~new_SUB_1605_U49;
  assign new_SUB_1605_U238 = ~new_SUB_1605_U237 | ~new_SUB_1605_U178;
  assign new_SUB_1605_U239 = ~P1_DATAO_REG_17_ | ~new_SUB_1605_U48;
  assign new_SUB_1605_U240 = ~new_SUB_1605_U177;
  assign new_SUB_1605_U241 = ~P2_DATAO_REG_18_ | ~new_SUB_1605_U51;
  assign new_SUB_1605_U242 = ~new_SUB_1605_U241 | ~new_SUB_1605_U177;
  assign new_SUB_1605_U243 = ~P1_DATAO_REG_18_ | ~new_SUB_1605_U50;
  assign new_SUB_1605_U244 = ~new_SUB_1605_U176;
  assign new_SUB_1605_U245 = ~P2_DATAO_REG_19_ | ~new_SUB_1605_U53;
  assign new_SUB_1605_U246 = ~new_SUB_1605_U245 | ~new_SUB_1605_U176;
  assign new_SUB_1605_U247 = ~P1_DATAO_REG_19_ | ~new_SUB_1605_U52;
  assign new_SUB_1605_U248 = ~new_SUB_1605_U173;
  assign new_SUB_1605_U249 = ~P2_DATAO_REG_20_ | ~new_SUB_1605_U55;
  assign new_SUB_1605_U250 = ~new_SUB_1605_U249 | ~new_SUB_1605_U173;
  assign new_SUB_1605_U251 = ~P1_DATAO_REG_20_ | ~new_SUB_1605_U54;
  assign new_SUB_1605_U252 = ~new_SUB_1605_U172;
  assign new_SUB_1605_U253 = ~P2_DATAO_REG_21_ | ~new_SUB_1605_U57;
  assign new_SUB_1605_U254 = ~new_SUB_1605_U253 | ~new_SUB_1605_U172;
  assign new_SUB_1605_U255 = ~P1_DATAO_REG_21_ | ~new_SUB_1605_U56;
  assign new_SUB_1605_U256 = ~new_SUB_1605_U171;
  assign new_SUB_1605_U257 = ~P2_DATAO_REG_22_ | ~new_SUB_1605_U59;
  assign new_SUB_1605_U258 = ~new_SUB_1605_U257 | ~new_SUB_1605_U171;
  assign new_SUB_1605_U259 = ~P1_DATAO_REG_22_ | ~new_SUB_1605_U58;
  assign new_SUB_1605_U260 = ~new_SUB_1605_U170;
  assign new_SUB_1605_U261 = ~P2_DATAO_REG_23_ | ~new_SUB_1605_U61;
  assign new_SUB_1605_U262 = ~new_SUB_1605_U261 | ~new_SUB_1605_U170;
  assign new_SUB_1605_U263 = ~P1_DATAO_REG_23_ | ~new_SUB_1605_U60;
  assign new_SUB_1605_U264 = ~new_SUB_1605_U169;
  assign new_SUB_1605_U265 = ~P2_DATAO_REG_24_ | ~new_SUB_1605_U63;
  assign new_SUB_1605_U266 = ~new_SUB_1605_U265 | ~new_SUB_1605_U169;
  assign new_SUB_1605_U267 = ~P1_DATAO_REG_24_ | ~new_SUB_1605_U62;
  assign new_SUB_1605_U268 = ~new_SUB_1605_U168;
  assign new_SUB_1605_U269 = ~P2_DATAO_REG_25_ | ~new_SUB_1605_U65;
  assign new_SUB_1605_U270 = ~new_SUB_1605_U269 | ~new_SUB_1605_U168;
  assign new_SUB_1605_U271 = ~P1_DATAO_REG_25_ | ~new_SUB_1605_U64;
  assign new_SUB_1605_U272 = ~new_SUB_1605_U167;
  assign new_SUB_1605_U273 = ~P2_DATAO_REG_26_ | ~new_SUB_1605_U67;
  assign new_SUB_1605_U274 = ~new_SUB_1605_U273 | ~new_SUB_1605_U167;
  assign new_SUB_1605_U275 = ~P1_DATAO_REG_26_ | ~new_SUB_1605_U66;
  assign new_SUB_1605_U276 = ~new_SUB_1605_U166;
  assign new_SUB_1605_U277 = ~P2_DATAO_REG_27_ | ~new_SUB_1605_U69;
  assign new_SUB_1605_U278 = ~new_SUB_1605_U277 | ~new_SUB_1605_U166;
  assign new_SUB_1605_U279 = ~P1_DATAO_REG_27_ | ~new_SUB_1605_U68;
  assign new_SUB_1605_U280 = ~new_SUB_1605_U165;
  assign new_SUB_1605_U281 = ~P2_DATAO_REG_28_ | ~new_SUB_1605_U71;
  assign new_SUB_1605_U282 = ~new_SUB_1605_U281 | ~new_SUB_1605_U165;
  assign new_SUB_1605_U283 = ~P1_DATAO_REG_28_ | ~new_SUB_1605_U70;
  assign new_SUB_1605_U284 = ~new_SUB_1605_U164;
  assign new_SUB_1605_U285 = ~P2_DATAO_REG_29_ | ~new_SUB_1605_U73;
  assign new_SUB_1605_U286 = ~new_SUB_1605_U285 | ~new_SUB_1605_U164;
  assign new_SUB_1605_U287 = ~P1_DATAO_REG_29_ | ~new_SUB_1605_U72;
  assign new_SUB_1605_U288 = ~new_SUB_1605_U162;
  assign new_SUB_1605_U289 = ~P2_DATAO_REG_30_ | ~new_SUB_1605_U74;
  assign new_SUB_1605_U290 = ~P1_DATAO_REG_30_ | ~new_SUB_1605_U75;
  assign new_SUB_1605_U291 = ~P1_DATAO_REG_0_ | ~new_SUB_1605_U23;
  assign new_SUB_1605_U292 = ~P1_DATAO_REG_1_ | ~new_SUB_1605_U174;
  assign new_SUB_1605_U293 = ~new_SUB_1605_U286 | ~new_SUB_1605_U126;
  assign new_SUB_1605_U294 = ~new_SUB_1605_U6 | ~new_SUB_1605_U163;
  assign new_SUB_1605_U295 = ~new_SUB_1605_U195 | ~new_SUB_1605_U192;
  assign new_SUB_1605_U296 = ~new_SUB_1605_U295 | ~new_SUB_1605_U299;
  assign new_SUB_1605_U297 = ~new_SUB_1605_U111 | ~new_SUB_1605_U163;
  assign new_SUB_1605_U298 = ~new_SUB_1605_U112 | ~new_SUB_1605_U295;
  assign new_SUB_1605_U299 = ~P2_DATAO_REG_3_ | ~new_SUB_1605_U29;
  assign new_SUB_1605_U300 = ~new_SUB_1605_U109 | ~new_SUB_1605_U202;
  assign new_SUB_1605_U301 = ~new_SUB_1605_U21;
  assign new_SUB_1605_U302 = ~new_SUB_1605_U301 | ~new_SUB_1605_U206;
  assign new_SUB_1605_U303 = ~new_SUB_1605_U110 | ~new_SUB_1605_U300;
  assign new_SUB_1605_U304 = ~new_SUB_1605_U9 | ~new_SUB_1605_U152;
  assign new_SUB_1605_U305 = ~new_SUB_1605_U210 | ~new_SUB_1605_U212;
  assign new_SUB_1605_U306 = ~new_SUB_1605_U77;
  assign new_SUB_1605_U307 = ~new_SUB_1605_U10 | ~new_SUB_1605_U152;
  assign new_SUB_1605_U308 = ~new_SUB_1605_U77 | ~new_SUB_1605_U215;
  assign new_SUB_1605_U309 = ~new_SUB_1605_U76;
  assign new_SUB_1605_U310 = ~new_SUB_1605_U124 | ~new_SUB_1605_U152;
  assign new_SUB_1605_U311 = ~new_SUB_1605_U76 | ~new_SUB_1605_U218;
  assign new_SUB_1605_U312 = ~new_SUB_1605_U314 | ~new_SUB_1605_U313 | ~new_SUB_1605_U292;
  assign new_SUB_1605_U313 = ~P1_DATAO_REG_1_ | ~new_SUB_1605_U175;
  assign new_SUB_1605_U314 = ~new_SUB_1605_U175 | ~new_SUB_1605_U174;
  assign new_SUB_1605_U315 = ~new_SUB_1605_U200 | ~new_SUB_1605_U156;
  assign new_SUB_1605_U316 = ~new_SUB_1605_U155;
  assign new_SUB_1605_U317 = ~new_SUB_1605_U7 | ~new_SUB_1605_U156;
  assign new_SUB_1605_U318 = ~new_SUB_1605_U154;
  assign new_SUB_1605_U319 = ~new_SUB_1605_U8 | ~new_SUB_1605_U156;
  assign new_SUB_1605_U320 = ~new_SUB_1605_U153;
  assign new_SUB_1605_U321 = ~new_SUB_1605_U114 | ~new_SUB_1605_U156;
  assign new_SUB_1605_U322 = ~new_SUB_1605_U152;
  assign new_SUB_1605_U323 = ~new_SUB_1605_U127 | ~new_SUB_1605_U162;
  assign new_SUB_1605_U324 = ~P2_DATAO_REG_9_ | ~new_SUB_1605_U32;
  assign new_SUB_1605_U325 = ~P1_DATAO_REG_9_ | ~new_SUB_1605_U31;
  assign new_SUB_1605_U326 = ~new_SUB_1605_U116;
  assign new_SUB_1605_U327 = ~new_SUB_1605_U322 | ~new_SUB_1605_U326;
  assign new_SUB_1605_U328 = ~new_SUB_1605_U116 | ~new_SUB_1605_U152;
  assign new_SUB_1605_U329 = ~P2_DATAO_REG_8_ | ~new_SUB_1605_U14;
  assign new_SUB_1605_U330 = ~P1_DATAO_REG_8_ | ~new_SUB_1605_U15;
  assign new_SUB_1605_U331 = ~new_SUB_1605_U117;
  assign new_SUB_1605_U332 = ~new_SUB_1605_U320 | ~new_SUB_1605_U331;
  assign new_SUB_1605_U333 = ~new_SUB_1605_U117 | ~new_SUB_1605_U153;
  assign new_SUB_1605_U334 = ~P2_DATAO_REG_7_ | ~new_SUB_1605_U18;
  assign new_SUB_1605_U335 = ~P1_DATAO_REG_7_ | ~new_SUB_1605_U16;
  assign new_SUB_1605_U336 = ~new_SUB_1605_U119;
  assign new_SUB_1605_U337 = ~new_SUB_1605_U318 | ~new_SUB_1605_U336;
  assign new_SUB_1605_U338 = ~new_SUB_1605_U119 | ~new_SUB_1605_U154;
  assign new_SUB_1605_U339 = ~P2_DATAO_REG_6_ | ~new_SUB_1605_U17;
  assign new_SUB_1605_U340 = ~P1_DATAO_REG_6_ | ~new_SUB_1605_U19;
  assign new_SUB_1605_U341 = ~new_SUB_1605_U120;
  assign new_SUB_1605_U342 = ~new_SUB_1605_U316 | ~new_SUB_1605_U341;
  assign new_SUB_1605_U343 = ~new_SUB_1605_U120 | ~new_SUB_1605_U155;
  assign new_SUB_1605_U344 = ~P2_DATAO_REG_5_ | ~new_SUB_1605_U20;
  assign new_SUB_1605_U345 = ~P1_DATAO_REG_5_ | ~new_SUB_1605_U30;
  assign new_SUB_1605_U346 = ~new_SUB_1605_U121;
  assign new_SUB_1605_U347 = ~new_SUB_1605_U199 | ~new_SUB_1605_U346;
  assign new_SUB_1605_U348 = ~new_SUB_1605_U121 | ~new_SUB_1605_U156;
  assign new_SUB_1605_U349 = ~P2_DATAO_REG_4_ | ~new_SUB_1605_U22;
  assign new_SUB_1605_U350 = ~P1_DATAO_REG_4_ | ~new_SUB_1605_U25;
  assign new_SUB_1605_U351 = ~new_SUB_1605_U122;
  assign new_SUB_1605_U352 = ~new_SUB_1605_U196 | ~new_SUB_1605_U351;
  assign new_SUB_1605_U353 = ~new_SUB_1605_U122 | ~new_SUB_1605_U157;
  assign new_SUB_1605_U354 = ~P2_DATAO_REG_3_ | ~new_SUB_1605_U29;
  assign new_SUB_1605_U355 = ~P1_DATAO_REG_3_ | ~new_SUB_1605_U27;
  assign new_SUB_1605_U356 = ~new_SUB_1605_U123;
  assign new_SUB_1605_U357 = ~new_SUB_1605_U193 | ~new_SUB_1605_U356;
  assign new_SUB_1605_U358 = ~new_SUB_1605_U123 | ~new_SUB_1605_U158;
  assign new_SUB_1605_U359 = ~P2_DATAO_REG_31_ | ~new_SUB_1605_U160;
  assign new_SUB_1605_U360 = ~P1_DATAO_REG_31_ | ~new_SUB_1605_U159;
  assign new_SUB_1605_U361 = ~new_SUB_1605_U360 | ~new_SUB_1605_U359;
  assign new_SUB_1605_U362 = ~P2_DATAO_REG_31_ | ~new_SUB_1605_U160;
  assign new_SUB_1605_U363 = ~P1_DATAO_REG_31_ | ~new_SUB_1605_U159;
  assign new_SUB_1605_U364 = ~new_SUB_1605_U75 | ~P1_DATAO_REG_30_ | ~new_SUB_1605_U361;
  assign new_SUB_1605_U365 = ~P2_DATAO_REG_30_ | ~new_SUB_1605_U11 | ~new_SUB_1605_U74;
  assign new_SUB_1605_U366 = ~P2_DATAO_REG_30_ | ~new_SUB_1605_U74;
  assign new_SUB_1605_U367 = ~P1_DATAO_REG_30_ | ~new_SUB_1605_U75;
  assign new_SUB_1605_U368 = ~new_SUB_1605_U129;
  assign new_SUB_1605_U369 = ~new_SUB_1605_U288 | ~new_SUB_1605_U368;
  assign new_SUB_1605_U370 = ~new_SUB_1605_U129 | ~new_SUB_1605_U162;
  assign new_SUB_1605_U371 = ~P2_DATAO_REG_2_ | ~new_SUB_1605_U28;
  assign new_SUB_1605_U372 = ~P1_DATAO_REG_2_ | ~new_SUB_1605_U26;
  assign new_SUB_1605_U373 = ~new_SUB_1605_U130;
  assign new_SUB_1605_U374 = ~new_SUB_1605_U189 | ~new_SUB_1605_U373;
  assign new_SUB_1605_U375 = ~new_SUB_1605_U130 | ~new_SUB_1605_U163;
  assign new_SUB_1605_U376 = ~P2_DATAO_REG_29_ | ~new_SUB_1605_U73;
  assign new_SUB_1605_U377 = ~P1_DATAO_REG_29_ | ~new_SUB_1605_U72;
  assign new_SUB_1605_U378 = ~new_SUB_1605_U131;
  assign new_SUB_1605_U379 = ~new_SUB_1605_U284 | ~new_SUB_1605_U378;
  assign new_SUB_1605_U380 = ~new_SUB_1605_U131 | ~new_SUB_1605_U164;
  assign new_SUB_1605_U381 = ~P2_DATAO_REG_28_ | ~new_SUB_1605_U71;
  assign new_SUB_1605_U382 = ~P1_DATAO_REG_28_ | ~new_SUB_1605_U70;
  assign new_SUB_1605_U383 = ~new_SUB_1605_U132;
  assign new_SUB_1605_U384 = ~new_SUB_1605_U280 | ~new_SUB_1605_U383;
  assign new_SUB_1605_U385 = ~new_SUB_1605_U132 | ~new_SUB_1605_U165;
  assign new_SUB_1605_U386 = ~P2_DATAO_REG_27_ | ~new_SUB_1605_U69;
  assign new_SUB_1605_U387 = ~P1_DATAO_REG_27_ | ~new_SUB_1605_U68;
  assign new_SUB_1605_U388 = ~new_SUB_1605_U133;
  assign new_SUB_1605_U389 = ~new_SUB_1605_U276 | ~new_SUB_1605_U388;
  assign new_SUB_1605_U390 = ~new_SUB_1605_U133 | ~new_SUB_1605_U166;
  assign new_SUB_1605_U391 = ~P2_DATAO_REG_26_ | ~new_SUB_1605_U67;
  assign new_SUB_1605_U392 = ~P1_DATAO_REG_26_ | ~new_SUB_1605_U66;
  assign new_SUB_1605_U393 = ~new_SUB_1605_U134;
  assign new_SUB_1605_U394 = ~new_SUB_1605_U272 | ~new_SUB_1605_U393;
  assign new_SUB_1605_U395 = ~new_SUB_1605_U134 | ~new_SUB_1605_U167;
  assign new_SUB_1605_U396 = ~P2_DATAO_REG_25_ | ~new_SUB_1605_U65;
  assign new_SUB_1605_U397 = ~P1_DATAO_REG_25_ | ~new_SUB_1605_U64;
  assign new_SUB_1605_U398 = ~new_SUB_1605_U135;
  assign new_SUB_1605_U399 = ~new_SUB_1605_U268 | ~new_SUB_1605_U398;
  assign new_SUB_1605_U400 = ~new_SUB_1605_U135 | ~new_SUB_1605_U168;
  assign new_SUB_1605_U401 = ~P2_DATAO_REG_24_ | ~new_SUB_1605_U63;
  assign new_SUB_1605_U402 = ~P1_DATAO_REG_24_ | ~new_SUB_1605_U62;
  assign new_SUB_1605_U403 = ~new_SUB_1605_U136;
  assign new_SUB_1605_U404 = ~new_SUB_1605_U264 | ~new_SUB_1605_U403;
  assign new_SUB_1605_U405 = ~new_SUB_1605_U136 | ~new_SUB_1605_U169;
  assign new_SUB_1605_U406 = ~P2_DATAO_REG_23_ | ~new_SUB_1605_U61;
  assign new_SUB_1605_U407 = ~P1_DATAO_REG_23_ | ~new_SUB_1605_U60;
  assign new_SUB_1605_U408 = ~new_SUB_1605_U137;
  assign new_SUB_1605_U409 = ~new_SUB_1605_U260 | ~new_SUB_1605_U408;
  assign new_SUB_1605_U410 = ~new_SUB_1605_U137 | ~new_SUB_1605_U170;
  assign new_SUB_1605_U411 = ~P2_DATAO_REG_22_ | ~new_SUB_1605_U59;
  assign new_SUB_1605_U412 = ~P1_DATAO_REG_22_ | ~new_SUB_1605_U58;
  assign new_SUB_1605_U413 = ~new_SUB_1605_U138;
  assign new_SUB_1605_U414 = ~new_SUB_1605_U256 | ~new_SUB_1605_U413;
  assign new_SUB_1605_U415 = ~new_SUB_1605_U138 | ~new_SUB_1605_U171;
  assign new_SUB_1605_U416 = ~P2_DATAO_REG_21_ | ~new_SUB_1605_U57;
  assign new_SUB_1605_U417 = ~P1_DATAO_REG_21_ | ~new_SUB_1605_U56;
  assign new_SUB_1605_U418 = ~new_SUB_1605_U139;
  assign new_SUB_1605_U419 = ~new_SUB_1605_U252 | ~new_SUB_1605_U418;
  assign new_SUB_1605_U420 = ~new_SUB_1605_U139 | ~new_SUB_1605_U172;
  assign new_SUB_1605_U421 = ~P2_DATAO_REG_20_ | ~new_SUB_1605_U55;
  assign new_SUB_1605_U422 = ~P1_DATAO_REG_20_ | ~new_SUB_1605_U54;
  assign new_SUB_1605_U423 = ~new_SUB_1605_U140;
  assign new_SUB_1605_U424 = ~new_SUB_1605_U248 | ~new_SUB_1605_U423;
  assign new_SUB_1605_U425 = ~new_SUB_1605_U140 | ~new_SUB_1605_U173;
  assign new_SUB_1605_U426 = ~P2_DATAO_REG_1_ | ~new_SUB_1605_U24;
  assign new_SUB_1605_U427 = ~P1_DATAO_REG_1_ | ~new_SUB_1605_U174;
  assign new_SUB_1605_U428 = ~new_SUB_1605_U141;
  assign new_SUB_1605_U429 = ~new_SUB_1605_U187 | ~new_SUB_1605_U428;
  assign new_SUB_1605_U430 = ~new_SUB_1605_U141 | ~new_SUB_1605_U175;
  assign new_SUB_1605_U431 = ~P2_DATAO_REG_19_ | ~new_SUB_1605_U53;
  assign new_SUB_1605_U432 = ~P1_DATAO_REG_19_ | ~new_SUB_1605_U52;
  assign new_SUB_1605_U433 = ~new_SUB_1605_U142;
  assign new_SUB_1605_U434 = ~new_SUB_1605_U244 | ~new_SUB_1605_U433;
  assign new_SUB_1605_U435 = ~new_SUB_1605_U142 | ~new_SUB_1605_U176;
  assign new_SUB_1605_U436 = ~P2_DATAO_REG_18_ | ~new_SUB_1605_U51;
  assign new_SUB_1605_U437 = ~P1_DATAO_REG_18_ | ~new_SUB_1605_U50;
  assign new_SUB_1605_U438 = ~new_SUB_1605_U143;
  assign new_SUB_1605_U439 = ~new_SUB_1605_U240 | ~new_SUB_1605_U438;
  assign new_SUB_1605_U440 = ~new_SUB_1605_U143 | ~new_SUB_1605_U177;
  assign new_SUB_1605_U441 = ~P2_DATAO_REG_17_ | ~new_SUB_1605_U49;
  assign new_SUB_1605_U442 = ~P1_DATAO_REG_17_ | ~new_SUB_1605_U48;
  assign new_SUB_1605_U443 = ~new_SUB_1605_U144;
  assign new_SUB_1605_U444 = ~new_SUB_1605_U236 | ~new_SUB_1605_U443;
  assign new_SUB_1605_U445 = ~new_SUB_1605_U144 | ~new_SUB_1605_U178;
  assign new_SUB_1605_U446 = ~P2_DATAO_REG_16_ | ~new_SUB_1605_U47;
  assign new_SUB_1605_U447 = ~P1_DATAO_REG_16_ | ~new_SUB_1605_U46;
  assign new_SUB_1605_U448 = ~new_SUB_1605_U145;
  assign new_SUB_1605_U449 = ~new_SUB_1605_U232 | ~new_SUB_1605_U448;
  assign new_SUB_1605_U450 = ~new_SUB_1605_U145 | ~new_SUB_1605_U179;
  assign new_SUB_1605_U451 = ~P2_DATAO_REG_15_ | ~new_SUB_1605_U45;
  assign new_SUB_1605_U452 = ~P1_DATAO_REG_15_ | ~new_SUB_1605_U44;
  assign new_SUB_1605_U453 = ~new_SUB_1605_U146;
  assign new_SUB_1605_U454 = ~new_SUB_1605_U228 | ~new_SUB_1605_U453;
  assign new_SUB_1605_U455 = ~new_SUB_1605_U146 | ~new_SUB_1605_U180;
  assign new_SUB_1605_U456 = ~P2_DATAO_REG_14_ | ~new_SUB_1605_U43;
  assign new_SUB_1605_U457 = ~P1_DATAO_REG_14_ | ~new_SUB_1605_U42;
  assign new_SUB_1605_U458 = ~new_SUB_1605_U147;
  assign new_SUB_1605_U459 = ~new_SUB_1605_U224 | ~new_SUB_1605_U458;
  assign new_SUB_1605_U460 = ~new_SUB_1605_U147 | ~new_SUB_1605_U181;
  assign new_SUB_1605_U461 = ~P2_DATAO_REG_13_ | ~new_SUB_1605_U41;
  assign new_SUB_1605_U462 = ~P1_DATAO_REG_13_ | ~new_SUB_1605_U40;
  assign new_SUB_1605_U463 = ~new_SUB_1605_U148;
  assign new_SUB_1605_U464 = ~new_SUB_1605_U220 | ~new_SUB_1605_U463;
  assign new_SUB_1605_U465 = ~new_SUB_1605_U148 | ~new_SUB_1605_U182;
  assign new_SUB_1605_U466 = ~P2_DATAO_REG_12_ | ~new_SUB_1605_U33;
  assign new_SUB_1605_U467 = ~P1_DATAO_REG_12_ | ~new_SUB_1605_U34;
  assign new_SUB_1605_U468 = ~new_SUB_1605_U149;
  assign new_SUB_1605_U469 = ~new_SUB_1605_U217 | ~new_SUB_1605_U468;
  assign new_SUB_1605_U470 = ~new_SUB_1605_U149 | ~new_SUB_1605_U183;
  assign new_SUB_1605_U471 = ~P2_DATAO_REG_11_ | ~new_SUB_1605_U37;
  assign new_SUB_1605_U472 = ~P1_DATAO_REG_11_ | ~new_SUB_1605_U35;
  assign new_SUB_1605_U473 = ~new_SUB_1605_U150;
  assign new_SUB_1605_U474 = ~new_SUB_1605_U214 | ~new_SUB_1605_U473;
  assign new_SUB_1605_U475 = ~new_SUB_1605_U150 | ~new_SUB_1605_U184;
  assign new_SUB_1605_U476 = ~P2_DATAO_REG_10_ | ~new_SUB_1605_U38;
  assign new_SUB_1605_U477 = ~P1_DATAO_REG_10_ | ~new_SUB_1605_U36;
  assign new_SUB_1605_U478 = ~new_SUB_1605_U151;
  assign new_SUB_1605_U479 = ~new_SUB_1605_U211 | ~new_SUB_1605_U478;
  assign new_SUB_1605_U480 = ~new_SUB_1605_U151 | ~new_SUB_1605_U185;
  assign new_R152_U4 = new_R152_U206 & new_R152_U202;
  assign new_R152_U5 = new_R152_U214 & new_R152_U212;
  assign new_R152_U6 = new_R152_U5 & new_R152_U216;
  assign new_R152_U7 = new_R152_U222 & new_R152_U220;
  assign new_R152_U8 = new_R152_U7 & new_R152_U224;
  assign new_R152_U9 = new_R152_U8 & new_R152_U226;
  assign new_R152_U10 = new_R152_U199 & new_R152_U196;
  assign new_R152_U11 = new_R152_U391 & new_R152_U390;
  assign new_R152_U12 = new_R152_U128 & new_R152_U193;
  assign new_R152_U13 = ~new_R152_U172 | ~new_R152_U337;
  assign new_R152_U14 = ~SI_8_;
  assign new_R152_U15 = ~new_U127;
  assign new_R152_U16 = ~SI_7_;
  assign new_R152_U17 = ~new_U128;
  assign new_R152_U18 = ~new_U128 | ~SI_7_;
  assign new_R152_U19 = ~SI_6_;
  assign new_R152_U20 = ~new_U129;
  assign new_R152_U21 = ~SI_3_;
  assign new_R152_U22 = ~new_U134;
  assign new_R152_U23 = ~SI_1_;
  assign new_R152_U24 = ~SI_0_;
  assign new_R152_U25 = ~new_U157;
  assign new_R152_U26 = ~new_U156;
  assign new_R152_U27 = ~SI_2_;
  assign new_R152_U28 = ~new_U145;
  assign new_R152_U29 = ~new_U145 | ~SI_2_;
  assign new_R152_U30 = ~SI_5_;
  assign new_R152_U31 = ~new_U130;
  assign new_R152_U32 = ~SI_4_;
  assign new_R152_U33 = ~new_U131;
  assign new_R152_U34 = ~new_U131 | ~SI_4_;
  assign new_R152_U35 = ~new_U126;
  assign new_R152_U36 = ~SI_9_;
  assign new_R152_U37 = ~new_R152_U294 | ~new_R152_U207;
  assign new_R152_U38 = ~SI_15_;
  assign new_R152_U39 = ~new_U150;
  assign new_R152_U40 = ~SI_14_;
  assign new_R152_U41 = ~new_U151;
  assign new_R152_U42 = ~SI_13_;
  assign new_R152_U43 = ~new_U152;
  assign new_R152_U44 = ~SI_12_;
  assign new_R152_U45 = ~new_U153;
  assign new_R152_U46 = ~SI_11_;
  assign new_R152_U47 = ~new_U154;
  assign new_R152_U48 = ~new_U154 | ~SI_11_;
  assign new_R152_U49 = ~SI_10_;
  assign new_R152_U50 = ~new_U155;
  assign new_R152_U51 = ~SI_16_;
  assign new_R152_U52 = ~new_U149;
  assign new_R152_U53 = ~SI_17_;
  assign new_R152_U54 = ~new_U148;
  assign new_R152_U55 = ~SI_18_;
  assign new_R152_U56 = ~new_U147;
  assign new_R152_U57 = ~SI_19_;
  assign new_R152_U58 = ~new_U146;
  assign new_R152_U59 = ~SI_20_;
  assign new_R152_U60 = ~new_U144;
  assign new_R152_U61 = ~SI_21_;
  assign new_R152_U62 = ~new_U143;
  assign new_R152_U63 = ~SI_22_;
  assign new_R152_U64 = ~new_U142;
  assign new_R152_U65 = ~SI_23_;
  assign new_R152_U66 = ~new_U141;
  assign new_R152_U67 = ~SI_24_;
  assign new_R152_U68 = ~new_U140;
  assign new_R152_U69 = ~SI_25_;
  assign new_R152_U70 = ~new_U139;
  assign new_R152_U71 = ~SI_26_;
  assign new_R152_U72 = ~new_U138;
  assign new_R152_U73 = ~SI_27_;
  assign new_R152_U74 = ~new_U137;
  assign new_R152_U75 = ~SI_28_;
  assign new_R152_U76 = ~new_U136;
  assign new_R152_U77 = ~SI_29_;
  assign new_R152_U78 = ~new_U135;
  assign new_R152_U79 = ~SI_30_;
  assign new_R152_U80 = ~new_U133;
  assign new_R152_U81 = ~new_R152_U307 | ~new_R152_U227;
  assign new_R152_U82 = ~new_R152_U305 | ~new_R152_U225;
  assign new_R152_U83 = ~new_R152_U300 | ~new_R152_U217;
  assign new_R152_U84 = ~new_R152_U554 | ~new_R152_U553;
  assign new_R152_U85 = ~new_R152_U344 | ~new_R152_U343;
  assign new_R152_U86 = ~new_R152_U351 | ~new_R152_U350;
  assign new_R152_U87 = ~new_R152_U358 | ~new_R152_U357;
  assign new_R152_U88 = ~new_R152_U365 | ~new_R152_U364;
  assign new_R152_U89 = ~new_R152_U372 | ~new_R152_U371;
  assign new_R152_U90 = ~new_R152_U379 | ~new_R152_U378;
  assign new_R152_U91 = ~new_R152_U386 | ~new_R152_U385;
  assign new_R152_U92 = ~new_R152_U400 | ~new_R152_U399;
  assign new_R152_U93 = ~new_R152_U407 | ~new_R152_U406;
  assign new_R152_U94 = ~new_R152_U414 | ~new_R152_U413;
  assign new_R152_U95 = ~new_R152_U421 | ~new_R152_U420;
  assign new_R152_U96 = ~new_R152_U428 | ~new_R152_U427;
  assign new_R152_U97 = ~new_R152_U435 | ~new_R152_U434;
  assign new_R152_U98 = ~new_R152_U442 | ~new_R152_U441;
  assign new_R152_U99 = ~new_R152_U449 | ~new_R152_U448;
  assign new_R152_U100 = ~new_R152_U456 | ~new_R152_U455;
  assign new_R152_U101 = ~new_R152_U463 | ~new_R152_U462;
  assign new_R152_U102 = ~new_R152_U470 | ~new_R152_U469;
  assign new_R152_U103 = ~new_R152_U477 | ~new_R152_U476;
  assign new_R152_U104 = ~new_R152_U489 | ~new_R152_U488;
  assign new_R152_U105 = ~new_R152_U496 | ~new_R152_U495;
  assign new_R152_U106 = ~new_R152_U503 | ~new_R152_U502;
  assign new_R152_U107 = ~new_R152_U510 | ~new_R152_U509;
  assign new_R152_U108 = ~new_R152_U517 | ~new_R152_U516;
  assign new_R152_U109 = ~new_R152_U524 | ~new_R152_U523;
  assign new_R152_U110 = ~new_R152_U531 | ~new_R152_U530;
  assign new_R152_U111 = ~new_R152_U538 | ~new_R152_U537;
  assign new_R152_U112 = ~new_R152_U545 | ~new_R152_U544;
  assign new_R152_U113 = ~new_R152_U552 | ~new_R152_U551;
  assign new_R152_U114 = new_R152_U292 & new_R152_U200;
  assign new_R152_U115 = new_R152_U209 & new_R152_U4;
  assign new_R152_U116 = new_R152_U297 & new_R152_U210;
  assign new_R152_U117 = new_R152_U298 & new_R152_U215;
  assign new_R152_U118 = new_R152_U292 & new_R152_U200;
  assign new_R152_U119 = new_U156 & new_U157;
  assign new_R152_U120 = new_U157 & SI_0_;
  assign new_R152_U121 = SI_1_ & new_U156;
  assign new_R152_U122 = new_R152_U218 & new_R152_U6;
  assign new_R152_U123 = new_R152_U302 & new_R152_U219;
  assign new_R152_U124 = new_R152_U9 & new_R152_U228;
  assign new_R152_U125 = new_R152_U309 & new_R152_U229;
  assign new_R152_U126 = new_R152_U287 & new_R152_U389;
  assign new_R152_U127 = new_R152_U284 & new_R152_U11 & new_R152_U286;
  assign new_R152_U128 = new_R152_U288 & new_R152_U146;
  assign new_R152_U129 = new_R152_U303 & new_R152_U223;
  assign new_R152_U130 = new_R152_U339 & new_R152_U338;
  assign new_R152_U131 = ~new_R152_U117 | ~new_R152_U331;
  assign new_R152_U132 = new_R152_U346 & new_R152_U345;
  assign new_R152_U133 = ~new_R152_U329 | ~new_R152_U18;
  assign new_R152_U134 = new_R152_U353 & new_R152_U352;
  assign new_R152_U135 = ~new_R152_U116 | ~new_R152_U296;
  assign new_R152_U136 = new_R152_U360 & new_R152_U359;
  assign new_R152_U137 = ~new_R152_U295 | ~new_R152_U293;
  assign new_R152_U138 = new_R152_U367 & new_R152_U366;
  assign new_R152_U139 = ~new_R152_U34 | ~new_R152_U203;
  assign new_R152_U140 = new_R152_U374 & new_R152_U373;
  assign new_R152_U141 = ~new_R152_U118 | ~new_R152_U315;
  assign new_R152_U142 = new_R152_U381 & new_R152_U380;
  assign new_R152_U143 = ~new_R152_U29 | ~new_R152_U310 | ~new_R152_U312 | ~new_R152_U311;
  assign new_R152_U144 = ~new_U132;
  assign new_R152_U145 = ~SI_31_;
  assign new_R152_U146 = new_R152_U393 & new_R152_U392;
  assign new_R152_U147 = new_R152_U395 & new_R152_U394;
  assign new_R152_U148 = ~new_R152_U284 | ~new_R152_U283;
  assign new_R152_U149 = ~new_R152_U289 | ~new_R152_U290 | ~new_R152_U171;
  assign new_R152_U150 = new_R152_U409 & new_R152_U408;
  assign new_R152_U151 = ~new_R152_U280 | ~new_R152_U279;
  assign new_R152_U152 = new_R152_U416 & new_R152_U415;
  assign new_R152_U153 = ~new_R152_U276 | ~new_R152_U275;
  assign new_R152_U154 = new_R152_U423 & new_R152_U422;
  assign new_R152_U155 = ~new_R152_U272 | ~new_R152_U271;
  assign new_R152_U156 = new_R152_U430 & new_R152_U429;
  assign new_R152_U157 = ~new_R152_U268 | ~new_R152_U267;
  assign new_R152_U158 = new_R152_U437 & new_R152_U436;
  assign new_R152_U159 = ~new_R152_U264 | ~new_R152_U263;
  assign new_R152_U160 = new_R152_U444 & new_R152_U443;
  assign new_R152_U161 = ~new_R152_U260 | ~new_R152_U259;
  assign new_R152_U162 = new_R152_U451 & new_R152_U450;
  assign new_R152_U163 = ~new_R152_U256 | ~new_R152_U255;
  assign new_R152_U164 = new_R152_U458 & new_R152_U457;
  assign new_R152_U165 = ~new_R152_U252 | ~new_R152_U251;
  assign new_R152_U166 = new_R152_U465 & new_R152_U464;
  assign new_R152_U167 = ~new_R152_U248 | ~new_R152_U247;
  assign new_R152_U168 = new_R152_U472 & new_R152_U471;
  assign new_R152_U169 = ~new_R152_U244 | ~new_R152_U243;
  assign new_R152_U170 = ~new_U157 | ~SI_0_;
  assign new_R152_U171 = ~new_U157 | ~SI_0_ | ~SI_1_;
  assign new_R152_U172 = new_R152_U482 & new_R152_U481;
  assign new_R152_U173 = new_R152_U484 & new_R152_U483;
  assign new_R152_U174 = ~new_R152_U240 | ~new_R152_U239;
  assign new_R152_U175 = new_R152_U491 & new_R152_U490;
  assign new_R152_U176 = ~new_R152_U236 | ~new_R152_U235;
  assign new_R152_U177 = new_R152_U498 & new_R152_U497;
  assign new_R152_U178 = ~new_R152_U232 | ~new_R152_U231;
  assign new_R152_U179 = new_R152_U505 & new_R152_U504;
  assign new_R152_U180 = ~new_R152_U125 | ~new_R152_U327;
  assign new_R152_U181 = new_R152_U512 & new_R152_U511;
  assign new_R152_U182 = ~new_R152_U308 | ~new_R152_U325;
  assign new_R152_U183 = new_R152_U519 & new_R152_U518;
  assign new_R152_U184 = ~new_R152_U306 | ~new_R152_U323;
  assign new_R152_U185 = new_R152_U526 & new_R152_U525;
  assign new_R152_U186 = ~new_R152_U129 | ~new_R152_U321;
  assign new_R152_U187 = new_R152_U533 & new_R152_U532;
  assign new_R152_U188 = ~new_R152_U319 | ~new_R152_U48;
  assign new_R152_U189 = new_R152_U540 & new_R152_U539;
  assign new_R152_U190 = ~new_R152_U123 | ~new_R152_U335;
  assign new_R152_U191 = new_R152_U547 & new_R152_U546;
  assign new_R152_U192 = ~new_R152_U301 | ~new_R152_U333;
  assign new_R152_U193 = ~new_R152_U126 | ~new_R152_U148;
  assign new_R152_U194 = ~new_R152_U171;
  assign new_R152_U195 = ~new_R152_U149;
  assign new_R152_U196 = SI_2_ | new_U145;
  assign new_R152_U197 = ~new_R152_U29;
  assign new_R152_U198 = ~new_R152_U143;
  assign new_R152_U199 = SI_3_ | new_U134;
  assign new_R152_U200 = ~new_U134 | ~SI_3_;
  assign new_R152_U201 = ~new_R152_U114 | ~new_R152_U291;
  assign new_R152_U202 = SI_4_ | new_U131;
  assign new_R152_U203 = ~new_R152_U202 | ~new_R152_U201;
  assign new_R152_U204 = ~new_R152_U34;
  assign new_R152_U205 = ~new_R152_U139;
  assign new_R152_U206 = SI_5_ | new_U130;
  assign new_R152_U207 = ~new_U130 | ~SI_5_;
  assign new_R152_U208 = ~new_R152_U137;
  assign new_R152_U209 = SI_6_ | new_U129;
  assign new_R152_U210 = ~new_U129 | ~SI_6_;
  assign new_R152_U211 = ~new_R152_U135;
  assign new_R152_U212 = SI_7_ | new_U128;
  assign new_R152_U213 = ~new_R152_U18;
  assign new_R152_U214 = SI_8_ | new_U127;
  assign new_R152_U215 = ~new_U127 | ~SI_8_;
  assign new_R152_U216 = SI_9_ | new_U126;
  assign new_R152_U217 = ~SI_9_ | ~new_U126;
  assign new_R152_U218 = SI_10_ | new_U155;
  assign new_R152_U219 = ~new_U155 | ~SI_10_;
  assign new_R152_U220 = SI_11_ | new_U154;
  assign new_R152_U221 = ~new_R152_U48;
  assign new_R152_U222 = SI_12_ | new_U153;
  assign new_R152_U223 = ~new_U153 | ~SI_12_;
  assign new_R152_U224 = SI_13_ | new_U152;
  assign new_R152_U225 = ~new_U152 | ~SI_13_;
  assign new_R152_U226 = SI_14_ | new_U151;
  assign new_R152_U227 = ~new_U151 | ~SI_14_;
  assign new_R152_U228 = SI_15_ | new_U150;
  assign new_R152_U229 = ~new_U150 | ~SI_15_;
  assign new_R152_U230 = SI_16_ | new_U149;
  assign new_R152_U231 = ~new_R152_U230 | ~new_R152_U180;
  assign new_R152_U232 = ~new_U149 | ~SI_16_;
  assign new_R152_U233 = ~new_R152_U178;
  assign new_R152_U234 = SI_17_ | new_U148;
  assign new_R152_U235 = ~new_R152_U234 | ~new_R152_U178;
  assign new_R152_U236 = ~new_U148 | ~SI_17_;
  assign new_R152_U237 = ~new_R152_U176;
  assign new_R152_U238 = SI_18_ | new_U147;
  assign new_R152_U239 = ~new_R152_U238 | ~new_R152_U176;
  assign new_R152_U240 = ~new_U147 | ~SI_18_;
  assign new_R152_U241 = ~new_R152_U174;
  assign new_R152_U242 = SI_19_ | new_U146;
  assign new_R152_U243 = ~new_R152_U242 | ~new_R152_U174;
  assign new_R152_U244 = ~new_U146 | ~SI_19_;
  assign new_R152_U245 = ~new_R152_U169;
  assign new_R152_U246 = SI_20_ | new_U144;
  assign new_R152_U247 = ~new_R152_U246 | ~new_R152_U169;
  assign new_R152_U248 = ~new_U144 | ~SI_20_;
  assign new_R152_U249 = ~new_R152_U167;
  assign new_R152_U250 = SI_21_ | new_U143;
  assign new_R152_U251 = ~new_R152_U250 | ~new_R152_U167;
  assign new_R152_U252 = ~new_U143 | ~SI_21_;
  assign new_R152_U253 = ~new_R152_U165;
  assign new_R152_U254 = SI_22_ | new_U142;
  assign new_R152_U255 = ~new_R152_U254 | ~new_R152_U165;
  assign new_R152_U256 = ~new_U142 | ~SI_22_;
  assign new_R152_U257 = ~new_R152_U163;
  assign new_R152_U258 = SI_23_ | new_U141;
  assign new_R152_U259 = ~new_R152_U258 | ~new_R152_U163;
  assign new_R152_U260 = ~new_U141 | ~SI_23_;
  assign new_R152_U261 = ~new_R152_U161;
  assign new_R152_U262 = SI_24_ | new_U140;
  assign new_R152_U263 = ~new_R152_U262 | ~new_R152_U161;
  assign new_R152_U264 = ~new_U140 | ~SI_24_;
  assign new_R152_U265 = ~new_R152_U159;
  assign new_R152_U266 = SI_25_ | new_U139;
  assign new_R152_U267 = ~new_R152_U266 | ~new_R152_U159;
  assign new_R152_U268 = ~new_U139 | ~SI_25_;
  assign new_R152_U269 = ~new_R152_U157;
  assign new_R152_U270 = SI_26_ | new_U138;
  assign new_R152_U271 = ~new_R152_U270 | ~new_R152_U157;
  assign new_R152_U272 = ~new_U138 | ~SI_26_;
  assign new_R152_U273 = ~new_R152_U155;
  assign new_R152_U274 = SI_27_ | new_U137;
  assign new_R152_U275 = ~new_R152_U274 | ~new_R152_U155;
  assign new_R152_U276 = ~new_U137 | ~SI_27_;
  assign new_R152_U277 = ~new_R152_U153;
  assign new_R152_U278 = SI_28_ | new_U136;
  assign new_R152_U279 = ~new_R152_U278 | ~new_R152_U153;
  assign new_R152_U280 = ~new_U136 | ~SI_28_;
  assign new_R152_U281 = ~new_R152_U151;
  assign new_R152_U282 = SI_29_ | new_U135;
  assign new_R152_U283 = ~new_R152_U282 | ~new_R152_U151;
  assign new_R152_U284 = ~new_U135 | ~SI_29_;
  assign new_R152_U285 = ~new_R152_U148;
  assign new_R152_U286 = ~new_U133 | ~SI_30_;
  assign new_R152_U287 = new_U133 | SI_30_;
  assign new_R152_U288 = ~new_R152_U283 | ~new_R152_U127;
  assign new_R152_U289 = ~new_U156 | ~new_U157 | ~SI_0_;
  assign new_R152_U290 = ~new_U156 | ~SI_1_;
  assign new_R152_U291 = ~new_R152_U10 | ~new_R152_U313;
  assign new_R152_U292 = ~new_R152_U197 | ~new_R152_U199;
  assign new_R152_U293 = ~new_R152_U4 | ~new_R152_U201;
  assign new_R152_U294 = ~new_R152_U204 | ~new_R152_U206;
  assign new_R152_U295 = ~new_R152_U37;
  assign new_R152_U296 = ~new_R152_U115 | ~new_R152_U201;
  assign new_R152_U297 = ~new_R152_U37 | ~new_R152_U209;
  assign new_R152_U298 = ~new_R152_U213 | ~new_R152_U214;
  assign new_R152_U299 = ~new_R152_U298 | ~new_R152_U215;
  assign new_R152_U300 = ~new_R152_U299 | ~new_R152_U216;
  assign new_R152_U301 = ~new_R152_U83;
  assign new_R152_U302 = ~new_R152_U83 | ~new_R152_U218;
  assign new_R152_U303 = ~new_R152_U221 | ~new_R152_U222;
  assign new_R152_U304 = ~new_R152_U303 | ~new_R152_U223;
  assign new_R152_U305 = ~new_R152_U304 | ~new_R152_U224;
  assign new_R152_U306 = ~new_R152_U82;
  assign new_R152_U307 = ~new_R152_U82 | ~new_R152_U226;
  assign new_R152_U308 = ~new_R152_U81;
  assign new_R152_U309 = ~new_R152_U81 | ~new_R152_U228;
  assign new_R152_U310 = ~new_R152_U119 | ~SI_0_ | ~new_R152_U196;
  assign new_R152_U311 = ~new_R152_U120 | ~SI_1_ | ~new_R152_U196;
  assign new_R152_U312 = ~new_R152_U121 | ~new_R152_U196;
  assign new_R152_U313 = ~new_R152_U289 | ~new_R152_U290 | ~new_R152_U171;
  assign new_R152_U314 = ~new_R152_U141;
  assign new_R152_U315 = ~new_R152_U10 | ~new_R152_U316;
  assign new_R152_U316 = ~new_R152_U317 | ~new_R152_U318 | ~new_R152_U290;
  assign new_R152_U317 = ~new_U156 | ~new_U157 | ~SI_0_;
  assign new_R152_U318 = ~new_U157 | ~SI_0_ | ~SI_1_;
  assign new_R152_U319 = ~new_R152_U220 | ~new_R152_U190;
  assign new_R152_U320 = ~new_R152_U188;
  assign new_R152_U321 = ~new_R152_U7 | ~new_R152_U190;
  assign new_R152_U322 = ~new_R152_U186;
  assign new_R152_U323 = ~new_R152_U8 | ~new_R152_U190;
  assign new_R152_U324 = ~new_R152_U184;
  assign new_R152_U325 = ~new_R152_U9 | ~new_R152_U190;
  assign new_R152_U326 = ~new_R152_U182;
  assign new_R152_U327 = ~new_R152_U124 | ~new_R152_U190;
  assign new_R152_U328 = ~new_R152_U180;
  assign new_R152_U329 = ~new_R152_U212 | ~new_R152_U135;
  assign new_R152_U330 = ~new_R152_U133;
  assign new_R152_U331 = ~new_R152_U5 | ~new_R152_U135;
  assign new_R152_U332 = ~new_R152_U131;
  assign new_R152_U333 = ~new_R152_U6 | ~new_R152_U135;
  assign new_R152_U334 = ~new_R152_U192;
  assign new_R152_U335 = ~new_R152_U122 | ~new_R152_U135;
  assign new_R152_U336 = ~new_R152_U190;
  assign new_R152_U337 = ~new_R152_U480 | ~new_R152_U23;
  assign new_R152_U338 = ~new_U126 | ~new_R152_U36;
  assign new_R152_U339 = ~SI_9_ | ~new_R152_U35;
  assign new_R152_U340 = ~new_U126 | ~new_R152_U36;
  assign new_R152_U341 = ~SI_9_ | ~new_R152_U35;
  assign new_R152_U342 = ~new_R152_U341 | ~new_R152_U340;
  assign new_R152_U343 = ~new_R152_U130 | ~new_R152_U131;
  assign new_R152_U344 = ~new_R152_U332 | ~new_R152_U342;
  assign new_R152_U345 = ~new_U127 | ~new_R152_U14;
  assign new_R152_U346 = ~SI_8_ | ~new_R152_U15;
  assign new_R152_U347 = ~new_U127 | ~new_R152_U14;
  assign new_R152_U348 = ~SI_8_ | ~new_R152_U15;
  assign new_R152_U349 = ~new_R152_U348 | ~new_R152_U347;
  assign new_R152_U350 = ~new_R152_U132 | ~new_R152_U133;
  assign new_R152_U351 = ~new_R152_U330 | ~new_R152_U349;
  assign new_R152_U352 = ~new_U128 | ~new_R152_U16;
  assign new_R152_U353 = ~SI_7_ | ~new_R152_U17;
  assign new_R152_U354 = ~new_U128 | ~new_R152_U16;
  assign new_R152_U355 = ~SI_7_ | ~new_R152_U17;
  assign new_R152_U356 = ~new_R152_U355 | ~new_R152_U354;
  assign new_R152_U357 = ~new_R152_U134 | ~new_R152_U135;
  assign new_R152_U358 = ~new_R152_U211 | ~new_R152_U356;
  assign new_R152_U359 = ~new_U129 | ~new_R152_U19;
  assign new_R152_U360 = ~SI_6_ | ~new_R152_U20;
  assign new_R152_U361 = ~new_U129 | ~new_R152_U19;
  assign new_R152_U362 = ~SI_6_ | ~new_R152_U20;
  assign new_R152_U363 = ~new_R152_U362 | ~new_R152_U361;
  assign new_R152_U364 = ~new_R152_U136 | ~new_R152_U137;
  assign new_R152_U365 = ~new_R152_U208 | ~new_R152_U363;
  assign new_R152_U366 = ~new_U130 | ~new_R152_U30;
  assign new_R152_U367 = ~SI_5_ | ~new_R152_U31;
  assign new_R152_U368 = ~new_U130 | ~new_R152_U30;
  assign new_R152_U369 = ~SI_5_ | ~new_R152_U31;
  assign new_R152_U370 = ~new_R152_U369 | ~new_R152_U368;
  assign new_R152_U371 = ~new_R152_U138 | ~new_R152_U139;
  assign new_R152_U372 = ~new_R152_U205 | ~new_R152_U370;
  assign new_R152_U373 = ~new_U131 | ~new_R152_U32;
  assign new_R152_U374 = ~SI_4_ | ~new_R152_U33;
  assign new_R152_U375 = ~new_U131 | ~new_R152_U32;
  assign new_R152_U376 = ~SI_4_ | ~new_R152_U33;
  assign new_R152_U377 = ~new_R152_U376 | ~new_R152_U375;
  assign new_R152_U378 = ~new_R152_U140 | ~new_R152_U141;
  assign new_R152_U379 = ~new_R152_U314 | ~new_R152_U377;
  assign new_R152_U380 = ~new_U134 | ~new_R152_U21;
  assign new_R152_U381 = ~SI_3_ | ~new_R152_U22;
  assign new_R152_U382 = ~new_U134 | ~new_R152_U21;
  assign new_R152_U383 = ~SI_3_ | ~new_R152_U22;
  assign new_R152_U384 = ~new_R152_U383 | ~new_R152_U382;
  assign new_R152_U385 = ~new_R152_U142 | ~new_R152_U143;
  assign new_R152_U386 = ~new_R152_U198 | ~new_R152_U384;
  assign new_R152_U387 = ~new_U132 | ~new_R152_U145;
  assign new_R152_U388 = ~SI_31_ | ~new_R152_U144;
  assign new_R152_U389 = ~new_R152_U388 | ~new_R152_U387;
  assign new_R152_U390 = ~new_U132 | ~new_R152_U145;
  assign new_R152_U391 = ~SI_31_ | ~new_R152_U144;
  assign new_R152_U392 = ~new_R152_U80 | ~new_R152_U11 | ~new_R152_U79;
  assign new_R152_U393 = ~new_U133 | ~SI_30_ | ~new_R152_U389;
  assign new_R152_U394 = ~new_U133 | ~new_R152_U79;
  assign new_R152_U395 = ~SI_30_ | ~new_R152_U80;
  assign new_R152_U396 = ~new_U133 | ~new_R152_U79;
  assign new_R152_U397 = ~SI_30_ | ~new_R152_U80;
  assign new_R152_U398 = ~new_R152_U397 | ~new_R152_U396;
  assign new_R152_U399 = ~new_R152_U147 | ~new_R152_U148;
  assign new_R152_U400 = ~new_R152_U285 | ~new_R152_U398;
  assign new_R152_U401 = ~new_U145 | ~new_R152_U27;
  assign new_R152_U402 = ~SI_2_ | ~new_R152_U28;
  assign new_R152_U403 = ~new_U145 | ~new_R152_U27;
  assign new_R152_U404 = ~SI_2_ | ~new_R152_U28;
  assign new_R152_U405 = ~new_R152_U404 | ~new_R152_U403;
  assign new_R152_U406 = ~new_R152_U149 | ~new_R152_U402 | ~new_R152_U401;
  assign new_R152_U407 = ~new_R152_U195 | ~new_R152_U405;
  assign new_R152_U408 = ~new_U135 | ~new_R152_U77;
  assign new_R152_U409 = ~SI_29_ | ~new_R152_U78;
  assign new_R152_U410 = ~new_U135 | ~new_R152_U77;
  assign new_R152_U411 = ~SI_29_ | ~new_R152_U78;
  assign new_R152_U412 = ~new_R152_U411 | ~new_R152_U410;
  assign new_R152_U413 = ~new_R152_U150 | ~new_R152_U151;
  assign new_R152_U414 = ~new_R152_U281 | ~new_R152_U412;
  assign new_R152_U415 = ~new_U136 | ~new_R152_U75;
  assign new_R152_U416 = ~SI_28_ | ~new_R152_U76;
  assign new_R152_U417 = ~new_U136 | ~new_R152_U75;
  assign new_R152_U418 = ~SI_28_ | ~new_R152_U76;
  assign new_R152_U419 = ~new_R152_U418 | ~new_R152_U417;
  assign new_R152_U420 = ~new_R152_U152 | ~new_R152_U153;
  assign new_R152_U421 = ~new_R152_U277 | ~new_R152_U419;
  assign new_R152_U422 = ~new_U137 | ~new_R152_U73;
  assign new_R152_U423 = ~SI_27_ | ~new_R152_U74;
  assign new_R152_U424 = ~new_U137 | ~new_R152_U73;
  assign new_R152_U425 = ~SI_27_ | ~new_R152_U74;
  assign new_R152_U426 = ~new_R152_U425 | ~new_R152_U424;
  assign new_R152_U427 = ~new_R152_U154 | ~new_R152_U155;
  assign new_R152_U428 = ~new_R152_U273 | ~new_R152_U426;
  assign new_R152_U429 = ~new_U138 | ~new_R152_U71;
  assign new_R152_U430 = ~SI_26_ | ~new_R152_U72;
  assign new_R152_U431 = ~new_U138 | ~new_R152_U71;
  assign new_R152_U432 = ~SI_26_ | ~new_R152_U72;
  assign new_R152_U433 = ~new_R152_U432 | ~new_R152_U431;
  assign new_R152_U434 = ~new_R152_U156 | ~new_R152_U157;
  assign new_R152_U435 = ~new_R152_U269 | ~new_R152_U433;
  assign new_R152_U436 = ~new_U139 | ~new_R152_U69;
  assign new_R152_U437 = ~SI_25_ | ~new_R152_U70;
  assign new_R152_U438 = ~new_U139 | ~new_R152_U69;
  assign new_R152_U439 = ~SI_25_ | ~new_R152_U70;
  assign new_R152_U440 = ~new_R152_U439 | ~new_R152_U438;
  assign new_R152_U441 = ~new_R152_U158 | ~new_R152_U159;
  assign new_R152_U442 = ~new_R152_U265 | ~new_R152_U440;
  assign new_R152_U443 = ~new_U140 | ~new_R152_U67;
  assign new_R152_U444 = ~SI_24_ | ~new_R152_U68;
  assign new_R152_U445 = ~new_U140 | ~new_R152_U67;
  assign new_R152_U446 = ~SI_24_ | ~new_R152_U68;
  assign new_R152_U447 = ~new_R152_U446 | ~new_R152_U445;
  assign new_R152_U448 = ~new_R152_U160 | ~new_R152_U161;
  assign new_R152_U449 = ~new_R152_U261 | ~new_R152_U447;
  assign new_R152_U450 = ~new_U141 | ~new_R152_U65;
  assign new_R152_U451 = ~SI_23_ | ~new_R152_U66;
  assign new_R152_U452 = ~new_U141 | ~new_R152_U65;
  assign new_R152_U453 = ~SI_23_ | ~new_R152_U66;
  assign new_R152_U454 = ~new_R152_U453 | ~new_R152_U452;
  assign new_R152_U455 = ~new_R152_U162 | ~new_R152_U163;
  assign new_R152_U456 = ~new_R152_U257 | ~new_R152_U454;
  assign new_R152_U457 = ~new_U142 | ~new_R152_U63;
  assign new_R152_U458 = ~SI_22_ | ~new_R152_U64;
  assign new_R152_U459 = ~new_U142 | ~new_R152_U63;
  assign new_R152_U460 = ~SI_22_ | ~new_R152_U64;
  assign new_R152_U461 = ~new_R152_U460 | ~new_R152_U459;
  assign new_R152_U462 = ~new_R152_U164 | ~new_R152_U165;
  assign new_R152_U463 = ~new_R152_U253 | ~new_R152_U461;
  assign new_R152_U464 = ~new_U143 | ~new_R152_U61;
  assign new_R152_U465 = ~SI_21_ | ~new_R152_U62;
  assign new_R152_U466 = ~new_U143 | ~new_R152_U61;
  assign new_R152_U467 = ~SI_21_ | ~new_R152_U62;
  assign new_R152_U468 = ~new_R152_U467 | ~new_R152_U466;
  assign new_R152_U469 = ~new_R152_U166 | ~new_R152_U167;
  assign new_R152_U470 = ~new_R152_U249 | ~new_R152_U468;
  assign new_R152_U471 = ~new_U144 | ~new_R152_U59;
  assign new_R152_U472 = ~SI_20_ | ~new_R152_U60;
  assign new_R152_U473 = ~new_U144 | ~new_R152_U59;
  assign new_R152_U474 = ~SI_20_ | ~new_R152_U60;
  assign new_R152_U475 = ~new_R152_U474 | ~new_R152_U473;
  assign new_R152_U476 = ~new_R152_U168 | ~new_R152_U169;
  assign new_R152_U477 = ~new_R152_U245 | ~new_R152_U475;
  assign new_R152_U478 = ~new_U156 | ~new_R152_U170;
  assign new_R152_U479 = ~new_R152_U120 | ~new_R152_U26;
  assign new_R152_U480 = ~new_R152_U479 | ~new_R152_U478;
  assign new_R152_U481 = ~new_R152_U26 | ~SI_1_ | ~new_R152_U170;
  assign new_R152_U482 = ~new_R152_U194 | ~new_U156;
  assign new_R152_U483 = ~new_U146 | ~new_R152_U57;
  assign new_R152_U484 = ~SI_19_ | ~new_R152_U58;
  assign new_R152_U485 = ~new_U146 | ~new_R152_U57;
  assign new_R152_U486 = ~SI_19_ | ~new_R152_U58;
  assign new_R152_U487 = ~new_R152_U486 | ~new_R152_U485;
  assign new_R152_U488 = ~new_R152_U173 | ~new_R152_U174;
  assign new_R152_U489 = ~new_R152_U241 | ~new_R152_U487;
  assign new_R152_U490 = ~new_U147 | ~new_R152_U55;
  assign new_R152_U491 = ~SI_18_ | ~new_R152_U56;
  assign new_R152_U492 = ~new_U147 | ~new_R152_U55;
  assign new_R152_U493 = ~SI_18_ | ~new_R152_U56;
  assign new_R152_U494 = ~new_R152_U493 | ~new_R152_U492;
  assign new_R152_U495 = ~new_R152_U175 | ~new_R152_U176;
  assign new_R152_U496 = ~new_R152_U237 | ~new_R152_U494;
  assign new_R152_U497 = ~new_U148 | ~new_R152_U53;
  assign new_R152_U498 = ~SI_17_ | ~new_R152_U54;
  assign new_R152_U499 = ~new_U148 | ~new_R152_U53;
  assign new_R152_U500 = ~SI_17_ | ~new_R152_U54;
  assign new_R152_U501 = ~new_R152_U500 | ~new_R152_U499;
  assign new_R152_U502 = ~new_R152_U177 | ~new_R152_U178;
  assign new_R152_U503 = ~new_R152_U233 | ~new_R152_U501;
  assign new_R152_U504 = ~new_U149 | ~new_R152_U51;
  assign new_R152_U505 = ~SI_16_ | ~new_R152_U52;
  assign new_R152_U506 = ~new_U149 | ~new_R152_U51;
  assign new_R152_U507 = ~SI_16_ | ~new_R152_U52;
  assign new_R152_U508 = ~new_R152_U507 | ~new_R152_U506;
  assign new_R152_U509 = ~new_R152_U179 | ~new_R152_U180;
  assign new_R152_U510 = ~new_R152_U328 | ~new_R152_U508;
  assign new_R152_U511 = ~new_U150 | ~new_R152_U38;
  assign new_R152_U512 = ~SI_15_ | ~new_R152_U39;
  assign new_R152_U513 = ~new_U150 | ~new_R152_U38;
  assign new_R152_U514 = ~SI_15_ | ~new_R152_U39;
  assign new_R152_U515 = ~new_R152_U514 | ~new_R152_U513;
  assign new_R152_U516 = ~new_R152_U181 | ~new_R152_U182;
  assign new_R152_U517 = ~new_R152_U326 | ~new_R152_U515;
  assign new_R152_U518 = ~new_U151 | ~new_R152_U40;
  assign new_R152_U519 = ~SI_14_ | ~new_R152_U41;
  assign new_R152_U520 = ~new_U151 | ~new_R152_U40;
  assign new_R152_U521 = ~SI_14_ | ~new_R152_U41;
  assign new_R152_U522 = ~new_R152_U521 | ~new_R152_U520;
  assign new_R152_U523 = ~new_R152_U183 | ~new_R152_U184;
  assign new_R152_U524 = ~new_R152_U324 | ~new_R152_U522;
  assign new_R152_U525 = ~new_U152 | ~new_R152_U42;
  assign new_R152_U526 = ~SI_13_ | ~new_R152_U43;
  assign new_R152_U527 = ~new_U152 | ~new_R152_U42;
  assign new_R152_U528 = ~SI_13_ | ~new_R152_U43;
  assign new_R152_U529 = ~new_R152_U528 | ~new_R152_U527;
  assign new_R152_U530 = ~new_R152_U185 | ~new_R152_U186;
  assign new_R152_U531 = ~new_R152_U322 | ~new_R152_U529;
  assign new_R152_U532 = ~new_U153 | ~new_R152_U44;
  assign new_R152_U533 = ~SI_12_ | ~new_R152_U45;
  assign new_R152_U534 = ~new_U153 | ~new_R152_U44;
  assign new_R152_U535 = ~SI_12_ | ~new_R152_U45;
  assign new_R152_U536 = ~new_R152_U535 | ~new_R152_U534;
  assign new_R152_U537 = ~new_R152_U187 | ~new_R152_U188;
  assign new_R152_U538 = ~new_R152_U320 | ~new_R152_U536;
  assign new_R152_U539 = ~new_U154 | ~new_R152_U46;
  assign new_R152_U540 = ~SI_11_ | ~new_R152_U47;
  assign new_R152_U541 = ~new_U154 | ~new_R152_U46;
  assign new_R152_U542 = ~SI_11_ | ~new_R152_U47;
  assign new_R152_U543 = ~new_R152_U542 | ~new_R152_U541;
  assign new_R152_U544 = ~new_R152_U189 | ~new_R152_U190;
  assign new_R152_U545 = ~new_R152_U336 | ~new_R152_U543;
  assign new_R152_U546 = ~new_U155 | ~new_R152_U49;
  assign new_R152_U547 = ~SI_10_ | ~new_R152_U50;
  assign new_R152_U548 = ~new_U155 | ~new_R152_U49;
  assign new_R152_U549 = ~SI_10_ | ~new_R152_U50;
  assign new_R152_U550 = ~new_R152_U549 | ~new_R152_U548;
  assign new_R152_U551 = ~new_R152_U191 | ~new_R152_U192;
  assign new_R152_U552 = ~new_R152_U334 | ~new_R152_U550;
  assign new_R152_U553 = ~new_U157 | ~new_R152_U24;
  assign new_R152_U554 = ~SI_0_ | ~new_R152_U25;
  assign new_LT_1602_U6 = ~P3_ADDR_REG_19_;
  assign new_LT_1601_U6 = ~P1_ADDR_REG_19_;
  assign SUB_1596_U4 = new_SUB_1596_U159 & new_SUB_1596_U155;
  assign SUB_1596_U5 = ~new_SUB_1596_U160 | ~new_SUB_1596_U221 | ~new_SUB_1596_U220;
  assign new_SUB_1596_U6 = ~new_ADD_1596_U7;
  assign new_SUB_1596_U7 = ~P2_ADDR_REG_0_;
  assign new_SUB_1596_U8 = ~P2_ADDR_REG_1_;
  assign new_SUB_1596_U9 = ~P2_ADDR_REG_0_ | ~new_ADD_1596_U7;
  assign new_SUB_1596_U10 = ~new_ADD_1596_U55;
  assign new_SUB_1596_U11 = ~new_ADD_1596_U54;
  assign new_SUB_1596_U12 = ~P2_ADDR_REG_2_;
  assign new_SUB_1596_U13 = ~new_SUB_1596_U90 | ~new_SUB_1596_U89;
  assign new_SUB_1596_U14 = ~new_ADD_1596_U53;
  assign new_SUB_1596_U15 = ~P2_ADDR_REG_3_;
  assign new_SUB_1596_U16 = ~new_ADD_1596_U52;
  assign new_SUB_1596_U17 = ~P2_ADDR_REG_4_;
  assign new_SUB_1596_U18 = ~new_SUB_1596_U98 | ~new_SUB_1596_U97;
  assign new_SUB_1596_U19 = ~new_ADD_1596_U51;
  assign new_SUB_1596_U20 = ~P2_ADDR_REG_5_;
  assign new_SUB_1596_U21 = ~new_ADD_1596_U50;
  assign new_SUB_1596_U22 = ~P2_ADDR_REG_6_;
  assign new_SUB_1596_U23 = ~new_ADD_1596_U49;
  assign new_SUB_1596_U24 = ~P2_ADDR_REG_7_;
  assign new_SUB_1596_U25 = ~new_SUB_1596_U110 | ~new_SUB_1596_U109;
  assign new_SUB_1596_U26 = ~new_ADD_1596_U48;
  assign new_SUB_1596_U27 = ~P2_ADDR_REG_8_;
  assign new_SUB_1596_U28 = ~P2_ADDR_REG_9_;
  assign new_SUB_1596_U29 = ~new_ADD_1596_U47;
  assign new_SUB_1596_U30 = ~new_SUB_1596_U118 | ~new_SUB_1596_U117;
  assign new_SUB_1596_U31 = ~new_ADD_1596_U64;
  assign new_SUB_1596_U32 = ~P2_ADDR_REG_10_;
  assign new_SUB_1596_U33 = ~new_ADD_1596_U63;
  assign new_SUB_1596_U34 = ~P2_ADDR_REG_11_;
  assign new_SUB_1596_U35 = ~new_ADD_1596_U62;
  assign new_SUB_1596_U36 = ~P2_ADDR_REG_12_;
  assign new_SUB_1596_U37 = ~new_SUB_1596_U130 | ~new_SUB_1596_U129;
  assign new_SUB_1596_U38 = ~new_ADD_1596_U61;
  assign new_SUB_1596_U39 = ~P2_ADDR_REG_13_;
  assign new_SUB_1596_U40 = ~new_SUB_1596_U134 | ~new_SUB_1596_U133;
  assign new_SUB_1596_U41 = ~new_ADD_1596_U60;
  assign new_SUB_1596_U42 = ~P2_ADDR_REG_14_;
  assign new_SUB_1596_U43 = ~new_SUB_1596_U138 | ~new_SUB_1596_U137;
  assign new_SUB_1596_U44 = ~new_ADD_1596_U59;
  assign new_SUB_1596_U45 = ~P2_ADDR_REG_15_;
  assign new_SUB_1596_U46 = ~new_ADD_1596_U58;
  assign new_SUB_1596_U47 = ~P2_ADDR_REG_16_;
  assign new_SUB_1596_U48 = ~new_ADD_1596_U57;
  assign new_SUB_1596_U49 = ~P2_ADDR_REG_17_;
  assign new_SUB_1596_U50 = ~new_SUB_1596_U150 | ~new_SUB_1596_U149;
  assign new_SUB_1596_U51 = ~new_ADD_1596_U56;
  assign new_SUB_1596_U52 = ~P2_ADDR_REG_18_;
  assign SUB_1596_U53 = ~new_SUB_1596_U291 | ~new_SUB_1596_U290;
  assign SUB_1596_U54 = ~new_SUB_1596_U167 | ~new_SUB_1596_U166;
  assign SUB_1596_U55 = ~new_SUB_1596_U174 | ~new_SUB_1596_U173;
  assign SUB_1596_U56 = ~new_SUB_1596_U181 | ~new_SUB_1596_U180;
  assign SUB_1596_U57 = ~new_SUB_1596_U188 | ~new_SUB_1596_U187;
  assign SUB_1596_U58 = ~new_SUB_1596_U195 | ~new_SUB_1596_U194;
  assign SUB_1596_U59 = ~new_SUB_1596_U202 | ~new_SUB_1596_U201;
  assign SUB_1596_U60 = ~new_SUB_1596_U209 | ~new_SUB_1596_U208;
  assign SUB_1596_U61 = ~new_SUB_1596_U216 | ~new_SUB_1596_U215;
  assign SUB_1596_U62 = ~new_SUB_1596_U233 | ~new_SUB_1596_U232;
  assign SUB_1596_U63 = ~new_SUB_1596_U240 | ~new_SUB_1596_U239;
  assign SUB_1596_U64 = ~new_SUB_1596_U247 | ~new_SUB_1596_U246;
  assign SUB_1596_U65 = ~new_SUB_1596_U254 | ~new_SUB_1596_U253;
  assign SUB_1596_U66 = ~new_SUB_1596_U261 | ~new_SUB_1596_U260;
  assign SUB_1596_U67 = ~new_SUB_1596_U268 | ~new_SUB_1596_U267;
  assign SUB_1596_U68 = ~new_SUB_1596_U275 | ~new_SUB_1596_U274;
  assign SUB_1596_U69 = ~new_SUB_1596_U282 | ~new_SUB_1596_U281;
  assign SUB_1596_U70 = ~new_SUB_1596_U289 | ~new_SUB_1596_U288;
  assign new_SUB_1596_U71 = ~new_SUB_1596_U114 | ~new_SUB_1596_U113;
  assign new_SUB_1596_U72 = ~new_SUB_1596_U106 | ~new_SUB_1596_U105;
  assign new_SUB_1596_U73 = ~new_SUB_1596_U102 | ~new_SUB_1596_U101;
  assign new_SUB_1596_U74 = ~new_SUB_1596_U94 | ~new_SUB_1596_U93;
  assign new_SUB_1596_U75 = ~new_SUB_1596_U76 | ~new_SUB_1596_U86;
  assign new_SUB_1596_U76 = ~new_ADD_1596_U55 | ~new_SUB_1596_U84;
  assign new_SUB_1596_U77 = ~P2_ADDR_REG_19_;
  assign new_SUB_1596_U78 = ~new_ADD_1596_U6;
  assign new_SUB_1596_U79 = ~new_SUB_1596_U146 | ~new_SUB_1596_U145;
  assign new_SUB_1596_U80 = ~new_SUB_1596_U142 | ~new_SUB_1596_U141;
  assign new_SUB_1596_U81 = ~new_SUB_1596_U126 | ~new_SUB_1596_U125;
  assign new_SUB_1596_U82 = ~new_SUB_1596_U122 | ~new_SUB_1596_U121;
  assign new_SUB_1596_U83 = ~new_SUB_1596_U76;
  assign new_SUB_1596_U84 = ~new_SUB_1596_U9;
  assign new_SUB_1596_U85 = ~new_SUB_1596_U10 | ~new_SUB_1596_U9;
  assign new_SUB_1596_U86 = ~P2_ADDR_REG_1_ | ~new_SUB_1596_U85;
  assign new_SUB_1596_U87 = ~new_SUB_1596_U75;
  assign new_SUB_1596_U88 = new_ADD_1596_U54 | P2_ADDR_REG_2_;
  assign new_SUB_1596_U89 = ~new_SUB_1596_U88 | ~new_SUB_1596_U75;
  assign new_SUB_1596_U90 = ~P2_ADDR_REG_2_ | ~new_ADD_1596_U54;
  assign new_SUB_1596_U91 = ~new_SUB_1596_U13;
  assign new_SUB_1596_U92 = ~new_SUB_1596_U91 | ~new_SUB_1596_U15;
  assign new_SUB_1596_U93 = ~new_ADD_1596_U53 | ~new_SUB_1596_U92;
  assign new_SUB_1596_U94 = ~P2_ADDR_REG_3_ | ~new_SUB_1596_U13;
  assign new_SUB_1596_U95 = ~new_SUB_1596_U74;
  assign new_SUB_1596_U96 = new_ADD_1596_U52 | P2_ADDR_REG_4_;
  assign new_SUB_1596_U97 = ~new_SUB_1596_U96 | ~new_SUB_1596_U74;
  assign new_SUB_1596_U98 = ~P2_ADDR_REG_4_ | ~new_ADD_1596_U52;
  assign new_SUB_1596_U99 = ~new_SUB_1596_U18;
  assign new_SUB_1596_U100 = ~new_SUB_1596_U99 | ~new_SUB_1596_U20;
  assign new_SUB_1596_U101 = ~new_ADD_1596_U51 | ~new_SUB_1596_U100;
  assign new_SUB_1596_U102 = ~P2_ADDR_REG_5_ | ~new_SUB_1596_U18;
  assign new_SUB_1596_U103 = ~new_SUB_1596_U73;
  assign new_SUB_1596_U104 = new_ADD_1596_U50 | P2_ADDR_REG_6_;
  assign new_SUB_1596_U105 = ~new_SUB_1596_U104 | ~new_SUB_1596_U73;
  assign new_SUB_1596_U106 = ~P2_ADDR_REG_6_ | ~new_ADD_1596_U50;
  assign new_SUB_1596_U107 = ~new_SUB_1596_U72;
  assign new_SUB_1596_U108 = new_ADD_1596_U49 | P2_ADDR_REG_7_;
  assign new_SUB_1596_U109 = ~new_SUB_1596_U108 | ~new_SUB_1596_U72;
  assign new_SUB_1596_U110 = ~P2_ADDR_REG_7_ | ~new_ADD_1596_U49;
  assign new_SUB_1596_U111 = ~new_SUB_1596_U25;
  assign new_SUB_1596_U112 = ~new_SUB_1596_U111 | ~new_SUB_1596_U27;
  assign new_SUB_1596_U113 = ~new_ADD_1596_U48 | ~new_SUB_1596_U112;
  assign new_SUB_1596_U114 = ~P2_ADDR_REG_8_ | ~new_SUB_1596_U25;
  assign new_SUB_1596_U115 = ~new_SUB_1596_U71;
  assign new_SUB_1596_U116 = new_ADD_1596_U47 | P2_ADDR_REG_9_;
  assign new_SUB_1596_U117 = ~new_SUB_1596_U116 | ~new_SUB_1596_U71;
  assign new_SUB_1596_U118 = ~new_ADD_1596_U47 | ~P2_ADDR_REG_9_;
  assign new_SUB_1596_U119 = ~new_SUB_1596_U30;
  assign new_SUB_1596_U120 = ~new_SUB_1596_U119 | ~new_SUB_1596_U32;
  assign new_SUB_1596_U121 = ~new_ADD_1596_U64 | ~new_SUB_1596_U120;
  assign new_SUB_1596_U122 = ~P2_ADDR_REG_10_ | ~new_SUB_1596_U30;
  assign new_SUB_1596_U123 = ~new_SUB_1596_U82;
  assign new_SUB_1596_U124 = new_ADD_1596_U63 | P2_ADDR_REG_11_;
  assign new_SUB_1596_U125 = ~new_SUB_1596_U124 | ~new_SUB_1596_U82;
  assign new_SUB_1596_U126 = ~P2_ADDR_REG_11_ | ~new_ADD_1596_U63;
  assign new_SUB_1596_U127 = ~new_SUB_1596_U81;
  assign new_SUB_1596_U128 = new_ADD_1596_U62 | P2_ADDR_REG_12_;
  assign new_SUB_1596_U129 = ~new_SUB_1596_U128 | ~new_SUB_1596_U81;
  assign new_SUB_1596_U130 = ~P2_ADDR_REG_12_ | ~new_ADD_1596_U62;
  assign new_SUB_1596_U131 = ~new_SUB_1596_U37;
  assign new_SUB_1596_U132 = ~new_SUB_1596_U131 | ~new_SUB_1596_U39;
  assign new_SUB_1596_U133 = ~new_ADD_1596_U61 | ~new_SUB_1596_U132;
  assign new_SUB_1596_U134 = ~P2_ADDR_REG_13_ | ~new_SUB_1596_U37;
  assign new_SUB_1596_U135 = ~new_SUB_1596_U40;
  assign new_SUB_1596_U136 = ~new_SUB_1596_U135 | ~new_SUB_1596_U42;
  assign new_SUB_1596_U137 = ~new_ADD_1596_U60 | ~new_SUB_1596_U136;
  assign new_SUB_1596_U138 = ~P2_ADDR_REG_14_ | ~new_SUB_1596_U40;
  assign new_SUB_1596_U139 = ~new_SUB_1596_U43;
  assign new_SUB_1596_U140 = ~new_SUB_1596_U139 | ~new_SUB_1596_U45;
  assign new_SUB_1596_U141 = ~new_ADD_1596_U59 | ~new_SUB_1596_U140;
  assign new_SUB_1596_U142 = ~P2_ADDR_REG_15_ | ~new_SUB_1596_U43;
  assign new_SUB_1596_U143 = ~new_SUB_1596_U80;
  assign new_SUB_1596_U144 = new_ADD_1596_U58 | P2_ADDR_REG_16_;
  assign new_SUB_1596_U145 = ~new_SUB_1596_U144 | ~new_SUB_1596_U80;
  assign new_SUB_1596_U146 = ~P2_ADDR_REG_16_ | ~new_ADD_1596_U58;
  assign new_SUB_1596_U147 = ~new_SUB_1596_U79;
  assign new_SUB_1596_U148 = new_ADD_1596_U57 | P2_ADDR_REG_17_;
  assign new_SUB_1596_U149 = ~new_SUB_1596_U148 | ~new_SUB_1596_U79;
  assign new_SUB_1596_U150 = ~P2_ADDR_REG_17_ | ~new_ADD_1596_U57;
  assign new_SUB_1596_U151 = ~new_SUB_1596_U50;
  assign new_SUB_1596_U152 = ~new_SUB_1596_U151 | ~new_SUB_1596_U52;
  assign new_SUB_1596_U153 = ~new_ADD_1596_U56 | ~new_SUB_1596_U152;
  assign new_SUB_1596_U154 = ~P2_ADDR_REG_18_ | ~new_SUB_1596_U50;
  assign new_SUB_1596_U155 = ~new_SUB_1596_U222 | ~new_SUB_1596_U223 | ~new_SUB_1596_U154 | ~new_SUB_1596_U153;
  assign new_SUB_1596_U156 = ~P2_ADDR_REG_18_ | ~new_SUB_1596_U50;
  assign new_SUB_1596_U157 = ~new_SUB_1596_U156 | ~new_SUB_1596_U51;
  assign new_SUB_1596_U158 = ~new_SUB_1596_U151 | ~new_SUB_1596_U52;
  assign new_SUB_1596_U159 = ~new_SUB_1596_U226 | ~new_SUB_1596_U158 | ~new_SUB_1596_U157;
  assign new_SUB_1596_U160 = ~new_SUB_1596_U219 | ~new_SUB_1596_U10;
  assign new_SUB_1596_U161 = ~P2_ADDR_REG_9_ | ~new_SUB_1596_U29;
  assign new_SUB_1596_U162 = ~new_ADD_1596_U47 | ~new_SUB_1596_U28;
  assign new_SUB_1596_U163 = ~P2_ADDR_REG_9_ | ~new_SUB_1596_U29;
  assign new_SUB_1596_U164 = ~new_ADD_1596_U47 | ~new_SUB_1596_U28;
  assign new_SUB_1596_U165 = ~new_SUB_1596_U164 | ~new_SUB_1596_U163;
  assign new_SUB_1596_U166 = ~new_SUB_1596_U71 | ~new_SUB_1596_U162 | ~new_SUB_1596_U161;
  assign new_SUB_1596_U167 = ~new_SUB_1596_U115 | ~new_SUB_1596_U165;
  assign new_SUB_1596_U168 = ~P2_ADDR_REG_8_ | ~new_SUB_1596_U25;
  assign new_SUB_1596_U169 = ~new_SUB_1596_U111 | ~new_SUB_1596_U27;
  assign new_SUB_1596_U170 = ~P2_ADDR_REG_8_ | ~new_SUB_1596_U25;
  assign new_SUB_1596_U171 = ~new_SUB_1596_U111 | ~new_SUB_1596_U27;
  assign new_SUB_1596_U172 = ~new_SUB_1596_U171 | ~new_SUB_1596_U170;
  assign new_SUB_1596_U173 = ~new_SUB_1596_U26 | ~new_SUB_1596_U169 | ~new_SUB_1596_U168;
  assign new_SUB_1596_U174 = ~new_SUB_1596_U172 | ~new_ADD_1596_U48;
  assign new_SUB_1596_U175 = ~P2_ADDR_REG_7_ | ~new_SUB_1596_U23;
  assign new_SUB_1596_U176 = ~new_ADD_1596_U49 | ~new_SUB_1596_U24;
  assign new_SUB_1596_U177 = ~P2_ADDR_REG_7_ | ~new_SUB_1596_U23;
  assign new_SUB_1596_U178 = ~new_ADD_1596_U49 | ~new_SUB_1596_U24;
  assign new_SUB_1596_U179 = ~new_SUB_1596_U178 | ~new_SUB_1596_U177;
  assign new_SUB_1596_U180 = ~new_SUB_1596_U72 | ~new_SUB_1596_U176 | ~new_SUB_1596_U175;
  assign new_SUB_1596_U181 = ~new_SUB_1596_U107 | ~new_SUB_1596_U179;
  assign new_SUB_1596_U182 = ~P2_ADDR_REG_6_ | ~new_SUB_1596_U21;
  assign new_SUB_1596_U183 = ~new_ADD_1596_U50 | ~new_SUB_1596_U22;
  assign new_SUB_1596_U184 = ~P2_ADDR_REG_6_ | ~new_SUB_1596_U21;
  assign new_SUB_1596_U185 = ~new_ADD_1596_U50 | ~new_SUB_1596_U22;
  assign new_SUB_1596_U186 = ~new_SUB_1596_U185 | ~new_SUB_1596_U184;
  assign new_SUB_1596_U187 = ~new_SUB_1596_U73 | ~new_SUB_1596_U183 | ~new_SUB_1596_U182;
  assign new_SUB_1596_U188 = ~new_SUB_1596_U103 | ~new_SUB_1596_U186;
  assign new_SUB_1596_U189 = ~P2_ADDR_REG_5_ | ~new_SUB_1596_U18;
  assign new_SUB_1596_U190 = ~new_SUB_1596_U99 | ~new_SUB_1596_U20;
  assign new_SUB_1596_U191 = ~P2_ADDR_REG_5_ | ~new_SUB_1596_U18;
  assign new_SUB_1596_U192 = ~new_SUB_1596_U99 | ~new_SUB_1596_U20;
  assign new_SUB_1596_U193 = ~new_SUB_1596_U192 | ~new_SUB_1596_U191;
  assign new_SUB_1596_U194 = ~new_SUB_1596_U19 | ~new_SUB_1596_U190 | ~new_SUB_1596_U189;
  assign new_SUB_1596_U195 = ~new_SUB_1596_U193 | ~new_ADD_1596_U51;
  assign new_SUB_1596_U196 = ~P2_ADDR_REG_4_ | ~new_SUB_1596_U16;
  assign new_SUB_1596_U197 = ~new_ADD_1596_U52 | ~new_SUB_1596_U17;
  assign new_SUB_1596_U198 = ~P2_ADDR_REG_4_ | ~new_SUB_1596_U16;
  assign new_SUB_1596_U199 = ~new_ADD_1596_U52 | ~new_SUB_1596_U17;
  assign new_SUB_1596_U200 = ~new_SUB_1596_U199 | ~new_SUB_1596_U198;
  assign new_SUB_1596_U201 = ~new_SUB_1596_U74 | ~new_SUB_1596_U197 | ~new_SUB_1596_U196;
  assign new_SUB_1596_U202 = ~new_SUB_1596_U95 | ~new_SUB_1596_U200;
  assign new_SUB_1596_U203 = ~P2_ADDR_REG_3_ | ~new_SUB_1596_U13;
  assign new_SUB_1596_U204 = ~new_SUB_1596_U91 | ~new_SUB_1596_U15;
  assign new_SUB_1596_U205 = ~P2_ADDR_REG_3_ | ~new_SUB_1596_U13;
  assign new_SUB_1596_U206 = ~new_SUB_1596_U91 | ~new_SUB_1596_U15;
  assign new_SUB_1596_U207 = ~new_SUB_1596_U206 | ~new_SUB_1596_U205;
  assign new_SUB_1596_U208 = ~new_SUB_1596_U14 | ~new_SUB_1596_U204 | ~new_SUB_1596_U203;
  assign new_SUB_1596_U209 = ~new_SUB_1596_U207 | ~new_ADD_1596_U53;
  assign new_SUB_1596_U210 = ~P2_ADDR_REG_2_ | ~new_SUB_1596_U11;
  assign new_SUB_1596_U211 = ~new_ADD_1596_U54 | ~new_SUB_1596_U12;
  assign new_SUB_1596_U212 = ~P2_ADDR_REG_2_ | ~new_SUB_1596_U11;
  assign new_SUB_1596_U213 = ~new_ADD_1596_U54 | ~new_SUB_1596_U12;
  assign new_SUB_1596_U214 = ~new_SUB_1596_U213 | ~new_SUB_1596_U212;
  assign new_SUB_1596_U215 = ~new_SUB_1596_U75 | ~new_SUB_1596_U211 | ~new_SUB_1596_U210;
  assign new_SUB_1596_U216 = ~new_SUB_1596_U87 | ~new_SUB_1596_U214;
  assign new_SUB_1596_U217 = ~P2_ADDR_REG_1_ | ~new_SUB_1596_U9;
  assign new_SUB_1596_U218 = ~new_SUB_1596_U84 | ~new_SUB_1596_U8;
  assign new_SUB_1596_U219 = ~new_SUB_1596_U218 | ~new_SUB_1596_U217;
  assign new_SUB_1596_U220 = ~new_SUB_1596_U8 | ~new_ADD_1596_U55 | ~new_SUB_1596_U9;
  assign new_SUB_1596_U221 = ~new_SUB_1596_U83 | ~P2_ADDR_REG_1_;
  assign new_SUB_1596_U222 = ~P2_ADDR_REG_19_ | ~new_SUB_1596_U78;
  assign new_SUB_1596_U223 = ~new_ADD_1596_U6 | ~new_SUB_1596_U77;
  assign new_SUB_1596_U224 = ~P2_ADDR_REG_19_ | ~new_SUB_1596_U78;
  assign new_SUB_1596_U225 = ~new_ADD_1596_U6 | ~new_SUB_1596_U77;
  assign new_SUB_1596_U226 = ~new_SUB_1596_U225 | ~new_SUB_1596_U224;
  assign new_SUB_1596_U227 = ~P2_ADDR_REG_18_ | ~new_SUB_1596_U50;
  assign new_SUB_1596_U228 = ~new_SUB_1596_U151 | ~new_SUB_1596_U52;
  assign new_SUB_1596_U229 = ~P2_ADDR_REG_18_ | ~new_SUB_1596_U50;
  assign new_SUB_1596_U230 = ~new_SUB_1596_U151 | ~new_SUB_1596_U52;
  assign new_SUB_1596_U231 = ~new_SUB_1596_U230 | ~new_SUB_1596_U229;
  assign new_SUB_1596_U232 = ~new_SUB_1596_U51 | ~new_SUB_1596_U228 | ~new_SUB_1596_U227;
  assign new_SUB_1596_U233 = ~new_SUB_1596_U231 | ~new_ADD_1596_U56;
  assign new_SUB_1596_U234 = ~P2_ADDR_REG_17_ | ~new_SUB_1596_U48;
  assign new_SUB_1596_U235 = ~new_ADD_1596_U57 | ~new_SUB_1596_U49;
  assign new_SUB_1596_U236 = ~P2_ADDR_REG_17_ | ~new_SUB_1596_U48;
  assign new_SUB_1596_U237 = ~new_ADD_1596_U57 | ~new_SUB_1596_U49;
  assign new_SUB_1596_U238 = ~new_SUB_1596_U237 | ~new_SUB_1596_U236;
  assign new_SUB_1596_U239 = ~new_SUB_1596_U79 | ~new_SUB_1596_U235 | ~new_SUB_1596_U234;
  assign new_SUB_1596_U240 = ~new_SUB_1596_U147 | ~new_SUB_1596_U238;
  assign new_SUB_1596_U241 = ~P2_ADDR_REG_16_ | ~new_SUB_1596_U46;
  assign new_SUB_1596_U242 = ~new_ADD_1596_U58 | ~new_SUB_1596_U47;
  assign new_SUB_1596_U243 = ~P2_ADDR_REG_16_ | ~new_SUB_1596_U46;
  assign new_SUB_1596_U244 = ~new_ADD_1596_U58 | ~new_SUB_1596_U47;
  assign new_SUB_1596_U245 = ~new_SUB_1596_U244 | ~new_SUB_1596_U243;
  assign new_SUB_1596_U246 = ~new_SUB_1596_U80 | ~new_SUB_1596_U242 | ~new_SUB_1596_U241;
  assign new_SUB_1596_U247 = ~new_SUB_1596_U143 | ~new_SUB_1596_U245;
  assign new_SUB_1596_U248 = ~P2_ADDR_REG_15_ | ~new_SUB_1596_U43;
  assign new_SUB_1596_U249 = ~new_SUB_1596_U139 | ~new_SUB_1596_U45;
  assign new_SUB_1596_U250 = ~P2_ADDR_REG_15_ | ~new_SUB_1596_U43;
  assign new_SUB_1596_U251 = ~new_SUB_1596_U139 | ~new_SUB_1596_U45;
  assign new_SUB_1596_U252 = ~new_SUB_1596_U251 | ~new_SUB_1596_U250;
  assign new_SUB_1596_U253 = ~new_SUB_1596_U44 | ~new_SUB_1596_U249 | ~new_SUB_1596_U248;
  assign new_SUB_1596_U254 = ~new_SUB_1596_U252 | ~new_ADD_1596_U59;
  assign new_SUB_1596_U255 = ~P2_ADDR_REG_14_ | ~new_SUB_1596_U40;
  assign new_SUB_1596_U256 = ~new_SUB_1596_U135 | ~new_SUB_1596_U42;
  assign new_SUB_1596_U257 = ~P2_ADDR_REG_14_ | ~new_SUB_1596_U40;
  assign new_SUB_1596_U258 = ~new_SUB_1596_U135 | ~new_SUB_1596_U42;
  assign new_SUB_1596_U259 = ~new_SUB_1596_U258 | ~new_SUB_1596_U257;
  assign new_SUB_1596_U260 = ~new_SUB_1596_U41 | ~new_SUB_1596_U256 | ~new_SUB_1596_U255;
  assign new_SUB_1596_U261 = ~new_SUB_1596_U259 | ~new_ADD_1596_U60;
  assign new_SUB_1596_U262 = ~P2_ADDR_REG_13_ | ~new_SUB_1596_U37;
  assign new_SUB_1596_U263 = ~new_SUB_1596_U131 | ~new_SUB_1596_U39;
  assign new_SUB_1596_U264 = ~P2_ADDR_REG_13_ | ~new_SUB_1596_U37;
  assign new_SUB_1596_U265 = ~new_SUB_1596_U131 | ~new_SUB_1596_U39;
  assign new_SUB_1596_U266 = ~new_SUB_1596_U265 | ~new_SUB_1596_U264;
  assign new_SUB_1596_U267 = ~new_SUB_1596_U38 | ~new_SUB_1596_U263 | ~new_SUB_1596_U262;
  assign new_SUB_1596_U268 = ~new_SUB_1596_U266 | ~new_ADD_1596_U61;
  assign new_SUB_1596_U269 = ~P2_ADDR_REG_12_ | ~new_SUB_1596_U35;
  assign new_SUB_1596_U270 = ~new_ADD_1596_U62 | ~new_SUB_1596_U36;
  assign new_SUB_1596_U271 = ~P2_ADDR_REG_12_ | ~new_SUB_1596_U35;
  assign new_SUB_1596_U272 = ~new_ADD_1596_U62 | ~new_SUB_1596_U36;
  assign new_SUB_1596_U273 = ~new_SUB_1596_U272 | ~new_SUB_1596_U271;
  assign new_SUB_1596_U274 = ~new_SUB_1596_U81 | ~new_SUB_1596_U270 | ~new_SUB_1596_U269;
  assign new_SUB_1596_U275 = ~new_SUB_1596_U127 | ~new_SUB_1596_U273;
  assign new_SUB_1596_U276 = ~P2_ADDR_REG_11_ | ~new_SUB_1596_U33;
  assign new_SUB_1596_U277 = ~new_ADD_1596_U63 | ~new_SUB_1596_U34;
  assign new_SUB_1596_U278 = ~P2_ADDR_REG_11_ | ~new_SUB_1596_U33;
  assign new_SUB_1596_U279 = ~new_ADD_1596_U63 | ~new_SUB_1596_U34;
  assign new_SUB_1596_U280 = ~new_SUB_1596_U279 | ~new_SUB_1596_U278;
  assign new_SUB_1596_U281 = ~new_SUB_1596_U82 | ~new_SUB_1596_U277 | ~new_SUB_1596_U276;
  assign new_SUB_1596_U282 = ~new_SUB_1596_U123 | ~new_SUB_1596_U280;
  assign new_SUB_1596_U283 = ~P2_ADDR_REG_10_ | ~new_SUB_1596_U30;
  assign new_SUB_1596_U284 = ~new_SUB_1596_U119 | ~new_SUB_1596_U32;
  assign new_SUB_1596_U285 = ~P2_ADDR_REG_10_ | ~new_SUB_1596_U30;
  assign new_SUB_1596_U286 = ~new_SUB_1596_U119 | ~new_SUB_1596_U32;
  assign new_SUB_1596_U287 = ~new_SUB_1596_U286 | ~new_SUB_1596_U285;
  assign new_SUB_1596_U288 = ~new_SUB_1596_U31 | ~new_SUB_1596_U284 | ~new_SUB_1596_U283;
  assign new_SUB_1596_U289 = ~new_SUB_1596_U287 | ~new_ADD_1596_U64;
  assign new_SUB_1596_U290 = ~P2_ADDR_REG_0_ | ~new_SUB_1596_U6;
  assign new_SUB_1596_U291 = ~new_ADD_1596_U7 | ~new_SUB_1596_U7;
  assign new_ADD_1596_U6 = ~new_ADD_1596_U174 | ~new_ADD_1596_U178;
  assign new_ADD_1596_U7 = ~new_ADD_1596_U9 | ~new_ADD_1596_U179;
  assign new_ADD_1596_U8 = ~P3_ADDR_REG_0_;
  assign new_ADD_1596_U9 = ~P3_ADDR_REG_0_ | ~new_ADD_1596_U46;
  assign new_ADD_1596_U10 = ~P1_ADDR_REG_1_;
  assign new_ADD_1596_U11 = ~P3_ADDR_REG_2_;
  assign new_ADD_1596_U12 = ~P1_ADDR_REG_2_;
  assign new_ADD_1596_U13 = ~P3_ADDR_REG_3_;
  assign new_ADD_1596_U14 = ~P1_ADDR_REG_3_;
  assign new_ADD_1596_U15 = ~P3_ADDR_REG_4_;
  assign new_ADD_1596_U16 = ~P1_ADDR_REG_4_;
  assign new_ADD_1596_U17 = ~P3_ADDR_REG_5_;
  assign new_ADD_1596_U18 = ~P1_ADDR_REG_5_;
  assign new_ADD_1596_U19 = ~P3_ADDR_REG_6_;
  assign new_ADD_1596_U20 = ~P1_ADDR_REG_6_;
  assign new_ADD_1596_U21 = ~P3_ADDR_REG_7_;
  assign new_ADD_1596_U22 = ~P1_ADDR_REG_7_;
  assign new_ADD_1596_U23 = ~P3_ADDR_REG_8_;
  assign new_ADD_1596_U24 = ~P1_ADDR_REG_8_;
  assign new_ADD_1596_U25 = ~P3_ADDR_REG_9_;
  assign new_ADD_1596_U26 = ~P1_ADDR_REG_9_;
  assign new_ADD_1596_U27 = ~P3_ADDR_REG_10_;
  assign new_ADD_1596_U28 = ~P1_ADDR_REG_10_;
  assign new_ADD_1596_U29 = ~P3_ADDR_REG_11_;
  assign new_ADD_1596_U30 = ~P1_ADDR_REG_11_;
  assign new_ADD_1596_U31 = ~P3_ADDR_REG_12_;
  assign new_ADD_1596_U32 = ~P1_ADDR_REG_12_;
  assign new_ADD_1596_U33 = ~P3_ADDR_REG_13_;
  assign new_ADD_1596_U34 = ~P1_ADDR_REG_13_;
  assign new_ADD_1596_U35 = ~P3_ADDR_REG_14_;
  assign new_ADD_1596_U36 = ~P1_ADDR_REG_14_;
  assign new_ADD_1596_U37 = ~P3_ADDR_REG_15_;
  assign new_ADD_1596_U38 = ~P1_ADDR_REG_15_;
  assign new_ADD_1596_U39 = ~P3_ADDR_REG_16_;
  assign new_ADD_1596_U40 = ~P1_ADDR_REG_16_;
  assign new_ADD_1596_U41 = ~P3_ADDR_REG_17_;
  assign new_ADD_1596_U42 = ~P1_ADDR_REG_17_;
  assign new_ADD_1596_U43 = ~P3_ADDR_REG_18_;
  assign new_ADD_1596_U44 = ~P1_ADDR_REG_18_;
  assign new_ADD_1596_U45 = ~new_ADD_1596_U169 | ~new_ADD_1596_U168;
  assign new_ADD_1596_U46 = ~P1_ADDR_REG_0_;
  assign new_ADD_1596_U47 = ~new_ADD_1596_U184 | ~new_ADD_1596_U183;
  assign new_ADD_1596_U48 = ~new_ADD_1596_U189 | ~new_ADD_1596_U188;
  assign new_ADD_1596_U49 = ~new_ADD_1596_U194 | ~new_ADD_1596_U193;
  assign new_ADD_1596_U50 = ~new_ADD_1596_U199 | ~new_ADD_1596_U198;
  assign new_ADD_1596_U51 = ~new_ADD_1596_U204 | ~new_ADD_1596_U203;
  assign new_ADD_1596_U52 = ~new_ADD_1596_U209 | ~new_ADD_1596_U208;
  assign new_ADD_1596_U53 = ~new_ADD_1596_U214 | ~new_ADD_1596_U213;
  assign new_ADD_1596_U54 = ~new_ADD_1596_U219 | ~new_ADD_1596_U218;
  assign new_ADD_1596_U55 = ~new_ADD_1596_U224 | ~new_ADD_1596_U223;
  assign new_ADD_1596_U56 = ~new_ADD_1596_U234 | ~new_ADD_1596_U233;
  assign new_ADD_1596_U57 = ~new_ADD_1596_U239 | ~new_ADD_1596_U238;
  assign new_ADD_1596_U58 = ~new_ADD_1596_U244 | ~new_ADD_1596_U243;
  assign new_ADD_1596_U59 = ~new_ADD_1596_U249 | ~new_ADD_1596_U248;
  assign new_ADD_1596_U60 = ~new_ADD_1596_U254 | ~new_ADD_1596_U253;
  assign new_ADD_1596_U61 = ~new_ADD_1596_U259 | ~new_ADD_1596_U258;
  assign new_ADD_1596_U62 = ~new_ADD_1596_U264 | ~new_ADD_1596_U263;
  assign new_ADD_1596_U63 = ~new_ADD_1596_U269 | ~new_ADD_1596_U268;
  assign new_ADD_1596_U64 = ~new_ADD_1596_U274 | ~new_ADD_1596_U273;
  assign new_ADD_1596_U65 = ~new_ADD_1596_U181 | ~new_ADD_1596_U180;
  assign new_ADD_1596_U66 = ~new_ADD_1596_U186 | ~new_ADD_1596_U185;
  assign new_ADD_1596_U67 = ~new_ADD_1596_U191 | ~new_ADD_1596_U190;
  assign new_ADD_1596_U68 = ~new_ADD_1596_U196 | ~new_ADD_1596_U195;
  assign new_ADD_1596_U69 = ~new_ADD_1596_U201 | ~new_ADD_1596_U200;
  assign new_ADD_1596_U70 = ~new_ADD_1596_U206 | ~new_ADD_1596_U205;
  assign new_ADD_1596_U71 = ~new_ADD_1596_U211 | ~new_ADD_1596_U210;
  assign new_ADD_1596_U72 = ~new_ADD_1596_U216 | ~new_ADD_1596_U215;
  assign new_ADD_1596_U73 = ~new_ADD_1596_U221 | ~new_ADD_1596_U220;
  assign new_ADD_1596_U74 = ~new_ADD_1596_U231 | ~new_ADD_1596_U230;
  assign new_ADD_1596_U75 = ~new_ADD_1596_U236 | ~new_ADD_1596_U235;
  assign new_ADD_1596_U76 = ~new_ADD_1596_U241 | ~new_ADD_1596_U240;
  assign new_ADD_1596_U77 = ~new_ADD_1596_U246 | ~new_ADD_1596_U245;
  assign new_ADD_1596_U78 = ~new_ADD_1596_U251 | ~new_ADD_1596_U250;
  assign new_ADD_1596_U79 = ~new_ADD_1596_U256 | ~new_ADD_1596_U255;
  assign new_ADD_1596_U80 = ~new_ADD_1596_U261 | ~new_ADD_1596_U260;
  assign new_ADD_1596_U81 = ~new_ADD_1596_U266 | ~new_ADD_1596_U265;
  assign new_ADD_1596_U82 = ~new_ADD_1596_U271 | ~new_ADD_1596_U270;
  assign new_ADD_1596_U83 = ~new_ADD_1596_U133 | ~new_ADD_1596_U132;
  assign new_ADD_1596_U84 = ~new_ADD_1596_U129 | ~new_ADD_1596_U128;
  assign new_ADD_1596_U85 = ~new_ADD_1596_U125 | ~new_ADD_1596_U124;
  assign new_ADD_1596_U86 = ~new_ADD_1596_U121 | ~new_ADD_1596_U120;
  assign new_ADD_1596_U87 = ~new_ADD_1596_U117 | ~new_ADD_1596_U116;
  assign new_ADD_1596_U88 = ~new_ADD_1596_U113 | ~new_ADD_1596_U112;
  assign new_ADD_1596_U89 = ~new_ADD_1596_U109 | ~new_ADD_1596_U108;
  assign new_ADD_1596_U90 = ~new_ADD_1596_U105 | ~new_ADD_1596_U104;
  assign new_ADD_1596_U91 = ~P3_ADDR_REG_1_;
  assign new_ADD_1596_U92 = ~P3_ADDR_REG_19_;
  assign new_ADD_1596_U93 = ~P1_ADDR_REG_19_;
  assign new_ADD_1596_U94 = ~new_ADD_1596_U165 | ~new_ADD_1596_U164;
  assign new_ADD_1596_U95 = ~new_ADD_1596_U161 | ~new_ADD_1596_U160;
  assign new_ADD_1596_U96 = ~new_ADD_1596_U157 | ~new_ADD_1596_U156;
  assign new_ADD_1596_U97 = ~new_ADD_1596_U153 | ~new_ADD_1596_U152;
  assign new_ADD_1596_U98 = ~new_ADD_1596_U149 | ~new_ADD_1596_U148;
  assign new_ADD_1596_U99 = ~new_ADD_1596_U145 | ~new_ADD_1596_U144;
  assign new_ADD_1596_U100 = ~new_ADD_1596_U141 | ~new_ADD_1596_U140;
  assign new_ADD_1596_U101 = ~new_ADD_1596_U137 | ~new_ADD_1596_U136;
  assign new_ADD_1596_U102 = ~new_ADD_1596_U9;
  assign new_ADD_1596_U103 = ~new_ADD_1596_U102 | ~new_ADD_1596_U10;
  assign new_ADD_1596_U104 = ~new_ADD_1596_U103 | ~new_ADD_1596_U91;
  assign new_ADD_1596_U105 = ~P1_ADDR_REG_1_ | ~new_ADD_1596_U9;
  assign new_ADD_1596_U106 = ~new_ADD_1596_U90;
  assign new_ADD_1596_U107 = ~P3_ADDR_REG_2_ | ~new_ADD_1596_U12;
  assign new_ADD_1596_U108 = ~new_ADD_1596_U107 | ~new_ADD_1596_U90;
  assign new_ADD_1596_U109 = ~P1_ADDR_REG_2_ | ~new_ADD_1596_U11;
  assign new_ADD_1596_U110 = ~new_ADD_1596_U89;
  assign new_ADD_1596_U111 = ~P3_ADDR_REG_3_ | ~new_ADD_1596_U14;
  assign new_ADD_1596_U112 = ~new_ADD_1596_U111 | ~new_ADD_1596_U89;
  assign new_ADD_1596_U113 = ~P1_ADDR_REG_3_ | ~new_ADD_1596_U13;
  assign new_ADD_1596_U114 = ~new_ADD_1596_U88;
  assign new_ADD_1596_U115 = ~P3_ADDR_REG_4_ | ~new_ADD_1596_U16;
  assign new_ADD_1596_U116 = ~new_ADD_1596_U115 | ~new_ADD_1596_U88;
  assign new_ADD_1596_U117 = ~P1_ADDR_REG_4_ | ~new_ADD_1596_U15;
  assign new_ADD_1596_U118 = ~new_ADD_1596_U87;
  assign new_ADD_1596_U119 = ~P3_ADDR_REG_5_ | ~new_ADD_1596_U18;
  assign new_ADD_1596_U120 = ~new_ADD_1596_U119 | ~new_ADD_1596_U87;
  assign new_ADD_1596_U121 = ~P1_ADDR_REG_5_ | ~new_ADD_1596_U17;
  assign new_ADD_1596_U122 = ~new_ADD_1596_U86;
  assign new_ADD_1596_U123 = ~P3_ADDR_REG_6_ | ~new_ADD_1596_U20;
  assign new_ADD_1596_U124 = ~new_ADD_1596_U123 | ~new_ADD_1596_U86;
  assign new_ADD_1596_U125 = ~P1_ADDR_REG_6_ | ~new_ADD_1596_U19;
  assign new_ADD_1596_U126 = ~new_ADD_1596_U85;
  assign new_ADD_1596_U127 = ~P3_ADDR_REG_7_ | ~new_ADD_1596_U22;
  assign new_ADD_1596_U128 = ~new_ADD_1596_U127 | ~new_ADD_1596_U85;
  assign new_ADD_1596_U129 = ~P1_ADDR_REG_7_ | ~new_ADD_1596_U21;
  assign new_ADD_1596_U130 = ~new_ADD_1596_U84;
  assign new_ADD_1596_U131 = ~P3_ADDR_REG_8_ | ~new_ADD_1596_U24;
  assign new_ADD_1596_U132 = ~new_ADD_1596_U131 | ~new_ADD_1596_U84;
  assign new_ADD_1596_U133 = ~P1_ADDR_REG_8_ | ~new_ADD_1596_U23;
  assign new_ADD_1596_U134 = ~new_ADD_1596_U83;
  assign new_ADD_1596_U135 = ~P3_ADDR_REG_9_ | ~new_ADD_1596_U26;
  assign new_ADD_1596_U136 = ~new_ADD_1596_U135 | ~new_ADD_1596_U83;
  assign new_ADD_1596_U137 = ~P1_ADDR_REG_9_ | ~new_ADD_1596_U25;
  assign new_ADD_1596_U138 = ~new_ADD_1596_U101;
  assign new_ADD_1596_U139 = ~P3_ADDR_REG_10_ | ~new_ADD_1596_U28;
  assign new_ADD_1596_U140 = ~new_ADD_1596_U139 | ~new_ADD_1596_U101;
  assign new_ADD_1596_U141 = ~P1_ADDR_REG_10_ | ~new_ADD_1596_U27;
  assign new_ADD_1596_U142 = ~new_ADD_1596_U100;
  assign new_ADD_1596_U143 = ~P3_ADDR_REG_11_ | ~new_ADD_1596_U30;
  assign new_ADD_1596_U144 = ~new_ADD_1596_U143 | ~new_ADD_1596_U100;
  assign new_ADD_1596_U145 = ~P1_ADDR_REG_11_ | ~new_ADD_1596_U29;
  assign new_ADD_1596_U146 = ~new_ADD_1596_U99;
  assign new_ADD_1596_U147 = ~P3_ADDR_REG_12_ | ~new_ADD_1596_U32;
  assign new_ADD_1596_U148 = ~new_ADD_1596_U147 | ~new_ADD_1596_U99;
  assign new_ADD_1596_U149 = ~P1_ADDR_REG_12_ | ~new_ADD_1596_U31;
  assign new_ADD_1596_U150 = ~new_ADD_1596_U98;
  assign new_ADD_1596_U151 = ~P3_ADDR_REG_13_ | ~new_ADD_1596_U34;
  assign new_ADD_1596_U152 = ~new_ADD_1596_U151 | ~new_ADD_1596_U98;
  assign new_ADD_1596_U153 = ~P1_ADDR_REG_13_ | ~new_ADD_1596_U33;
  assign new_ADD_1596_U154 = ~new_ADD_1596_U97;
  assign new_ADD_1596_U155 = ~P3_ADDR_REG_14_ | ~new_ADD_1596_U36;
  assign new_ADD_1596_U156 = ~new_ADD_1596_U155 | ~new_ADD_1596_U97;
  assign new_ADD_1596_U157 = ~P1_ADDR_REG_14_ | ~new_ADD_1596_U35;
  assign new_ADD_1596_U158 = ~new_ADD_1596_U96;
  assign new_ADD_1596_U159 = ~P3_ADDR_REG_15_ | ~new_ADD_1596_U38;
  assign new_ADD_1596_U160 = ~new_ADD_1596_U159 | ~new_ADD_1596_U96;
  assign new_ADD_1596_U161 = ~P1_ADDR_REG_15_ | ~new_ADD_1596_U37;
  assign new_ADD_1596_U162 = ~new_ADD_1596_U95;
  assign new_ADD_1596_U163 = ~P3_ADDR_REG_16_ | ~new_ADD_1596_U40;
  assign new_ADD_1596_U164 = ~new_ADD_1596_U163 | ~new_ADD_1596_U95;
  assign new_ADD_1596_U165 = ~P1_ADDR_REG_16_ | ~new_ADD_1596_U39;
  assign new_ADD_1596_U166 = ~new_ADD_1596_U94;
  assign new_ADD_1596_U167 = ~P3_ADDR_REG_17_ | ~new_ADD_1596_U42;
  assign new_ADD_1596_U168 = ~new_ADD_1596_U167 | ~new_ADD_1596_U94;
  assign new_ADD_1596_U169 = ~P1_ADDR_REG_17_ | ~new_ADD_1596_U41;
  assign new_ADD_1596_U170 = ~new_ADD_1596_U45;
  assign new_ADD_1596_U171 = ~P1_ADDR_REG_18_ | ~new_ADD_1596_U43;
  assign new_ADD_1596_U172 = ~new_ADD_1596_U170 | ~new_ADD_1596_U171;
  assign new_ADD_1596_U173 = ~P3_ADDR_REG_18_ | ~new_ADD_1596_U44;
  assign new_ADD_1596_U174 = ~new_ADD_1596_U172 | ~new_ADD_1596_U173 | ~new_ADD_1596_U229;
  assign new_ADD_1596_U175 = ~P3_ADDR_REG_18_ | ~new_ADD_1596_U44;
  assign new_ADD_1596_U176 = ~new_ADD_1596_U175 | ~new_ADD_1596_U45;
  assign new_ADD_1596_U177 = ~P1_ADDR_REG_18_ | ~new_ADD_1596_U43;
  assign new_ADD_1596_U178 = ~new_ADD_1596_U176 | ~new_ADD_1596_U177 | ~new_ADD_1596_U226 | ~new_ADD_1596_U225;
  assign new_ADD_1596_U179 = ~P1_ADDR_REG_0_ | ~new_ADD_1596_U8;
  assign new_ADD_1596_U180 = ~P3_ADDR_REG_9_ | ~new_ADD_1596_U26;
  assign new_ADD_1596_U181 = ~P1_ADDR_REG_9_ | ~new_ADD_1596_U25;
  assign new_ADD_1596_U182 = ~new_ADD_1596_U65;
  assign new_ADD_1596_U183 = ~new_ADD_1596_U134 | ~new_ADD_1596_U182;
  assign new_ADD_1596_U184 = ~new_ADD_1596_U65 | ~new_ADD_1596_U83;
  assign new_ADD_1596_U185 = ~P3_ADDR_REG_8_ | ~new_ADD_1596_U24;
  assign new_ADD_1596_U186 = ~P1_ADDR_REG_8_ | ~new_ADD_1596_U23;
  assign new_ADD_1596_U187 = ~new_ADD_1596_U66;
  assign new_ADD_1596_U188 = ~new_ADD_1596_U130 | ~new_ADD_1596_U187;
  assign new_ADD_1596_U189 = ~new_ADD_1596_U66 | ~new_ADD_1596_U84;
  assign new_ADD_1596_U190 = ~P3_ADDR_REG_7_ | ~new_ADD_1596_U22;
  assign new_ADD_1596_U191 = ~P1_ADDR_REG_7_ | ~new_ADD_1596_U21;
  assign new_ADD_1596_U192 = ~new_ADD_1596_U67;
  assign new_ADD_1596_U193 = ~new_ADD_1596_U126 | ~new_ADD_1596_U192;
  assign new_ADD_1596_U194 = ~new_ADD_1596_U67 | ~new_ADD_1596_U85;
  assign new_ADD_1596_U195 = ~P3_ADDR_REG_6_ | ~new_ADD_1596_U20;
  assign new_ADD_1596_U196 = ~P1_ADDR_REG_6_ | ~new_ADD_1596_U19;
  assign new_ADD_1596_U197 = ~new_ADD_1596_U68;
  assign new_ADD_1596_U198 = ~new_ADD_1596_U122 | ~new_ADD_1596_U197;
  assign new_ADD_1596_U199 = ~new_ADD_1596_U68 | ~new_ADD_1596_U86;
  assign new_ADD_1596_U200 = ~P3_ADDR_REG_5_ | ~new_ADD_1596_U18;
  assign new_ADD_1596_U201 = ~P1_ADDR_REG_5_ | ~new_ADD_1596_U17;
  assign new_ADD_1596_U202 = ~new_ADD_1596_U69;
  assign new_ADD_1596_U203 = ~new_ADD_1596_U118 | ~new_ADD_1596_U202;
  assign new_ADD_1596_U204 = ~new_ADD_1596_U69 | ~new_ADD_1596_U87;
  assign new_ADD_1596_U205 = ~P3_ADDR_REG_4_ | ~new_ADD_1596_U16;
  assign new_ADD_1596_U206 = ~P1_ADDR_REG_4_ | ~new_ADD_1596_U15;
  assign new_ADD_1596_U207 = ~new_ADD_1596_U70;
  assign new_ADD_1596_U208 = ~new_ADD_1596_U114 | ~new_ADD_1596_U207;
  assign new_ADD_1596_U209 = ~new_ADD_1596_U70 | ~new_ADD_1596_U88;
  assign new_ADD_1596_U210 = ~P3_ADDR_REG_3_ | ~new_ADD_1596_U14;
  assign new_ADD_1596_U211 = ~P1_ADDR_REG_3_ | ~new_ADD_1596_U13;
  assign new_ADD_1596_U212 = ~new_ADD_1596_U71;
  assign new_ADD_1596_U213 = ~new_ADD_1596_U110 | ~new_ADD_1596_U212;
  assign new_ADD_1596_U214 = ~new_ADD_1596_U71 | ~new_ADD_1596_U89;
  assign new_ADD_1596_U215 = ~P3_ADDR_REG_2_ | ~new_ADD_1596_U12;
  assign new_ADD_1596_U216 = ~P1_ADDR_REG_2_ | ~new_ADD_1596_U11;
  assign new_ADD_1596_U217 = ~new_ADD_1596_U72;
  assign new_ADD_1596_U218 = ~new_ADD_1596_U106 | ~new_ADD_1596_U217;
  assign new_ADD_1596_U219 = ~new_ADD_1596_U72 | ~new_ADD_1596_U90;
  assign new_ADD_1596_U220 = ~P3_ADDR_REG_1_ | ~new_ADD_1596_U10;
  assign new_ADD_1596_U221 = ~P1_ADDR_REG_1_ | ~new_ADD_1596_U91;
  assign new_ADD_1596_U222 = ~new_ADD_1596_U73;
  assign new_ADD_1596_U223 = ~new_ADD_1596_U222 | ~new_ADD_1596_U102;
  assign new_ADD_1596_U224 = ~new_ADD_1596_U73 | ~new_ADD_1596_U9;
  assign new_ADD_1596_U225 = ~P3_ADDR_REG_19_ | ~new_ADD_1596_U93;
  assign new_ADD_1596_U226 = ~P1_ADDR_REG_19_ | ~new_ADD_1596_U92;
  assign new_ADD_1596_U227 = ~P3_ADDR_REG_19_ | ~new_ADD_1596_U93;
  assign new_ADD_1596_U228 = ~P1_ADDR_REG_19_ | ~new_ADD_1596_U92;
  assign new_ADD_1596_U229 = ~new_ADD_1596_U228 | ~new_ADD_1596_U227;
  assign new_ADD_1596_U230 = ~P3_ADDR_REG_18_ | ~new_ADD_1596_U44;
  assign new_ADD_1596_U231 = ~P1_ADDR_REG_18_ | ~new_ADD_1596_U43;
  assign new_ADD_1596_U232 = ~new_ADD_1596_U74;
  assign new_ADD_1596_U233 = ~new_ADD_1596_U232 | ~new_ADD_1596_U170;
  assign new_ADD_1596_U234 = ~new_ADD_1596_U74 | ~new_ADD_1596_U45;
  assign new_ADD_1596_U235 = ~P3_ADDR_REG_17_ | ~new_ADD_1596_U42;
  assign new_ADD_1596_U236 = ~P1_ADDR_REG_17_ | ~new_ADD_1596_U41;
  assign new_ADD_1596_U237 = ~new_ADD_1596_U75;
  assign new_ADD_1596_U238 = ~new_ADD_1596_U166 | ~new_ADD_1596_U237;
  assign new_ADD_1596_U239 = ~new_ADD_1596_U75 | ~new_ADD_1596_U94;
  assign new_ADD_1596_U240 = ~P3_ADDR_REG_16_ | ~new_ADD_1596_U40;
  assign new_ADD_1596_U241 = ~P1_ADDR_REG_16_ | ~new_ADD_1596_U39;
  assign new_ADD_1596_U242 = ~new_ADD_1596_U76;
  assign new_ADD_1596_U243 = ~new_ADD_1596_U162 | ~new_ADD_1596_U242;
  assign new_ADD_1596_U244 = ~new_ADD_1596_U76 | ~new_ADD_1596_U95;
  assign new_ADD_1596_U245 = ~P3_ADDR_REG_15_ | ~new_ADD_1596_U38;
  assign new_ADD_1596_U246 = ~P1_ADDR_REG_15_ | ~new_ADD_1596_U37;
  assign new_ADD_1596_U247 = ~new_ADD_1596_U77;
  assign new_ADD_1596_U248 = ~new_ADD_1596_U158 | ~new_ADD_1596_U247;
  assign new_ADD_1596_U249 = ~new_ADD_1596_U77 | ~new_ADD_1596_U96;
  assign new_ADD_1596_U250 = ~P3_ADDR_REG_14_ | ~new_ADD_1596_U36;
  assign new_ADD_1596_U251 = ~P1_ADDR_REG_14_ | ~new_ADD_1596_U35;
  assign new_ADD_1596_U252 = ~new_ADD_1596_U78;
  assign new_ADD_1596_U253 = ~new_ADD_1596_U154 | ~new_ADD_1596_U252;
  assign new_ADD_1596_U254 = ~new_ADD_1596_U78 | ~new_ADD_1596_U97;
  assign new_ADD_1596_U255 = ~P3_ADDR_REG_13_ | ~new_ADD_1596_U34;
  assign new_ADD_1596_U256 = ~P1_ADDR_REG_13_ | ~new_ADD_1596_U33;
  assign new_ADD_1596_U257 = ~new_ADD_1596_U79;
  assign new_ADD_1596_U258 = ~new_ADD_1596_U150 | ~new_ADD_1596_U257;
  assign new_ADD_1596_U259 = ~new_ADD_1596_U79 | ~new_ADD_1596_U98;
  assign new_ADD_1596_U260 = ~P3_ADDR_REG_12_ | ~new_ADD_1596_U32;
  assign new_ADD_1596_U261 = ~P1_ADDR_REG_12_ | ~new_ADD_1596_U31;
  assign new_ADD_1596_U262 = ~new_ADD_1596_U80;
  assign new_ADD_1596_U263 = ~new_ADD_1596_U146 | ~new_ADD_1596_U262;
  assign new_ADD_1596_U264 = ~new_ADD_1596_U80 | ~new_ADD_1596_U99;
  assign new_ADD_1596_U265 = ~P3_ADDR_REG_11_ | ~new_ADD_1596_U30;
  assign new_ADD_1596_U266 = ~P1_ADDR_REG_11_ | ~new_ADD_1596_U29;
  assign new_ADD_1596_U267 = ~new_ADD_1596_U81;
  assign new_ADD_1596_U268 = ~new_ADD_1596_U142 | ~new_ADD_1596_U267;
  assign new_ADD_1596_U269 = ~new_ADD_1596_U81 | ~new_ADD_1596_U100;
  assign new_ADD_1596_U270 = ~P3_ADDR_REG_10_ | ~new_ADD_1596_U28;
  assign new_ADD_1596_U271 = ~P1_ADDR_REG_10_ | ~new_ADD_1596_U27;
  assign new_ADD_1596_U272 = ~new_ADD_1596_U82;
  assign new_ADD_1596_U273 = ~new_ADD_1596_U138 | ~new_ADD_1596_U272;
  assign new_ADD_1596_U274 = ~new_ADD_1596_U82 | ~new_ADD_1596_U101;
  assign new_LT_1601_21_U6 = ~P2_ADDR_REG_19_;
  assign new_P1_ADD_99_U4 = ~P1_REG3_REG_3_;
  assign new_P1_ADD_99_U5 = new_P1_ADD_99_U102 & P1_REG3_REG_28_ & P1_REG3_REG_27_;
  assign new_P1_ADD_99_U6 = ~P1_REG3_REG_4_;
  assign new_P1_ADD_99_U7 = ~P1_REG3_REG_4_ | ~P1_REG3_REG_3_;
  assign new_P1_ADD_99_U8 = ~P1_REG3_REG_5_;
  assign new_P1_ADD_99_U9 = ~P1_REG3_REG_5_ | ~new_P1_ADD_99_U80;
  assign new_P1_ADD_99_U10 = ~P1_REG3_REG_6_;
  assign new_P1_ADD_99_U11 = ~P1_REG3_REG_6_ | ~new_P1_ADD_99_U81;
  assign new_P1_ADD_99_U12 = ~P1_REG3_REG_7_;
  assign new_P1_ADD_99_U13 = ~P1_REG3_REG_7_ | ~new_P1_ADD_99_U82;
  assign new_P1_ADD_99_U14 = ~P1_REG3_REG_8_;
  assign new_P1_ADD_99_U15 = ~P1_REG3_REG_9_;
  assign new_P1_ADD_99_U16 = ~P1_REG3_REG_8_ | ~new_P1_ADD_99_U83;
  assign new_P1_ADD_99_U17 = ~new_P1_ADD_99_U84 | ~P1_REG3_REG_9_;
  assign new_P1_ADD_99_U18 = ~P1_REG3_REG_10_;
  assign new_P1_ADD_99_U19 = ~P1_REG3_REG_10_ | ~new_P1_ADD_99_U85;
  assign new_P1_ADD_99_U20 = ~P1_REG3_REG_11_;
  assign new_P1_ADD_99_U21 = ~P1_REG3_REG_11_ | ~new_P1_ADD_99_U86;
  assign new_P1_ADD_99_U22 = ~P1_REG3_REG_12_;
  assign new_P1_ADD_99_U23 = ~P1_REG3_REG_12_ | ~new_P1_ADD_99_U87;
  assign new_P1_ADD_99_U24 = ~P1_REG3_REG_13_;
  assign new_P1_ADD_99_U25 = ~P1_REG3_REG_13_ | ~new_P1_ADD_99_U88;
  assign new_P1_ADD_99_U26 = ~P1_REG3_REG_14_;
  assign new_P1_ADD_99_U27 = ~P1_REG3_REG_14_ | ~new_P1_ADD_99_U89;
  assign new_P1_ADD_99_U28 = ~P1_REG3_REG_15_;
  assign new_P1_ADD_99_U29 = ~P1_REG3_REG_15_ | ~new_P1_ADD_99_U90;
  assign new_P1_ADD_99_U30 = ~P1_REG3_REG_16_;
  assign new_P1_ADD_99_U31 = ~P1_REG3_REG_16_ | ~new_P1_ADD_99_U91;
  assign new_P1_ADD_99_U32 = ~P1_REG3_REG_17_;
  assign new_P1_ADD_99_U33 = ~P1_REG3_REG_17_ | ~new_P1_ADD_99_U92;
  assign new_P1_ADD_99_U34 = ~P1_REG3_REG_18_;
  assign new_P1_ADD_99_U35 = ~P1_REG3_REG_18_ | ~new_P1_ADD_99_U93;
  assign new_P1_ADD_99_U36 = ~P1_REG3_REG_19_;
  assign new_P1_ADD_99_U37 = ~P1_REG3_REG_19_ | ~new_P1_ADD_99_U94;
  assign new_P1_ADD_99_U38 = ~P1_REG3_REG_20_;
  assign new_P1_ADD_99_U39 = ~P1_REG3_REG_20_ | ~new_P1_ADD_99_U95;
  assign new_P1_ADD_99_U40 = ~P1_REG3_REG_21_;
  assign new_P1_ADD_99_U41 = ~P1_REG3_REG_21_ | ~new_P1_ADD_99_U96;
  assign new_P1_ADD_99_U42 = ~P1_REG3_REG_22_;
  assign new_P1_ADD_99_U43 = ~P1_REG3_REG_22_ | ~new_P1_ADD_99_U97;
  assign new_P1_ADD_99_U44 = ~P1_REG3_REG_23_;
  assign new_P1_ADD_99_U45 = ~P1_REG3_REG_23_ | ~new_P1_ADD_99_U98;
  assign new_P1_ADD_99_U46 = ~P1_REG3_REG_24_;
  assign new_P1_ADD_99_U47 = ~P1_REG3_REG_24_ | ~new_P1_ADD_99_U99;
  assign new_P1_ADD_99_U48 = ~P1_REG3_REG_25_;
  assign new_P1_ADD_99_U49 = ~P1_REG3_REG_25_ | ~new_P1_ADD_99_U100;
  assign new_P1_ADD_99_U50 = ~P1_REG3_REG_26_;
  assign new_P1_ADD_99_U51 = ~P1_REG3_REG_26_ | ~new_P1_ADD_99_U101;
  assign new_P1_ADD_99_U52 = ~P1_REG3_REG_28_;
  assign new_P1_ADD_99_U53 = ~P1_REG3_REG_27_;
  assign new_P1_ADD_99_U54 = ~new_P1_ADD_99_U105 | ~new_P1_ADD_99_U104;
  assign new_P1_ADD_99_U55 = ~new_P1_ADD_99_U107 | ~new_P1_ADD_99_U106;
  assign new_P1_ADD_99_U56 = ~new_P1_ADD_99_U109 | ~new_P1_ADD_99_U108;
  assign new_P1_ADD_99_U57 = ~new_P1_ADD_99_U111 | ~new_P1_ADD_99_U110;
  assign new_P1_ADD_99_U58 = ~new_P1_ADD_99_U113 | ~new_P1_ADD_99_U112;
  assign new_P1_ADD_99_U59 = ~new_P1_ADD_99_U115 | ~new_P1_ADD_99_U114;
  assign new_P1_ADD_99_U60 = ~new_P1_ADD_99_U117 | ~new_P1_ADD_99_U116;
  assign new_P1_ADD_99_U61 = ~new_P1_ADD_99_U119 | ~new_P1_ADD_99_U118;
  assign new_P1_ADD_99_U62 = ~new_P1_ADD_99_U121 | ~new_P1_ADD_99_U120;
  assign new_P1_ADD_99_U63 = ~new_P1_ADD_99_U123 | ~new_P1_ADD_99_U122;
  assign new_P1_ADD_99_U64 = ~new_P1_ADD_99_U125 | ~new_P1_ADD_99_U124;
  assign new_P1_ADD_99_U65 = ~new_P1_ADD_99_U127 | ~new_P1_ADD_99_U126;
  assign new_P1_ADD_99_U66 = ~new_P1_ADD_99_U129 | ~new_P1_ADD_99_U128;
  assign new_P1_ADD_99_U67 = ~new_P1_ADD_99_U131 | ~new_P1_ADD_99_U130;
  assign new_P1_ADD_99_U68 = ~new_P1_ADD_99_U133 | ~new_P1_ADD_99_U132;
  assign new_P1_ADD_99_U69 = ~new_P1_ADD_99_U135 | ~new_P1_ADD_99_U134;
  assign new_P1_ADD_99_U70 = ~new_P1_ADD_99_U137 | ~new_P1_ADD_99_U136;
  assign new_P1_ADD_99_U71 = ~new_P1_ADD_99_U139 | ~new_P1_ADD_99_U138;
  assign new_P1_ADD_99_U72 = ~new_P1_ADD_99_U141 | ~new_P1_ADD_99_U140;
  assign new_P1_ADD_99_U73 = ~new_P1_ADD_99_U143 | ~new_P1_ADD_99_U142;
  assign new_P1_ADD_99_U74 = ~new_P1_ADD_99_U145 | ~new_P1_ADD_99_U144;
  assign new_P1_ADD_99_U75 = ~new_P1_ADD_99_U147 | ~new_P1_ADD_99_U146;
  assign new_P1_ADD_99_U76 = ~new_P1_ADD_99_U149 | ~new_P1_ADD_99_U148;
  assign new_P1_ADD_99_U77 = ~new_P1_ADD_99_U151 | ~new_P1_ADD_99_U150;
  assign new_P1_ADD_99_U78 = ~new_P1_ADD_99_U153 | ~new_P1_ADD_99_U152;
  assign new_P1_ADD_99_U79 = ~P1_REG3_REG_27_ | ~new_P1_ADD_99_U102;
  assign new_P1_ADD_99_U80 = ~new_P1_ADD_99_U7;
  assign new_P1_ADD_99_U81 = ~new_P1_ADD_99_U9;
  assign new_P1_ADD_99_U82 = ~new_P1_ADD_99_U11;
  assign new_P1_ADD_99_U83 = ~new_P1_ADD_99_U13;
  assign new_P1_ADD_99_U84 = ~new_P1_ADD_99_U16;
  assign new_P1_ADD_99_U85 = ~new_P1_ADD_99_U17;
  assign new_P1_ADD_99_U86 = ~new_P1_ADD_99_U19;
  assign new_P1_ADD_99_U87 = ~new_P1_ADD_99_U21;
  assign new_P1_ADD_99_U88 = ~new_P1_ADD_99_U23;
  assign new_P1_ADD_99_U89 = ~new_P1_ADD_99_U25;
  assign new_P1_ADD_99_U90 = ~new_P1_ADD_99_U27;
  assign new_P1_ADD_99_U91 = ~new_P1_ADD_99_U29;
  assign new_P1_ADD_99_U92 = ~new_P1_ADD_99_U31;
  assign new_P1_ADD_99_U93 = ~new_P1_ADD_99_U33;
  assign new_P1_ADD_99_U94 = ~new_P1_ADD_99_U35;
  assign new_P1_ADD_99_U95 = ~new_P1_ADD_99_U37;
  assign new_P1_ADD_99_U96 = ~new_P1_ADD_99_U39;
  assign new_P1_ADD_99_U97 = ~new_P1_ADD_99_U41;
  assign new_P1_ADD_99_U98 = ~new_P1_ADD_99_U43;
  assign new_P1_ADD_99_U99 = ~new_P1_ADD_99_U45;
  assign new_P1_ADD_99_U100 = ~new_P1_ADD_99_U47;
  assign new_P1_ADD_99_U101 = ~new_P1_ADD_99_U49;
  assign new_P1_ADD_99_U102 = ~new_P1_ADD_99_U51;
  assign new_P1_ADD_99_U103 = ~new_P1_ADD_99_U79;
  assign new_P1_ADD_99_U104 = ~P1_REG3_REG_9_ | ~new_P1_ADD_99_U16;
  assign new_P1_ADD_99_U105 = ~new_P1_ADD_99_U84 | ~new_P1_ADD_99_U15;
  assign new_P1_ADD_99_U106 = ~P1_REG3_REG_8_ | ~new_P1_ADD_99_U13;
  assign new_P1_ADD_99_U107 = ~new_P1_ADD_99_U83 | ~new_P1_ADD_99_U14;
  assign new_P1_ADD_99_U108 = ~P1_REG3_REG_7_ | ~new_P1_ADD_99_U11;
  assign new_P1_ADD_99_U109 = ~new_P1_ADD_99_U82 | ~new_P1_ADD_99_U12;
  assign new_P1_ADD_99_U110 = ~P1_REG3_REG_6_ | ~new_P1_ADD_99_U9;
  assign new_P1_ADD_99_U111 = ~new_P1_ADD_99_U81 | ~new_P1_ADD_99_U10;
  assign new_P1_ADD_99_U112 = ~P1_REG3_REG_5_ | ~new_P1_ADD_99_U7;
  assign new_P1_ADD_99_U113 = ~new_P1_ADD_99_U80 | ~new_P1_ADD_99_U8;
  assign new_P1_ADD_99_U114 = ~P1_REG3_REG_4_ | ~new_P1_ADD_99_U4;
  assign new_P1_ADD_99_U115 = ~P1_REG3_REG_3_ | ~new_P1_ADD_99_U6;
  assign new_P1_ADD_99_U116 = ~P1_REG3_REG_28_ | ~new_P1_ADD_99_U79;
  assign new_P1_ADD_99_U117 = ~new_P1_ADD_99_U103 | ~new_P1_ADD_99_U52;
  assign new_P1_ADD_99_U118 = ~P1_REG3_REG_27_ | ~new_P1_ADD_99_U51;
  assign new_P1_ADD_99_U119 = ~new_P1_ADD_99_U102 | ~new_P1_ADD_99_U53;
  assign new_P1_ADD_99_U120 = ~P1_REG3_REG_26_ | ~new_P1_ADD_99_U49;
  assign new_P1_ADD_99_U121 = ~new_P1_ADD_99_U101 | ~new_P1_ADD_99_U50;
  assign new_P1_ADD_99_U122 = ~P1_REG3_REG_25_ | ~new_P1_ADD_99_U47;
  assign new_P1_ADD_99_U123 = ~new_P1_ADD_99_U100 | ~new_P1_ADD_99_U48;
  assign new_P1_ADD_99_U124 = ~P1_REG3_REG_24_ | ~new_P1_ADD_99_U45;
  assign new_P1_ADD_99_U125 = ~new_P1_ADD_99_U99 | ~new_P1_ADD_99_U46;
  assign new_P1_ADD_99_U126 = ~P1_REG3_REG_23_ | ~new_P1_ADD_99_U43;
  assign new_P1_ADD_99_U127 = ~new_P1_ADD_99_U98 | ~new_P1_ADD_99_U44;
  assign new_P1_ADD_99_U128 = ~P1_REG3_REG_22_ | ~new_P1_ADD_99_U41;
  assign new_P1_ADD_99_U129 = ~new_P1_ADD_99_U97 | ~new_P1_ADD_99_U42;
  assign new_P1_ADD_99_U130 = ~P1_REG3_REG_21_ | ~new_P1_ADD_99_U39;
  assign new_P1_ADD_99_U131 = ~new_P1_ADD_99_U96 | ~new_P1_ADD_99_U40;
  assign new_P1_ADD_99_U132 = ~P1_REG3_REG_20_ | ~new_P1_ADD_99_U37;
  assign new_P1_ADD_99_U133 = ~new_P1_ADD_99_U95 | ~new_P1_ADD_99_U38;
  assign new_P1_ADD_99_U134 = ~P1_REG3_REG_19_ | ~new_P1_ADD_99_U35;
  assign new_P1_ADD_99_U135 = ~new_P1_ADD_99_U94 | ~new_P1_ADD_99_U36;
  assign new_P1_ADD_99_U136 = ~P1_REG3_REG_18_ | ~new_P1_ADD_99_U33;
  assign new_P1_ADD_99_U137 = ~new_P1_ADD_99_U93 | ~new_P1_ADD_99_U34;
  assign new_P1_ADD_99_U138 = ~P1_REG3_REG_17_ | ~new_P1_ADD_99_U31;
  assign new_P1_ADD_99_U139 = ~new_P1_ADD_99_U92 | ~new_P1_ADD_99_U32;
  assign new_P1_ADD_99_U140 = ~P1_REG3_REG_16_ | ~new_P1_ADD_99_U29;
  assign new_P1_ADD_99_U141 = ~new_P1_ADD_99_U91 | ~new_P1_ADD_99_U30;
  assign new_P1_ADD_99_U142 = ~P1_REG3_REG_15_ | ~new_P1_ADD_99_U27;
  assign new_P1_ADD_99_U143 = ~new_P1_ADD_99_U90 | ~new_P1_ADD_99_U28;
  assign new_P1_ADD_99_U144 = ~P1_REG3_REG_14_ | ~new_P1_ADD_99_U25;
  assign new_P1_ADD_99_U145 = ~new_P1_ADD_99_U89 | ~new_P1_ADD_99_U26;
  assign new_P1_ADD_99_U146 = ~P1_REG3_REG_13_ | ~new_P1_ADD_99_U23;
  assign new_P1_ADD_99_U147 = ~new_P1_ADD_99_U88 | ~new_P1_ADD_99_U24;
  assign new_P1_ADD_99_U148 = ~P1_REG3_REG_12_ | ~new_P1_ADD_99_U21;
  assign new_P1_ADD_99_U149 = ~new_P1_ADD_99_U87 | ~new_P1_ADD_99_U22;
  assign new_P1_ADD_99_U150 = ~P1_REG3_REG_11_ | ~new_P1_ADD_99_U19;
  assign new_P1_ADD_99_U151 = ~new_P1_ADD_99_U86 | ~new_P1_ADD_99_U20;
  assign new_P1_ADD_99_U152 = ~P1_REG3_REG_10_ | ~new_P1_ADD_99_U17;
  assign new_P1_ADD_99_U153 = ~new_P1_ADD_99_U85 | ~new_P1_ADD_99_U18;
  assign new_P1_R1105_U4 = new_P1_R1105_U95 & new_P1_R1105_U94;
  assign new_P1_R1105_U5 = new_P1_R1105_U96 & new_P1_R1105_U97;
  assign new_P1_R1105_U6 = new_P1_R1105_U113 & new_P1_R1105_U112;
  assign new_P1_R1105_U7 = new_P1_R1105_U155 & new_P1_R1105_U154;
  assign new_P1_R1105_U8 = new_P1_R1105_U164 & new_P1_R1105_U163;
  assign new_P1_R1105_U9 = new_P1_R1105_U182 & new_P1_R1105_U181;
  assign new_P1_R1105_U10 = new_P1_R1105_U218 & new_P1_R1105_U215;
  assign new_P1_R1105_U11 = new_P1_R1105_U211 & new_P1_R1105_U208;
  assign new_P1_R1105_U12 = new_P1_R1105_U202 & new_P1_R1105_U199;
  assign new_P1_R1105_U13 = new_P1_R1105_U196 & new_P1_R1105_U192;
  assign new_P1_R1105_U14 = new_P1_R1105_U151 & new_P1_R1105_U148;
  assign new_P1_R1105_U15 = new_P1_R1105_U143 & new_P1_R1105_U140;
  assign new_P1_R1105_U16 = new_P1_R1105_U129 & new_P1_R1105_U126;
  assign new_P1_R1105_U17 = ~P1_REG2_REG_6_;
  assign new_P1_R1105_U18 = ~new_P1_U3475;
  assign new_P1_R1105_U19 = ~new_P1_U3478;
  assign new_P1_R1105_U20 = ~new_P1_U3475 | ~P1_REG2_REG_6_;
  assign new_P1_R1105_U21 = ~P1_REG2_REG_7_;
  assign new_P1_R1105_U22 = ~P1_REG2_REG_4_;
  assign new_P1_R1105_U23 = ~new_P1_U3469;
  assign new_P1_R1105_U24 = ~new_P1_U3472;
  assign new_P1_R1105_U25 = ~P1_REG2_REG_2_;
  assign new_P1_R1105_U26 = ~new_P1_U3463;
  assign new_P1_R1105_U27 = ~P1_REG2_REG_0_;
  assign new_P1_R1105_U28 = ~new_P1_U3454;
  assign new_P1_R1105_U29 = ~new_P1_U3454 | ~P1_REG2_REG_0_;
  assign new_P1_R1105_U30 = ~P1_REG2_REG_3_;
  assign new_P1_R1105_U31 = ~new_P1_U3466;
  assign new_P1_R1105_U32 = ~new_P1_U3469 | ~P1_REG2_REG_4_;
  assign new_P1_R1105_U33 = ~P1_REG2_REG_5_;
  assign new_P1_R1105_U34 = ~P1_REG2_REG_8_;
  assign new_P1_R1105_U35 = ~new_P1_U3481;
  assign new_P1_R1105_U36 = ~new_P1_U3484;
  assign new_P1_R1105_U37 = ~P1_REG2_REG_9_;
  assign new_P1_R1105_U38 = ~new_P1_R1105_U49 | ~new_P1_R1105_U121;
  assign new_P1_R1105_U39 = ~new_P1_R1105_U109 | ~new_P1_R1105_U110 | ~new_P1_R1105_U108;
  assign new_P1_R1105_U40 = ~new_P1_R1105_U98 | ~new_P1_R1105_U99;
  assign new_P1_R1105_U41 = ~P1_REG2_REG_1_ | ~new_P1_U3460;
  assign new_P1_R1105_U42 = ~new_P1_R1105_U135 | ~new_P1_R1105_U136 | ~new_P1_R1105_U134;
  assign new_P1_R1105_U43 = ~new_P1_R1105_U132 | ~new_P1_R1105_U131;
  assign new_P1_R1105_U44 = ~P1_REG2_REG_16_;
  assign new_P1_R1105_U45 = ~new_P1_U3505;
  assign new_P1_R1105_U46 = ~new_P1_U3508;
  assign new_P1_R1105_U47 = ~new_P1_U3505 | ~P1_REG2_REG_16_;
  assign new_P1_R1105_U48 = ~P1_REG2_REG_17_;
  assign new_P1_R1105_U49 = ~new_P1_U3481 | ~P1_REG2_REG_8_;
  assign new_P1_R1105_U50 = ~P1_REG2_REG_10_;
  assign new_P1_R1105_U51 = ~new_P1_U3487;
  assign new_P1_R1105_U52 = ~P1_REG2_REG_12_;
  assign new_P1_R1105_U53 = ~new_P1_U3493;
  assign new_P1_R1105_U54 = ~P1_REG2_REG_11_;
  assign new_P1_R1105_U55 = ~new_P1_U3490;
  assign new_P1_R1105_U56 = ~new_P1_U3490 | ~P1_REG2_REG_11_;
  assign new_P1_R1105_U57 = ~P1_REG2_REG_13_;
  assign new_P1_R1105_U58 = ~new_P1_U3496;
  assign new_P1_R1105_U59 = ~P1_REG2_REG_14_;
  assign new_P1_R1105_U60 = ~new_P1_U3499;
  assign new_P1_R1105_U61 = ~P1_REG2_REG_15_;
  assign new_P1_R1105_U62 = ~new_P1_U3502;
  assign new_P1_R1105_U63 = ~P1_REG2_REG_18_;
  assign new_P1_R1105_U64 = ~new_P1_U3511;
  assign new_P1_R1105_U65 = ~new_P1_R1105_U187 | ~new_P1_R1105_U186 | ~new_P1_R1105_U185;
  assign new_P1_R1105_U66 = ~new_P1_R1105_U179 | ~new_P1_R1105_U178;
  assign new_P1_R1105_U67 = ~new_P1_R1105_U56 | ~new_P1_R1105_U204;
  assign new_P1_R1105_U68 = ~new_P1_R1105_U259 | ~new_P1_R1105_U258;
  assign new_P1_R1105_U69 = ~new_P1_R1105_U308 | ~new_P1_R1105_U307;
  assign new_P1_R1105_U70 = ~new_P1_R1105_U231 | ~new_P1_R1105_U230;
  assign new_P1_R1105_U71 = ~new_P1_R1105_U236 | ~new_P1_R1105_U235;
  assign new_P1_R1105_U72 = ~new_P1_R1105_U243 | ~new_P1_R1105_U242;
  assign new_P1_R1105_U73 = ~new_P1_R1105_U250 | ~new_P1_R1105_U249;
  assign new_P1_R1105_U74 = ~new_P1_R1105_U255 | ~new_P1_R1105_U254;
  assign new_P1_R1105_U75 = ~new_P1_R1105_U271 | ~new_P1_R1105_U270;
  assign new_P1_R1105_U76 = ~new_P1_R1105_U278 | ~new_P1_R1105_U277;
  assign new_P1_R1105_U77 = ~new_P1_R1105_U285 | ~new_P1_R1105_U284;
  assign new_P1_R1105_U78 = ~new_P1_R1105_U292 | ~new_P1_R1105_U291;
  assign new_P1_R1105_U79 = ~new_P1_R1105_U299 | ~new_P1_R1105_U298;
  assign new_P1_R1105_U80 = ~new_P1_R1105_U304 | ~new_P1_R1105_U303;
  assign new_P1_R1105_U81 = ~new_P1_R1105_U118 | ~new_P1_R1105_U117 | ~new_P1_R1105_U116;
  assign new_P1_R1105_U82 = ~new_P1_R1105_U133 | ~new_P1_R1105_U145;
  assign new_P1_R1105_U83 = ~new_P1_R1105_U41 | ~new_P1_R1105_U152;
  assign new_P1_R1105_U84 = ~new_P1_U3452;
  assign new_P1_R1105_U85 = ~P1_REG2_REG_19_;
  assign new_P1_R1105_U86 = ~new_P1_R1105_U175 | ~new_P1_R1105_U174;
  assign new_P1_R1105_U87 = ~new_P1_R1105_U171 | ~new_P1_R1105_U170;
  assign new_P1_R1105_U88 = ~new_P1_R1105_U161 | ~new_P1_R1105_U160;
  assign new_P1_R1105_U89 = ~new_P1_R1105_U32;
  assign new_P1_R1105_U90 = ~P1_REG2_REG_9_ | ~new_P1_U3484;
  assign new_P1_R1105_U91 = ~new_P1_U3493 | ~P1_REG2_REG_12_;
  assign new_P1_R1105_U92 = ~new_P1_R1105_U56;
  assign new_P1_R1105_U93 = ~new_P1_R1105_U49;
  assign new_P1_R1105_U94 = new_P1_U3472 | P1_REG2_REG_5_;
  assign new_P1_R1105_U95 = new_P1_U3469 | P1_REG2_REG_4_;
  assign new_P1_R1105_U96 = P1_REG2_REG_3_ | new_P1_U3466;
  assign new_P1_R1105_U97 = P1_REG2_REG_2_ | new_P1_U3463;
  assign new_P1_R1105_U98 = ~new_P1_R1105_U29;
  assign new_P1_R1105_U99 = P1_REG2_REG_1_ | new_P1_U3460;
  assign new_P1_R1105_U100 = ~new_P1_R1105_U40;
  assign new_P1_R1105_U101 = ~new_P1_R1105_U41;
  assign new_P1_R1105_U102 = ~new_P1_R1105_U40 | ~new_P1_R1105_U41;
  assign new_P1_R1105_U103 = ~new_P1_R1105_U96 | ~P1_REG2_REG_2_ | ~new_P1_U3463;
  assign new_P1_R1105_U104 = ~new_P1_R1105_U5 | ~new_P1_R1105_U102;
  assign new_P1_R1105_U105 = ~new_P1_U3466 | ~P1_REG2_REG_3_;
  assign new_P1_R1105_U106 = ~new_P1_R1105_U104 | ~new_P1_R1105_U105 | ~new_P1_R1105_U103;
  assign new_P1_R1105_U107 = ~new_P1_R1105_U33 | ~new_P1_R1105_U32;
  assign new_P1_R1105_U108 = ~new_P1_U3472 | ~new_P1_R1105_U107;
  assign new_P1_R1105_U109 = ~new_P1_R1105_U4 | ~new_P1_R1105_U106;
  assign new_P1_R1105_U110 = ~P1_REG2_REG_5_ | ~new_P1_R1105_U89;
  assign new_P1_R1105_U111 = ~new_P1_R1105_U39;
  assign new_P1_R1105_U112 = new_P1_U3478 | P1_REG2_REG_7_;
  assign new_P1_R1105_U113 = new_P1_U3475 | P1_REG2_REG_6_;
  assign new_P1_R1105_U114 = ~new_P1_R1105_U20;
  assign new_P1_R1105_U115 = ~new_P1_R1105_U21 | ~new_P1_R1105_U20;
  assign new_P1_R1105_U116 = ~new_P1_U3478 | ~new_P1_R1105_U115;
  assign new_P1_R1105_U117 = ~P1_REG2_REG_7_ | ~new_P1_R1105_U114;
  assign new_P1_R1105_U118 = ~new_P1_R1105_U6 | ~new_P1_R1105_U39;
  assign new_P1_R1105_U119 = ~new_P1_R1105_U81;
  assign new_P1_R1105_U120 = P1_REG2_REG_8_ | new_P1_U3481;
  assign new_P1_R1105_U121 = ~new_P1_R1105_U120 | ~new_P1_R1105_U81;
  assign new_P1_R1105_U122 = ~new_P1_R1105_U38;
  assign new_P1_R1105_U123 = new_P1_U3484 | P1_REG2_REG_9_;
  assign new_P1_R1105_U124 = P1_REG2_REG_6_ | new_P1_U3475;
  assign new_P1_R1105_U125 = ~new_P1_R1105_U124 | ~new_P1_R1105_U39;
  assign new_P1_R1105_U126 = ~new_P1_R1105_U125 | ~new_P1_R1105_U20 | ~new_P1_R1105_U238 | ~new_P1_R1105_U237;
  assign new_P1_R1105_U127 = ~new_P1_R1105_U111 | ~new_P1_R1105_U20;
  assign new_P1_R1105_U128 = ~P1_REG2_REG_7_ | ~new_P1_U3478;
  assign new_P1_R1105_U129 = ~new_P1_R1105_U127 | ~new_P1_R1105_U128 | ~new_P1_R1105_U6;
  assign new_P1_R1105_U130 = new_P1_U3475 | P1_REG2_REG_6_;
  assign new_P1_R1105_U131 = ~new_P1_R1105_U101 | ~new_P1_R1105_U97;
  assign new_P1_R1105_U132 = ~new_P1_U3463 | ~P1_REG2_REG_2_;
  assign new_P1_R1105_U133 = ~new_P1_R1105_U43;
  assign new_P1_R1105_U134 = ~new_P1_R1105_U100 | ~new_P1_R1105_U5;
  assign new_P1_R1105_U135 = ~new_P1_R1105_U43 | ~new_P1_R1105_U96;
  assign new_P1_R1105_U136 = ~new_P1_U3466 | ~P1_REG2_REG_3_;
  assign new_P1_R1105_U137 = ~new_P1_R1105_U42;
  assign new_P1_R1105_U138 = P1_REG2_REG_4_ | new_P1_U3469;
  assign new_P1_R1105_U139 = ~new_P1_R1105_U138 | ~new_P1_R1105_U42;
  assign new_P1_R1105_U140 = ~new_P1_R1105_U139 | ~new_P1_R1105_U32 | ~new_P1_R1105_U245 | ~new_P1_R1105_U244;
  assign new_P1_R1105_U141 = ~new_P1_R1105_U137 | ~new_P1_R1105_U32;
  assign new_P1_R1105_U142 = ~P1_REG2_REG_5_ | ~new_P1_U3472;
  assign new_P1_R1105_U143 = ~new_P1_R1105_U141 | ~new_P1_R1105_U142 | ~new_P1_R1105_U4;
  assign new_P1_R1105_U144 = new_P1_U3469 | P1_REG2_REG_4_;
  assign new_P1_R1105_U145 = ~new_P1_R1105_U100 | ~new_P1_R1105_U97;
  assign new_P1_R1105_U146 = ~new_P1_R1105_U82;
  assign new_P1_R1105_U147 = ~new_P1_U3466 | ~P1_REG2_REG_3_;
  assign new_P1_R1105_U148 = ~new_P1_R1105_U256 | ~new_P1_R1105_U257 | ~new_P1_R1105_U41 | ~new_P1_R1105_U40;
  assign new_P1_R1105_U149 = ~new_P1_R1105_U41 | ~new_P1_R1105_U40;
  assign new_P1_R1105_U150 = ~new_P1_U3463 | ~P1_REG2_REG_2_;
  assign new_P1_R1105_U151 = ~new_P1_R1105_U149 | ~new_P1_R1105_U150 | ~new_P1_R1105_U97;
  assign new_P1_R1105_U152 = P1_REG2_REG_1_ | new_P1_U3460;
  assign new_P1_R1105_U153 = ~new_P1_R1105_U83;
  assign new_P1_R1105_U154 = new_P1_U3484 | P1_REG2_REG_9_;
  assign new_P1_R1105_U155 = new_P1_U3487 | P1_REG2_REG_10_;
  assign new_P1_R1105_U156 = ~new_P1_R1105_U93 | ~new_P1_R1105_U7;
  assign new_P1_R1105_U157 = ~new_P1_U3487 | ~P1_REG2_REG_10_;
  assign new_P1_R1105_U158 = ~new_P1_R1105_U156 | ~new_P1_R1105_U157 | ~new_P1_R1105_U90;
  assign new_P1_R1105_U159 = P1_REG2_REG_10_ | new_P1_U3487;
  assign new_P1_R1105_U160 = ~new_P1_R1105_U81 | ~new_P1_R1105_U120 | ~new_P1_R1105_U7;
  assign new_P1_R1105_U161 = ~new_P1_R1105_U159 | ~new_P1_R1105_U158;
  assign new_P1_R1105_U162 = ~new_P1_R1105_U88;
  assign new_P1_R1105_U163 = new_P1_U3496 | P1_REG2_REG_13_;
  assign new_P1_R1105_U164 = new_P1_U3493 | P1_REG2_REG_12_;
  assign new_P1_R1105_U165 = ~new_P1_R1105_U92 | ~new_P1_R1105_U8;
  assign new_P1_R1105_U166 = ~new_P1_U3496 | ~P1_REG2_REG_13_;
  assign new_P1_R1105_U167 = ~new_P1_R1105_U165 | ~new_P1_R1105_U166 | ~new_P1_R1105_U91;
  assign new_P1_R1105_U168 = P1_REG2_REG_11_ | new_P1_U3490;
  assign new_P1_R1105_U169 = P1_REG2_REG_13_ | new_P1_U3496;
  assign new_P1_R1105_U170 = ~new_P1_R1105_U88 | ~new_P1_R1105_U168 | ~new_P1_R1105_U8;
  assign new_P1_R1105_U171 = ~new_P1_R1105_U169 | ~new_P1_R1105_U167;
  assign new_P1_R1105_U172 = ~new_P1_R1105_U87;
  assign new_P1_R1105_U173 = P1_REG2_REG_14_ | new_P1_U3499;
  assign new_P1_R1105_U174 = ~new_P1_R1105_U173 | ~new_P1_R1105_U87;
  assign new_P1_R1105_U175 = ~new_P1_U3499 | ~P1_REG2_REG_14_;
  assign new_P1_R1105_U176 = ~new_P1_R1105_U86;
  assign new_P1_R1105_U177 = P1_REG2_REG_15_ | new_P1_U3502;
  assign new_P1_R1105_U178 = ~new_P1_R1105_U177 | ~new_P1_R1105_U86;
  assign new_P1_R1105_U179 = ~new_P1_U3502 | ~P1_REG2_REG_15_;
  assign new_P1_R1105_U180 = ~new_P1_R1105_U66;
  assign new_P1_R1105_U181 = new_P1_U3508 | P1_REG2_REG_17_;
  assign new_P1_R1105_U182 = new_P1_U3505 | P1_REG2_REG_16_;
  assign new_P1_R1105_U183 = ~new_P1_R1105_U47;
  assign new_P1_R1105_U184 = ~new_P1_R1105_U48 | ~new_P1_R1105_U47;
  assign new_P1_R1105_U185 = ~new_P1_U3508 | ~new_P1_R1105_U184;
  assign new_P1_R1105_U186 = ~P1_REG2_REG_17_ | ~new_P1_R1105_U183;
  assign new_P1_R1105_U187 = ~new_P1_R1105_U9 | ~new_P1_R1105_U66;
  assign new_P1_R1105_U188 = ~new_P1_R1105_U65;
  assign new_P1_R1105_U189 = P1_REG2_REG_18_ | new_P1_U3511;
  assign new_P1_R1105_U190 = ~new_P1_R1105_U189 | ~new_P1_R1105_U65;
  assign new_P1_R1105_U191 = ~new_P1_U3511 | ~P1_REG2_REG_18_;
  assign new_P1_R1105_U192 = ~new_P1_R1105_U190 | ~new_P1_R1105_U191 | ~new_P1_R1105_U261 | ~new_P1_R1105_U260;
  assign new_P1_R1105_U193 = ~new_P1_U3511 | ~P1_REG2_REG_18_;
  assign new_P1_R1105_U194 = ~new_P1_R1105_U188 | ~new_P1_R1105_U193;
  assign new_P1_R1105_U195 = new_P1_U3511 | P1_REG2_REG_18_;
  assign new_P1_R1105_U196 = ~new_P1_R1105_U194 | ~new_P1_R1105_U195 | ~new_P1_R1105_U264;
  assign new_P1_R1105_U197 = P1_REG2_REG_16_ | new_P1_U3505;
  assign new_P1_R1105_U198 = ~new_P1_R1105_U197 | ~new_P1_R1105_U66;
  assign new_P1_R1105_U199 = ~new_P1_R1105_U198 | ~new_P1_R1105_U47 | ~new_P1_R1105_U273 | ~new_P1_R1105_U272;
  assign new_P1_R1105_U200 = ~new_P1_R1105_U180 | ~new_P1_R1105_U47;
  assign new_P1_R1105_U201 = ~P1_REG2_REG_17_ | ~new_P1_U3508;
  assign new_P1_R1105_U202 = ~new_P1_R1105_U200 | ~new_P1_R1105_U201 | ~new_P1_R1105_U9;
  assign new_P1_R1105_U203 = new_P1_U3505 | P1_REG2_REG_16_;
  assign new_P1_R1105_U204 = ~new_P1_R1105_U168 | ~new_P1_R1105_U88;
  assign new_P1_R1105_U205 = ~new_P1_R1105_U67;
  assign new_P1_R1105_U206 = P1_REG2_REG_12_ | new_P1_U3493;
  assign new_P1_R1105_U207 = ~new_P1_R1105_U206 | ~new_P1_R1105_U67;
  assign new_P1_R1105_U208 = ~new_P1_R1105_U207 | ~new_P1_R1105_U91 | ~new_P1_R1105_U294 | ~new_P1_R1105_U293;
  assign new_P1_R1105_U209 = ~new_P1_R1105_U205 | ~new_P1_R1105_U91;
  assign new_P1_R1105_U210 = ~new_P1_U3496 | ~P1_REG2_REG_13_;
  assign new_P1_R1105_U211 = ~new_P1_R1105_U209 | ~new_P1_R1105_U210 | ~new_P1_R1105_U8;
  assign new_P1_R1105_U212 = new_P1_U3493 | P1_REG2_REG_12_;
  assign new_P1_R1105_U213 = P1_REG2_REG_9_ | new_P1_U3484;
  assign new_P1_R1105_U214 = ~new_P1_R1105_U213 | ~new_P1_R1105_U38;
  assign new_P1_R1105_U215 = ~new_P1_R1105_U214 | ~new_P1_R1105_U90 | ~new_P1_R1105_U306 | ~new_P1_R1105_U305;
  assign new_P1_R1105_U216 = ~new_P1_R1105_U122 | ~new_P1_R1105_U90;
  assign new_P1_R1105_U217 = ~new_P1_U3487 | ~P1_REG2_REG_10_;
  assign new_P1_R1105_U218 = ~new_P1_R1105_U216 | ~new_P1_R1105_U217 | ~new_P1_R1105_U7;
  assign new_P1_R1105_U219 = ~new_P1_R1105_U123 | ~new_P1_R1105_U90;
  assign new_P1_R1105_U220 = ~new_P1_R1105_U120 | ~new_P1_R1105_U49;
  assign new_P1_R1105_U221 = ~new_P1_R1105_U130 | ~new_P1_R1105_U20;
  assign new_P1_R1105_U222 = ~new_P1_R1105_U144 | ~new_P1_R1105_U32;
  assign new_P1_R1105_U223 = ~new_P1_R1105_U147 | ~new_P1_R1105_U96;
  assign new_P1_R1105_U224 = ~new_P1_R1105_U203 | ~new_P1_R1105_U47;
  assign new_P1_R1105_U225 = ~new_P1_R1105_U212 | ~new_P1_R1105_U91;
  assign new_P1_R1105_U226 = ~new_P1_R1105_U168 | ~new_P1_R1105_U56;
  assign new_P1_R1105_U227 = ~new_P1_U3484 | ~new_P1_R1105_U37;
  assign new_P1_R1105_U228 = ~P1_REG2_REG_9_ | ~new_P1_R1105_U36;
  assign new_P1_R1105_U229 = ~new_P1_R1105_U228 | ~new_P1_R1105_U227;
  assign new_P1_R1105_U230 = ~new_P1_R1105_U219 | ~new_P1_R1105_U38;
  assign new_P1_R1105_U231 = ~new_P1_R1105_U229 | ~new_P1_R1105_U122;
  assign new_P1_R1105_U232 = ~new_P1_U3481 | ~new_P1_R1105_U34;
  assign new_P1_R1105_U233 = ~P1_REG2_REG_8_ | ~new_P1_R1105_U35;
  assign new_P1_R1105_U234 = ~new_P1_R1105_U233 | ~new_P1_R1105_U232;
  assign new_P1_R1105_U235 = ~new_P1_R1105_U220 | ~new_P1_R1105_U81;
  assign new_P1_R1105_U236 = ~new_P1_R1105_U119 | ~new_P1_R1105_U234;
  assign new_P1_R1105_U237 = ~new_P1_U3478 | ~new_P1_R1105_U21;
  assign new_P1_R1105_U238 = ~P1_REG2_REG_7_ | ~new_P1_R1105_U19;
  assign new_P1_R1105_U239 = ~new_P1_U3475 | ~new_P1_R1105_U17;
  assign new_P1_R1105_U240 = ~P1_REG2_REG_6_ | ~new_P1_R1105_U18;
  assign new_P1_R1105_U241 = ~new_P1_R1105_U240 | ~new_P1_R1105_U239;
  assign new_P1_R1105_U242 = ~new_P1_R1105_U221 | ~new_P1_R1105_U39;
  assign new_P1_R1105_U243 = ~new_P1_R1105_U241 | ~new_P1_R1105_U111;
  assign new_P1_R1105_U244 = ~new_P1_U3472 | ~new_P1_R1105_U33;
  assign new_P1_R1105_U245 = ~P1_REG2_REG_5_ | ~new_P1_R1105_U24;
  assign new_P1_R1105_U246 = ~new_P1_U3469 | ~new_P1_R1105_U22;
  assign new_P1_R1105_U247 = ~P1_REG2_REG_4_ | ~new_P1_R1105_U23;
  assign new_P1_R1105_U248 = ~new_P1_R1105_U247 | ~new_P1_R1105_U246;
  assign new_P1_R1105_U249 = ~new_P1_R1105_U222 | ~new_P1_R1105_U42;
  assign new_P1_R1105_U250 = ~new_P1_R1105_U248 | ~new_P1_R1105_U137;
  assign new_P1_R1105_U251 = ~new_P1_U3466 | ~new_P1_R1105_U30;
  assign new_P1_R1105_U252 = ~P1_REG2_REG_3_ | ~new_P1_R1105_U31;
  assign new_P1_R1105_U253 = ~new_P1_R1105_U252 | ~new_P1_R1105_U251;
  assign new_P1_R1105_U254 = ~new_P1_R1105_U223 | ~new_P1_R1105_U82;
  assign new_P1_R1105_U255 = ~new_P1_R1105_U146 | ~new_P1_R1105_U253;
  assign new_P1_R1105_U256 = ~new_P1_U3463 | ~new_P1_R1105_U25;
  assign new_P1_R1105_U257 = ~P1_REG2_REG_2_ | ~new_P1_R1105_U26;
  assign new_P1_R1105_U258 = ~new_P1_R1105_U98 | ~new_P1_R1105_U83;
  assign new_P1_R1105_U259 = ~new_P1_R1105_U153 | ~new_P1_R1105_U29;
  assign new_P1_R1105_U260 = ~new_P1_U3452 | ~new_P1_R1105_U85;
  assign new_P1_R1105_U261 = ~P1_REG2_REG_19_ | ~new_P1_R1105_U84;
  assign new_P1_R1105_U262 = ~new_P1_U3452 | ~new_P1_R1105_U85;
  assign new_P1_R1105_U263 = ~P1_REG2_REG_19_ | ~new_P1_R1105_U84;
  assign new_P1_R1105_U264 = ~new_P1_R1105_U263 | ~new_P1_R1105_U262;
  assign new_P1_R1105_U265 = ~new_P1_U3511 | ~new_P1_R1105_U63;
  assign new_P1_R1105_U266 = ~P1_REG2_REG_18_ | ~new_P1_R1105_U64;
  assign new_P1_R1105_U267 = ~new_P1_U3511 | ~new_P1_R1105_U63;
  assign new_P1_R1105_U268 = ~P1_REG2_REG_18_ | ~new_P1_R1105_U64;
  assign new_P1_R1105_U269 = ~new_P1_R1105_U268 | ~new_P1_R1105_U267;
  assign new_P1_R1105_U270 = ~new_P1_R1105_U65 | ~new_P1_R1105_U266 | ~new_P1_R1105_U265;
  assign new_P1_R1105_U271 = ~new_P1_R1105_U269 | ~new_P1_R1105_U188;
  assign new_P1_R1105_U272 = ~new_P1_U3508 | ~new_P1_R1105_U48;
  assign new_P1_R1105_U273 = ~P1_REG2_REG_17_ | ~new_P1_R1105_U46;
  assign new_P1_R1105_U274 = ~new_P1_U3505 | ~new_P1_R1105_U44;
  assign new_P1_R1105_U275 = ~P1_REG2_REG_16_ | ~new_P1_R1105_U45;
  assign new_P1_R1105_U276 = ~new_P1_R1105_U275 | ~new_P1_R1105_U274;
  assign new_P1_R1105_U277 = ~new_P1_R1105_U224 | ~new_P1_R1105_U66;
  assign new_P1_R1105_U278 = ~new_P1_R1105_U276 | ~new_P1_R1105_U180;
  assign new_P1_R1105_U279 = ~new_P1_U3502 | ~new_P1_R1105_U61;
  assign new_P1_R1105_U280 = ~P1_REG2_REG_15_ | ~new_P1_R1105_U62;
  assign new_P1_R1105_U281 = ~new_P1_U3502 | ~new_P1_R1105_U61;
  assign new_P1_R1105_U282 = ~P1_REG2_REG_15_ | ~new_P1_R1105_U62;
  assign new_P1_R1105_U283 = ~new_P1_R1105_U282 | ~new_P1_R1105_U281;
  assign new_P1_R1105_U284 = ~new_P1_R1105_U86 | ~new_P1_R1105_U280 | ~new_P1_R1105_U279;
  assign new_P1_R1105_U285 = ~new_P1_R1105_U176 | ~new_P1_R1105_U283;
  assign new_P1_R1105_U286 = ~new_P1_U3499 | ~new_P1_R1105_U59;
  assign new_P1_R1105_U287 = ~P1_REG2_REG_14_ | ~new_P1_R1105_U60;
  assign new_P1_R1105_U288 = ~new_P1_U3499 | ~new_P1_R1105_U59;
  assign new_P1_R1105_U289 = ~P1_REG2_REG_14_ | ~new_P1_R1105_U60;
  assign new_P1_R1105_U290 = ~new_P1_R1105_U289 | ~new_P1_R1105_U288;
  assign new_P1_R1105_U291 = ~new_P1_R1105_U87 | ~new_P1_R1105_U287 | ~new_P1_R1105_U286;
  assign new_P1_R1105_U292 = ~new_P1_R1105_U172 | ~new_P1_R1105_U290;
  assign new_P1_R1105_U293 = ~new_P1_U3496 | ~new_P1_R1105_U57;
  assign new_P1_R1105_U294 = ~P1_REG2_REG_13_ | ~new_P1_R1105_U58;
  assign new_P1_R1105_U295 = ~new_P1_U3493 | ~new_P1_R1105_U52;
  assign new_P1_R1105_U296 = ~P1_REG2_REG_12_ | ~new_P1_R1105_U53;
  assign new_P1_R1105_U297 = ~new_P1_R1105_U296 | ~new_P1_R1105_U295;
  assign new_P1_R1105_U298 = ~new_P1_R1105_U225 | ~new_P1_R1105_U67;
  assign new_P1_R1105_U299 = ~new_P1_R1105_U297 | ~new_P1_R1105_U205;
  assign new_P1_R1105_U300 = ~new_P1_U3490 | ~new_P1_R1105_U54;
  assign new_P1_R1105_U301 = ~P1_REG2_REG_11_ | ~new_P1_R1105_U55;
  assign new_P1_R1105_U302 = ~new_P1_R1105_U301 | ~new_P1_R1105_U300;
  assign new_P1_R1105_U303 = ~new_P1_R1105_U226 | ~new_P1_R1105_U88;
  assign new_P1_R1105_U304 = ~new_P1_R1105_U162 | ~new_P1_R1105_U302;
  assign new_P1_R1105_U305 = ~new_P1_U3487 | ~new_P1_R1105_U50;
  assign new_P1_R1105_U306 = ~P1_REG2_REG_10_ | ~new_P1_R1105_U51;
  assign new_P1_R1105_U307 = ~new_P1_U3454 | ~new_P1_R1105_U27;
  assign new_P1_R1105_U308 = ~P1_REG2_REG_0_ | ~new_P1_R1105_U28;
  assign new_P1_SUB_88_U6 = new_P1_SUB_88_U227 & new_P1_SUB_88_U38;
  assign new_P1_SUB_88_U7 = new_P1_SUB_88_U225 & new_P1_SUB_88_U192;
  assign new_P1_SUB_88_U8 = new_P1_SUB_88_U224 & new_P1_SUB_88_U35;
  assign new_P1_SUB_88_U9 = new_P1_SUB_88_U223 & new_P1_SUB_88_U36;
  assign new_P1_SUB_88_U10 = new_P1_SUB_88_U221 & new_P1_SUB_88_U195;
  assign new_P1_SUB_88_U11 = new_P1_SUB_88_U220 & new_P1_SUB_88_U34;
  assign new_P1_SUB_88_U12 = new_P1_SUB_88_U219 & new_P1_SUB_88_U197;
  assign new_P1_SUB_88_U13 = new_P1_SUB_88_U217 & new_P1_SUB_88_U198;
  assign new_P1_SUB_88_U14 = new_P1_SUB_88_U216 & new_P1_SUB_88_U172;
  assign new_P1_SUB_88_U15 = new_P1_SUB_88_U215 & new_P1_SUB_88_U200;
  assign new_P1_SUB_88_U16 = new_P1_SUB_88_U213 & new_P1_SUB_88_U201;
  assign new_P1_SUB_88_U17 = new_P1_SUB_88_U212 & new_P1_SUB_88_U169;
  assign new_P1_SUB_88_U18 = new_P1_SUB_88_U211 & new_P1_SUB_88_U167;
  assign new_P1_SUB_88_U19 = new_P1_SUB_88_U209 & new_P1_SUB_88_U204;
  assign new_P1_SUB_88_U20 = new_P1_SUB_88_U208 & new_P1_SUB_88_U33;
  assign new_P1_SUB_88_U21 = new_P1_SUB_88_U207 & new_P1_SUB_88_U27;
  assign new_P1_SUB_88_U22 = new_P1_SUB_88_U190 & new_P1_SUB_88_U180;
  assign new_P1_SUB_88_U23 = new_P1_SUB_88_U189 & new_P1_SUB_88_U29;
  assign new_P1_SUB_88_U24 = new_P1_SUB_88_U188 & new_P1_SUB_88_U30;
  assign new_P1_SUB_88_U25 = new_P1_SUB_88_U186 & new_P1_SUB_88_U183;
  assign new_P1_SUB_88_U26 = new_P1_SUB_88_U185 & new_P1_SUB_88_U28;
  assign new_P1_SUB_88_U27 = P1_IR_REG_2_ | P1_IR_REG_1_ | P1_IR_REG_0_;
  assign new_P1_SUB_88_U28 = ~new_P1_SUB_88_U43 | ~new_P1_SUB_88_U44 | ~new_P1_SUB_88_U230;
  assign new_P1_SUB_88_U29 = ~new_P1_SUB_88_U45 | ~new_P1_SUB_88_U230;
  assign new_P1_SUB_88_U30 = ~new_P1_SUB_88_U46 | ~new_P1_SUB_88_U181;
  assign new_P1_SUB_88_U31 = ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U32 = ~P1_IR_REG_3_;
  assign new_P1_SUB_88_U33 = ~new_P1_SUB_88_U56 | ~new_P1_SUB_88_U51;
  assign new_P1_SUB_88_U34 = ~new_P1_SUB_88_U127 | ~new_P1_SUB_88_U128 | ~new_P1_SUB_88_U130 | ~new_P1_SUB_88_U129;
  assign new_P1_SUB_88_U35 = ~new_P1_SUB_88_U156 | ~new_P1_SUB_88_U184;
  assign new_P1_SUB_88_U36 = ~new_P1_SUB_88_U157 | ~new_P1_SUB_88_U193;
  assign new_P1_SUB_88_U37 = ~P1_IR_REG_15_;
  assign new_P1_SUB_88_U38 = ~new_P1_SUB_88_U158 | ~new_P1_SUB_88_U184;
  assign new_P1_SUB_88_U39 = ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U40 = ~new_P1_SUB_88_U247 | ~new_P1_SUB_88_U246;
  assign new_P1_SUB_88_U41 = ~new_P1_SUB_88_U237 | ~new_P1_SUB_88_U236;
  assign new_P1_SUB_88_U42 = ~new_P1_SUB_88_U241 | ~new_P1_SUB_88_U240;
  assign new_P1_SUB_88_U43 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U44 = ~P1_IR_REG_7_ & ~P1_IR_REG_8_;
  assign new_P1_SUB_88_U45 = ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U46 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_;
  assign new_P1_SUB_88_U47 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U48 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_ & ~P1_IR_REG_15_;
  assign new_P1_SUB_88_U49 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_88_U50 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_88_U51 = new_P1_SUB_88_U47 & new_P1_SUB_88_U48 & new_P1_SUB_88_U50 & new_P1_SUB_88_U49;
  assign new_P1_SUB_88_U52 = ~P1_IR_REG_26_ & ~P1_IR_REG_25_ & ~P1_IR_REG_23_ & ~P1_IR_REG_24_;
  assign new_P1_SUB_88_U53 = ~P1_IR_REG_2_ & ~P1_IR_REG_29_ & ~P1_IR_REG_27_ & ~P1_IR_REG_28_;
  assign new_P1_SUB_88_U54 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U55 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U56 = new_P1_SUB_88_U52 & new_P1_SUB_88_U53 & new_P1_SUB_88_U55 & new_P1_SUB_88_U54;
  assign new_P1_SUB_88_U57 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U58 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_ & ~P1_IR_REG_15_;
  assign new_P1_SUB_88_U59 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_88_U60 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_88_U61 = new_P1_SUB_88_U57 & new_P1_SUB_88_U58 & new_P1_SUB_88_U60 & new_P1_SUB_88_U59;
  assign new_P1_SUB_88_U62 = ~P1_IR_REG_26_ & ~P1_IR_REG_25_ & ~P1_IR_REG_23_ & ~P1_IR_REG_24_;
  assign new_P1_SUB_88_U63 = ~P1_IR_REG_28_ & ~P1_IR_REG_2_ & ~P1_IR_REG_27_;
  assign new_P1_SUB_88_U64 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U65 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U66 = new_P1_SUB_88_U62 & new_P1_SUB_88_U63 & new_P1_SUB_88_U65 & new_P1_SUB_88_U64;
  assign new_P1_SUB_88_U67 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U68 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U69 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_88_U70 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_88_U71 = new_P1_SUB_88_U67 & new_P1_SUB_88_U68 & new_P1_SUB_88_U70 & new_P1_SUB_88_U69;
  assign new_P1_SUB_88_U72 = ~P1_IR_REG_25_ & ~P1_IR_REG_24_ & ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_88_U73 = ~P1_IR_REG_27_ & ~P1_IR_REG_2_ & ~P1_IR_REG_26_;
  assign new_P1_SUB_88_U74 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U75 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U76 = new_P1_SUB_88_U72 & new_P1_SUB_88_U73 & new_P1_SUB_88_U75 & new_P1_SUB_88_U74;
  assign new_P1_SUB_88_U77 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U78 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U79 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_88_U80 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_88_U81 = new_P1_SUB_88_U77 & new_P1_SUB_88_U78 & new_P1_SUB_88_U80 & new_P1_SUB_88_U79;
  assign new_P1_SUB_88_U82 = ~P1_IR_REG_25_ & ~P1_IR_REG_24_ & ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_88_U83 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_26_;
  assign new_P1_SUB_88_U84 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U85 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U86 = new_P1_SUB_88_U82 & new_P1_SUB_88_U83 & new_P1_SUB_88_U85 & new_P1_SUB_88_U84;
  assign new_P1_SUB_88_U87 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U88 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U89 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_88_U90 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_88_U91 = new_P1_SUB_88_U87 & new_P1_SUB_88_U88 & new_P1_SUB_88_U90 & new_P1_SUB_88_U89;
  assign new_P1_SUB_88_U92 = ~P1_IR_REG_25_ & ~P1_IR_REG_24_ & ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_88_U93 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_26_;
  assign new_P1_SUB_88_U94 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U95 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U96 = new_P1_SUB_88_U92 & new_P1_SUB_88_U93 & new_P1_SUB_88_U95 & new_P1_SUB_88_U94;
  assign new_P1_SUB_88_U97 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U98 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U99 = ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_;
  assign new_P1_SUB_88_U100 = ~P1_IR_REG_0_ & ~P1_IR_REG_20_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_88_U101 = new_P1_SUB_88_U97 & new_P1_SUB_88_U98 & new_P1_SUB_88_U100 & new_P1_SUB_88_U99;
  assign new_P1_SUB_88_U102 = ~P1_IR_REG_24_ & ~P1_IR_REG_23_ & ~P1_IR_REG_21_ & ~P1_IR_REG_22_;
  assign new_P1_SUB_88_U103 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_25_;
  assign new_P1_SUB_88_U104 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U105 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U106 = new_P1_SUB_88_U102 & new_P1_SUB_88_U103 & new_P1_SUB_88_U105 & new_P1_SUB_88_U104;
  assign new_P1_SUB_88_U107 = ~P1_IR_REG_13_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U108 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U109 = ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_17_;
  assign new_P1_SUB_88_U110 = ~P1_IR_REG_0_ & ~P1_IR_REG_20_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_88_U111 = new_P1_SUB_88_U107 & new_P1_SUB_88_U108 & new_P1_SUB_88_U110 & new_P1_SUB_88_U109;
  assign new_P1_SUB_88_U112 = ~P1_IR_REG_22_ & ~P1_IR_REG_23_ & ~P1_IR_REG_21_;
  assign new_P1_SUB_88_U113 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_24_;
  assign new_P1_SUB_88_U114 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U115 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U116 = new_P1_SUB_88_U112 & new_P1_SUB_88_U113 & new_P1_SUB_88_U115 & new_P1_SUB_88_U114;
  assign new_P1_SUB_88_U117 = ~P1_IR_REG_11_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_;
  assign new_P1_SUB_88_U118 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_ & ~P1_IR_REG_13_;
  assign new_P1_SUB_88_U119 = ~P1_IR_REG_17_ & ~P1_IR_REG_18_ & ~P1_IR_REG_16_;
  assign new_P1_SUB_88_U120 = ~P1_IR_REG_1_ & ~P1_IR_REG_0_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_88_U121 = new_P1_SUB_88_U117 & new_P1_SUB_88_U118 & new_P1_SUB_88_U120 & new_P1_SUB_88_U119;
  assign new_P1_SUB_88_U122 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_88_U123 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_23_;
  assign new_P1_SUB_88_U124 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U125 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U126 = new_P1_SUB_88_U122 & new_P1_SUB_88_U123 & new_P1_SUB_88_U125 & new_P1_SUB_88_U124;
  assign new_P1_SUB_88_U127 = ~P1_IR_REG_11_ & ~P1_IR_REG_10_ & ~P1_IR_REG_12_ & ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U128 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_15_ & ~P1_IR_REG_16_;
  assign new_P1_SUB_88_U129 = ~P1_IR_REG_5_ & ~P1_IR_REG_4_ & ~P1_IR_REG_2_ & ~P1_IR_REG_3_;
  assign new_P1_SUB_88_U130 = ~P1_IR_REG_9_ & ~P1_IR_REG_8_ & ~P1_IR_REG_6_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U131 = ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign new_P1_SUB_88_U132 = ~P1_IR_REG_19_ & ~P1_IR_REG_20_;
  assign new_P1_SUB_88_U133 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_;
  assign new_P1_SUB_88_U134 = new_P1_SUB_88_U133 & new_P1_SUB_88_U132 & new_P1_SUB_88_U131;
  assign new_P1_SUB_88_U135 = ~P1_IR_REG_11_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_;
  assign new_P1_SUB_88_U136 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_ & ~P1_IR_REG_13_;
  assign new_P1_SUB_88_U137 = new_P1_SUB_88_U136 & new_P1_SUB_88_U135;
  assign new_P1_SUB_88_U138 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_88_U139 = ~P1_IR_REG_20_ & ~P1_IR_REG_21_ & ~P1_IR_REG_0_;
  assign new_P1_SUB_88_U140 = ~P1_IR_REG_3_ & ~P1_IR_REG_4_ & ~P1_IR_REG_2_;
  assign new_P1_SUB_88_U141 = new_P1_SUB_88_U140 & new_P1_SUB_88_U139;
  assign new_P1_SUB_88_U142 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_7_ & ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_88_U143 = ~P1_IR_REG_11_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_;
  assign new_P1_SUB_88_U144 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_ & ~P1_IR_REG_13_;
  assign new_P1_SUB_88_U145 = ~P1_IR_REG_17_ & ~P1_IR_REG_16_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_88_U146 = ~P1_IR_REG_20_ & ~P1_IR_REG_0_ & ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U147 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_7_ & ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_88_U148 = ~P1_IR_REG_11_ & ~P1_IR_REG_10_ & ~P1_IR_REG_12_ & ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U149 = ~P1_IR_REG_16_ & ~P1_IR_REG_15_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign new_P1_SUB_88_U150 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_ & ~P1_IR_REG_2_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign new_P1_SUB_88_U151 = ~P1_IR_REG_6_ & ~P1_IR_REG_5_ & ~P1_IR_REG_7_ & ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_88_U152 = ~P1_IR_REG_11_ & ~P1_IR_REG_10_ & ~P1_IR_REG_12_ & ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U153 = ~P1_IR_REG_16_ & ~P1_IR_REG_15_ & ~P1_IR_REG_17_ & ~P1_IR_REG_18_ & ~P1_IR_REG_1_;
  assign new_P1_SUB_88_U154 = ~P1_IR_REG_2_ & ~P1_IR_REG_0_ & ~P1_IR_REG_3_ & ~P1_IR_REG_4_ & ~P1_IR_REG_5_;
  assign new_P1_SUB_88_U155 = ~P1_IR_REG_9_ & ~P1_IR_REG_8_ & ~P1_IR_REG_6_ & ~P1_IR_REG_7_;
  assign new_P1_SUB_88_U156 = ~P1_IR_REG_9_ & ~P1_IR_REG_12_ & ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign new_P1_SUB_88_U157 = ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign new_P1_SUB_88_U158 = ~P1_IR_REG_10_ & ~P1_IR_REG_9_;
  assign new_P1_SUB_88_U159 = ~P1_IR_REG_9_;
  assign new_P1_SUB_88_U160 = new_P1_SUB_88_U233 & new_P1_SUB_88_U232;
  assign new_P1_SUB_88_U161 = ~P1_IR_REG_5_;
  assign new_P1_SUB_88_U162 = new_P1_SUB_88_U235 & new_P1_SUB_88_U234;
  assign new_P1_SUB_88_U163 = ~P1_IR_REG_31_;
  assign new_P1_SUB_88_U164 = ~P1_IR_REG_30_;
  assign new_P1_SUB_88_U165 = new_P1_SUB_88_U239 & new_P1_SUB_88_U238;
  assign new_P1_SUB_88_U166 = ~P1_IR_REG_27_;
  assign new_P1_SUB_88_U167 = ~new_P1_SUB_88_U96 | ~new_P1_SUB_88_U91;
  assign new_P1_SUB_88_U168 = ~P1_IR_REG_25_;
  assign new_P1_SUB_88_U169 = ~new_P1_SUB_88_U116 | ~new_P1_SUB_88_U111;
  assign new_P1_SUB_88_U170 = new_P1_SUB_88_U243 & new_P1_SUB_88_U242;
  assign new_P1_SUB_88_U171 = ~P1_IR_REG_21_;
  assign new_P1_SUB_88_U172 = ~new_P1_SUB_88_U146 | ~new_P1_SUB_88_U147 | ~new_P1_SUB_88_U145 | ~new_P1_SUB_88_U144 | ~new_P1_SUB_88_U143;
  assign new_P1_SUB_88_U173 = new_P1_SUB_88_U245 & new_P1_SUB_88_U244;
  assign new_P1_SUB_88_U174 = ~P1_IR_REG_1_;
  assign new_P1_SUB_88_U175 = ~P1_IR_REG_0_;
  assign new_P1_SUB_88_U176 = ~P1_IR_REG_17_;
  assign new_P1_SUB_88_U177 = new_P1_SUB_88_U249 & new_P1_SUB_88_U248;
  assign new_P1_SUB_88_U178 = ~P1_IR_REG_13_;
  assign new_P1_SUB_88_U179 = new_P1_SUB_88_U251 & new_P1_SUB_88_U250;
  assign new_P1_SUB_88_U180 = ~new_P1_SUB_88_U230 | ~new_P1_SUB_88_U32;
  assign new_P1_SUB_88_U181 = ~new_P1_SUB_88_U29;
  assign new_P1_SUB_88_U182 = ~new_P1_SUB_88_U30;
  assign new_P1_SUB_88_U183 = ~new_P1_SUB_88_U182 | ~new_P1_SUB_88_U31;
  assign new_P1_SUB_88_U184 = ~new_P1_SUB_88_U28;
  assign new_P1_SUB_88_U185 = ~P1_IR_REG_8_ | ~new_P1_SUB_88_U183;
  assign new_P1_SUB_88_U186 = ~P1_IR_REG_7_ | ~new_P1_SUB_88_U30;
  assign new_P1_SUB_88_U187 = ~new_P1_SUB_88_U181 | ~new_P1_SUB_88_U161;
  assign new_P1_SUB_88_U188 = ~P1_IR_REG_6_ | ~new_P1_SUB_88_U187;
  assign new_P1_SUB_88_U189 = ~P1_IR_REG_4_ | ~new_P1_SUB_88_U180;
  assign new_P1_SUB_88_U190 = ~P1_IR_REG_3_ | ~new_P1_SUB_88_U27;
  assign new_P1_SUB_88_U191 = ~new_P1_SUB_88_U38;
  assign new_P1_SUB_88_U192 = ~new_P1_SUB_88_U191 | ~new_P1_SUB_88_U39;
  assign new_P1_SUB_88_U193 = ~new_P1_SUB_88_U35;
  assign new_P1_SUB_88_U194 = ~new_P1_SUB_88_U36;
  assign new_P1_SUB_88_U195 = ~new_P1_SUB_88_U194 | ~new_P1_SUB_88_U37;
  assign new_P1_SUB_88_U196 = ~new_P1_SUB_88_U34;
  assign new_P1_SUB_88_U197 = ~new_P1_SUB_88_U152 | ~new_P1_SUB_88_U153 | ~new_P1_SUB_88_U155 | ~new_P1_SUB_88_U154;
  assign new_P1_SUB_88_U198 = ~new_P1_SUB_88_U148 | ~new_P1_SUB_88_U149 | ~new_P1_SUB_88_U151 | ~new_P1_SUB_88_U150;
  assign new_P1_SUB_88_U199 = ~new_P1_SUB_88_U172;
  assign new_P1_SUB_88_U200 = ~new_P1_SUB_88_U134 | ~new_P1_SUB_88_U196;
  assign new_P1_SUB_88_U201 = ~new_P1_SUB_88_U126 | ~new_P1_SUB_88_U121;
  assign new_P1_SUB_88_U202 = ~new_P1_SUB_88_U169;
  assign new_P1_SUB_88_U203 = ~new_P1_SUB_88_U167;
  assign new_P1_SUB_88_U204 = ~new_P1_SUB_88_U66 | ~new_P1_SUB_88_U61;
  assign new_P1_SUB_88_U205 = ~new_P1_SUB_88_U33;
  assign new_P1_SUB_88_U206 = P1_IR_REG_1_ | P1_IR_REG_0_;
  assign new_P1_SUB_88_U207 = ~P1_IR_REG_2_ | ~new_P1_SUB_88_U206;
  assign new_P1_SUB_88_U208 = ~P1_IR_REG_29_ | ~new_P1_SUB_88_U204;
  assign new_P1_SUB_88_U209 = ~P1_IR_REG_28_ | ~new_P1_SUB_88_U229;
  assign new_P1_SUB_88_U210 = ~new_P1_SUB_88_U106 | ~new_P1_SUB_88_U101;
  assign new_P1_SUB_88_U211 = ~P1_IR_REG_26_ | ~new_P1_SUB_88_U210;
  assign new_P1_SUB_88_U212 = ~P1_IR_REG_24_ | ~new_P1_SUB_88_U201;
  assign new_P1_SUB_88_U213 = ~P1_IR_REG_23_ | ~new_P1_SUB_88_U200;
  assign new_P1_SUB_88_U214 = ~new_P1_SUB_88_U137 | ~new_P1_SUB_88_U138 | ~new_P1_SUB_88_U142 | ~new_P1_SUB_88_U141;
  assign new_P1_SUB_88_U215 = ~P1_IR_REG_22_ | ~new_P1_SUB_88_U214;
  assign new_P1_SUB_88_U216 = ~P1_IR_REG_20_ | ~new_P1_SUB_88_U198;
  assign new_P1_SUB_88_U217 = ~P1_IR_REG_19_ | ~new_P1_SUB_88_U197;
  assign new_P1_SUB_88_U218 = ~new_P1_SUB_88_U196 | ~new_P1_SUB_88_U176;
  assign new_P1_SUB_88_U219 = ~P1_IR_REG_18_ | ~new_P1_SUB_88_U218;
  assign new_P1_SUB_88_U220 = ~P1_IR_REG_16_ | ~new_P1_SUB_88_U195;
  assign new_P1_SUB_88_U221 = ~P1_IR_REG_15_ | ~new_P1_SUB_88_U36;
  assign new_P1_SUB_88_U222 = ~new_P1_SUB_88_U193 | ~new_P1_SUB_88_U178;
  assign new_P1_SUB_88_U223 = ~P1_IR_REG_14_ | ~new_P1_SUB_88_U222;
  assign new_P1_SUB_88_U224 = ~P1_IR_REG_12_ | ~new_P1_SUB_88_U192;
  assign new_P1_SUB_88_U225 = ~P1_IR_REG_11_ | ~new_P1_SUB_88_U38;
  assign new_P1_SUB_88_U226 = ~new_P1_SUB_88_U184 | ~new_P1_SUB_88_U159;
  assign new_P1_SUB_88_U227 = ~P1_IR_REG_10_ | ~new_P1_SUB_88_U226;
  assign new_P1_SUB_88_U228 = ~new_P1_SUB_88_U205 | ~new_P1_SUB_88_U164;
  assign new_P1_SUB_88_U229 = ~new_P1_SUB_88_U76 | ~new_P1_SUB_88_U71;
  assign new_P1_SUB_88_U230 = ~new_P1_SUB_88_U27;
  assign new_P1_SUB_88_U231 = ~new_P1_SUB_88_U86 | ~new_P1_SUB_88_U81;
  assign new_P1_SUB_88_U232 = ~P1_IR_REG_9_ | ~new_P1_SUB_88_U28;
  assign new_P1_SUB_88_U233 = ~new_P1_SUB_88_U184 | ~new_P1_SUB_88_U159;
  assign new_P1_SUB_88_U234 = ~P1_IR_REG_5_ | ~new_P1_SUB_88_U29;
  assign new_P1_SUB_88_U235 = ~new_P1_SUB_88_U181 | ~new_P1_SUB_88_U161;
  assign new_P1_SUB_88_U236 = ~new_P1_SUB_88_U228 | ~new_P1_SUB_88_U163;
  assign new_P1_SUB_88_U237 = ~P1_IR_REG_31_ | ~new_P1_SUB_88_U205 | ~new_P1_SUB_88_U164;
  assign new_P1_SUB_88_U238 = ~P1_IR_REG_30_ | ~new_P1_SUB_88_U33;
  assign new_P1_SUB_88_U239 = ~new_P1_SUB_88_U205 | ~new_P1_SUB_88_U164;
  assign new_P1_SUB_88_U240 = ~new_P1_SUB_88_U203 | ~P1_IR_REG_27_;
  assign new_P1_SUB_88_U241 = ~new_P1_SUB_88_U231 | ~new_P1_SUB_88_U166;
  assign new_P1_SUB_88_U242 = ~P1_IR_REG_25_ | ~new_P1_SUB_88_U169;
  assign new_P1_SUB_88_U243 = ~new_P1_SUB_88_U202 | ~new_P1_SUB_88_U168;
  assign new_P1_SUB_88_U244 = ~P1_IR_REG_21_ | ~new_P1_SUB_88_U172;
  assign new_P1_SUB_88_U245 = ~new_P1_SUB_88_U199 | ~new_P1_SUB_88_U171;
  assign new_P1_SUB_88_U246 = ~P1_IR_REG_1_ | ~new_P1_SUB_88_U175;
  assign new_P1_SUB_88_U247 = ~P1_IR_REG_0_ | ~new_P1_SUB_88_U174;
  assign new_P1_SUB_88_U248 = ~P1_IR_REG_17_ | ~new_P1_SUB_88_U34;
  assign new_P1_SUB_88_U249 = ~new_P1_SUB_88_U196 | ~new_P1_SUB_88_U176;
  assign new_P1_SUB_88_U250 = ~P1_IR_REG_13_ | ~new_P1_SUB_88_U35;
  assign new_P1_SUB_88_U251 = ~new_P1_SUB_88_U193 | ~new_P1_SUB_88_U178;
  assign new_P1_R1309_U6 = ~new_P1_U3059;
  assign new_P1_R1309_U7 = ~new_P1_U3056;
  assign new_P1_R1309_U8 = new_P1_R1309_U10 & new_P1_R1309_U9;
  assign new_P1_R1309_U9 = ~new_P1_U3056 | ~new_P1_R1309_U6;
  assign new_P1_R1309_U10 = ~new_P1_U3059 | ~new_P1_R1309_U7;
  assign new_P1_R1282_U6 = new_P1_R1282_U135 & new_P1_R1282_U35;
  assign new_P1_R1282_U7 = new_P1_R1282_U133 & new_P1_R1282_U36;
  assign new_P1_R1282_U8 = new_P1_R1282_U132 & new_P1_R1282_U37;
  assign new_P1_R1282_U9 = new_P1_R1282_U131 & new_P1_R1282_U38;
  assign new_P1_R1282_U10 = new_P1_R1282_U129 & new_P1_R1282_U39;
  assign new_P1_R1282_U11 = new_P1_R1282_U128 & new_P1_R1282_U40;
  assign new_P1_R1282_U12 = new_P1_R1282_U127 & new_P1_R1282_U41;
  assign new_P1_R1282_U13 = new_P1_R1282_U125 & new_P1_R1282_U42;
  assign new_P1_R1282_U14 = new_P1_R1282_U123 & new_P1_R1282_U43;
  assign new_P1_R1282_U15 = new_P1_R1282_U121 & new_P1_R1282_U44;
  assign new_P1_R1282_U16 = new_P1_R1282_U119 & new_P1_R1282_U45;
  assign new_P1_R1282_U17 = new_P1_R1282_U117 & new_P1_R1282_U46;
  assign new_P1_R1282_U18 = new_P1_R1282_U115 & new_P1_R1282_U25;
  assign new_P1_R1282_U19 = new_P1_R1282_U113 & new_P1_R1282_U67;
  assign new_P1_R1282_U20 = new_P1_R1282_U98 & new_P1_R1282_U26;
  assign new_P1_R1282_U21 = new_P1_R1282_U97 & new_P1_R1282_U27;
  assign new_P1_R1282_U22 = new_P1_R1282_U96 & new_P1_R1282_U28;
  assign new_P1_R1282_U23 = new_P1_R1282_U94 & new_P1_R1282_U29;
  assign new_P1_R1282_U24 = new_P1_R1282_U93 & new_P1_R1282_U30;
  assign new_P1_R1282_U25 = new_P1_U3464 | new_P1_U3461 | new_P1_U3456;
  assign new_P1_R1282_U26 = ~new_P1_R1282_U87 | ~new_P1_R1282_U34;
  assign new_P1_R1282_U27 = ~new_P1_R1282_U88 | ~new_P1_R1282_U33;
  assign new_P1_R1282_U28 = ~new_P1_R1282_U57 | ~new_P1_R1282_U89;
  assign new_P1_R1282_U29 = ~new_P1_R1282_U90 | ~new_P1_R1282_U32;
  assign new_P1_R1282_U30 = ~new_P1_R1282_U91 | ~new_P1_R1282_U31;
  assign new_P1_R1282_U31 = ~new_P1_U3482;
  assign new_P1_R1282_U32 = ~new_P1_U3479;
  assign new_P1_R1282_U33 = ~new_P1_U3470;
  assign new_P1_R1282_U34 = ~new_P1_U3467;
  assign new_P1_R1282_U35 = ~new_P1_R1282_U58 | ~new_P1_R1282_U92;
  assign new_P1_R1282_U36 = ~new_P1_R1282_U99 | ~new_P1_R1282_U55;
  assign new_P1_R1282_U37 = ~new_P1_R1282_U100 | ~new_P1_R1282_U54;
  assign new_P1_R1282_U38 = ~new_P1_R1282_U59 | ~new_P1_R1282_U101;
  assign new_P1_R1282_U39 = ~new_P1_R1282_U102 | ~new_P1_R1282_U53;
  assign new_P1_R1282_U40 = ~new_P1_R1282_U103 | ~new_P1_R1282_U52;
  assign new_P1_R1282_U41 = ~new_P1_R1282_U60 | ~new_P1_R1282_U104;
  assign new_P1_R1282_U42 = ~new_P1_R1282_U61 | ~new_P1_R1282_U105;
  assign new_P1_R1282_U43 = ~new_P1_R1282_U51 | ~new_P1_R1282_U106 | ~new_P1_R1282_U77;
  assign new_P1_R1282_U44 = ~new_P1_R1282_U50 | ~new_P1_R1282_U107 | ~new_P1_R1282_U75;
  assign new_P1_R1282_U45 = ~new_P1_R1282_U49 | ~new_P1_R1282_U108 | ~new_P1_R1282_U73;
  assign new_P1_R1282_U46 = ~new_P1_R1282_U48 | ~new_P1_R1282_U109 | ~new_P1_R1282_U71;
  assign new_P1_R1282_U47 = ~new_P1_U4027;
  assign new_P1_R1282_U48 = ~new_P1_U4017;
  assign new_P1_R1282_U49 = ~new_P1_U4019;
  assign new_P1_R1282_U50 = ~new_P1_U4021;
  assign new_P1_R1282_U51 = ~new_P1_U4023;
  assign new_P1_R1282_U52 = ~new_P1_U3506;
  assign new_P1_R1282_U53 = ~new_P1_U3503;
  assign new_P1_R1282_U54 = ~new_P1_U3494;
  assign new_P1_R1282_U55 = ~new_P1_U3491;
  assign new_P1_R1282_U56 = ~new_P1_R1282_U153 | ~new_P1_R1282_U152;
  assign new_P1_R1282_U57 = ~new_P1_U3473 & ~new_P1_U3476;
  assign new_P1_R1282_U58 = ~new_P1_U3488 & ~new_P1_U3485;
  assign new_P1_R1282_U59 = ~new_P1_U3497 & ~new_P1_U3500;
  assign new_P1_R1282_U60 = ~new_P1_U3509 & ~new_P1_U3512;
  assign new_P1_R1282_U61 = ~new_P1_U3514 & ~new_P1_U4025;
  assign new_P1_R1282_U62 = ~new_P1_U3485;
  assign new_P1_R1282_U63 = new_P1_R1282_U137 & new_P1_R1282_U136;
  assign new_P1_R1282_U64 = ~new_P1_U3473;
  assign new_P1_R1282_U65 = new_P1_R1282_U139 & new_P1_R1282_U138;
  assign new_P1_R1282_U66 = ~new_P1_U4026;
  assign new_P1_R1282_U67 = ~new_P1_R1282_U47 | ~new_P1_R1282_U110 | ~new_P1_R1282_U69;
  assign new_P1_R1282_U68 = new_P1_R1282_U141 & new_P1_R1282_U140;
  assign new_P1_R1282_U69 = ~new_P1_U4028;
  assign new_P1_R1282_U70 = new_P1_R1282_U143 & new_P1_R1282_U142;
  assign new_P1_R1282_U71 = ~new_P1_U4018;
  assign new_P1_R1282_U72 = new_P1_R1282_U145 & new_P1_R1282_U144;
  assign new_P1_R1282_U73 = ~new_P1_U4020;
  assign new_P1_R1282_U74 = new_P1_R1282_U147 & new_P1_R1282_U146;
  assign new_P1_R1282_U75 = ~new_P1_U4022;
  assign new_P1_R1282_U76 = new_P1_R1282_U149 & new_P1_R1282_U148;
  assign new_P1_R1282_U77 = ~new_P1_U4024;
  assign new_P1_R1282_U78 = new_P1_R1282_U151 & new_P1_R1282_U150;
  assign new_P1_R1282_U79 = ~new_P1_U3461;
  assign new_P1_R1282_U80 = ~new_P1_U3456;
  assign new_P1_R1282_U81 = ~new_P1_U3514;
  assign new_P1_R1282_U82 = new_P1_R1282_U155 & new_P1_R1282_U154;
  assign new_P1_R1282_U83 = ~new_P1_U3509;
  assign new_P1_R1282_U84 = new_P1_R1282_U157 & new_P1_R1282_U156;
  assign new_P1_R1282_U85 = ~new_P1_U3497;
  assign new_P1_R1282_U86 = new_P1_R1282_U159 & new_P1_R1282_U158;
  assign new_P1_R1282_U87 = ~new_P1_R1282_U25;
  assign new_P1_R1282_U88 = ~new_P1_R1282_U26;
  assign new_P1_R1282_U89 = ~new_P1_R1282_U27;
  assign new_P1_R1282_U90 = ~new_P1_R1282_U28;
  assign new_P1_R1282_U91 = ~new_P1_R1282_U29;
  assign new_P1_R1282_U92 = ~new_P1_R1282_U30;
  assign new_P1_R1282_U93 = ~new_P1_U3482 | ~new_P1_R1282_U29;
  assign new_P1_R1282_U94 = ~new_P1_U3479 | ~new_P1_R1282_U28;
  assign new_P1_R1282_U95 = ~new_P1_R1282_U89 | ~new_P1_R1282_U64;
  assign new_P1_R1282_U96 = ~new_P1_U3476 | ~new_P1_R1282_U95;
  assign new_P1_R1282_U97 = ~new_P1_U3470 | ~new_P1_R1282_U26;
  assign new_P1_R1282_U98 = ~new_P1_U3467 | ~new_P1_R1282_U25;
  assign new_P1_R1282_U99 = ~new_P1_R1282_U35;
  assign new_P1_R1282_U100 = ~new_P1_R1282_U36;
  assign new_P1_R1282_U101 = ~new_P1_R1282_U37;
  assign new_P1_R1282_U102 = ~new_P1_R1282_U38;
  assign new_P1_R1282_U103 = ~new_P1_R1282_U39;
  assign new_P1_R1282_U104 = ~new_P1_R1282_U40;
  assign new_P1_R1282_U105 = ~new_P1_R1282_U41;
  assign new_P1_R1282_U106 = ~new_P1_R1282_U42;
  assign new_P1_R1282_U107 = ~new_P1_R1282_U43;
  assign new_P1_R1282_U108 = ~new_P1_R1282_U44;
  assign new_P1_R1282_U109 = ~new_P1_R1282_U45;
  assign new_P1_R1282_U110 = ~new_P1_R1282_U46;
  assign new_P1_R1282_U111 = ~new_P1_R1282_U67;
  assign new_P1_R1282_U112 = ~new_P1_R1282_U110 | ~new_P1_R1282_U69;
  assign new_P1_R1282_U113 = ~new_P1_U4027 | ~new_P1_R1282_U112;
  assign new_P1_R1282_U114 = new_P1_U3461 | new_P1_U3456;
  assign new_P1_R1282_U115 = ~new_P1_U3464 | ~new_P1_R1282_U114;
  assign new_P1_R1282_U116 = ~new_P1_R1282_U109 | ~new_P1_R1282_U71;
  assign new_P1_R1282_U117 = ~new_P1_U4017 | ~new_P1_R1282_U116;
  assign new_P1_R1282_U118 = ~new_P1_R1282_U108 | ~new_P1_R1282_U73;
  assign new_P1_R1282_U119 = ~new_P1_U4019 | ~new_P1_R1282_U118;
  assign new_P1_R1282_U120 = ~new_P1_R1282_U107 | ~new_P1_R1282_U75;
  assign new_P1_R1282_U121 = ~new_P1_U4021 | ~new_P1_R1282_U120;
  assign new_P1_R1282_U122 = ~new_P1_R1282_U106 | ~new_P1_R1282_U77;
  assign new_P1_R1282_U123 = ~new_P1_U4023 | ~new_P1_R1282_U122;
  assign new_P1_R1282_U124 = ~new_P1_R1282_U105 | ~new_P1_R1282_U81;
  assign new_P1_R1282_U125 = ~new_P1_U4025 | ~new_P1_R1282_U124;
  assign new_P1_R1282_U126 = ~new_P1_R1282_U104 | ~new_P1_R1282_U83;
  assign new_P1_R1282_U127 = ~new_P1_U3512 | ~new_P1_R1282_U126;
  assign new_P1_R1282_U128 = ~new_P1_U3506 | ~new_P1_R1282_U39;
  assign new_P1_R1282_U129 = ~new_P1_U3503 | ~new_P1_R1282_U38;
  assign new_P1_R1282_U130 = ~new_P1_R1282_U101 | ~new_P1_R1282_U85;
  assign new_P1_R1282_U131 = ~new_P1_U3500 | ~new_P1_R1282_U130;
  assign new_P1_R1282_U132 = ~new_P1_U3494 | ~new_P1_R1282_U36;
  assign new_P1_R1282_U133 = ~new_P1_U3491 | ~new_P1_R1282_U35;
  assign new_P1_R1282_U134 = ~new_P1_R1282_U92 | ~new_P1_R1282_U62;
  assign new_P1_R1282_U135 = ~new_P1_U3488 | ~new_P1_R1282_U134;
  assign new_P1_R1282_U136 = ~new_P1_U3485 | ~new_P1_R1282_U30;
  assign new_P1_R1282_U137 = ~new_P1_R1282_U92 | ~new_P1_R1282_U62;
  assign new_P1_R1282_U138 = ~new_P1_U3473 | ~new_P1_R1282_U27;
  assign new_P1_R1282_U139 = ~new_P1_R1282_U89 | ~new_P1_R1282_U64;
  assign new_P1_R1282_U140 = ~new_P1_U4026 | ~new_P1_R1282_U67;
  assign new_P1_R1282_U141 = ~new_P1_R1282_U111 | ~new_P1_R1282_U66;
  assign new_P1_R1282_U142 = ~new_P1_U4028 | ~new_P1_R1282_U46;
  assign new_P1_R1282_U143 = ~new_P1_R1282_U110 | ~new_P1_R1282_U69;
  assign new_P1_R1282_U144 = ~new_P1_U4018 | ~new_P1_R1282_U45;
  assign new_P1_R1282_U145 = ~new_P1_R1282_U109 | ~new_P1_R1282_U71;
  assign new_P1_R1282_U146 = ~new_P1_U4020 | ~new_P1_R1282_U44;
  assign new_P1_R1282_U147 = ~new_P1_R1282_U108 | ~new_P1_R1282_U73;
  assign new_P1_R1282_U148 = ~new_P1_U4022 | ~new_P1_R1282_U43;
  assign new_P1_R1282_U149 = ~new_P1_R1282_U107 | ~new_P1_R1282_U75;
  assign new_P1_R1282_U150 = ~new_P1_U4024 | ~new_P1_R1282_U42;
  assign new_P1_R1282_U151 = ~new_P1_R1282_U106 | ~new_P1_R1282_U77;
  assign new_P1_R1282_U152 = ~new_P1_U3461 | ~new_P1_R1282_U80;
  assign new_P1_R1282_U153 = ~new_P1_U3456 | ~new_P1_R1282_U79;
  assign new_P1_R1282_U154 = ~new_P1_U3514 | ~new_P1_R1282_U41;
  assign new_P1_R1282_U155 = ~new_P1_R1282_U105 | ~new_P1_R1282_U81;
  assign new_P1_R1282_U156 = ~new_P1_U3509 | ~new_P1_R1282_U40;
  assign new_P1_R1282_U157 = ~new_P1_R1282_U104 | ~new_P1_R1282_U83;
  assign new_P1_R1282_U158 = ~new_P1_U3497 | ~new_P1_R1282_U37;
  assign new_P1_R1282_U159 = ~new_P1_R1282_U101 | ~new_P1_R1282_U85;
  assign new_P1_R1240_U4 = new_P1_R1240_U176 & new_P1_R1240_U175;
  assign new_P1_R1240_U5 = new_P1_R1240_U177 & new_P1_R1240_U178;
  assign new_P1_R1240_U6 = new_P1_R1240_U194 & new_P1_R1240_U193;
  assign new_P1_R1240_U7 = new_P1_R1240_U234 & new_P1_R1240_U233;
  assign new_P1_R1240_U8 = new_P1_R1240_U243 & new_P1_R1240_U242;
  assign new_P1_R1240_U9 = new_P1_R1240_U261 & new_P1_R1240_U260;
  assign new_P1_R1240_U10 = new_P1_R1240_U269 & new_P1_R1240_U268;
  assign new_P1_R1240_U11 = new_P1_R1240_U348 & new_P1_R1240_U345;
  assign new_P1_R1240_U12 = new_P1_R1240_U341 & new_P1_R1240_U338;
  assign new_P1_R1240_U13 = new_P1_R1240_U332 & new_P1_R1240_U329;
  assign new_P1_R1240_U14 = new_P1_R1240_U323 & new_P1_R1240_U320;
  assign new_P1_R1240_U15 = new_P1_R1240_U317 & new_P1_R1240_U315;
  assign new_P1_R1240_U16 = new_P1_R1240_U310 & new_P1_R1240_U307;
  assign new_P1_R1240_U17 = new_P1_R1240_U232 & new_P1_R1240_U229;
  assign new_P1_R1240_U18 = new_P1_R1240_U224 & new_P1_R1240_U221;
  assign new_P1_R1240_U19 = new_P1_R1240_U210 & new_P1_R1240_U207;
  assign new_P1_R1240_U20 = ~new_P1_U3476;
  assign new_P1_R1240_U21 = ~new_P1_U3071;
  assign new_P1_R1240_U22 = ~new_P1_U3070;
  assign new_P1_R1240_U23 = ~new_P1_U3071 | ~new_P1_U3476;
  assign new_P1_R1240_U24 = ~new_P1_U3479;
  assign new_P1_R1240_U25 = ~new_P1_U3470;
  assign new_P1_R1240_U26 = ~new_P1_U3060;
  assign new_P1_R1240_U27 = ~new_P1_U3067;
  assign new_P1_R1240_U28 = ~new_P1_U3464;
  assign new_P1_R1240_U29 = ~new_P1_U3068;
  assign new_P1_R1240_U30 = ~new_P1_U3456;
  assign new_P1_R1240_U31 = ~new_P1_U3077;
  assign new_P1_R1240_U32 = ~new_P1_U3077 | ~new_P1_U3456;
  assign new_P1_R1240_U33 = ~new_P1_U3467;
  assign new_P1_R1240_U34 = ~new_P1_U3064;
  assign new_P1_R1240_U35 = ~new_P1_U3060 | ~new_P1_U3470;
  assign new_P1_R1240_U36 = ~new_P1_U3473;
  assign new_P1_R1240_U37 = ~new_P1_U3482;
  assign new_P1_R1240_U38 = ~new_P1_U3084;
  assign new_P1_R1240_U39 = ~new_P1_U3083;
  assign new_P1_R1240_U40 = ~new_P1_U3485;
  assign new_P1_R1240_U41 = ~new_P1_R1240_U62 | ~new_P1_R1240_U202;
  assign new_P1_R1240_U42 = ~new_P1_R1240_U118 | ~new_P1_R1240_U190;
  assign new_P1_R1240_U43 = ~new_P1_R1240_U179 | ~new_P1_R1240_U180;
  assign new_P1_R1240_U44 = ~new_P1_U3461 | ~new_P1_U3078;
  assign new_P1_R1240_U45 = ~new_P1_R1240_U122 | ~new_P1_R1240_U216;
  assign new_P1_R1240_U46 = ~new_P1_R1240_U213 | ~new_P1_R1240_U212;
  assign new_P1_R1240_U47 = ~new_P1_U4018;
  assign new_P1_R1240_U48 = ~new_P1_U3053;
  assign new_P1_R1240_U49 = ~new_P1_U3057;
  assign new_P1_R1240_U50 = ~new_P1_U4019;
  assign new_P1_R1240_U51 = ~new_P1_U4020;
  assign new_P1_R1240_U52 = ~new_P1_U3058;
  assign new_P1_R1240_U53 = ~new_P1_U4021;
  assign new_P1_R1240_U54 = ~new_P1_U3065;
  assign new_P1_R1240_U55 = ~new_P1_U4024;
  assign new_P1_R1240_U56 = ~new_P1_U3075;
  assign new_P1_R1240_U57 = ~new_P1_U3506;
  assign new_P1_R1240_U58 = ~new_P1_U3073;
  assign new_P1_R1240_U59 = ~new_P1_U3069;
  assign new_P1_R1240_U60 = ~new_P1_U3073 | ~new_P1_U3506;
  assign new_P1_R1240_U61 = ~new_P1_U3509;
  assign new_P1_R1240_U62 = ~new_P1_U3084 | ~new_P1_U3482;
  assign new_P1_R1240_U63 = ~new_P1_U3488;
  assign new_P1_R1240_U64 = ~new_P1_U3062;
  assign new_P1_R1240_U65 = ~new_P1_U3494;
  assign new_P1_R1240_U66 = ~new_P1_U3072;
  assign new_P1_R1240_U67 = ~new_P1_U3491;
  assign new_P1_R1240_U68 = ~new_P1_U3063;
  assign new_P1_R1240_U69 = ~new_P1_U3063 | ~new_P1_U3491;
  assign new_P1_R1240_U70 = ~new_P1_U3497;
  assign new_P1_R1240_U71 = ~new_P1_U3080;
  assign new_P1_R1240_U72 = ~new_P1_U3500;
  assign new_P1_R1240_U73 = ~new_P1_U3079;
  assign new_P1_R1240_U74 = ~new_P1_U3503;
  assign new_P1_R1240_U75 = ~new_P1_U3074;
  assign new_P1_R1240_U76 = ~new_P1_U3512;
  assign new_P1_R1240_U77 = ~new_P1_U3082;
  assign new_P1_R1240_U78 = ~new_P1_U3082 | ~new_P1_U3512;
  assign new_P1_R1240_U79 = ~new_P1_U3514;
  assign new_P1_R1240_U80 = ~new_P1_U3081;
  assign new_P1_R1240_U81 = ~new_P1_U3081 | ~new_P1_U3514;
  assign new_P1_R1240_U82 = ~new_P1_U4025;
  assign new_P1_R1240_U83 = ~new_P1_U4023;
  assign new_P1_R1240_U84 = ~new_P1_U3061;
  assign new_P1_R1240_U85 = ~new_P1_U4022;
  assign new_P1_R1240_U86 = ~new_P1_U3066;
  assign new_P1_R1240_U87 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1240_U88 = ~new_P1_U3054;
  assign new_P1_R1240_U89 = ~new_P1_U4017;
  assign new_P1_R1240_U90 = ~new_P1_R1240_U303 | ~new_P1_R1240_U173;
  assign new_P1_R1240_U91 = ~new_P1_U3076;
  assign new_P1_R1240_U92 = ~new_P1_R1240_U78 | ~new_P1_R1240_U312;
  assign new_P1_R1240_U93 = ~new_P1_R1240_U258 | ~new_P1_R1240_U257;
  assign new_P1_R1240_U94 = ~new_P1_R1240_U69 | ~new_P1_R1240_U334;
  assign new_P1_R1240_U95 = ~new_P1_R1240_U454 | ~new_P1_R1240_U453;
  assign new_P1_R1240_U96 = ~new_P1_R1240_U501 | ~new_P1_R1240_U500;
  assign new_P1_R1240_U97 = ~new_P1_R1240_U372 | ~new_P1_R1240_U371;
  assign new_P1_R1240_U98 = ~new_P1_R1240_U377 | ~new_P1_R1240_U376;
  assign new_P1_R1240_U99 = ~new_P1_R1240_U384 | ~new_P1_R1240_U383;
  assign new_P1_R1240_U100 = ~new_P1_R1240_U391 | ~new_P1_R1240_U390;
  assign new_P1_R1240_U101 = ~new_P1_R1240_U396 | ~new_P1_R1240_U395;
  assign new_P1_R1240_U102 = ~new_P1_R1240_U405 | ~new_P1_R1240_U404;
  assign new_P1_R1240_U103 = ~new_P1_R1240_U412 | ~new_P1_R1240_U411;
  assign new_P1_R1240_U104 = ~new_P1_R1240_U419 | ~new_P1_R1240_U418;
  assign new_P1_R1240_U105 = ~new_P1_R1240_U426 | ~new_P1_R1240_U425;
  assign new_P1_R1240_U106 = ~new_P1_R1240_U431 | ~new_P1_R1240_U430;
  assign new_P1_R1240_U107 = ~new_P1_R1240_U438 | ~new_P1_R1240_U437;
  assign new_P1_R1240_U108 = ~new_P1_R1240_U445 | ~new_P1_R1240_U444;
  assign new_P1_R1240_U109 = ~new_P1_R1240_U459 | ~new_P1_R1240_U458;
  assign new_P1_R1240_U110 = ~new_P1_R1240_U464 | ~new_P1_R1240_U463;
  assign new_P1_R1240_U111 = ~new_P1_R1240_U471 | ~new_P1_R1240_U470;
  assign new_P1_R1240_U112 = ~new_P1_R1240_U478 | ~new_P1_R1240_U477;
  assign new_P1_R1240_U113 = ~new_P1_R1240_U485 | ~new_P1_R1240_U484;
  assign new_P1_R1240_U114 = ~new_P1_R1240_U492 | ~new_P1_R1240_U491;
  assign new_P1_R1240_U115 = ~new_P1_R1240_U497 | ~new_P1_R1240_U496;
  assign new_P1_R1240_U116 = new_P1_U3464 & new_P1_U3068;
  assign new_P1_R1240_U117 = new_P1_R1240_U186 & new_P1_R1240_U184;
  assign new_P1_R1240_U118 = new_P1_R1240_U191 & new_P1_R1240_U189;
  assign new_P1_R1240_U119 = new_P1_R1240_U198 & new_P1_R1240_U197;
  assign new_P1_R1240_U120 = new_P1_R1240_U23 & new_P1_R1240_U379 & new_P1_R1240_U378;
  assign new_P1_R1240_U121 = new_P1_R1240_U209 & new_P1_R1240_U6;
  assign new_P1_R1240_U122 = new_P1_R1240_U217 & new_P1_R1240_U215;
  assign new_P1_R1240_U123 = new_P1_R1240_U35 & new_P1_R1240_U386 & new_P1_R1240_U385;
  assign new_P1_R1240_U124 = new_P1_R1240_U223 & new_P1_R1240_U4;
  assign new_P1_R1240_U125 = new_P1_R1240_U231 & new_P1_R1240_U178;
  assign new_P1_R1240_U126 = new_P1_R1240_U201 & new_P1_R1240_U7;
  assign new_P1_R1240_U127 = new_P1_R1240_U236 & new_P1_R1240_U168;
  assign new_P1_R1240_U128 = new_P1_R1240_U245 & new_P1_R1240_U169;
  assign new_P1_R1240_U129 = new_P1_R1240_U265 & new_P1_R1240_U264;
  assign new_P1_R1240_U130 = new_P1_R1240_U10 & new_P1_R1240_U279;
  assign new_P1_R1240_U131 = new_P1_R1240_U282 & new_P1_R1240_U277;
  assign new_P1_R1240_U132 = new_P1_R1240_U298 & new_P1_R1240_U295;
  assign new_P1_R1240_U133 = new_P1_R1240_U365 & new_P1_R1240_U299;
  assign new_P1_R1240_U134 = new_P1_R1240_U156 & new_P1_R1240_U275;
  assign new_P1_R1240_U135 = new_P1_R1240_U60 & new_P1_R1240_U466 & new_P1_R1240_U465;
  assign new_P1_R1240_U136 = new_P1_R1240_U169 & new_P1_R1240_U487 & new_P1_R1240_U486;
  assign new_P1_R1240_U137 = new_P1_R1240_U340 & new_P1_R1240_U8;
  assign new_P1_R1240_U138 = new_P1_R1240_U168 & new_P1_R1240_U499 & new_P1_R1240_U498;
  assign new_P1_R1240_U139 = new_P1_R1240_U347 & new_P1_R1240_U7;
  assign new_P1_R1240_U140 = ~new_P1_R1240_U119 | ~new_P1_R1240_U199;
  assign new_P1_R1240_U141 = ~new_P1_R1240_U214 | ~new_P1_R1240_U226;
  assign new_P1_R1240_U142 = ~new_P1_U3055;
  assign new_P1_R1240_U143 = ~new_P1_U4028;
  assign new_P1_R1240_U144 = new_P1_R1240_U400 & new_P1_R1240_U399;
  assign new_P1_R1240_U145 = ~new_P1_R1240_U361 | ~new_P1_R1240_U301 | ~new_P1_R1240_U166;
  assign new_P1_R1240_U146 = new_P1_R1240_U407 & new_P1_R1240_U406;
  assign new_P1_R1240_U147 = ~new_P1_R1240_U133 | ~new_P1_R1240_U367 | ~new_P1_R1240_U366;
  assign new_P1_R1240_U148 = new_P1_R1240_U414 & new_P1_R1240_U413;
  assign new_P1_R1240_U149 = ~new_P1_R1240_U87 | ~new_P1_R1240_U362 | ~new_P1_R1240_U296;
  assign new_P1_R1240_U150 = new_P1_R1240_U421 & new_P1_R1240_U420;
  assign new_P1_R1240_U151 = ~new_P1_R1240_U290 | ~new_P1_R1240_U289;
  assign new_P1_R1240_U152 = new_P1_R1240_U433 & new_P1_R1240_U432;
  assign new_P1_R1240_U153 = ~new_P1_R1240_U286 | ~new_P1_R1240_U285;
  assign new_P1_R1240_U154 = new_P1_R1240_U440 & new_P1_R1240_U439;
  assign new_P1_R1240_U155 = ~new_P1_R1240_U131 | ~new_P1_R1240_U281;
  assign new_P1_R1240_U156 = new_P1_R1240_U447 & new_P1_R1240_U446;
  assign new_P1_R1240_U157 = new_P1_R1240_U452 & new_P1_R1240_U451;
  assign new_P1_R1240_U158 = ~new_P1_R1240_U44 | ~new_P1_R1240_U324;
  assign new_P1_R1240_U159 = ~new_P1_R1240_U129 | ~new_P1_R1240_U266;
  assign new_P1_R1240_U160 = new_P1_R1240_U473 & new_P1_R1240_U472;
  assign new_P1_R1240_U161 = ~new_P1_R1240_U254 | ~new_P1_R1240_U253;
  assign new_P1_R1240_U162 = new_P1_R1240_U480 & new_P1_R1240_U479;
  assign new_P1_R1240_U163 = ~new_P1_R1240_U250 | ~new_P1_R1240_U249;
  assign new_P1_R1240_U164 = ~new_P1_R1240_U240 | ~new_P1_R1240_U239;
  assign new_P1_R1240_U165 = ~new_P1_R1240_U364 | ~new_P1_R1240_U363;
  assign new_P1_R1240_U166 = ~new_P1_U3054 | ~new_P1_R1240_U147;
  assign new_P1_R1240_U167 = ~new_P1_R1240_U35;
  assign new_P1_R1240_U168 = ~new_P1_U3485 | ~new_P1_U3083;
  assign new_P1_R1240_U169 = ~new_P1_U3072 | ~new_P1_U3494;
  assign new_P1_R1240_U170 = ~new_P1_U3058 | ~new_P1_U4020;
  assign new_P1_R1240_U171 = ~new_P1_R1240_U69;
  assign new_P1_R1240_U172 = ~new_P1_R1240_U78;
  assign new_P1_R1240_U173 = ~new_P1_U3065 | ~new_P1_U4021;
  assign new_P1_R1240_U174 = ~new_P1_R1240_U62;
  assign new_P1_R1240_U175 = new_P1_U3067 | new_P1_U3473;
  assign new_P1_R1240_U176 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1240_U177 = new_P1_U3467 | new_P1_U3064;
  assign new_P1_R1240_U178 = new_P1_U3464 | new_P1_U3068;
  assign new_P1_R1240_U179 = ~new_P1_R1240_U32;
  assign new_P1_R1240_U180 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1240_U181 = ~new_P1_R1240_U43;
  assign new_P1_R1240_U182 = ~new_P1_R1240_U44;
  assign new_P1_R1240_U183 = ~new_P1_R1240_U43 | ~new_P1_R1240_U44;
  assign new_P1_R1240_U184 = ~new_P1_R1240_U116 | ~new_P1_R1240_U177;
  assign new_P1_R1240_U185 = ~new_P1_R1240_U5 | ~new_P1_R1240_U183;
  assign new_P1_R1240_U186 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1240_U187 = ~new_P1_R1240_U117 | ~new_P1_R1240_U185;
  assign new_P1_R1240_U188 = ~new_P1_R1240_U36 | ~new_P1_R1240_U35;
  assign new_P1_R1240_U189 = ~new_P1_U3067 | ~new_P1_R1240_U188;
  assign new_P1_R1240_U190 = ~new_P1_R1240_U4 | ~new_P1_R1240_U187;
  assign new_P1_R1240_U191 = ~new_P1_U3473 | ~new_P1_R1240_U167;
  assign new_P1_R1240_U192 = ~new_P1_R1240_U42;
  assign new_P1_R1240_U193 = new_P1_U3070 | new_P1_U3479;
  assign new_P1_R1240_U194 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1240_U195 = ~new_P1_R1240_U23;
  assign new_P1_R1240_U196 = ~new_P1_R1240_U24 | ~new_P1_R1240_U23;
  assign new_P1_R1240_U197 = ~new_P1_U3070 | ~new_P1_R1240_U196;
  assign new_P1_R1240_U198 = ~new_P1_U3479 | ~new_P1_R1240_U195;
  assign new_P1_R1240_U199 = ~new_P1_R1240_U6 | ~new_P1_R1240_U42;
  assign new_P1_R1240_U200 = ~new_P1_R1240_U140;
  assign new_P1_R1240_U201 = new_P1_U3482 | new_P1_U3084;
  assign new_P1_R1240_U202 = ~new_P1_R1240_U201 | ~new_P1_R1240_U140;
  assign new_P1_R1240_U203 = ~new_P1_R1240_U41;
  assign new_P1_R1240_U204 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1240_U205 = new_P1_U3476 | new_P1_U3071;
  assign new_P1_R1240_U206 = ~new_P1_R1240_U205 | ~new_P1_R1240_U42;
  assign new_P1_R1240_U207 = ~new_P1_R1240_U120 | ~new_P1_R1240_U206;
  assign new_P1_R1240_U208 = ~new_P1_R1240_U192 | ~new_P1_R1240_U23;
  assign new_P1_R1240_U209 = ~new_P1_U3479 | ~new_P1_U3070;
  assign new_P1_R1240_U210 = ~new_P1_R1240_U121 | ~new_P1_R1240_U208;
  assign new_P1_R1240_U211 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1240_U212 = ~new_P1_R1240_U182 | ~new_P1_R1240_U178;
  assign new_P1_R1240_U213 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1240_U214 = ~new_P1_R1240_U46;
  assign new_P1_R1240_U215 = ~new_P1_R1240_U181 | ~new_P1_R1240_U5;
  assign new_P1_R1240_U216 = ~new_P1_R1240_U46 | ~new_P1_R1240_U177;
  assign new_P1_R1240_U217 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1240_U218 = ~new_P1_R1240_U45;
  assign new_P1_R1240_U219 = new_P1_U3470 | new_P1_U3060;
  assign new_P1_R1240_U220 = ~new_P1_R1240_U219 | ~new_P1_R1240_U45;
  assign new_P1_R1240_U221 = ~new_P1_R1240_U123 | ~new_P1_R1240_U220;
  assign new_P1_R1240_U222 = ~new_P1_R1240_U218 | ~new_P1_R1240_U35;
  assign new_P1_R1240_U223 = ~new_P1_U3473 | ~new_P1_U3067;
  assign new_P1_R1240_U224 = ~new_P1_R1240_U124 | ~new_P1_R1240_U222;
  assign new_P1_R1240_U225 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1240_U226 = ~new_P1_R1240_U181 | ~new_P1_R1240_U178;
  assign new_P1_R1240_U227 = ~new_P1_R1240_U141;
  assign new_P1_R1240_U228 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1240_U229 = ~new_P1_R1240_U43 | ~new_P1_R1240_U44 | ~new_P1_R1240_U398 | ~new_P1_R1240_U397;
  assign new_P1_R1240_U230 = ~new_P1_R1240_U44 | ~new_P1_R1240_U43;
  assign new_P1_R1240_U231 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1240_U232 = ~new_P1_R1240_U125 | ~new_P1_R1240_U230;
  assign new_P1_R1240_U233 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1240_U234 = new_P1_U3062 | new_P1_U3488;
  assign new_P1_R1240_U235 = ~new_P1_R1240_U174 | ~new_P1_R1240_U7;
  assign new_P1_R1240_U236 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1240_U237 = ~new_P1_R1240_U127 | ~new_P1_R1240_U235;
  assign new_P1_R1240_U238 = new_P1_U3488 | new_P1_U3062;
  assign new_P1_R1240_U239 = ~new_P1_R1240_U126 | ~new_P1_R1240_U140;
  assign new_P1_R1240_U240 = ~new_P1_R1240_U238 | ~new_P1_R1240_U237;
  assign new_P1_R1240_U241 = ~new_P1_R1240_U164;
  assign new_P1_R1240_U242 = new_P1_U3080 | new_P1_U3497;
  assign new_P1_R1240_U243 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1240_U244 = ~new_P1_R1240_U171 | ~new_P1_R1240_U8;
  assign new_P1_R1240_U245 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1240_U246 = ~new_P1_R1240_U128 | ~new_P1_R1240_U244;
  assign new_P1_R1240_U247 = new_P1_U3491 | new_P1_U3063;
  assign new_P1_R1240_U248 = new_P1_U3497 | new_P1_U3080;
  assign new_P1_R1240_U249 = ~new_P1_R1240_U8 | ~new_P1_R1240_U247 | ~new_P1_R1240_U164;
  assign new_P1_R1240_U250 = ~new_P1_R1240_U248 | ~new_P1_R1240_U246;
  assign new_P1_R1240_U251 = ~new_P1_R1240_U163;
  assign new_P1_R1240_U252 = new_P1_U3500 | new_P1_U3079;
  assign new_P1_R1240_U253 = ~new_P1_R1240_U252 | ~new_P1_R1240_U163;
  assign new_P1_R1240_U254 = ~new_P1_U3079 | ~new_P1_U3500;
  assign new_P1_R1240_U255 = ~new_P1_R1240_U161;
  assign new_P1_R1240_U256 = new_P1_U3503 | new_P1_U3074;
  assign new_P1_R1240_U257 = ~new_P1_R1240_U256 | ~new_P1_R1240_U161;
  assign new_P1_R1240_U258 = ~new_P1_U3074 | ~new_P1_U3503;
  assign new_P1_R1240_U259 = ~new_P1_R1240_U93;
  assign new_P1_R1240_U260 = new_P1_U3069 | new_P1_U3509;
  assign new_P1_R1240_U261 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1240_U262 = ~new_P1_R1240_U60;
  assign new_P1_R1240_U263 = ~new_P1_R1240_U61 | ~new_P1_R1240_U60;
  assign new_P1_R1240_U264 = ~new_P1_U3069 | ~new_P1_R1240_U263;
  assign new_P1_R1240_U265 = ~new_P1_U3509 | ~new_P1_R1240_U262;
  assign new_P1_R1240_U266 = ~new_P1_R1240_U9 | ~new_P1_R1240_U93;
  assign new_P1_R1240_U267 = ~new_P1_R1240_U159;
  assign new_P1_R1240_U268 = new_P1_U3076 | new_P1_U4025;
  assign new_P1_R1240_U269 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1240_U270 = new_P1_U3075 | new_P1_U4024;
  assign new_P1_R1240_U271 = ~new_P1_R1240_U81;
  assign new_P1_R1240_U272 = ~new_P1_U4025 | ~new_P1_R1240_U271;
  assign new_P1_R1240_U273 = ~new_P1_R1240_U272 | ~new_P1_R1240_U91;
  assign new_P1_R1240_U274 = ~new_P1_R1240_U81 | ~new_P1_R1240_U82;
  assign new_P1_R1240_U275 = ~new_P1_R1240_U274 | ~new_P1_R1240_U273;
  assign new_P1_R1240_U276 = ~new_P1_R1240_U172 | ~new_P1_R1240_U10;
  assign new_P1_R1240_U277 = ~new_P1_U3075 | ~new_P1_U4024;
  assign new_P1_R1240_U278 = ~new_P1_R1240_U275 | ~new_P1_R1240_U276;
  assign new_P1_R1240_U279 = new_P1_U3512 | new_P1_U3082;
  assign new_P1_R1240_U280 = new_P1_U4024 | new_P1_U3075;
  assign new_P1_R1240_U281 = ~new_P1_R1240_U130 | ~new_P1_R1240_U270 | ~new_P1_R1240_U159;
  assign new_P1_R1240_U282 = ~new_P1_R1240_U280 | ~new_P1_R1240_U278;
  assign new_P1_R1240_U283 = ~new_P1_R1240_U155;
  assign new_P1_R1240_U284 = new_P1_U4023 | new_P1_U3061;
  assign new_P1_R1240_U285 = ~new_P1_R1240_U284 | ~new_P1_R1240_U155;
  assign new_P1_R1240_U286 = ~new_P1_U3061 | ~new_P1_U4023;
  assign new_P1_R1240_U287 = ~new_P1_R1240_U153;
  assign new_P1_R1240_U288 = new_P1_U4022 | new_P1_U3066;
  assign new_P1_R1240_U289 = ~new_P1_R1240_U288 | ~new_P1_R1240_U153;
  assign new_P1_R1240_U290 = ~new_P1_U3066 | ~new_P1_U4022;
  assign new_P1_R1240_U291 = ~new_P1_R1240_U151;
  assign new_P1_R1240_U292 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1240_U293 = ~new_P1_R1240_U173 | ~new_P1_R1240_U170;
  assign new_P1_R1240_U294 = ~new_P1_R1240_U87;
  assign new_P1_R1240_U295 = new_P1_U4021 | new_P1_U3065;
  assign new_P1_R1240_U296 = ~new_P1_R1240_U165 | ~new_P1_R1240_U151 | ~new_P1_R1240_U295;
  assign new_P1_R1240_U297 = ~new_P1_R1240_U149;
  assign new_P1_R1240_U298 = new_P1_U4018 | new_P1_U3053;
  assign new_P1_R1240_U299 = ~new_P1_U3053 | ~new_P1_U4018;
  assign new_P1_R1240_U300 = ~new_P1_R1240_U147;
  assign new_P1_R1240_U301 = ~new_P1_U4017 | ~new_P1_R1240_U147;
  assign new_P1_R1240_U302 = ~new_P1_R1240_U145;
  assign new_P1_R1240_U303 = ~new_P1_R1240_U295 | ~new_P1_R1240_U151;
  assign new_P1_R1240_U304 = ~new_P1_R1240_U90;
  assign new_P1_R1240_U305 = new_P1_U4020 | new_P1_U3058;
  assign new_P1_R1240_U306 = ~new_P1_R1240_U305 | ~new_P1_R1240_U90;
  assign new_P1_R1240_U307 = ~new_P1_R1240_U150 | ~new_P1_R1240_U306 | ~new_P1_R1240_U170;
  assign new_P1_R1240_U308 = ~new_P1_R1240_U304 | ~new_P1_R1240_U170;
  assign new_P1_R1240_U309 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1240_U310 = ~new_P1_R1240_U165 | ~new_P1_R1240_U308 | ~new_P1_R1240_U309;
  assign new_P1_R1240_U311 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1240_U312 = ~new_P1_R1240_U279 | ~new_P1_R1240_U159;
  assign new_P1_R1240_U313 = ~new_P1_R1240_U92;
  assign new_P1_R1240_U314 = ~new_P1_R1240_U10 | ~new_P1_R1240_U92;
  assign new_P1_R1240_U315 = ~new_P1_R1240_U134 | ~new_P1_R1240_U314;
  assign new_P1_R1240_U316 = ~new_P1_R1240_U314 | ~new_P1_R1240_U275;
  assign new_P1_R1240_U317 = ~new_P1_R1240_U450 | ~new_P1_R1240_U316;
  assign new_P1_R1240_U318 = new_P1_U3514 | new_P1_U3081;
  assign new_P1_R1240_U319 = ~new_P1_R1240_U318 | ~new_P1_R1240_U92;
  assign new_P1_R1240_U320 = ~new_P1_R1240_U157 | ~new_P1_R1240_U319 | ~new_P1_R1240_U81;
  assign new_P1_R1240_U321 = ~new_P1_R1240_U313 | ~new_P1_R1240_U81;
  assign new_P1_R1240_U322 = ~new_P1_U3076 | ~new_P1_U4025;
  assign new_P1_R1240_U323 = ~new_P1_R1240_U10 | ~new_P1_R1240_U322 | ~new_P1_R1240_U321;
  assign new_P1_R1240_U324 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1240_U325 = ~new_P1_R1240_U158;
  assign new_P1_R1240_U326 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1240_U327 = new_P1_U3506 | new_P1_U3073;
  assign new_P1_R1240_U328 = ~new_P1_R1240_U327 | ~new_P1_R1240_U93;
  assign new_P1_R1240_U329 = ~new_P1_R1240_U135 | ~new_P1_R1240_U328;
  assign new_P1_R1240_U330 = ~new_P1_R1240_U259 | ~new_P1_R1240_U60;
  assign new_P1_R1240_U331 = ~new_P1_U3509 | ~new_P1_U3069;
  assign new_P1_R1240_U332 = ~new_P1_R1240_U9 | ~new_P1_R1240_U331 | ~new_P1_R1240_U330;
  assign new_P1_R1240_U333 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1240_U334 = ~new_P1_R1240_U247 | ~new_P1_R1240_U164;
  assign new_P1_R1240_U335 = ~new_P1_R1240_U94;
  assign new_P1_R1240_U336 = new_P1_U3494 | new_P1_U3072;
  assign new_P1_R1240_U337 = ~new_P1_R1240_U336 | ~new_P1_R1240_U94;
  assign new_P1_R1240_U338 = ~new_P1_R1240_U136 | ~new_P1_R1240_U337;
  assign new_P1_R1240_U339 = ~new_P1_R1240_U335 | ~new_P1_R1240_U169;
  assign new_P1_R1240_U340 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1240_U341 = ~new_P1_R1240_U137 | ~new_P1_R1240_U339;
  assign new_P1_R1240_U342 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1240_U343 = new_P1_U3485 | new_P1_U3083;
  assign new_P1_R1240_U344 = ~new_P1_R1240_U343 | ~new_P1_R1240_U41;
  assign new_P1_R1240_U345 = ~new_P1_R1240_U138 | ~new_P1_R1240_U344;
  assign new_P1_R1240_U346 = ~new_P1_R1240_U203 | ~new_P1_R1240_U168;
  assign new_P1_R1240_U347 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1240_U348 = ~new_P1_R1240_U139 | ~new_P1_R1240_U346;
  assign new_P1_R1240_U349 = ~new_P1_R1240_U204 | ~new_P1_R1240_U168;
  assign new_P1_R1240_U350 = ~new_P1_R1240_U201 | ~new_P1_R1240_U62;
  assign new_P1_R1240_U351 = ~new_P1_R1240_U211 | ~new_P1_R1240_U23;
  assign new_P1_R1240_U352 = ~new_P1_R1240_U225 | ~new_P1_R1240_U35;
  assign new_P1_R1240_U353 = ~new_P1_R1240_U228 | ~new_P1_R1240_U177;
  assign new_P1_R1240_U354 = ~new_P1_R1240_U311 | ~new_P1_R1240_U170;
  assign new_P1_R1240_U355 = ~new_P1_R1240_U295 | ~new_P1_R1240_U173;
  assign new_P1_R1240_U356 = ~new_P1_R1240_U326 | ~new_P1_R1240_U81;
  assign new_P1_R1240_U357 = ~new_P1_R1240_U279 | ~new_P1_R1240_U78;
  assign new_P1_R1240_U358 = ~new_P1_R1240_U333 | ~new_P1_R1240_U60;
  assign new_P1_R1240_U359 = ~new_P1_R1240_U342 | ~new_P1_R1240_U169;
  assign new_P1_R1240_U360 = ~new_P1_R1240_U247 | ~new_P1_R1240_U69;
  assign new_P1_R1240_U361 = ~new_P1_U4017 | ~new_P1_U3054;
  assign new_P1_R1240_U362 = ~new_P1_R1240_U293 | ~new_P1_R1240_U165;
  assign new_P1_R1240_U363 = ~new_P1_U3057 | ~new_P1_R1240_U292;
  assign new_P1_R1240_U364 = ~new_P1_U4019 | ~new_P1_R1240_U292;
  assign new_P1_R1240_U365 = ~new_P1_R1240_U298 | ~new_P1_R1240_U293 | ~new_P1_R1240_U165;
  assign new_P1_R1240_U366 = ~new_P1_R1240_U132 | ~new_P1_R1240_U151 | ~new_P1_R1240_U165;
  assign new_P1_R1240_U367 = ~new_P1_R1240_U294 | ~new_P1_R1240_U298;
  assign new_P1_R1240_U368 = ~new_P1_U3083 | ~new_P1_R1240_U40;
  assign new_P1_R1240_U369 = ~new_P1_U3485 | ~new_P1_R1240_U39;
  assign new_P1_R1240_U370 = ~new_P1_R1240_U369 | ~new_P1_R1240_U368;
  assign new_P1_R1240_U371 = ~new_P1_R1240_U349 | ~new_P1_R1240_U41;
  assign new_P1_R1240_U372 = ~new_P1_R1240_U370 | ~new_P1_R1240_U203;
  assign new_P1_R1240_U373 = ~new_P1_U3084 | ~new_P1_R1240_U37;
  assign new_P1_R1240_U374 = ~new_P1_U3482 | ~new_P1_R1240_U38;
  assign new_P1_R1240_U375 = ~new_P1_R1240_U374 | ~new_P1_R1240_U373;
  assign new_P1_R1240_U376 = ~new_P1_R1240_U350 | ~new_P1_R1240_U140;
  assign new_P1_R1240_U377 = ~new_P1_R1240_U200 | ~new_P1_R1240_U375;
  assign new_P1_R1240_U378 = ~new_P1_U3070 | ~new_P1_R1240_U24;
  assign new_P1_R1240_U379 = ~new_P1_U3479 | ~new_P1_R1240_U22;
  assign new_P1_R1240_U380 = ~new_P1_U3071 | ~new_P1_R1240_U20;
  assign new_P1_R1240_U381 = ~new_P1_U3476 | ~new_P1_R1240_U21;
  assign new_P1_R1240_U382 = ~new_P1_R1240_U381 | ~new_P1_R1240_U380;
  assign new_P1_R1240_U383 = ~new_P1_R1240_U351 | ~new_P1_R1240_U42;
  assign new_P1_R1240_U384 = ~new_P1_R1240_U382 | ~new_P1_R1240_U192;
  assign new_P1_R1240_U385 = ~new_P1_U3067 | ~new_P1_R1240_U36;
  assign new_P1_R1240_U386 = ~new_P1_U3473 | ~new_P1_R1240_U27;
  assign new_P1_R1240_U387 = ~new_P1_U3060 | ~new_P1_R1240_U25;
  assign new_P1_R1240_U388 = ~new_P1_U3470 | ~new_P1_R1240_U26;
  assign new_P1_R1240_U389 = ~new_P1_R1240_U388 | ~new_P1_R1240_U387;
  assign new_P1_R1240_U390 = ~new_P1_R1240_U352 | ~new_P1_R1240_U45;
  assign new_P1_R1240_U391 = ~new_P1_R1240_U389 | ~new_P1_R1240_U218;
  assign new_P1_R1240_U392 = ~new_P1_U3064 | ~new_P1_R1240_U33;
  assign new_P1_R1240_U393 = ~new_P1_U3467 | ~new_P1_R1240_U34;
  assign new_P1_R1240_U394 = ~new_P1_R1240_U393 | ~new_P1_R1240_U392;
  assign new_P1_R1240_U395 = ~new_P1_R1240_U353 | ~new_P1_R1240_U141;
  assign new_P1_R1240_U396 = ~new_P1_R1240_U227 | ~new_P1_R1240_U394;
  assign new_P1_R1240_U397 = ~new_P1_U3068 | ~new_P1_R1240_U28;
  assign new_P1_R1240_U398 = ~new_P1_U3464 | ~new_P1_R1240_U29;
  assign new_P1_R1240_U399 = ~new_P1_U3055 | ~new_P1_R1240_U143;
  assign new_P1_R1240_U400 = ~new_P1_U4028 | ~new_P1_R1240_U142;
  assign new_P1_R1240_U401 = ~new_P1_U3055 | ~new_P1_R1240_U143;
  assign new_P1_R1240_U402 = ~new_P1_U4028 | ~new_P1_R1240_U142;
  assign new_P1_R1240_U403 = ~new_P1_R1240_U402 | ~new_P1_R1240_U401;
  assign new_P1_R1240_U404 = ~new_P1_R1240_U144 | ~new_P1_R1240_U145;
  assign new_P1_R1240_U405 = ~new_P1_R1240_U302 | ~new_P1_R1240_U403;
  assign new_P1_R1240_U406 = ~new_P1_U3054 | ~new_P1_R1240_U89;
  assign new_P1_R1240_U407 = ~new_P1_U4017 | ~new_P1_R1240_U88;
  assign new_P1_R1240_U408 = ~new_P1_U3054 | ~new_P1_R1240_U89;
  assign new_P1_R1240_U409 = ~new_P1_U4017 | ~new_P1_R1240_U88;
  assign new_P1_R1240_U410 = ~new_P1_R1240_U409 | ~new_P1_R1240_U408;
  assign new_P1_R1240_U411 = ~new_P1_R1240_U146 | ~new_P1_R1240_U147;
  assign new_P1_R1240_U412 = ~new_P1_R1240_U300 | ~new_P1_R1240_U410;
  assign new_P1_R1240_U413 = ~new_P1_U3053 | ~new_P1_R1240_U47;
  assign new_P1_R1240_U414 = ~new_P1_U4018 | ~new_P1_R1240_U48;
  assign new_P1_R1240_U415 = ~new_P1_U3053 | ~new_P1_R1240_U47;
  assign new_P1_R1240_U416 = ~new_P1_U4018 | ~new_P1_R1240_U48;
  assign new_P1_R1240_U417 = ~new_P1_R1240_U416 | ~new_P1_R1240_U415;
  assign new_P1_R1240_U418 = ~new_P1_R1240_U148 | ~new_P1_R1240_U149;
  assign new_P1_R1240_U419 = ~new_P1_R1240_U297 | ~new_P1_R1240_U417;
  assign new_P1_R1240_U420 = ~new_P1_U3057 | ~new_P1_R1240_U50;
  assign new_P1_R1240_U421 = ~new_P1_U4019 | ~new_P1_R1240_U49;
  assign new_P1_R1240_U422 = ~new_P1_U3058 | ~new_P1_R1240_U51;
  assign new_P1_R1240_U423 = ~new_P1_U4020 | ~new_P1_R1240_U52;
  assign new_P1_R1240_U424 = ~new_P1_R1240_U423 | ~new_P1_R1240_U422;
  assign new_P1_R1240_U425 = ~new_P1_R1240_U354 | ~new_P1_R1240_U90;
  assign new_P1_R1240_U426 = ~new_P1_R1240_U424 | ~new_P1_R1240_U304;
  assign new_P1_R1240_U427 = ~new_P1_U3065 | ~new_P1_R1240_U53;
  assign new_P1_R1240_U428 = ~new_P1_U4021 | ~new_P1_R1240_U54;
  assign new_P1_R1240_U429 = ~new_P1_R1240_U428 | ~new_P1_R1240_U427;
  assign new_P1_R1240_U430 = ~new_P1_R1240_U355 | ~new_P1_R1240_U151;
  assign new_P1_R1240_U431 = ~new_P1_R1240_U291 | ~new_P1_R1240_U429;
  assign new_P1_R1240_U432 = ~new_P1_U3066 | ~new_P1_R1240_U85;
  assign new_P1_R1240_U433 = ~new_P1_U4022 | ~new_P1_R1240_U86;
  assign new_P1_R1240_U434 = ~new_P1_U3066 | ~new_P1_R1240_U85;
  assign new_P1_R1240_U435 = ~new_P1_U4022 | ~new_P1_R1240_U86;
  assign new_P1_R1240_U436 = ~new_P1_R1240_U435 | ~new_P1_R1240_U434;
  assign new_P1_R1240_U437 = ~new_P1_R1240_U152 | ~new_P1_R1240_U153;
  assign new_P1_R1240_U438 = ~new_P1_R1240_U287 | ~new_P1_R1240_U436;
  assign new_P1_R1240_U439 = ~new_P1_U3061 | ~new_P1_R1240_U83;
  assign new_P1_R1240_U440 = ~new_P1_U4023 | ~new_P1_R1240_U84;
  assign new_P1_R1240_U441 = ~new_P1_U3061 | ~new_P1_R1240_U83;
  assign new_P1_R1240_U442 = ~new_P1_U4023 | ~new_P1_R1240_U84;
  assign new_P1_R1240_U443 = ~new_P1_R1240_U442 | ~new_P1_R1240_U441;
  assign new_P1_R1240_U444 = ~new_P1_R1240_U154 | ~new_P1_R1240_U155;
  assign new_P1_R1240_U445 = ~new_P1_R1240_U283 | ~new_P1_R1240_U443;
  assign new_P1_R1240_U446 = ~new_P1_U3075 | ~new_P1_R1240_U55;
  assign new_P1_R1240_U447 = ~new_P1_U4024 | ~new_P1_R1240_U56;
  assign new_P1_R1240_U448 = ~new_P1_U3075 | ~new_P1_R1240_U55;
  assign new_P1_R1240_U449 = ~new_P1_U4024 | ~new_P1_R1240_U56;
  assign new_P1_R1240_U450 = ~new_P1_R1240_U449 | ~new_P1_R1240_U448;
  assign new_P1_R1240_U451 = ~new_P1_U3076 | ~new_P1_R1240_U82;
  assign new_P1_R1240_U452 = ~new_P1_U4025 | ~new_P1_R1240_U91;
  assign new_P1_R1240_U453 = ~new_P1_R1240_U179 | ~new_P1_R1240_U158;
  assign new_P1_R1240_U454 = ~new_P1_R1240_U325 | ~new_P1_R1240_U32;
  assign new_P1_R1240_U455 = ~new_P1_U3081 | ~new_P1_R1240_U79;
  assign new_P1_R1240_U456 = ~new_P1_U3514 | ~new_P1_R1240_U80;
  assign new_P1_R1240_U457 = ~new_P1_R1240_U456 | ~new_P1_R1240_U455;
  assign new_P1_R1240_U458 = ~new_P1_R1240_U356 | ~new_P1_R1240_U92;
  assign new_P1_R1240_U459 = ~new_P1_R1240_U457 | ~new_P1_R1240_U313;
  assign new_P1_R1240_U460 = ~new_P1_U3082 | ~new_P1_R1240_U76;
  assign new_P1_R1240_U461 = ~new_P1_U3512 | ~new_P1_R1240_U77;
  assign new_P1_R1240_U462 = ~new_P1_R1240_U461 | ~new_P1_R1240_U460;
  assign new_P1_R1240_U463 = ~new_P1_R1240_U357 | ~new_P1_R1240_U159;
  assign new_P1_R1240_U464 = ~new_P1_R1240_U267 | ~new_P1_R1240_U462;
  assign new_P1_R1240_U465 = ~new_P1_U3069 | ~new_P1_R1240_U61;
  assign new_P1_R1240_U466 = ~new_P1_U3509 | ~new_P1_R1240_U59;
  assign new_P1_R1240_U467 = ~new_P1_U3073 | ~new_P1_R1240_U57;
  assign new_P1_R1240_U468 = ~new_P1_U3506 | ~new_P1_R1240_U58;
  assign new_P1_R1240_U469 = ~new_P1_R1240_U468 | ~new_P1_R1240_U467;
  assign new_P1_R1240_U470 = ~new_P1_R1240_U358 | ~new_P1_R1240_U93;
  assign new_P1_R1240_U471 = ~new_P1_R1240_U469 | ~new_P1_R1240_U259;
  assign new_P1_R1240_U472 = ~new_P1_U3074 | ~new_P1_R1240_U74;
  assign new_P1_R1240_U473 = ~new_P1_U3503 | ~new_P1_R1240_U75;
  assign new_P1_R1240_U474 = ~new_P1_U3074 | ~new_P1_R1240_U74;
  assign new_P1_R1240_U475 = ~new_P1_U3503 | ~new_P1_R1240_U75;
  assign new_P1_R1240_U476 = ~new_P1_R1240_U475 | ~new_P1_R1240_U474;
  assign new_P1_R1240_U477 = ~new_P1_R1240_U160 | ~new_P1_R1240_U161;
  assign new_P1_R1240_U478 = ~new_P1_R1240_U255 | ~new_P1_R1240_U476;
  assign new_P1_R1240_U479 = ~new_P1_U3079 | ~new_P1_R1240_U72;
  assign new_P1_R1240_U480 = ~new_P1_U3500 | ~new_P1_R1240_U73;
  assign new_P1_R1240_U481 = ~new_P1_U3079 | ~new_P1_R1240_U72;
  assign new_P1_R1240_U482 = ~new_P1_U3500 | ~new_P1_R1240_U73;
  assign new_P1_R1240_U483 = ~new_P1_R1240_U482 | ~new_P1_R1240_U481;
  assign new_P1_R1240_U484 = ~new_P1_R1240_U162 | ~new_P1_R1240_U163;
  assign new_P1_R1240_U485 = ~new_P1_R1240_U251 | ~new_P1_R1240_U483;
  assign new_P1_R1240_U486 = ~new_P1_U3080 | ~new_P1_R1240_U70;
  assign new_P1_R1240_U487 = ~new_P1_U3497 | ~new_P1_R1240_U71;
  assign new_P1_R1240_U488 = ~new_P1_U3072 | ~new_P1_R1240_U65;
  assign new_P1_R1240_U489 = ~new_P1_U3494 | ~new_P1_R1240_U66;
  assign new_P1_R1240_U490 = ~new_P1_R1240_U489 | ~new_P1_R1240_U488;
  assign new_P1_R1240_U491 = ~new_P1_R1240_U359 | ~new_P1_R1240_U94;
  assign new_P1_R1240_U492 = ~new_P1_R1240_U490 | ~new_P1_R1240_U335;
  assign new_P1_R1240_U493 = ~new_P1_U3063 | ~new_P1_R1240_U67;
  assign new_P1_R1240_U494 = ~new_P1_U3491 | ~new_P1_R1240_U68;
  assign new_P1_R1240_U495 = ~new_P1_R1240_U494 | ~new_P1_R1240_U493;
  assign new_P1_R1240_U496 = ~new_P1_R1240_U360 | ~new_P1_R1240_U164;
  assign new_P1_R1240_U497 = ~new_P1_R1240_U241 | ~new_P1_R1240_U495;
  assign new_P1_R1240_U498 = ~new_P1_U3062 | ~new_P1_R1240_U63;
  assign new_P1_R1240_U499 = ~new_P1_U3488 | ~new_P1_R1240_U64;
  assign new_P1_R1240_U500 = ~new_P1_U3077 | ~new_P1_R1240_U30;
  assign new_P1_R1240_U501 = ~new_P1_U3456 | ~new_P1_R1240_U31;
  assign new_P1_R1162_U4 = new_P1_R1162_U95 & new_P1_R1162_U94;
  assign new_P1_R1162_U5 = new_P1_R1162_U96 & new_P1_R1162_U97;
  assign new_P1_R1162_U6 = new_P1_R1162_U113 & new_P1_R1162_U112;
  assign new_P1_R1162_U7 = new_P1_R1162_U155 & new_P1_R1162_U154;
  assign new_P1_R1162_U8 = new_P1_R1162_U164 & new_P1_R1162_U163;
  assign new_P1_R1162_U9 = new_P1_R1162_U182 & new_P1_R1162_U181;
  assign new_P1_R1162_U10 = new_P1_R1162_U218 & new_P1_R1162_U215;
  assign new_P1_R1162_U11 = new_P1_R1162_U211 & new_P1_R1162_U208;
  assign new_P1_R1162_U12 = new_P1_R1162_U202 & new_P1_R1162_U199;
  assign new_P1_R1162_U13 = new_P1_R1162_U196 & new_P1_R1162_U192;
  assign new_P1_R1162_U14 = new_P1_R1162_U151 & new_P1_R1162_U148;
  assign new_P1_R1162_U15 = new_P1_R1162_U143 & new_P1_R1162_U140;
  assign new_P1_R1162_U16 = new_P1_R1162_U129 & new_P1_R1162_U126;
  assign new_P1_R1162_U17 = ~P1_REG1_REG_6_;
  assign new_P1_R1162_U18 = ~new_P1_U3475;
  assign new_P1_R1162_U19 = ~new_P1_U3478;
  assign new_P1_R1162_U20 = ~new_P1_U3475 | ~P1_REG1_REG_6_;
  assign new_P1_R1162_U21 = ~P1_REG1_REG_7_;
  assign new_P1_R1162_U22 = ~P1_REG1_REG_4_;
  assign new_P1_R1162_U23 = ~new_P1_U3469;
  assign new_P1_R1162_U24 = ~new_P1_U3472;
  assign new_P1_R1162_U25 = ~P1_REG1_REG_2_;
  assign new_P1_R1162_U26 = ~new_P1_U3463;
  assign new_P1_R1162_U27 = ~P1_REG1_REG_0_;
  assign new_P1_R1162_U28 = ~new_P1_U3454;
  assign new_P1_R1162_U29 = ~new_P1_U3454 | ~P1_REG1_REG_0_;
  assign new_P1_R1162_U30 = ~P1_REG1_REG_3_;
  assign new_P1_R1162_U31 = ~new_P1_U3466;
  assign new_P1_R1162_U32 = ~new_P1_U3469 | ~P1_REG1_REG_4_;
  assign new_P1_R1162_U33 = ~P1_REG1_REG_5_;
  assign new_P1_R1162_U34 = ~P1_REG1_REG_8_;
  assign new_P1_R1162_U35 = ~new_P1_U3481;
  assign new_P1_R1162_U36 = ~new_P1_U3484;
  assign new_P1_R1162_U37 = ~P1_REG1_REG_9_;
  assign new_P1_R1162_U38 = ~new_P1_R1162_U49 | ~new_P1_R1162_U121;
  assign new_P1_R1162_U39 = ~new_P1_R1162_U109 | ~new_P1_R1162_U110 | ~new_P1_R1162_U108;
  assign new_P1_R1162_U40 = ~new_P1_R1162_U98 | ~new_P1_R1162_U99;
  assign new_P1_R1162_U41 = ~P1_REG1_REG_1_ | ~new_P1_U3460;
  assign new_P1_R1162_U42 = ~new_P1_R1162_U135 | ~new_P1_R1162_U136 | ~new_P1_R1162_U134;
  assign new_P1_R1162_U43 = ~new_P1_R1162_U132 | ~new_P1_R1162_U131;
  assign new_P1_R1162_U44 = ~P1_REG1_REG_16_;
  assign new_P1_R1162_U45 = ~new_P1_U3505;
  assign new_P1_R1162_U46 = ~new_P1_U3508;
  assign new_P1_R1162_U47 = ~new_P1_U3505 | ~P1_REG1_REG_16_;
  assign new_P1_R1162_U48 = ~P1_REG1_REG_17_;
  assign new_P1_R1162_U49 = ~new_P1_U3481 | ~P1_REG1_REG_8_;
  assign new_P1_R1162_U50 = ~P1_REG1_REG_10_;
  assign new_P1_R1162_U51 = ~new_P1_U3487;
  assign new_P1_R1162_U52 = ~P1_REG1_REG_12_;
  assign new_P1_R1162_U53 = ~new_P1_U3493;
  assign new_P1_R1162_U54 = ~P1_REG1_REG_11_;
  assign new_P1_R1162_U55 = ~new_P1_U3490;
  assign new_P1_R1162_U56 = ~new_P1_U3490 | ~P1_REG1_REG_11_;
  assign new_P1_R1162_U57 = ~P1_REG1_REG_13_;
  assign new_P1_R1162_U58 = ~new_P1_U3496;
  assign new_P1_R1162_U59 = ~P1_REG1_REG_14_;
  assign new_P1_R1162_U60 = ~new_P1_U3499;
  assign new_P1_R1162_U61 = ~P1_REG1_REG_15_;
  assign new_P1_R1162_U62 = ~new_P1_U3502;
  assign new_P1_R1162_U63 = ~P1_REG1_REG_18_;
  assign new_P1_R1162_U64 = ~new_P1_U3511;
  assign new_P1_R1162_U65 = ~new_P1_R1162_U187 | ~new_P1_R1162_U186 | ~new_P1_R1162_U185;
  assign new_P1_R1162_U66 = ~new_P1_R1162_U179 | ~new_P1_R1162_U178;
  assign new_P1_R1162_U67 = ~new_P1_R1162_U56 | ~new_P1_R1162_U204;
  assign new_P1_R1162_U68 = ~new_P1_R1162_U259 | ~new_P1_R1162_U258;
  assign new_P1_R1162_U69 = ~new_P1_R1162_U308 | ~new_P1_R1162_U307;
  assign new_P1_R1162_U70 = ~new_P1_R1162_U231 | ~new_P1_R1162_U230;
  assign new_P1_R1162_U71 = ~new_P1_R1162_U236 | ~new_P1_R1162_U235;
  assign new_P1_R1162_U72 = ~new_P1_R1162_U243 | ~new_P1_R1162_U242;
  assign new_P1_R1162_U73 = ~new_P1_R1162_U250 | ~new_P1_R1162_U249;
  assign new_P1_R1162_U74 = ~new_P1_R1162_U255 | ~new_P1_R1162_U254;
  assign new_P1_R1162_U75 = ~new_P1_R1162_U271 | ~new_P1_R1162_U270;
  assign new_P1_R1162_U76 = ~new_P1_R1162_U278 | ~new_P1_R1162_U277;
  assign new_P1_R1162_U77 = ~new_P1_R1162_U285 | ~new_P1_R1162_U284;
  assign new_P1_R1162_U78 = ~new_P1_R1162_U292 | ~new_P1_R1162_U291;
  assign new_P1_R1162_U79 = ~new_P1_R1162_U299 | ~new_P1_R1162_U298;
  assign new_P1_R1162_U80 = ~new_P1_R1162_U304 | ~new_P1_R1162_U303;
  assign new_P1_R1162_U81 = ~new_P1_R1162_U118 | ~new_P1_R1162_U117 | ~new_P1_R1162_U116;
  assign new_P1_R1162_U82 = ~new_P1_R1162_U133 | ~new_P1_R1162_U145;
  assign new_P1_R1162_U83 = ~new_P1_R1162_U41 | ~new_P1_R1162_U152;
  assign new_P1_R1162_U84 = ~new_P1_U3452;
  assign new_P1_R1162_U85 = ~P1_REG1_REG_19_;
  assign new_P1_R1162_U86 = ~new_P1_R1162_U175 | ~new_P1_R1162_U174;
  assign new_P1_R1162_U87 = ~new_P1_R1162_U171 | ~new_P1_R1162_U170;
  assign new_P1_R1162_U88 = ~new_P1_R1162_U161 | ~new_P1_R1162_U160;
  assign new_P1_R1162_U89 = ~new_P1_R1162_U32;
  assign new_P1_R1162_U90 = ~P1_REG1_REG_9_ | ~new_P1_U3484;
  assign new_P1_R1162_U91 = ~new_P1_U3493 | ~P1_REG1_REG_12_;
  assign new_P1_R1162_U92 = ~new_P1_R1162_U56;
  assign new_P1_R1162_U93 = ~new_P1_R1162_U49;
  assign new_P1_R1162_U94 = new_P1_U3472 | P1_REG1_REG_5_;
  assign new_P1_R1162_U95 = new_P1_U3469 | P1_REG1_REG_4_;
  assign new_P1_R1162_U96 = P1_REG1_REG_3_ | new_P1_U3466;
  assign new_P1_R1162_U97 = P1_REG1_REG_2_ | new_P1_U3463;
  assign new_P1_R1162_U98 = ~new_P1_R1162_U29;
  assign new_P1_R1162_U99 = P1_REG1_REG_1_ | new_P1_U3460;
  assign new_P1_R1162_U100 = ~new_P1_R1162_U40;
  assign new_P1_R1162_U101 = ~new_P1_R1162_U41;
  assign new_P1_R1162_U102 = ~new_P1_R1162_U40 | ~new_P1_R1162_U41;
  assign new_P1_R1162_U103 = ~new_P1_R1162_U96 | ~P1_REG1_REG_2_ | ~new_P1_U3463;
  assign new_P1_R1162_U104 = ~new_P1_R1162_U5 | ~new_P1_R1162_U102;
  assign new_P1_R1162_U105 = ~new_P1_U3466 | ~P1_REG1_REG_3_;
  assign new_P1_R1162_U106 = ~new_P1_R1162_U104 | ~new_P1_R1162_U105 | ~new_P1_R1162_U103;
  assign new_P1_R1162_U107 = ~new_P1_R1162_U33 | ~new_P1_R1162_U32;
  assign new_P1_R1162_U108 = ~new_P1_U3472 | ~new_P1_R1162_U107;
  assign new_P1_R1162_U109 = ~new_P1_R1162_U4 | ~new_P1_R1162_U106;
  assign new_P1_R1162_U110 = ~P1_REG1_REG_5_ | ~new_P1_R1162_U89;
  assign new_P1_R1162_U111 = ~new_P1_R1162_U39;
  assign new_P1_R1162_U112 = new_P1_U3478 | P1_REG1_REG_7_;
  assign new_P1_R1162_U113 = new_P1_U3475 | P1_REG1_REG_6_;
  assign new_P1_R1162_U114 = ~new_P1_R1162_U20;
  assign new_P1_R1162_U115 = ~new_P1_R1162_U21 | ~new_P1_R1162_U20;
  assign new_P1_R1162_U116 = ~new_P1_U3478 | ~new_P1_R1162_U115;
  assign new_P1_R1162_U117 = ~P1_REG1_REG_7_ | ~new_P1_R1162_U114;
  assign new_P1_R1162_U118 = ~new_P1_R1162_U6 | ~new_P1_R1162_U39;
  assign new_P1_R1162_U119 = ~new_P1_R1162_U81;
  assign new_P1_R1162_U120 = P1_REG1_REG_8_ | new_P1_U3481;
  assign new_P1_R1162_U121 = ~new_P1_R1162_U120 | ~new_P1_R1162_U81;
  assign new_P1_R1162_U122 = ~new_P1_R1162_U38;
  assign new_P1_R1162_U123 = new_P1_U3484 | P1_REG1_REG_9_;
  assign new_P1_R1162_U124 = P1_REG1_REG_6_ | new_P1_U3475;
  assign new_P1_R1162_U125 = ~new_P1_R1162_U124 | ~new_P1_R1162_U39;
  assign new_P1_R1162_U126 = ~new_P1_R1162_U125 | ~new_P1_R1162_U20 | ~new_P1_R1162_U238 | ~new_P1_R1162_U237;
  assign new_P1_R1162_U127 = ~new_P1_R1162_U111 | ~new_P1_R1162_U20;
  assign new_P1_R1162_U128 = ~P1_REG1_REG_7_ | ~new_P1_U3478;
  assign new_P1_R1162_U129 = ~new_P1_R1162_U127 | ~new_P1_R1162_U128 | ~new_P1_R1162_U6;
  assign new_P1_R1162_U130 = new_P1_U3475 | P1_REG1_REG_6_;
  assign new_P1_R1162_U131 = ~new_P1_R1162_U101 | ~new_P1_R1162_U97;
  assign new_P1_R1162_U132 = ~new_P1_U3463 | ~P1_REG1_REG_2_;
  assign new_P1_R1162_U133 = ~new_P1_R1162_U43;
  assign new_P1_R1162_U134 = ~new_P1_R1162_U100 | ~new_P1_R1162_U5;
  assign new_P1_R1162_U135 = ~new_P1_R1162_U43 | ~new_P1_R1162_U96;
  assign new_P1_R1162_U136 = ~new_P1_U3466 | ~P1_REG1_REG_3_;
  assign new_P1_R1162_U137 = ~new_P1_R1162_U42;
  assign new_P1_R1162_U138 = P1_REG1_REG_4_ | new_P1_U3469;
  assign new_P1_R1162_U139 = ~new_P1_R1162_U138 | ~new_P1_R1162_U42;
  assign new_P1_R1162_U140 = ~new_P1_R1162_U139 | ~new_P1_R1162_U32 | ~new_P1_R1162_U245 | ~new_P1_R1162_U244;
  assign new_P1_R1162_U141 = ~new_P1_R1162_U137 | ~new_P1_R1162_U32;
  assign new_P1_R1162_U142 = ~P1_REG1_REG_5_ | ~new_P1_U3472;
  assign new_P1_R1162_U143 = ~new_P1_R1162_U141 | ~new_P1_R1162_U142 | ~new_P1_R1162_U4;
  assign new_P1_R1162_U144 = new_P1_U3469 | P1_REG1_REG_4_;
  assign new_P1_R1162_U145 = ~new_P1_R1162_U100 | ~new_P1_R1162_U97;
  assign new_P1_R1162_U146 = ~new_P1_R1162_U82;
  assign new_P1_R1162_U147 = ~new_P1_U3466 | ~P1_REG1_REG_3_;
  assign new_P1_R1162_U148 = ~new_P1_R1162_U40 | ~new_P1_R1162_U41 | ~new_P1_R1162_U257 | ~new_P1_R1162_U256;
  assign new_P1_R1162_U149 = ~new_P1_R1162_U41 | ~new_P1_R1162_U40;
  assign new_P1_R1162_U150 = ~new_P1_U3463 | ~P1_REG1_REG_2_;
  assign new_P1_R1162_U151 = ~new_P1_R1162_U149 | ~new_P1_R1162_U150 | ~new_P1_R1162_U97;
  assign new_P1_R1162_U152 = P1_REG1_REG_1_ | new_P1_U3460;
  assign new_P1_R1162_U153 = ~new_P1_R1162_U83;
  assign new_P1_R1162_U154 = new_P1_U3484 | P1_REG1_REG_9_;
  assign new_P1_R1162_U155 = new_P1_U3487 | P1_REG1_REG_10_;
  assign new_P1_R1162_U156 = ~new_P1_R1162_U93 | ~new_P1_R1162_U7;
  assign new_P1_R1162_U157 = ~new_P1_U3487 | ~P1_REG1_REG_10_;
  assign new_P1_R1162_U158 = ~new_P1_R1162_U156 | ~new_P1_R1162_U157 | ~new_P1_R1162_U90;
  assign new_P1_R1162_U159 = P1_REG1_REG_10_ | new_P1_U3487;
  assign new_P1_R1162_U160 = ~new_P1_R1162_U81 | ~new_P1_R1162_U120 | ~new_P1_R1162_U7;
  assign new_P1_R1162_U161 = ~new_P1_R1162_U159 | ~new_P1_R1162_U158;
  assign new_P1_R1162_U162 = ~new_P1_R1162_U88;
  assign new_P1_R1162_U163 = new_P1_U3496 | P1_REG1_REG_13_;
  assign new_P1_R1162_U164 = new_P1_U3493 | P1_REG1_REG_12_;
  assign new_P1_R1162_U165 = ~new_P1_R1162_U92 | ~new_P1_R1162_U8;
  assign new_P1_R1162_U166 = ~new_P1_U3496 | ~P1_REG1_REG_13_;
  assign new_P1_R1162_U167 = ~new_P1_R1162_U165 | ~new_P1_R1162_U166 | ~new_P1_R1162_U91;
  assign new_P1_R1162_U168 = P1_REG1_REG_11_ | new_P1_U3490;
  assign new_P1_R1162_U169 = P1_REG1_REG_13_ | new_P1_U3496;
  assign new_P1_R1162_U170 = ~new_P1_R1162_U88 | ~new_P1_R1162_U168 | ~new_P1_R1162_U8;
  assign new_P1_R1162_U171 = ~new_P1_R1162_U169 | ~new_P1_R1162_U167;
  assign new_P1_R1162_U172 = ~new_P1_R1162_U87;
  assign new_P1_R1162_U173 = P1_REG1_REG_14_ | new_P1_U3499;
  assign new_P1_R1162_U174 = ~new_P1_R1162_U173 | ~new_P1_R1162_U87;
  assign new_P1_R1162_U175 = ~new_P1_U3499 | ~P1_REG1_REG_14_;
  assign new_P1_R1162_U176 = ~new_P1_R1162_U86;
  assign new_P1_R1162_U177 = P1_REG1_REG_15_ | new_P1_U3502;
  assign new_P1_R1162_U178 = ~new_P1_R1162_U177 | ~new_P1_R1162_U86;
  assign new_P1_R1162_U179 = ~new_P1_U3502 | ~P1_REG1_REG_15_;
  assign new_P1_R1162_U180 = ~new_P1_R1162_U66;
  assign new_P1_R1162_U181 = new_P1_U3508 | P1_REG1_REG_17_;
  assign new_P1_R1162_U182 = new_P1_U3505 | P1_REG1_REG_16_;
  assign new_P1_R1162_U183 = ~new_P1_R1162_U47;
  assign new_P1_R1162_U184 = ~new_P1_R1162_U48 | ~new_P1_R1162_U47;
  assign new_P1_R1162_U185 = ~new_P1_U3508 | ~new_P1_R1162_U184;
  assign new_P1_R1162_U186 = ~P1_REG1_REG_17_ | ~new_P1_R1162_U183;
  assign new_P1_R1162_U187 = ~new_P1_R1162_U9 | ~new_P1_R1162_U66;
  assign new_P1_R1162_U188 = ~new_P1_R1162_U65;
  assign new_P1_R1162_U189 = P1_REG1_REG_18_ | new_P1_U3511;
  assign new_P1_R1162_U190 = ~new_P1_R1162_U189 | ~new_P1_R1162_U65;
  assign new_P1_R1162_U191 = ~new_P1_U3511 | ~P1_REG1_REG_18_;
  assign new_P1_R1162_U192 = ~new_P1_R1162_U190 | ~new_P1_R1162_U191 | ~new_P1_R1162_U261 | ~new_P1_R1162_U260;
  assign new_P1_R1162_U193 = ~new_P1_U3511 | ~P1_REG1_REG_18_;
  assign new_P1_R1162_U194 = ~new_P1_R1162_U188 | ~new_P1_R1162_U193;
  assign new_P1_R1162_U195 = new_P1_U3511 | P1_REG1_REG_18_;
  assign new_P1_R1162_U196 = ~new_P1_R1162_U194 | ~new_P1_R1162_U195 | ~new_P1_R1162_U264;
  assign new_P1_R1162_U197 = P1_REG1_REG_16_ | new_P1_U3505;
  assign new_P1_R1162_U198 = ~new_P1_R1162_U197 | ~new_P1_R1162_U66;
  assign new_P1_R1162_U199 = ~new_P1_R1162_U198 | ~new_P1_R1162_U47 | ~new_P1_R1162_U273 | ~new_P1_R1162_U272;
  assign new_P1_R1162_U200 = ~new_P1_R1162_U180 | ~new_P1_R1162_U47;
  assign new_P1_R1162_U201 = ~P1_REG1_REG_17_ | ~new_P1_U3508;
  assign new_P1_R1162_U202 = ~new_P1_R1162_U200 | ~new_P1_R1162_U201 | ~new_P1_R1162_U9;
  assign new_P1_R1162_U203 = new_P1_U3505 | P1_REG1_REG_16_;
  assign new_P1_R1162_U204 = ~new_P1_R1162_U168 | ~new_P1_R1162_U88;
  assign new_P1_R1162_U205 = ~new_P1_R1162_U67;
  assign new_P1_R1162_U206 = P1_REG1_REG_12_ | new_P1_U3493;
  assign new_P1_R1162_U207 = ~new_P1_R1162_U206 | ~new_P1_R1162_U67;
  assign new_P1_R1162_U208 = ~new_P1_R1162_U207 | ~new_P1_R1162_U91 | ~new_P1_R1162_U294 | ~new_P1_R1162_U293;
  assign new_P1_R1162_U209 = ~new_P1_R1162_U205 | ~new_P1_R1162_U91;
  assign new_P1_R1162_U210 = ~new_P1_U3496 | ~P1_REG1_REG_13_;
  assign new_P1_R1162_U211 = ~new_P1_R1162_U209 | ~new_P1_R1162_U210 | ~new_P1_R1162_U8;
  assign new_P1_R1162_U212 = new_P1_U3493 | P1_REG1_REG_12_;
  assign new_P1_R1162_U213 = P1_REG1_REG_9_ | new_P1_U3484;
  assign new_P1_R1162_U214 = ~new_P1_R1162_U213 | ~new_P1_R1162_U38;
  assign new_P1_R1162_U215 = ~new_P1_R1162_U214 | ~new_P1_R1162_U90 | ~new_P1_R1162_U306 | ~new_P1_R1162_U305;
  assign new_P1_R1162_U216 = ~new_P1_R1162_U122 | ~new_P1_R1162_U90;
  assign new_P1_R1162_U217 = ~new_P1_U3487 | ~P1_REG1_REG_10_;
  assign new_P1_R1162_U218 = ~new_P1_R1162_U216 | ~new_P1_R1162_U217 | ~new_P1_R1162_U7;
  assign new_P1_R1162_U219 = ~new_P1_R1162_U123 | ~new_P1_R1162_U90;
  assign new_P1_R1162_U220 = ~new_P1_R1162_U120 | ~new_P1_R1162_U49;
  assign new_P1_R1162_U221 = ~new_P1_R1162_U130 | ~new_P1_R1162_U20;
  assign new_P1_R1162_U222 = ~new_P1_R1162_U144 | ~new_P1_R1162_U32;
  assign new_P1_R1162_U223 = ~new_P1_R1162_U147 | ~new_P1_R1162_U96;
  assign new_P1_R1162_U224 = ~new_P1_R1162_U203 | ~new_P1_R1162_U47;
  assign new_P1_R1162_U225 = ~new_P1_R1162_U212 | ~new_P1_R1162_U91;
  assign new_P1_R1162_U226 = ~new_P1_R1162_U168 | ~new_P1_R1162_U56;
  assign new_P1_R1162_U227 = ~new_P1_U3484 | ~new_P1_R1162_U37;
  assign new_P1_R1162_U228 = ~P1_REG1_REG_9_ | ~new_P1_R1162_U36;
  assign new_P1_R1162_U229 = ~new_P1_R1162_U228 | ~new_P1_R1162_U227;
  assign new_P1_R1162_U230 = ~new_P1_R1162_U219 | ~new_P1_R1162_U38;
  assign new_P1_R1162_U231 = ~new_P1_R1162_U229 | ~new_P1_R1162_U122;
  assign new_P1_R1162_U232 = ~new_P1_U3481 | ~new_P1_R1162_U34;
  assign new_P1_R1162_U233 = ~P1_REG1_REG_8_ | ~new_P1_R1162_U35;
  assign new_P1_R1162_U234 = ~new_P1_R1162_U233 | ~new_P1_R1162_U232;
  assign new_P1_R1162_U235 = ~new_P1_R1162_U220 | ~new_P1_R1162_U81;
  assign new_P1_R1162_U236 = ~new_P1_R1162_U119 | ~new_P1_R1162_U234;
  assign new_P1_R1162_U237 = ~new_P1_U3478 | ~new_P1_R1162_U21;
  assign new_P1_R1162_U238 = ~P1_REG1_REG_7_ | ~new_P1_R1162_U19;
  assign new_P1_R1162_U239 = ~new_P1_U3475 | ~new_P1_R1162_U17;
  assign new_P1_R1162_U240 = ~P1_REG1_REG_6_ | ~new_P1_R1162_U18;
  assign new_P1_R1162_U241 = ~new_P1_R1162_U240 | ~new_P1_R1162_U239;
  assign new_P1_R1162_U242 = ~new_P1_R1162_U221 | ~new_P1_R1162_U39;
  assign new_P1_R1162_U243 = ~new_P1_R1162_U241 | ~new_P1_R1162_U111;
  assign new_P1_R1162_U244 = ~new_P1_U3472 | ~new_P1_R1162_U33;
  assign new_P1_R1162_U245 = ~P1_REG1_REG_5_ | ~new_P1_R1162_U24;
  assign new_P1_R1162_U246 = ~new_P1_U3469 | ~new_P1_R1162_U22;
  assign new_P1_R1162_U247 = ~P1_REG1_REG_4_ | ~new_P1_R1162_U23;
  assign new_P1_R1162_U248 = ~new_P1_R1162_U247 | ~new_P1_R1162_U246;
  assign new_P1_R1162_U249 = ~new_P1_R1162_U222 | ~new_P1_R1162_U42;
  assign new_P1_R1162_U250 = ~new_P1_R1162_U248 | ~new_P1_R1162_U137;
  assign new_P1_R1162_U251 = ~new_P1_U3466 | ~new_P1_R1162_U30;
  assign new_P1_R1162_U252 = ~P1_REG1_REG_3_ | ~new_P1_R1162_U31;
  assign new_P1_R1162_U253 = ~new_P1_R1162_U252 | ~new_P1_R1162_U251;
  assign new_P1_R1162_U254 = ~new_P1_R1162_U223 | ~new_P1_R1162_U82;
  assign new_P1_R1162_U255 = ~new_P1_R1162_U146 | ~new_P1_R1162_U253;
  assign new_P1_R1162_U256 = ~new_P1_U3463 | ~new_P1_R1162_U25;
  assign new_P1_R1162_U257 = ~P1_REG1_REG_2_ | ~new_P1_R1162_U26;
  assign new_P1_R1162_U258 = ~new_P1_R1162_U98 | ~new_P1_R1162_U83;
  assign new_P1_R1162_U259 = ~new_P1_R1162_U153 | ~new_P1_R1162_U29;
  assign new_P1_R1162_U260 = ~new_P1_U3452 | ~new_P1_R1162_U85;
  assign new_P1_R1162_U261 = ~P1_REG1_REG_19_ | ~new_P1_R1162_U84;
  assign new_P1_R1162_U262 = ~new_P1_U3452 | ~new_P1_R1162_U85;
  assign new_P1_R1162_U263 = ~P1_REG1_REG_19_ | ~new_P1_R1162_U84;
  assign new_P1_R1162_U264 = ~new_P1_R1162_U263 | ~new_P1_R1162_U262;
  assign new_P1_R1162_U265 = ~new_P1_U3511 | ~new_P1_R1162_U63;
  assign new_P1_R1162_U266 = ~P1_REG1_REG_18_ | ~new_P1_R1162_U64;
  assign new_P1_R1162_U267 = ~new_P1_U3511 | ~new_P1_R1162_U63;
  assign new_P1_R1162_U268 = ~P1_REG1_REG_18_ | ~new_P1_R1162_U64;
  assign new_P1_R1162_U269 = ~new_P1_R1162_U268 | ~new_P1_R1162_U267;
  assign new_P1_R1162_U270 = ~new_P1_R1162_U65 | ~new_P1_R1162_U266 | ~new_P1_R1162_U265;
  assign new_P1_R1162_U271 = ~new_P1_R1162_U269 | ~new_P1_R1162_U188;
  assign new_P1_R1162_U272 = ~new_P1_U3508 | ~new_P1_R1162_U48;
  assign new_P1_R1162_U273 = ~P1_REG1_REG_17_ | ~new_P1_R1162_U46;
  assign new_P1_R1162_U274 = ~new_P1_U3505 | ~new_P1_R1162_U44;
  assign new_P1_R1162_U275 = ~P1_REG1_REG_16_ | ~new_P1_R1162_U45;
  assign new_P1_R1162_U276 = ~new_P1_R1162_U275 | ~new_P1_R1162_U274;
  assign new_P1_R1162_U277 = ~new_P1_R1162_U224 | ~new_P1_R1162_U66;
  assign new_P1_R1162_U278 = ~new_P1_R1162_U276 | ~new_P1_R1162_U180;
  assign new_P1_R1162_U279 = ~new_P1_U3502 | ~new_P1_R1162_U61;
  assign new_P1_R1162_U280 = ~P1_REG1_REG_15_ | ~new_P1_R1162_U62;
  assign new_P1_R1162_U281 = ~new_P1_U3502 | ~new_P1_R1162_U61;
  assign new_P1_R1162_U282 = ~P1_REG1_REG_15_ | ~new_P1_R1162_U62;
  assign new_P1_R1162_U283 = ~new_P1_R1162_U282 | ~new_P1_R1162_U281;
  assign new_P1_R1162_U284 = ~new_P1_R1162_U86 | ~new_P1_R1162_U280 | ~new_P1_R1162_U279;
  assign new_P1_R1162_U285 = ~new_P1_R1162_U176 | ~new_P1_R1162_U283;
  assign new_P1_R1162_U286 = ~new_P1_U3499 | ~new_P1_R1162_U59;
  assign new_P1_R1162_U287 = ~P1_REG1_REG_14_ | ~new_P1_R1162_U60;
  assign new_P1_R1162_U288 = ~new_P1_U3499 | ~new_P1_R1162_U59;
  assign new_P1_R1162_U289 = ~P1_REG1_REG_14_ | ~new_P1_R1162_U60;
  assign new_P1_R1162_U290 = ~new_P1_R1162_U289 | ~new_P1_R1162_U288;
  assign new_P1_R1162_U291 = ~new_P1_R1162_U87 | ~new_P1_R1162_U287 | ~new_P1_R1162_U286;
  assign new_P1_R1162_U292 = ~new_P1_R1162_U172 | ~new_P1_R1162_U290;
  assign new_P1_R1162_U293 = ~new_P1_U3496 | ~new_P1_R1162_U57;
  assign new_P1_R1162_U294 = ~P1_REG1_REG_13_ | ~new_P1_R1162_U58;
  assign new_P1_R1162_U295 = ~new_P1_U3493 | ~new_P1_R1162_U52;
  assign new_P1_R1162_U296 = ~P1_REG1_REG_12_ | ~new_P1_R1162_U53;
  assign new_P1_R1162_U297 = ~new_P1_R1162_U296 | ~new_P1_R1162_U295;
  assign new_P1_R1162_U298 = ~new_P1_R1162_U225 | ~new_P1_R1162_U67;
  assign new_P1_R1162_U299 = ~new_P1_R1162_U297 | ~new_P1_R1162_U205;
  assign new_P1_R1162_U300 = ~new_P1_U3490 | ~new_P1_R1162_U54;
  assign new_P1_R1162_U301 = ~P1_REG1_REG_11_ | ~new_P1_R1162_U55;
  assign new_P1_R1162_U302 = ~new_P1_R1162_U301 | ~new_P1_R1162_U300;
  assign new_P1_R1162_U303 = ~new_P1_R1162_U226 | ~new_P1_R1162_U88;
  assign new_P1_R1162_U304 = ~new_P1_R1162_U162 | ~new_P1_R1162_U302;
  assign new_P1_R1162_U305 = ~new_P1_U3487 | ~new_P1_R1162_U50;
  assign new_P1_R1162_U306 = ~P1_REG1_REG_10_ | ~new_P1_R1162_U51;
  assign new_P1_R1162_U307 = ~new_P1_U3454 | ~new_P1_R1162_U27;
  assign new_P1_R1162_U308 = ~P1_REG1_REG_0_ | ~new_P1_R1162_U28;
  assign new_P1_R1117_U6 = new_P1_R1117_U184 & new_P1_R1117_U201;
  assign new_P1_R1117_U7 = new_P1_R1117_U203 & new_P1_R1117_U202;
  assign new_P1_R1117_U8 = new_P1_R1117_U179 & new_P1_R1117_U240;
  assign new_P1_R1117_U9 = new_P1_R1117_U242 & new_P1_R1117_U241;
  assign new_P1_R1117_U10 = new_P1_R1117_U259 & new_P1_R1117_U258;
  assign new_P1_R1117_U11 = new_P1_R1117_U285 & new_P1_R1117_U284;
  assign new_P1_R1117_U12 = new_P1_R1117_U383 & new_P1_R1117_U382;
  assign new_P1_R1117_U13 = ~new_P1_R1117_U340 | ~new_P1_R1117_U343;
  assign new_P1_R1117_U14 = ~new_P1_R1117_U329 | ~new_P1_R1117_U332;
  assign new_P1_R1117_U15 = ~new_P1_R1117_U318 | ~new_P1_R1117_U321;
  assign new_P1_R1117_U16 = ~new_P1_R1117_U310 | ~new_P1_R1117_U312;
  assign new_P1_R1117_U17 = ~new_P1_R1117_U348 | ~new_P1_R1117_U156 | ~new_P1_R1117_U175;
  assign new_P1_R1117_U18 = ~new_P1_R1117_U236 | ~new_P1_R1117_U238;
  assign new_P1_R1117_U19 = ~new_P1_R1117_U228 | ~new_P1_R1117_U231;
  assign new_P1_R1117_U20 = ~new_P1_R1117_U220 | ~new_P1_R1117_U222;
  assign new_P1_R1117_U21 = ~new_P1_R1117_U25 | ~new_P1_R1117_U346;
  assign new_P1_R1117_U22 = ~new_P1_U3479;
  assign new_P1_R1117_U23 = ~new_P1_U3464;
  assign new_P1_R1117_U24 = ~new_P1_U3456;
  assign new_P1_R1117_U25 = ~new_P1_U3456 | ~new_P1_R1117_U93;
  assign new_P1_R1117_U26 = ~new_P1_U3078;
  assign new_P1_R1117_U27 = ~new_P1_U3467;
  assign new_P1_R1117_U28 = ~new_P1_U3068;
  assign new_P1_R1117_U29 = ~new_P1_U3068 | ~new_P1_R1117_U23;
  assign new_P1_R1117_U30 = ~new_P1_U3064;
  assign new_P1_R1117_U31 = ~new_P1_U3476;
  assign new_P1_R1117_U32 = ~new_P1_U3473;
  assign new_P1_R1117_U33 = ~new_P1_U3470;
  assign new_P1_R1117_U34 = ~new_P1_U3071;
  assign new_P1_R1117_U35 = ~new_P1_U3067;
  assign new_P1_R1117_U36 = ~new_P1_U3060;
  assign new_P1_R1117_U37 = ~new_P1_U3060 | ~new_P1_R1117_U33;
  assign new_P1_R1117_U38 = ~new_P1_U3482;
  assign new_P1_R1117_U39 = ~new_P1_U3070;
  assign new_P1_R1117_U40 = ~new_P1_U3070 | ~new_P1_R1117_U22;
  assign new_P1_R1117_U41 = ~new_P1_U3084;
  assign new_P1_R1117_U42 = ~new_P1_U3485;
  assign new_P1_R1117_U43 = ~new_P1_U3083;
  assign new_P1_R1117_U44 = ~new_P1_R1117_U209 | ~new_P1_R1117_U208;
  assign new_P1_R1117_U45 = ~new_P1_R1117_U37 | ~new_P1_R1117_U224;
  assign new_P1_R1117_U46 = ~new_P1_R1117_U193 | ~new_P1_R1117_U192;
  assign new_P1_R1117_U47 = ~new_P1_U4019;
  assign new_P1_R1117_U48 = ~new_P1_U4023;
  assign new_P1_R1117_U49 = ~new_P1_U3503;
  assign new_P1_R1117_U50 = ~new_P1_U3491;
  assign new_P1_R1117_U51 = ~new_P1_U3488;
  assign new_P1_R1117_U52 = ~new_P1_U3063;
  assign new_P1_R1117_U53 = ~new_P1_U3062;
  assign new_P1_R1117_U54 = ~new_P1_U3083 | ~new_P1_R1117_U42;
  assign new_P1_R1117_U55 = ~new_P1_U3494;
  assign new_P1_R1117_U56 = ~new_P1_U3072;
  assign new_P1_R1117_U57 = ~new_P1_U3497;
  assign new_P1_R1117_U58 = ~new_P1_U3080;
  assign new_P1_R1117_U59 = ~new_P1_U3506;
  assign new_P1_R1117_U60 = ~new_P1_U3500;
  assign new_P1_R1117_U61 = ~new_P1_U3073;
  assign new_P1_R1117_U62 = ~new_P1_U3074;
  assign new_P1_R1117_U63 = ~new_P1_U3079;
  assign new_P1_R1117_U64 = ~new_P1_U3079 | ~new_P1_R1117_U60;
  assign new_P1_R1117_U65 = ~new_P1_U3509;
  assign new_P1_R1117_U66 = ~new_P1_U3069;
  assign new_P1_R1117_U67 = ~new_P1_R1117_U269 | ~new_P1_R1117_U268;
  assign new_P1_R1117_U68 = ~new_P1_U3082;
  assign new_P1_R1117_U69 = ~new_P1_U3514;
  assign new_P1_R1117_U70 = ~new_P1_U3081;
  assign new_P1_R1117_U71 = ~new_P1_U4025;
  assign new_P1_R1117_U72 = ~new_P1_U3076;
  assign new_P1_R1117_U73 = ~new_P1_U4022;
  assign new_P1_R1117_U74 = ~new_P1_U4024;
  assign new_P1_R1117_U75 = ~new_P1_U3066;
  assign new_P1_R1117_U76 = ~new_P1_U3061;
  assign new_P1_R1117_U77 = ~new_P1_U3075;
  assign new_P1_R1117_U78 = ~new_P1_U3075 | ~new_P1_R1117_U74;
  assign new_P1_R1117_U79 = ~new_P1_U4021;
  assign new_P1_R1117_U80 = ~new_P1_U3065;
  assign new_P1_R1117_U81 = ~new_P1_U4020;
  assign new_P1_R1117_U82 = ~new_P1_U3058;
  assign new_P1_R1117_U83 = ~new_P1_U4018;
  assign new_P1_R1117_U84 = ~new_P1_U3057;
  assign new_P1_R1117_U85 = ~new_P1_U3057 | ~new_P1_R1117_U47;
  assign new_P1_R1117_U86 = ~new_P1_U3053;
  assign new_P1_R1117_U87 = ~new_P1_U4017;
  assign new_P1_R1117_U88 = ~new_P1_U3054;
  assign new_P1_R1117_U89 = ~new_P1_R1117_U299 | ~new_P1_R1117_U298;
  assign new_P1_R1117_U90 = ~new_P1_R1117_U78 | ~new_P1_R1117_U314;
  assign new_P1_R1117_U91 = ~new_P1_R1117_U64 | ~new_P1_R1117_U325;
  assign new_P1_R1117_U92 = ~new_P1_R1117_U54 | ~new_P1_R1117_U336;
  assign new_P1_R1117_U93 = ~new_P1_U3077;
  assign new_P1_R1117_U94 = ~new_P1_R1117_U393 | ~new_P1_R1117_U392;
  assign new_P1_R1117_U95 = ~new_P1_R1117_U407 | ~new_P1_R1117_U406;
  assign new_P1_R1117_U96 = ~new_P1_R1117_U412 | ~new_P1_R1117_U411;
  assign new_P1_R1117_U97 = ~new_P1_R1117_U428 | ~new_P1_R1117_U427;
  assign new_P1_R1117_U98 = ~new_P1_R1117_U433 | ~new_P1_R1117_U432;
  assign new_P1_R1117_U99 = ~new_P1_R1117_U438 | ~new_P1_R1117_U437;
  assign new_P1_R1117_U100 = ~new_P1_R1117_U443 | ~new_P1_R1117_U442;
  assign new_P1_R1117_U101 = ~new_P1_R1117_U448 | ~new_P1_R1117_U447;
  assign new_P1_R1117_U102 = ~new_P1_R1117_U464 | ~new_P1_R1117_U463;
  assign new_P1_R1117_U103 = ~new_P1_R1117_U469 | ~new_P1_R1117_U468;
  assign new_P1_R1117_U104 = ~new_P1_R1117_U352 | ~new_P1_R1117_U351;
  assign new_P1_R1117_U105 = ~new_P1_R1117_U361 | ~new_P1_R1117_U360;
  assign new_P1_R1117_U106 = ~new_P1_R1117_U368 | ~new_P1_R1117_U367;
  assign new_P1_R1117_U107 = ~new_P1_R1117_U372 | ~new_P1_R1117_U371;
  assign new_P1_R1117_U108 = ~new_P1_R1117_U381 | ~new_P1_R1117_U380;
  assign new_P1_R1117_U109 = ~new_P1_R1117_U402 | ~new_P1_R1117_U401;
  assign new_P1_R1117_U110 = ~new_P1_R1117_U419 | ~new_P1_R1117_U418;
  assign new_P1_R1117_U111 = ~new_P1_R1117_U423 | ~new_P1_R1117_U422;
  assign new_P1_R1117_U112 = ~new_P1_R1117_U455 | ~new_P1_R1117_U454;
  assign new_P1_R1117_U113 = ~new_P1_R1117_U459 | ~new_P1_R1117_U458;
  assign new_P1_R1117_U114 = ~new_P1_R1117_U476 | ~new_P1_R1117_U475;
  assign new_P1_R1117_U115 = new_P1_R1117_U195 & new_P1_R1117_U183;
  assign new_P1_R1117_U116 = new_P1_R1117_U198 & new_P1_R1117_U199;
  assign new_P1_R1117_U117 = new_P1_R1117_U211 & new_P1_R1117_U185;
  assign new_P1_R1117_U118 = new_P1_R1117_U214 & new_P1_R1117_U215;
  assign new_P1_R1117_U119 = new_P1_R1117_U40 & new_P1_R1117_U354 & new_P1_R1117_U353;
  assign new_P1_R1117_U120 = new_P1_R1117_U357 & new_P1_R1117_U185;
  assign new_P1_R1117_U121 = new_P1_R1117_U230 & new_P1_R1117_U7;
  assign new_P1_R1117_U122 = new_P1_R1117_U364 & new_P1_R1117_U184;
  assign new_P1_R1117_U123 = new_P1_R1117_U29 & new_P1_R1117_U374 & new_P1_R1117_U373;
  assign new_P1_R1117_U124 = new_P1_R1117_U377 & new_P1_R1117_U183;
  assign new_P1_R1117_U125 = new_P1_R1117_U217 & new_P1_R1117_U8;
  assign new_P1_R1117_U126 = new_P1_R1117_U262 & new_P1_R1117_U180;
  assign new_P1_R1117_U127 = new_P1_R1117_U288 & new_P1_R1117_U181;
  assign new_P1_R1117_U128 = new_P1_R1117_U304 & new_P1_R1117_U305;
  assign new_P1_R1117_U129 = new_P1_R1117_U307 & new_P1_R1117_U386;
  assign new_P1_R1117_U130 = new_P1_R1117_U308 & new_P1_R1117_U305 & new_P1_R1117_U304;
  assign new_P1_R1117_U131 = ~new_P1_R1117_U390 | ~new_P1_R1117_U389;
  assign new_P1_R1117_U132 = new_P1_R1117_U85 & new_P1_R1117_U395 & new_P1_R1117_U394;
  assign new_P1_R1117_U133 = new_P1_R1117_U398 & new_P1_R1117_U182;
  assign new_P1_R1117_U134 = ~new_P1_R1117_U404 | ~new_P1_R1117_U403;
  assign new_P1_R1117_U135 = ~new_P1_R1117_U409 | ~new_P1_R1117_U408;
  assign new_P1_R1117_U136 = new_P1_R1117_U415 & new_P1_R1117_U181;
  assign new_P1_R1117_U137 = ~new_P1_R1117_U425 | ~new_P1_R1117_U424;
  assign new_P1_R1117_U138 = ~new_P1_R1117_U430 | ~new_P1_R1117_U429;
  assign new_P1_R1117_U139 = ~new_P1_R1117_U435 | ~new_P1_R1117_U434;
  assign new_P1_R1117_U140 = ~new_P1_R1117_U440 | ~new_P1_R1117_U439;
  assign new_P1_R1117_U141 = ~new_P1_R1117_U445 | ~new_P1_R1117_U444;
  assign new_P1_R1117_U142 = new_P1_R1117_U451 & new_P1_R1117_U180;
  assign new_P1_R1117_U143 = ~new_P1_R1117_U461 | ~new_P1_R1117_U460;
  assign new_P1_R1117_U144 = ~new_P1_R1117_U466 | ~new_P1_R1117_U465;
  assign new_P1_R1117_U145 = new_P1_R1117_U342 & new_P1_R1117_U9;
  assign new_P1_R1117_U146 = new_P1_R1117_U472 & new_P1_R1117_U179;
  assign new_P1_R1117_U147 = new_P1_R1117_U350 & new_P1_R1117_U349;
  assign new_P1_R1117_U148 = ~new_P1_R1117_U118 | ~new_P1_R1117_U212;
  assign new_P1_R1117_U149 = new_P1_R1117_U359 & new_P1_R1117_U358;
  assign new_P1_R1117_U150 = new_P1_R1117_U366 & new_P1_R1117_U365;
  assign new_P1_R1117_U151 = new_P1_R1117_U370 & new_P1_R1117_U369;
  assign new_P1_R1117_U152 = ~new_P1_R1117_U116 | ~new_P1_R1117_U196;
  assign new_P1_R1117_U153 = new_P1_R1117_U379 & new_P1_R1117_U378;
  assign new_P1_R1117_U154 = ~new_P1_U4028;
  assign new_P1_R1117_U155 = ~new_P1_U3055;
  assign new_P1_R1117_U156 = new_P1_R1117_U388 & new_P1_R1117_U387;
  assign new_P1_R1117_U157 = ~new_P1_R1117_U128 | ~new_P1_R1117_U302;
  assign new_P1_R1117_U158 = new_P1_R1117_U400 & new_P1_R1117_U399;
  assign new_P1_R1117_U159 = ~new_P1_R1117_U295 | ~new_P1_R1117_U294;
  assign new_P1_R1117_U160 = ~new_P1_R1117_U291 | ~new_P1_R1117_U290;
  assign new_P1_R1117_U161 = new_P1_R1117_U417 & new_P1_R1117_U416;
  assign new_P1_R1117_U162 = new_P1_R1117_U421 & new_P1_R1117_U420;
  assign new_P1_R1117_U163 = ~new_P1_R1117_U281 | ~new_P1_R1117_U280;
  assign new_P1_R1117_U164 = ~new_P1_R1117_U277 | ~new_P1_R1117_U276;
  assign new_P1_R1117_U165 = ~new_P1_U3461;
  assign new_P1_R1117_U166 = ~new_P1_R1117_U273 | ~new_P1_R1117_U272;
  assign new_P1_R1117_U167 = ~new_P1_U3512;
  assign new_P1_R1117_U168 = ~new_P1_R1117_U265 | ~new_P1_R1117_U264;
  assign new_P1_R1117_U169 = new_P1_R1117_U453 & new_P1_R1117_U452;
  assign new_P1_R1117_U170 = new_P1_R1117_U457 & new_P1_R1117_U456;
  assign new_P1_R1117_U171 = ~new_P1_R1117_U255 | ~new_P1_R1117_U254;
  assign new_P1_R1117_U172 = ~new_P1_R1117_U251 | ~new_P1_R1117_U250;
  assign new_P1_R1117_U173 = ~new_P1_R1117_U247 | ~new_P1_R1117_U246;
  assign new_P1_R1117_U174 = new_P1_R1117_U474 & new_P1_R1117_U473;
  assign new_P1_R1117_U175 = ~new_P1_R1117_U129 | ~new_P1_R1117_U157;
  assign new_P1_R1117_U176 = ~new_P1_R1117_U85;
  assign new_P1_R1117_U177 = ~new_P1_R1117_U29;
  assign new_P1_R1117_U178 = ~new_P1_R1117_U40;
  assign new_P1_R1117_U179 = ~new_P1_U3488 | ~new_P1_R1117_U53;
  assign new_P1_R1117_U180 = ~new_P1_U3503 | ~new_P1_R1117_U62;
  assign new_P1_R1117_U181 = ~new_P1_U4023 | ~new_P1_R1117_U76;
  assign new_P1_R1117_U182 = ~new_P1_U4019 | ~new_P1_R1117_U84;
  assign new_P1_R1117_U183 = ~new_P1_U3464 | ~new_P1_R1117_U28;
  assign new_P1_R1117_U184 = ~new_P1_U3473 | ~new_P1_R1117_U35;
  assign new_P1_R1117_U185 = ~new_P1_U3479 | ~new_P1_R1117_U39;
  assign new_P1_R1117_U186 = ~new_P1_R1117_U64;
  assign new_P1_R1117_U187 = ~new_P1_R1117_U78;
  assign new_P1_R1117_U188 = ~new_P1_R1117_U37;
  assign new_P1_R1117_U189 = ~new_P1_R1117_U54;
  assign new_P1_R1117_U190 = ~new_P1_R1117_U25;
  assign new_P1_R1117_U191 = ~new_P1_R1117_U190 | ~new_P1_R1117_U26;
  assign new_P1_R1117_U192 = ~new_P1_R1117_U191 | ~new_P1_R1117_U165;
  assign new_P1_R1117_U193 = ~new_P1_U3078 | ~new_P1_R1117_U25;
  assign new_P1_R1117_U194 = ~new_P1_R1117_U46;
  assign new_P1_R1117_U195 = ~new_P1_U3467 | ~new_P1_R1117_U30;
  assign new_P1_R1117_U196 = ~new_P1_R1117_U115 | ~new_P1_R1117_U46;
  assign new_P1_R1117_U197 = ~new_P1_R1117_U30 | ~new_P1_R1117_U29;
  assign new_P1_R1117_U198 = ~new_P1_R1117_U197 | ~new_P1_R1117_U27;
  assign new_P1_R1117_U199 = ~new_P1_U3064 | ~new_P1_R1117_U177;
  assign new_P1_R1117_U200 = ~new_P1_R1117_U152;
  assign new_P1_R1117_U201 = ~new_P1_U3476 | ~new_P1_R1117_U34;
  assign new_P1_R1117_U202 = ~new_P1_U3071 | ~new_P1_R1117_U31;
  assign new_P1_R1117_U203 = ~new_P1_U3067 | ~new_P1_R1117_U32;
  assign new_P1_R1117_U204 = ~new_P1_R1117_U188 | ~new_P1_R1117_U6;
  assign new_P1_R1117_U205 = ~new_P1_R1117_U7 | ~new_P1_R1117_U204;
  assign new_P1_R1117_U206 = ~new_P1_U3470 | ~new_P1_R1117_U36;
  assign new_P1_R1117_U207 = ~new_P1_U3476 | ~new_P1_R1117_U34;
  assign new_P1_R1117_U208 = ~new_P1_R1117_U6 | ~new_P1_R1117_U206 | ~new_P1_R1117_U152;
  assign new_P1_R1117_U209 = ~new_P1_R1117_U207 | ~new_P1_R1117_U205;
  assign new_P1_R1117_U210 = ~new_P1_R1117_U44;
  assign new_P1_R1117_U211 = ~new_P1_U3482 | ~new_P1_R1117_U41;
  assign new_P1_R1117_U212 = ~new_P1_R1117_U117 | ~new_P1_R1117_U44;
  assign new_P1_R1117_U213 = ~new_P1_R1117_U41 | ~new_P1_R1117_U40;
  assign new_P1_R1117_U214 = ~new_P1_R1117_U213 | ~new_P1_R1117_U38;
  assign new_P1_R1117_U215 = ~new_P1_U3084 | ~new_P1_R1117_U178;
  assign new_P1_R1117_U216 = ~new_P1_R1117_U148;
  assign new_P1_R1117_U217 = ~new_P1_U3485 | ~new_P1_R1117_U43;
  assign new_P1_R1117_U218 = ~new_P1_R1117_U217 | ~new_P1_R1117_U54;
  assign new_P1_R1117_U219 = ~new_P1_R1117_U210 | ~new_P1_R1117_U40;
  assign new_P1_R1117_U220 = ~new_P1_R1117_U120 | ~new_P1_R1117_U219;
  assign new_P1_R1117_U221 = ~new_P1_R1117_U44 | ~new_P1_R1117_U185;
  assign new_P1_R1117_U222 = ~new_P1_R1117_U119 | ~new_P1_R1117_U221;
  assign new_P1_R1117_U223 = ~new_P1_R1117_U40 | ~new_P1_R1117_U185;
  assign new_P1_R1117_U224 = ~new_P1_R1117_U206 | ~new_P1_R1117_U152;
  assign new_P1_R1117_U225 = ~new_P1_R1117_U45;
  assign new_P1_R1117_U226 = ~new_P1_U3067 | ~new_P1_R1117_U32;
  assign new_P1_R1117_U227 = ~new_P1_R1117_U225 | ~new_P1_R1117_U226;
  assign new_P1_R1117_U228 = ~new_P1_R1117_U122 | ~new_P1_R1117_U227;
  assign new_P1_R1117_U229 = ~new_P1_R1117_U45 | ~new_P1_R1117_U184;
  assign new_P1_R1117_U230 = ~new_P1_U3476 | ~new_P1_R1117_U34;
  assign new_P1_R1117_U231 = ~new_P1_R1117_U121 | ~new_P1_R1117_U229;
  assign new_P1_R1117_U232 = ~new_P1_U3067 | ~new_P1_R1117_U32;
  assign new_P1_R1117_U233 = ~new_P1_R1117_U184 | ~new_P1_R1117_U232;
  assign new_P1_R1117_U234 = ~new_P1_R1117_U206 | ~new_P1_R1117_U37;
  assign new_P1_R1117_U235 = ~new_P1_R1117_U194 | ~new_P1_R1117_U29;
  assign new_P1_R1117_U236 = ~new_P1_R1117_U124 | ~new_P1_R1117_U235;
  assign new_P1_R1117_U237 = ~new_P1_R1117_U46 | ~new_P1_R1117_U183;
  assign new_P1_R1117_U238 = ~new_P1_R1117_U123 | ~new_P1_R1117_U237;
  assign new_P1_R1117_U239 = ~new_P1_R1117_U29 | ~new_P1_R1117_U183;
  assign new_P1_R1117_U240 = ~new_P1_U3491 | ~new_P1_R1117_U52;
  assign new_P1_R1117_U241 = ~new_P1_U3063 | ~new_P1_R1117_U50;
  assign new_P1_R1117_U242 = ~new_P1_U3062 | ~new_P1_R1117_U51;
  assign new_P1_R1117_U243 = ~new_P1_R1117_U189 | ~new_P1_R1117_U8;
  assign new_P1_R1117_U244 = ~new_P1_R1117_U9 | ~new_P1_R1117_U243;
  assign new_P1_R1117_U245 = ~new_P1_U3491 | ~new_P1_R1117_U52;
  assign new_P1_R1117_U246 = ~new_P1_R1117_U125 | ~new_P1_R1117_U148;
  assign new_P1_R1117_U247 = ~new_P1_R1117_U245 | ~new_P1_R1117_U244;
  assign new_P1_R1117_U248 = ~new_P1_R1117_U173;
  assign new_P1_R1117_U249 = ~new_P1_U3494 | ~new_P1_R1117_U56;
  assign new_P1_R1117_U250 = ~new_P1_R1117_U249 | ~new_P1_R1117_U173;
  assign new_P1_R1117_U251 = ~new_P1_U3072 | ~new_P1_R1117_U55;
  assign new_P1_R1117_U252 = ~new_P1_R1117_U172;
  assign new_P1_R1117_U253 = ~new_P1_U3497 | ~new_P1_R1117_U58;
  assign new_P1_R1117_U254 = ~new_P1_R1117_U253 | ~new_P1_R1117_U172;
  assign new_P1_R1117_U255 = ~new_P1_U3080 | ~new_P1_R1117_U57;
  assign new_P1_R1117_U256 = ~new_P1_R1117_U171;
  assign new_P1_R1117_U257 = ~new_P1_U3506 | ~new_P1_R1117_U61;
  assign new_P1_R1117_U258 = ~new_P1_U3073 | ~new_P1_R1117_U59;
  assign new_P1_R1117_U259 = ~new_P1_U3074 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U260 = ~new_P1_R1117_U186 | ~new_P1_R1117_U180;
  assign new_P1_R1117_U261 = ~new_P1_R1117_U10 | ~new_P1_R1117_U260;
  assign new_P1_R1117_U262 = ~new_P1_U3500 | ~new_P1_R1117_U63;
  assign new_P1_R1117_U263 = ~new_P1_U3506 | ~new_P1_R1117_U61;
  assign new_P1_R1117_U264 = ~new_P1_R1117_U257 | ~new_P1_R1117_U171 | ~new_P1_R1117_U126;
  assign new_P1_R1117_U265 = ~new_P1_R1117_U263 | ~new_P1_R1117_U261;
  assign new_P1_R1117_U266 = ~new_P1_R1117_U168;
  assign new_P1_R1117_U267 = ~new_P1_U3509 | ~new_P1_R1117_U66;
  assign new_P1_R1117_U268 = ~new_P1_R1117_U267 | ~new_P1_R1117_U168;
  assign new_P1_R1117_U269 = ~new_P1_U3069 | ~new_P1_R1117_U65;
  assign new_P1_R1117_U270 = ~new_P1_R1117_U67;
  assign new_P1_R1117_U271 = ~new_P1_R1117_U270 | ~new_P1_R1117_U68;
  assign new_P1_R1117_U272 = ~new_P1_R1117_U271 | ~new_P1_R1117_U167;
  assign new_P1_R1117_U273 = ~new_P1_U3082 | ~new_P1_R1117_U67;
  assign new_P1_R1117_U274 = ~new_P1_R1117_U166;
  assign new_P1_R1117_U275 = ~new_P1_U3514 | ~new_P1_R1117_U70;
  assign new_P1_R1117_U276 = ~new_P1_R1117_U275 | ~new_P1_R1117_U166;
  assign new_P1_R1117_U277 = ~new_P1_U3081 | ~new_P1_R1117_U69;
  assign new_P1_R1117_U278 = ~new_P1_R1117_U164;
  assign new_P1_R1117_U279 = ~new_P1_U4025 | ~new_P1_R1117_U72;
  assign new_P1_R1117_U280 = ~new_P1_R1117_U279 | ~new_P1_R1117_U164;
  assign new_P1_R1117_U281 = ~new_P1_U3076 | ~new_P1_R1117_U71;
  assign new_P1_R1117_U282 = ~new_P1_R1117_U163;
  assign new_P1_R1117_U283 = ~new_P1_U4022 | ~new_P1_R1117_U75;
  assign new_P1_R1117_U284 = ~new_P1_U3066 | ~new_P1_R1117_U73;
  assign new_P1_R1117_U285 = ~new_P1_U3061 | ~new_P1_R1117_U48;
  assign new_P1_R1117_U286 = ~new_P1_R1117_U187 | ~new_P1_R1117_U181;
  assign new_P1_R1117_U287 = ~new_P1_R1117_U11 | ~new_P1_R1117_U286;
  assign new_P1_R1117_U288 = ~new_P1_U4024 | ~new_P1_R1117_U77;
  assign new_P1_R1117_U289 = ~new_P1_U4022 | ~new_P1_R1117_U75;
  assign new_P1_R1117_U290 = ~new_P1_R1117_U283 | ~new_P1_R1117_U163 | ~new_P1_R1117_U127;
  assign new_P1_R1117_U291 = ~new_P1_R1117_U289 | ~new_P1_R1117_U287;
  assign new_P1_R1117_U292 = ~new_P1_R1117_U160;
  assign new_P1_R1117_U293 = ~new_P1_U4021 | ~new_P1_R1117_U80;
  assign new_P1_R1117_U294 = ~new_P1_R1117_U293 | ~new_P1_R1117_U160;
  assign new_P1_R1117_U295 = ~new_P1_U3065 | ~new_P1_R1117_U79;
  assign new_P1_R1117_U296 = ~new_P1_R1117_U159;
  assign new_P1_R1117_U297 = ~new_P1_U4020 | ~new_P1_R1117_U82;
  assign new_P1_R1117_U298 = ~new_P1_R1117_U297 | ~new_P1_R1117_U159;
  assign new_P1_R1117_U299 = ~new_P1_U3058 | ~new_P1_R1117_U81;
  assign new_P1_R1117_U300 = ~new_P1_R1117_U89;
  assign new_P1_R1117_U301 = ~new_P1_U4018 | ~new_P1_R1117_U86;
  assign new_P1_R1117_U302 = ~new_P1_R1117_U301 | ~new_P1_R1117_U89 | ~new_P1_R1117_U182;
  assign new_P1_R1117_U303 = ~new_P1_R1117_U86 | ~new_P1_R1117_U85;
  assign new_P1_R1117_U304 = ~new_P1_R1117_U303 | ~new_P1_R1117_U83;
  assign new_P1_R1117_U305 = ~new_P1_U3053 | ~new_P1_R1117_U176;
  assign new_P1_R1117_U306 = ~new_P1_R1117_U157;
  assign new_P1_R1117_U307 = ~new_P1_U4017 | ~new_P1_R1117_U88;
  assign new_P1_R1117_U308 = ~new_P1_U3054 | ~new_P1_R1117_U87;
  assign new_P1_R1117_U309 = ~new_P1_R1117_U300 | ~new_P1_R1117_U85;
  assign new_P1_R1117_U310 = ~new_P1_R1117_U133 | ~new_P1_R1117_U309;
  assign new_P1_R1117_U311 = ~new_P1_R1117_U89 | ~new_P1_R1117_U182;
  assign new_P1_R1117_U312 = ~new_P1_R1117_U132 | ~new_P1_R1117_U311;
  assign new_P1_R1117_U313 = ~new_P1_R1117_U85 | ~new_P1_R1117_U182;
  assign new_P1_R1117_U314 = ~new_P1_R1117_U288 | ~new_P1_R1117_U163;
  assign new_P1_R1117_U315 = ~new_P1_R1117_U90;
  assign new_P1_R1117_U316 = ~new_P1_U3061 | ~new_P1_R1117_U48;
  assign new_P1_R1117_U317 = ~new_P1_R1117_U315 | ~new_P1_R1117_U316;
  assign new_P1_R1117_U318 = ~new_P1_R1117_U136 | ~new_P1_R1117_U317;
  assign new_P1_R1117_U319 = ~new_P1_R1117_U90 | ~new_P1_R1117_U181;
  assign new_P1_R1117_U320 = ~new_P1_U4022 | ~new_P1_R1117_U75;
  assign new_P1_R1117_U321 = ~new_P1_R1117_U11 | ~new_P1_R1117_U320 | ~new_P1_R1117_U319;
  assign new_P1_R1117_U322 = ~new_P1_U3061 | ~new_P1_R1117_U48;
  assign new_P1_R1117_U323 = ~new_P1_R1117_U181 | ~new_P1_R1117_U322;
  assign new_P1_R1117_U324 = ~new_P1_R1117_U288 | ~new_P1_R1117_U78;
  assign new_P1_R1117_U325 = ~new_P1_R1117_U262 | ~new_P1_R1117_U171;
  assign new_P1_R1117_U326 = ~new_P1_R1117_U91;
  assign new_P1_R1117_U327 = ~new_P1_U3074 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U328 = ~new_P1_R1117_U326 | ~new_P1_R1117_U327;
  assign new_P1_R1117_U329 = ~new_P1_R1117_U142 | ~new_P1_R1117_U328;
  assign new_P1_R1117_U330 = ~new_P1_R1117_U91 | ~new_P1_R1117_U180;
  assign new_P1_R1117_U331 = ~new_P1_U3506 | ~new_P1_R1117_U61;
  assign new_P1_R1117_U332 = ~new_P1_R1117_U10 | ~new_P1_R1117_U331 | ~new_P1_R1117_U330;
  assign new_P1_R1117_U333 = ~new_P1_U3074 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U334 = ~new_P1_R1117_U180 | ~new_P1_R1117_U333;
  assign new_P1_R1117_U335 = ~new_P1_R1117_U262 | ~new_P1_R1117_U64;
  assign new_P1_R1117_U336 = ~new_P1_R1117_U217 | ~new_P1_R1117_U148;
  assign new_P1_R1117_U337 = ~new_P1_R1117_U92;
  assign new_P1_R1117_U338 = ~new_P1_U3062 | ~new_P1_R1117_U51;
  assign new_P1_R1117_U339 = ~new_P1_R1117_U337 | ~new_P1_R1117_U338;
  assign new_P1_R1117_U340 = ~new_P1_R1117_U146 | ~new_P1_R1117_U339;
  assign new_P1_R1117_U341 = ~new_P1_R1117_U92 | ~new_P1_R1117_U179;
  assign new_P1_R1117_U342 = ~new_P1_U3491 | ~new_P1_R1117_U52;
  assign new_P1_R1117_U343 = ~new_P1_R1117_U145 | ~new_P1_R1117_U341;
  assign new_P1_R1117_U344 = ~new_P1_U3062 | ~new_P1_R1117_U51;
  assign new_P1_R1117_U345 = ~new_P1_R1117_U179 | ~new_P1_R1117_U344;
  assign new_P1_R1117_U346 = ~new_P1_U3077 | ~new_P1_R1117_U24;
  assign new_P1_R1117_U347 = ~new_P1_R1117_U301 | ~new_P1_R1117_U89 | ~new_P1_R1117_U182;
  assign new_P1_R1117_U348 = ~new_P1_R1117_U130 | ~new_P1_R1117_U12 | ~new_P1_R1117_U347;
  assign new_P1_R1117_U349 = ~new_P1_U3485 | ~new_P1_R1117_U43;
  assign new_P1_R1117_U350 = ~new_P1_U3083 | ~new_P1_R1117_U42;
  assign new_P1_R1117_U351 = ~new_P1_R1117_U218 | ~new_P1_R1117_U148;
  assign new_P1_R1117_U352 = ~new_P1_R1117_U216 | ~new_P1_R1117_U147;
  assign new_P1_R1117_U353 = ~new_P1_U3482 | ~new_P1_R1117_U41;
  assign new_P1_R1117_U354 = ~new_P1_U3084 | ~new_P1_R1117_U38;
  assign new_P1_R1117_U355 = ~new_P1_U3482 | ~new_P1_R1117_U41;
  assign new_P1_R1117_U356 = ~new_P1_U3084 | ~new_P1_R1117_U38;
  assign new_P1_R1117_U357 = ~new_P1_R1117_U356 | ~new_P1_R1117_U355;
  assign new_P1_R1117_U358 = ~new_P1_U3479 | ~new_P1_R1117_U39;
  assign new_P1_R1117_U359 = ~new_P1_U3070 | ~new_P1_R1117_U22;
  assign new_P1_R1117_U360 = ~new_P1_R1117_U223 | ~new_P1_R1117_U44;
  assign new_P1_R1117_U361 = ~new_P1_R1117_U149 | ~new_P1_R1117_U210;
  assign new_P1_R1117_U362 = ~new_P1_U3476 | ~new_P1_R1117_U34;
  assign new_P1_R1117_U363 = ~new_P1_U3071 | ~new_P1_R1117_U31;
  assign new_P1_R1117_U364 = ~new_P1_R1117_U363 | ~new_P1_R1117_U362;
  assign new_P1_R1117_U365 = ~new_P1_U3473 | ~new_P1_R1117_U35;
  assign new_P1_R1117_U366 = ~new_P1_U3067 | ~new_P1_R1117_U32;
  assign new_P1_R1117_U367 = ~new_P1_R1117_U233 | ~new_P1_R1117_U45;
  assign new_P1_R1117_U368 = ~new_P1_R1117_U150 | ~new_P1_R1117_U225;
  assign new_P1_R1117_U369 = ~new_P1_U3470 | ~new_P1_R1117_U36;
  assign new_P1_R1117_U370 = ~new_P1_U3060 | ~new_P1_R1117_U33;
  assign new_P1_R1117_U371 = ~new_P1_R1117_U234 | ~new_P1_R1117_U152;
  assign new_P1_R1117_U372 = ~new_P1_R1117_U200 | ~new_P1_R1117_U151;
  assign new_P1_R1117_U373 = ~new_P1_U3467 | ~new_P1_R1117_U30;
  assign new_P1_R1117_U374 = ~new_P1_U3064 | ~new_P1_R1117_U27;
  assign new_P1_R1117_U375 = ~new_P1_U3467 | ~new_P1_R1117_U30;
  assign new_P1_R1117_U376 = ~new_P1_U3064 | ~new_P1_R1117_U27;
  assign new_P1_R1117_U377 = ~new_P1_R1117_U376 | ~new_P1_R1117_U375;
  assign new_P1_R1117_U378 = ~new_P1_U3464 | ~new_P1_R1117_U28;
  assign new_P1_R1117_U379 = ~new_P1_U3068 | ~new_P1_R1117_U23;
  assign new_P1_R1117_U380 = ~new_P1_R1117_U239 | ~new_P1_R1117_U46;
  assign new_P1_R1117_U381 = ~new_P1_R1117_U153 | ~new_P1_R1117_U194;
  assign new_P1_R1117_U382 = ~new_P1_U4028 | ~new_P1_R1117_U155;
  assign new_P1_R1117_U383 = ~new_P1_U3055 | ~new_P1_R1117_U154;
  assign new_P1_R1117_U384 = ~new_P1_U4028 | ~new_P1_R1117_U155;
  assign new_P1_R1117_U385 = ~new_P1_U3055 | ~new_P1_R1117_U154;
  assign new_P1_R1117_U386 = ~new_P1_R1117_U385 | ~new_P1_R1117_U384;
  assign new_P1_R1117_U387 = ~new_P1_R1117_U87 | ~new_P1_U3054 | ~new_P1_R1117_U386;
  assign new_P1_R1117_U388 = ~new_P1_U4017 | ~new_P1_R1117_U12 | ~new_P1_R1117_U88;
  assign new_P1_R1117_U389 = ~new_P1_U4017 | ~new_P1_R1117_U88;
  assign new_P1_R1117_U390 = ~new_P1_U3054 | ~new_P1_R1117_U87;
  assign new_P1_R1117_U391 = ~new_P1_R1117_U131;
  assign new_P1_R1117_U392 = ~new_P1_R1117_U306 | ~new_P1_R1117_U391;
  assign new_P1_R1117_U393 = ~new_P1_R1117_U131 | ~new_P1_R1117_U157;
  assign new_P1_R1117_U394 = ~new_P1_U4018 | ~new_P1_R1117_U86;
  assign new_P1_R1117_U395 = ~new_P1_U3053 | ~new_P1_R1117_U83;
  assign new_P1_R1117_U396 = ~new_P1_U4018 | ~new_P1_R1117_U86;
  assign new_P1_R1117_U397 = ~new_P1_U3053 | ~new_P1_R1117_U83;
  assign new_P1_R1117_U398 = ~new_P1_R1117_U397 | ~new_P1_R1117_U396;
  assign new_P1_R1117_U399 = ~new_P1_U4019 | ~new_P1_R1117_U84;
  assign new_P1_R1117_U400 = ~new_P1_U3057 | ~new_P1_R1117_U47;
  assign new_P1_R1117_U401 = ~new_P1_R1117_U313 | ~new_P1_R1117_U89;
  assign new_P1_R1117_U402 = ~new_P1_R1117_U158 | ~new_P1_R1117_U300;
  assign new_P1_R1117_U403 = ~new_P1_U4020 | ~new_P1_R1117_U82;
  assign new_P1_R1117_U404 = ~new_P1_U3058 | ~new_P1_R1117_U81;
  assign new_P1_R1117_U405 = ~new_P1_R1117_U134;
  assign new_P1_R1117_U406 = ~new_P1_R1117_U296 | ~new_P1_R1117_U405;
  assign new_P1_R1117_U407 = ~new_P1_R1117_U134 | ~new_P1_R1117_U159;
  assign new_P1_R1117_U408 = ~new_P1_U4021 | ~new_P1_R1117_U80;
  assign new_P1_R1117_U409 = ~new_P1_U3065 | ~new_P1_R1117_U79;
  assign new_P1_R1117_U410 = ~new_P1_R1117_U135;
  assign new_P1_R1117_U411 = ~new_P1_R1117_U292 | ~new_P1_R1117_U410;
  assign new_P1_R1117_U412 = ~new_P1_R1117_U135 | ~new_P1_R1117_U160;
  assign new_P1_R1117_U413 = ~new_P1_U4022 | ~new_P1_R1117_U75;
  assign new_P1_R1117_U414 = ~new_P1_U3066 | ~new_P1_R1117_U73;
  assign new_P1_R1117_U415 = ~new_P1_R1117_U414 | ~new_P1_R1117_U413;
  assign new_P1_R1117_U416 = ~new_P1_U4023 | ~new_P1_R1117_U76;
  assign new_P1_R1117_U417 = ~new_P1_U3061 | ~new_P1_R1117_U48;
  assign new_P1_R1117_U418 = ~new_P1_R1117_U323 | ~new_P1_R1117_U90;
  assign new_P1_R1117_U419 = ~new_P1_R1117_U161 | ~new_P1_R1117_U315;
  assign new_P1_R1117_U420 = ~new_P1_U4024 | ~new_P1_R1117_U77;
  assign new_P1_R1117_U421 = ~new_P1_U3075 | ~new_P1_R1117_U74;
  assign new_P1_R1117_U422 = ~new_P1_R1117_U324 | ~new_P1_R1117_U163;
  assign new_P1_R1117_U423 = ~new_P1_R1117_U282 | ~new_P1_R1117_U162;
  assign new_P1_R1117_U424 = ~new_P1_U4025 | ~new_P1_R1117_U72;
  assign new_P1_R1117_U425 = ~new_P1_U3076 | ~new_P1_R1117_U71;
  assign new_P1_R1117_U426 = ~new_P1_R1117_U137;
  assign new_P1_R1117_U427 = ~new_P1_R1117_U278 | ~new_P1_R1117_U426;
  assign new_P1_R1117_U428 = ~new_P1_R1117_U137 | ~new_P1_R1117_U164;
  assign new_P1_R1117_U429 = ~new_P1_U3461 | ~new_P1_R1117_U26;
  assign new_P1_R1117_U430 = ~new_P1_U3078 | ~new_P1_R1117_U165;
  assign new_P1_R1117_U431 = ~new_P1_R1117_U138;
  assign new_P1_R1117_U432 = ~new_P1_R1117_U431 | ~new_P1_R1117_U190;
  assign new_P1_R1117_U433 = ~new_P1_R1117_U138 | ~new_P1_R1117_U25;
  assign new_P1_R1117_U434 = ~new_P1_U3514 | ~new_P1_R1117_U70;
  assign new_P1_R1117_U435 = ~new_P1_U3081 | ~new_P1_R1117_U69;
  assign new_P1_R1117_U436 = ~new_P1_R1117_U139;
  assign new_P1_R1117_U437 = ~new_P1_R1117_U274 | ~new_P1_R1117_U436;
  assign new_P1_R1117_U438 = ~new_P1_R1117_U139 | ~new_P1_R1117_U166;
  assign new_P1_R1117_U439 = ~new_P1_U3512 | ~new_P1_R1117_U68;
  assign new_P1_R1117_U440 = ~new_P1_U3082 | ~new_P1_R1117_U167;
  assign new_P1_R1117_U441 = ~new_P1_R1117_U140;
  assign new_P1_R1117_U442 = ~new_P1_R1117_U441 | ~new_P1_R1117_U270;
  assign new_P1_R1117_U443 = ~new_P1_R1117_U140 | ~new_P1_R1117_U67;
  assign new_P1_R1117_U444 = ~new_P1_U3509 | ~new_P1_R1117_U66;
  assign new_P1_R1117_U445 = ~new_P1_U3069 | ~new_P1_R1117_U65;
  assign new_P1_R1117_U446 = ~new_P1_R1117_U141;
  assign new_P1_R1117_U447 = ~new_P1_R1117_U266 | ~new_P1_R1117_U446;
  assign new_P1_R1117_U448 = ~new_P1_R1117_U141 | ~new_P1_R1117_U168;
  assign new_P1_R1117_U449 = ~new_P1_U3506 | ~new_P1_R1117_U61;
  assign new_P1_R1117_U450 = ~new_P1_U3073 | ~new_P1_R1117_U59;
  assign new_P1_R1117_U451 = ~new_P1_R1117_U450 | ~new_P1_R1117_U449;
  assign new_P1_R1117_U452 = ~new_P1_U3503 | ~new_P1_R1117_U62;
  assign new_P1_R1117_U453 = ~new_P1_U3074 | ~new_P1_R1117_U49;
  assign new_P1_R1117_U454 = ~new_P1_R1117_U334 | ~new_P1_R1117_U91;
  assign new_P1_R1117_U455 = ~new_P1_R1117_U169 | ~new_P1_R1117_U326;
  assign new_P1_R1117_U456 = ~new_P1_U3500 | ~new_P1_R1117_U63;
  assign new_P1_R1117_U457 = ~new_P1_U3079 | ~new_P1_R1117_U60;
  assign new_P1_R1117_U458 = ~new_P1_R1117_U335 | ~new_P1_R1117_U171;
  assign new_P1_R1117_U459 = ~new_P1_R1117_U256 | ~new_P1_R1117_U170;
  assign new_P1_R1117_U460 = ~new_P1_U3497 | ~new_P1_R1117_U58;
  assign new_P1_R1117_U461 = ~new_P1_U3080 | ~new_P1_R1117_U57;
  assign new_P1_R1117_U462 = ~new_P1_R1117_U143;
  assign new_P1_R1117_U463 = ~new_P1_R1117_U252 | ~new_P1_R1117_U462;
  assign new_P1_R1117_U464 = ~new_P1_R1117_U143 | ~new_P1_R1117_U172;
  assign new_P1_R1117_U465 = ~new_P1_U3494 | ~new_P1_R1117_U56;
  assign new_P1_R1117_U466 = ~new_P1_U3072 | ~new_P1_R1117_U55;
  assign new_P1_R1117_U467 = ~new_P1_R1117_U144;
  assign new_P1_R1117_U468 = ~new_P1_R1117_U248 | ~new_P1_R1117_U467;
  assign new_P1_R1117_U469 = ~new_P1_R1117_U144 | ~new_P1_R1117_U173;
  assign new_P1_R1117_U470 = ~new_P1_U3491 | ~new_P1_R1117_U52;
  assign new_P1_R1117_U471 = ~new_P1_U3063 | ~new_P1_R1117_U50;
  assign new_P1_R1117_U472 = ~new_P1_R1117_U471 | ~new_P1_R1117_U470;
  assign new_P1_R1117_U473 = ~new_P1_U3488 | ~new_P1_R1117_U53;
  assign new_P1_R1117_U474 = ~new_P1_U3062 | ~new_P1_R1117_U51;
  assign new_P1_R1117_U475 = ~new_P1_R1117_U345 | ~new_P1_R1117_U92;
  assign new_P1_R1117_U476 = ~new_P1_R1117_U174 | ~new_P1_R1117_U337;
  assign new_P1_R1375_U6 = new_P1_R1375_U8 & new_P1_R1375_U191;
  assign new_P1_R1375_U7 = new_P1_R1375_U189 & new_P1_R1375_U190 & new_P1_R1375_U100;
  assign new_P1_R1375_U8 = new_P1_R1375_U195 & new_P1_R1375_U194;
  assign new_P1_R1375_U9 = ~new_P1_R1375_U7 | ~new_P1_R1375_U192;
  assign new_P1_R1375_U10 = ~new_P1_U3088;
  assign new_P1_R1375_U11 = ~new_P1_U3087;
  assign new_P1_R1375_U12 = ~new_P1_U3121;
  assign new_P1_R1375_U13 = ~new_P1_U3120;
  assign new_P1_R1375_U14 = ~new_P1_U3152;
  assign new_P1_R1375_U15 = ~new_P1_U3117;
  assign new_P1_R1375_U16 = ~new_P1_U3149;
  assign new_P1_R1375_U17 = ~new_P1_U3148;
  assign new_P1_R1375_U18 = ~new_P1_U3116;
  assign new_P1_R1375_U19 = ~new_P1_U3115;
  assign new_P1_R1375_U20 = ~new_P1_U3147;
  assign new_P1_R1375_U21 = ~new_P1_U3146;
  assign new_P1_R1375_U22 = ~new_P1_U3114;
  assign new_P1_R1375_U23 = ~new_P1_U3113;
  assign new_P1_R1375_U24 = ~new_P1_U3145;
  assign new_P1_R1375_U25 = ~new_P1_U3144;
  assign new_P1_R1375_U26 = ~new_P1_U3112;
  assign new_P1_R1375_U27 = ~new_P1_U3111;
  assign new_P1_R1375_U28 = ~new_P1_U3143;
  assign new_P1_R1375_U29 = ~new_P1_U3142;
  assign new_P1_R1375_U30 = ~new_P1_U3110;
  assign new_P1_R1375_U31 = ~new_P1_U3109;
  assign new_P1_R1375_U32 = ~new_P1_U3141;
  assign new_P1_R1375_U33 = ~new_P1_U3140;
  assign new_P1_R1375_U34 = ~new_P1_U3108;
  assign new_P1_R1375_U35 = ~new_P1_U3107;
  assign new_P1_R1375_U36 = ~new_P1_U3139;
  assign new_P1_R1375_U37 = ~new_P1_U3138;
  assign new_P1_R1375_U38 = ~new_P1_U3106;
  assign new_P1_R1375_U39 = ~new_P1_U3105;
  assign new_P1_R1375_U40 = ~new_P1_U3137;
  assign new_P1_R1375_U41 = ~new_P1_U3136;
  assign new_P1_R1375_U42 = ~new_P1_U3104;
  assign new_P1_R1375_U43 = ~new_P1_U3103;
  assign new_P1_R1375_U44 = ~new_P1_U3135;
  assign new_P1_R1375_U45 = ~new_P1_U3134;
  assign new_P1_R1375_U46 = ~new_P1_U3102;
  assign new_P1_R1375_U47 = ~new_P1_U3101;
  assign new_P1_R1375_U48 = ~new_P1_U3133;
  assign new_P1_R1375_U49 = ~new_P1_U3132;
  assign new_P1_R1375_U50 = ~new_P1_U3100;
  assign new_P1_R1375_U51 = ~new_P1_U3099;
  assign new_P1_R1375_U52 = ~new_P1_U3131;
  assign new_P1_R1375_U53 = ~new_P1_U3130;
  assign new_P1_R1375_U54 = ~new_P1_U3098;
  assign new_P1_R1375_U55 = ~new_P1_U3097;
  assign new_P1_R1375_U56 = ~new_P1_U3129;
  assign new_P1_R1375_U57 = ~new_P1_U3128;
  assign new_P1_R1375_U58 = ~new_P1_U3096;
  assign new_P1_R1375_U59 = ~new_P1_U3095;
  assign new_P1_R1375_U60 = ~new_P1_U3127;
  assign new_P1_R1375_U61 = ~new_P1_U3126;
  assign new_P1_R1375_U62 = ~new_P1_U3094;
  assign new_P1_R1375_U63 = ~new_P1_U3093;
  assign new_P1_R1375_U64 = ~new_P1_U3125;
  assign new_P1_R1375_U65 = ~new_P1_U3124;
  assign new_P1_R1375_U66 = ~new_P1_U3092;
  assign new_P1_R1375_U67 = ~new_P1_U3091;
  assign new_P1_R1375_U68 = ~new_P1_U3123;
  assign new_P1_R1375_U69 = ~new_P1_U3089;
  assign new_P1_R1375_U70 = new_P1_R1375_U107 & new_P1_R1375_U108;
  assign new_P1_R1375_U71 = new_P1_R1375_U110 & new_P1_R1375_U111;
  assign new_P1_R1375_U72 = new_P1_R1375_U113 & new_P1_R1375_U114;
  assign new_P1_R1375_U73 = new_P1_R1375_U116 & new_P1_R1375_U117;
  assign new_P1_R1375_U74 = new_P1_R1375_U119 & new_P1_R1375_U120;
  assign new_P1_R1375_U75 = new_P1_R1375_U122 & new_P1_R1375_U123;
  assign new_P1_R1375_U76 = new_P1_R1375_U125 & new_P1_R1375_U126;
  assign new_P1_R1375_U77 = new_P1_R1375_U128 & new_P1_R1375_U129;
  assign new_P1_R1375_U78 = new_P1_R1375_U131 & new_P1_R1375_U132;
  assign new_P1_R1375_U79 = new_P1_R1375_U134 & new_P1_R1375_U135;
  assign new_P1_R1375_U80 = new_P1_R1375_U137 & new_P1_R1375_U138;
  assign new_P1_R1375_U81 = new_P1_R1375_U140 & new_P1_R1375_U141;
  assign new_P1_R1375_U82 = new_P1_R1375_U143 & new_P1_R1375_U144;
  assign new_P1_R1375_U83 = new_P1_R1375_U146 & new_P1_R1375_U147;
  assign new_P1_R1375_U84 = new_P1_R1375_U149 & new_P1_R1375_U150;
  assign new_P1_R1375_U85 = new_P1_R1375_U152 & new_P1_R1375_U153;
  assign new_P1_R1375_U86 = new_P1_R1375_U155 & new_P1_R1375_U156;
  assign new_P1_R1375_U87 = new_P1_R1375_U158 & new_P1_R1375_U159;
  assign new_P1_R1375_U88 = new_P1_R1375_U161 & new_P1_R1375_U162;
  assign new_P1_R1375_U89 = new_P1_R1375_U164 & new_P1_R1375_U165;
  assign new_P1_R1375_U90 = new_P1_R1375_U167 & new_P1_R1375_U168;
  assign new_P1_R1375_U91 = new_P1_R1375_U170 & new_P1_R1375_U171;
  assign new_P1_R1375_U92 = new_P1_R1375_U173 & new_P1_R1375_U174;
  assign new_P1_R1375_U93 = new_P1_R1375_U176 & new_P1_R1375_U177;
  assign new_P1_R1375_U94 = new_P1_R1375_U179 & new_P1_R1375_U180;
  assign new_P1_R1375_U95 = new_P1_R1375_U182 & new_P1_R1375_U183;
  assign new_P1_R1375_U96 = new_P1_R1375_U186 & new_P1_R1375_U101;
  assign new_P1_R1375_U97 = new_P1_R1375_U186 & new_P1_U3090;
  assign new_P1_R1375_U98 = new_P1_R1375_U187 & new_P1_R1375_U188;
  assign new_P1_R1375_U99 = ~new_P1_U3119;
  assign new_P1_R1375_U100 = new_P1_R1375_U197 & new_P1_R1375_U196;
  assign new_P1_R1375_U101 = ~new_P1_U3122;
  assign new_P1_R1375_U102 = ~new_P1_U3150 | ~new_P1_U3151;
  assign new_P1_R1375_U103 = ~new_P1_U3118 | ~new_P1_R1375_U102;
  assign new_P1_R1375_U104 = new_P1_U3150 | new_P1_U3151;
  assign new_P1_R1375_U105 = ~new_P1_U3117 | ~new_P1_R1375_U16;
  assign new_P1_R1375_U106 = ~new_P1_R1375_U103 | ~new_P1_R1375_U104 | ~new_P1_R1375_U105;
  assign new_P1_R1375_U107 = ~new_P1_U3149 | ~new_P1_R1375_U15;
  assign new_P1_R1375_U108 = ~new_P1_U3148 | ~new_P1_R1375_U18;
  assign new_P1_R1375_U109 = ~new_P1_R1375_U70 | ~new_P1_R1375_U106;
  assign new_P1_R1375_U110 = ~new_P1_U3116 | ~new_P1_R1375_U17;
  assign new_P1_R1375_U111 = ~new_P1_U3115 | ~new_P1_R1375_U20;
  assign new_P1_R1375_U112 = ~new_P1_R1375_U71 | ~new_P1_R1375_U109;
  assign new_P1_R1375_U113 = ~new_P1_U3147 | ~new_P1_R1375_U19;
  assign new_P1_R1375_U114 = ~new_P1_U3146 | ~new_P1_R1375_U22;
  assign new_P1_R1375_U115 = ~new_P1_R1375_U72 | ~new_P1_R1375_U112;
  assign new_P1_R1375_U116 = ~new_P1_U3114 | ~new_P1_R1375_U21;
  assign new_P1_R1375_U117 = ~new_P1_U3113 | ~new_P1_R1375_U24;
  assign new_P1_R1375_U118 = ~new_P1_R1375_U73 | ~new_P1_R1375_U115;
  assign new_P1_R1375_U119 = ~new_P1_U3145 | ~new_P1_R1375_U23;
  assign new_P1_R1375_U120 = ~new_P1_U3144 | ~new_P1_R1375_U26;
  assign new_P1_R1375_U121 = ~new_P1_R1375_U74 | ~new_P1_R1375_U118;
  assign new_P1_R1375_U122 = ~new_P1_U3112 | ~new_P1_R1375_U25;
  assign new_P1_R1375_U123 = ~new_P1_U3111 | ~new_P1_R1375_U28;
  assign new_P1_R1375_U124 = ~new_P1_R1375_U75 | ~new_P1_R1375_U121;
  assign new_P1_R1375_U125 = ~new_P1_U3143 | ~new_P1_R1375_U27;
  assign new_P1_R1375_U126 = ~new_P1_U3142 | ~new_P1_R1375_U30;
  assign new_P1_R1375_U127 = ~new_P1_R1375_U76 | ~new_P1_R1375_U124;
  assign new_P1_R1375_U128 = ~new_P1_U3110 | ~new_P1_R1375_U29;
  assign new_P1_R1375_U129 = ~new_P1_U3109 | ~new_P1_R1375_U32;
  assign new_P1_R1375_U130 = ~new_P1_R1375_U77 | ~new_P1_R1375_U127;
  assign new_P1_R1375_U131 = ~new_P1_U3141 | ~new_P1_R1375_U31;
  assign new_P1_R1375_U132 = ~new_P1_U3140 | ~new_P1_R1375_U34;
  assign new_P1_R1375_U133 = ~new_P1_R1375_U78 | ~new_P1_R1375_U130;
  assign new_P1_R1375_U134 = ~new_P1_U3108 | ~new_P1_R1375_U33;
  assign new_P1_R1375_U135 = ~new_P1_U3107 | ~new_P1_R1375_U36;
  assign new_P1_R1375_U136 = ~new_P1_R1375_U79 | ~new_P1_R1375_U133;
  assign new_P1_R1375_U137 = ~new_P1_U3139 | ~new_P1_R1375_U35;
  assign new_P1_R1375_U138 = ~new_P1_U3138 | ~new_P1_R1375_U38;
  assign new_P1_R1375_U139 = ~new_P1_R1375_U80 | ~new_P1_R1375_U136;
  assign new_P1_R1375_U140 = ~new_P1_U3106 | ~new_P1_R1375_U37;
  assign new_P1_R1375_U141 = ~new_P1_U3105 | ~new_P1_R1375_U40;
  assign new_P1_R1375_U142 = ~new_P1_R1375_U81 | ~new_P1_R1375_U139;
  assign new_P1_R1375_U143 = ~new_P1_U3137 | ~new_P1_R1375_U39;
  assign new_P1_R1375_U144 = ~new_P1_U3136 | ~new_P1_R1375_U42;
  assign new_P1_R1375_U145 = ~new_P1_R1375_U82 | ~new_P1_R1375_U142;
  assign new_P1_R1375_U146 = ~new_P1_U3104 | ~new_P1_R1375_U41;
  assign new_P1_R1375_U147 = ~new_P1_U3103 | ~new_P1_R1375_U44;
  assign new_P1_R1375_U148 = ~new_P1_R1375_U83 | ~new_P1_R1375_U145;
  assign new_P1_R1375_U149 = ~new_P1_U3135 | ~new_P1_R1375_U43;
  assign new_P1_R1375_U150 = ~new_P1_U3134 | ~new_P1_R1375_U46;
  assign new_P1_R1375_U151 = ~new_P1_R1375_U84 | ~new_P1_R1375_U148;
  assign new_P1_R1375_U152 = ~new_P1_U3102 | ~new_P1_R1375_U45;
  assign new_P1_R1375_U153 = ~new_P1_U3101 | ~new_P1_R1375_U48;
  assign new_P1_R1375_U154 = ~new_P1_R1375_U85 | ~new_P1_R1375_U151;
  assign new_P1_R1375_U155 = ~new_P1_U3133 | ~new_P1_R1375_U47;
  assign new_P1_R1375_U156 = ~new_P1_U3132 | ~new_P1_R1375_U50;
  assign new_P1_R1375_U157 = ~new_P1_R1375_U86 | ~new_P1_R1375_U154;
  assign new_P1_R1375_U158 = ~new_P1_U3100 | ~new_P1_R1375_U49;
  assign new_P1_R1375_U159 = ~new_P1_U3099 | ~new_P1_R1375_U52;
  assign new_P1_R1375_U160 = ~new_P1_R1375_U87 | ~new_P1_R1375_U157;
  assign new_P1_R1375_U161 = ~new_P1_U3131 | ~new_P1_R1375_U51;
  assign new_P1_R1375_U162 = ~new_P1_U3130 | ~new_P1_R1375_U54;
  assign new_P1_R1375_U163 = ~new_P1_R1375_U88 | ~new_P1_R1375_U160;
  assign new_P1_R1375_U164 = ~new_P1_U3098 | ~new_P1_R1375_U53;
  assign new_P1_R1375_U165 = ~new_P1_U3097 | ~new_P1_R1375_U56;
  assign new_P1_R1375_U166 = ~new_P1_R1375_U89 | ~new_P1_R1375_U163;
  assign new_P1_R1375_U167 = ~new_P1_U3129 | ~new_P1_R1375_U55;
  assign new_P1_R1375_U168 = ~new_P1_U3128 | ~new_P1_R1375_U58;
  assign new_P1_R1375_U169 = ~new_P1_R1375_U90 | ~new_P1_R1375_U166;
  assign new_P1_R1375_U170 = ~new_P1_U3096 | ~new_P1_R1375_U57;
  assign new_P1_R1375_U171 = ~new_P1_U3095 | ~new_P1_R1375_U60;
  assign new_P1_R1375_U172 = ~new_P1_R1375_U91 | ~new_P1_R1375_U169;
  assign new_P1_R1375_U173 = ~new_P1_U3127 | ~new_P1_R1375_U59;
  assign new_P1_R1375_U174 = ~new_P1_U3126 | ~new_P1_R1375_U62;
  assign new_P1_R1375_U175 = ~new_P1_R1375_U92 | ~new_P1_R1375_U172;
  assign new_P1_R1375_U176 = ~new_P1_U3094 | ~new_P1_R1375_U61;
  assign new_P1_R1375_U177 = ~new_P1_U3093 | ~new_P1_R1375_U64;
  assign new_P1_R1375_U178 = ~new_P1_R1375_U93 | ~new_P1_R1375_U175;
  assign new_P1_R1375_U179 = ~new_P1_U3125 | ~new_P1_R1375_U63;
  assign new_P1_R1375_U180 = ~new_P1_U3124 | ~new_P1_R1375_U66;
  assign new_P1_R1375_U181 = ~new_P1_R1375_U94 | ~new_P1_R1375_U178;
  assign new_P1_R1375_U182 = ~new_P1_U3092 | ~new_P1_R1375_U65;
  assign new_P1_R1375_U183 = ~new_P1_U3091 | ~new_P1_R1375_U68;
  assign new_P1_R1375_U184 = ~new_P1_R1375_U95 | ~new_P1_R1375_U181;
  assign new_P1_R1375_U185 = ~new_P1_R1375_U96 | ~new_P1_R1375_U184;
  assign new_P1_R1375_U186 = ~new_P1_U3123 | ~new_P1_R1375_U67;
  assign new_P1_R1375_U187 = ~new_P1_U3090 | ~new_P1_R1375_U101;
  assign new_P1_R1375_U188 = ~new_P1_U3089 | ~new_P1_R1375_U12;
  assign new_P1_R1375_U189 = ~new_P1_R1375_U69 | ~new_P1_U3121 | ~new_P1_R1375_U8 | ~new_P1_R1375_U191;
  assign new_P1_R1375_U190 = ~new_P1_U3120 | ~new_P1_R1375_U8 | ~new_P1_R1375_U10;
  assign new_P1_R1375_U191 = ~new_P1_U3088 | ~new_P1_R1375_U13;
  assign new_P1_R1375_U192 = ~new_P1_R1375_U185 | ~new_P1_R1375_U98 | ~new_P1_R1375_U6 | ~new_P1_R1375_U193;
  assign new_P1_R1375_U193 = ~new_P1_R1375_U97 | ~new_P1_R1375_U184;
  assign new_P1_R1375_U194 = ~new_P1_U3087 | ~new_P1_R1375_U99;
  assign new_P1_R1375_U195 = ~new_P1_U3119 | ~new_P1_R1375_U11;
  assign new_P1_R1375_U196 = ~new_P1_R1375_U99 | ~new_P1_U3152 | ~new_P1_U3087;
  assign new_P1_R1375_U197 = ~new_P1_U3119 | ~new_P1_R1375_U14 | ~new_P1_R1375_U11;
  assign new_P1_R1352_U6 = new_P1_U3059 & new_P1_R1352_U7;
  assign new_P1_R1352_U7 = ~new_P1_U3056;
  assign new_P1_R1207_U6 = new_P1_R1207_U184 & new_P1_R1207_U201;
  assign new_P1_R1207_U7 = new_P1_R1207_U203 & new_P1_R1207_U202;
  assign new_P1_R1207_U8 = new_P1_R1207_U179 & new_P1_R1207_U240;
  assign new_P1_R1207_U9 = new_P1_R1207_U242 & new_P1_R1207_U241;
  assign new_P1_R1207_U10 = new_P1_R1207_U259 & new_P1_R1207_U258;
  assign new_P1_R1207_U11 = new_P1_R1207_U285 & new_P1_R1207_U284;
  assign new_P1_R1207_U12 = new_P1_R1207_U383 & new_P1_R1207_U382;
  assign new_P1_R1207_U13 = ~new_P1_R1207_U340 | ~new_P1_R1207_U343;
  assign new_P1_R1207_U14 = ~new_P1_R1207_U329 | ~new_P1_R1207_U332;
  assign new_P1_R1207_U15 = ~new_P1_R1207_U318 | ~new_P1_R1207_U321;
  assign new_P1_R1207_U16 = ~new_P1_R1207_U310 | ~new_P1_R1207_U312;
  assign new_P1_R1207_U17 = ~new_P1_R1207_U348 | ~new_P1_R1207_U156 | ~new_P1_R1207_U175;
  assign new_P1_R1207_U18 = ~new_P1_R1207_U236 | ~new_P1_R1207_U238;
  assign new_P1_R1207_U19 = ~new_P1_R1207_U228 | ~new_P1_R1207_U231;
  assign new_P1_R1207_U20 = ~new_P1_R1207_U220 | ~new_P1_R1207_U222;
  assign new_P1_R1207_U21 = ~new_P1_R1207_U25 | ~new_P1_R1207_U346;
  assign new_P1_R1207_U22 = ~new_P1_U3479;
  assign new_P1_R1207_U23 = ~new_P1_U3464;
  assign new_P1_R1207_U24 = ~new_P1_U3456;
  assign new_P1_R1207_U25 = ~new_P1_U3456 | ~new_P1_R1207_U93;
  assign new_P1_R1207_U26 = ~new_P1_U3078;
  assign new_P1_R1207_U27 = ~new_P1_U3467;
  assign new_P1_R1207_U28 = ~new_P1_U3068;
  assign new_P1_R1207_U29 = ~new_P1_U3068 | ~new_P1_R1207_U23;
  assign new_P1_R1207_U30 = ~new_P1_U3064;
  assign new_P1_R1207_U31 = ~new_P1_U3476;
  assign new_P1_R1207_U32 = ~new_P1_U3473;
  assign new_P1_R1207_U33 = ~new_P1_U3470;
  assign new_P1_R1207_U34 = ~new_P1_U3071;
  assign new_P1_R1207_U35 = ~new_P1_U3067;
  assign new_P1_R1207_U36 = ~new_P1_U3060;
  assign new_P1_R1207_U37 = ~new_P1_U3060 | ~new_P1_R1207_U33;
  assign new_P1_R1207_U38 = ~new_P1_U3482;
  assign new_P1_R1207_U39 = ~new_P1_U3070;
  assign new_P1_R1207_U40 = ~new_P1_U3070 | ~new_P1_R1207_U22;
  assign new_P1_R1207_U41 = ~new_P1_U3084;
  assign new_P1_R1207_U42 = ~new_P1_U3485;
  assign new_P1_R1207_U43 = ~new_P1_U3083;
  assign new_P1_R1207_U44 = ~new_P1_R1207_U209 | ~new_P1_R1207_U208;
  assign new_P1_R1207_U45 = ~new_P1_R1207_U37 | ~new_P1_R1207_U224;
  assign new_P1_R1207_U46 = ~new_P1_R1207_U193 | ~new_P1_R1207_U192;
  assign new_P1_R1207_U47 = ~new_P1_U4019;
  assign new_P1_R1207_U48 = ~new_P1_U4023;
  assign new_P1_R1207_U49 = ~new_P1_U3503;
  assign new_P1_R1207_U50 = ~new_P1_U3491;
  assign new_P1_R1207_U51 = ~new_P1_U3488;
  assign new_P1_R1207_U52 = ~new_P1_U3063;
  assign new_P1_R1207_U53 = ~new_P1_U3062;
  assign new_P1_R1207_U54 = ~new_P1_U3083 | ~new_P1_R1207_U42;
  assign new_P1_R1207_U55 = ~new_P1_U3494;
  assign new_P1_R1207_U56 = ~new_P1_U3072;
  assign new_P1_R1207_U57 = ~new_P1_U3497;
  assign new_P1_R1207_U58 = ~new_P1_U3080;
  assign new_P1_R1207_U59 = ~new_P1_U3506;
  assign new_P1_R1207_U60 = ~new_P1_U3500;
  assign new_P1_R1207_U61 = ~new_P1_U3073;
  assign new_P1_R1207_U62 = ~new_P1_U3074;
  assign new_P1_R1207_U63 = ~new_P1_U3079;
  assign new_P1_R1207_U64 = ~new_P1_U3079 | ~new_P1_R1207_U60;
  assign new_P1_R1207_U65 = ~new_P1_U3509;
  assign new_P1_R1207_U66 = ~new_P1_U3069;
  assign new_P1_R1207_U67 = ~new_P1_R1207_U269 | ~new_P1_R1207_U268;
  assign new_P1_R1207_U68 = ~new_P1_U3082;
  assign new_P1_R1207_U69 = ~new_P1_U3514;
  assign new_P1_R1207_U70 = ~new_P1_U3081;
  assign new_P1_R1207_U71 = ~new_P1_U4025;
  assign new_P1_R1207_U72 = ~new_P1_U3076;
  assign new_P1_R1207_U73 = ~new_P1_U4022;
  assign new_P1_R1207_U74 = ~new_P1_U4024;
  assign new_P1_R1207_U75 = ~new_P1_U3066;
  assign new_P1_R1207_U76 = ~new_P1_U3061;
  assign new_P1_R1207_U77 = ~new_P1_U3075;
  assign new_P1_R1207_U78 = ~new_P1_U3075 | ~new_P1_R1207_U74;
  assign new_P1_R1207_U79 = ~new_P1_U4021;
  assign new_P1_R1207_U80 = ~new_P1_U3065;
  assign new_P1_R1207_U81 = ~new_P1_U4020;
  assign new_P1_R1207_U82 = ~new_P1_U3058;
  assign new_P1_R1207_U83 = ~new_P1_U4018;
  assign new_P1_R1207_U84 = ~new_P1_U3057;
  assign new_P1_R1207_U85 = ~new_P1_U3057 | ~new_P1_R1207_U47;
  assign new_P1_R1207_U86 = ~new_P1_U3053;
  assign new_P1_R1207_U87 = ~new_P1_U4017;
  assign new_P1_R1207_U88 = ~new_P1_U3054;
  assign new_P1_R1207_U89 = ~new_P1_R1207_U299 | ~new_P1_R1207_U298;
  assign new_P1_R1207_U90 = ~new_P1_R1207_U78 | ~new_P1_R1207_U314;
  assign new_P1_R1207_U91 = ~new_P1_R1207_U64 | ~new_P1_R1207_U325;
  assign new_P1_R1207_U92 = ~new_P1_R1207_U54 | ~new_P1_R1207_U336;
  assign new_P1_R1207_U93 = ~new_P1_U3077;
  assign new_P1_R1207_U94 = ~new_P1_R1207_U393 | ~new_P1_R1207_U392;
  assign new_P1_R1207_U95 = ~new_P1_R1207_U407 | ~new_P1_R1207_U406;
  assign new_P1_R1207_U96 = ~new_P1_R1207_U412 | ~new_P1_R1207_U411;
  assign new_P1_R1207_U97 = ~new_P1_R1207_U428 | ~new_P1_R1207_U427;
  assign new_P1_R1207_U98 = ~new_P1_R1207_U433 | ~new_P1_R1207_U432;
  assign new_P1_R1207_U99 = ~new_P1_R1207_U438 | ~new_P1_R1207_U437;
  assign new_P1_R1207_U100 = ~new_P1_R1207_U443 | ~new_P1_R1207_U442;
  assign new_P1_R1207_U101 = ~new_P1_R1207_U448 | ~new_P1_R1207_U447;
  assign new_P1_R1207_U102 = ~new_P1_R1207_U464 | ~new_P1_R1207_U463;
  assign new_P1_R1207_U103 = ~new_P1_R1207_U469 | ~new_P1_R1207_U468;
  assign new_P1_R1207_U104 = ~new_P1_R1207_U352 | ~new_P1_R1207_U351;
  assign new_P1_R1207_U105 = ~new_P1_R1207_U361 | ~new_P1_R1207_U360;
  assign new_P1_R1207_U106 = ~new_P1_R1207_U368 | ~new_P1_R1207_U367;
  assign new_P1_R1207_U107 = ~new_P1_R1207_U372 | ~new_P1_R1207_U371;
  assign new_P1_R1207_U108 = ~new_P1_R1207_U381 | ~new_P1_R1207_U380;
  assign new_P1_R1207_U109 = ~new_P1_R1207_U402 | ~new_P1_R1207_U401;
  assign new_P1_R1207_U110 = ~new_P1_R1207_U419 | ~new_P1_R1207_U418;
  assign new_P1_R1207_U111 = ~new_P1_R1207_U423 | ~new_P1_R1207_U422;
  assign new_P1_R1207_U112 = ~new_P1_R1207_U455 | ~new_P1_R1207_U454;
  assign new_P1_R1207_U113 = ~new_P1_R1207_U459 | ~new_P1_R1207_U458;
  assign new_P1_R1207_U114 = ~new_P1_R1207_U476 | ~new_P1_R1207_U475;
  assign new_P1_R1207_U115 = new_P1_R1207_U195 & new_P1_R1207_U183;
  assign new_P1_R1207_U116 = new_P1_R1207_U198 & new_P1_R1207_U199;
  assign new_P1_R1207_U117 = new_P1_R1207_U211 & new_P1_R1207_U185;
  assign new_P1_R1207_U118 = new_P1_R1207_U214 & new_P1_R1207_U215;
  assign new_P1_R1207_U119 = new_P1_R1207_U40 & new_P1_R1207_U354 & new_P1_R1207_U353;
  assign new_P1_R1207_U120 = new_P1_R1207_U357 & new_P1_R1207_U185;
  assign new_P1_R1207_U121 = new_P1_R1207_U230 & new_P1_R1207_U7;
  assign new_P1_R1207_U122 = new_P1_R1207_U364 & new_P1_R1207_U184;
  assign new_P1_R1207_U123 = new_P1_R1207_U29 & new_P1_R1207_U374 & new_P1_R1207_U373;
  assign new_P1_R1207_U124 = new_P1_R1207_U377 & new_P1_R1207_U183;
  assign new_P1_R1207_U125 = new_P1_R1207_U217 & new_P1_R1207_U8;
  assign new_P1_R1207_U126 = new_P1_R1207_U262 & new_P1_R1207_U180;
  assign new_P1_R1207_U127 = new_P1_R1207_U288 & new_P1_R1207_U181;
  assign new_P1_R1207_U128 = new_P1_R1207_U304 & new_P1_R1207_U305;
  assign new_P1_R1207_U129 = new_P1_R1207_U307 & new_P1_R1207_U386;
  assign new_P1_R1207_U130 = new_P1_R1207_U308 & new_P1_R1207_U305 & new_P1_R1207_U304;
  assign new_P1_R1207_U131 = ~new_P1_R1207_U390 | ~new_P1_R1207_U389;
  assign new_P1_R1207_U132 = new_P1_R1207_U85 & new_P1_R1207_U395 & new_P1_R1207_U394;
  assign new_P1_R1207_U133 = new_P1_R1207_U398 & new_P1_R1207_U182;
  assign new_P1_R1207_U134 = ~new_P1_R1207_U404 | ~new_P1_R1207_U403;
  assign new_P1_R1207_U135 = ~new_P1_R1207_U409 | ~new_P1_R1207_U408;
  assign new_P1_R1207_U136 = new_P1_R1207_U415 & new_P1_R1207_U181;
  assign new_P1_R1207_U137 = ~new_P1_R1207_U425 | ~new_P1_R1207_U424;
  assign new_P1_R1207_U138 = ~new_P1_R1207_U430 | ~new_P1_R1207_U429;
  assign new_P1_R1207_U139 = ~new_P1_R1207_U435 | ~new_P1_R1207_U434;
  assign new_P1_R1207_U140 = ~new_P1_R1207_U440 | ~new_P1_R1207_U439;
  assign new_P1_R1207_U141 = ~new_P1_R1207_U445 | ~new_P1_R1207_U444;
  assign new_P1_R1207_U142 = new_P1_R1207_U451 & new_P1_R1207_U180;
  assign new_P1_R1207_U143 = ~new_P1_R1207_U461 | ~new_P1_R1207_U460;
  assign new_P1_R1207_U144 = ~new_P1_R1207_U466 | ~new_P1_R1207_U465;
  assign new_P1_R1207_U145 = new_P1_R1207_U342 & new_P1_R1207_U9;
  assign new_P1_R1207_U146 = new_P1_R1207_U472 & new_P1_R1207_U179;
  assign new_P1_R1207_U147 = new_P1_R1207_U350 & new_P1_R1207_U349;
  assign new_P1_R1207_U148 = ~new_P1_R1207_U118 | ~new_P1_R1207_U212;
  assign new_P1_R1207_U149 = new_P1_R1207_U359 & new_P1_R1207_U358;
  assign new_P1_R1207_U150 = new_P1_R1207_U366 & new_P1_R1207_U365;
  assign new_P1_R1207_U151 = new_P1_R1207_U370 & new_P1_R1207_U369;
  assign new_P1_R1207_U152 = ~new_P1_R1207_U116 | ~new_P1_R1207_U196;
  assign new_P1_R1207_U153 = new_P1_R1207_U379 & new_P1_R1207_U378;
  assign new_P1_R1207_U154 = ~new_P1_U4028;
  assign new_P1_R1207_U155 = ~new_P1_U3055;
  assign new_P1_R1207_U156 = new_P1_R1207_U388 & new_P1_R1207_U387;
  assign new_P1_R1207_U157 = ~new_P1_R1207_U128 | ~new_P1_R1207_U302;
  assign new_P1_R1207_U158 = new_P1_R1207_U400 & new_P1_R1207_U399;
  assign new_P1_R1207_U159 = ~new_P1_R1207_U295 | ~new_P1_R1207_U294;
  assign new_P1_R1207_U160 = ~new_P1_R1207_U291 | ~new_P1_R1207_U290;
  assign new_P1_R1207_U161 = new_P1_R1207_U417 & new_P1_R1207_U416;
  assign new_P1_R1207_U162 = new_P1_R1207_U421 & new_P1_R1207_U420;
  assign new_P1_R1207_U163 = ~new_P1_R1207_U281 | ~new_P1_R1207_U280;
  assign new_P1_R1207_U164 = ~new_P1_R1207_U277 | ~new_P1_R1207_U276;
  assign new_P1_R1207_U165 = ~new_P1_U3461;
  assign new_P1_R1207_U166 = ~new_P1_R1207_U273 | ~new_P1_R1207_U272;
  assign new_P1_R1207_U167 = ~new_P1_U3512;
  assign new_P1_R1207_U168 = ~new_P1_R1207_U265 | ~new_P1_R1207_U264;
  assign new_P1_R1207_U169 = new_P1_R1207_U453 & new_P1_R1207_U452;
  assign new_P1_R1207_U170 = new_P1_R1207_U457 & new_P1_R1207_U456;
  assign new_P1_R1207_U171 = ~new_P1_R1207_U255 | ~new_P1_R1207_U254;
  assign new_P1_R1207_U172 = ~new_P1_R1207_U251 | ~new_P1_R1207_U250;
  assign new_P1_R1207_U173 = ~new_P1_R1207_U247 | ~new_P1_R1207_U246;
  assign new_P1_R1207_U174 = new_P1_R1207_U474 & new_P1_R1207_U473;
  assign new_P1_R1207_U175 = ~new_P1_R1207_U129 | ~new_P1_R1207_U157;
  assign new_P1_R1207_U176 = ~new_P1_R1207_U85;
  assign new_P1_R1207_U177 = ~new_P1_R1207_U29;
  assign new_P1_R1207_U178 = ~new_P1_R1207_U40;
  assign new_P1_R1207_U179 = ~new_P1_U3488 | ~new_P1_R1207_U53;
  assign new_P1_R1207_U180 = ~new_P1_U3503 | ~new_P1_R1207_U62;
  assign new_P1_R1207_U181 = ~new_P1_U4023 | ~new_P1_R1207_U76;
  assign new_P1_R1207_U182 = ~new_P1_U4019 | ~new_P1_R1207_U84;
  assign new_P1_R1207_U183 = ~new_P1_U3464 | ~new_P1_R1207_U28;
  assign new_P1_R1207_U184 = ~new_P1_U3473 | ~new_P1_R1207_U35;
  assign new_P1_R1207_U185 = ~new_P1_U3479 | ~new_P1_R1207_U39;
  assign new_P1_R1207_U186 = ~new_P1_R1207_U64;
  assign new_P1_R1207_U187 = ~new_P1_R1207_U78;
  assign new_P1_R1207_U188 = ~new_P1_R1207_U37;
  assign new_P1_R1207_U189 = ~new_P1_R1207_U54;
  assign new_P1_R1207_U190 = ~new_P1_R1207_U25;
  assign new_P1_R1207_U191 = ~new_P1_R1207_U190 | ~new_P1_R1207_U26;
  assign new_P1_R1207_U192 = ~new_P1_R1207_U191 | ~new_P1_R1207_U165;
  assign new_P1_R1207_U193 = ~new_P1_U3078 | ~new_P1_R1207_U25;
  assign new_P1_R1207_U194 = ~new_P1_R1207_U46;
  assign new_P1_R1207_U195 = ~new_P1_U3467 | ~new_P1_R1207_U30;
  assign new_P1_R1207_U196 = ~new_P1_R1207_U115 | ~new_P1_R1207_U46;
  assign new_P1_R1207_U197 = ~new_P1_R1207_U30 | ~new_P1_R1207_U29;
  assign new_P1_R1207_U198 = ~new_P1_R1207_U197 | ~new_P1_R1207_U27;
  assign new_P1_R1207_U199 = ~new_P1_U3064 | ~new_P1_R1207_U177;
  assign new_P1_R1207_U200 = ~new_P1_R1207_U152;
  assign new_P1_R1207_U201 = ~new_P1_U3476 | ~new_P1_R1207_U34;
  assign new_P1_R1207_U202 = ~new_P1_U3071 | ~new_P1_R1207_U31;
  assign new_P1_R1207_U203 = ~new_P1_U3067 | ~new_P1_R1207_U32;
  assign new_P1_R1207_U204 = ~new_P1_R1207_U188 | ~new_P1_R1207_U6;
  assign new_P1_R1207_U205 = ~new_P1_R1207_U7 | ~new_P1_R1207_U204;
  assign new_P1_R1207_U206 = ~new_P1_U3470 | ~new_P1_R1207_U36;
  assign new_P1_R1207_U207 = ~new_P1_U3476 | ~new_P1_R1207_U34;
  assign new_P1_R1207_U208 = ~new_P1_R1207_U6 | ~new_P1_R1207_U206 | ~new_P1_R1207_U152;
  assign new_P1_R1207_U209 = ~new_P1_R1207_U207 | ~new_P1_R1207_U205;
  assign new_P1_R1207_U210 = ~new_P1_R1207_U44;
  assign new_P1_R1207_U211 = ~new_P1_U3482 | ~new_P1_R1207_U41;
  assign new_P1_R1207_U212 = ~new_P1_R1207_U117 | ~new_P1_R1207_U44;
  assign new_P1_R1207_U213 = ~new_P1_R1207_U41 | ~new_P1_R1207_U40;
  assign new_P1_R1207_U214 = ~new_P1_R1207_U213 | ~new_P1_R1207_U38;
  assign new_P1_R1207_U215 = ~new_P1_U3084 | ~new_P1_R1207_U178;
  assign new_P1_R1207_U216 = ~new_P1_R1207_U148;
  assign new_P1_R1207_U217 = ~new_P1_U3485 | ~new_P1_R1207_U43;
  assign new_P1_R1207_U218 = ~new_P1_R1207_U217 | ~new_P1_R1207_U54;
  assign new_P1_R1207_U219 = ~new_P1_R1207_U210 | ~new_P1_R1207_U40;
  assign new_P1_R1207_U220 = ~new_P1_R1207_U120 | ~new_P1_R1207_U219;
  assign new_P1_R1207_U221 = ~new_P1_R1207_U44 | ~new_P1_R1207_U185;
  assign new_P1_R1207_U222 = ~new_P1_R1207_U119 | ~new_P1_R1207_U221;
  assign new_P1_R1207_U223 = ~new_P1_R1207_U40 | ~new_P1_R1207_U185;
  assign new_P1_R1207_U224 = ~new_P1_R1207_U206 | ~new_P1_R1207_U152;
  assign new_P1_R1207_U225 = ~new_P1_R1207_U45;
  assign new_P1_R1207_U226 = ~new_P1_U3067 | ~new_P1_R1207_U32;
  assign new_P1_R1207_U227 = ~new_P1_R1207_U225 | ~new_P1_R1207_U226;
  assign new_P1_R1207_U228 = ~new_P1_R1207_U122 | ~new_P1_R1207_U227;
  assign new_P1_R1207_U229 = ~new_P1_R1207_U45 | ~new_P1_R1207_U184;
  assign new_P1_R1207_U230 = ~new_P1_U3476 | ~new_P1_R1207_U34;
  assign new_P1_R1207_U231 = ~new_P1_R1207_U121 | ~new_P1_R1207_U229;
  assign new_P1_R1207_U232 = ~new_P1_U3067 | ~new_P1_R1207_U32;
  assign new_P1_R1207_U233 = ~new_P1_R1207_U184 | ~new_P1_R1207_U232;
  assign new_P1_R1207_U234 = ~new_P1_R1207_U206 | ~new_P1_R1207_U37;
  assign new_P1_R1207_U235 = ~new_P1_R1207_U194 | ~new_P1_R1207_U29;
  assign new_P1_R1207_U236 = ~new_P1_R1207_U124 | ~new_P1_R1207_U235;
  assign new_P1_R1207_U237 = ~new_P1_R1207_U46 | ~new_P1_R1207_U183;
  assign new_P1_R1207_U238 = ~new_P1_R1207_U123 | ~new_P1_R1207_U237;
  assign new_P1_R1207_U239 = ~new_P1_R1207_U29 | ~new_P1_R1207_U183;
  assign new_P1_R1207_U240 = ~new_P1_U3491 | ~new_P1_R1207_U52;
  assign new_P1_R1207_U241 = ~new_P1_U3063 | ~new_P1_R1207_U50;
  assign new_P1_R1207_U242 = ~new_P1_U3062 | ~new_P1_R1207_U51;
  assign new_P1_R1207_U243 = ~new_P1_R1207_U189 | ~new_P1_R1207_U8;
  assign new_P1_R1207_U244 = ~new_P1_R1207_U9 | ~new_P1_R1207_U243;
  assign new_P1_R1207_U245 = ~new_P1_U3491 | ~new_P1_R1207_U52;
  assign new_P1_R1207_U246 = ~new_P1_R1207_U125 | ~new_P1_R1207_U148;
  assign new_P1_R1207_U247 = ~new_P1_R1207_U245 | ~new_P1_R1207_U244;
  assign new_P1_R1207_U248 = ~new_P1_R1207_U173;
  assign new_P1_R1207_U249 = ~new_P1_U3494 | ~new_P1_R1207_U56;
  assign new_P1_R1207_U250 = ~new_P1_R1207_U249 | ~new_P1_R1207_U173;
  assign new_P1_R1207_U251 = ~new_P1_U3072 | ~new_P1_R1207_U55;
  assign new_P1_R1207_U252 = ~new_P1_R1207_U172;
  assign new_P1_R1207_U253 = ~new_P1_U3497 | ~new_P1_R1207_U58;
  assign new_P1_R1207_U254 = ~new_P1_R1207_U253 | ~new_P1_R1207_U172;
  assign new_P1_R1207_U255 = ~new_P1_U3080 | ~new_P1_R1207_U57;
  assign new_P1_R1207_U256 = ~new_P1_R1207_U171;
  assign new_P1_R1207_U257 = ~new_P1_U3506 | ~new_P1_R1207_U61;
  assign new_P1_R1207_U258 = ~new_P1_U3073 | ~new_P1_R1207_U59;
  assign new_P1_R1207_U259 = ~new_P1_U3074 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U260 = ~new_P1_R1207_U186 | ~new_P1_R1207_U180;
  assign new_P1_R1207_U261 = ~new_P1_R1207_U10 | ~new_P1_R1207_U260;
  assign new_P1_R1207_U262 = ~new_P1_U3500 | ~new_P1_R1207_U63;
  assign new_P1_R1207_U263 = ~new_P1_U3506 | ~new_P1_R1207_U61;
  assign new_P1_R1207_U264 = ~new_P1_R1207_U257 | ~new_P1_R1207_U171 | ~new_P1_R1207_U126;
  assign new_P1_R1207_U265 = ~new_P1_R1207_U263 | ~new_P1_R1207_U261;
  assign new_P1_R1207_U266 = ~new_P1_R1207_U168;
  assign new_P1_R1207_U267 = ~new_P1_U3509 | ~new_P1_R1207_U66;
  assign new_P1_R1207_U268 = ~new_P1_R1207_U267 | ~new_P1_R1207_U168;
  assign new_P1_R1207_U269 = ~new_P1_U3069 | ~new_P1_R1207_U65;
  assign new_P1_R1207_U270 = ~new_P1_R1207_U67;
  assign new_P1_R1207_U271 = ~new_P1_R1207_U270 | ~new_P1_R1207_U68;
  assign new_P1_R1207_U272 = ~new_P1_R1207_U271 | ~new_P1_R1207_U167;
  assign new_P1_R1207_U273 = ~new_P1_U3082 | ~new_P1_R1207_U67;
  assign new_P1_R1207_U274 = ~new_P1_R1207_U166;
  assign new_P1_R1207_U275 = ~new_P1_U3514 | ~new_P1_R1207_U70;
  assign new_P1_R1207_U276 = ~new_P1_R1207_U275 | ~new_P1_R1207_U166;
  assign new_P1_R1207_U277 = ~new_P1_U3081 | ~new_P1_R1207_U69;
  assign new_P1_R1207_U278 = ~new_P1_R1207_U164;
  assign new_P1_R1207_U279 = ~new_P1_U4025 | ~new_P1_R1207_U72;
  assign new_P1_R1207_U280 = ~new_P1_R1207_U279 | ~new_P1_R1207_U164;
  assign new_P1_R1207_U281 = ~new_P1_U3076 | ~new_P1_R1207_U71;
  assign new_P1_R1207_U282 = ~new_P1_R1207_U163;
  assign new_P1_R1207_U283 = ~new_P1_U4022 | ~new_P1_R1207_U75;
  assign new_P1_R1207_U284 = ~new_P1_U3066 | ~new_P1_R1207_U73;
  assign new_P1_R1207_U285 = ~new_P1_U3061 | ~new_P1_R1207_U48;
  assign new_P1_R1207_U286 = ~new_P1_R1207_U187 | ~new_P1_R1207_U181;
  assign new_P1_R1207_U287 = ~new_P1_R1207_U11 | ~new_P1_R1207_U286;
  assign new_P1_R1207_U288 = ~new_P1_U4024 | ~new_P1_R1207_U77;
  assign new_P1_R1207_U289 = ~new_P1_U4022 | ~new_P1_R1207_U75;
  assign new_P1_R1207_U290 = ~new_P1_R1207_U283 | ~new_P1_R1207_U163 | ~new_P1_R1207_U127;
  assign new_P1_R1207_U291 = ~new_P1_R1207_U289 | ~new_P1_R1207_U287;
  assign new_P1_R1207_U292 = ~new_P1_R1207_U160;
  assign new_P1_R1207_U293 = ~new_P1_U4021 | ~new_P1_R1207_U80;
  assign new_P1_R1207_U294 = ~new_P1_R1207_U293 | ~new_P1_R1207_U160;
  assign new_P1_R1207_U295 = ~new_P1_U3065 | ~new_P1_R1207_U79;
  assign new_P1_R1207_U296 = ~new_P1_R1207_U159;
  assign new_P1_R1207_U297 = ~new_P1_U4020 | ~new_P1_R1207_U82;
  assign new_P1_R1207_U298 = ~new_P1_R1207_U297 | ~new_P1_R1207_U159;
  assign new_P1_R1207_U299 = ~new_P1_U3058 | ~new_P1_R1207_U81;
  assign new_P1_R1207_U300 = ~new_P1_R1207_U89;
  assign new_P1_R1207_U301 = ~new_P1_U4018 | ~new_P1_R1207_U86;
  assign new_P1_R1207_U302 = ~new_P1_R1207_U301 | ~new_P1_R1207_U89 | ~new_P1_R1207_U182;
  assign new_P1_R1207_U303 = ~new_P1_R1207_U86 | ~new_P1_R1207_U85;
  assign new_P1_R1207_U304 = ~new_P1_R1207_U303 | ~new_P1_R1207_U83;
  assign new_P1_R1207_U305 = ~new_P1_U3053 | ~new_P1_R1207_U176;
  assign new_P1_R1207_U306 = ~new_P1_R1207_U157;
  assign new_P1_R1207_U307 = ~new_P1_U4017 | ~new_P1_R1207_U88;
  assign new_P1_R1207_U308 = ~new_P1_U3054 | ~new_P1_R1207_U87;
  assign new_P1_R1207_U309 = ~new_P1_R1207_U300 | ~new_P1_R1207_U85;
  assign new_P1_R1207_U310 = ~new_P1_R1207_U133 | ~new_P1_R1207_U309;
  assign new_P1_R1207_U311 = ~new_P1_R1207_U89 | ~new_P1_R1207_U182;
  assign new_P1_R1207_U312 = ~new_P1_R1207_U132 | ~new_P1_R1207_U311;
  assign new_P1_R1207_U313 = ~new_P1_R1207_U85 | ~new_P1_R1207_U182;
  assign new_P1_R1207_U314 = ~new_P1_R1207_U288 | ~new_P1_R1207_U163;
  assign new_P1_R1207_U315 = ~new_P1_R1207_U90;
  assign new_P1_R1207_U316 = ~new_P1_U3061 | ~new_P1_R1207_U48;
  assign new_P1_R1207_U317 = ~new_P1_R1207_U315 | ~new_P1_R1207_U316;
  assign new_P1_R1207_U318 = ~new_P1_R1207_U136 | ~new_P1_R1207_U317;
  assign new_P1_R1207_U319 = ~new_P1_R1207_U90 | ~new_P1_R1207_U181;
  assign new_P1_R1207_U320 = ~new_P1_U4022 | ~new_P1_R1207_U75;
  assign new_P1_R1207_U321 = ~new_P1_R1207_U11 | ~new_P1_R1207_U320 | ~new_P1_R1207_U319;
  assign new_P1_R1207_U322 = ~new_P1_U3061 | ~new_P1_R1207_U48;
  assign new_P1_R1207_U323 = ~new_P1_R1207_U181 | ~new_P1_R1207_U322;
  assign new_P1_R1207_U324 = ~new_P1_R1207_U288 | ~new_P1_R1207_U78;
  assign new_P1_R1207_U325 = ~new_P1_R1207_U262 | ~new_P1_R1207_U171;
  assign new_P1_R1207_U326 = ~new_P1_R1207_U91;
  assign new_P1_R1207_U327 = ~new_P1_U3074 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U328 = ~new_P1_R1207_U326 | ~new_P1_R1207_U327;
  assign new_P1_R1207_U329 = ~new_P1_R1207_U142 | ~new_P1_R1207_U328;
  assign new_P1_R1207_U330 = ~new_P1_R1207_U91 | ~new_P1_R1207_U180;
  assign new_P1_R1207_U331 = ~new_P1_U3506 | ~new_P1_R1207_U61;
  assign new_P1_R1207_U332 = ~new_P1_R1207_U10 | ~new_P1_R1207_U331 | ~new_P1_R1207_U330;
  assign new_P1_R1207_U333 = ~new_P1_U3074 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U334 = ~new_P1_R1207_U180 | ~new_P1_R1207_U333;
  assign new_P1_R1207_U335 = ~new_P1_R1207_U262 | ~new_P1_R1207_U64;
  assign new_P1_R1207_U336 = ~new_P1_R1207_U217 | ~new_P1_R1207_U148;
  assign new_P1_R1207_U337 = ~new_P1_R1207_U92;
  assign new_P1_R1207_U338 = ~new_P1_U3062 | ~new_P1_R1207_U51;
  assign new_P1_R1207_U339 = ~new_P1_R1207_U337 | ~new_P1_R1207_U338;
  assign new_P1_R1207_U340 = ~new_P1_R1207_U146 | ~new_P1_R1207_U339;
  assign new_P1_R1207_U341 = ~new_P1_R1207_U92 | ~new_P1_R1207_U179;
  assign new_P1_R1207_U342 = ~new_P1_U3491 | ~new_P1_R1207_U52;
  assign new_P1_R1207_U343 = ~new_P1_R1207_U145 | ~new_P1_R1207_U341;
  assign new_P1_R1207_U344 = ~new_P1_U3062 | ~new_P1_R1207_U51;
  assign new_P1_R1207_U345 = ~new_P1_R1207_U179 | ~new_P1_R1207_U344;
  assign new_P1_R1207_U346 = ~new_P1_U3077 | ~new_P1_R1207_U24;
  assign new_P1_R1207_U347 = ~new_P1_R1207_U301 | ~new_P1_R1207_U89 | ~new_P1_R1207_U182;
  assign new_P1_R1207_U348 = ~new_P1_R1207_U130 | ~new_P1_R1207_U12 | ~new_P1_R1207_U347;
  assign new_P1_R1207_U349 = ~new_P1_U3485 | ~new_P1_R1207_U43;
  assign new_P1_R1207_U350 = ~new_P1_U3083 | ~new_P1_R1207_U42;
  assign new_P1_R1207_U351 = ~new_P1_R1207_U218 | ~new_P1_R1207_U148;
  assign new_P1_R1207_U352 = ~new_P1_R1207_U216 | ~new_P1_R1207_U147;
  assign new_P1_R1207_U353 = ~new_P1_U3482 | ~new_P1_R1207_U41;
  assign new_P1_R1207_U354 = ~new_P1_U3084 | ~new_P1_R1207_U38;
  assign new_P1_R1207_U355 = ~new_P1_U3482 | ~new_P1_R1207_U41;
  assign new_P1_R1207_U356 = ~new_P1_U3084 | ~new_P1_R1207_U38;
  assign new_P1_R1207_U357 = ~new_P1_R1207_U356 | ~new_P1_R1207_U355;
  assign new_P1_R1207_U358 = ~new_P1_U3479 | ~new_P1_R1207_U39;
  assign new_P1_R1207_U359 = ~new_P1_U3070 | ~new_P1_R1207_U22;
  assign new_P1_R1207_U360 = ~new_P1_R1207_U223 | ~new_P1_R1207_U44;
  assign new_P1_R1207_U361 = ~new_P1_R1207_U149 | ~new_P1_R1207_U210;
  assign new_P1_R1207_U362 = ~new_P1_U3476 | ~new_P1_R1207_U34;
  assign new_P1_R1207_U363 = ~new_P1_U3071 | ~new_P1_R1207_U31;
  assign new_P1_R1207_U364 = ~new_P1_R1207_U363 | ~new_P1_R1207_U362;
  assign new_P1_R1207_U365 = ~new_P1_U3473 | ~new_P1_R1207_U35;
  assign new_P1_R1207_U366 = ~new_P1_U3067 | ~new_P1_R1207_U32;
  assign new_P1_R1207_U367 = ~new_P1_R1207_U233 | ~new_P1_R1207_U45;
  assign new_P1_R1207_U368 = ~new_P1_R1207_U150 | ~new_P1_R1207_U225;
  assign new_P1_R1207_U369 = ~new_P1_U3470 | ~new_P1_R1207_U36;
  assign new_P1_R1207_U370 = ~new_P1_U3060 | ~new_P1_R1207_U33;
  assign new_P1_R1207_U371 = ~new_P1_R1207_U234 | ~new_P1_R1207_U152;
  assign new_P1_R1207_U372 = ~new_P1_R1207_U200 | ~new_P1_R1207_U151;
  assign new_P1_R1207_U373 = ~new_P1_U3467 | ~new_P1_R1207_U30;
  assign new_P1_R1207_U374 = ~new_P1_U3064 | ~new_P1_R1207_U27;
  assign new_P1_R1207_U375 = ~new_P1_U3467 | ~new_P1_R1207_U30;
  assign new_P1_R1207_U376 = ~new_P1_U3064 | ~new_P1_R1207_U27;
  assign new_P1_R1207_U377 = ~new_P1_R1207_U376 | ~new_P1_R1207_U375;
  assign new_P1_R1207_U378 = ~new_P1_U3464 | ~new_P1_R1207_U28;
  assign new_P1_R1207_U379 = ~new_P1_U3068 | ~new_P1_R1207_U23;
  assign new_P1_R1207_U380 = ~new_P1_R1207_U239 | ~new_P1_R1207_U46;
  assign new_P1_R1207_U381 = ~new_P1_R1207_U153 | ~new_P1_R1207_U194;
  assign new_P1_R1207_U382 = ~new_P1_U4028 | ~new_P1_R1207_U155;
  assign new_P1_R1207_U383 = ~new_P1_U3055 | ~new_P1_R1207_U154;
  assign new_P1_R1207_U384 = ~new_P1_U4028 | ~new_P1_R1207_U155;
  assign new_P1_R1207_U385 = ~new_P1_U3055 | ~new_P1_R1207_U154;
  assign new_P1_R1207_U386 = ~new_P1_R1207_U385 | ~new_P1_R1207_U384;
  assign new_P1_R1207_U387 = ~new_P1_R1207_U87 | ~new_P1_U3054 | ~new_P1_R1207_U386;
  assign new_P1_R1207_U388 = ~new_P1_U4017 | ~new_P1_R1207_U12 | ~new_P1_R1207_U88;
  assign new_P1_R1207_U389 = ~new_P1_U4017 | ~new_P1_R1207_U88;
  assign new_P1_R1207_U390 = ~new_P1_U3054 | ~new_P1_R1207_U87;
  assign new_P1_R1207_U391 = ~new_P1_R1207_U131;
  assign new_P1_R1207_U392 = ~new_P1_R1207_U306 | ~new_P1_R1207_U391;
  assign new_P1_R1207_U393 = ~new_P1_R1207_U131 | ~new_P1_R1207_U157;
  assign new_P1_R1207_U394 = ~new_P1_U4018 | ~new_P1_R1207_U86;
  assign new_P1_R1207_U395 = ~new_P1_U3053 | ~new_P1_R1207_U83;
  assign new_P1_R1207_U396 = ~new_P1_U4018 | ~new_P1_R1207_U86;
  assign new_P1_R1207_U397 = ~new_P1_U3053 | ~new_P1_R1207_U83;
  assign new_P1_R1207_U398 = ~new_P1_R1207_U397 | ~new_P1_R1207_U396;
  assign new_P1_R1207_U399 = ~new_P1_U4019 | ~new_P1_R1207_U84;
  assign new_P1_R1207_U400 = ~new_P1_U3057 | ~new_P1_R1207_U47;
  assign new_P1_R1207_U401 = ~new_P1_R1207_U313 | ~new_P1_R1207_U89;
  assign new_P1_R1207_U402 = ~new_P1_R1207_U158 | ~new_P1_R1207_U300;
  assign new_P1_R1207_U403 = ~new_P1_U4020 | ~new_P1_R1207_U82;
  assign new_P1_R1207_U404 = ~new_P1_U3058 | ~new_P1_R1207_U81;
  assign new_P1_R1207_U405 = ~new_P1_R1207_U134;
  assign new_P1_R1207_U406 = ~new_P1_R1207_U296 | ~new_P1_R1207_U405;
  assign new_P1_R1207_U407 = ~new_P1_R1207_U134 | ~new_P1_R1207_U159;
  assign new_P1_R1207_U408 = ~new_P1_U4021 | ~new_P1_R1207_U80;
  assign new_P1_R1207_U409 = ~new_P1_U3065 | ~new_P1_R1207_U79;
  assign new_P1_R1207_U410 = ~new_P1_R1207_U135;
  assign new_P1_R1207_U411 = ~new_P1_R1207_U292 | ~new_P1_R1207_U410;
  assign new_P1_R1207_U412 = ~new_P1_R1207_U135 | ~new_P1_R1207_U160;
  assign new_P1_R1207_U413 = ~new_P1_U4022 | ~new_P1_R1207_U75;
  assign new_P1_R1207_U414 = ~new_P1_U3066 | ~new_P1_R1207_U73;
  assign new_P1_R1207_U415 = ~new_P1_R1207_U414 | ~new_P1_R1207_U413;
  assign new_P1_R1207_U416 = ~new_P1_U4023 | ~new_P1_R1207_U76;
  assign new_P1_R1207_U417 = ~new_P1_U3061 | ~new_P1_R1207_U48;
  assign new_P1_R1207_U418 = ~new_P1_R1207_U323 | ~new_P1_R1207_U90;
  assign new_P1_R1207_U419 = ~new_P1_R1207_U161 | ~new_P1_R1207_U315;
  assign new_P1_R1207_U420 = ~new_P1_U4024 | ~new_P1_R1207_U77;
  assign new_P1_R1207_U421 = ~new_P1_U3075 | ~new_P1_R1207_U74;
  assign new_P1_R1207_U422 = ~new_P1_R1207_U324 | ~new_P1_R1207_U163;
  assign new_P1_R1207_U423 = ~new_P1_R1207_U282 | ~new_P1_R1207_U162;
  assign new_P1_R1207_U424 = ~new_P1_U4025 | ~new_P1_R1207_U72;
  assign new_P1_R1207_U425 = ~new_P1_U3076 | ~new_P1_R1207_U71;
  assign new_P1_R1207_U426 = ~new_P1_R1207_U137;
  assign new_P1_R1207_U427 = ~new_P1_R1207_U278 | ~new_P1_R1207_U426;
  assign new_P1_R1207_U428 = ~new_P1_R1207_U137 | ~new_P1_R1207_U164;
  assign new_P1_R1207_U429 = ~new_P1_U3461 | ~new_P1_R1207_U26;
  assign new_P1_R1207_U430 = ~new_P1_U3078 | ~new_P1_R1207_U165;
  assign new_P1_R1207_U431 = ~new_P1_R1207_U138;
  assign new_P1_R1207_U432 = ~new_P1_R1207_U431 | ~new_P1_R1207_U190;
  assign new_P1_R1207_U433 = ~new_P1_R1207_U138 | ~new_P1_R1207_U25;
  assign new_P1_R1207_U434 = ~new_P1_U3514 | ~new_P1_R1207_U70;
  assign new_P1_R1207_U435 = ~new_P1_U3081 | ~new_P1_R1207_U69;
  assign new_P1_R1207_U436 = ~new_P1_R1207_U139;
  assign new_P1_R1207_U437 = ~new_P1_R1207_U274 | ~new_P1_R1207_U436;
  assign new_P1_R1207_U438 = ~new_P1_R1207_U139 | ~new_P1_R1207_U166;
  assign new_P1_R1207_U439 = ~new_P1_U3512 | ~new_P1_R1207_U68;
  assign new_P1_R1207_U440 = ~new_P1_U3082 | ~new_P1_R1207_U167;
  assign new_P1_R1207_U441 = ~new_P1_R1207_U140;
  assign new_P1_R1207_U442 = ~new_P1_R1207_U441 | ~new_P1_R1207_U270;
  assign new_P1_R1207_U443 = ~new_P1_R1207_U140 | ~new_P1_R1207_U67;
  assign new_P1_R1207_U444 = ~new_P1_U3509 | ~new_P1_R1207_U66;
  assign new_P1_R1207_U445 = ~new_P1_U3069 | ~new_P1_R1207_U65;
  assign new_P1_R1207_U446 = ~new_P1_R1207_U141;
  assign new_P1_R1207_U447 = ~new_P1_R1207_U266 | ~new_P1_R1207_U446;
  assign new_P1_R1207_U448 = ~new_P1_R1207_U141 | ~new_P1_R1207_U168;
  assign new_P1_R1207_U449 = ~new_P1_U3506 | ~new_P1_R1207_U61;
  assign new_P1_R1207_U450 = ~new_P1_U3073 | ~new_P1_R1207_U59;
  assign new_P1_R1207_U451 = ~new_P1_R1207_U450 | ~new_P1_R1207_U449;
  assign new_P1_R1207_U452 = ~new_P1_U3503 | ~new_P1_R1207_U62;
  assign new_P1_R1207_U453 = ~new_P1_U3074 | ~new_P1_R1207_U49;
  assign new_P1_R1207_U454 = ~new_P1_R1207_U334 | ~new_P1_R1207_U91;
  assign new_P1_R1207_U455 = ~new_P1_R1207_U169 | ~new_P1_R1207_U326;
  assign new_P1_R1207_U456 = ~new_P1_U3500 | ~new_P1_R1207_U63;
  assign new_P1_R1207_U457 = ~new_P1_U3079 | ~new_P1_R1207_U60;
  assign new_P1_R1207_U458 = ~new_P1_R1207_U335 | ~new_P1_R1207_U171;
  assign new_P1_R1207_U459 = ~new_P1_R1207_U256 | ~new_P1_R1207_U170;
  assign new_P1_R1207_U460 = ~new_P1_U3497 | ~new_P1_R1207_U58;
  assign new_P1_R1207_U461 = ~new_P1_U3080 | ~new_P1_R1207_U57;
  assign new_P1_R1207_U462 = ~new_P1_R1207_U143;
  assign new_P1_R1207_U463 = ~new_P1_R1207_U252 | ~new_P1_R1207_U462;
  assign new_P1_R1207_U464 = ~new_P1_R1207_U143 | ~new_P1_R1207_U172;
  assign new_P1_R1207_U465 = ~new_P1_U3494 | ~new_P1_R1207_U56;
  assign new_P1_R1207_U466 = ~new_P1_U3072 | ~new_P1_R1207_U55;
  assign new_P1_R1207_U467 = ~new_P1_R1207_U144;
  assign new_P1_R1207_U468 = ~new_P1_R1207_U248 | ~new_P1_R1207_U467;
  assign new_P1_R1207_U469 = ~new_P1_R1207_U144 | ~new_P1_R1207_U173;
  assign new_P1_R1207_U470 = ~new_P1_U3491 | ~new_P1_R1207_U52;
  assign new_P1_R1207_U471 = ~new_P1_U3063 | ~new_P1_R1207_U50;
  assign new_P1_R1207_U472 = ~new_P1_R1207_U471 | ~new_P1_R1207_U470;
  assign new_P1_R1207_U473 = ~new_P1_U3488 | ~new_P1_R1207_U53;
  assign new_P1_R1207_U474 = ~new_P1_U3062 | ~new_P1_R1207_U51;
  assign new_P1_R1207_U475 = ~new_P1_R1207_U345 | ~new_P1_R1207_U92;
  assign new_P1_R1207_U476 = ~new_P1_R1207_U174 | ~new_P1_R1207_U337;
  assign new_P1_R1165_U4 = new_P1_R1165_U202 & new_P1_R1165_U201;
  assign new_P1_R1165_U5 = new_P1_R1165_U217 & new_P1_R1165_U216;
  assign new_P1_R1165_U6 = new_P1_R1165_U251 & new_P1_R1165_U250;
  assign new_P1_R1165_U7 = new_P1_R1165_U269 & new_P1_R1165_U268;
  assign new_P1_R1165_U8 = new_P1_R1165_U281 & new_P1_R1165_U280;
  assign new_P1_R1165_U9 = new_P1_R1165_U339 & new_P1_R1165_U336;
  assign new_P1_R1165_U10 = new_P1_R1165_U330 & new_P1_R1165_U327;
  assign new_P1_R1165_U11 = new_P1_R1165_U323 & new_P1_R1165_U320;
  assign new_P1_R1165_U12 = new_P1_R1165_U314 & new_P1_R1165_U311;
  assign new_P1_R1165_U13 = new_P1_R1165_U240 & new_P1_R1165_U237;
  assign new_P1_R1165_U14 = new_P1_R1165_U233 & new_P1_R1165_U230;
  assign new_P1_R1165_U15 = ~new_P1_U3211;
  assign new_P1_R1165_U16 = ~new_P1_U3175;
  assign new_P1_R1165_U17 = ~new_P1_U3175 | ~new_P1_R1165_U59;
  assign new_P1_R1165_U18 = ~new_P1_U3174;
  assign new_P1_R1165_U19 = ~new_P1_U3179;
  assign new_P1_R1165_U20 = ~new_P1_U3179 | ~new_P1_R1165_U61;
  assign new_P1_R1165_U21 = ~new_P1_U3178;
  assign new_P1_R1165_U22 = ~new_P1_U3181;
  assign new_P1_R1165_U23 = ~new_P1_U3180;
  assign new_P1_R1165_U24 = ~new_P1_R1165_U110 | ~new_P1_R1165_U206;
  assign new_P1_R1165_U25 = ~new_P1_U3177;
  assign new_P1_R1165_U26 = ~new_P1_U3176;
  assign new_P1_R1165_U27 = ~new_P1_U3173;
  assign new_P1_R1165_U28 = ~new_P1_U3172;
  assign new_P1_R1165_U29 = ~new_P1_R1165_U226 | ~new_P1_R1165_U225;
  assign new_P1_R1165_U30 = ~new_P1_R1165_U214 | ~new_P1_R1165_U213;
  assign new_P1_R1165_U31 = ~new_P1_R1165_U199 | ~new_P1_R1165_U198;
  assign new_P1_R1165_U32 = ~new_P1_U3154;
  assign new_P1_R1165_U33 = ~new_P1_U3155;
  assign new_P1_R1165_U34 = ~new_P1_U3156;
  assign new_P1_R1165_U35 = ~new_P1_U3157;
  assign new_P1_R1165_U36 = ~new_P1_U3160;
  assign new_P1_R1165_U37 = ~new_P1_U3165;
  assign new_P1_R1165_U38 = ~new_P1_U3165 | ~new_P1_R1165_U73;
  assign new_P1_R1165_U39 = ~new_P1_U3164;
  assign new_P1_R1165_U40 = ~new_P1_U3171;
  assign new_P1_R1165_U41 = ~new_P1_U3169;
  assign new_P1_R1165_U42 = ~new_P1_U3170;
  assign new_P1_R1165_U43 = ~new_P1_U3170 | ~new_P1_R1165_U76;
  assign new_P1_R1165_U44 = ~new_P1_U3168;
  assign new_P1_R1165_U45 = ~new_P1_U3167;
  assign new_P1_R1165_U46 = ~new_P1_U3166;
  assign new_P1_R1165_U47 = ~new_P1_U3163;
  assign new_P1_R1165_U48 = ~new_P1_U3162;
  assign new_P1_R1165_U49 = ~new_P1_U3162 | ~new_P1_R1165_U82;
  assign new_P1_R1165_U50 = ~new_P1_U3161;
  assign new_P1_R1165_U51 = ~new_P1_U3159;
  assign new_P1_R1165_U52 = ~new_P1_U3158;
  assign new_P1_R1165_U53 = ~new_P1_U3155 | ~new_P1_R1165_U70;
  assign new_P1_R1165_U54 = ~new_P1_R1165_U192 | ~new_P1_R1165_U307;
  assign new_P1_R1165_U55 = ~new_P1_R1165_U49 | ~new_P1_R1165_U316;
  assign new_P1_R1165_U56 = ~new_P1_R1165_U266 | ~new_P1_R1165_U265;
  assign new_P1_R1165_U57 = ~new_P1_R1165_U43 | ~new_P1_R1165_U332;
  assign new_P1_R1165_U58 = ~new_P1_R1165_U359 | ~new_P1_R1165_U358;
  assign new_P1_R1165_U59 = ~new_P1_R1165_U388 | ~new_P1_R1165_U387;
  assign new_P1_R1165_U60 = ~new_P1_R1165_U385 | ~new_P1_R1165_U384;
  assign new_P1_R1165_U61 = ~new_P1_R1165_U376 | ~new_P1_R1165_U375;
  assign new_P1_R1165_U62 = ~new_P1_R1165_U373 | ~new_P1_R1165_U372;
  assign new_P1_R1165_U63 = ~new_P1_R1165_U367 | ~new_P1_R1165_U366;
  assign new_P1_R1165_U64 = ~new_P1_R1165_U370 | ~new_P1_R1165_U369;
  assign new_P1_R1165_U65 = ~new_P1_R1165_U379 | ~new_P1_R1165_U378;
  assign new_P1_R1165_U66 = ~new_P1_R1165_U382 | ~new_P1_R1165_U381;
  assign new_P1_R1165_U67 = ~new_P1_R1165_U391 | ~new_P1_R1165_U390;
  assign new_P1_R1165_U68 = ~new_P1_R1165_U431 | ~new_P1_R1165_U430;
  assign new_P1_R1165_U69 = ~new_P1_R1165_U434 | ~new_P1_R1165_U433;
  assign new_P1_R1165_U70 = ~new_P1_R1165_U437 | ~new_P1_R1165_U436;
  assign new_P1_R1165_U71 = ~new_P1_R1165_U440 | ~new_P1_R1165_U439;
  assign new_P1_R1165_U72 = ~new_P1_R1165_U443 | ~new_P1_R1165_U442;
  assign new_P1_R1165_U73 = ~new_P1_R1165_U473 | ~new_P1_R1165_U472;
  assign new_P1_R1165_U74 = ~new_P1_R1165_U470 | ~new_P1_R1165_U469;
  assign new_P1_R1165_U75 = ~new_P1_R1165_U452 | ~new_P1_R1165_U451;
  assign new_P1_R1165_U76 = ~new_P1_R1165_U461 | ~new_P1_R1165_U460;
  assign new_P1_R1165_U77 = ~new_P1_R1165_U455 | ~new_P1_R1165_U454;
  assign new_P1_R1165_U78 = ~new_P1_R1165_U458 | ~new_P1_R1165_U457;
  assign new_P1_R1165_U79 = ~new_P1_R1165_U464 | ~new_P1_R1165_U463;
  assign new_P1_R1165_U80 = ~new_P1_R1165_U467 | ~new_P1_R1165_U466;
  assign new_P1_R1165_U81 = ~new_P1_R1165_U476 | ~new_P1_R1165_U475;
  assign new_P1_R1165_U82 = ~new_P1_R1165_U449 | ~new_P1_R1165_U448;
  assign new_P1_R1165_U83 = ~new_P1_R1165_U446 | ~new_P1_R1165_U445;
  assign new_P1_R1165_U84 = ~new_P1_R1165_U479 | ~new_P1_R1165_U478;
  assign new_P1_R1165_U85 = ~new_P1_R1165_U482 | ~new_P1_R1165_U481;
  assign new_P1_R1165_U86 = ~new_P1_R1165_U488 | ~new_P1_R1165_U487;
  assign new_P1_R1165_U87 = ~new_P1_R1165_U595 | ~new_P1_R1165_U594;
  assign new_P1_R1165_U88 = ~new_P1_R1165_U394 | ~new_P1_R1165_U393;
  assign new_P1_R1165_U89 = ~new_P1_R1165_U401 | ~new_P1_R1165_U400;
  assign new_P1_R1165_U90 = ~new_P1_R1165_U408 | ~new_P1_R1165_U407;
  assign new_P1_R1165_U91 = ~new_P1_R1165_U415 | ~new_P1_R1165_U414;
  assign new_P1_R1165_U92 = ~new_P1_R1165_U422 | ~new_P1_R1165_U421;
  assign new_P1_R1165_U93 = ~new_P1_R1165_U429 | ~new_P1_R1165_U428;
  assign new_P1_R1165_U94 = ~new_P1_R1165_U491 | ~new_P1_R1165_U490;
  assign new_P1_R1165_U95 = ~new_P1_R1165_U498 | ~new_P1_R1165_U497;
  assign new_P1_R1165_U96 = ~new_P1_R1165_U505 | ~new_P1_R1165_U504;
  assign new_P1_R1165_U97 = ~new_P1_R1165_U510 | ~new_P1_R1165_U509;
  assign new_P1_R1165_U98 = ~new_P1_R1165_U517 | ~new_P1_R1165_U516;
  assign new_P1_R1165_U99 = ~new_P1_R1165_U524 | ~new_P1_R1165_U523;
  assign new_P1_R1165_U100 = ~new_P1_R1165_U531 | ~new_P1_R1165_U530;
  assign new_P1_R1165_U101 = ~new_P1_R1165_U538 | ~new_P1_R1165_U537;
  assign new_P1_R1165_U102 = ~new_P1_R1165_U543 | ~new_P1_R1165_U542;
  assign new_P1_R1165_U103 = ~new_P1_R1165_U550 | ~new_P1_R1165_U549;
  assign new_P1_R1165_U104 = ~new_P1_R1165_U557 | ~new_P1_R1165_U556;
  assign new_P1_R1165_U105 = ~new_P1_R1165_U564 | ~new_P1_R1165_U563;
  assign new_P1_R1165_U106 = ~new_P1_R1165_U571 | ~new_P1_R1165_U570;
  assign new_P1_R1165_U107 = ~new_P1_R1165_U578 | ~new_P1_R1165_U577;
  assign new_P1_R1165_U108 = ~new_P1_R1165_U583 | ~new_P1_R1165_U582;
  assign new_P1_R1165_U109 = ~new_P1_R1165_U590 | ~new_P1_R1165_U589;
  assign new_P1_R1165_U110 = new_P1_R1165_U205 & new_P1_R1165_U204;
  assign new_P1_R1165_U111 = new_P1_R1165_U221 & new_P1_R1165_U220;
  assign new_P1_R1165_U112 = new_P1_R1165_U17 & new_P1_R1165_U403 & new_P1_R1165_U402;
  assign new_P1_R1165_U113 = new_P1_R1165_U232 & new_P1_R1165_U5;
  assign new_P1_R1165_U114 = new_P1_R1165_U20 & new_P1_R1165_U424 & new_P1_R1165_U423;
  assign new_P1_R1165_U115 = new_P1_R1165_U239 & new_P1_R1165_U4;
  assign new_P1_R1165_U116 = new_P1_R1165_U255 & new_P1_R1165_U6;
  assign new_P1_R1165_U117 = new_P1_R1165_U253 & new_P1_R1165_U187;
  assign new_P1_R1165_U118 = new_P1_R1165_U273 & new_P1_R1165_U272;
  assign new_P1_R1165_U119 = new_P1_R1165_U357 & new_P1_R1165_U53;
  assign new_P1_R1165_U120 = new_P1_R1165_U306 & new_P1_R1165_U301;
  assign new_P1_R1165_U121 = new_P1_R1165_U354 & new_P1_R1165_U305;
  assign new_P1_R1165_U122 = ~new_P1_R1165_U485 | ~new_P1_R1165_U484;
  assign new_P1_R1165_U123 = new_P1_R1165_U189 & new_P1_R1165_U500 & new_P1_R1165_U499;
  assign new_P1_R1165_U124 = new_P1_R1165_U188 & new_P1_R1165_U526 & new_P1_R1165_U525;
  assign new_P1_R1165_U125 = new_P1_R1165_U38 & new_P1_R1165_U552 & new_P1_R1165_U551;
  assign new_P1_R1165_U126 = new_P1_R1165_U329 & new_P1_R1165_U7;
  assign new_P1_R1165_U127 = new_P1_R1165_U187 & new_P1_R1165_U573 & new_P1_R1165_U572;
  assign new_P1_R1165_U128 = new_P1_R1165_U338 & new_P1_R1165_U6;
  assign new_P1_R1165_U129 = ~new_P1_R1165_U592 | ~new_P1_R1165_U591;
  assign new_P1_R1165_U130 = ~new_P1_U3201;
  assign new_P1_R1165_U131 = new_P1_R1165_U362 & new_P1_R1165_U361;
  assign new_P1_R1165_U132 = ~new_P1_U3210;
  assign new_P1_R1165_U133 = ~new_P1_U3209;
  assign new_P1_R1165_U134 = ~new_P1_U3207;
  assign new_P1_R1165_U135 = ~new_P1_U3208;
  assign new_P1_R1165_U136 = ~new_P1_U3206;
  assign new_P1_R1165_U137 = ~new_P1_U3205;
  assign new_P1_R1165_U138 = ~new_P1_U3203;
  assign new_P1_R1165_U139 = ~new_P1_U3204;
  assign new_P1_R1165_U140 = ~new_P1_U3202;
  assign new_P1_R1165_U141 = new_P1_R1165_U396 & new_P1_R1165_U395;
  assign new_P1_R1165_U142 = ~new_P1_R1165_U111 | ~new_P1_R1165_U222;
  assign new_P1_R1165_U143 = new_P1_R1165_U410 & new_P1_R1165_U409;
  assign new_P1_R1165_U144 = ~new_P1_R1165_U210 | ~new_P1_R1165_U209;
  assign new_P1_R1165_U145 = new_P1_R1165_U417 & new_P1_R1165_U416;
  assign new_P1_R1165_U146 = ~new_P1_U3183;
  assign new_P1_R1165_U147 = ~new_P1_U3185;
  assign new_P1_R1165_U148 = ~new_P1_U3184;
  assign new_P1_R1165_U149 = ~new_P1_U3186;
  assign new_P1_R1165_U150 = ~new_P1_U3189;
  assign new_P1_R1165_U151 = ~new_P1_U3190;
  assign new_P1_R1165_U152 = ~new_P1_U3191;
  assign new_P1_R1165_U153 = ~new_P1_U3200;
  assign new_P1_R1165_U154 = ~new_P1_U3197;
  assign new_P1_R1165_U155 = ~new_P1_U3198;
  assign new_P1_R1165_U156 = ~new_P1_U3199;
  assign new_P1_R1165_U157 = ~new_P1_U3196;
  assign new_P1_R1165_U158 = ~new_P1_U3195;
  assign new_P1_R1165_U159 = ~new_P1_U3193;
  assign new_P1_R1165_U160 = ~new_P1_U3194;
  assign new_P1_R1165_U161 = ~new_P1_U3192;
  assign new_P1_R1165_U162 = ~new_P1_U3188;
  assign new_P1_R1165_U163 = ~new_P1_U3187;
  assign new_P1_R1165_U164 = ~new_P1_U3153;
  assign new_P1_R1165_U165 = ~new_P1_U3182;
  assign new_P1_R1165_U166 = new_P1_R1165_U493 & new_P1_R1165_U492;
  assign new_P1_R1165_U167 = ~new_P1_R1165_U53 | ~new_P1_R1165_U351 | ~new_P1_R1165_U302;
  assign new_P1_R1165_U168 = ~new_P1_R1165_U296 | ~new_P1_R1165_U295;
  assign new_P1_R1165_U169 = new_P1_R1165_U512 & new_P1_R1165_U511;
  assign new_P1_R1165_U170 = ~new_P1_R1165_U292 | ~new_P1_R1165_U291;
  assign new_P1_R1165_U171 = new_P1_R1165_U519 & new_P1_R1165_U518;
  assign new_P1_R1165_U172 = ~new_P1_R1165_U288 | ~new_P1_R1165_U287 | ~new_P1_R1165_U283;
  assign new_P1_R1165_U173 = new_P1_R1165_U533 & new_P1_R1165_U532;
  assign new_P1_R1165_U174 = ~new_P1_R1165_U195 | ~new_P1_R1165_U194;
  assign new_P1_R1165_U175 = ~new_P1_R1165_U278 | ~new_P1_R1165_U277;
  assign new_P1_R1165_U176 = new_P1_R1165_U545 & new_P1_R1165_U544;
  assign new_P1_R1165_U177 = ~new_P1_R1165_U118 | ~new_P1_R1165_U274;
  assign new_P1_R1165_U178 = new_P1_R1165_U559 & new_P1_R1165_U558;
  assign new_P1_R1165_U179 = ~new_P1_R1165_U262 | ~new_P1_R1165_U261;
  assign new_P1_R1165_U180 = new_P1_R1165_U566 & new_P1_R1165_U565;
  assign new_P1_R1165_U181 = ~new_P1_R1165_U258 | ~new_P1_R1165_U257;
  assign new_P1_R1165_U182 = ~new_P1_R1165_U248 | ~new_P1_R1165_U247;
  assign new_P1_R1165_U183 = new_P1_R1165_U585 & new_P1_R1165_U584;
  assign new_P1_R1165_U184 = ~new_P1_R1165_U244 | ~new_P1_R1165_U243;
  assign new_P1_R1165_U185 = ~new_P1_R1165_U353 | ~new_P1_R1165_U352;
  assign new_P1_R1165_U186 = ~new_P1_R1165_U20;
  assign new_P1_R1165_U187 = ~new_P1_U3169 | ~new_P1_R1165_U78;
  assign new_P1_R1165_U188 = ~new_P1_U3161 | ~new_P1_R1165_U83;
  assign new_P1_R1165_U189 = ~new_P1_U3156 | ~new_P1_R1165_U69;
  assign new_P1_R1165_U190 = ~new_P1_R1165_U43;
  assign new_P1_R1165_U191 = ~new_P1_R1165_U49;
  assign new_P1_R1165_U192 = ~new_P1_U3157 | ~new_P1_R1165_U71;
  assign new_P1_R1165_U193 = new_P1_U3211 | new_P1_U3181;
  assign new_P1_R1165_U194 = ~new_P1_R1165_U63 | ~new_P1_R1165_U193;
  assign new_P1_R1165_U195 = ~new_P1_U3181 | ~new_P1_U3211;
  assign new_P1_R1165_U196 = ~new_P1_R1165_U174;
  assign new_P1_R1165_U197 = ~new_P1_R1165_U371 | ~new_P1_R1165_U23;
  assign new_P1_R1165_U198 = ~new_P1_R1165_U197 | ~new_P1_R1165_U174;
  assign new_P1_R1165_U199 = ~new_P1_U3180 | ~new_P1_R1165_U64;
  assign new_P1_R1165_U200 = ~new_P1_R1165_U31;
  assign new_P1_R1165_U201 = ~new_P1_R1165_U374 | ~new_P1_R1165_U21;
  assign new_P1_R1165_U202 = ~new_P1_R1165_U377 | ~new_P1_R1165_U19;
  assign new_P1_R1165_U203 = ~new_P1_R1165_U21 | ~new_P1_R1165_U20;
  assign new_P1_R1165_U204 = ~new_P1_R1165_U62 | ~new_P1_R1165_U203;
  assign new_P1_R1165_U205 = ~new_P1_U3178 | ~new_P1_R1165_U186;
  assign new_P1_R1165_U206 = ~new_P1_R1165_U4 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U207 = ~new_P1_R1165_U24;
  assign new_P1_R1165_U208 = ~new_P1_R1165_U207 | ~new_P1_R1165_U25;
  assign new_P1_R1165_U209 = ~new_P1_R1165_U65 | ~new_P1_R1165_U208;
  assign new_P1_R1165_U210 = ~new_P1_U3177 | ~new_P1_R1165_U24;
  assign new_P1_R1165_U211 = ~new_P1_R1165_U144;
  assign new_P1_R1165_U212 = ~new_P1_R1165_U383 | ~new_P1_R1165_U26;
  assign new_P1_R1165_U213 = ~new_P1_R1165_U212 | ~new_P1_R1165_U144;
  assign new_P1_R1165_U214 = ~new_P1_U3176 | ~new_P1_R1165_U66;
  assign new_P1_R1165_U215 = ~new_P1_R1165_U30;
  assign new_P1_R1165_U216 = ~new_P1_R1165_U386 | ~new_P1_R1165_U18;
  assign new_P1_R1165_U217 = ~new_P1_R1165_U389 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U218 = ~new_P1_R1165_U17;
  assign new_P1_R1165_U219 = ~new_P1_R1165_U18 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U220 = ~new_P1_R1165_U60 | ~new_P1_R1165_U219;
  assign new_P1_R1165_U221 = ~new_P1_U3174 | ~new_P1_R1165_U218;
  assign new_P1_R1165_U222 = ~new_P1_R1165_U5 | ~new_P1_R1165_U30;
  assign new_P1_R1165_U223 = ~new_P1_R1165_U142;
  assign new_P1_R1165_U224 = ~new_P1_R1165_U392 | ~new_P1_R1165_U27;
  assign new_P1_R1165_U225 = ~new_P1_R1165_U224 | ~new_P1_R1165_U142;
  assign new_P1_R1165_U226 = ~new_P1_U3173 | ~new_P1_R1165_U67;
  assign new_P1_R1165_U227 = ~new_P1_R1165_U29;
  assign new_P1_R1165_U228 = ~new_P1_R1165_U389 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U229 = ~new_P1_R1165_U228 | ~new_P1_R1165_U30;
  assign new_P1_R1165_U230 = ~new_P1_R1165_U112 | ~new_P1_R1165_U229;
  assign new_P1_R1165_U231 = ~new_P1_R1165_U215 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U232 = ~new_P1_U3174 | ~new_P1_R1165_U60;
  assign new_P1_R1165_U233 = ~new_P1_R1165_U113 | ~new_P1_R1165_U231;
  assign new_P1_R1165_U234 = ~new_P1_R1165_U389 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U235 = ~new_P1_R1165_U377 | ~new_P1_R1165_U19;
  assign new_P1_R1165_U236 = ~new_P1_R1165_U235 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U237 = ~new_P1_R1165_U114 | ~new_P1_R1165_U236;
  assign new_P1_R1165_U238 = ~new_P1_R1165_U200 | ~new_P1_R1165_U20;
  assign new_P1_R1165_U239 = ~new_P1_U3178 | ~new_P1_R1165_U62;
  assign new_P1_R1165_U240 = ~new_P1_R1165_U115 | ~new_P1_R1165_U238;
  assign new_P1_R1165_U241 = ~new_P1_R1165_U377 | ~new_P1_R1165_U19;
  assign new_P1_R1165_U242 = ~new_P1_R1165_U227 | ~new_P1_R1165_U28;
  assign new_P1_R1165_U243 = ~new_P1_R1165_U58 | ~new_P1_R1165_U242;
  assign new_P1_R1165_U244 = ~new_P1_U3172 | ~new_P1_R1165_U29;
  assign new_P1_R1165_U245 = ~new_P1_R1165_U184;
  assign new_P1_R1165_U246 = ~new_P1_R1165_U453 | ~new_P1_R1165_U40;
  assign new_P1_R1165_U247 = ~new_P1_R1165_U246 | ~new_P1_R1165_U184;
  assign new_P1_R1165_U248 = ~new_P1_U3171 | ~new_P1_R1165_U75;
  assign new_P1_R1165_U249 = ~new_P1_R1165_U182;
  assign new_P1_R1165_U250 = ~new_P1_R1165_U456 | ~new_P1_R1165_U44;
  assign new_P1_R1165_U251 = ~new_P1_R1165_U459 | ~new_P1_R1165_U41;
  assign new_P1_R1165_U252 = ~new_P1_R1165_U190 | ~new_P1_R1165_U6;
  assign new_P1_R1165_U253 = ~new_P1_U3168 | ~new_P1_R1165_U77;
  assign new_P1_R1165_U254 = ~new_P1_R1165_U117 | ~new_P1_R1165_U252;
  assign new_P1_R1165_U255 = ~new_P1_R1165_U462 | ~new_P1_R1165_U42;
  assign new_P1_R1165_U256 = ~new_P1_R1165_U456 | ~new_P1_R1165_U44;
  assign new_P1_R1165_U257 = ~new_P1_R1165_U116 | ~new_P1_R1165_U182;
  assign new_P1_R1165_U258 = ~new_P1_R1165_U256 | ~new_P1_R1165_U254;
  assign new_P1_R1165_U259 = ~new_P1_R1165_U181;
  assign new_P1_R1165_U260 = ~new_P1_R1165_U465 | ~new_P1_R1165_U45;
  assign new_P1_R1165_U261 = ~new_P1_R1165_U260 | ~new_P1_R1165_U181;
  assign new_P1_R1165_U262 = ~new_P1_U3167 | ~new_P1_R1165_U79;
  assign new_P1_R1165_U263 = ~new_P1_R1165_U179;
  assign new_P1_R1165_U264 = ~new_P1_R1165_U468 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U265 = ~new_P1_R1165_U264 | ~new_P1_R1165_U179;
  assign new_P1_R1165_U266 = ~new_P1_U3166 | ~new_P1_R1165_U80;
  assign new_P1_R1165_U267 = ~new_P1_R1165_U56;
  assign new_P1_R1165_U268 = ~new_P1_R1165_U471 | ~new_P1_R1165_U39;
  assign new_P1_R1165_U269 = ~new_P1_R1165_U474 | ~new_P1_R1165_U37;
  assign new_P1_R1165_U270 = ~new_P1_R1165_U38;
  assign new_P1_R1165_U271 = ~new_P1_R1165_U39 | ~new_P1_R1165_U38;
  assign new_P1_R1165_U272 = ~new_P1_R1165_U74 | ~new_P1_R1165_U271;
  assign new_P1_R1165_U273 = ~new_P1_U3164 | ~new_P1_R1165_U270;
  assign new_P1_R1165_U274 = ~new_P1_R1165_U7 | ~new_P1_R1165_U56;
  assign new_P1_R1165_U275 = ~new_P1_R1165_U177;
  assign new_P1_R1165_U276 = ~new_P1_R1165_U477 | ~new_P1_R1165_U47;
  assign new_P1_R1165_U277 = ~new_P1_R1165_U276 | ~new_P1_R1165_U177;
  assign new_P1_R1165_U278 = ~new_P1_U3163 | ~new_P1_R1165_U81;
  assign new_P1_R1165_U279 = ~new_P1_R1165_U175;
  assign new_P1_R1165_U280 = ~new_P1_R1165_U444 | ~new_P1_R1165_U36;
  assign new_P1_R1165_U281 = ~new_P1_R1165_U447 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U282 = ~new_P1_R1165_U191 | ~new_P1_R1165_U8;
  assign new_P1_R1165_U283 = ~new_P1_U3160 | ~new_P1_R1165_U72;
  assign new_P1_R1165_U284 = ~new_P1_R1165_U188 | ~new_P1_R1165_U282;
  assign new_P1_R1165_U285 = ~new_P1_R1165_U450 | ~new_P1_R1165_U48;
  assign new_P1_R1165_U286 = ~new_P1_R1165_U444 | ~new_P1_R1165_U36;
  assign new_P1_R1165_U287 = ~new_P1_R1165_U8 | ~new_P1_R1165_U285 | ~new_P1_R1165_U175;
  assign new_P1_R1165_U288 = ~new_P1_R1165_U286 | ~new_P1_R1165_U284;
  assign new_P1_R1165_U289 = ~new_P1_R1165_U172;
  assign new_P1_R1165_U290 = ~new_P1_R1165_U480 | ~new_P1_R1165_U51;
  assign new_P1_R1165_U291 = ~new_P1_R1165_U290 | ~new_P1_R1165_U172;
  assign new_P1_R1165_U292 = ~new_P1_U3159 | ~new_P1_R1165_U84;
  assign new_P1_R1165_U293 = ~new_P1_R1165_U170;
  assign new_P1_R1165_U294 = ~new_P1_R1165_U483 | ~new_P1_R1165_U52;
  assign new_P1_R1165_U295 = ~new_P1_R1165_U294 | ~new_P1_R1165_U170;
  assign new_P1_R1165_U296 = ~new_P1_U3158 | ~new_P1_R1165_U85;
  assign new_P1_R1165_U297 = ~new_P1_R1165_U168;
  assign new_P1_R1165_U298 = ~new_P1_R1165_U435 | ~new_P1_R1165_U34;
  assign new_P1_R1165_U299 = ~new_P1_R1165_U192 | ~new_P1_R1165_U189;
  assign new_P1_R1165_U300 = ~new_P1_R1165_U53;
  assign new_P1_R1165_U301 = ~new_P1_R1165_U441 | ~new_P1_R1165_U35;
  assign new_P1_R1165_U302 = ~new_P1_R1165_U185 | ~new_P1_R1165_U168 | ~new_P1_R1165_U301;
  assign new_P1_R1165_U303 = ~new_P1_R1165_U167;
  assign new_P1_R1165_U304 = ~new_P1_R1165_U432 | ~new_P1_R1165_U32;
  assign new_P1_R1165_U305 = ~new_P1_U3154 | ~new_P1_R1165_U68;
  assign new_P1_R1165_U306 = ~new_P1_R1165_U432 | ~new_P1_R1165_U32;
  assign new_P1_R1165_U307 = ~new_P1_R1165_U301 | ~new_P1_R1165_U168;
  assign new_P1_R1165_U308 = ~new_P1_R1165_U54;
  assign new_P1_R1165_U309 = ~new_P1_R1165_U435 | ~new_P1_R1165_U34;
  assign new_P1_R1165_U310 = ~new_P1_R1165_U309 | ~new_P1_R1165_U54;
  assign new_P1_R1165_U311 = ~new_P1_R1165_U123 | ~new_P1_R1165_U310;
  assign new_P1_R1165_U312 = ~new_P1_R1165_U308 | ~new_P1_R1165_U189;
  assign new_P1_R1165_U313 = ~new_P1_U3155 | ~new_P1_R1165_U70;
  assign new_P1_R1165_U314 = ~new_P1_R1165_U185 | ~new_P1_R1165_U312 | ~new_P1_R1165_U313;
  assign new_P1_R1165_U315 = ~new_P1_R1165_U435 | ~new_P1_R1165_U34;
  assign new_P1_R1165_U316 = ~new_P1_R1165_U285 | ~new_P1_R1165_U175;
  assign new_P1_R1165_U317 = ~new_P1_R1165_U55;
  assign new_P1_R1165_U318 = ~new_P1_R1165_U447 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U319 = ~new_P1_R1165_U318 | ~new_P1_R1165_U55;
  assign new_P1_R1165_U320 = ~new_P1_R1165_U124 | ~new_P1_R1165_U319;
  assign new_P1_R1165_U321 = ~new_P1_R1165_U317 | ~new_P1_R1165_U188;
  assign new_P1_R1165_U322 = ~new_P1_U3160 | ~new_P1_R1165_U72;
  assign new_P1_R1165_U323 = ~new_P1_R1165_U8 | ~new_P1_R1165_U322 | ~new_P1_R1165_U321;
  assign new_P1_R1165_U324 = ~new_P1_R1165_U447 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U325 = ~new_P1_R1165_U474 | ~new_P1_R1165_U37;
  assign new_P1_R1165_U326 = ~new_P1_R1165_U325 | ~new_P1_R1165_U56;
  assign new_P1_R1165_U327 = ~new_P1_R1165_U125 | ~new_P1_R1165_U326;
  assign new_P1_R1165_U328 = ~new_P1_R1165_U267 | ~new_P1_R1165_U38;
  assign new_P1_R1165_U329 = ~new_P1_U3164 | ~new_P1_R1165_U74;
  assign new_P1_R1165_U330 = ~new_P1_R1165_U126 | ~new_P1_R1165_U328;
  assign new_P1_R1165_U331 = ~new_P1_R1165_U474 | ~new_P1_R1165_U37;
  assign new_P1_R1165_U332 = ~new_P1_R1165_U255 | ~new_P1_R1165_U182;
  assign new_P1_R1165_U333 = ~new_P1_R1165_U57;
  assign new_P1_R1165_U334 = ~new_P1_R1165_U459 | ~new_P1_R1165_U41;
  assign new_P1_R1165_U335 = ~new_P1_R1165_U334 | ~new_P1_R1165_U57;
  assign new_P1_R1165_U336 = ~new_P1_R1165_U127 | ~new_P1_R1165_U335;
  assign new_P1_R1165_U337 = ~new_P1_R1165_U333 | ~new_P1_R1165_U187;
  assign new_P1_R1165_U338 = ~new_P1_U3168 | ~new_P1_R1165_U77;
  assign new_P1_R1165_U339 = ~new_P1_R1165_U128 | ~new_P1_R1165_U337;
  assign new_P1_R1165_U340 = ~new_P1_R1165_U459 | ~new_P1_R1165_U41;
  assign new_P1_R1165_U341 = ~new_P1_R1165_U234 | ~new_P1_R1165_U17;
  assign new_P1_R1165_U342 = ~new_P1_R1165_U241 | ~new_P1_R1165_U20;
  assign new_P1_R1165_U343 = ~new_P1_R1165_U315 | ~new_P1_R1165_U189;
  assign new_P1_R1165_U344 = ~new_P1_R1165_U301 | ~new_P1_R1165_U192;
  assign new_P1_R1165_U345 = ~new_P1_R1165_U324 | ~new_P1_R1165_U188;
  assign new_P1_R1165_U346 = ~new_P1_R1165_U285 | ~new_P1_R1165_U49;
  assign new_P1_R1165_U347 = ~new_P1_R1165_U331 | ~new_P1_R1165_U38;
  assign new_P1_R1165_U348 = ~new_P1_R1165_U340 | ~new_P1_R1165_U187;
  assign new_P1_R1165_U349 = ~new_P1_R1165_U255 | ~new_P1_R1165_U43;
  assign new_P1_R1165_U350 = ~new_P1_R1165_U119 | ~new_P1_R1165_U351 | ~new_P1_R1165_U302;
  assign new_P1_R1165_U351 = ~new_P1_R1165_U299 | ~new_P1_R1165_U185;
  assign new_P1_R1165_U352 = ~new_P1_R1165_U70 | ~new_P1_R1165_U298;
  assign new_P1_R1165_U353 = ~new_P1_U3155 | ~new_P1_R1165_U298;
  assign new_P1_R1165_U354 = ~new_P1_R1165_U306 | ~new_P1_R1165_U299 | ~new_P1_R1165_U185;
  assign new_P1_R1165_U355 = ~new_P1_R1165_U120 | ~new_P1_R1165_U168 | ~new_P1_R1165_U185;
  assign new_P1_R1165_U356 = ~new_P1_R1165_U300 | ~new_P1_R1165_U306;
  assign new_P1_R1165_U357 = ~new_P1_U3154 | ~new_P1_R1165_U68;
  assign new_P1_R1165_U358 = ~new_P1_U3211 | ~new_P1_R1165_U130;
  assign new_P1_R1165_U359 = ~new_P1_U3201 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U360 = ~new_P1_R1165_U58;
  assign new_P1_R1165_U361 = ~new_P1_R1165_U360 | ~new_P1_U3172;
  assign new_P1_R1165_U362 = ~new_P1_R1165_U58 | ~new_P1_R1165_U28;
  assign new_P1_R1165_U363 = ~new_P1_R1165_U360 | ~new_P1_U3172;
  assign new_P1_R1165_U364 = ~new_P1_R1165_U58 | ~new_P1_R1165_U28;
  assign new_P1_R1165_U365 = ~new_P1_R1165_U364 | ~new_P1_R1165_U363;
  assign new_P1_R1165_U366 = ~new_P1_U3211 | ~new_P1_R1165_U132;
  assign new_P1_R1165_U367 = ~new_P1_U3210 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U368 = ~new_P1_R1165_U63;
  assign new_P1_R1165_U369 = ~new_P1_U3211 | ~new_P1_R1165_U133;
  assign new_P1_R1165_U370 = ~new_P1_U3209 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U371 = ~new_P1_R1165_U64;
  assign new_P1_R1165_U372 = ~new_P1_U3211 | ~new_P1_R1165_U134;
  assign new_P1_R1165_U373 = ~new_P1_U3207 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U374 = ~new_P1_R1165_U62;
  assign new_P1_R1165_U375 = ~new_P1_U3211 | ~new_P1_R1165_U135;
  assign new_P1_R1165_U376 = ~new_P1_U3208 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U377 = ~new_P1_R1165_U61;
  assign new_P1_R1165_U378 = ~new_P1_U3211 | ~new_P1_R1165_U136;
  assign new_P1_R1165_U379 = ~new_P1_U3206 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U380 = ~new_P1_R1165_U65;
  assign new_P1_R1165_U381 = ~new_P1_U3211 | ~new_P1_R1165_U137;
  assign new_P1_R1165_U382 = ~new_P1_U3205 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U383 = ~new_P1_R1165_U66;
  assign new_P1_R1165_U384 = ~new_P1_U3211 | ~new_P1_R1165_U138;
  assign new_P1_R1165_U385 = ~new_P1_U3203 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U386 = ~new_P1_R1165_U60;
  assign new_P1_R1165_U387 = ~new_P1_U3211 | ~new_P1_R1165_U139;
  assign new_P1_R1165_U388 = ~new_P1_U3204 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U389 = ~new_P1_R1165_U59;
  assign new_P1_R1165_U390 = ~new_P1_U3211 | ~new_P1_R1165_U140;
  assign new_P1_R1165_U391 = ~new_P1_U3202 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U392 = ~new_P1_R1165_U67;
  assign new_P1_R1165_U393 = ~new_P1_R1165_U131 | ~new_P1_R1165_U29;
  assign new_P1_R1165_U394 = ~new_P1_R1165_U365 | ~new_P1_R1165_U227;
  assign new_P1_R1165_U395 = ~new_P1_R1165_U392 | ~new_P1_U3173;
  assign new_P1_R1165_U396 = ~new_P1_R1165_U67 | ~new_P1_R1165_U27;
  assign new_P1_R1165_U397 = ~new_P1_R1165_U392 | ~new_P1_U3173;
  assign new_P1_R1165_U398 = ~new_P1_R1165_U67 | ~new_P1_R1165_U27;
  assign new_P1_R1165_U399 = ~new_P1_R1165_U398 | ~new_P1_R1165_U397;
  assign new_P1_R1165_U400 = ~new_P1_R1165_U141 | ~new_P1_R1165_U142;
  assign new_P1_R1165_U401 = ~new_P1_R1165_U223 | ~new_P1_R1165_U399;
  assign new_P1_R1165_U402 = ~new_P1_R1165_U386 | ~new_P1_U3174;
  assign new_P1_R1165_U403 = ~new_P1_R1165_U60 | ~new_P1_R1165_U18;
  assign new_P1_R1165_U404 = ~new_P1_R1165_U389 | ~new_P1_U3175;
  assign new_P1_R1165_U405 = ~new_P1_R1165_U59 | ~new_P1_R1165_U16;
  assign new_P1_R1165_U406 = ~new_P1_R1165_U405 | ~new_P1_R1165_U404;
  assign new_P1_R1165_U407 = ~new_P1_R1165_U341 | ~new_P1_R1165_U30;
  assign new_P1_R1165_U408 = ~new_P1_R1165_U406 | ~new_P1_R1165_U215;
  assign new_P1_R1165_U409 = ~new_P1_R1165_U383 | ~new_P1_U3176;
  assign new_P1_R1165_U410 = ~new_P1_R1165_U66 | ~new_P1_R1165_U26;
  assign new_P1_R1165_U411 = ~new_P1_R1165_U383 | ~new_P1_U3176;
  assign new_P1_R1165_U412 = ~new_P1_R1165_U66 | ~new_P1_R1165_U26;
  assign new_P1_R1165_U413 = ~new_P1_R1165_U412 | ~new_P1_R1165_U411;
  assign new_P1_R1165_U414 = ~new_P1_R1165_U143 | ~new_P1_R1165_U144;
  assign new_P1_R1165_U415 = ~new_P1_R1165_U211 | ~new_P1_R1165_U413;
  assign new_P1_R1165_U416 = ~new_P1_R1165_U380 | ~new_P1_U3177;
  assign new_P1_R1165_U417 = ~new_P1_R1165_U65 | ~new_P1_R1165_U25;
  assign new_P1_R1165_U418 = ~new_P1_R1165_U380 | ~new_P1_U3177;
  assign new_P1_R1165_U419 = ~new_P1_R1165_U65 | ~new_P1_R1165_U25;
  assign new_P1_R1165_U420 = ~new_P1_R1165_U419 | ~new_P1_R1165_U418;
  assign new_P1_R1165_U421 = ~new_P1_R1165_U145 | ~new_P1_R1165_U24;
  assign new_P1_R1165_U422 = ~new_P1_R1165_U420 | ~new_P1_R1165_U207;
  assign new_P1_R1165_U423 = ~new_P1_R1165_U374 | ~new_P1_U3178;
  assign new_P1_R1165_U424 = ~new_P1_R1165_U62 | ~new_P1_R1165_U21;
  assign new_P1_R1165_U425 = ~new_P1_R1165_U377 | ~new_P1_U3179;
  assign new_P1_R1165_U426 = ~new_P1_R1165_U61 | ~new_P1_R1165_U19;
  assign new_P1_R1165_U427 = ~new_P1_R1165_U426 | ~new_P1_R1165_U425;
  assign new_P1_R1165_U428 = ~new_P1_R1165_U342 | ~new_P1_R1165_U31;
  assign new_P1_R1165_U429 = ~new_P1_R1165_U427 | ~new_P1_R1165_U200;
  assign new_P1_R1165_U430 = ~new_P1_U3211 | ~new_P1_R1165_U146;
  assign new_P1_R1165_U431 = ~new_P1_U3183 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U432 = ~new_P1_R1165_U68;
  assign new_P1_R1165_U433 = ~new_P1_U3211 | ~new_P1_R1165_U147;
  assign new_P1_R1165_U434 = ~new_P1_U3185 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U435 = ~new_P1_R1165_U69;
  assign new_P1_R1165_U436 = ~new_P1_U3211 | ~new_P1_R1165_U148;
  assign new_P1_R1165_U437 = ~new_P1_U3184 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U438 = ~new_P1_R1165_U70;
  assign new_P1_R1165_U439 = ~new_P1_U3211 | ~new_P1_R1165_U149;
  assign new_P1_R1165_U440 = ~new_P1_U3186 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U441 = ~new_P1_R1165_U71;
  assign new_P1_R1165_U442 = ~new_P1_U3211 | ~new_P1_R1165_U150;
  assign new_P1_R1165_U443 = ~new_P1_U3189 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U444 = ~new_P1_R1165_U72;
  assign new_P1_R1165_U445 = ~new_P1_U3211 | ~new_P1_R1165_U151;
  assign new_P1_R1165_U446 = ~new_P1_U3190 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U447 = ~new_P1_R1165_U83;
  assign new_P1_R1165_U448 = ~new_P1_U3211 | ~new_P1_R1165_U152;
  assign new_P1_R1165_U449 = ~new_P1_U3191 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U450 = ~new_P1_R1165_U82;
  assign new_P1_R1165_U451 = ~new_P1_U3211 | ~new_P1_R1165_U153;
  assign new_P1_R1165_U452 = ~new_P1_U3200 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U453 = ~new_P1_R1165_U75;
  assign new_P1_R1165_U454 = ~new_P1_U3211 | ~new_P1_R1165_U154;
  assign new_P1_R1165_U455 = ~new_P1_U3197 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U456 = ~new_P1_R1165_U77;
  assign new_P1_R1165_U457 = ~new_P1_U3211 | ~new_P1_R1165_U155;
  assign new_P1_R1165_U458 = ~new_P1_U3198 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U459 = ~new_P1_R1165_U78;
  assign new_P1_R1165_U460 = ~new_P1_U3211 | ~new_P1_R1165_U156;
  assign new_P1_R1165_U461 = ~new_P1_U3199 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U462 = ~new_P1_R1165_U76;
  assign new_P1_R1165_U463 = ~new_P1_U3211 | ~new_P1_R1165_U157;
  assign new_P1_R1165_U464 = ~new_P1_U3196 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U465 = ~new_P1_R1165_U79;
  assign new_P1_R1165_U466 = ~new_P1_U3211 | ~new_P1_R1165_U158;
  assign new_P1_R1165_U467 = ~new_P1_U3195 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U468 = ~new_P1_R1165_U80;
  assign new_P1_R1165_U469 = ~new_P1_U3211 | ~new_P1_R1165_U159;
  assign new_P1_R1165_U470 = ~new_P1_U3193 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U471 = ~new_P1_R1165_U74;
  assign new_P1_R1165_U472 = ~new_P1_U3211 | ~new_P1_R1165_U160;
  assign new_P1_R1165_U473 = ~new_P1_U3194 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U474 = ~new_P1_R1165_U73;
  assign new_P1_R1165_U475 = ~new_P1_U3211 | ~new_P1_R1165_U161;
  assign new_P1_R1165_U476 = ~new_P1_U3192 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U477 = ~new_P1_R1165_U81;
  assign new_P1_R1165_U478 = ~new_P1_U3211 | ~new_P1_R1165_U162;
  assign new_P1_R1165_U479 = ~new_P1_U3188 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U480 = ~new_P1_R1165_U84;
  assign new_P1_R1165_U481 = ~new_P1_U3211 | ~new_P1_R1165_U163;
  assign new_P1_R1165_U482 = ~new_P1_U3187 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U483 = ~new_P1_R1165_U85;
  assign new_P1_R1165_U484 = ~new_P1_U3211 | ~new_P1_R1165_U164;
  assign new_P1_R1165_U485 = ~new_P1_U3153 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U486 = ~new_P1_R1165_U122;
  assign new_P1_R1165_U487 = ~new_P1_U3182 | ~new_P1_R1165_U486;
  assign new_P1_R1165_U488 = ~new_P1_R1165_U122 | ~new_P1_R1165_U165;
  assign new_P1_R1165_U489 = ~new_P1_R1165_U86;
  assign new_P1_R1165_U490 = ~new_P1_R1165_U489 | ~new_P1_R1165_U350 | ~new_P1_R1165_U304;
  assign new_P1_R1165_U491 = ~new_P1_R1165_U86 | ~new_P1_R1165_U121 | ~new_P1_R1165_U356 | ~new_P1_R1165_U355;
  assign new_P1_R1165_U492 = ~new_P1_R1165_U432 | ~new_P1_U3154;
  assign new_P1_R1165_U493 = ~new_P1_R1165_U68 | ~new_P1_R1165_U32;
  assign new_P1_R1165_U494 = ~new_P1_R1165_U432 | ~new_P1_U3154;
  assign new_P1_R1165_U495 = ~new_P1_R1165_U68 | ~new_P1_R1165_U32;
  assign new_P1_R1165_U496 = ~new_P1_R1165_U495 | ~new_P1_R1165_U494;
  assign new_P1_R1165_U497 = ~new_P1_R1165_U166 | ~new_P1_R1165_U167;
  assign new_P1_R1165_U498 = ~new_P1_R1165_U303 | ~new_P1_R1165_U496;
  assign new_P1_R1165_U499 = ~new_P1_R1165_U438 | ~new_P1_U3155;
  assign new_P1_R1165_U500 = ~new_P1_R1165_U70 | ~new_P1_R1165_U33;
  assign new_P1_R1165_U501 = ~new_P1_R1165_U435 | ~new_P1_U3156;
  assign new_P1_R1165_U502 = ~new_P1_R1165_U69 | ~new_P1_R1165_U34;
  assign new_P1_R1165_U503 = ~new_P1_R1165_U502 | ~new_P1_R1165_U501;
  assign new_P1_R1165_U504 = ~new_P1_R1165_U343 | ~new_P1_R1165_U54;
  assign new_P1_R1165_U505 = ~new_P1_R1165_U503 | ~new_P1_R1165_U308;
  assign new_P1_R1165_U506 = ~new_P1_R1165_U441 | ~new_P1_U3157;
  assign new_P1_R1165_U507 = ~new_P1_R1165_U71 | ~new_P1_R1165_U35;
  assign new_P1_R1165_U508 = ~new_P1_R1165_U507 | ~new_P1_R1165_U506;
  assign new_P1_R1165_U509 = ~new_P1_R1165_U344 | ~new_P1_R1165_U168;
  assign new_P1_R1165_U510 = ~new_P1_R1165_U297 | ~new_P1_R1165_U508;
  assign new_P1_R1165_U511 = ~new_P1_R1165_U483 | ~new_P1_U3158;
  assign new_P1_R1165_U512 = ~new_P1_R1165_U85 | ~new_P1_R1165_U52;
  assign new_P1_R1165_U513 = ~new_P1_R1165_U483 | ~new_P1_U3158;
  assign new_P1_R1165_U514 = ~new_P1_R1165_U85 | ~new_P1_R1165_U52;
  assign new_P1_R1165_U515 = ~new_P1_R1165_U514 | ~new_P1_R1165_U513;
  assign new_P1_R1165_U516 = ~new_P1_R1165_U169 | ~new_P1_R1165_U170;
  assign new_P1_R1165_U517 = ~new_P1_R1165_U293 | ~new_P1_R1165_U515;
  assign new_P1_R1165_U518 = ~new_P1_R1165_U480 | ~new_P1_U3159;
  assign new_P1_R1165_U519 = ~new_P1_R1165_U84 | ~new_P1_R1165_U51;
  assign new_P1_R1165_U520 = ~new_P1_R1165_U480 | ~new_P1_U3159;
  assign new_P1_R1165_U521 = ~new_P1_R1165_U84 | ~new_P1_R1165_U51;
  assign new_P1_R1165_U522 = ~new_P1_R1165_U521 | ~new_P1_R1165_U520;
  assign new_P1_R1165_U523 = ~new_P1_R1165_U171 | ~new_P1_R1165_U172;
  assign new_P1_R1165_U524 = ~new_P1_R1165_U289 | ~new_P1_R1165_U522;
  assign new_P1_R1165_U525 = ~new_P1_R1165_U444 | ~new_P1_U3160;
  assign new_P1_R1165_U526 = ~new_P1_R1165_U72 | ~new_P1_R1165_U36;
  assign new_P1_R1165_U527 = ~new_P1_R1165_U447 | ~new_P1_U3161;
  assign new_P1_R1165_U528 = ~new_P1_R1165_U83 | ~new_P1_R1165_U50;
  assign new_P1_R1165_U529 = ~new_P1_R1165_U528 | ~new_P1_R1165_U527;
  assign new_P1_R1165_U530 = ~new_P1_R1165_U345 | ~new_P1_R1165_U55;
  assign new_P1_R1165_U531 = ~new_P1_R1165_U529 | ~new_P1_R1165_U317;
  assign new_P1_R1165_U532 = ~new_P1_R1165_U371 | ~new_P1_U3180;
  assign new_P1_R1165_U533 = ~new_P1_R1165_U64 | ~new_P1_R1165_U23;
  assign new_P1_R1165_U534 = ~new_P1_R1165_U371 | ~new_P1_U3180;
  assign new_P1_R1165_U535 = ~new_P1_R1165_U64 | ~new_P1_R1165_U23;
  assign new_P1_R1165_U536 = ~new_P1_R1165_U535 | ~new_P1_R1165_U534;
  assign new_P1_R1165_U537 = ~new_P1_R1165_U173 | ~new_P1_R1165_U174;
  assign new_P1_R1165_U538 = ~new_P1_R1165_U196 | ~new_P1_R1165_U536;
  assign new_P1_R1165_U539 = ~new_P1_R1165_U450 | ~new_P1_U3162;
  assign new_P1_R1165_U540 = ~new_P1_R1165_U82 | ~new_P1_R1165_U48;
  assign new_P1_R1165_U541 = ~new_P1_R1165_U540 | ~new_P1_R1165_U539;
  assign new_P1_R1165_U542 = ~new_P1_R1165_U346 | ~new_P1_R1165_U175;
  assign new_P1_R1165_U543 = ~new_P1_R1165_U279 | ~new_P1_R1165_U541;
  assign new_P1_R1165_U544 = ~new_P1_R1165_U477 | ~new_P1_U3163;
  assign new_P1_R1165_U545 = ~new_P1_R1165_U81 | ~new_P1_R1165_U47;
  assign new_P1_R1165_U546 = ~new_P1_R1165_U477 | ~new_P1_U3163;
  assign new_P1_R1165_U547 = ~new_P1_R1165_U81 | ~new_P1_R1165_U47;
  assign new_P1_R1165_U548 = ~new_P1_R1165_U547 | ~new_P1_R1165_U546;
  assign new_P1_R1165_U549 = ~new_P1_R1165_U176 | ~new_P1_R1165_U177;
  assign new_P1_R1165_U550 = ~new_P1_R1165_U275 | ~new_P1_R1165_U548;
  assign new_P1_R1165_U551 = ~new_P1_R1165_U471 | ~new_P1_U3164;
  assign new_P1_R1165_U552 = ~new_P1_R1165_U74 | ~new_P1_R1165_U39;
  assign new_P1_R1165_U553 = ~new_P1_R1165_U474 | ~new_P1_U3165;
  assign new_P1_R1165_U554 = ~new_P1_R1165_U73 | ~new_P1_R1165_U37;
  assign new_P1_R1165_U555 = ~new_P1_R1165_U554 | ~new_P1_R1165_U553;
  assign new_P1_R1165_U556 = ~new_P1_R1165_U347 | ~new_P1_R1165_U56;
  assign new_P1_R1165_U557 = ~new_P1_R1165_U555 | ~new_P1_R1165_U267;
  assign new_P1_R1165_U558 = ~new_P1_R1165_U468 | ~new_P1_U3166;
  assign new_P1_R1165_U559 = ~new_P1_R1165_U80 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U560 = ~new_P1_R1165_U468 | ~new_P1_U3166;
  assign new_P1_R1165_U561 = ~new_P1_R1165_U80 | ~new_P1_R1165_U46;
  assign new_P1_R1165_U562 = ~new_P1_R1165_U561 | ~new_P1_R1165_U560;
  assign new_P1_R1165_U563 = ~new_P1_R1165_U178 | ~new_P1_R1165_U179;
  assign new_P1_R1165_U564 = ~new_P1_R1165_U263 | ~new_P1_R1165_U562;
  assign new_P1_R1165_U565 = ~new_P1_R1165_U465 | ~new_P1_U3167;
  assign new_P1_R1165_U566 = ~new_P1_R1165_U79 | ~new_P1_R1165_U45;
  assign new_P1_R1165_U567 = ~new_P1_R1165_U465 | ~new_P1_U3167;
  assign new_P1_R1165_U568 = ~new_P1_R1165_U79 | ~new_P1_R1165_U45;
  assign new_P1_R1165_U569 = ~new_P1_R1165_U568 | ~new_P1_R1165_U567;
  assign new_P1_R1165_U570 = ~new_P1_R1165_U180 | ~new_P1_R1165_U181;
  assign new_P1_R1165_U571 = ~new_P1_R1165_U259 | ~new_P1_R1165_U569;
  assign new_P1_R1165_U572 = ~new_P1_R1165_U456 | ~new_P1_U3168;
  assign new_P1_R1165_U573 = ~new_P1_R1165_U77 | ~new_P1_R1165_U44;
  assign new_P1_R1165_U574 = ~new_P1_R1165_U459 | ~new_P1_U3169;
  assign new_P1_R1165_U575 = ~new_P1_R1165_U78 | ~new_P1_R1165_U41;
  assign new_P1_R1165_U576 = ~new_P1_R1165_U575 | ~new_P1_R1165_U574;
  assign new_P1_R1165_U577 = ~new_P1_R1165_U348 | ~new_P1_R1165_U57;
  assign new_P1_R1165_U578 = ~new_P1_R1165_U576 | ~new_P1_R1165_U333;
  assign new_P1_R1165_U579 = ~new_P1_R1165_U462 | ~new_P1_U3170;
  assign new_P1_R1165_U580 = ~new_P1_R1165_U76 | ~new_P1_R1165_U42;
  assign new_P1_R1165_U581 = ~new_P1_R1165_U580 | ~new_P1_R1165_U579;
  assign new_P1_R1165_U582 = ~new_P1_R1165_U349 | ~new_P1_R1165_U182;
  assign new_P1_R1165_U583 = ~new_P1_R1165_U249 | ~new_P1_R1165_U581;
  assign new_P1_R1165_U584 = ~new_P1_R1165_U453 | ~new_P1_U3171;
  assign new_P1_R1165_U585 = ~new_P1_R1165_U75 | ~new_P1_R1165_U40;
  assign new_P1_R1165_U586 = ~new_P1_R1165_U453 | ~new_P1_U3171;
  assign new_P1_R1165_U587 = ~new_P1_R1165_U75 | ~new_P1_R1165_U40;
  assign new_P1_R1165_U588 = ~new_P1_R1165_U587 | ~new_P1_R1165_U586;
  assign new_P1_R1165_U589 = ~new_P1_R1165_U183 | ~new_P1_R1165_U184;
  assign new_P1_R1165_U590 = ~new_P1_R1165_U245 | ~new_P1_R1165_U588;
  assign new_P1_R1165_U591 = ~new_P1_U3181 | ~new_P1_R1165_U15;
  assign new_P1_R1165_U592 = ~new_P1_U3211 | ~new_P1_R1165_U22;
  assign new_P1_R1165_U593 = ~new_P1_R1165_U129;
  assign new_P1_R1165_U594 = ~new_P1_R1165_U63 | ~new_P1_R1165_U593;
  assign new_P1_R1165_U595 = ~new_P1_R1165_U129 | ~new_P1_R1165_U368;
  assign new_P1_R1150_U6 = new_P1_R1150_U184 & new_P1_R1150_U201;
  assign new_P1_R1150_U7 = new_P1_R1150_U203 & new_P1_R1150_U202;
  assign new_P1_R1150_U8 = new_P1_R1150_U179 & new_P1_R1150_U240;
  assign new_P1_R1150_U9 = new_P1_R1150_U242 & new_P1_R1150_U241;
  assign new_P1_R1150_U10 = new_P1_R1150_U259 & new_P1_R1150_U258;
  assign new_P1_R1150_U11 = new_P1_R1150_U285 & new_P1_R1150_U284;
  assign new_P1_R1150_U12 = new_P1_R1150_U383 & new_P1_R1150_U382;
  assign new_P1_R1150_U13 = ~new_P1_R1150_U340 | ~new_P1_R1150_U343;
  assign new_P1_R1150_U14 = ~new_P1_R1150_U329 | ~new_P1_R1150_U332;
  assign new_P1_R1150_U15 = ~new_P1_R1150_U318 | ~new_P1_R1150_U321;
  assign new_P1_R1150_U16 = ~new_P1_R1150_U310 | ~new_P1_R1150_U312;
  assign new_P1_R1150_U17 = ~new_P1_R1150_U348 | ~new_P1_R1150_U156 | ~new_P1_R1150_U175;
  assign new_P1_R1150_U18 = ~new_P1_R1150_U236 | ~new_P1_R1150_U238;
  assign new_P1_R1150_U19 = ~new_P1_R1150_U228 | ~new_P1_R1150_U231;
  assign new_P1_R1150_U20 = ~new_P1_R1150_U220 | ~new_P1_R1150_U222;
  assign new_P1_R1150_U21 = ~new_P1_R1150_U25 | ~new_P1_R1150_U346;
  assign new_P1_R1150_U22 = ~new_P1_U3479;
  assign new_P1_R1150_U23 = ~new_P1_U3464;
  assign new_P1_R1150_U24 = ~new_P1_U3456;
  assign new_P1_R1150_U25 = ~new_P1_U3456 | ~new_P1_R1150_U93;
  assign new_P1_R1150_U26 = ~new_P1_U3078;
  assign new_P1_R1150_U27 = ~new_P1_U3467;
  assign new_P1_R1150_U28 = ~new_P1_U3068;
  assign new_P1_R1150_U29 = ~new_P1_U3068 | ~new_P1_R1150_U23;
  assign new_P1_R1150_U30 = ~new_P1_U3064;
  assign new_P1_R1150_U31 = ~new_P1_U3476;
  assign new_P1_R1150_U32 = ~new_P1_U3473;
  assign new_P1_R1150_U33 = ~new_P1_U3470;
  assign new_P1_R1150_U34 = ~new_P1_U3071;
  assign new_P1_R1150_U35 = ~new_P1_U3067;
  assign new_P1_R1150_U36 = ~new_P1_U3060;
  assign new_P1_R1150_U37 = ~new_P1_U3060 | ~new_P1_R1150_U33;
  assign new_P1_R1150_U38 = ~new_P1_U3482;
  assign new_P1_R1150_U39 = ~new_P1_U3070;
  assign new_P1_R1150_U40 = ~new_P1_U3070 | ~new_P1_R1150_U22;
  assign new_P1_R1150_U41 = ~new_P1_U3084;
  assign new_P1_R1150_U42 = ~new_P1_U3485;
  assign new_P1_R1150_U43 = ~new_P1_U3083;
  assign new_P1_R1150_U44 = ~new_P1_R1150_U209 | ~new_P1_R1150_U208;
  assign new_P1_R1150_U45 = ~new_P1_R1150_U37 | ~new_P1_R1150_U224;
  assign new_P1_R1150_U46 = ~new_P1_R1150_U193 | ~new_P1_R1150_U192;
  assign new_P1_R1150_U47 = ~new_P1_U4019;
  assign new_P1_R1150_U48 = ~new_P1_U4023;
  assign new_P1_R1150_U49 = ~new_P1_U3503;
  assign new_P1_R1150_U50 = ~new_P1_U3491;
  assign new_P1_R1150_U51 = ~new_P1_U3488;
  assign new_P1_R1150_U52 = ~new_P1_U3063;
  assign new_P1_R1150_U53 = ~new_P1_U3062;
  assign new_P1_R1150_U54 = ~new_P1_U3083 | ~new_P1_R1150_U42;
  assign new_P1_R1150_U55 = ~new_P1_U3494;
  assign new_P1_R1150_U56 = ~new_P1_U3072;
  assign new_P1_R1150_U57 = ~new_P1_U3497;
  assign new_P1_R1150_U58 = ~new_P1_U3080;
  assign new_P1_R1150_U59 = ~new_P1_U3506;
  assign new_P1_R1150_U60 = ~new_P1_U3500;
  assign new_P1_R1150_U61 = ~new_P1_U3073;
  assign new_P1_R1150_U62 = ~new_P1_U3074;
  assign new_P1_R1150_U63 = ~new_P1_U3079;
  assign new_P1_R1150_U64 = ~new_P1_U3079 | ~new_P1_R1150_U60;
  assign new_P1_R1150_U65 = ~new_P1_U3509;
  assign new_P1_R1150_U66 = ~new_P1_U3069;
  assign new_P1_R1150_U67 = ~new_P1_R1150_U269 | ~new_P1_R1150_U268;
  assign new_P1_R1150_U68 = ~new_P1_U3082;
  assign new_P1_R1150_U69 = ~new_P1_U3514;
  assign new_P1_R1150_U70 = ~new_P1_U3081;
  assign new_P1_R1150_U71 = ~new_P1_U4025;
  assign new_P1_R1150_U72 = ~new_P1_U3076;
  assign new_P1_R1150_U73 = ~new_P1_U4022;
  assign new_P1_R1150_U74 = ~new_P1_U4024;
  assign new_P1_R1150_U75 = ~new_P1_U3066;
  assign new_P1_R1150_U76 = ~new_P1_U3061;
  assign new_P1_R1150_U77 = ~new_P1_U3075;
  assign new_P1_R1150_U78 = ~new_P1_U3075 | ~new_P1_R1150_U74;
  assign new_P1_R1150_U79 = ~new_P1_U4021;
  assign new_P1_R1150_U80 = ~new_P1_U3065;
  assign new_P1_R1150_U81 = ~new_P1_U4020;
  assign new_P1_R1150_U82 = ~new_P1_U3058;
  assign new_P1_R1150_U83 = ~new_P1_U4018;
  assign new_P1_R1150_U84 = ~new_P1_U3057;
  assign new_P1_R1150_U85 = ~new_P1_U3057 | ~new_P1_R1150_U47;
  assign new_P1_R1150_U86 = ~new_P1_U3053;
  assign new_P1_R1150_U87 = ~new_P1_U4017;
  assign new_P1_R1150_U88 = ~new_P1_U3054;
  assign new_P1_R1150_U89 = ~new_P1_R1150_U299 | ~new_P1_R1150_U298;
  assign new_P1_R1150_U90 = ~new_P1_R1150_U78 | ~new_P1_R1150_U314;
  assign new_P1_R1150_U91 = ~new_P1_R1150_U64 | ~new_P1_R1150_U325;
  assign new_P1_R1150_U92 = ~new_P1_R1150_U54 | ~new_P1_R1150_U336;
  assign new_P1_R1150_U93 = ~new_P1_U3077;
  assign new_P1_R1150_U94 = ~new_P1_R1150_U393 | ~new_P1_R1150_U392;
  assign new_P1_R1150_U95 = ~new_P1_R1150_U407 | ~new_P1_R1150_U406;
  assign new_P1_R1150_U96 = ~new_P1_R1150_U412 | ~new_P1_R1150_U411;
  assign new_P1_R1150_U97 = ~new_P1_R1150_U428 | ~new_P1_R1150_U427;
  assign new_P1_R1150_U98 = ~new_P1_R1150_U433 | ~new_P1_R1150_U432;
  assign new_P1_R1150_U99 = ~new_P1_R1150_U438 | ~new_P1_R1150_U437;
  assign new_P1_R1150_U100 = ~new_P1_R1150_U443 | ~new_P1_R1150_U442;
  assign new_P1_R1150_U101 = ~new_P1_R1150_U448 | ~new_P1_R1150_U447;
  assign new_P1_R1150_U102 = ~new_P1_R1150_U464 | ~new_P1_R1150_U463;
  assign new_P1_R1150_U103 = ~new_P1_R1150_U469 | ~new_P1_R1150_U468;
  assign new_P1_R1150_U104 = ~new_P1_R1150_U352 | ~new_P1_R1150_U351;
  assign new_P1_R1150_U105 = ~new_P1_R1150_U361 | ~new_P1_R1150_U360;
  assign new_P1_R1150_U106 = ~new_P1_R1150_U368 | ~new_P1_R1150_U367;
  assign new_P1_R1150_U107 = ~new_P1_R1150_U372 | ~new_P1_R1150_U371;
  assign new_P1_R1150_U108 = ~new_P1_R1150_U381 | ~new_P1_R1150_U380;
  assign new_P1_R1150_U109 = ~new_P1_R1150_U402 | ~new_P1_R1150_U401;
  assign new_P1_R1150_U110 = ~new_P1_R1150_U419 | ~new_P1_R1150_U418;
  assign new_P1_R1150_U111 = ~new_P1_R1150_U423 | ~new_P1_R1150_U422;
  assign new_P1_R1150_U112 = ~new_P1_R1150_U455 | ~new_P1_R1150_U454;
  assign new_P1_R1150_U113 = ~new_P1_R1150_U459 | ~new_P1_R1150_U458;
  assign new_P1_R1150_U114 = ~new_P1_R1150_U476 | ~new_P1_R1150_U475;
  assign new_P1_R1150_U115 = new_P1_R1150_U195 & new_P1_R1150_U183;
  assign new_P1_R1150_U116 = new_P1_R1150_U198 & new_P1_R1150_U199;
  assign new_P1_R1150_U117 = new_P1_R1150_U211 & new_P1_R1150_U185;
  assign new_P1_R1150_U118 = new_P1_R1150_U214 & new_P1_R1150_U215;
  assign new_P1_R1150_U119 = new_P1_R1150_U40 & new_P1_R1150_U354 & new_P1_R1150_U353;
  assign new_P1_R1150_U120 = new_P1_R1150_U357 & new_P1_R1150_U185;
  assign new_P1_R1150_U121 = new_P1_R1150_U230 & new_P1_R1150_U7;
  assign new_P1_R1150_U122 = new_P1_R1150_U364 & new_P1_R1150_U184;
  assign new_P1_R1150_U123 = new_P1_R1150_U29 & new_P1_R1150_U374 & new_P1_R1150_U373;
  assign new_P1_R1150_U124 = new_P1_R1150_U377 & new_P1_R1150_U183;
  assign new_P1_R1150_U125 = new_P1_R1150_U217 & new_P1_R1150_U8;
  assign new_P1_R1150_U126 = new_P1_R1150_U262 & new_P1_R1150_U180;
  assign new_P1_R1150_U127 = new_P1_R1150_U288 & new_P1_R1150_U181;
  assign new_P1_R1150_U128 = new_P1_R1150_U304 & new_P1_R1150_U305;
  assign new_P1_R1150_U129 = new_P1_R1150_U307 & new_P1_R1150_U386;
  assign new_P1_R1150_U130 = new_P1_R1150_U308 & new_P1_R1150_U305 & new_P1_R1150_U304;
  assign new_P1_R1150_U131 = ~new_P1_R1150_U390 | ~new_P1_R1150_U389;
  assign new_P1_R1150_U132 = new_P1_R1150_U85 & new_P1_R1150_U395 & new_P1_R1150_U394;
  assign new_P1_R1150_U133 = new_P1_R1150_U398 & new_P1_R1150_U182;
  assign new_P1_R1150_U134 = ~new_P1_R1150_U404 | ~new_P1_R1150_U403;
  assign new_P1_R1150_U135 = ~new_P1_R1150_U409 | ~new_P1_R1150_U408;
  assign new_P1_R1150_U136 = new_P1_R1150_U415 & new_P1_R1150_U181;
  assign new_P1_R1150_U137 = ~new_P1_R1150_U425 | ~new_P1_R1150_U424;
  assign new_P1_R1150_U138 = ~new_P1_R1150_U430 | ~new_P1_R1150_U429;
  assign new_P1_R1150_U139 = ~new_P1_R1150_U435 | ~new_P1_R1150_U434;
  assign new_P1_R1150_U140 = ~new_P1_R1150_U440 | ~new_P1_R1150_U439;
  assign new_P1_R1150_U141 = ~new_P1_R1150_U445 | ~new_P1_R1150_U444;
  assign new_P1_R1150_U142 = new_P1_R1150_U451 & new_P1_R1150_U180;
  assign new_P1_R1150_U143 = ~new_P1_R1150_U461 | ~new_P1_R1150_U460;
  assign new_P1_R1150_U144 = ~new_P1_R1150_U466 | ~new_P1_R1150_U465;
  assign new_P1_R1150_U145 = new_P1_R1150_U342 & new_P1_R1150_U9;
  assign new_P1_R1150_U146 = new_P1_R1150_U472 & new_P1_R1150_U179;
  assign new_P1_R1150_U147 = new_P1_R1150_U350 & new_P1_R1150_U349;
  assign new_P1_R1150_U148 = ~new_P1_R1150_U118 | ~new_P1_R1150_U212;
  assign new_P1_R1150_U149 = new_P1_R1150_U359 & new_P1_R1150_U358;
  assign new_P1_R1150_U150 = new_P1_R1150_U366 & new_P1_R1150_U365;
  assign new_P1_R1150_U151 = new_P1_R1150_U370 & new_P1_R1150_U369;
  assign new_P1_R1150_U152 = ~new_P1_R1150_U116 | ~new_P1_R1150_U196;
  assign new_P1_R1150_U153 = new_P1_R1150_U379 & new_P1_R1150_U378;
  assign new_P1_R1150_U154 = ~new_P1_U4028;
  assign new_P1_R1150_U155 = ~new_P1_U3055;
  assign new_P1_R1150_U156 = new_P1_R1150_U388 & new_P1_R1150_U387;
  assign new_P1_R1150_U157 = ~new_P1_R1150_U128 | ~new_P1_R1150_U302;
  assign new_P1_R1150_U158 = new_P1_R1150_U400 & new_P1_R1150_U399;
  assign new_P1_R1150_U159 = ~new_P1_R1150_U295 | ~new_P1_R1150_U294;
  assign new_P1_R1150_U160 = ~new_P1_R1150_U291 | ~new_P1_R1150_U290;
  assign new_P1_R1150_U161 = new_P1_R1150_U417 & new_P1_R1150_U416;
  assign new_P1_R1150_U162 = new_P1_R1150_U421 & new_P1_R1150_U420;
  assign new_P1_R1150_U163 = ~new_P1_R1150_U281 | ~new_P1_R1150_U280;
  assign new_P1_R1150_U164 = ~new_P1_R1150_U277 | ~new_P1_R1150_U276;
  assign new_P1_R1150_U165 = ~new_P1_U3461;
  assign new_P1_R1150_U166 = ~new_P1_R1150_U273 | ~new_P1_R1150_U272;
  assign new_P1_R1150_U167 = ~new_P1_U3512;
  assign new_P1_R1150_U168 = ~new_P1_R1150_U265 | ~new_P1_R1150_U264;
  assign new_P1_R1150_U169 = new_P1_R1150_U453 & new_P1_R1150_U452;
  assign new_P1_R1150_U170 = new_P1_R1150_U457 & new_P1_R1150_U456;
  assign new_P1_R1150_U171 = ~new_P1_R1150_U255 | ~new_P1_R1150_U254;
  assign new_P1_R1150_U172 = ~new_P1_R1150_U251 | ~new_P1_R1150_U250;
  assign new_P1_R1150_U173 = ~new_P1_R1150_U247 | ~new_P1_R1150_U246;
  assign new_P1_R1150_U174 = new_P1_R1150_U474 & new_P1_R1150_U473;
  assign new_P1_R1150_U175 = ~new_P1_R1150_U129 | ~new_P1_R1150_U157;
  assign new_P1_R1150_U176 = ~new_P1_R1150_U85;
  assign new_P1_R1150_U177 = ~new_P1_R1150_U29;
  assign new_P1_R1150_U178 = ~new_P1_R1150_U40;
  assign new_P1_R1150_U179 = ~new_P1_U3488 | ~new_P1_R1150_U53;
  assign new_P1_R1150_U180 = ~new_P1_U3503 | ~new_P1_R1150_U62;
  assign new_P1_R1150_U181 = ~new_P1_U4023 | ~new_P1_R1150_U76;
  assign new_P1_R1150_U182 = ~new_P1_U4019 | ~new_P1_R1150_U84;
  assign new_P1_R1150_U183 = ~new_P1_U3464 | ~new_P1_R1150_U28;
  assign new_P1_R1150_U184 = ~new_P1_U3473 | ~new_P1_R1150_U35;
  assign new_P1_R1150_U185 = ~new_P1_U3479 | ~new_P1_R1150_U39;
  assign new_P1_R1150_U186 = ~new_P1_R1150_U64;
  assign new_P1_R1150_U187 = ~new_P1_R1150_U78;
  assign new_P1_R1150_U188 = ~new_P1_R1150_U37;
  assign new_P1_R1150_U189 = ~new_P1_R1150_U54;
  assign new_P1_R1150_U190 = ~new_P1_R1150_U25;
  assign new_P1_R1150_U191 = ~new_P1_R1150_U190 | ~new_P1_R1150_U26;
  assign new_P1_R1150_U192 = ~new_P1_R1150_U191 | ~new_P1_R1150_U165;
  assign new_P1_R1150_U193 = ~new_P1_U3078 | ~new_P1_R1150_U25;
  assign new_P1_R1150_U194 = ~new_P1_R1150_U46;
  assign new_P1_R1150_U195 = ~new_P1_U3467 | ~new_P1_R1150_U30;
  assign new_P1_R1150_U196 = ~new_P1_R1150_U115 | ~new_P1_R1150_U46;
  assign new_P1_R1150_U197 = ~new_P1_R1150_U30 | ~new_P1_R1150_U29;
  assign new_P1_R1150_U198 = ~new_P1_R1150_U197 | ~new_P1_R1150_U27;
  assign new_P1_R1150_U199 = ~new_P1_U3064 | ~new_P1_R1150_U177;
  assign new_P1_R1150_U200 = ~new_P1_R1150_U152;
  assign new_P1_R1150_U201 = ~new_P1_U3476 | ~new_P1_R1150_U34;
  assign new_P1_R1150_U202 = ~new_P1_U3071 | ~new_P1_R1150_U31;
  assign new_P1_R1150_U203 = ~new_P1_U3067 | ~new_P1_R1150_U32;
  assign new_P1_R1150_U204 = ~new_P1_R1150_U188 | ~new_P1_R1150_U6;
  assign new_P1_R1150_U205 = ~new_P1_R1150_U7 | ~new_P1_R1150_U204;
  assign new_P1_R1150_U206 = ~new_P1_U3470 | ~new_P1_R1150_U36;
  assign new_P1_R1150_U207 = ~new_P1_U3476 | ~new_P1_R1150_U34;
  assign new_P1_R1150_U208 = ~new_P1_R1150_U6 | ~new_P1_R1150_U206 | ~new_P1_R1150_U152;
  assign new_P1_R1150_U209 = ~new_P1_R1150_U207 | ~new_P1_R1150_U205;
  assign new_P1_R1150_U210 = ~new_P1_R1150_U44;
  assign new_P1_R1150_U211 = ~new_P1_U3482 | ~new_P1_R1150_U41;
  assign new_P1_R1150_U212 = ~new_P1_R1150_U117 | ~new_P1_R1150_U44;
  assign new_P1_R1150_U213 = ~new_P1_R1150_U41 | ~new_P1_R1150_U40;
  assign new_P1_R1150_U214 = ~new_P1_R1150_U213 | ~new_P1_R1150_U38;
  assign new_P1_R1150_U215 = ~new_P1_U3084 | ~new_P1_R1150_U178;
  assign new_P1_R1150_U216 = ~new_P1_R1150_U148;
  assign new_P1_R1150_U217 = ~new_P1_U3485 | ~new_P1_R1150_U43;
  assign new_P1_R1150_U218 = ~new_P1_R1150_U217 | ~new_P1_R1150_U54;
  assign new_P1_R1150_U219 = ~new_P1_R1150_U210 | ~new_P1_R1150_U40;
  assign new_P1_R1150_U220 = ~new_P1_R1150_U120 | ~new_P1_R1150_U219;
  assign new_P1_R1150_U221 = ~new_P1_R1150_U44 | ~new_P1_R1150_U185;
  assign new_P1_R1150_U222 = ~new_P1_R1150_U119 | ~new_P1_R1150_U221;
  assign new_P1_R1150_U223 = ~new_P1_R1150_U40 | ~new_P1_R1150_U185;
  assign new_P1_R1150_U224 = ~new_P1_R1150_U206 | ~new_P1_R1150_U152;
  assign new_P1_R1150_U225 = ~new_P1_R1150_U45;
  assign new_P1_R1150_U226 = ~new_P1_U3067 | ~new_P1_R1150_U32;
  assign new_P1_R1150_U227 = ~new_P1_R1150_U225 | ~new_P1_R1150_U226;
  assign new_P1_R1150_U228 = ~new_P1_R1150_U122 | ~new_P1_R1150_U227;
  assign new_P1_R1150_U229 = ~new_P1_R1150_U45 | ~new_P1_R1150_U184;
  assign new_P1_R1150_U230 = ~new_P1_U3476 | ~new_P1_R1150_U34;
  assign new_P1_R1150_U231 = ~new_P1_R1150_U121 | ~new_P1_R1150_U229;
  assign new_P1_R1150_U232 = ~new_P1_U3067 | ~new_P1_R1150_U32;
  assign new_P1_R1150_U233 = ~new_P1_R1150_U184 | ~new_P1_R1150_U232;
  assign new_P1_R1150_U234 = ~new_P1_R1150_U206 | ~new_P1_R1150_U37;
  assign new_P1_R1150_U235 = ~new_P1_R1150_U194 | ~new_P1_R1150_U29;
  assign new_P1_R1150_U236 = ~new_P1_R1150_U124 | ~new_P1_R1150_U235;
  assign new_P1_R1150_U237 = ~new_P1_R1150_U46 | ~new_P1_R1150_U183;
  assign new_P1_R1150_U238 = ~new_P1_R1150_U123 | ~new_P1_R1150_U237;
  assign new_P1_R1150_U239 = ~new_P1_R1150_U29 | ~new_P1_R1150_U183;
  assign new_P1_R1150_U240 = ~new_P1_U3491 | ~new_P1_R1150_U52;
  assign new_P1_R1150_U241 = ~new_P1_U3063 | ~new_P1_R1150_U50;
  assign new_P1_R1150_U242 = ~new_P1_U3062 | ~new_P1_R1150_U51;
  assign new_P1_R1150_U243 = ~new_P1_R1150_U189 | ~new_P1_R1150_U8;
  assign new_P1_R1150_U244 = ~new_P1_R1150_U9 | ~new_P1_R1150_U243;
  assign new_P1_R1150_U245 = ~new_P1_U3491 | ~new_P1_R1150_U52;
  assign new_P1_R1150_U246 = ~new_P1_R1150_U125 | ~new_P1_R1150_U148;
  assign new_P1_R1150_U247 = ~new_P1_R1150_U245 | ~new_P1_R1150_U244;
  assign new_P1_R1150_U248 = ~new_P1_R1150_U173;
  assign new_P1_R1150_U249 = ~new_P1_U3494 | ~new_P1_R1150_U56;
  assign new_P1_R1150_U250 = ~new_P1_R1150_U249 | ~new_P1_R1150_U173;
  assign new_P1_R1150_U251 = ~new_P1_U3072 | ~new_P1_R1150_U55;
  assign new_P1_R1150_U252 = ~new_P1_R1150_U172;
  assign new_P1_R1150_U253 = ~new_P1_U3497 | ~new_P1_R1150_U58;
  assign new_P1_R1150_U254 = ~new_P1_R1150_U253 | ~new_P1_R1150_U172;
  assign new_P1_R1150_U255 = ~new_P1_U3080 | ~new_P1_R1150_U57;
  assign new_P1_R1150_U256 = ~new_P1_R1150_U171;
  assign new_P1_R1150_U257 = ~new_P1_U3506 | ~new_P1_R1150_U61;
  assign new_P1_R1150_U258 = ~new_P1_U3073 | ~new_P1_R1150_U59;
  assign new_P1_R1150_U259 = ~new_P1_U3074 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U260 = ~new_P1_R1150_U186 | ~new_P1_R1150_U180;
  assign new_P1_R1150_U261 = ~new_P1_R1150_U10 | ~new_P1_R1150_U260;
  assign new_P1_R1150_U262 = ~new_P1_U3500 | ~new_P1_R1150_U63;
  assign new_P1_R1150_U263 = ~new_P1_U3506 | ~new_P1_R1150_U61;
  assign new_P1_R1150_U264 = ~new_P1_R1150_U257 | ~new_P1_R1150_U171 | ~new_P1_R1150_U126;
  assign new_P1_R1150_U265 = ~new_P1_R1150_U263 | ~new_P1_R1150_U261;
  assign new_P1_R1150_U266 = ~new_P1_R1150_U168;
  assign new_P1_R1150_U267 = ~new_P1_U3509 | ~new_P1_R1150_U66;
  assign new_P1_R1150_U268 = ~new_P1_R1150_U267 | ~new_P1_R1150_U168;
  assign new_P1_R1150_U269 = ~new_P1_U3069 | ~new_P1_R1150_U65;
  assign new_P1_R1150_U270 = ~new_P1_R1150_U67;
  assign new_P1_R1150_U271 = ~new_P1_R1150_U270 | ~new_P1_R1150_U68;
  assign new_P1_R1150_U272 = ~new_P1_R1150_U271 | ~new_P1_R1150_U167;
  assign new_P1_R1150_U273 = ~new_P1_U3082 | ~new_P1_R1150_U67;
  assign new_P1_R1150_U274 = ~new_P1_R1150_U166;
  assign new_P1_R1150_U275 = ~new_P1_U3514 | ~new_P1_R1150_U70;
  assign new_P1_R1150_U276 = ~new_P1_R1150_U275 | ~new_P1_R1150_U166;
  assign new_P1_R1150_U277 = ~new_P1_U3081 | ~new_P1_R1150_U69;
  assign new_P1_R1150_U278 = ~new_P1_R1150_U164;
  assign new_P1_R1150_U279 = ~new_P1_U4025 | ~new_P1_R1150_U72;
  assign new_P1_R1150_U280 = ~new_P1_R1150_U279 | ~new_P1_R1150_U164;
  assign new_P1_R1150_U281 = ~new_P1_U3076 | ~new_P1_R1150_U71;
  assign new_P1_R1150_U282 = ~new_P1_R1150_U163;
  assign new_P1_R1150_U283 = ~new_P1_U4022 | ~new_P1_R1150_U75;
  assign new_P1_R1150_U284 = ~new_P1_U3066 | ~new_P1_R1150_U73;
  assign new_P1_R1150_U285 = ~new_P1_U3061 | ~new_P1_R1150_U48;
  assign new_P1_R1150_U286 = ~new_P1_R1150_U187 | ~new_P1_R1150_U181;
  assign new_P1_R1150_U287 = ~new_P1_R1150_U11 | ~new_P1_R1150_U286;
  assign new_P1_R1150_U288 = ~new_P1_U4024 | ~new_P1_R1150_U77;
  assign new_P1_R1150_U289 = ~new_P1_U4022 | ~new_P1_R1150_U75;
  assign new_P1_R1150_U290 = ~new_P1_R1150_U283 | ~new_P1_R1150_U163 | ~new_P1_R1150_U127;
  assign new_P1_R1150_U291 = ~new_P1_R1150_U289 | ~new_P1_R1150_U287;
  assign new_P1_R1150_U292 = ~new_P1_R1150_U160;
  assign new_P1_R1150_U293 = ~new_P1_U4021 | ~new_P1_R1150_U80;
  assign new_P1_R1150_U294 = ~new_P1_R1150_U293 | ~new_P1_R1150_U160;
  assign new_P1_R1150_U295 = ~new_P1_U3065 | ~new_P1_R1150_U79;
  assign new_P1_R1150_U296 = ~new_P1_R1150_U159;
  assign new_P1_R1150_U297 = ~new_P1_U4020 | ~new_P1_R1150_U82;
  assign new_P1_R1150_U298 = ~new_P1_R1150_U297 | ~new_P1_R1150_U159;
  assign new_P1_R1150_U299 = ~new_P1_U3058 | ~new_P1_R1150_U81;
  assign new_P1_R1150_U300 = ~new_P1_R1150_U89;
  assign new_P1_R1150_U301 = ~new_P1_U4018 | ~new_P1_R1150_U86;
  assign new_P1_R1150_U302 = ~new_P1_R1150_U301 | ~new_P1_R1150_U89 | ~new_P1_R1150_U182;
  assign new_P1_R1150_U303 = ~new_P1_R1150_U86 | ~new_P1_R1150_U85;
  assign new_P1_R1150_U304 = ~new_P1_R1150_U303 | ~new_P1_R1150_U83;
  assign new_P1_R1150_U305 = ~new_P1_U3053 | ~new_P1_R1150_U176;
  assign new_P1_R1150_U306 = ~new_P1_R1150_U157;
  assign new_P1_R1150_U307 = ~new_P1_U4017 | ~new_P1_R1150_U88;
  assign new_P1_R1150_U308 = ~new_P1_U3054 | ~new_P1_R1150_U87;
  assign new_P1_R1150_U309 = ~new_P1_R1150_U300 | ~new_P1_R1150_U85;
  assign new_P1_R1150_U310 = ~new_P1_R1150_U133 | ~new_P1_R1150_U309;
  assign new_P1_R1150_U311 = ~new_P1_R1150_U89 | ~new_P1_R1150_U182;
  assign new_P1_R1150_U312 = ~new_P1_R1150_U132 | ~new_P1_R1150_U311;
  assign new_P1_R1150_U313 = ~new_P1_R1150_U85 | ~new_P1_R1150_U182;
  assign new_P1_R1150_U314 = ~new_P1_R1150_U288 | ~new_P1_R1150_U163;
  assign new_P1_R1150_U315 = ~new_P1_R1150_U90;
  assign new_P1_R1150_U316 = ~new_P1_U3061 | ~new_P1_R1150_U48;
  assign new_P1_R1150_U317 = ~new_P1_R1150_U315 | ~new_P1_R1150_U316;
  assign new_P1_R1150_U318 = ~new_P1_R1150_U136 | ~new_P1_R1150_U317;
  assign new_P1_R1150_U319 = ~new_P1_R1150_U90 | ~new_P1_R1150_U181;
  assign new_P1_R1150_U320 = ~new_P1_U4022 | ~new_P1_R1150_U75;
  assign new_P1_R1150_U321 = ~new_P1_R1150_U11 | ~new_P1_R1150_U320 | ~new_P1_R1150_U319;
  assign new_P1_R1150_U322 = ~new_P1_U3061 | ~new_P1_R1150_U48;
  assign new_P1_R1150_U323 = ~new_P1_R1150_U181 | ~new_P1_R1150_U322;
  assign new_P1_R1150_U324 = ~new_P1_R1150_U288 | ~new_P1_R1150_U78;
  assign new_P1_R1150_U325 = ~new_P1_R1150_U262 | ~new_P1_R1150_U171;
  assign new_P1_R1150_U326 = ~new_P1_R1150_U91;
  assign new_P1_R1150_U327 = ~new_P1_U3074 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U328 = ~new_P1_R1150_U326 | ~new_P1_R1150_U327;
  assign new_P1_R1150_U329 = ~new_P1_R1150_U142 | ~new_P1_R1150_U328;
  assign new_P1_R1150_U330 = ~new_P1_R1150_U91 | ~new_P1_R1150_U180;
  assign new_P1_R1150_U331 = ~new_P1_U3506 | ~new_P1_R1150_U61;
  assign new_P1_R1150_U332 = ~new_P1_R1150_U10 | ~new_P1_R1150_U331 | ~new_P1_R1150_U330;
  assign new_P1_R1150_U333 = ~new_P1_U3074 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U334 = ~new_P1_R1150_U180 | ~new_P1_R1150_U333;
  assign new_P1_R1150_U335 = ~new_P1_R1150_U262 | ~new_P1_R1150_U64;
  assign new_P1_R1150_U336 = ~new_P1_R1150_U217 | ~new_P1_R1150_U148;
  assign new_P1_R1150_U337 = ~new_P1_R1150_U92;
  assign new_P1_R1150_U338 = ~new_P1_U3062 | ~new_P1_R1150_U51;
  assign new_P1_R1150_U339 = ~new_P1_R1150_U337 | ~new_P1_R1150_U338;
  assign new_P1_R1150_U340 = ~new_P1_R1150_U146 | ~new_P1_R1150_U339;
  assign new_P1_R1150_U341 = ~new_P1_R1150_U92 | ~new_P1_R1150_U179;
  assign new_P1_R1150_U342 = ~new_P1_U3491 | ~new_P1_R1150_U52;
  assign new_P1_R1150_U343 = ~new_P1_R1150_U145 | ~new_P1_R1150_U341;
  assign new_P1_R1150_U344 = ~new_P1_U3062 | ~new_P1_R1150_U51;
  assign new_P1_R1150_U345 = ~new_P1_R1150_U179 | ~new_P1_R1150_U344;
  assign new_P1_R1150_U346 = ~new_P1_U3077 | ~new_P1_R1150_U24;
  assign new_P1_R1150_U347 = ~new_P1_R1150_U301 | ~new_P1_R1150_U89 | ~new_P1_R1150_U182;
  assign new_P1_R1150_U348 = ~new_P1_R1150_U130 | ~new_P1_R1150_U12 | ~new_P1_R1150_U347;
  assign new_P1_R1150_U349 = ~new_P1_U3485 | ~new_P1_R1150_U43;
  assign new_P1_R1150_U350 = ~new_P1_U3083 | ~new_P1_R1150_U42;
  assign new_P1_R1150_U351 = ~new_P1_R1150_U218 | ~new_P1_R1150_U148;
  assign new_P1_R1150_U352 = ~new_P1_R1150_U216 | ~new_P1_R1150_U147;
  assign new_P1_R1150_U353 = ~new_P1_U3482 | ~new_P1_R1150_U41;
  assign new_P1_R1150_U354 = ~new_P1_U3084 | ~new_P1_R1150_U38;
  assign new_P1_R1150_U355 = ~new_P1_U3482 | ~new_P1_R1150_U41;
  assign new_P1_R1150_U356 = ~new_P1_U3084 | ~new_P1_R1150_U38;
  assign new_P1_R1150_U357 = ~new_P1_R1150_U356 | ~new_P1_R1150_U355;
  assign new_P1_R1150_U358 = ~new_P1_U3479 | ~new_P1_R1150_U39;
  assign new_P1_R1150_U359 = ~new_P1_U3070 | ~new_P1_R1150_U22;
  assign new_P1_R1150_U360 = ~new_P1_R1150_U223 | ~new_P1_R1150_U44;
  assign new_P1_R1150_U361 = ~new_P1_R1150_U149 | ~new_P1_R1150_U210;
  assign new_P1_R1150_U362 = ~new_P1_U3476 | ~new_P1_R1150_U34;
  assign new_P1_R1150_U363 = ~new_P1_U3071 | ~new_P1_R1150_U31;
  assign new_P1_R1150_U364 = ~new_P1_R1150_U363 | ~new_P1_R1150_U362;
  assign new_P1_R1150_U365 = ~new_P1_U3473 | ~new_P1_R1150_U35;
  assign new_P1_R1150_U366 = ~new_P1_U3067 | ~new_P1_R1150_U32;
  assign new_P1_R1150_U367 = ~new_P1_R1150_U233 | ~new_P1_R1150_U45;
  assign new_P1_R1150_U368 = ~new_P1_R1150_U150 | ~new_P1_R1150_U225;
  assign new_P1_R1150_U369 = ~new_P1_U3470 | ~new_P1_R1150_U36;
  assign new_P1_R1150_U370 = ~new_P1_U3060 | ~new_P1_R1150_U33;
  assign new_P1_R1150_U371 = ~new_P1_R1150_U234 | ~new_P1_R1150_U152;
  assign new_P1_R1150_U372 = ~new_P1_R1150_U200 | ~new_P1_R1150_U151;
  assign new_P1_R1150_U373 = ~new_P1_U3467 | ~new_P1_R1150_U30;
  assign new_P1_R1150_U374 = ~new_P1_U3064 | ~new_P1_R1150_U27;
  assign new_P1_R1150_U375 = ~new_P1_U3467 | ~new_P1_R1150_U30;
  assign new_P1_R1150_U376 = ~new_P1_U3064 | ~new_P1_R1150_U27;
  assign new_P1_R1150_U377 = ~new_P1_R1150_U376 | ~new_P1_R1150_U375;
  assign new_P1_R1150_U378 = ~new_P1_U3464 | ~new_P1_R1150_U28;
  assign new_P1_R1150_U379 = ~new_P1_U3068 | ~new_P1_R1150_U23;
  assign new_P1_R1150_U380 = ~new_P1_R1150_U239 | ~new_P1_R1150_U46;
  assign new_P1_R1150_U381 = ~new_P1_R1150_U153 | ~new_P1_R1150_U194;
  assign new_P1_R1150_U382 = ~new_P1_U4028 | ~new_P1_R1150_U155;
  assign new_P1_R1150_U383 = ~new_P1_U3055 | ~new_P1_R1150_U154;
  assign new_P1_R1150_U384 = ~new_P1_U4028 | ~new_P1_R1150_U155;
  assign new_P1_R1150_U385 = ~new_P1_U3055 | ~new_P1_R1150_U154;
  assign new_P1_R1150_U386 = ~new_P1_R1150_U385 | ~new_P1_R1150_U384;
  assign new_P1_R1150_U387 = ~new_P1_R1150_U87 | ~new_P1_U3054 | ~new_P1_R1150_U386;
  assign new_P1_R1150_U388 = ~new_P1_U4017 | ~new_P1_R1150_U12 | ~new_P1_R1150_U88;
  assign new_P1_R1150_U389 = ~new_P1_U4017 | ~new_P1_R1150_U88;
  assign new_P1_R1150_U390 = ~new_P1_U3054 | ~new_P1_R1150_U87;
  assign new_P1_R1150_U391 = ~new_P1_R1150_U131;
  assign new_P1_R1150_U392 = ~new_P1_R1150_U306 | ~new_P1_R1150_U391;
  assign new_P1_R1150_U393 = ~new_P1_R1150_U131 | ~new_P1_R1150_U157;
  assign new_P1_R1150_U394 = ~new_P1_U4018 | ~new_P1_R1150_U86;
  assign new_P1_R1150_U395 = ~new_P1_U3053 | ~new_P1_R1150_U83;
  assign new_P1_R1150_U396 = ~new_P1_U4018 | ~new_P1_R1150_U86;
  assign new_P1_R1150_U397 = ~new_P1_U3053 | ~new_P1_R1150_U83;
  assign new_P1_R1150_U398 = ~new_P1_R1150_U397 | ~new_P1_R1150_U396;
  assign new_P1_R1150_U399 = ~new_P1_U4019 | ~new_P1_R1150_U84;
  assign new_P1_R1150_U400 = ~new_P1_U3057 | ~new_P1_R1150_U47;
  assign new_P1_R1150_U401 = ~new_P1_R1150_U313 | ~new_P1_R1150_U89;
  assign new_P1_R1150_U402 = ~new_P1_R1150_U158 | ~new_P1_R1150_U300;
  assign new_P1_R1150_U403 = ~new_P1_U4020 | ~new_P1_R1150_U82;
  assign new_P1_R1150_U404 = ~new_P1_U3058 | ~new_P1_R1150_U81;
  assign new_P1_R1150_U405 = ~new_P1_R1150_U134;
  assign new_P1_R1150_U406 = ~new_P1_R1150_U296 | ~new_P1_R1150_U405;
  assign new_P1_R1150_U407 = ~new_P1_R1150_U134 | ~new_P1_R1150_U159;
  assign new_P1_R1150_U408 = ~new_P1_U4021 | ~new_P1_R1150_U80;
  assign new_P1_R1150_U409 = ~new_P1_U3065 | ~new_P1_R1150_U79;
  assign new_P1_R1150_U410 = ~new_P1_R1150_U135;
  assign new_P1_R1150_U411 = ~new_P1_R1150_U292 | ~new_P1_R1150_U410;
  assign new_P1_R1150_U412 = ~new_P1_R1150_U135 | ~new_P1_R1150_U160;
  assign new_P1_R1150_U413 = ~new_P1_U4022 | ~new_P1_R1150_U75;
  assign new_P1_R1150_U414 = ~new_P1_U3066 | ~new_P1_R1150_U73;
  assign new_P1_R1150_U415 = ~new_P1_R1150_U414 | ~new_P1_R1150_U413;
  assign new_P1_R1150_U416 = ~new_P1_U4023 | ~new_P1_R1150_U76;
  assign new_P1_R1150_U417 = ~new_P1_U3061 | ~new_P1_R1150_U48;
  assign new_P1_R1150_U418 = ~new_P1_R1150_U323 | ~new_P1_R1150_U90;
  assign new_P1_R1150_U419 = ~new_P1_R1150_U161 | ~new_P1_R1150_U315;
  assign new_P1_R1150_U420 = ~new_P1_U4024 | ~new_P1_R1150_U77;
  assign new_P1_R1150_U421 = ~new_P1_U3075 | ~new_P1_R1150_U74;
  assign new_P1_R1150_U422 = ~new_P1_R1150_U324 | ~new_P1_R1150_U163;
  assign new_P1_R1150_U423 = ~new_P1_R1150_U282 | ~new_P1_R1150_U162;
  assign new_P1_R1150_U424 = ~new_P1_U4025 | ~new_P1_R1150_U72;
  assign new_P1_R1150_U425 = ~new_P1_U3076 | ~new_P1_R1150_U71;
  assign new_P1_R1150_U426 = ~new_P1_R1150_U137;
  assign new_P1_R1150_U427 = ~new_P1_R1150_U278 | ~new_P1_R1150_U426;
  assign new_P1_R1150_U428 = ~new_P1_R1150_U137 | ~new_P1_R1150_U164;
  assign new_P1_R1150_U429 = ~new_P1_U3461 | ~new_P1_R1150_U26;
  assign new_P1_R1150_U430 = ~new_P1_U3078 | ~new_P1_R1150_U165;
  assign new_P1_R1150_U431 = ~new_P1_R1150_U138;
  assign new_P1_R1150_U432 = ~new_P1_R1150_U431 | ~new_P1_R1150_U190;
  assign new_P1_R1150_U433 = ~new_P1_R1150_U138 | ~new_P1_R1150_U25;
  assign new_P1_R1150_U434 = ~new_P1_U3514 | ~new_P1_R1150_U70;
  assign new_P1_R1150_U435 = ~new_P1_U3081 | ~new_P1_R1150_U69;
  assign new_P1_R1150_U436 = ~new_P1_R1150_U139;
  assign new_P1_R1150_U437 = ~new_P1_R1150_U274 | ~new_P1_R1150_U436;
  assign new_P1_R1150_U438 = ~new_P1_R1150_U139 | ~new_P1_R1150_U166;
  assign new_P1_R1150_U439 = ~new_P1_U3512 | ~new_P1_R1150_U68;
  assign new_P1_R1150_U440 = ~new_P1_U3082 | ~new_P1_R1150_U167;
  assign new_P1_R1150_U441 = ~new_P1_R1150_U140;
  assign new_P1_R1150_U442 = ~new_P1_R1150_U441 | ~new_P1_R1150_U270;
  assign new_P1_R1150_U443 = ~new_P1_R1150_U140 | ~new_P1_R1150_U67;
  assign new_P1_R1150_U444 = ~new_P1_U3509 | ~new_P1_R1150_U66;
  assign new_P1_R1150_U445 = ~new_P1_U3069 | ~new_P1_R1150_U65;
  assign new_P1_R1150_U446 = ~new_P1_R1150_U141;
  assign new_P1_R1150_U447 = ~new_P1_R1150_U266 | ~new_P1_R1150_U446;
  assign new_P1_R1150_U448 = ~new_P1_R1150_U141 | ~new_P1_R1150_U168;
  assign new_P1_R1150_U449 = ~new_P1_U3506 | ~new_P1_R1150_U61;
  assign new_P1_R1150_U450 = ~new_P1_U3073 | ~new_P1_R1150_U59;
  assign new_P1_R1150_U451 = ~new_P1_R1150_U450 | ~new_P1_R1150_U449;
  assign new_P1_R1150_U452 = ~new_P1_U3503 | ~new_P1_R1150_U62;
  assign new_P1_R1150_U453 = ~new_P1_U3074 | ~new_P1_R1150_U49;
  assign new_P1_R1150_U454 = ~new_P1_R1150_U334 | ~new_P1_R1150_U91;
  assign new_P1_R1150_U455 = ~new_P1_R1150_U169 | ~new_P1_R1150_U326;
  assign new_P1_R1150_U456 = ~new_P1_U3500 | ~new_P1_R1150_U63;
  assign new_P1_R1150_U457 = ~new_P1_U3079 | ~new_P1_R1150_U60;
  assign new_P1_R1150_U458 = ~new_P1_R1150_U335 | ~new_P1_R1150_U171;
  assign new_P1_R1150_U459 = ~new_P1_R1150_U256 | ~new_P1_R1150_U170;
  assign new_P1_R1150_U460 = ~new_P1_U3497 | ~new_P1_R1150_U58;
  assign new_P1_R1150_U461 = ~new_P1_U3080 | ~new_P1_R1150_U57;
  assign new_P1_R1150_U462 = ~new_P1_R1150_U143;
  assign new_P1_R1150_U463 = ~new_P1_R1150_U252 | ~new_P1_R1150_U462;
  assign new_P1_R1150_U464 = ~new_P1_R1150_U143 | ~new_P1_R1150_U172;
  assign new_P1_R1150_U465 = ~new_P1_U3494 | ~new_P1_R1150_U56;
  assign new_P1_R1150_U466 = ~new_P1_U3072 | ~new_P1_R1150_U55;
  assign new_P1_R1150_U467 = ~new_P1_R1150_U144;
  assign new_P1_R1150_U468 = ~new_P1_R1150_U248 | ~new_P1_R1150_U467;
  assign new_P1_R1150_U469 = ~new_P1_R1150_U144 | ~new_P1_R1150_U173;
  assign new_P1_R1150_U470 = ~new_P1_U3491 | ~new_P1_R1150_U52;
  assign new_P1_R1150_U471 = ~new_P1_U3063 | ~new_P1_R1150_U50;
  assign new_P1_R1150_U472 = ~new_P1_R1150_U471 | ~new_P1_R1150_U470;
  assign new_P1_R1150_U473 = ~new_P1_U3488 | ~new_P1_R1150_U53;
  assign new_P1_R1150_U474 = ~new_P1_U3062 | ~new_P1_R1150_U51;
  assign new_P1_R1150_U475 = ~new_P1_R1150_U345 | ~new_P1_R1150_U92;
  assign new_P1_R1150_U476 = ~new_P1_R1150_U174 | ~new_P1_R1150_U337;
  assign new_P1_R1192_U6 = new_P1_R1192_U184 & new_P1_R1192_U201;
  assign new_P1_R1192_U7 = new_P1_R1192_U203 & new_P1_R1192_U202;
  assign new_P1_R1192_U8 = new_P1_R1192_U179 & new_P1_R1192_U240;
  assign new_P1_R1192_U9 = new_P1_R1192_U242 & new_P1_R1192_U241;
  assign new_P1_R1192_U10 = new_P1_R1192_U259 & new_P1_R1192_U258;
  assign new_P1_R1192_U11 = new_P1_R1192_U285 & new_P1_R1192_U284;
  assign new_P1_R1192_U12 = new_P1_R1192_U383 & new_P1_R1192_U382;
  assign new_P1_R1192_U13 = ~new_P1_R1192_U340 | ~new_P1_R1192_U343;
  assign new_P1_R1192_U14 = ~new_P1_R1192_U329 | ~new_P1_R1192_U332;
  assign new_P1_R1192_U15 = ~new_P1_R1192_U318 | ~new_P1_R1192_U321;
  assign new_P1_R1192_U16 = ~new_P1_R1192_U310 | ~new_P1_R1192_U312;
  assign new_P1_R1192_U17 = ~new_P1_R1192_U348 | ~new_P1_R1192_U156 | ~new_P1_R1192_U175;
  assign new_P1_R1192_U18 = ~new_P1_R1192_U236 | ~new_P1_R1192_U238;
  assign new_P1_R1192_U19 = ~new_P1_R1192_U228 | ~new_P1_R1192_U231;
  assign new_P1_R1192_U20 = ~new_P1_R1192_U220 | ~new_P1_R1192_U222;
  assign new_P1_R1192_U21 = ~new_P1_R1192_U25 | ~new_P1_R1192_U346;
  assign new_P1_R1192_U22 = ~new_P1_U3479;
  assign new_P1_R1192_U23 = ~new_P1_U3464;
  assign new_P1_R1192_U24 = ~new_P1_U3456;
  assign new_P1_R1192_U25 = ~new_P1_U3456 | ~new_P1_R1192_U93;
  assign new_P1_R1192_U26 = ~new_P1_U3078;
  assign new_P1_R1192_U27 = ~new_P1_U3467;
  assign new_P1_R1192_U28 = ~new_P1_U3068;
  assign new_P1_R1192_U29 = ~new_P1_U3068 | ~new_P1_R1192_U23;
  assign new_P1_R1192_U30 = ~new_P1_U3064;
  assign new_P1_R1192_U31 = ~new_P1_U3476;
  assign new_P1_R1192_U32 = ~new_P1_U3473;
  assign new_P1_R1192_U33 = ~new_P1_U3470;
  assign new_P1_R1192_U34 = ~new_P1_U3071;
  assign new_P1_R1192_U35 = ~new_P1_U3067;
  assign new_P1_R1192_U36 = ~new_P1_U3060;
  assign new_P1_R1192_U37 = ~new_P1_U3060 | ~new_P1_R1192_U33;
  assign new_P1_R1192_U38 = ~new_P1_U3482;
  assign new_P1_R1192_U39 = ~new_P1_U3070;
  assign new_P1_R1192_U40 = ~new_P1_U3070 | ~new_P1_R1192_U22;
  assign new_P1_R1192_U41 = ~new_P1_U3084;
  assign new_P1_R1192_U42 = ~new_P1_U3485;
  assign new_P1_R1192_U43 = ~new_P1_U3083;
  assign new_P1_R1192_U44 = ~new_P1_R1192_U209 | ~new_P1_R1192_U208;
  assign new_P1_R1192_U45 = ~new_P1_R1192_U37 | ~new_P1_R1192_U224;
  assign new_P1_R1192_U46 = ~new_P1_R1192_U193 | ~new_P1_R1192_U192;
  assign new_P1_R1192_U47 = ~new_P1_U4019;
  assign new_P1_R1192_U48 = ~new_P1_U4023;
  assign new_P1_R1192_U49 = ~new_P1_U3503;
  assign new_P1_R1192_U50 = ~new_P1_U3491;
  assign new_P1_R1192_U51 = ~new_P1_U3488;
  assign new_P1_R1192_U52 = ~new_P1_U3063;
  assign new_P1_R1192_U53 = ~new_P1_U3062;
  assign new_P1_R1192_U54 = ~new_P1_U3083 | ~new_P1_R1192_U42;
  assign new_P1_R1192_U55 = ~new_P1_U3494;
  assign new_P1_R1192_U56 = ~new_P1_U3072;
  assign new_P1_R1192_U57 = ~new_P1_U3497;
  assign new_P1_R1192_U58 = ~new_P1_U3080;
  assign new_P1_R1192_U59 = ~new_P1_U3506;
  assign new_P1_R1192_U60 = ~new_P1_U3500;
  assign new_P1_R1192_U61 = ~new_P1_U3073;
  assign new_P1_R1192_U62 = ~new_P1_U3074;
  assign new_P1_R1192_U63 = ~new_P1_U3079;
  assign new_P1_R1192_U64 = ~new_P1_U3079 | ~new_P1_R1192_U60;
  assign new_P1_R1192_U65 = ~new_P1_U3509;
  assign new_P1_R1192_U66 = ~new_P1_U3069;
  assign new_P1_R1192_U67 = ~new_P1_R1192_U269 | ~new_P1_R1192_U268;
  assign new_P1_R1192_U68 = ~new_P1_U3082;
  assign new_P1_R1192_U69 = ~new_P1_U3514;
  assign new_P1_R1192_U70 = ~new_P1_U3081;
  assign new_P1_R1192_U71 = ~new_P1_U4025;
  assign new_P1_R1192_U72 = ~new_P1_U3076;
  assign new_P1_R1192_U73 = ~new_P1_U4022;
  assign new_P1_R1192_U74 = ~new_P1_U4024;
  assign new_P1_R1192_U75 = ~new_P1_U3066;
  assign new_P1_R1192_U76 = ~new_P1_U3061;
  assign new_P1_R1192_U77 = ~new_P1_U3075;
  assign new_P1_R1192_U78 = ~new_P1_U3075 | ~new_P1_R1192_U74;
  assign new_P1_R1192_U79 = ~new_P1_U4021;
  assign new_P1_R1192_U80 = ~new_P1_U3065;
  assign new_P1_R1192_U81 = ~new_P1_U4020;
  assign new_P1_R1192_U82 = ~new_P1_U3058;
  assign new_P1_R1192_U83 = ~new_P1_U4018;
  assign new_P1_R1192_U84 = ~new_P1_U3057;
  assign new_P1_R1192_U85 = ~new_P1_U3057 | ~new_P1_R1192_U47;
  assign new_P1_R1192_U86 = ~new_P1_U3053;
  assign new_P1_R1192_U87 = ~new_P1_U4017;
  assign new_P1_R1192_U88 = ~new_P1_U3054;
  assign new_P1_R1192_U89 = ~new_P1_R1192_U299 | ~new_P1_R1192_U298;
  assign new_P1_R1192_U90 = ~new_P1_R1192_U78 | ~new_P1_R1192_U314;
  assign new_P1_R1192_U91 = ~new_P1_R1192_U64 | ~new_P1_R1192_U325;
  assign new_P1_R1192_U92 = ~new_P1_R1192_U54 | ~new_P1_R1192_U336;
  assign new_P1_R1192_U93 = ~new_P1_U3077;
  assign new_P1_R1192_U94 = ~new_P1_R1192_U393 | ~new_P1_R1192_U392;
  assign new_P1_R1192_U95 = ~new_P1_R1192_U407 | ~new_P1_R1192_U406;
  assign new_P1_R1192_U96 = ~new_P1_R1192_U412 | ~new_P1_R1192_U411;
  assign new_P1_R1192_U97 = ~new_P1_R1192_U428 | ~new_P1_R1192_U427;
  assign new_P1_R1192_U98 = ~new_P1_R1192_U433 | ~new_P1_R1192_U432;
  assign new_P1_R1192_U99 = ~new_P1_R1192_U438 | ~new_P1_R1192_U437;
  assign new_P1_R1192_U100 = ~new_P1_R1192_U443 | ~new_P1_R1192_U442;
  assign new_P1_R1192_U101 = ~new_P1_R1192_U448 | ~new_P1_R1192_U447;
  assign new_P1_R1192_U102 = ~new_P1_R1192_U464 | ~new_P1_R1192_U463;
  assign new_P1_R1192_U103 = ~new_P1_R1192_U469 | ~new_P1_R1192_U468;
  assign new_P1_R1192_U104 = ~new_P1_R1192_U352 | ~new_P1_R1192_U351;
  assign new_P1_R1192_U105 = ~new_P1_R1192_U361 | ~new_P1_R1192_U360;
  assign new_P1_R1192_U106 = ~new_P1_R1192_U368 | ~new_P1_R1192_U367;
  assign new_P1_R1192_U107 = ~new_P1_R1192_U372 | ~new_P1_R1192_U371;
  assign new_P1_R1192_U108 = ~new_P1_R1192_U381 | ~new_P1_R1192_U380;
  assign new_P1_R1192_U109 = ~new_P1_R1192_U402 | ~new_P1_R1192_U401;
  assign new_P1_R1192_U110 = ~new_P1_R1192_U419 | ~new_P1_R1192_U418;
  assign new_P1_R1192_U111 = ~new_P1_R1192_U423 | ~new_P1_R1192_U422;
  assign new_P1_R1192_U112 = ~new_P1_R1192_U455 | ~new_P1_R1192_U454;
  assign new_P1_R1192_U113 = ~new_P1_R1192_U459 | ~new_P1_R1192_U458;
  assign new_P1_R1192_U114 = ~new_P1_R1192_U476 | ~new_P1_R1192_U475;
  assign new_P1_R1192_U115 = new_P1_R1192_U195 & new_P1_R1192_U183;
  assign new_P1_R1192_U116 = new_P1_R1192_U198 & new_P1_R1192_U199;
  assign new_P1_R1192_U117 = new_P1_R1192_U211 & new_P1_R1192_U185;
  assign new_P1_R1192_U118 = new_P1_R1192_U214 & new_P1_R1192_U215;
  assign new_P1_R1192_U119 = new_P1_R1192_U40 & new_P1_R1192_U354 & new_P1_R1192_U353;
  assign new_P1_R1192_U120 = new_P1_R1192_U357 & new_P1_R1192_U185;
  assign new_P1_R1192_U121 = new_P1_R1192_U230 & new_P1_R1192_U7;
  assign new_P1_R1192_U122 = new_P1_R1192_U364 & new_P1_R1192_U184;
  assign new_P1_R1192_U123 = new_P1_R1192_U29 & new_P1_R1192_U374 & new_P1_R1192_U373;
  assign new_P1_R1192_U124 = new_P1_R1192_U377 & new_P1_R1192_U183;
  assign new_P1_R1192_U125 = new_P1_R1192_U217 & new_P1_R1192_U8;
  assign new_P1_R1192_U126 = new_P1_R1192_U262 & new_P1_R1192_U180;
  assign new_P1_R1192_U127 = new_P1_R1192_U288 & new_P1_R1192_U181;
  assign new_P1_R1192_U128 = new_P1_R1192_U304 & new_P1_R1192_U305;
  assign new_P1_R1192_U129 = new_P1_R1192_U307 & new_P1_R1192_U386;
  assign new_P1_R1192_U130 = new_P1_R1192_U308 & new_P1_R1192_U305 & new_P1_R1192_U304;
  assign new_P1_R1192_U131 = ~new_P1_R1192_U390 | ~new_P1_R1192_U389;
  assign new_P1_R1192_U132 = new_P1_R1192_U85 & new_P1_R1192_U395 & new_P1_R1192_U394;
  assign new_P1_R1192_U133 = new_P1_R1192_U398 & new_P1_R1192_U182;
  assign new_P1_R1192_U134 = ~new_P1_R1192_U404 | ~new_P1_R1192_U403;
  assign new_P1_R1192_U135 = ~new_P1_R1192_U409 | ~new_P1_R1192_U408;
  assign new_P1_R1192_U136 = new_P1_R1192_U415 & new_P1_R1192_U181;
  assign new_P1_R1192_U137 = ~new_P1_R1192_U425 | ~new_P1_R1192_U424;
  assign new_P1_R1192_U138 = ~new_P1_R1192_U430 | ~new_P1_R1192_U429;
  assign new_P1_R1192_U139 = ~new_P1_R1192_U435 | ~new_P1_R1192_U434;
  assign new_P1_R1192_U140 = ~new_P1_R1192_U440 | ~new_P1_R1192_U439;
  assign new_P1_R1192_U141 = ~new_P1_R1192_U445 | ~new_P1_R1192_U444;
  assign new_P1_R1192_U142 = new_P1_R1192_U451 & new_P1_R1192_U180;
  assign new_P1_R1192_U143 = ~new_P1_R1192_U461 | ~new_P1_R1192_U460;
  assign new_P1_R1192_U144 = ~new_P1_R1192_U466 | ~new_P1_R1192_U465;
  assign new_P1_R1192_U145 = new_P1_R1192_U342 & new_P1_R1192_U9;
  assign new_P1_R1192_U146 = new_P1_R1192_U472 & new_P1_R1192_U179;
  assign new_P1_R1192_U147 = new_P1_R1192_U350 & new_P1_R1192_U349;
  assign new_P1_R1192_U148 = ~new_P1_R1192_U118 | ~new_P1_R1192_U212;
  assign new_P1_R1192_U149 = new_P1_R1192_U359 & new_P1_R1192_U358;
  assign new_P1_R1192_U150 = new_P1_R1192_U366 & new_P1_R1192_U365;
  assign new_P1_R1192_U151 = new_P1_R1192_U370 & new_P1_R1192_U369;
  assign new_P1_R1192_U152 = ~new_P1_R1192_U116 | ~new_P1_R1192_U196;
  assign new_P1_R1192_U153 = new_P1_R1192_U379 & new_P1_R1192_U378;
  assign new_P1_R1192_U154 = ~new_P1_U4028;
  assign new_P1_R1192_U155 = ~new_P1_U3055;
  assign new_P1_R1192_U156 = new_P1_R1192_U388 & new_P1_R1192_U387;
  assign new_P1_R1192_U157 = ~new_P1_R1192_U128 | ~new_P1_R1192_U302;
  assign new_P1_R1192_U158 = new_P1_R1192_U400 & new_P1_R1192_U399;
  assign new_P1_R1192_U159 = ~new_P1_R1192_U295 | ~new_P1_R1192_U294;
  assign new_P1_R1192_U160 = ~new_P1_R1192_U291 | ~new_P1_R1192_U290;
  assign new_P1_R1192_U161 = new_P1_R1192_U417 & new_P1_R1192_U416;
  assign new_P1_R1192_U162 = new_P1_R1192_U421 & new_P1_R1192_U420;
  assign new_P1_R1192_U163 = ~new_P1_R1192_U281 | ~new_P1_R1192_U280;
  assign new_P1_R1192_U164 = ~new_P1_R1192_U277 | ~new_P1_R1192_U276;
  assign new_P1_R1192_U165 = ~new_P1_U3461;
  assign new_P1_R1192_U166 = ~new_P1_R1192_U273 | ~new_P1_R1192_U272;
  assign new_P1_R1192_U167 = ~new_P1_U3512;
  assign new_P1_R1192_U168 = ~new_P1_R1192_U265 | ~new_P1_R1192_U264;
  assign new_P1_R1192_U169 = new_P1_R1192_U453 & new_P1_R1192_U452;
  assign new_P1_R1192_U170 = new_P1_R1192_U457 & new_P1_R1192_U456;
  assign new_P1_R1192_U171 = ~new_P1_R1192_U255 | ~new_P1_R1192_U254;
  assign new_P1_R1192_U172 = ~new_P1_R1192_U251 | ~new_P1_R1192_U250;
  assign new_P1_R1192_U173 = ~new_P1_R1192_U247 | ~new_P1_R1192_U246;
  assign new_P1_R1192_U174 = new_P1_R1192_U474 & new_P1_R1192_U473;
  assign new_P1_R1192_U175 = ~new_P1_R1192_U129 | ~new_P1_R1192_U157;
  assign new_P1_R1192_U176 = ~new_P1_R1192_U85;
  assign new_P1_R1192_U177 = ~new_P1_R1192_U29;
  assign new_P1_R1192_U178 = ~new_P1_R1192_U40;
  assign new_P1_R1192_U179 = ~new_P1_U3488 | ~new_P1_R1192_U53;
  assign new_P1_R1192_U180 = ~new_P1_U3503 | ~new_P1_R1192_U62;
  assign new_P1_R1192_U181 = ~new_P1_U4023 | ~new_P1_R1192_U76;
  assign new_P1_R1192_U182 = ~new_P1_U4019 | ~new_P1_R1192_U84;
  assign new_P1_R1192_U183 = ~new_P1_U3464 | ~new_P1_R1192_U28;
  assign new_P1_R1192_U184 = ~new_P1_U3473 | ~new_P1_R1192_U35;
  assign new_P1_R1192_U185 = ~new_P1_U3479 | ~new_P1_R1192_U39;
  assign new_P1_R1192_U186 = ~new_P1_R1192_U64;
  assign new_P1_R1192_U187 = ~new_P1_R1192_U78;
  assign new_P1_R1192_U188 = ~new_P1_R1192_U37;
  assign new_P1_R1192_U189 = ~new_P1_R1192_U54;
  assign new_P1_R1192_U190 = ~new_P1_R1192_U25;
  assign new_P1_R1192_U191 = ~new_P1_R1192_U190 | ~new_P1_R1192_U26;
  assign new_P1_R1192_U192 = ~new_P1_R1192_U191 | ~new_P1_R1192_U165;
  assign new_P1_R1192_U193 = ~new_P1_U3078 | ~new_P1_R1192_U25;
  assign new_P1_R1192_U194 = ~new_P1_R1192_U46;
  assign new_P1_R1192_U195 = ~new_P1_U3467 | ~new_P1_R1192_U30;
  assign new_P1_R1192_U196 = ~new_P1_R1192_U115 | ~new_P1_R1192_U46;
  assign new_P1_R1192_U197 = ~new_P1_R1192_U30 | ~new_P1_R1192_U29;
  assign new_P1_R1192_U198 = ~new_P1_R1192_U197 | ~new_P1_R1192_U27;
  assign new_P1_R1192_U199 = ~new_P1_U3064 | ~new_P1_R1192_U177;
  assign new_P1_R1192_U200 = ~new_P1_R1192_U152;
  assign new_P1_R1192_U201 = ~new_P1_U3476 | ~new_P1_R1192_U34;
  assign new_P1_R1192_U202 = ~new_P1_U3071 | ~new_P1_R1192_U31;
  assign new_P1_R1192_U203 = ~new_P1_U3067 | ~new_P1_R1192_U32;
  assign new_P1_R1192_U204 = ~new_P1_R1192_U188 | ~new_P1_R1192_U6;
  assign new_P1_R1192_U205 = ~new_P1_R1192_U7 | ~new_P1_R1192_U204;
  assign new_P1_R1192_U206 = ~new_P1_U3470 | ~new_P1_R1192_U36;
  assign new_P1_R1192_U207 = ~new_P1_U3476 | ~new_P1_R1192_U34;
  assign new_P1_R1192_U208 = ~new_P1_R1192_U6 | ~new_P1_R1192_U206 | ~new_P1_R1192_U152;
  assign new_P1_R1192_U209 = ~new_P1_R1192_U207 | ~new_P1_R1192_U205;
  assign new_P1_R1192_U210 = ~new_P1_R1192_U44;
  assign new_P1_R1192_U211 = ~new_P1_U3482 | ~new_P1_R1192_U41;
  assign new_P1_R1192_U212 = ~new_P1_R1192_U117 | ~new_P1_R1192_U44;
  assign new_P1_R1192_U213 = ~new_P1_R1192_U41 | ~new_P1_R1192_U40;
  assign new_P1_R1192_U214 = ~new_P1_R1192_U213 | ~new_P1_R1192_U38;
  assign new_P1_R1192_U215 = ~new_P1_U3084 | ~new_P1_R1192_U178;
  assign new_P1_R1192_U216 = ~new_P1_R1192_U148;
  assign new_P1_R1192_U217 = ~new_P1_U3485 | ~new_P1_R1192_U43;
  assign new_P1_R1192_U218 = ~new_P1_R1192_U217 | ~new_P1_R1192_U54;
  assign new_P1_R1192_U219 = ~new_P1_R1192_U210 | ~new_P1_R1192_U40;
  assign new_P1_R1192_U220 = ~new_P1_R1192_U120 | ~new_P1_R1192_U219;
  assign new_P1_R1192_U221 = ~new_P1_R1192_U44 | ~new_P1_R1192_U185;
  assign new_P1_R1192_U222 = ~new_P1_R1192_U119 | ~new_P1_R1192_U221;
  assign new_P1_R1192_U223 = ~new_P1_R1192_U40 | ~new_P1_R1192_U185;
  assign new_P1_R1192_U224 = ~new_P1_R1192_U206 | ~new_P1_R1192_U152;
  assign new_P1_R1192_U225 = ~new_P1_R1192_U45;
  assign new_P1_R1192_U226 = ~new_P1_U3067 | ~new_P1_R1192_U32;
  assign new_P1_R1192_U227 = ~new_P1_R1192_U225 | ~new_P1_R1192_U226;
  assign new_P1_R1192_U228 = ~new_P1_R1192_U122 | ~new_P1_R1192_U227;
  assign new_P1_R1192_U229 = ~new_P1_R1192_U45 | ~new_P1_R1192_U184;
  assign new_P1_R1192_U230 = ~new_P1_U3476 | ~new_P1_R1192_U34;
  assign new_P1_R1192_U231 = ~new_P1_R1192_U121 | ~new_P1_R1192_U229;
  assign new_P1_R1192_U232 = ~new_P1_U3067 | ~new_P1_R1192_U32;
  assign new_P1_R1192_U233 = ~new_P1_R1192_U184 | ~new_P1_R1192_U232;
  assign new_P1_R1192_U234 = ~new_P1_R1192_U206 | ~new_P1_R1192_U37;
  assign new_P1_R1192_U235 = ~new_P1_R1192_U194 | ~new_P1_R1192_U29;
  assign new_P1_R1192_U236 = ~new_P1_R1192_U124 | ~new_P1_R1192_U235;
  assign new_P1_R1192_U237 = ~new_P1_R1192_U46 | ~new_P1_R1192_U183;
  assign new_P1_R1192_U238 = ~new_P1_R1192_U123 | ~new_P1_R1192_U237;
  assign new_P1_R1192_U239 = ~new_P1_R1192_U29 | ~new_P1_R1192_U183;
  assign new_P1_R1192_U240 = ~new_P1_U3491 | ~new_P1_R1192_U52;
  assign new_P1_R1192_U241 = ~new_P1_U3063 | ~new_P1_R1192_U50;
  assign new_P1_R1192_U242 = ~new_P1_U3062 | ~new_P1_R1192_U51;
  assign new_P1_R1192_U243 = ~new_P1_R1192_U189 | ~new_P1_R1192_U8;
  assign new_P1_R1192_U244 = ~new_P1_R1192_U9 | ~new_P1_R1192_U243;
  assign new_P1_R1192_U245 = ~new_P1_U3491 | ~new_P1_R1192_U52;
  assign new_P1_R1192_U246 = ~new_P1_R1192_U125 | ~new_P1_R1192_U148;
  assign new_P1_R1192_U247 = ~new_P1_R1192_U245 | ~new_P1_R1192_U244;
  assign new_P1_R1192_U248 = ~new_P1_R1192_U173;
  assign new_P1_R1192_U249 = ~new_P1_U3494 | ~new_P1_R1192_U56;
  assign new_P1_R1192_U250 = ~new_P1_R1192_U249 | ~new_P1_R1192_U173;
  assign new_P1_R1192_U251 = ~new_P1_U3072 | ~new_P1_R1192_U55;
  assign new_P1_R1192_U252 = ~new_P1_R1192_U172;
  assign new_P1_R1192_U253 = ~new_P1_U3497 | ~new_P1_R1192_U58;
  assign new_P1_R1192_U254 = ~new_P1_R1192_U253 | ~new_P1_R1192_U172;
  assign new_P1_R1192_U255 = ~new_P1_U3080 | ~new_P1_R1192_U57;
  assign new_P1_R1192_U256 = ~new_P1_R1192_U171;
  assign new_P1_R1192_U257 = ~new_P1_U3506 | ~new_P1_R1192_U61;
  assign new_P1_R1192_U258 = ~new_P1_U3073 | ~new_P1_R1192_U59;
  assign new_P1_R1192_U259 = ~new_P1_U3074 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U260 = ~new_P1_R1192_U186 | ~new_P1_R1192_U180;
  assign new_P1_R1192_U261 = ~new_P1_R1192_U10 | ~new_P1_R1192_U260;
  assign new_P1_R1192_U262 = ~new_P1_U3500 | ~new_P1_R1192_U63;
  assign new_P1_R1192_U263 = ~new_P1_U3506 | ~new_P1_R1192_U61;
  assign new_P1_R1192_U264 = ~new_P1_R1192_U257 | ~new_P1_R1192_U171 | ~new_P1_R1192_U126;
  assign new_P1_R1192_U265 = ~new_P1_R1192_U263 | ~new_P1_R1192_U261;
  assign new_P1_R1192_U266 = ~new_P1_R1192_U168;
  assign new_P1_R1192_U267 = ~new_P1_U3509 | ~new_P1_R1192_U66;
  assign new_P1_R1192_U268 = ~new_P1_R1192_U267 | ~new_P1_R1192_U168;
  assign new_P1_R1192_U269 = ~new_P1_U3069 | ~new_P1_R1192_U65;
  assign new_P1_R1192_U270 = ~new_P1_R1192_U67;
  assign new_P1_R1192_U271 = ~new_P1_R1192_U270 | ~new_P1_R1192_U68;
  assign new_P1_R1192_U272 = ~new_P1_R1192_U271 | ~new_P1_R1192_U167;
  assign new_P1_R1192_U273 = ~new_P1_U3082 | ~new_P1_R1192_U67;
  assign new_P1_R1192_U274 = ~new_P1_R1192_U166;
  assign new_P1_R1192_U275 = ~new_P1_U3514 | ~new_P1_R1192_U70;
  assign new_P1_R1192_U276 = ~new_P1_R1192_U275 | ~new_P1_R1192_U166;
  assign new_P1_R1192_U277 = ~new_P1_U3081 | ~new_P1_R1192_U69;
  assign new_P1_R1192_U278 = ~new_P1_R1192_U164;
  assign new_P1_R1192_U279 = ~new_P1_U4025 | ~new_P1_R1192_U72;
  assign new_P1_R1192_U280 = ~new_P1_R1192_U279 | ~new_P1_R1192_U164;
  assign new_P1_R1192_U281 = ~new_P1_U3076 | ~new_P1_R1192_U71;
  assign new_P1_R1192_U282 = ~new_P1_R1192_U163;
  assign new_P1_R1192_U283 = ~new_P1_U4022 | ~new_P1_R1192_U75;
  assign new_P1_R1192_U284 = ~new_P1_U3066 | ~new_P1_R1192_U73;
  assign new_P1_R1192_U285 = ~new_P1_U3061 | ~new_P1_R1192_U48;
  assign new_P1_R1192_U286 = ~new_P1_R1192_U187 | ~new_P1_R1192_U181;
  assign new_P1_R1192_U287 = ~new_P1_R1192_U11 | ~new_P1_R1192_U286;
  assign new_P1_R1192_U288 = ~new_P1_U4024 | ~new_P1_R1192_U77;
  assign new_P1_R1192_U289 = ~new_P1_U4022 | ~new_P1_R1192_U75;
  assign new_P1_R1192_U290 = ~new_P1_R1192_U283 | ~new_P1_R1192_U163 | ~new_P1_R1192_U127;
  assign new_P1_R1192_U291 = ~new_P1_R1192_U289 | ~new_P1_R1192_U287;
  assign new_P1_R1192_U292 = ~new_P1_R1192_U160;
  assign new_P1_R1192_U293 = ~new_P1_U4021 | ~new_P1_R1192_U80;
  assign new_P1_R1192_U294 = ~new_P1_R1192_U293 | ~new_P1_R1192_U160;
  assign new_P1_R1192_U295 = ~new_P1_U3065 | ~new_P1_R1192_U79;
  assign new_P1_R1192_U296 = ~new_P1_R1192_U159;
  assign new_P1_R1192_U297 = ~new_P1_U4020 | ~new_P1_R1192_U82;
  assign new_P1_R1192_U298 = ~new_P1_R1192_U297 | ~new_P1_R1192_U159;
  assign new_P1_R1192_U299 = ~new_P1_U3058 | ~new_P1_R1192_U81;
  assign new_P1_R1192_U300 = ~new_P1_R1192_U89;
  assign new_P1_R1192_U301 = ~new_P1_U4018 | ~new_P1_R1192_U86;
  assign new_P1_R1192_U302 = ~new_P1_R1192_U301 | ~new_P1_R1192_U89 | ~new_P1_R1192_U182;
  assign new_P1_R1192_U303 = ~new_P1_R1192_U86 | ~new_P1_R1192_U85;
  assign new_P1_R1192_U304 = ~new_P1_R1192_U303 | ~new_P1_R1192_U83;
  assign new_P1_R1192_U305 = ~new_P1_U3053 | ~new_P1_R1192_U176;
  assign new_P1_R1192_U306 = ~new_P1_R1192_U157;
  assign new_P1_R1192_U307 = ~new_P1_U4017 | ~new_P1_R1192_U88;
  assign new_P1_R1192_U308 = ~new_P1_U3054 | ~new_P1_R1192_U87;
  assign new_P1_R1192_U309 = ~new_P1_R1192_U300 | ~new_P1_R1192_U85;
  assign new_P1_R1192_U310 = ~new_P1_R1192_U133 | ~new_P1_R1192_U309;
  assign new_P1_R1192_U311 = ~new_P1_R1192_U89 | ~new_P1_R1192_U182;
  assign new_P1_R1192_U312 = ~new_P1_R1192_U132 | ~new_P1_R1192_U311;
  assign new_P1_R1192_U313 = ~new_P1_R1192_U85 | ~new_P1_R1192_U182;
  assign new_P1_R1192_U314 = ~new_P1_R1192_U288 | ~new_P1_R1192_U163;
  assign new_P1_R1192_U315 = ~new_P1_R1192_U90;
  assign new_P1_R1192_U316 = ~new_P1_U3061 | ~new_P1_R1192_U48;
  assign new_P1_R1192_U317 = ~new_P1_R1192_U315 | ~new_P1_R1192_U316;
  assign new_P1_R1192_U318 = ~new_P1_R1192_U136 | ~new_P1_R1192_U317;
  assign new_P1_R1192_U319 = ~new_P1_R1192_U90 | ~new_P1_R1192_U181;
  assign new_P1_R1192_U320 = ~new_P1_U4022 | ~new_P1_R1192_U75;
  assign new_P1_R1192_U321 = ~new_P1_R1192_U11 | ~new_P1_R1192_U320 | ~new_P1_R1192_U319;
  assign new_P1_R1192_U322 = ~new_P1_U3061 | ~new_P1_R1192_U48;
  assign new_P1_R1192_U323 = ~new_P1_R1192_U181 | ~new_P1_R1192_U322;
  assign new_P1_R1192_U324 = ~new_P1_R1192_U288 | ~new_P1_R1192_U78;
  assign new_P1_R1192_U325 = ~new_P1_R1192_U262 | ~new_P1_R1192_U171;
  assign new_P1_R1192_U326 = ~new_P1_R1192_U91;
  assign new_P1_R1192_U327 = ~new_P1_U3074 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U328 = ~new_P1_R1192_U326 | ~new_P1_R1192_U327;
  assign new_P1_R1192_U329 = ~new_P1_R1192_U142 | ~new_P1_R1192_U328;
  assign new_P1_R1192_U330 = ~new_P1_R1192_U91 | ~new_P1_R1192_U180;
  assign new_P1_R1192_U331 = ~new_P1_U3506 | ~new_P1_R1192_U61;
  assign new_P1_R1192_U332 = ~new_P1_R1192_U10 | ~new_P1_R1192_U331 | ~new_P1_R1192_U330;
  assign new_P1_R1192_U333 = ~new_P1_U3074 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U334 = ~new_P1_R1192_U180 | ~new_P1_R1192_U333;
  assign new_P1_R1192_U335 = ~new_P1_R1192_U262 | ~new_P1_R1192_U64;
  assign new_P1_R1192_U336 = ~new_P1_R1192_U217 | ~new_P1_R1192_U148;
  assign new_P1_R1192_U337 = ~new_P1_R1192_U92;
  assign new_P1_R1192_U338 = ~new_P1_U3062 | ~new_P1_R1192_U51;
  assign new_P1_R1192_U339 = ~new_P1_R1192_U337 | ~new_P1_R1192_U338;
  assign new_P1_R1192_U340 = ~new_P1_R1192_U146 | ~new_P1_R1192_U339;
  assign new_P1_R1192_U341 = ~new_P1_R1192_U92 | ~new_P1_R1192_U179;
  assign new_P1_R1192_U342 = ~new_P1_U3491 | ~new_P1_R1192_U52;
  assign new_P1_R1192_U343 = ~new_P1_R1192_U145 | ~new_P1_R1192_U341;
  assign new_P1_R1192_U344 = ~new_P1_U3062 | ~new_P1_R1192_U51;
  assign new_P1_R1192_U345 = ~new_P1_R1192_U179 | ~new_P1_R1192_U344;
  assign new_P1_R1192_U346 = ~new_P1_U3077 | ~new_P1_R1192_U24;
  assign new_P1_R1192_U347 = ~new_P1_R1192_U301 | ~new_P1_R1192_U89 | ~new_P1_R1192_U182;
  assign new_P1_R1192_U348 = ~new_P1_R1192_U130 | ~new_P1_R1192_U12 | ~new_P1_R1192_U347;
  assign new_P1_R1192_U349 = ~new_P1_U3485 | ~new_P1_R1192_U43;
  assign new_P1_R1192_U350 = ~new_P1_U3083 | ~new_P1_R1192_U42;
  assign new_P1_R1192_U351 = ~new_P1_R1192_U218 | ~new_P1_R1192_U148;
  assign new_P1_R1192_U352 = ~new_P1_R1192_U216 | ~new_P1_R1192_U147;
  assign new_P1_R1192_U353 = ~new_P1_U3482 | ~new_P1_R1192_U41;
  assign new_P1_R1192_U354 = ~new_P1_U3084 | ~new_P1_R1192_U38;
  assign new_P1_R1192_U355 = ~new_P1_U3482 | ~new_P1_R1192_U41;
  assign new_P1_R1192_U356 = ~new_P1_U3084 | ~new_P1_R1192_U38;
  assign new_P1_R1192_U357 = ~new_P1_R1192_U356 | ~new_P1_R1192_U355;
  assign new_P1_R1192_U358 = ~new_P1_U3479 | ~new_P1_R1192_U39;
  assign new_P1_R1192_U359 = ~new_P1_U3070 | ~new_P1_R1192_U22;
  assign new_P1_R1192_U360 = ~new_P1_R1192_U223 | ~new_P1_R1192_U44;
  assign new_P1_R1192_U361 = ~new_P1_R1192_U149 | ~new_P1_R1192_U210;
  assign new_P1_R1192_U362 = ~new_P1_U3476 | ~new_P1_R1192_U34;
  assign new_P1_R1192_U363 = ~new_P1_U3071 | ~new_P1_R1192_U31;
  assign new_P1_R1192_U364 = ~new_P1_R1192_U363 | ~new_P1_R1192_U362;
  assign new_P1_R1192_U365 = ~new_P1_U3473 | ~new_P1_R1192_U35;
  assign new_P1_R1192_U366 = ~new_P1_U3067 | ~new_P1_R1192_U32;
  assign new_P1_R1192_U367 = ~new_P1_R1192_U233 | ~new_P1_R1192_U45;
  assign new_P1_R1192_U368 = ~new_P1_R1192_U150 | ~new_P1_R1192_U225;
  assign new_P1_R1192_U369 = ~new_P1_U3470 | ~new_P1_R1192_U36;
  assign new_P1_R1192_U370 = ~new_P1_U3060 | ~new_P1_R1192_U33;
  assign new_P1_R1192_U371 = ~new_P1_R1192_U234 | ~new_P1_R1192_U152;
  assign new_P1_R1192_U372 = ~new_P1_R1192_U200 | ~new_P1_R1192_U151;
  assign new_P1_R1192_U373 = ~new_P1_U3467 | ~new_P1_R1192_U30;
  assign new_P1_R1192_U374 = ~new_P1_U3064 | ~new_P1_R1192_U27;
  assign new_P1_R1192_U375 = ~new_P1_U3467 | ~new_P1_R1192_U30;
  assign new_P1_R1192_U376 = ~new_P1_U3064 | ~new_P1_R1192_U27;
  assign new_P1_R1192_U377 = ~new_P1_R1192_U376 | ~new_P1_R1192_U375;
  assign new_P1_R1192_U378 = ~new_P1_U3464 | ~new_P1_R1192_U28;
  assign new_P1_R1192_U379 = ~new_P1_U3068 | ~new_P1_R1192_U23;
  assign new_P1_R1192_U380 = ~new_P1_R1192_U239 | ~new_P1_R1192_U46;
  assign new_P1_R1192_U381 = ~new_P1_R1192_U153 | ~new_P1_R1192_U194;
  assign new_P1_R1192_U382 = ~new_P1_U4028 | ~new_P1_R1192_U155;
  assign new_P1_R1192_U383 = ~new_P1_U3055 | ~new_P1_R1192_U154;
  assign new_P1_R1192_U384 = ~new_P1_U4028 | ~new_P1_R1192_U155;
  assign new_P1_R1192_U385 = ~new_P1_U3055 | ~new_P1_R1192_U154;
  assign new_P1_R1192_U386 = ~new_P1_R1192_U385 | ~new_P1_R1192_U384;
  assign new_P1_R1192_U387 = ~new_P1_R1192_U87 | ~new_P1_U3054 | ~new_P1_R1192_U386;
  assign new_P1_R1192_U388 = ~new_P1_U4017 | ~new_P1_R1192_U12 | ~new_P1_R1192_U88;
  assign new_P1_R1192_U389 = ~new_P1_U4017 | ~new_P1_R1192_U88;
  assign new_P1_R1192_U390 = ~new_P1_U3054 | ~new_P1_R1192_U87;
  assign new_P1_R1192_U391 = ~new_P1_R1192_U131;
  assign new_P1_R1192_U392 = ~new_P1_R1192_U306 | ~new_P1_R1192_U391;
  assign new_P1_R1192_U393 = ~new_P1_R1192_U131 | ~new_P1_R1192_U157;
  assign new_P1_R1192_U394 = ~new_P1_U4018 | ~new_P1_R1192_U86;
  assign new_P1_R1192_U395 = ~new_P1_U3053 | ~new_P1_R1192_U83;
  assign new_P1_R1192_U396 = ~new_P1_U4018 | ~new_P1_R1192_U86;
  assign new_P1_R1192_U397 = ~new_P1_U3053 | ~new_P1_R1192_U83;
  assign new_P1_R1192_U398 = ~new_P1_R1192_U397 | ~new_P1_R1192_U396;
  assign new_P1_R1192_U399 = ~new_P1_U4019 | ~new_P1_R1192_U84;
  assign new_P1_R1192_U400 = ~new_P1_U3057 | ~new_P1_R1192_U47;
  assign new_P1_R1192_U401 = ~new_P1_R1192_U313 | ~new_P1_R1192_U89;
  assign new_P1_R1192_U402 = ~new_P1_R1192_U158 | ~new_P1_R1192_U300;
  assign new_P1_R1192_U403 = ~new_P1_U4020 | ~new_P1_R1192_U82;
  assign new_P1_R1192_U404 = ~new_P1_U3058 | ~new_P1_R1192_U81;
  assign new_P1_R1192_U405 = ~new_P1_R1192_U134;
  assign new_P1_R1192_U406 = ~new_P1_R1192_U296 | ~new_P1_R1192_U405;
  assign new_P1_R1192_U407 = ~new_P1_R1192_U134 | ~new_P1_R1192_U159;
  assign new_P1_R1192_U408 = ~new_P1_U4021 | ~new_P1_R1192_U80;
  assign new_P1_R1192_U409 = ~new_P1_U3065 | ~new_P1_R1192_U79;
  assign new_P1_R1192_U410 = ~new_P1_R1192_U135;
  assign new_P1_R1192_U411 = ~new_P1_R1192_U292 | ~new_P1_R1192_U410;
  assign new_P1_R1192_U412 = ~new_P1_R1192_U135 | ~new_P1_R1192_U160;
  assign new_P1_R1192_U413 = ~new_P1_U4022 | ~new_P1_R1192_U75;
  assign new_P1_R1192_U414 = ~new_P1_U3066 | ~new_P1_R1192_U73;
  assign new_P1_R1192_U415 = ~new_P1_R1192_U414 | ~new_P1_R1192_U413;
  assign new_P1_R1192_U416 = ~new_P1_U4023 | ~new_P1_R1192_U76;
  assign new_P1_R1192_U417 = ~new_P1_U3061 | ~new_P1_R1192_U48;
  assign new_P1_R1192_U418 = ~new_P1_R1192_U323 | ~new_P1_R1192_U90;
  assign new_P1_R1192_U419 = ~new_P1_R1192_U161 | ~new_P1_R1192_U315;
  assign new_P1_R1192_U420 = ~new_P1_U4024 | ~new_P1_R1192_U77;
  assign new_P1_R1192_U421 = ~new_P1_U3075 | ~new_P1_R1192_U74;
  assign new_P1_R1192_U422 = ~new_P1_R1192_U324 | ~new_P1_R1192_U163;
  assign new_P1_R1192_U423 = ~new_P1_R1192_U282 | ~new_P1_R1192_U162;
  assign new_P1_R1192_U424 = ~new_P1_U4025 | ~new_P1_R1192_U72;
  assign new_P1_R1192_U425 = ~new_P1_U3076 | ~new_P1_R1192_U71;
  assign new_P1_R1192_U426 = ~new_P1_R1192_U137;
  assign new_P1_R1192_U427 = ~new_P1_R1192_U278 | ~new_P1_R1192_U426;
  assign new_P1_R1192_U428 = ~new_P1_R1192_U137 | ~new_P1_R1192_U164;
  assign new_P1_R1192_U429 = ~new_P1_U3461 | ~new_P1_R1192_U26;
  assign new_P1_R1192_U430 = ~new_P1_U3078 | ~new_P1_R1192_U165;
  assign new_P1_R1192_U431 = ~new_P1_R1192_U138;
  assign new_P1_R1192_U432 = ~new_P1_R1192_U431 | ~new_P1_R1192_U190;
  assign new_P1_R1192_U433 = ~new_P1_R1192_U138 | ~new_P1_R1192_U25;
  assign new_P1_R1192_U434 = ~new_P1_U3514 | ~new_P1_R1192_U70;
  assign new_P1_R1192_U435 = ~new_P1_U3081 | ~new_P1_R1192_U69;
  assign new_P1_R1192_U436 = ~new_P1_R1192_U139;
  assign new_P1_R1192_U437 = ~new_P1_R1192_U274 | ~new_P1_R1192_U436;
  assign new_P1_R1192_U438 = ~new_P1_R1192_U139 | ~new_P1_R1192_U166;
  assign new_P1_R1192_U439 = ~new_P1_U3512 | ~new_P1_R1192_U68;
  assign new_P1_R1192_U440 = ~new_P1_U3082 | ~new_P1_R1192_U167;
  assign new_P1_R1192_U441 = ~new_P1_R1192_U140;
  assign new_P1_R1192_U442 = ~new_P1_R1192_U441 | ~new_P1_R1192_U270;
  assign new_P1_R1192_U443 = ~new_P1_R1192_U140 | ~new_P1_R1192_U67;
  assign new_P1_R1192_U444 = ~new_P1_U3509 | ~new_P1_R1192_U66;
  assign new_P1_R1192_U445 = ~new_P1_U3069 | ~new_P1_R1192_U65;
  assign new_P1_R1192_U446 = ~new_P1_R1192_U141;
  assign new_P1_R1192_U447 = ~new_P1_R1192_U266 | ~new_P1_R1192_U446;
  assign new_P1_R1192_U448 = ~new_P1_R1192_U141 | ~new_P1_R1192_U168;
  assign new_P1_R1192_U449 = ~new_P1_U3506 | ~new_P1_R1192_U61;
  assign new_P1_R1192_U450 = ~new_P1_U3073 | ~new_P1_R1192_U59;
  assign new_P1_R1192_U451 = ~new_P1_R1192_U450 | ~new_P1_R1192_U449;
  assign new_P1_R1192_U452 = ~new_P1_U3503 | ~new_P1_R1192_U62;
  assign new_P1_R1192_U453 = ~new_P1_U3074 | ~new_P1_R1192_U49;
  assign new_P1_R1192_U454 = ~new_P1_R1192_U334 | ~new_P1_R1192_U91;
  assign new_P1_R1192_U455 = ~new_P1_R1192_U169 | ~new_P1_R1192_U326;
  assign new_P1_R1192_U456 = ~new_P1_U3500 | ~new_P1_R1192_U63;
  assign new_P1_R1192_U457 = ~new_P1_U3079 | ~new_P1_R1192_U60;
  assign new_P1_R1192_U458 = ~new_P1_R1192_U335 | ~new_P1_R1192_U171;
  assign new_P1_R1192_U459 = ~new_P1_R1192_U256 | ~new_P1_R1192_U170;
  assign new_P1_R1192_U460 = ~new_P1_U3497 | ~new_P1_R1192_U58;
  assign new_P1_R1192_U461 = ~new_P1_U3080 | ~new_P1_R1192_U57;
  assign new_P1_R1192_U462 = ~new_P1_R1192_U143;
  assign new_P1_R1192_U463 = ~new_P1_R1192_U252 | ~new_P1_R1192_U462;
  assign new_P1_R1192_U464 = ~new_P1_R1192_U143 | ~new_P1_R1192_U172;
  assign new_P1_R1192_U465 = ~new_P1_U3494 | ~new_P1_R1192_U56;
  assign new_P1_R1192_U466 = ~new_P1_U3072 | ~new_P1_R1192_U55;
  assign new_P1_R1192_U467 = ~new_P1_R1192_U144;
  assign new_P1_R1192_U468 = ~new_P1_R1192_U248 | ~new_P1_R1192_U467;
  assign new_P1_R1192_U469 = ~new_P1_R1192_U144 | ~new_P1_R1192_U173;
  assign new_P1_R1192_U470 = ~new_P1_U3491 | ~new_P1_R1192_U52;
  assign new_P1_R1192_U471 = ~new_P1_U3063 | ~new_P1_R1192_U50;
  assign new_P1_R1192_U472 = ~new_P1_R1192_U471 | ~new_P1_R1192_U470;
  assign new_P1_R1192_U473 = ~new_P1_U3488 | ~new_P1_R1192_U53;
  assign new_P1_R1192_U474 = ~new_P1_U3062 | ~new_P1_R1192_U51;
  assign new_P1_R1192_U475 = ~new_P1_R1192_U345 | ~new_P1_R1192_U92;
  assign new_P1_R1192_U476 = ~new_P1_R1192_U174 | ~new_P1_R1192_U337;
  assign new_P1_R1171_U4 = new_P1_R1171_U176 & new_P1_R1171_U175;
  assign new_P1_R1171_U5 = new_P1_R1171_U177 & new_P1_R1171_U178;
  assign new_P1_R1171_U6 = new_P1_R1171_U194 & new_P1_R1171_U193;
  assign new_P1_R1171_U7 = new_P1_R1171_U234 & new_P1_R1171_U233;
  assign new_P1_R1171_U8 = new_P1_R1171_U243 & new_P1_R1171_U242;
  assign new_P1_R1171_U9 = new_P1_R1171_U261 & new_P1_R1171_U260;
  assign new_P1_R1171_U10 = new_P1_R1171_U269 & new_P1_R1171_U268;
  assign new_P1_R1171_U11 = new_P1_R1171_U348 & new_P1_R1171_U345;
  assign new_P1_R1171_U12 = new_P1_R1171_U341 & new_P1_R1171_U338;
  assign new_P1_R1171_U13 = new_P1_R1171_U332 & new_P1_R1171_U329;
  assign new_P1_R1171_U14 = new_P1_R1171_U323 & new_P1_R1171_U320;
  assign new_P1_R1171_U15 = new_P1_R1171_U317 & new_P1_R1171_U315;
  assign new_P1_R1171_U16 = new_P1_R1171_U310 & new_P1_R1171_U307;
  assign new_P1_R1171_U17 = new_P1_R1171_U232 & new_P1_R1171_U229;
  assign new_P1_R1171_U18 = new_P1_R1171_U224 & new_P1_R1171_U221;
  assign new_P1_R1171_U19 = new_P1_R1171_U210 & new_P1_R1171_U207;
  assign new_P1_R1171_U20 = ~new_P1_U3476;
  assign new_P1_R1171_U21 = ~new_P1_U3071;
  assign new_P1_R1171_U22 = ~new_P1_U3070;
  assign new_P1_R1171_U23 = ~new_P1_U3071 | ~new_P1_U3476;
  assign new_P1_R1171_U24 = ~new_P1_U3479;
  assign new_P1_R1171_U25 = ~new_P1_U3470;
  assign new_P1_R1171_U26 = ~new_P1_U3060;
  assign new_P1_R1171_U27 = ~new_P1_U3067;
  assign new_P1_R1171_U28 = ~new_P1_U3464;
  assign new_P1_R1171_U29 = ~new_P1_U3068;
  assign new_P1_R1171_U30 = ~new_P1_U3456;
  assign new_P1_R1171_U31 = ~new_P1_U3077;
  assign new_P1_R1171_U32 = ~new_P1_U3077 | ~new_P1_U3456;
  assign new_P1_R1171_U33 = ~new_P1_U3467;
  assign new_P1_R1171_U34 = ~new_P1_U3064;
  assign new_P1_R1171_U35 = ~new_P1_U3060 | ~new_P1_U3470;
  assign new_P1_R1171_U36 = ~new_P1_U3473;
  assign new_P1_R1171_U37 = ~new_P1_U3482;
  assign new_P1_R1171_U38 = ~new_P1_U3084;
  assign new_P1_R1171_U39 = ~new_P1_U3083;
  assign new_P1_R1171_U40 = ~new_P1_U3485;
  assign new_P1_R1171_U41 = ~new_P1_R1171_U62 | ~new_P1_R1171_U202;
  assign new_P1_R1171_U42 = ~new_P1_R1171_U118 | ~new_P1_R1171_U190;
  assign new_P1_R1171_U43 = ~new_P1_R1171_U179 | ~new_P1_R1171_U180;
  assign new_P1_R1171_U44 = ~new_P1_U3461 | ~new_P1_U3078;
  assign new_P1_R1171_U45 = ~new_P1_R1171_U122 | ~new_P1_R1171_U216;
  assign new_P1_R1171_U46 = ~new_P1_R1171_U213 | ~new_P1_R1171_U212;
  assign new_P1_R1171_U47 = ~new_P1_U4018;
  assign new_P1_R1171_U48 = ~new_P1_U3053;
  assign new_P1_R1171_U49 = ~new_P1_U3057;
  assign new_P1_R1171_U50 = ~new_P1_U4019;
  assign new_P1_R1171_U51 = ~new_P1_U4020;
  assign new_P1_R1171_U52 = ~new_P1_U3058;
  assign new_P1_R1171_U53 = ~new_P1_U4021;
  assign new_P1_R1171_U54 = ~new_P1_U3065;
  assign new_P1_R1171_U55 = ~new_P1_U4024;
  assign new_P1_R1171_U56 = ~new_P1_U3075;
  assign new_P1_R1171_U57 = ~new_P1_U3506;
  assign new_P1_R1171_U58 = ~new_P1_U3073;
  assign new_P1_R1171_U59 = ~new_P1_U3069;
  assign new_P1_R1171_U60 = ~new_P1_U3073 | ~new_P1_U3506;
  assign new_P1_R1171_U61 = ~new_P1_U3509;
  assign new_P1_R1171_U62 = ~new_P1_U3084 | ~new_P1_U3482;
  assign new_P1_R1171_U63 = ~new_P1_U3488;
  assign new_P1_R1171_U64 = ~new_P1_U3062;
  assign new_P1_R1171_U65 = ~new_P1_U3494;
  assign new_P1_R1171_U66 = ~new_P1_U3072;
  assign new_P1_R1171_U67 = ~new_P1_U3491;
  assign new_P1_R1171_U68 = ~new_P1_U3063;
  assign new_P1_R1171_U69 = ~new_P1_U3063 | ~new_P1_U3491;
  assign new_P1_R1171_U70 = ~new_P1_U3497;
  assign new_P1_R1171_U71 = ~new_P1_U3080;
  assign new_P1_R1171_U72 = ~new_P1_U3500;
  assign new_P1_R1171_U73 = ~new_P1_U3079;
  assign new_P1_R1171_U74 = ~new_P1_U3503;
  assign new_P1_R1171_U75 = ~new_P1_U3074;
  assign new_P1_R1171_U76 = ~new_P1_U3512;
  assign new_P1_R1171_U77 = ~new_P1_U3082;
  assign new_P1_R1171_U78 = ~new_P1_U3082 | ~new_P1_U3512;
  assign new_P1_R1171_U79 = ~new_P1_U3514;
  assign new_P1_R1171_U80 = ~new_P1_U3081;
  assign new_P1_R1171_U81 = ~new_P1_U3081 | ~new_P1_U3514;
  assign new_P1_R1171_U82 = ~new_P1_U4025;
  assign new_P1_R1171_U83 = ~new_P1_U4023;
  assign new_P1_R1171_U84 = ~new_P1_U3061;
  assign new_P1_R1171_U85 = ~new_P1_U4022;
  assign new_P1_R1171_U86 = ~new_P1_U3066;
  assign new_P1_R1171_U87 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1171_U88 = ~new_P1_U3054;
  assign new_P1_R1171_U89 = ~new_P1_U4017;
  assign new_P1_R1171_U90 = ~new_P1_R1171_U303 | ~new_P1_R1171_U173;
  assign new_P1_R1171_U91 = ~new_P1_U3076;
  assign new_P1_R1171_U92 = ~new_P1_R1171_U78 | ~new_P1_R1171_U312;
  assign new_P1_R1171_U93 = ~new_P1_R1171_U258 | ~new_P1_R1171_U257;
  assign new_P1_R1171_U94 = ~new_P1_R1171_U69 | ~new_P1_R1171_U334;
  assign new_P1_R1171_U95 = ~new_P1_R1171_U454 | ~new_P1_R1171_U453;
  assign new_P1_R1171_U96 = ~new_P1_R1171_U501 | ~new_P1_R1171_U500;
  assign new_P1_R1171_U97 = ~new_P1_R1171_U372 | ~new_P1_R1171_U371;
  assign new_P1_R1171_U98 = ~new_P1_R1171_U377 | ~new_P1_R1171_U376;
  assign new_P1_R1171_U99 = ~new_P1_R1171_U384 | ~new_P1_R1171_U383;
  assign new_P1_R1171_U100 = ~new_P1_R1171_U391 | ~new_P1_R1171_U390;
  assign new_P1_R1171_U101 = ~new_P1_R1171_U396 | ~new_P1_R1171_U395;
  assign new_P1_R1171_U102 = ~new_P1_R1171_U405 | ~new_P1_R1171_U404;
  assign new_P1_R1171_U103 = ~new_P1_R1171_U412 | ~new_P1_R1171_U411;
  assign new_P1_R1171_U104 = ~new_P1_R1171_U419 | ~new_P1_R1171_U418;
  assign new_P1_R1171_U105 = ~new_P1_R1171_U426 | ~new_P1_R1171_U425;
  assign new_P1_R1171_U106 = ~new_P1_R1171_U431 | ~new_P1_R1171_U430;
  assign new_P1_R1171_U107 = ~new_P1_R1171_U438 | ~new_P1_R1171_U437;
  assign new_P1_R1171_U108 = ~new_P1_R1171_U445 | ~new_P1_R1171_U444;
  assign new_P1_R1171_U109 = ~new_P1_R1171_U459 | ~new_P1_R1171_U458;
  assign new_P1_R1171_U110 = ~new_P1_R1171_U464 | ~new_P1_R1171_U463;
  assign new_P1_R1171_U111 = ~new_P1_R1171_U471 | ~new_P1_R1171_U470;
  assign new_P1_R1171_U112 = ~new_P1_R1171_U478 | ~new_P1_R1171_U477;
  assign new_P1_R1171_U113 = ~new_P1_R1171_U485 | ~new_P1_R1171_U484;
  assign new_P1_R1171_U114 = ~new_P1_R1171_U492 | ~new_P1_R1171_U491;
  assign new_P1_R1171_U115 = ~new_P1_R1171_U497 | ~new_P1_R1171_U496;
  assign new_P1_R1171_U116 = new_P1_U3464 & new_P1_U3068;
  assign new_P1_R1171_U117 = new_P1_R1171_U186 & new_P1_R1171_U184;
  assign new_P1_R1171_U118 = new_P1_R1171_U191 & new_P1_R1171_U189;
  assign new_P1_R1171_U119 = new_P1_R1171_U198 & new_P1_R1171_U197;
  assign new_P1_R1171_U120 = new_P1_R1171_U23 & new_P1_R1171_U379 & new_P1_R1171_U378;
  assign new_P1_R1171_U121 = new_P1_R1171_U209 & new_P1_R1171_U6;
  assign new_P1_R1171_U122 = new_P1_R1171_U217 & new_P1_R1171_U215;
  assign new_P1_R1171_U123 = new_P1_R1171_U35 & new_P1_R1171_U386 & new_P1_R1171_U385;
  assign new_P1_R1171_U124 = new_P1_R1171_U223 & new_P1_R1171_U4;
  assign new_P1_R1171_U125 = new_P1_R1171_U231 & new_P1_R1171_U178;
  assign new_P1_R1171_U126 = new_P1_R1171_U201 & new_P1_R1171_U7;
  assign new_P1_R1171_U127 = new_P1_R1171_U236 & new_P1_R1171_U168;
  assign new_P1_R1171_U128 = new_P1_R1171_U245 & new_P1_R1171_U169;
  assign new_P1_R1171_U129 = new_P1_R1171_U265 & new_P1_R1171_U264;
  assign new_P1_R1171_U130 = new_P1_R1171_U10 & new_P1_R1171_U279;
  assign new_P1_R1171_U131 = new_P1_R1171_U282 & new_P1_R1171_U277;
  assign new_P1_R1171_U132 = new_P1_R1171_U298 & new_P1_R1171_U295;
  assign new_P1_R1171_U133 = new_P1_R1171_U365 & new_P1_R1171_U299;
  assign new_P1_R1171_U134 = new_P1_R1171_U156 & new_P1_R1171_U275;
  assign new_P1_R1171_U135 = new_P1_R1171_U60 & new_P1_R1171_U466 & new_P1_R1171_U465;
  assign new_P1_R1171_U136 = new_P1_R1171_U169 & new_P1_R1171_U487 & new_P1_R1171_U486;
  assign new_P1_R1171_U137 = new_P1_R1171_U340 & new_P1_R1171_U8;
  assign new_P1_R1171_U138 = new_P1_R1171_U168 & new_P1_R1171_U499 & new_P1_R1171_U498;
  assign new_P1_R1171_U139 = new_P1_R1171_U347 & new_P1_R1171_U7;
  assign new_P1_R1171_U140 = ~new_P1_R1171_U119 | ~new_P1_R1171_U199;
  assign new_P1_R1171_U141 = ~new_P1_R1171_U214 | ~new_P1_R1171_U226;
  assign new_P1_R1171_U142 = ~new_P1_U3055;
  assign new_P1_R1171_U143 = ~new_P1_U4028;
  assign new_P1_R1171_U144 = new_P1_R1171_U400 & new_P1_R1171_U399;
  assign new_P1_R1171_U145 = ~new_P1_R1171_U361 | ~new_P1_R1171_U301 | ~new_P1_R1171_U166;
  assign new_P1_R1171_U146 = new_P1_R1171_U407 & new_P1_R1171_U406;
  assign new_P1_R1171_U147 = ~new_P1_R1171_U133 | ~new_P1_R1171_U367 | ~new_P1_R1171_U366;
  assign new_P1_R1171_U148 = new_P1_R1171_U414 & new_P1_R1171_U413;
  assign new_P1_R1171_U149 = ~new_P1_R1171_U87 | ~new_P1_R1171_U362 | ~new_P1_R1171_U296;
  assign new_P1_R1171_U150 = new_P1_R1171_U421 & new_P1_R1171_U420;
  assign new_P1_R1171_U151 = ~new_P1_R1171_U290 | ~new_P1_R1171_U289;
  assign new_P1_R1171_U152 = new_P1_R1171_U433 & new_P1_R1171_U432;
  assign new_P1_R1171_U153 = ~new_P1_R1171_U286 | ~new_P1_R1171_U285;
  assign new_P1_R1171_U154 = new_P1_R1171_U440 & new_P1_R1171_U439;
  assign new_P1_R1171_U155 = ~new_P1_R1171_U131 | ~new_P1_R1171_U281;
  assign new_P1_R1171_U156 = new_P1_R1171_U447 & new_P1_R1171_U446;
  assign new_P1_R1171_U157 = new_P1_R1171_U452 & new_P1_R1171_U451;
  assign new_P1_R1171_U158 = ~new_P1_R1171_U44 | ~new_P1_R1171_U324;
  assign new_P1_R1171_U159 = ~new_P1_R1171_U129 | ~new_P1_R1171_U266;
  assign new_P1_R1171_U160 = new_P1_R1171_U473 & new_P1_R1171_U472;
  assign new_P1_R1171_U161 = ~new_P1_R1171_U254 | ~new_P1_R1171_U253;
  assign new_P1_R1171_U162 = new_P1_R1171_U480 & new_P1_R1171_U479;
  assign new_P1_R1171_U163 = ~new_P1_R1171_U250 | ~new_P1_R1171_U249;
  assign new_P1_R1171_U164 = ~new_P1_R1171_U240 | ~new_P1_R1171_U239;
  assign new_P1_R1171_U165 = ~new_P1_R1171_U364 | ~new_P1_R1171_U363;
  assign new_P1_R1171_U166 = ~new_P1_U3054 | ~new_P1_R1171_U147;
  assign new_P1_R1171_U167 = ~new_P1_R1171_U35;
  assign new_P1_R1171_U168 = ~new_P1_U3485 | ~new_P1_U3083;
  assign new_P1_R1171_U169 = ~new_P1_U3072 | ~new_P1_U3494;
  assign new_P1_R1171_U170 = ~new_P1_U3058 | ~new_P1_U4020;
  assign new_P1_R1171_U171 = ~new_P1_R1171_U69;
  assign new_P1_R1171_U172 = ~new_P1_R1171_U78;
  assign new_P1_R1171_U173 = ~new_P1_U3065 | ~new_P1_U4021;
  assign new_P1_R1171_U174 = ~new_P1_R1171_U62;
  assign new_P1_R1171_U175 = new_P1_U3067 | new_P1_U3473;
  assign new_P1_R1171_U176 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1171_U177 = new_P1_U3467 | new_P1_U3064;
  assign new_P1_R1171_U178 = new_P1_U3464 | new_P1_U3068;
  assign new_P1_R1171_U179 = ~new_P1_R1171_U32;
  assign new_P1_R1171_U180 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1171_U181 = ~new_P1_R1171_U43;
  assign new_P1_R1171_U182 = ~new_P1_R1171_U44;
  assign new_P1_R1171_U183 = ~new_P1_R1171_U43 | ~new_P1_R1171_U44;
  assign new_P1_R1171_U184 = ~new_P1_R1171_U116 | ~new_P1_R1171_U177;
  assign new_P1_R1171_U185 = ~new_P1_R1171_U5 | ~new_P1_R1171_U183;
  assign new_P1_R1171_U186 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1171_U187 = ~new_P1_R1171_U117 | ~new_P1_R1171_U185;
  assign new_P1_R1171_U188 = ~new_P1_R1171_U36 | ~new_P1_R1171_U35;
  assign new_P1_R1171_U189 = ~new_P1_U3067 | ~new_P1_R1171_U188;
  assign new_P1_R1171_U190 = ~new_P1_R1171_U4 | ~new_P1_R1171_U187;
  assign new_P1_R1171_U191 = ~new_P1_U3473 | ~new_P1_R1171_U167;
  assign new_P1_R1171_U192 = ~new_P1_R1171_U42;
  assign new_P1_R1171_U193 = new_P1_U3070 | new_P1_U3479;
  assign new_P1_R1171_U194 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1171_U195 = ~new_P1_R1171_U23;
  assign new_P1_R1171_U196 = ~new_P1_R1171_U24 | ~new_P1_R1171_U23;
  assign new_P1_R1171_U197 = ~new_P1_U3070 | ~new_P1_R1171_U196;
  assign new_P1_R1171_U198 = ~new_P1_U3479 | ~new_P1_R1171_U195;
  assign new_P1_R1171_U199 = ~new_P1_R1171_U6 | ~new_P1_R1171_U42;
  assign new_P1_R1171_U200 = ~new_P1_R1171_U140;
  assign new_P1_R1171_U201 = new_P1_U3482 | new_P1_U3084;
  assign new_P1_R1171_U202 = ~new_P1_R1171_U201 | ~new_P1_R1171_U140;
  assign new_P1_R1171_U203 = ~new_P1_R1171_U41;
  assign new_P1_R1171_U204 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1171_U205 = new_P1_U3476 | new_P1_U3071;
  assign new_P1_R1171_U206 = ~new_P1_R1171_U205 | ~new_P1_R1171_U42;
  assign new_P1_R1171_U207 = ~new_P1_R1171_U120 | ~new_P1_R1171_U206;
  assign new_P1_R1171_U208 = ~new_P1_R1171_U192 | ~new_P1_R1171_U23;
  assign new_P1_R1171_U209 = ~new_P1_U3479 | ~new_P1_U3070;
  assign new_P1_R1171_U210 = ~new_P1_R1171_U121 | ~new_P1_R1171_U208;
  assign new_P1_R1171_U211 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1171_U212 = ~new_P1_R1171_U182 | ~new_P1_R1171_U178;
  assign new_P1_R1171_U213 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1171_U214 = ~new_P1_R1171_U46;
  assign new_P1_R1171_U215 = ~new_P1_R1171_U181 | ~new_P1_R1171_U5;
  assign new_P1_R1171_U216 = ~new_P1_R1171_U46 | ~new_P1_R1171_U177;
  assign new_P1_R1171_U217 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1171_U218 = ~new_P1_R1171_U45;
  assign new_P1_R1171_U219 = new_P1_U3470 | new_P1_U3060;
  assign new_P1_R1171_U220 = ~new_P1_R1171_U219 | ~new_P1_R1171_U45;
  assign new_P1_R1171_U221 = ~new_P1_R1171_U123 | ~new_P1_R1171_U220;
  assign new_P1_R1171_U222 = ~new_P1_R1171_U218 | ~new_P1_R1171_U35;
  assign new_P1_R1171_U223 = ~new_P1_U3473 | ~new_P1_U3067;
  assign new_P1_R1171_U224 = ~new_P1_R1171_U124 | ~new_P1_R1171_U222;
  assign new_P1_R1171_U225 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1171_U226 = ~new_P1_R1171_U181 | ~new_P1_R1171_U178;
  assign new_P1_R1171_U227 = ~new_P1_R1171_U141;
  assign new_P1_R1171_U228 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1171_U229 = ~new_P1_R1171_U43 | ~new_P1_R1171_U44 | ~new_P1_R1171_U398 | ~new_P1_R1171_U397;
  assign new_P1_R1171_U230 = ~new_P1_R1171_U44 | ~new_P1_R1171_U43;
  assign new_P1_R1171_U231 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1171_U232 = ~new_P1_R1171_U125 | ~new_P1_R1171_U230;
  assign new_P1_R1171_U233 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1171_U234 = new_P1_U3062 | new_P1_U3488;
  assign new_P1_R1171_U235 = ~new_P1_R1171_U174 | ~new_P1_R1171_U7;
  assign new_P1_R1171_U236 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1171_U237 = ~new_P1_R1171_U127 | ~new_P1_R1171_U235;
  assign new_P1_R1171_U238 = new_P1_U3488 | new_P1_U3062;
  assign new_P1_R1171_U239 = ~new_P1_R1171_U126 | ~new_P1_R1171_U140;
  assign new_P1_R1171_U240 = ~new_P1_R1171_U238 | ~new_P1_R1171_U237;
  assign new_P1_R1171_U241 = ~new_P1_R1171_U164;
  assign new_P1_R1171_U242 = new_P1_U3080 | new_P1_U3497;
  assign new_P1_R1171_U243 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1171_U244 = ~new_P1_R1171_U171 | ~new_P1_R1171_U8;
  assign new_P1_R1171_U245 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1171_U246 = ~new_P1_R1171_U128 | ~new_P1_R1171_U244;
  assign new_P1_R1171_U247 = new_P1_U3491 | new_P1_U3063;
  assign new_P1_R1171_U248 = new_P1_U3497 | new_P1_U3080;
  assign new_P1_R1171_U249 = ~new_P1_R1171_U8 | ~new_P1_R1171_U247 | ~new_P1_R1171_U164;
  assign new_P1_R1171_U250 = ~new_P1_R1171_U248 | ~new_P1_R1171_U246;
  assign new_P1_R1171_U251 = ~new_P1_R1171_U163;
  assign new_P1_R1171_U252 = new_P1_U3500 | new_P1_U3079;
  assign new_P1_R1171_U253 = ~new_P1_R1171_U252 | ~new_P1_R1171_U163;
  assign new_P1_R1171_U254 = ~new_P1_U3079 | ~new_P1_U3500;
  assign new_P1_R1171_U255 = ~new_P1_R1171_U161;
  assign new_P1_R1171_U256 = new_P1_U3503 | new_P1_U3074;
  assign new_P1_R1171_U257 = ~new_P1_R1171_U256 | ~new_P1_R1171_U161;
  assign new_P1_R1171_U258 = ~new_P1_U3074 | ~new_P1_U3503;
  assign new_P1_R1171_U259 = ~new_P1_R1171_U93;
  assign new_P1_R1171_U260 = new_P1_U3069 | new_P1_U3509;
  assign new_P1_R1171_U261 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1171_U262 = ~new_P1_R1171_U60;
  assign new_P1_R1171_U263 = ~new_P1_R1171_U61 | ~new_P1_R1171_U60;
  assign new_P1_R1171_U264 = ~new_P1_U3069 | ~new_P1_R1171_U263;
  assign new_P1_R1171_U265 = ~new_P1_U3509 | ~new_P1_R1171_U262;
  assign new_P1_R1171_U266 = ~new_P1_R1171_U9 | ~new_P1_R1171_U93;
  assign new_P1_R1171_U267 = ~new_P1_R1171_U159;
  assign new_P1_R1171_U268 = new_P1_U3076 | new_P1_U4025;
  assign new_P1_R1171_U269 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1171_U270 = new_P1_U3075 | new_P1_U4024;
  assign new_P1_R1171_U271 = ~new_P1_R1171_U81;
  assign new_P1_R1171_U272 = ~new_P1_U4025 | ~new_P1_R1171_U271;
  assign new_P1_R1171_U273 = ~new_P1_R1171_U272 | ~new_P1_R1171_U91;
  assign new_P1_R1171_U274 = ~new_P1_R1171_U81 | ~new_P1_R1171_U82;
  assign new_P1_R1171_U275 = ~new_P1_R1171_U274 | ~new_P1_R1171_U273;
  assign new_P1_R1171_U276 = ~new_P1_R1171_U172 | ~new_P1_R1171_U10;
  assign new_P1_R1171_U277 = ~new_P1_U3075 | ~new_P1_U4024;
  assign new_P1_R1171_U278 = ~new_P1_R1171_U275 | ~new_P1_R1171_U276;
  assign new_P1_R1171_U279 = new_P1_U3512 | new_P1_U3082;
  assign new_P1_R1171_U280 = new_P1_U4024 | new_P1_U3075;
  assign new_P1_R1171_U281 = ~new_P1_R1171_U130 | ~new_P1_R1171_U270 | ~new_P1_R1171_U159;
  assign new_P1_R1171_U282 = ~new_P1_R1171_U280 | ~new_P1_R1171_U278;
  assign new_P1_R1171_U283 = ~new_P1_R1171_U155;
  assign new_P1_R1171_U284 = new_P1_U4023 | new_P1_U3061;
  assign new_P1_R1171_U285 = ~new_P1_R1171_U284 | ~new_P1_R1171_U155;
  assign new_P1_R1171_U286 = ~new_P1_U3061 | ~new_P1_U4023;
  assign new_P1_R1171_U287 = ~new_P1_R1171_U153;
  assign new_P1_R1171_U288 = new_P1_U4022 | new_P1_U3066;
  assign new_P1_R1171_U289 = ~new_P1_R1171_U288 | ~new_P1_R1171_U153;
  assign new_P1_R1171_U290 = ~new_P1_U3066 | ~new_P1_U4022;
  assign new_P1_R1171_U291 = ~new_P1_R1171_U151;
  assign new_P1_R1171_U292 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1171_U293 = ~new_P1_R1171_U173 | ~new_P1_R1171_U170;
  assign new_P1_R1171_U294 = ~new_P1_R1171_U87;
  assign new_P1_R1171_U295 = new_P1_U4021 | new_P1_U3065;
  assign new_P1_R1171_U296 = ~new_P1_R1171_U165 | ~new_P1_R1171_U151 | ~new_P1_R1171_U295;
  assign new_P1_R1171_U297 = ~new_P1_R1171_U149;
  assign new_P1_R1171_U298 = new_P1_U4018 | new_P1_U3053;
  assign new_P1_R1171_U299 = ~new_P1_U3053 | ~new_P1_U4018;
  assign new_P1_R1171_U300 = ~new_P1_R1171_U147;
  assign new_P1_R1171_U301 = ~new_P1_U4017 | ~new_P1_R1171_U147;
  assign new_P1_R1171_U302 = ~new_P1_R1171_U145;
  assign new_P1_R1171_U303 = ~new_P1_R1171_U295 | ~new_P1_R1171_U151;
  assign new_P1_R1171_U304 = ~new_P1_R1171_U90;
  assign new_P1_R1171_U305 = new_P1_U4020 | new_P1_U3058;
  assign new_P1_R1171_U306 = ~new_P1_R1171_U305 | ~new_P1_R1171_U90;
  assign new_P1_R1171_U307 = ~new_P1_R1171_U150 | ~new_P1_R1171_U306 | ~new_P1_R1171_U170;
  assign new_P1_R1171_U308 = ~new_P1_R1171_U304 | ~new_P1_R1171_U170;
  assign new_P1_R1171_U309 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1171_U310 = ~new_P1_R1171_U165 | ~new_P1_R1171_U308 | ~new_P1_R1171_U309;
  assign new_P1_R1171_U311 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1171_U312 = ~new_P1_R1171_U279 | ~new_P1_R1171_U159;
  assign new_P1_R1171_U313 = ~new_P1_R1171_U92;
  assign new_P1_R1171_U314 = ~new_P1_R1171_U10 | ~new_P1_R1171_U92;
  assign new_P1_R1171_U315 = ~new_P1_R1171_U134 | ~new_P1_R1171_U314;
  assign new_P1_R1171_U316 = ~new_P1_R1171_U314 | ~new_P1_R1171_U275;
  assign new_P1_R1171_U317 = ~new_P1_R1171_U450 | ~new_P1_R1171_U316;
  assign new_P1_R1171_U318 = new_P1_U3514 | new_P1_U3081;
  assign new_P1_R1171_U319 = ~new_P1_R1171_U318 | ~new_P1_R1171_U92;
  assign new_P1_R1171_U320 = ~new_P1_R1171_U157 | ~new_P1_R1171_U319 | ~new_P1_R1171_U81;
  assign new_P1_R1171_U321 = ~new_P1_R1171_U313 | ~new_P1_R1171_U81;
  assign new_P1_R1171_U322 = ~new_P1_U3076 | ~new_P1_U4025;
  assign new_P1_R1171_U323 = ~new_P1_R1171_U10 | ~new_P1_R1171_U322 | ~new_P1_R1171_U321;
  assign new_P1_R1171_U324 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1171_U325 = ~new_P1_R1171_U158;
  assign new_P1_R1171_U326 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1171_U327 = new_P1_U3506 | new_P1_U3073;
  assign new_P1_R1171_U328 = ~new_P1_R1171_U327 | ~new_P1_R1171_U93;
  assign new_P1_R1171_U329 = ~new_P1_R1171_U135 | ~new_P1_R1171_U328;
  assign new_P1_R1171_U330 = ~new_P1_R1171_U259 | ~new_P1_R1171_U60;
  assign new_P1_R1171_U331 = ~new_P1_U3509 | ~new_P1_U3069;
  assign new_P1_R1171_U332 = ~new_P1_R1171_U9 | ~new_P1_R1171_U331 | ~new_P1_R1171_U330;
  assign new_P1_R1171_U333 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1171_U334 = ~new_P1_R1171_U247 | ~new_P1_R1171_U164;
  assign new_P1_R1171_U335 = ~new_P1_R1171_U94;
  assign new_P1_R1171_U336 = new_P1_U3494 | new_P1_U3072;
  assign new_P1_R1171_U337 = ~new_P1_R1171_U336 | ~new_P1_R1171_U94;
  assign new_P1_R1171_U338 = ~new_P1_R1171_U136 | ~new_P1_R1171_U337;
  assign new_P1_R1171_U339 = ~new_P1_R1171_U335 | ~new_P1_R1171_U169;
  assign new_P1_R1171_U340 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1171_U341 = ~new_P1_R1171_U137 | ~new_P1_R1171_U339;
  assign new_P1_R1171_U342 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1171_U343 = new_P1_U3485 | new_P1_U3083;
  assign new_P1_R1171_U344 = ~new_P1_R1171_U343 | ~new_P1_R1171_U41;
  assign new_P1_R1171_U345 = ~new_P1_R1171_U138 | ~new_P1_R1171_U344;
  assign new_P1_R1171_U346 = ~new_P1_R1171_U203 | ~new_P1_R1171_U168;
  assign new_P1_R1171_U347 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1171_U348 = ~new_P1_R1171_U139 | ~new_P1_R1171_U346;
  assign new_P1_R1171_U349 = ~new_P1_R1171_U204 | ~new_P1_R1171_U168;
  assign new_P1_R1171_U350 = ~new_P1_R1171_U201 | ~new_P1_R1171_U62;
  assign new_P1_R1171_U351 = ~new_P1_R1171_U211 | ~new_P1_R1171_U23;
  assign new_P1_R1171_U352 = ~new_P1_R1171_U225 | ~new_P1_R1171_U35;
  assign new_P1_R1171_U353 = ~new_P1_R1171_U228 | ~new_P1_R1171_U177;
  assign new_P1_R1171_U354 = ~new_P1_R1171_U311 | ~new_P1_R1171_U170;
  assign new_P1_R1171_U355 = ~new_P1_R1171_U295 | ~new_P1_R1171_U173;
  assign new_P1_R1171_U356 = ~new_P1_R1171_U326 | ~new_P1_R1171_U81;
  assign new_P1_R1171_U357 = ~new_P1_R1171_U279 | ~new_P1_R1171_U78;
  assign new_P1_R1171_U358 = ~new_P1_R1171_U333 | ~new_P1_R1171_U60;
  assign new_P1_R1171_U359 = ~new_P1_R1171_U342 | ~new_P1_R1171_U169;
  assign new_P1_R1171_U360 = ~new_P1_R1171_U247 | ~new_P1_R1171_U69;
  assign new_P1_R1171_U361 = ~new_P1_U4017 | ~new_P1_U3054;
  assign new_P1_R1171_U362 = ~new_P1_R1171_U293 | ~new_P1_R1171_U165;
  assign new_P1_R1171_U363 = ~new_P1_U3057 | ~new_P1_R1171_U292;
  assign new_P1_R1171_U364 = ~new_P1_U4019 | ~new_P1_R1171_U292;
  assign new_P1_R1171_U365 = ~new_P1_R1171_U298 | ~new_P1_R1171_U293 | ~new_P1_R1171_U165;
  assign new_P1_R1171_U366 = ~new_P1_R1171_U132 | ~new_P1_R1171_U151 | ~new_P1_R1171_U165;
  assign new_P1_R1171_U367 = ~new_P1_R1171_U294 | ~new_P1_R1171_U298;
  assign new_P1_R1171_U368 = ~new_P1_U3083 | ~new_P1_R1171_U40;
  assign new_P1_R1171_U369 = ~new_P1_U3485 | ~new_P1_R1171_U39;
  assign new_P1_R1171_U370 = ~new_P1_R1171_U369 | ~new_P1_R1171_U368;
  assign new_P1_R1171_U371 = ~new_P1_R1171_U349 | ~new_P1_R1171_U41;
  assign new_P1_R1171_U372 = ~new_P1_R1171_U370 | ~new_P1_R1171_U203;
  assign new_P1_R1171_U373 = ~new_P1_U3084 | ~new_P1_R1171_U37;
  assign new_P1_R1171_U374 = ~new_P1_U3482 | ~new_P1_R1171_U38;
  assign new_P1_R1171_U375 = ~new_P1_R1171_U374 | ~new_P1_R1171_U373;
  assign new_P1_R1171_U376 = ~new_P1_R1171_U350 | ~new_P1_R1171_U140;
  assign new_P1_R1171_U377 = ~new_P1_R1171_U200 | ~new_P1_R1171_U375;
  assign new_P1_R1171_U378 = ~new_P1_U3070 | ~new_P1_R1171_U24;
  assign new_P1_R1171_U379 = ~new_P1_U3479 | ~new_P1_R1171_U22;
  assign new_P1_R1171_U380 = ~new_P1_U3071 | ~new_P1_R1171_U20;
  assign new_P1_R1171_U381 = ~new_P1_U3476 | ~new_P1_R1171_U21;
  assign new_P1_R1171_U382 = ~new_P1_R1171_U381 | ~new_P1_R1171_U380;
  assign new_P1_R1171_U383 = ~new_P1_R1171_U351 | ~new_P1_R1171_U42;
  assign new_P1_R1171_U384 = ~new_P1_R1171_U382 | ~new_P1_R1171_U192;
  assign new_P1_R1171_U385 = ~new_P1_U3067 | ~new_P1_R1171_U36;
  assign new_P1_R1171_U386 = ~new_P1_U3473 | ~new_P1_R1171_U27;
  assign new_P1_R1171_U387 = ~new_P1_U3060 | ~new_P1_R1171_U25;
  assign new_P1_R1171_U388 = ~new_P1_U3470 | ~new_P1_R1171_U26;
  assign new_P1_R1171_U389 = ~new_P1_R1171_U388 | ~new_P1_R1171_U387;
  assign new_P1_R1171_U390 = ~new_P1_R1171_U352 | ~new_P1_R1171_U45;
  assign new_P1_R1171_U391 = ~new_P1_R1171_U389 | ~new_P1_R1171_U218;
  assign new_P1_R1171_U392 = ~new_P1_U3064 | ~new_P1_R1171_U33;
  assign new_P1_R1171_U393 = ~new_P1_U3467 | ~new_P1_R1171_U34;
  assign new_P1_R1171_U394 = ~new_P1_R1171_U393 | ~new_P1_R1171_U392;
  assign new_P1_R1171_U395 = ~new_P1_R1171_U353 | ~new_P1_R1171_U141;
  assign new_P1_R1171_U396 = ~new_P1_R1171_U227 | ~new_P1_R1171_U394;
  assign new_P1_R1171_U397 = ~new_P1_U3068 | ~new_P1_R1171_U28;
  assign new_P1_R1171_U398 = ~new_P1_U3464 | ~new_P1_R1171_U29;
  assign new_P1_R1171_U399 = ~new_P1_U3055 | ~new_P1_R1171_U143;
  assign new_P1_R1171_U400 = ~new_P1_U4028 | ~new_P1_R1171_U142;
  assign new_P1_R1171_U401 = ~new_P1_U3055 | ~new_P1_R1171_U143;
  assign new_P1_R1171_U402 = ~new_P1_U4028 | ~new_P1_R1171_U142;
  assign new_P1_R1171_U403 = ~new_P1_R1171_U402 | ~new_P1_R1171_U401;
  assign new_P1_R1171_U404 = ~new_P1_R1171_U144 | ~new_P1_R1171_U145;
  assign new_P1_R1171_U405 = ~new_P1_R1171_U302 | ~new_P1_R1171_U403;
  assign new_P1_R1171_U406 = ~new_P1_U3054 | ~new_P1_R1171_U89;
  assign new_P1_R1171_U407 = ~new_P1_U4017 | ~new_P1_R1171_U88;
  assign new_P1_R1171_U408 = ~new_P1_U3054 | ~new_P1_R1171_U89;
  assign new_P1_R1171_U409 = ~new_P1_U4017 | ~new_P1_R1171_U88;
  assign new_P1_R1171_U410 = ~new_P1_R1171_U409 | ~new_P1_R1171_U408;
  assign new_P1_R1171_U411 = ~new_P1_R1171_U146 | ~new_P1_R1171_U147;
  assign new_P1_R1171_U412 = ~new_P1_R1171_U300 | ~new_P1_R1171_U410;
  assign new_P1_R1171_U413 = ~new_P1_U3053 | ~new_P1_R1171_U47;
  assign new_P1_R1171_U414 = ~new_P1_U4018 | ~new_P1_R1171_U48;
  assign new_P1_R1171_U415 = ~new_P1_U3053 | ~new_P1_R1171_U47;
  assign new_P1_R1171_U416 = ~new_P1_U4018 | ~new_P1_R1171_U48;
  assign new_P1_R1171_U417 = ~new_P1_R1171_U416 | ~new_P1_R1171_U415;
  assign new_P1_R1171_U418 = ~new_P1_R1171_U148 | ~new_P1_R1171_U149;
  assign new_P1_R1171_U419 = ~new_P1_R1171_U297 | ~new_P1_R1171_U417;
  assign new_P1_R1171_U420 = ~new_P1_U3057 | ~new_P1_R1171_U50;
  assign new_P1_R1171_U421 = ~new_P1_U4019 | ~new_P1_R1171_U49;
  assign new_P1_R1171_U422 = ~new_P1_U3058 | ~new_P1_R1171_U51;
  assign new_P1_R1171_U423 = ~new_P1_U4020 | ~new_P1_R1171_U52;
  assign new_P1_R1171_U424 = ~new_P1_R1171_U423 | ~new_P1_R1171_U422;
  assign new_P1_R1171_U425 = ~new_P1_R1171_U354 | ~new_P1_R1171_U90;
  assign new_P1_R1171_U426 = ~new_P1_R1171_U424 | ~new_P1_R1171_U304;
  assign new_P1_R1171_U427 = ~new_P1_U3065 | ~new_P1_R1171_U53;
  assign new_P1_R1171_U428 = ~new_P1_U4021 | ~new_P1_R1171_U54;
  assign new_P1_R1171_U429 = ~new_P1_R1171_U428 | ~new_P1_R1171_U427;
  assign new_P1_R1171_U430 = ~new_P1_R1171_U355 | ~new_P1_R1171_U151;
  assign new_P1_R1171_U431 = ~new_P1_R1171_U291 | ~new_P1_R1171_U429;
  assign new_P1_R1171_U432 = ~new_P1_U3066 | ~new_P1_R1171_U85;
  assign new_P1_R1171_U433 = ~new_P1_U4022 | ~new_P1_R1171_U86;
  assign new_P1_R1171_U434 = ~new_P1_U3066 | ~new_P1_R1171_U85;
  assign new_P1_R1171_U435 = ~new_P1_U4022 | ~new_P1_R1171_U86;
  assign new_P1_R1171_U436 = ~new_P1_R1171_U435 | ~new_P1_R1171_U434;
  assign new_P1_R1171_U437 = ~new_P1_R1171_U152 | ~new_P1_R1171_U153;
  assign new_P1_R1171_U438 = ~new_P1_R1171_U287 | ~new_P1_R1171_U436;
  assign new_P1_R1171_U439 = ~new_P1_U3061 | ~new_P1_R1171_U83;
  assign new_P1_R1171_U440 = ~new_P1_U4023 | ~new_P1_R1171_U84;
  assign new_P1_R1171_U441 = ~new_P1_U3061 | ~new_P1_R1171_U83;
  assign new_P1_R1171_U442 = ~new_P1_U4023 | ~new_P1_R1171_U84;
  assign new_P1_R1171_U443 = ~new_P1_R1171_U442 | ~new_P1_R1171_U441;
  assign new_P1_R1171_U444 = ~new_P1_R1171_U154 | ~new_P1_R1171_U155;
  assign new_P1_R1171_U445 = ~new_P1_R1171_U283 | ~new_P1_R1171_U443;
  assign new_P1_R1171_U446 = ~new_P1_U3075 | ~new_P1_R1171_U55;
  assign new_P1_R1171_U447 = ~new_P1_U4024 | ~new_P1_R1171_U56;
  assign new_P1_R1171_U448 = ~new_P1_U3075 | ~new_P1_R1171_U55;
  assign new_P1_R1171_U449 = ~new_P1_U4024 | ~new_P1_R1171_U56;
  assign new_P1_R1171_U450 = ~new_P1_R1171_U449 | ~new_P1_R1171_U448;
  assign new_P1_R1171_U451 = ~new_P1_U3076 | ~new_P1_R1171_U82;
  assign new_P1_R1171_U452 = ~new_P1_U4025 | ~new_P1_R1171_U91;
  assign new_P1_R1171_U453 = ~new_P1_R1171_U179 | ~new_P1_R1171_U158;
  assign new_P1_R1171_U454 = ~new_P1_R1171_U325 | ~new_P1_R1171_U32;
  assign new_P1_R1171_U455 = ~new_P1_U3081 | ~new_P1_R1171_U79;
  assign new_P1_R1171_U456 = ~new_P1_U3514 | ~new_P1_R1171_U80;
  assign new_P1_R1171_U457 = ~new_P1_R1171_U456 | ~new_P1_R1171_U455;
  assign new_P1_R1171_U458 = ~new_P1_R1171_U356 | ~new_P1_R1171_U92;
  assign new_P1_R1171_U459 = ~new_P1_R1171_U457 | ~new_P1_R1171_U313;
  assign new_P1_R1171_U460 = ~new_P1_U3082 | ~new_P1_R1171_U76;
  assign new_P1_R1171_U461 = ~new_P1_U3512 | ~new_P1_R1171_U77;
  assign new_P1_R1171_U462 = ~new_P1_R1171_U461 | ~new_P1_R1171_U460;
  assign new_P1_R1171_U463 = ~new_P1_R1171_U357 | ~new_P1_R1171_U159;
  assign new_P1_R1171_U464 = ~new_P1_R1171_U267 | ~new_P1_R1171_U462;
  assign new_P1_R1171_U465 = ~new_P1_U3069 | ~new_P1_R1171_U61;
  assign new_P1_R1171_U466 = ~new_P1_U3509 | ~new_P1_R1171_U59;
  assign new_P1_R1171_U467 = ~new_P1_U3073 | ~new_P1_R1171_U57;
  assign new_P1_R1171_U468 = ~new_P1_U3506 | ~new_P1_R1171_U58;
  assign new_P1_R1171_U469 = ~new_P1_R1171_U468 | ~new_P1_R1171_U467;
  assign new_P1_R1171_U470 = ~new_P1_R1171_U358 | ~new_P1_R1171_U93;
  assign new_P1_R1171_U471 = ~new_P1_R1171_U469 | ~new_P1_R1171_U259;
  assign new_P1_R1171_U472 = ~new_P1_U3074 | ~new_P1_R1171_U74;
  assign new_P1_R1171_U473 = ~new_P1_U3503 | ~new_P1_R1171_U75;
  assign new_P1_R1171_U474 = ~new_P1_U3074 | ~new_P1_R1171_U74;
  assign new_P1_R1171_U475 = ~new_P1_U3503 | ~new_P1_R1171_U75;
  assign new_P1_R1171_U476 = ~new_P1_R1171_U475 | ~new_P1_R1171_U474;
  assign new_P1_R1171_U477 = ~new_P1_R1171_U160 | ~new_P1_R1171_U161;
  assign new_P1_R1171_U478 = ~new_P1_R1171_U255 | ~new_P1_R1171_U476;
  assign new_P1_R1171_U479 = ~new_P1_U3079 | ~new_P1_R1171_U72;
  assign new_P1_R1171_U480 = ~new_P1_U3500 | ~new_P1_R1171_U73;
  assign new_P1_R1171_U481 = ~new_P1_U3079 | ~new_P1_R1171_U72;
  assign new_P1_R1171_U482 = ~new_P1_U3500 | ~new_P1_R1171_U73;
  assign new_P1_R1171_U483 = ~new_P1_R1171_U482 | ~new_P1_R1171_U481;
  assign new_P1_R1171_U484 = ~new_P1_R1171_U162 | ~new_P1_R1171_U163;
  assign new_P1_R1171_U485 = ~new_P1_R1171_U251 | ~new_P1_R1171_U483;
  assign new_P1_R1171_U486 = ~new_P1_U3080 | ~new_P1_R1171_U70;
  assign new_P1_R1171_U487 = ~new_P1_U3497 | ~new_P1_R1171_U71;
  assign new_P1_R1171_U488 = ~new_P1_U3072 | ~new_P1_R1171_U65;
  assign new_P1_R1171_U489 = ~new_P1_U3494 | ~new_P1_R1171_U66;
  assign new_P1_R1171_U490 = ~new_P1_R1171_U489 | ~new_P1_R1171_U488;
  assign new_P1_R1171_U491 = ~new_P1_R1171_U359 | ~new_P1_R1171_U94;
  assign new_P1_R1171_U492 = ~new_P1_R1171_U490 | ~new_P1_R1171_U335;
  assign new_P1_R1171_U493 = ~new_P1_U3063 | ~new_P1_R1171_U67;
  assign new_P1_R1171_U494 = ~new_P1_U3491 | ~new_P1_R1171_U68;
  assign new_P1_R1171_U495 = ~new_P1_R1171_U494 | ~new_P1_R1171_U493;
  assign new_P1_R1171_U496 = ~new_P1_R1171_U360 | ~new_P1_R1171_U164;
  assign new_P1_R1171_U497 = ~new_P1_R1171_U241 | ~new_P1_R1171_U495;
  assign new_P1_R1171_U498 = ~new_P1_U3062 | ~new_P1_R1171_U63;
  assign new_P1_R1171_U499 = ~new_P1_U3488 | ~new_P1_R1171_U64;
  assign new_P1_R1171_U500 = ~new_P1_U3077 | ~new_P1_R1171_U30;
  assign new_P1_R1171_U501 = ~new_P1_U3456 | ~new_P1_R1171_U31;
  assign new_P1_R1138_U4 = new_P1_R1138_U176 & new_P1_R1138_U175;
  assign new_P1_R1138_U5 = new_P1_R1138_U177 & new_P1_R1138_U178;
  assign new_P1_R1138_U6 = new_P1_R1138_U194 & new_P1_R1138_U193;
  assign new_P1_R1138_U7 = new_P1_R1138_U234 & new_P1_R1138_U233;
  assign new_P1_R1138_U8 = new_P1_R1138_U243 & new_P1_R1138_U242;
  assign new_P1_R1138_U9 = new_P1_R1138_U261 & new_P1_R1138_U260;
  assign new_P1_R1138_U10 = new_P1_R1138_U269 & new_P1_R1138_U268;
  assign new_P1_R1138_U11 = new_P1_R1138_U348 & new_P1_R1138_U345;
  assign new_P1_R1138_U12 = new_P1_R1138_U341 & new_P1_R1138_U338;
  assign new_P1_R1138_U13 = new_P1_R1138_U332 & new_P1_R1138_U329;
  assign new_P1_R1138_U14 = new_P1_R1138_U323 & new_P1_R1138_U320;
  assign new_P1_R1138_U15 = new_P1_R1138_U317 & new_P1_R1138_U315;
  assign new_P1_R1138_U16 = new_P1_R1138_U310 & new_P1_R1138_U307;
  assign new_P1_R1138_U17 = new_P1_R1138_U232 & new_P1_R1138_U229;
  assign new_P1_R1138_U18 = new_P1_R1138_U224 & new_P1_R1138_U221;
  assign new_P1_R1138_U19 = new_P1_R1138_U210 & new_P1_R1138_U207;
  assign new_P1_R1138_U20 = ~new_P1_U3476;
  assign new_P1_R1138_U21 = ~new_P1_U3071;
  assign new_P1_R1138_U22 = ~new_P1_U3070;
  assign new_P1_R1138_U23 = ~new_P1_U3071 | ~new_P1_U3476;
  assign new_P1_R1138_U24 = ~new_P1_U3479;
  assign new_P1_R1138_U25 = ~new_P1_U3470;
  assign new_P1_R1138_U26 = ~new_P1_U3060;
  assign new_P1_R1138_U27 = ~new_P1_U3067;
  assign new_P1_R1138_U28 = ~new_P1_U3464;
  assign new_P1_R1138_U29 = ~new_P1_U3068;
  assign new_P1_R1138_U30 = ~new_P1_U3456;
  assign new_P1_R1138_U31 = ~new_P1_U3077;
  assign new_P1_R1138_U32 = ~new_P1_U3077 | ~new_P1_U3456;
  assign new_P1_R1138_U33 = ~new_P1_U3467;
  assign new_P1_R1138_U34 = ~new_P1_U3064;
  assign new_P1_R1138_U35 = ~new_P1_U3060 | ~new_P1_U3470;
  assign new_P1_R1138_U36 = ~new_P1_U3473;
  assign new_P1_R1138_U37 = ~new_P1_U3482;
  assign new_P1_R1138_U38 = ~new_P1_U3084;
  assign new_P1_R1138_U39 = ~new_P1_U3083;
  assign new_P1_R1138_U40 = ~new_P1_U3485;
  assign new_P1_R1138_U41 = ~new_P1_R1138_U62 | ~new_P1_R1138_U202;
  assign new_P1_R1138_U42 = ~new_P1_R1138_U118 | ~new_P1_R1138_U190;
  assign new_P1_R1138_U43 = ~new_P1_R1138_U179 | ~new_P1_R1138_U180;
  assign new_P1_R1138_U44 = ~new_P1_U3461 | ~new_P1_U3078;
  assign new_P1_R1138_U45 = ~new_P1_R1138_U122 | ~new_P1_R1138_U216;
  assign new_P1_R1138_U46 = ~new_P1_R1138_U213 | ~new_P1_R1138_U212;
  assign new_P1_R1138_U47 = ~new_P1_U4018;
  assign new_P1_R1138_U48 = ~new_P1_U3053;
  assign new_P1_R1138_U49 = ~new_P1_U3057;
  assign new_P1_R1138_U50 = ~new_P1_U4019;
  assign new_P1_R1138_U51 = ~new_P1_U4020;
  assign new_P1_R1138_U52 = ~new_P1_U3058;
  assign new_P1_R1138_U53 = ~new_P1_U4021;
  assign new_P1_R1138_U54 = ~new_P1_U3065;
  assign new_P1_R1138_U55 = ~new_P1_U4024;
  assign new_P1_R1138_U56 = ~new_P1_U3075;
  assign new_P1_R1138_U57 = ~new_P1_U3506;
  assign new_P1_R1138_U58 = ~new_P1_U3073;
  assign new_P1_R1138_U59 = ~new_P1_U3069;
  assign new_P1_R1138_U60 = ~new_P1_U3073 | ~new_P1_U3506;
  assign new_P1_R1138_U61 = ~new_P1_U3509;
  assign new_P1_R1138_U62 = ~new_P1_U3084 | ~new_P1_U3482;
  assign new_P1_R1138_U63 = ~new_P1_U3488;
  assign new_P1_R1138_U64 = ~new_P1_U3062;
  assign new_P1_R1138_U65 = ~new_P1_U3494;
  assign new_P1_R1138_U66 = ~new_P1_U3072;
  assign new_P1_R1138_U67 = ~new_P1_U3491;
  assign new_P1_R1138_U68 = ~new_P1_U3063;
  assign new_P1_R1138_U69 = ~new_P1_U3063 | ~new_P1_U3491;
  assign new_P1_R1138_U70 = ~new_P1_U3497;
  assign new_P1_R1138_U71 = ~new_P1_U3080;
  assign new_P1_R1138_U72 = ~new_P1_U3500;
  assign new_P1_R1138_U73 = ~new_P1_U3079;
  assign new_P1_R1138_U74 = ~new_P1_U3503;
  assign new_P1_R1138_U75 = ~new_P1_U3074;
  assign new_P1_R1138_U76 = ~new_P1_U3512;
  assign new_P1_R1138_U77 = ~new_P1_U3082;
  assign new_P1_R1138_U78 = ~new_P1_U3082 | ~new_P1_U3512;
  assign new_P1_R1138_U79 = ~new_P1_U3514;
  assign new_P1_R1138_U80 = ~new_P1_U3081;
  assign new_P1_R1138_U81 = ~new_P1_U3081 | ~new_P1_U3514;
  assign new_P1_R1138_U82 = ~new_P1_U4025;
  assign new_P1_R1138_U83 = ~new_P1_U4023;
  assign new_P1_R1138_U84 = ~new_P1_U3061;
  assign new_P1_R1138_U85 = ~new_P1_U4022;
  assign new_P1_R1138_U86 = ~new_P1_U3066;
  assign new_P1_R1138_U87 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1138_U88 = ~new_P1_U3054;
  assign new_P1_R1138_U89 = ~new_P1_U4017;
  assign new_P1_R1138_U90 = ~new_P1_R1138_U303 | ~new_P1_R1138_U173;
  assign new_P1_R1138_U91 = ~new_P1_U3076;
  assign new_P1_R1138_U92 = ~new_P1_R1138_U78 | ~new_P1_R1138_U312;
  assign new_P1_R1138_U93 = ~new_P1_R1138_U258 | ~new_P1_R1138_U257;
  assign new_P1_R1138_U94 = ~new_P1_R1138_U69 | ~new_P1_R1138_U334;
  assign new_P1_R1138_U95 = ~new_P1_R1138_U454 | ~new_P1_R1138_U453;
  assign new_P1_R1138_U96 = ~new_P1_R1138_U501 | ~new_P1_R1138_U500;
  assign new_P1_R1138_U97 = ~new_P1_R1138_U372 | ~new_P1_R1138_U371;
  assign new_P1_R1138_U98 = ~new_P1_R1138_U377 | ~new_P1_R1138_U376;
  assign new_P1_R1138_U99 = ~new_P1_R1138_U384 | ~new_P1_R1138_U383;
  assign new_P1_R1138_U100 = ~new_P1_R1138_U391 | ~new_P1_R1138_U390;
  assign new_P1_R1138_U101 = ~new_P1_R1138_U396 | ~new_P1_R1138_U395;
  assign new_P1_R1138_U102 = ~new_P1_R1138_U405 | ~new_P1_R1138_U404;
  assign new_P1_R1138_U103 = ~new_P1_R1138_U412 | ~new_P1_R1138_U411;
  assign new_P1_R1138_U104 = ~new_P1_R1138_U419 | ~new_P1_R1138_U418;
  assign new_P1_R1138_U105 = ~new_P1_R1138_U426 | ~new_P1_R1138_U425;
  assign new_P1_R1138_U106 = ~new_P1_R1138_U431 | ~new_P1_R1138_U430;
  assign new_P1_R1138_U107 = ~new_P1_R1138_U438 | ~new_P1_R1138_U437;
  assign new_P1_R1138_U108 = ~new_P1_R1138_U445 | ~new_P1_R1138_U444;
  assign new_P1_R1138_U109 = ~new_P1_R1138_U459 | ~new_P1_R1138_U458;
  assign new_P1_R1138_U110 = ~new_P1_R1138_U464 | ~new_P1_R1138_U463;
  assign new_P1_R1138_U111 = ~new_P1_R1138_U471 | ~new_P1_R1138_U470;
  assign new_P1_R1138_U112 = ~new_P1_R1138_U478 | ~new_P1_R1138_U477;
  assign new_P1_R1138_U113 = ~new_P1_R1138_U485 | ~new_P1_R1138_U484;
  assign new_P1_R1138_U114 = ~new_P1_R1138_U492 | ~new_P1_R1138_U491;
  assign new_P1_R1138_U115 = ~new_P1_R1138_U497 | ~new_P1_R1138_U496;
  assign new_P1_R1138_U116 = new_P1_U3464 & new_P1_U3068;
  assign new_P1_R1138_U117 = new_P1_R1138_U186 & new_P1_R1138_U184;
  assign new_P1_R1138_U118 = new_P1_R1138_U191 & new_P1_R1138_U189;
  assign new_P1_R1138_U119 = new_P1_R1138_U198 & new_P1_R1138_U197;
  assign new_P1_R1138_U120 = new_P1_R1138_U23 & new_P1_R1138_U379 & new_P1_R1138_U378;
  assign new_P1_R1138_U121 = new_P1_R1138_U209 & new_P1_R1138_U6;
  assign new_P1_R1138_U122 = new_P1_R1138_U217 & new_P1_R1138_U215;
  assign new_P1_R1138_U123 = new_P1_R1138_U35 & new_P1_R1138_U386 & new_P1_R1138_U385;
  assign new_P1_R1138_U124 = new_P1_R1138_U223 & new_P1_R1138_U4;
  assign new_P1_R1138_U125 = new_P1_R1138_U231 & new_P1_R1138_U178;
  assign new_P1_R1138_U126 = new_P1_R1138_U201 & new_P1_R1138_U7;
  assign new_P1_R1138_U127 = new_P1_R1138_U236 & new_P1_R1138_U168;
  assign new_P1_R1138_U128 = new_P1_R1138_U245 & new_P1_R1138_U169;
  assign new_P1_R1138_U129 = new_P1_R1138_U265 & new_P1_R1138_U264;
  assign new_P1_R1138_U130 = new_P1_R1138_U10 & new_P1_R1138_U279;
  assign new_P1_R1138_U131 = new_P1_R1138_U282 & new_P1_R1138_U277;
  assign new_P1_R1138_U132 = new_P1_R1138_U298 & new_P1_R1138_U295;
  assign new_P1_R1138_U133 = new_P1_R1138_U365 & new_P1_R1138_U299;
  assign new_P1_R1138_U134 = new_P1_R1138_U156 & new_P1_R1138_U275;
  assign new_P1_R1138_U135 = new_P1_R1138_U60 & new_P1_R1138_U466 & new_P1_R1138_U465;
  assign new_P1_R1138_U136 = new_P1_R1138_U169 & new_P1_R1138_U487 & new_P1_R1138_U486;
  assign new_P1_R1138_U137 = new_P1_R1138_U340 & new_P1_R1138_U8;
  assign new_P1_R1138_U138 = new_P1_R1138_U168 & new_P1_R1138_U499 & new_P1_R1138_U498;
  assign new_P1_R1138_U139 = new_P1_R1138_U347 & new_P1_R1138_U7;
  assign new_P1_R1138_U140 = ~new_P1_R1138_U119 | ~new_P1_R1138_U199;
  assign new_P1_R1138_U141 = ~new_P1_R1138_U214 | ~new_P1_R1138_U226;
  assign new_P1_R1138_U142 = ~new_P1_U3055;
  assign new_P1_R1138_U143 = ~new_P1_U4028;
  assign new_P1_R1138_U144 = new_P1_R1138_U400 & new_P1_R1138_U399;
  assign new_P1_R1138_U145 = ~new_P1_R1138_U361 | ~new_P1_R1138_U301 | ~new_P1_R1138_U166;
  assign new_P1_R1138_U146 = new_P1_R1138_U407 & new_P1_R1138_U406;
  assign new_P1_R1138_U147 = ~new_P1_R1138_U133 | ~new_P1_R1138_U367 | ~new_P1_R1138_U366;
  assign new_P1_R1138_U148 = new_P1_R1138_U414 & new_P1_R1138_U413;
  assign new_P1_R1138_U149 = ~new_P1_R1138_U87 | ~new_P1_R1138_U362 | ~new_P1_R1138_U296;
  assign new_P1_R1138_U150 = new_P1_R1138_U421 & new_P1_R1138_U420;
  assign new_P1_R1138_U151 = ~new_P1_R1138_U290 | ~new_P1_R1138_U289;
  assign new_P1_R1138_U152 = new_P1_R1138_U433 & new_P1_R1138_U432;
  assign new_P1_R1138_U153 = ~new_P1_R1138_U286 | ~new_P1_R1138_U285;
  assign new_P1_R1138_U154 = new_P1_R1138_U440 & new_P1_R1138_U439;
  assign new_P1_R1138_U155 = ~new_P1_R1138_U131 | ~new_P1_R1138_U281;
  assign new_P1_R1138_U156 = new_P1_R1138_U447 & new_P1_R1138_U446;
  assign new_P1_R1138_U157 = new_P1_R1138_U452 & new_P1_R1138_U451;
  assign new_P1_R1138_U158 = ~new_P1_R1138_U44 | ~new_P1_R1138_U324;
  assign new_P1_R1138_U159 = ~new_P1_R1138_U129 | ~new_P1_R1138_U266;
  assign new_P1_R1138_U160 = new_P1_R1138_U473 & new_P1_R1138_U472;
  assign new_P1_R1138_U161 = ~new_P1_R1138_U254 | ~new_P1_R1138_U253;
  assign new_P1_R1138_U162 = new_P1_R1138_U480 & new_P1_R1138_U479;
  assign new_P1_R1138_U163 = ~new_P1_R1138_U250 | ~new_P1_R1138_U249;
  assign new_P1_R1138_U164 = ~new_P1_R1138_U240 | ~new_P1_R1138_U239;
  assign new_P1_R1138_U165 = ~new_P1_R1138_U364 | ~new_P1_R1138_U363;
  assign new_P1_R1138_U166 = ~new_P1_U3054 | ~new_P1_R1138_U147;
  assign new_P1_R1138_U167 = ~new_P1_R1138_U35;
  assign new_P1_R1138_U168 = ~new_P1_U3485 | ~new_P1_U3083;
  assign new_P1_R1138_U169 = ~new_P1_U3072 | ~new_P1_U3494;
  assign new_P1_R1138_U170 = ~new_P1_U3058 | ~new_P1_U4020;
  assign new_P1_R1138_U171 = ~new_P1_R1138_U69;
  assign new_P1_R1138_U172 = ~new_P1_R1138_U78;
  assign new_P1_R1138_U173 = ~new_P1_U3065 | ~new_P1_U4021;
  assign new_P1_R1138_U174 = ~new_P1_R1138_U62;
  assign new_P1_R1138_U175 = new_P1_U3067 | new_P1_U3473;
  assign new_P1_R1138_U176 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1138_U177 = new_P1_U3467 | new_P1_U3064;
  assign new_P1_R1138_U178 = new_P1_U3464 | new_P1_U3068;
  assign new_P1_R1138_U179 = ~new_P1_R1138_U32;
  assign new_P1_R1138_U180 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1138_U181 = ~new_P1_R1138_U43;
  assign new_P1_R1138_U182 = ~new_P1_R1138_U44;
  assign new_P1_R1138_U183 = ~new_P1_R1138_U43 | ~new_P1_R1138_U44;
  assign new_P1_R1138_U184 = ~new_P1_R1138_U116 | ~new_P1_R1138_U177;
  assign new_P1_R1138_U185 = ~new_P1_R1138_U5 | ~new_P1_R1138_U183;
  assign new_P1_R1138_U186 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1138_U187 = ~new_P1_R1138_U117 | ~new_P1_R1138_U185;
  assign new_P1_R1138_U188 = ~new_P1_R1138_U36 | ~new_P1_R1138_U35;
  assign new_P1_R1138_U189 = ~new_P1_U3067 | ~new_P1_R1138_U188;
  assign new_P1_R1138_U190 = ~new_P1_R1138_U4 | ~new_P1_R1138_U187;
  assign new_P1_R1138_U191 = ~new_P1_U3473 | ~new_P1_R1138_U167;
  assign new_P1_R1138_U192 = ~new_P1_R1138_U42;
  assign new_P1_R1138_U193 = new_P1_U3070 | new_P1_U3479;
  assign new_P1_R1138_U194 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1138_U195 = ~new_P1_R1138_U23;
  assign new_P1_R1138_U196 = ~new_P1_R1138_U24 | ~new_P1_R1138_U23;
  assign new_P1_R1138_U197 = ~new_P1_U3070 | ~new_P1_R1138_U196;
  assign new_P1_R1138_U198 = ~new_P1_U3479 | ~new_P1_R1138_U195;
  assign new_P1_R1138_U199 = ~new_P1_R1138_U6 | ~new_P1_R1138_U42;
  assign new_P1_R1138_U200 = ~new_P1_R1138_U140;
  assign new_P1_R1138_U201 = new_P1_U3482 | new_P1_U3084;
  assign new_P1_R1138_U202 = ~new_P1_R1138_U201 | ~new_P1_R1138_U140;
  assign new_P1_R1138_U203 = ~new_P1_R1138_U41;
  assign new_P1_R1138_U204 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1138_U205 = new_P1_U3476 | new_P1_U3071;
  assign new_P1_R1138_U206 = ~new_P1_R1138_U205 | ~new_P1_R1138_U42;
  assign new_P1_R1138_U207 = ~new_P1_R1138_U120 | ~new_P1_R1138_U206;
  assign new_P1_R1138_U208 = ~new_P1_R1138_U192 | ~new_P1_R1138_U23;
  assign new_P1_R1138_U209 = ~new_P1_U3479 | ~new_P1_U3070;
  assign new_P1_R1138_U210 = ~new_P1_R1138_U121 | ~new_P1_R1138_U208;
  assign new_P1_R1138_U211 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1138_U212 = ~new_P1_R1138_U182 | ~new_P1_R1138_U178;
  assign new_P1_R1138_U213 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1138_U214 = ~new_P1_R1138_U46;
  assign new_P1_R1138_U215 = ~new_P1_R1138_U181 | ~new_P1_R1138_U5;
  assign new_P1_R1138_U216 = ~new_P1_R1138_U46 | ~new_P1_R1138_U177;
  assign new_P1_R1138_U217 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1138_U218 = ~new_P1_R1138_U45;
  assign new_P1_R1138_U219 = new_P1_U3470 | new_P1_U3060;
  assign new_P1_R1138_U220 = ~new_P1_R1138_U219 | ~new_P1_R1138_U45;
  assign new_P1_R1138_U221 = ~new_P1_R1138_U123 | ~new_P1_R1138_U220;
  assign new_P1_R1138_U222 = ~new_P1_R1138_U218 | ~new_P1_R1138_U35;
  assign new_P1_R1138_U223 = ~new_P1_U3473 | ~new_P1_U3067;
  assign new_P1_R1138_U224 = ~new_P1_R1138_U124 | ~new_P1_R1138_U222;
  assign new_P1_R1138_U225 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1138_U226 = ~new_P1_R1138_U181 | ~new_P1_R1138_U178;
  assign new_P1_R1138_U227 = ~new_P1_R1138_U141;
  assign new_P1_R1138_U228 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1138_U229 = ~new_P1_R1138_U43 | ~new_P1_R1138_U44 | ~new_P1_R1138_U398 | ~new_P1_R1138_U397;
  assign new_P1_R1138_U230 = ~new_P1_R1138_U44 | ~new_P1_R1138_U43;
  assign new_P1_R1138_U231 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1138_U232 = ~new_P1_R1138_U125 | ~new_P1_R1138_U230;
  assign new_P1_R1138_U233 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1138_U234 = new_P1_U3062 | new_P1_U3488;
  assign new_P1_R1138_U235 = ~new_P1_R1138_U174 | ~new_P1_R1138_U7;
  assign new_P1_R1138_U236 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1138_U237 = ~new_P1_R1138_U127 | ~new_P1_R1138_U235;
  assign new_P1_R1138_U238 = new_P1_U3488 | new_P1_U3062;
  assign new_P1_R1138_U239 = ~new_P1_R1138_U126 | ~new_P1_R1138_U140;
  assign new_P1_R1138_U240 = ~new_P1_R1138_U238 | ~new_P1_R1138_U237;
  assign new_P1_R1138_U241 = ~new_P1_R1138_U164;
  assign new_P1_R1138_U242 = new_P1_U3080 | new_P1_U3497;
  assign new_P1_R1138_U243 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1138_U244 = ~new_P1_R1138_U171 | ~new_P1_R1138_U8;
  assign new_P1_R1138_U245 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1138_U246 = ~new_P1_R1138_U128 | ~new_P1_R1138_U244;
  assign new_P1_R1138_U247 = new_P1_U3491 | new_P1_U3063;
  assign new_P1_R1138_U248 = new_P1_U3497 | new_P1_U3080;
  assign new_P1_R1138_U249 = ~new_P1_R1138_U8 | ~new_P1_R1138_U247 | ~new_P1_R1138_U164;
  assign new_P1_R1138_U250 = ~new_P1_R1138_U248 | ~new_P1_R1138_U246;
  assign new_P1_R1138_U251 = ~new_P1_R1138_U163;
  assign new_P1_R1138_U252 = new_P1_U3500 | new_P1_U3079;
  assign new_P1_R1138_U253 = ~new_P1_R1138_U252 | ~new_P1_R1138_U163;
  assign new_P1_R1138_U254 = ~new_P1_U3079 | ~new_P1_U3500;
  assign new_P1_R1138_U255 = ~new_P1_R1138_U161;
  assign new_P1_R1138_U256 = new_P1_U3503 | new_P1_U3074;
  assign new_P1_R1138_U257 = ~new_P1_R1138_U256 | ~new_P1_R1138_U161;
  assign new_P1_R1138_U258 = ~new_P1_U3074 | ~new_P1_U3503;
  assign new_P1_R1138_U259 = ~new_P1_R1138_U93;
  assign new_P1_R1138_U260 = new_P1_U3069 | new_P1_U3509;
  assign new_P1_R1138_U261 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1138_U262 = ~new_P1_R1138_U60;
  assign new_P1_R1138_U263 = ~new_P1_R1138_U61 | ~new_P1_R1138_U60;
  assign new_P1_R1138_U264 = ~new_P1_U3069 | ~new_P1_R1138_U263;
  assign new_P1_R1138_U265 = ~new_P1_U3509 | ~new_P1_R1138_U262;
  assign new_P1_R1138_U266 = ~new_P1_R1138_U9 | ~new_P1_R1138_U93;
  assign new_P1_R1138_U267 = ~new_P1_R1138_U159;
  assign new_P1_R1138_U268 = new_P1_U3076 | new_P1_U4025;
  assign new_P1_R1138_U269 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1138_U270 = new_P1_U3075 | new_P1_U4024;
  assign new_P1_R1138_U271 = ~new_P1_R1138_U81;
  assign new_P1_R1138_U272 = ~new_P1_U4025 | ~new_P1_R1138_U271;
  assign new_P1_R1138_U273 = ~new_P1_R1138_U272 | ~new_P1_R1138_U91;
  assign new_P1_R1138_U274 = ~new_P1_R1138_U81 | ~new_P1_R1138_U82;
  assign new_P1_R1138_U275 = ~new_P1_R1138_U274 | ~new_P1_R1138_U273;
  assign new_P1_R1138_U276 = ~new_P1_R1138_U172 | ~new_P1_R1138_U10;
  assign new_P1_R1138_U277 = ~new_P1_U3075 | ~new_P1_U4024;
  assign new_P1_R1138_U278 = ~new_P1_R1138_U275 | ~new_P1_R1138_U276;
  assign new_P1_R1138_U279 = new_P1_U3512 | new_P1_U3082;
  assign new_P1_R1138_U280 = new_P1_U4024 | new_P1_U3075;
  assign new_P1_R1138_U281 = ~new_P1_R1138_U130 | ~new_P1_R1138_U270 | ~new_P1_R1138_U159;
  assign new_P1_R1138_U282 = ~new_P1_R1138_U280 | ~new_P1_R1138_U278;
  assign new_P1_R1138_U283 = ~new_P1_R1138_U155;
  assign new_P1_R1138_U284 = new_P1_U4023 | new_P1_U3061;
  assign new_P1_R1138_U285 = ~new_P1_R1138_U284 | ~new_P1_R1138_U155;
  assign new_P1_R1138_U286 = ~new_P1_U3061 | ~new_P1_U4023;
  assign new_P1_R1138_U287 = ~new_P1_R1138_U153;
  assign new_P1_R1138_U288 = new_P1_U4022 | new_P1_U3066;
  assign new_P1_R1138_U289 = ~new_P1_R1138_U288 | ~new_P1_R1138_U153;
  assign new_P1_R1138_U290 = ~new_P1_U3066 | ~new_P1_U4022;
  assign new_P1_R1138_U291 = ~new_P1_R1138_U151;
  assign new_P1_R1138_U292 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1138_U293 = ~new_P1_R1138_U173 | ~new_P1_R1138_U170;
  assign new_P1_R1138_U294 = ~new_P1_R1138_U87;
  assign new_P1_R1138_U295 = new_P1_U4021 | new_P1_U3065;
  assign new_P1_R1138_U296 = ~new_P1_R1138_U165 | ~new_P1_R1138_U151 | ~new_P1_R1138_U295;
  assign new_P1_R1138_U297 = ~new_P1_R1138_U149;
  assign new_P1_R1138_U298 = new_P1_U4018 | new_P1_U3053;
  assign new_P1_R1138_U299 = ~new_P1_U3053 | ~new_P1_U4018;
  assign new_P1_R1138_U300 = ~new_P1_R1138_U147;
  assign new_P1_R1138_U301 = ~new_P1_U4017 | ~new_P1_R1138_U147;
  assign new_P1_R1138_U302 = ~new_P1_R1138_U145;
  assign new_P1_R1138_U303 = ~new_P1_R1138_U295 | ~new_P1_R1138_U151;
  assign new_P1_R1138_U304 = ~new_P1_R1138_U90;
  assign new_P1_R1138_U305 = new_P1_U4020 | new_P1_U3058;
  assign new_P1_R1138_U306 = ~new_P1_R1138_U305 | ~new_P1_R1138_U90;
  assign new_P1_R1138_U307 = ~new_P1_R1138_U150 | ~new_P1_R1138_U306 | ~new_P1_R1138_U170;
  assign new_P1_R1138_U308 = ~new_P1_R1138_U304 | ~new_P1_R1138_U170;
  assign new_P1_R1138_U309 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1138_U310 = ~new_P1_R1138_U165 | ~new_P1_R1138_U308 | ~new_P1_R1138_U309;
  assign new_P1_R1138_U311 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1138_U312 = ~new_P1_R1138_U279 | ~new_P1_R1138_U159;
  assign new_P1_R1138_U313 = ~new_P1_R1138_U92;
  assign new_P1_R1138_U314 = ~new_P1_R1138_U10 | ~new_P1_R1138_U92;
  assign new_P1_R1138_U315 = ~new_P1_R1138_U134 | ~new_P1_R1138_U314;
  assign new_P1_R1138_U316 = ~new_P1_R1138_U314 | ~new_P1_R1138_U275;
  assign new_P1_R1138_U317 = ~new_P1_R1138_U450 | ~new_P1_R1138_U316;
  assign new_P1_R1138_U318 = new_P1_U3514 | new_P1_U3081;
  assign new_P1_R1138_U319 = ~new_P1_R1138_U318 | ~new_P1_R1138_U92;
  assign new_P1_R1138_U320 = ~new_P1_R1138_U157 | ~new_P1_R1138_U319 | ~new_P1_R1138_U81;
  assign new_P1_R1138_U321 = ~new_P1_R1138_U313 | ~new_P1_R1138_U81;
  assign new_P1_R1138_U322 = ~new_P1_U3076 | ~new_P1_U4025;
  assign new_P1_R1138_U323 = ~new_P1_R1138_U10 | ~new_P1_R1138_U322 | ~new_P1_R1138_U321;
  assign new_P1_R1138_U324 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1138_U325 = ~new_P1_R1138_U158;
  assign new_P1_R1138_U326 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1138_U327 = new_P1_U3506 | new_P1_U3073;
  assign new_P1_R1138_U328 = ~new_P1_R1138_U327 | ~new_P1_R1138_U93;
  assign new_P1_R1138_U329 = ~new_P1_R1138_U135 | ~new_P1_R1138_U328;
  assign new_P1_R1138_U330 = ~new_P1_R1138_U259 | ~new_P1_R1138_U60;
  assign new_P1_R1138_U331 = ~new_P1_U3509 | ~new_P1_U3069;
  assign new_P1_R1138_U332 = ~new_P1_R1138_U9 | ~new_P1_R1138_U331 | ~new_P1_R1138_U330;
  assign new_P1_R1138_U333 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1138_U334 = ~new_P1_R1138_U247 | ~new_P1_R1138_U164;
  assign new_P1_R1138_U335 = ~new_P1_R1138_U94;
  assign new_P1_R1138_U336 = new_P1_U3494 | new_P1_U3072;
  assign new_P1_R1138_U337 = ~new_P1_R1138_U336 | ~new_P1_R1138_U94;
  assign new_P1_R1138_U338 = ~new_P1_R1138_U136 | ~new_P1_R1138_U337;
  assign new_P1_R1138_U339 = ~new_P1_R1138_U335 | ~new_P1_R1138_U169;
  assign new_P1_R1138_U340 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1138_U341 = ~new_P1_R1138_U137 | ~new_P1_R1138_U339;
  assign new_P1_R1138_U342 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1138_U343 = new_P1_U3485 | new_P1_U3083;
  assign new_P1_R1138_U344 = ~new_P1_R1138_U343 | ~new_P1_R1138_U41;
  assign new_P1_R1138_U345 = ~new_P1_R1138_U138 | ~new_P1_R1138_U344;
  assign new_P1_R1138_U346 = ~new_P1_R1138_U203 | ~new_P1_R1138_U168;
  assign new_P1_R1138_U347 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1138_U348 = ~new_P1_R1138_U139 | ~new_P1_R1138_U346;
  assign new_P1_R1138_U349 = ~new_P1_R1138_U204 | ~new_P1_R1138_U168;
  assign new_P1_R1138_U350 = ~new_P1_R1138_U201 | ~new_P1_R1138_U62;
  assign new_P1_R1138_U351 = ~new_P1_R1138_U211 | ~new_P1_R1138_U23;
  assign new_P1_R1138_U352 = ~new_P1_R1138_U225 | ~new_P1_R1138_U35;
  assign new_P1_R1138_U353 = ~new_P1_R1138_U228 | ~new_P1_R1138_U177;
  assign new_P1_R1138_U354 = ~new_P1_R1138_U311 | ~new_P1_R1138_U170;
  assign new_P1_R1138_U355 = ~new_P1_R1138_U295 | ~new_P1_R1138_U173;
  assign new_P1_R1138_U356 = ~new_P1_R1138_U326 | ~new_P1_R1138_U81;
  assign new_P1_R1138_U357 = ~new_P1_R1138_U279 | ~new_P1_R1138_U78;
  assign new_P1_R1138_U358 = ~new_P1_R1138_U333 | ~new_P1_R1138_U60;
  assign new_P1_R1138_U359 = ~new_P1_R1138_U342 | ~new_P1_R1138_U169;
  assign new_P1_R1138_U360 = ~new_P1_R1138_U247 | ~new_P1_R1138_U69;
  assign new_P1_R1138_U361 = ~new_P1_U4017 | ~new_P1_U3054;
  assign new_P1_R1138_U362 = ~new_P1_R1138_U293 | ~new_P1_R1138_U165;
  assign new_P1_R1138_U363 = ~new_P1_U3057 | ~new_P1_R1138_U292;
  assign new_P1_R1138_U364 = ~new_P1_U4019 | ~new_P1_R1138_U292;
  assign new_P1_R1138_U365 = ~new_P1_R1138_U298 | ~new_P1_R1138_U293 | ~new_P1_R1138_U165;
  assign new_P1_R1138_U366 = ~new_P1_R1138_U132 | ~new_P1_R1138_U151 | ~new_P1_R1138_U165;
  assign new_P1_R1138_U367 = ~new_P1_R1138_U294 | ~new_P1_R1138_U298;
  assign new_P1_R1138_U368 = ~new_P1_U3083 | ~new_P1_R1138_U40;
  assign new_P1_R1138_U369 = ~new_P1_U3485 | ~new_P1_R1138_U39;
  assign new_P1_R1138_U370 = ~new_P1_R1138_U369 | ~new_P1_R1138_U368;
  assign new_P1_R1138_U371 = ~new_P1_R1138_U349 | ~new_P1_R1138_U41;
  assign new_P1_R1138_U372 = ~new_P1_R1138_U370 | ~new_P1_R1138_U203;
  assign new_P1_R1138_U373 = ~new_P1_U3084 | ~new_P1_R1138_U37;
  assign new_P1_R1138_U374 = ~new_P1_U3482 | ~new_P1_R1138_U38;
  assign new_P1_R1138_U375 = ~new_P1_R1138_U374 | ~new_P1_R1138_U373;
  assign new_P1_R1138_U376 = ~new_P1_R1138_U350 | ~new_P1_R1138_U140;
  assign new_P1_R1138_U377 = ~new_P1_R1138_U200 | ~new_P1_R1138_U375;
  assign new_P1_R1138_U378 = ~new_P1_U3070 | ~new_P1_R1138_U24;
  assign new_P1_R1138_U379 = ~new_P1_U3479 | ~new_P1_R1138_U22;
  assign new_P1_R1138_U380 = ~new_P1_U3071 | ~new_P1_R1138_U20;
  assign new_P1_R1138_U381 = ~new_P1_U3476 | ~new_P1_R1138_U21;
  assign new_P1_R1138_U382 = ~new_P1_R1138_U381 | ~new_P1_R1138_U380;
  assign new_P1_R1138_U383 = ~new_P1_R1138_U351 | ~new_P1_R1138_U42;
  assign new_P1_R1138_U384 = ~new_P1_R1138_U382 | ~new_P1_R1138_U192;
  assign new_P1_R1138_U385 = ~new_P1_U3067 | ~new_P1_R1138_U36;
  assign new_P1_R1138_U386 = ~new_P1_U3473 | ~new_P1_R1138_U27;
  assign new_P1_R1138_U387 = ~new_P1_U3060 | ~new_P1_R1138_U25;
  assign new_P1_R1138_U388 = ~new_P1_U3470 | ~new_P1_R1138_U26;
  assign new_P1_R1138_U389 = ~new_P1_R1138_U388 | ~new_P1_R1138_U387;
  assign new_P1_R1138_U390 = ~new_P1_R1138_U352 | ~new_P1_R1138_U45;
  assign new_P1_R1138_U391 = ~new_P1_R1138_U389 | ~new_P1_R1138_U218;
  assign new_P1_R1138_U392 = ~new_P1_U3064 | ~new_P1_R1138_U33;
  assign new_P1_R1138_U393 = ~new_P1_U3467 | ~new_P1_R1138_U34;
  assign new_P1_R1138_U394 = ~new_P1_R1138_U393 | ~new_P1_R1138_U392;
  assign new_P1_R1138_U395 = ~new_P1_R1138_U353 | ~new_P1_R1138_U141;
  assign new_P1_R1138_U396 = ~new_P1_R1138_U227 | ~new_P1_R1138_U394;
  assign new_P1_R1138_U397 = ~new_P1_U3068 | ~new_P1_R1138_U28;
  assign new_P1_R1138_U398 = ~new_P1_U3464 | ~new_P1_R1138_U29;
  assign new_P1_R1138_U399 = ~new_P1_U3055 | ~new_P1_R1138_U143;
  assign new_P1_R1138_U400 = ~new_P1_U4028 | ~new_P1_R1138_U142;
  assign new_P1_R1138_U401 = ~new_P1_U3055 | ~new_P1_R1138_U143;
  assign new_P1_R1138_U402 = ~new_P1_U4028 | ~new_P1_R1138_U142;
  assign new_P1_R1138_U403 = ~new_P1_R1138_U402 | ~new_P1_R1138_U401;
  assign new_P1_R1138_U404 = ~new_P1_R1138_U144 | ~new_P1_R1138_U145;
  assign new_P1_R1138_U405 = ~new_P1_R1138_U302 | ~new_P1_R1138_U403;
  assign new_P1_R1138_U406 = ~new_P1_U3054 | ~new_P1_R1138_U89;
  assign new_P1_R1138_U407 = ~new_P1_U4017 | ~new_P1_R1138_U88;
  assign new_P1_R1138_U408 = ~new_P1_U3054 | ~new_P1_R1138_U89;
  assign new_P1_R1138_U409 = ~new_P1_U4017 | ~new_P1_R1138_U88;
  assign new_P1_R1138_U410 = ~new_P1_R1138_U409 | ~new_P1_R1138_U408;
  assign new_P1_R1138_U411 = ~new_P1_R1138_U146 | ~new_P1_R1138_U147;
  assign new_P1_R1138_U412 = ~new_P1_R1138_U300 | ~new_P1_R1138_U410;
  assign new_P1_R1138_U413 = ~new_P1_U3053 | ~new_P1_R1138_U47;
  assign new_P1_R1138_U414 = ~new_P1_U4018 | ~new_P1_R1138_U48;
  assign new_P1_R1138_U415 = ~new_P1_U3053 | ~new_P1_R1138_U47;
  assign new_P1_R1138_U416 = ~new_P1_U4018 | ~new_P1_R1138_U48;
  assign new_P1_R1138_U417 = ~new_P1_R1138_U416 | ~new_P1_R1138_U415;
  assign new_P1_R1138_U418 = ~new_P1_R1138_U148 | ~new_P1_R1138_U149;
  assign new_P1_R1138_U419 = ~new_P1_R1138_U297 | ~new_P1_R1138_U417;
  assign new_P1_R1138_U420 = ~new_P1_U3057 | ~new_P1_R1138_U50;
  assign new_P1_R1138_U421 = ~new_P1_U4019 | ~new_P1_R1138_U49;
  assign new_P1_R1138_U422 = ~new_P1_U3058 | ~new_P1_R1138_U51;
  assign new_P1_R1138_U423 = ~new_P1_U4020 | ~new_P1_R1138_U52;
  assign new_P1_R1138_U424 = ~new_P1_R1138_U423 | ~new_P1_R1138_U422;
  assign new_P1_R1138_U425 = ~new_P1_R1138_U354 | ~new_P1_R1138_U90;
  assign new_P1_R1138_U426 = ~new_P1_R1138_U424 | ~new_P1_R1138_U304;
  assign new_P1_R1138_U427 = ~new_P1_U3065 | ~new_P1_R1138_U53;
  assign new_P1_R1138_U428 = ~new_P1_U4021 | ~new_P1_R1138_U54;
  assign new_P1_R1138_U429 = ~new_P1_R1138_U428 | ~new_P1_R1138_U427;
  assign new_P1_R1138_U430 = ~new_P1_R1138_U355 | ~new_P1_R1138_U151;
  assign new_P1_R1138_U431 = ~new_P1_R1138_U291 | ~new_P1_R1138_U429;
  assign new_P1_R1138_U432 = ~new_P1_U3066 | ~new_P1_R1138_U85;
  assign new_P1_R1138_U433 = ~new_P1_U4022 | ~new_P1_R1138_U86;
  assign new_P1_R1138_U434 = ~new_P1_U3066 | ~new_P1_R1138_U85;
  assign new_P1_R1138_U435 = ~new_P1_U4022 | ~new_P1_R1138_U86;
  assign new_P1_R1138_U436 = ~new_P1_R1138_U435 | ~new_P1_R1138_U434;
  assign new_P1_R1138_U437 = ~new_P1_R1138_U152 | ~new_P1_R1138_U153;
  assign new_P1_R1138_U438 = ~new_P1_R1138_U287 | ~new_P1_R1138_U436;
  assign new_P1_R1138_U439 = ~new_P1_U3061 | ~new_P1_R1138_U83;
  assign new_P1_R1138_U440 = ~new_P1_U4023 | ~new_P1_R1138_U84;
  assign new_P1_R1138_U441 = ~new_P1_U3061 | ~new_P1_R1138_U83;
  assign new_P1_R1138_U442 = ~new_P1_U4023 | ~new_P1_R1138_U84;
  assign new_P1_R1138_U443 = ~new_P1_R1138_U442 | ~new_P1_R1138_U441;
  assign new_P1_R1138_U444 = ~new_P1_R1138_U154 | ~new_P1_R1138_U155;
  assign new_P1_R1138_U445 = ~new_P1_R1138_U283 | ~new_P1_R1138_U443;
  assign new_P1_R1138_U446 = ~new_P1_U3075 | ~new_P1_R1138_U55;
  assign new_P1_R1138_U447 = ~new_P1_U4024 | ~new_P1_R1138_U56;
  assign new_P1_R1138_U448 = ~new_P1_U3075 | ~new_P1_R1138_U55;
  assign new_P1_R1138_U449 = ~new_P1_U4024 | ~new_P1_R1138_U56;
  assign new_P1_R1138_U450 = ~new_P1_R1138_U449 | ~new_P1_R1138_U448;
  assign new_P1_R1138_U451 = ~new_P1_U3076 | ~new_P1_R1138_U82;
  assign new_P1_R1138_U452 = ~new_P1_U4025 | ~new_P1_R1138_U91;
  assign new_P1_R1138_U453 = ~new_P1_R1138_U179 | ~new_P1_R1138_U158;
  assign new_P1_R1138_U454 = ~new_P1_R1138_U325 | ~new_P1_R1138_U32;
  assign new_P1_R1138_U455 = ~new_P1_U3081 | ~new_P1_R1138_U79;
  assign new_P1_R1138_U456 = ~new_P1_U3514 | ~new_P1_R1138_U80;
  assign new_P1_R1138_U457 = ~new_P1_R1138_U456 | ~new_P1_R1138_U455;
  assign new_P1_R1138_U458 = ~new_P1_R1138_U356 | ~new_P1_R1138_U92;
  assign new_P1_R1138_U459 = ~new_P1_R1138_U457 | ~new_P1_R1138_U313;
  assign new_P1_R1138_U460 = ~new_P1_U3082 | ~new_P1_R1138_U76;
  assign new_P1_R1138_U461 = ~new_P1_U3512 | ~new_P1_R1138_U77;
  assign new_P1_R1138_U462 = ~new_P1_R1138_U461 | ~new_P1_R1138_U460;
  assign new_P1_R1138_U463 = ~new_P1_R1138_U357 | ~new_P1_R1138_U159;
  assign new_P1_R1138_U464 = ~new_P1_R1138_U267 | ~new_P1_R1138_U462;
  assign new_P1_R1138_U465 = ~new_P1_U3069 | ~new_P1_R1138_U61;
  assign new_P1_R1138_U466 = ~new_P1_U3509 | ~new_P1_R1138_U59;
  assign new_P1_R1138_U467 = ~new_P1_U3073 | ~new_P1_R1138_U57;
  assign new_P1_R1138_U468 = ~new_P1_U3506 | ~new_P1_R1138_U58;
  assign new_P1_R1138_U469 = ~new_P1_R1138_U468 | ~new_P1_R1138_U467;
  assign new_P1_R1138_U470 = ~new_P1_R1138_U358 | ~new_P1_R1138_U93;
  assign new_P1_R1138_U471 = ~new_P1_R1138_U469 | ~new_P1_R1138_U259;
  assign new_P1_R1138_U472 = ~new_P1_U3074 | ~new_P1_R1138_U74;
  assign new_P1_R1138_U473 = ~new_P1_U3503 | ~new_P1_R1138_U75;
  assign new_P1_R1138_U474 = ~new_P1_U3074 | ~new_P1_R1138_U74;
  assign new_P1_R1138_U475 = ~new_P1_U3503 | ~new_P1_R1138_U75;
  assign new_P1_R1138_U476 = ~new_P1_R1138_U475 | ~new_P1_R1138_U474;
  assign new_P1_R1138_U477 = ~new_P1_R1138_U160 | ~new_P1_R1138_U161;
  assign new_P1_R1138_U478 = ~new_P1_R1138_U255 | ~new_P1_R1138_U476;
  assign new_P1_R1138_U479 = ~new_P1_U3079 | ~new_P1_R1138_U72;
  assign new_P1_R1138_U480 = ~new_P1_U3500 | ~new_P1_R1138_U73;
  assign new_P1_R1138_U481 = ~new_P1_U3079 | ~new_P1_R1138_U72;
  assign new_P1_R1138_U482 = ~new_P1_U3500 | ~new_P1_R1138_U73;
  assign new_P1_R1138_U483 = ~new_P1_R1138_U482 | ~new_P1_R1138_U481;
  assign new_P1_R1138_U484 = ~new_P1_R1138_U162 | ~new_P1_R1138_U163;
  assign new_P1_R1138_U485 = ~new_P1_R1138_U251 | ~new_P1_R1138_U483;
  assign new_P1_R1138_U486 = ~new_P1_U3080 | ~new_P1_R1138_U70;
  assign new_P1_R1138_U487 = ~new_P1_U3497 | ~new_P1_R1138_U71;
  assign new_P1_R1138_U488 = ~new_P1_U3072 | ~new_P1_R1138_U65;
  assign new_P1_R1138_U489 = ~new_P1_U3494 | ~new_P1_R1138_U66;
  assign new_P1_R1138_U490 = ~new_P1_R1138_U489 | ~new_P1_R1138_U488;
  assign new_P1_R1138_U491 = ~new_P1_R1138_U359 | ~new_P1_R1138_U94;
  assign new_P1_R1138_U492 = ~new_P1_R1138_U490 | ~new_P1_R1138_U335;
  assign new_P1_R1138_U493 = ~new_P1_U3063 | ~new_P1_R1138_U67;
  assign new_P1_R1138_U494 = ~new_P1_U3491 | ~new_P1_R1138_U68;
  assign new_P1_R1138_U495 = ~new_P1_R1138_U494 | ~new_P1_R1138_U493;
  assign new_P1_R1138_U496 = ~new_P1_R1138_U360 | ~new_P1_R1138_U164;
  assign new_P1_R1138_U497 = ~new_P1_R1138_U241 | ~new_P1_R1138_U495;
  assign new_P1_R1138_U498 = ~new_P1_U3062 | ~new_P1_R1138_U63;
  assign new_P1_R1138_U499 = ~new_P1_U3488 | ~new_P1_R1138_U64;
  assign new_P1_R1138_U500 = ~new_P1_U3077 | ~new_P1_R1138_U30;
  assign new_P1_R1138_U501 = ~new_P1_U3456 | ~new_P1_R1138_U31;
  assign new_P1_R1222_U4 = new_P1_R1222_U176 & new_P1_R1222_U175;
  assign new_P1_R1222_U5 = new_P1_R1222_U177 & new_P1_R1222_U178;
  assign new_P1_R1222_U6 = new_P1_R1222_U194 & new_P1_R1222_U193;
  assign new_P1_R1222_U7 = new_P1_R1222_U234 & new_P1_R1222_U233;
  assign new_P1_R1222_U8 = new_P1_R1222_U243 & new_P1_R1222_U242;
  assign new_P1_R1222_U9 = new_P1_R1222_U261 & new_P1_R1222_U260;
  assign new_P1_R1222_U10 = new_P1_R1222_U269 & new_P1_R1222_U268;
  assign new_P1_R1222_U11 = new_P1_R1222_U348 & new_P1_R1222_U345;
  assign new_P1_R1222_U12 = new_P1_R1222_U341 & new_P1_R1222_U338;
  assign new_P1_R1222_U13 = new_P1_R1222_U332 & new_P1_R1222_U329;
  assign new_P1_R1222_U14 = new_P1_R1222_U323 & new_P1_R1222_U320;
  assign new_P1_R1222_U15 = new_P1_R1222_U317 & new_P1_R1222_U315;
  assign new_P1_R1222_U16 = new_P1_R1222_U310 & new_P1_R1222_U307;
  assign new_P1_R1222_U17 = new_P1_R1222_U232 & new_P1_R1222_U229;
  assign new_P1_R1222_U18 = new_P1_R1222_U224 & new_P1_R1222_U221;
  assign new_P1_R1222_U19 = new_P1_R1222_U210 & new_P1_R1222_U207;
  assign new_P1_R1222_U20 = ~new_P1_U3476;
  assign new_P1_R1222_U21 = ~new_P1_U3071;
  assign new_P1_R1222_U22 = ~new_P1_U3070;
  assign new_P1_R1222_U23 = ~new_P1_U3071 | ~new_P1_U3476;
  assign new_P1_R1222_U24 = ~new_P1_U3479;
  assign new_P1_R1222_U25 = ~new_P1_U3470;
  assign new_P1_R1222_U26 = ~new_P1_U3060;
  assign new_P1_R1222_U27 = ~new_P1_U3067;
  assign new_P1_R1222_U28 = ~new_P1_U3464;
  assign new_P1_R1222_U29 = ~new_P1_U3068;
  assign new_P1_R1222_U30 = ~new_P1_U3456;
  assign new_P1_R1222_U31 = ~new_P1_U3077;
  assign new_P1_R1222_U32 = ~new_P1_U3077 | ~new_P1_U3456;
  assign new_P1_R1222_U33 = ~new_P1_U3467;
  assign new_P1_R1222_U34 = ~new_P1_U3064;
  assign new_P1_R1222_U35 = ~new_P1_U3060 | ~new_P1_U3470;
  assign new_P1_R1222_U36 = ~new_P1_U3473;
  assign new_P1_R1222_U37 = ~new_P1_U3482;
  assign new_P1_R1222_U38 = ~new_P1_U3084;
  assign new_P1_R1222_U39 = ~new_P1_U3083;
  assign new_P1_R1222_U40 = ~new_P1_U3485;
  assign new_P1_R1222_U41 = ~new_P1_R1222_U62 | ~new_P1_R1222_U202;
  assign new_P1_R1222_U42 = ~new_P1_R1222_U118 | ~new_P1_R1222_U190;
  assign new_P1_R1222_U43 = ~new_P1_R1222_U179 | ~new_P1_R1222_U180;
  assign new_P1_R1222_U44 = ~new_P1_U3461 | ~new_P1_U3078;
  assign new_P1_R1222_U45 = ~new_P1_R1222_U122 | ~new_P1_R1222_U216;
  assign new_P1_R1222_U46 = ~new_P1_R1222_U213 | ~new_P1_R1222_U212;
  assign new_P1_R1222_U47 = ~new_P1_U4018;
  assign new_P1_R1222_U48 = ~new_P1_U3053;
  assign new_P1_R1222_U49 = ~new_P1_U3057;
  assign new_P1_R1222_U50 = ~new_P1_U4019;
  assign new_P1_R1222_U51 = ~new_P1_U4020;
  assign new_P1_R1222_U52 = ~new_P1_U3058;
  assign new_P1_R1222_U53 = ~new_P1_U4021;
  assign new_P1_R1222_U54 = ~new_P1_U3065;
  assign new_P1_R1222_U55 = ~new_P1_U4024;
  assign new_P1_R1222_U56 = ~new_P1_U3075;
  assign new_P1_R1222_U57 = ~new_P1_U3506;
  assign new_P1_R1222_U58 = ~new_P1_U3073;
  assign new_P1_R1222_U59 = ~new_P1_U3069;
  assign new_P1_R1222_U60 = ~new_P1_U3073 | ~new_P1_U3506;
  assign new_P1_R1222_U61 = ~new_P1_U3509;
  assign new_P1_R1222_U62 = ~new_P1_U3084 | ~new_P1_U3482;
  assign new_P1_R1222_U63 = ~new_P1_U3488;
  assign new_P1_R1222_U64 = ~new_P1_U3062;
  assign new_P1_R1222_U65 = ~new_P1_U3494;
  assign new_P1_R1222_U66 = ~new_P1_U3072;
  assign new_P1_R1222_U67 = ~new_P1_U3491;
  assign new_P1_R1222_U68 = ~new_P1_U3063;
  assign new_P1_R1222_U69 = ~new_P1_U3063 | ~new_P1_U3491;
  assign new_P1_R1222_U70 = ~new_P1_U3497;
  assign new_P1_R1222_U71 = ~new_P1_U3080;
  assign new_P1_R1222_U72 = ~new_P1_U3500;
  assign new_P1_R1222_U73 = ~new_P1_U3079;
  assign new_P1_R1222_U74 = ~new_P1_U3503;
  assign new_P1_R1222_U75 = ~new_P1_U3074;
  assign new_P1_R1222_U76 = ~new_P1_U3512;
  assign new_P1_R1222_U77 = ~new_P1_U3082;
  assign new_P1_R1222_U78 = ~new_P1_U3082 | ~new_P1_U3512;
  assign new_P1_R1222_U79 = ~new_P1_U3514;
  assign new_P1_R1222_U80 = ~new_P1_U3081;
  assign new_P1_R1222_U81 = ~new_P1_U3081 | ~new_P1_U3514;
  assign new_P1_R1222_U82 = ~new_P1_U4025;
  assign new_P1_R1222_U83 = ~new_P1_U4023;
  assign new_P1_R1222_U84 = ~new_P1_U3061;
  assign new_P1_R1222_U85 = ~new_P1_U4022;
  assign new_P1_R1222_U86 = ~new_P1_U3066;
  assign new_P1_R1222_U87 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1222_U88 = ~new_P1_U3054;
  assign new_P1_R1222_U89 = ~new_P1_U4017;
  assign new_P1_R1222_U90 = ~new_P1_R1222_U303 | ~new_P1_R1222_U173;
  assign new_P1_R1222_U91 = ~new_P1_U3076;
  assign new_P1_R1222_U92 = ~new_P1_R1222_U78 | ~new_P1_R1222_U312;
  assign new_P1_R1222_U93 = ~new_P1_R1222_U258 | ~new_P1_R1222_U257;
  assign new_P1_R1222_U94 = ~new_P1_R1222_U69 | ~new_P1_R1222_U334;
  assign new_P1_R1222_U95 = ~new_P1_R1222_U454 | ~new_P1_R1222_U453;
  assign new_P1_R1222_U96 = ~new_P1_R1222_U501 | ~new_P1_R1222_U500;
  assign new_P1_R1222_U97 = ~new_P1_R1222_U372 | ~new_P1_R1222_U371;
  assign new_P1_R1222_U98 = ~new_P1_R1222_U377 | ~new_P1_R1222_U376;
  assign new_P1_R1222_U99 = ~new_P1_R1222_U384 | ~new_P1_R1222_U383;
  assign new_P1_R1222_U100 = ~new_P1_R1222_U391 | ~new_P1_R1222_U390;
  assign new_P1_R1222_U101 = ~new_P1_R1222_U396 | ~new_P1_R1222_U395;
  assign new_P1_R1222_U102 = ~new_P1_R1222_U405 | ~new_P1_R1222_U404;
  assign new_P1_R1222_U103 = ~new_P1_R1222_U412 | ~new_P1_R1222_U411;
  assign new_P1_R1222_U104 = ~new_P1_R1222_U419 | ~new_P1_R1222_U418;
  assign new_P1_R1222_U105 = ~new_P1_R1222_U426 | ~new_P1_R1222_U425;
  assign new_P1_R1222_U106 = ~new_P1_R1222_U431 | ~new_P1_R1222_U430;
  assign new_P1_R1222_U107 = ~new_P1_R1222_U438 | ~new_P1_R1222_U437;
  assign new_P1_R1222_U108 = ~new_P1_R1222_U445 | ~new_P1_R1222_U444;
  assign new_P1_R1222_U109 = ~new_P1_R1222_U459 | ~new_P1_R1222_U458;
  assign new_P1_R1222_U110 = ~new_P1_R1222_U464 | ~new_P1_R1222_U463;
  assign new_P1_R1222_U111 = ~new_P1_R1222_U471 | ~new_P1_R1222_U470;
  assign new_P1_R1222_U112 = ~new_P1_R1222_U478 | ~new_P1_R1222_U477;
  assign new_P1_R1222_U113 = ~new_P1_R1222_U485 | ~new_P1_R1222_U484;
  assign new_P1_R1222_U114 = ~new_P1_R1222_U492 | ~new_P1_R1222_U491;
  assign new_P1_R1222_U115 = ~new_P1_R1222_U497 | ~new_P1_R1222_U496;
  assign new_P1_R1222_U116 = new_P1_U3464 & new_P1_U3068;
  assign new_P1_R1222_U117 = new_P1_R1222_U186 & new_P1_R1222_U184;
  assign new_P1_R1222_U118 = new_P1_R1222_U191 & new_P1_R1222_U189;
  assign new_P1_R1222_U119 = new_P1_R1222_U198 & new_P1_R1222_U197;
  assign new_P1_R1222_U120 = new_P1_R1222_U23 & new_P1_R1222_U379 & new_P1_R1222_U378;
  assign new_P1_R1222_U121 = new_P1_R1222_U209 & new_P1_R1222_U6;
  assign new_P1_R1222_U122 = new_P1_R1222_U217 & new_P1_R1222_U215;
  assign new_P1_R1222_U123 = new_P1_R1222_U35 & new_P1_R1222_U386 & new_P1_R1222_U385;
  assign new_P1_R1222_U124 = new_P1_R1222_U223 & new_P1_R1222_U4;
  assign new_P1_R1222_U125 = new_P1_R1222_U231 & new_P1_R1222_U178;
  assign new_P1_R1222_U126 = new_P1_R1222_U201 & new_P1_R1222_U7;
  assign new_P1_R1222_U127 = new_P1_R1222_U236 & new_P1_R1222_U168;
  assign new_P1_R1222_U128 = new_P1_R1222_U245 & new_P1_R1222_U169;
  assign new_P1_R1222_U129 = new_P1_R1222_U265 & new_P1_R1222_U264;
  assign new_P1_R1222_U130 = new_P1_R1222_U10 & new_P1_R1222_U279;
  assign new_P1_R1222_U131 = new_P1_R1222_U282 & new_P1_R1222_U277;
  assign new_P1_R1222_U132 = new_P1_R1222_U298 & new_P1_R1222_U295;
  assign new_P1_R1222_U133 = new_P1_R1222_U365 & new_P1_R1222_U299;
  assign new_P1_R1222_U134 = new_P1_R1222_U156 & new_P1_R1222_U275;
  assign new_P1_R1222_U135 = new_P1_R1222_U60 & new_P1_R1222_U466 & new_P1_R1222_U465;
  assign new_P1_R1222_U136 = new_P1_R1222_U169 & new_P1_R1222_U487 & new_P1_R1222_U486;
  assign new_P1_R1222_U137 = new_P1_R1222_U340 & new_P1_R1222_U8;
  assign new_P1_R1222_U138 = new_P1_R1222_U168 & new_P1_R1222_U499 & new_P1_R1222_U498;
  assign new_P1_R1222_U139 = new_P1_R1222_U347 & new_P1_R1222_U7;
  assign new_P1_R1222_U140 = ~new_P1_R1222_U119 | ~new_P1_R1222_U199;
  assign new_P1_R1222_U141 = ~new_P1_R1222_U214 | ~new_P1_R1222_U226;
  assign new_P1_R1222_U142 = ~new_P1_U3055;
  assign new_P1_R1222_U143 = ~new_P1_U4028;
  assign new_P1_R1222_U144 = new_P1_R1222_U400 & new_P1_R1222_U399;
  assign new_P1_R1222_U145 = ~new_P1_R1222_U361 | ~new_P1_R1222_U301 | ~new_P1_R1222_U166;
  assign new_P1_R1222_U146 = new_P1_R1222_U407 & new_P1_R1222_U406;
  assign new_P1_R1222_U147 = ~new_P1_R1222_U133 | ~new_P1_R1222_U367 | ~new_P1_R1222_U366;
  assign new_P1_R1222_U148 = new_P1_R1222_U414 & new_P1_R1222_U413;
  assign new_P1_R1222_U149 = ~new_P1_R1222_U87 | ~new_P1_R1222_U362 | ~new_P1_R1222_U296;
  assign new_P1_R1222_U150 = new_P1_R1222_U421 & new_P1_R1222_U420;
  assign new_P1_R1222_U151 = ~new_P1_R1222_U290 | ~new_P1_R1222_U289;
  assign new_P1_R1222_U152 = new_P1_R1222_U433 & new_P1_R1222_U432;
  assign new_P1_R1222_U153 = ~new_P1_R1222_U286 | ~new_P1_R1222_U285;
  assign new_P1_R1222_U154 = new_P1_R1222_U440 & new_P1_R1222_U439;
  assign new_P1_R1222_U155 = ~new_P1_R1222_U131 | ~new_P1_R1222_U281;
  assign new_P1_R1222_U156 = new_P1_R1222_U447 & new_P1_R1222_U446;
  assign new_P1_R1222_U157 = new_P1_R1222_U452 & new_P1_R1222_U451;
  assign new_P1_R1222_U158 = ~new_P1_R1222_U44 | ~new_P1_R1222_U324;
  assign new_P1_R1222_U159 = ~new_P1_R1222_U129 | ~new_P1_R1222_U266;
  assign new_P1_R1222_U160 = new_P1_R1222_U473 & new_P1_R1222_U472;
  assign new_P1_R1222_U161 = ~new_P1_R1222_U254 | ~new_P1_R1222_U253;
  assign new_P1_R1222_U162 = new_P1_R1222_U480 & new_P1_R1222_U479;
  assign new_P1_R1222_U163 = ~new_P1_R1222_U250 | ~new_P1_R1222_U249;
  assign new_P1_R1222_U164 = ~new_P1_R1222_U240 | ~new_P1_R1222_U239;
  assign new_P1_R1222_U165 = ~new_P1_R1222_U364 | ~new_P1_R1222_U363;
  assign new_P1_R1222_U166 = ~new_P1_U3054 | ~new_P1_R1222_U147;
  assign new_P1_R1222_U167 = ~new_P1_R1222_U35;
  assign new_P1_R1222_U168 = ~new_P1_U3485 | ~new_P1_U3083;
  assign new_P1_R1222_U169 = ~new_P1_U3072 | ~new_P1_U3494;
  assign new_P1_R1222_U170 = ~new_P1_U3058 | ~new_P1_U4020;
  assign new_P1_R1222_U171 = ~new_P1_R1222_U69;
  assign new_P1_R1222_U172 = ~new_P1_R1222_U78;
  assign new_P1_R1222_U173 = ~new_P1_U3065 | ~new_P1_U4021;
  assign new_P1_R1222_U174 = ~new_P1_R1222_U62;
  assign new_P1_R1222_U175 = new_P1_U3067 | new_P1_U3473;
  assign new_P1_R1222_U176 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1222_U177 = new_P1_U3467 | new_P1_U3064;
  assign new_P1_R1222_U178 = new_P1_U3464 | new_P1_U3068;
  assign new_P1_R1222_U179 = ~new_P1_R1222_U32;
  assign new_P1_R1222_U180 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1222_U181 = ~new_P1_R1222_U43;
  assign new_P1_R1222_U182 = ~new_P1_R1222_U44;
  assign new_P1_R1222_U183 = ~new_P1_R1222_U43 | ~new_P1_R1222_U44;
  assign new_P1_R1222_U184 = ~new_P1_R1222_U116 | ~new_P1_R1222_U177;
  assign new_P1_R1222_U185 = ~new_P1_R1222_U5 | ~new_P1_R1222_U183;
  assign new_P1_R1222_U186 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1222_U187 = ~new_P1_R1222_U117 | ~new_P1_R1222_U185;
  assign new_P1_R1222_U188 = ~new_P1_R1222_U36 | ~new_P1_R1222_U35;
  assign new_P1_R1222_U189 = ~new_P1_U3067 | ~new_P1_R1222_U188;
  assign new_P1_R1222_U190 = ~new_P1_R1222_U4 | ~new_P1_R1222_U187;
  assign new_P1_R1222_U191 = ~new_P1_U3473 | ~new_P1_R1222_U167;
  assign new_P1_R1222_U192 = ~new_P1_R1222_U42;
  assign new_P1_R1222_U193 = new_P1_U3070 | new_P1_U3479;
  assign new_P1_R1222_U194 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1222_U195 = ~new_P1_R1222_U23;
  assign new_P1_R1222_U196 = ~new_P1_R1222_U24 | ~new_P1_R1222_U23;
  assign new_P1_R1222_U197 = ~new_P1_U3070 | ~new_P1_R1222_U196;
  assign new_P1_R1222_U198 = ~new_P1_U3479 | ~new_P1_R1222_U195;
  assign new_P1_R1222_U199 = ~new_P1_R1222_U6 | ~new_P1_R1222_U42;
  assign new_P1_R1222_U200 = ~new_P1_R1222_U140;
  assign new_P1_R1222_U201 = new_P1_U3482 | new_P1_U3084;
  assign new_P1_R1222_U202 = ~new_P1_R1222_U201 | ~new_P1_R1222_U140;
  assign new_P1_R1222_U203 = ~new_P1_R1222_U41;
  assign new_P1_R1222_U204 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1222_U205 = new_P1_U3476 | new_P1_U3071;
  assign new_P1_R1222_U206 = ~new_P1_R1222_U205 | ~new_P1_R1222_U42;
  assign new_P1_R1222_U207 = ~new_P1_R1222_U120 | ~new_P1_R1222_U206;
  assign new_P1_R1222_U208 = ~new_P1_R1222_U192 | ~new_P1_R1222_U23;
  assign new_P1_R1222_U209 = ~new_P1_U3479 | ~new_P1_U3070;
  assign new_P1_R1222_U210 = ~new_P1_R1222_U121 | ~new_P1_R1222_U208;
  assign new_P1_R1222_U211 = new_P1_U3071 | new_P1_U3476;
  assign new_P1_R1222_U212 = ~new_P1_R1222_U182 | ~new_P1_R1222_U178;
  assign new_P1_R1222_U213 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1222_U214 = ~new_P1_R1222_U46;
  assign new_P1_R1222_U215 = ~new_P1_R1222_U181 | ~new_P1_R1222_U5;
  assign new_P1_R1222_U216 = ~new_P1_R1222_U46 | ~new_P1_R1222_U177;
  assign new_P1_R1222_U217 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1222_U218 = ~new_P1_R1222_U45;
  assign new_P1_R1222_U219 = new_P1_U3470 | new_P1_U3060;
  assign new_P1_R1222_U220 = ~new_P1_R1222_U219 | ~new_P1_R1222_U45;
  assign new_P1_R1222_U221 = ~new_P1_R1222_U123 | ~new_P1_R1222_U220;
  assign new_P1_R1222_U222 = ~new_P1_R1222_U218 | ~new_P1_R1222_U35;
  assign new_P1_R1222_U223 = ~new_P1_U3473 | ~new_P1_U3067;
  assign new_P1_R1222_U224 = ~new_P1_R1222_U124 | ~new_P1_R1222_U222;
  assign new_P1_R1222_U225 = new_P1_U3060 | new_P1_U3470;
  assign new_P1_R1222_U226 = ~new_P1_R1222_U181 | ~new_P1_R1222_U178;
  assign new_P1_R1222_U227 = ~new_P1_R1222_U141;
  assign new_P1_R1222_U228 = ~new_P1_U3064 | ~new_P1_U3467;
  assign new_P1_R1222_U229 = ~new_P1_R1222_U43 | ~new_P1_R1222_U44 | ~new_P1_R1222_U398 | ~new_P1_R1222_U397;
  assign new_P1_R1222_U230 = ~new_P1_R1222_U44 | ~new_P1_R1222_U43;
  assign new_P1_R1222_U231 = ~new_P1_U3068 | ~new_P1_U3464;
  assign new_P1_R1222_U232 = ~new_P1_R1222_U125 | ~new_P1_R1222_U230;
  assign new_P1_R1222_U233 = new_P1_U3083 | new_P1_U3485;
  assign new_P1_R1222_U234 = new_P1_U3062 | new_P1_U3488;
  assign new_P1_R1222_U235 = ~new_P1_R1222_U174 | ~new_P1_R1222_U7;
  assign new_P1_R1222_U236 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1222_U237 = ~new_P1_R1222_U127 | ~new_P1_R1222_U235;
  assign new_P1_R1222_U238 = new_P1_U3488 | new_P1_U3062;
  assign new_P1_R1222_U239 = ~new_P1_R1222_U126 | ~new_P1_R1222_U140;
  assign new_P1_R1222_U240 = ~new_P1_R1222_U238 | ~new_P1_R1222_U237;
  assign new_P1_R1222_U241 = ~new_P1_R1222_U164;
  assign new_P1_R1222_U242 = new_P1_U3080 | new_P1_U3497;
  assign new_P1_R1222_U243 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1222_U244 = ~new_P1_R1222_U171 | ~new_P1_R1222_U8;
  assign new_P1_R1222_U245 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1222_U246 = ~new_P1_R1222_U128 | ~new_P1_R1222_U244;
  assign new_P1_R1222_U247 = new_P1_U3491 | new_P1_U3063;
  assign new_P1_R1222_U248 = new_P1_U3497 | new_P1_U3080;
  assign new_P1_R1222_U249 = ~new_P1_R1222_U8 | ~new_P1_R1222_U247 | ~new_P1_R1222_U164;
  assign new_P1_R1222_U250 = ~new_P1_R1222_U248 | ~new_P1_R1222_U246;
  assign new_P1_R1222_U251 = ~new_P1_R1222_U163;
  assign new_P1_R1222_U252 = new_P1_U3500 | new_P1_U3079;
  assign new_P1_R1222_U253 = ~new_P1_R1222_U252 | ~new_P1_R1222_U163;
  assign new_P1_R1222_U254 = ~new_P1_U3079 | ~new_P1_U3500;
  assign new_P1_R1222_U255 = ~new_P1_R1222_U161;
  assign new_P1_R1222_U256 = new_P1_U3503 | new_P1_U3074;
  assign new_P1_R1222_U257 = ~new_P1_R1222_U256 | ~new_P1_R1222_U161;
  assign new_P1_R1222_U258 = ~new_P1_U3074 | ~new_P1_U3503;
  assign new_P1_R1222_U259 = ~new_P1_R1222_U93;
  assign new_P1_R1222_U260 = new_P1_U3069 | new_P1_U3509;
  assign new_P1_R1222_U261 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1222_U262 = ~new_P1_R1222_U60;
  assign new_P1_R1222_U263 = ~new_P1_R1222_U61 | ~new_P1_R1222_U60;
  assign new_P1_R1222_U264 = ~new_P1_U3069 | ~new_P1_R1222_U263;
  assign new_P1_R1222_U265 = ~new_P1_U3509 | ~new_P1_R1222_U262;
  assign new_P1_R1222_U266 = ~new_P1_R1222_U9 | ~new_P1_R1222_U93;
  assign new_P1_R1222_U267 = ~new_P1_R1222_U159;
  assign new_P1_R1222_U268 = new_P1_U3076 | new_P1_U4025;
  assign new_P1_R1222_U269 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1222_U270 = new_P1_U3075 | new_P1_U4024;
  assign new_P1_R1222_U271 = ~new_P1_R1222_U81;
  assign new_P1_R1222_U272 = ~new_P1_U4025 | ~new_P1_R1222_U271;
  assign new_P1_R1222_U273 = ~new_P1_R1222_U272 | ~new_P1_R1222_U91;
  assign new_P1_R1222_U274 = ~new_P1_R1222_U81 | ~new_P1_R1222_U82;
  assign new_P1_R1222_U275 = ~new_P1_R1222_U274 | ~new_P1_R1222_U273;
  assign new_P1_R1222_U276 = ~new_P1_R1222_U172 | ~new_P1_R1222_U10;
  assign new_P1_R1222_U277 = ~new_P1_U3075 | ~new_P1_U4024;
  assign new_P1_R1222_U278 = ~new_P1_R1222_U275 | ~new_P1_R1222_U276;
  assign new_P1_R1222_U279 = new_P1_U3512 | new_P1_U3082;
  assign new_P1_R1222_U280 = new_P1_U4024 | new_P1_U3075;
  assign new_P1_R1222_U281 = ~new_P1_R1222_U130 | ~new_P1_R1222_U270 | ~new_P1_R1222_U159;
  assign new_P1_R1222_U282 = ~new_P1_R1222_U280 | ~new_P1_R1222_U278;
  assign new_P1_R1222_U283 = ~new_P1_R1222_U155;
  assign new_P1_R1222_U284 = new_P1_U4023 | new_P1_U3061;
  assign new_P1_R1222_U285 = ~new_P1_R1222_U284 | ~new_P1_R1222_U155;
  assign new_P1_R1222_U286 = ~new_P1_U3061 | ~new_P1_U4023;
  assign new_P1_R1222_U287 = ~new_P1_R1222_U153;
  assign new_P1_R1222_U288 = new_P1_U4022 | new_P1_U3066;
  assign new_P1_R1222_U289 = ~new_P1_R1222_U288 | ~new_P1_R1222_U153;
  assign new_P1_R1222_U290 = ~new_P1_U3066 | ~new_P1_U4022;
  assign new_P1_R1222_U291 = ~new_P1_R1222_U151;
  assign new_P1_R1222_U292 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1222_U293 = ~new_P1_R1222_U173 | ~new_P1_R1222_U170;
  assign new_P1_R1222_U294 = ~new_P1_R1222_U87;
  assign new_P1_R1222_U295 = new_P1_U4021 | new_P1_U3065;
  assign new_P1_R1222_U296 = ~new_P1_R1222_U165 | ~new_P1_R1222_U151 | ~new_P1_R1222_U295;
  assign new_P1_R1222_U297 = ~new_P1_R1222_U149;
  assign new_P1_R1222_U298 = new_P1_U4018 | new_P1_U3053;
  assign new_P1_R1222_U299 = ~new_P1_U3053 | ~new_P1_U4018;
  assign new_P1_R1222_U300 = ~new_P1_R1222_U147;
  assign new_P1_R1222_U301 = ~new_P1_U4017 | ~new_P1_R1222_U147;
  assign new_P1_R1222_U302 = ~new_P1_R1222_U145;
  assign new_P1_R1222_U303 = ~new_P1_R1222_U295 | ~new_P1_R1222_U151;
  assign new_P1_R1222_U304 = ~new_P1_R1222_U90;
  assign new_P1_R1222_U305 = new_P1_U4020 | new_P1_U3058;
  assign new_P1_R1222_U306 = ~new_P1_R1222_U305 | ~new_P1_R1222_U90;
  assign new_P1_R1222_U307 = ~new_P1_R1222_U150 | ~new_P1_R1222_U306 | ~new_P1_R1222_U170;
  assign new_P1_R1222_U308 = ~new_P1_R1222_U304 | ~new_P1_R1222_U170;
  assign new_P1_R1222_U309 = ~new_P1_U4019 | ~new_P1_U3057;
  assign new_P1_R1222_U310 = ~new_P1_R1222_U165 | ~new_P1_R1222_U308 | ~new_P1_R1222_U309;
  assign new_P1_R1222_U311 = new_P1_U3058 | new_P1_U4020;
  assign new_P1_R1222_U312 = ~new_P1_R1222_U279 | ~new_P1_R1222_U159;
  assign new_P1_R1222_U313 = ~new_P1_R1222_U92;
  assign new_P1_R1222_U314 = ~new_P1_R1222_U10 | ~new_P1_R1222_U92;
  assign new_P1_R1222_U315 = ~new_P1_R1222_U134 | ~new_P1_R1222_U314;
  assign new_P1_R1222_U316 = ~new_P1_R1222_U314 | ~new_P1_R1222_U275;
  assign new_P1_R1222_U317 = ~new_P1_R1222_U450 | ~new_P1_R1222_U316;
  assign new_P1_R1222_U318 = new_P1_U3514 | new_P1_U3081;
  assign new_P1_R1222_U319 = ~new_P1_R1222_U318 | ~new_P1_R1222_U92;
  assign new_P1_R1222_U320 = ~new_P1_R1222_U157 | ~new_P1_R1222_U319 | ~new_P1_R1222_U81;
  assign new_P1_R1222_U321 = ~new_P1_R1222_U313 | ~new_P1_R1222_U81;
  assign new_P1_R1222_U322 = ~new_P1_U3076 | ~new_P1_U4025;
  assign new_P1_R1222_U323 = ~new_P1_R1222_U10 | ~new_P1_R1222_U322 | ~new_P1_R1222_U321;
  assign new_P1_R1222_U324 = new_P1_U3461 | new_P1_U3078;
  assign new_P1_R1222_U325 = ~new_P1_R1222_U158;
  assign new_P1_R1222_U326 = new_P1_U3081 | new_P1_U3514;
  assign new_P1_R1222_U327 = new_P1_U3506 | new_P1_U3073;
  assign new_P1_R1222_U328 = ~new_P1_R1222_U327 | ~new_P1_R1222_U93;
  assign new_P1_R1222_U329 = ~new_P1_R1222_U135 | ~new_P1_R1222_U328;
  assign new_P1_R1222_U330 = ~new_P1_R1222_U259 | ~new_P1_R1222_U60;
  assign new_P1_R1222_U331 = ~new_P1_U3509 | ~new_P1_U3069;
  assign new_P1_R1222_U332 = ~new_P1_R1222_U9 | ~new_P1_R1222_U331 | ~new_P1_R1222_U330;
  assign new_P1_R1222_U333 = new_P1_U3073 | new_P1_U3506;
  assign new_P1_R1222_U334 = ~new_P1_R1222_U247 | ~new_P1_R1222_U164;
  assign new_P1_R1222_U335 = ~new_P1_R1222_U94;
  assign new_P1_R1222_U336 = new_P1_U3494 | new_P1_U3072;
  assign new_P1_R1222_U337 = ~new_P1_R1222_U336 | ~new_P1_R1222_U94;
  assign new_P1_R1222_U338 = ~new_P1_R1222_U136 | ~new_P1_R1222_U337;
  assign new_P1_R1222_U339 = ~new_P1_R1222_U335 | ~new_P1_R1222_U169;
  assign new_P1_R1222_U340 = ~new_P1_U3080 | ~new_P1_U3497;
  assign new_P1_R1222_U341 = ~new_P1_R1222_U137 | ~new_P1_R1222_U339;
  assign new_P1_R1222_U342 = new_P1_U3072 | new_P1_U3494;
  assign new_P1_R1222_U343 = new_P1_U3485 | new_P1_U3083;
  assign new_P1_R1222_U344 = ~new_P1_R1222_U343 | ~new_P1_R1222_U41;
  assign new_P1_R1222_U345 = ~new_P1_R1222_U138 | ~new_P1_R1222_U344;
  assign new_P1_R1222_U346 = ~new_P1_R1222_U203 | ~new_P1_R1222_U168;
  assign new_P1_R1222_U347 = ~new_P1_U3062 | ~new_P1_U3488;
  assign new_P1_R1222_U348 = ~new_P1_R1222_U139 | ~new_P1_R1222_U346;
  assign new_P1_R1222_U349 = ~new_P1_R1222_U204 | ~new_P1_R1222_U168;
  assign new_P1_R1222_U350 = ~new_P1_R1222_U201 | ~new_P1_R1222_U62;
  assign new_P1_R1222_U351 = ~new_P1_R1222_U211 | ~new_P1_R1222_U23;
  assign new_P1_R1222_U352 = ~new_P1_R1222_U225 | ~new_P1_R1222_U35;
  assign new_P1_R1222_U353 = ~new_P1_R1222_U228 | ~new_P1_R1222_U177;
  assign new_P1_R1222_U354 = ~new_P1_R1222_U311 | ~new_P1_R1222_U170;
  assign new_P1_R1222_U355 = ~new_P1_R1222_U295 | ~new_P1_R1222_U173;
  assign new_P1_R1222_U356 = ~new_P1_R1222_U326 | ~new_P1_R1222_U81;
  assign new_P1_R1222_U357 = ~new_P1_R1222_U279 | ~new_P1_R1222_U78;
  assign new_P1_R1222_U358 = ~new_P1_R1222_U333 | ~new_P1_R1222_U60;
  assign new_P1_R1222_U359 = ~new_P1_R1222_U342 | ~new_P1_R1222_U169;
  assign new_P1_R1222_U360 = ~new_P1_R1222_U247 | ~new_P1_R1222_U69;
  assign new_P1_R1222_U361 = ~new_P1_U4017 | ~new_P1_U3054;
  assign new_P1_R1222_U362 = ~new_P1_R1222_U293 | ~new_P1_R1222_U165;
  assign new_P1_R1222_U363 = ~new_P1_U3057 | ~new_P1_R1222_U292;
  assign new_P1_R1222_U364 = ~new_P1_U4019 | ~new_P1_R1222_U292;
  assign new_P1_R1222_U365 = ~new_P1_R1222_U298 | ~new_P1_R1222_U293 | ~new_P1_R1222_U165;
  assign new_P1_R1222_U366 = ~new_P1_R1222_U132 | ~new_P1_R1222_U151 | ~new_P1_R1222_U165;
  assign new_P1_R1222_U367 = ~new_P1_R1222_U294 | ~new_P1_R1222_U298;
  assign new_P1_R1222_U368 = ~new_P1_U3083 | ~new_P1_R1222_U40;
  assign new_P1_R1222_U369 = ~new_P1_U3485 | ~new_P1_R1222_U39;
  assign new_P1_R1222_U370 = ~new_P1_R1222_U369 | ~new_P1_R1222_U368;
  assign new_P1_R1222_U371 = ~new_P1_R1222_U349 | ~new_P1_R1222_U41;
  assign new_P1_R1222_U372 = ~new_P1_R1222_U370 | ~new_P1_R1222_U203;
  assign new_P1_R1222_U373 = ~new_P1_U3084 | ~new_P1_R1222_U37;
  assign new_P1_R1222_U374 = ~new_P1_U3482 | ~new_P1_R1222_U38;
  assign new_P1_R1222_U375 = ~new_P1_R1222_U374 | ~new_P1_R1222_U373;
  assign new_P1_R1222_U376 = ~new_P1_R1222_U350 | ~new_P1_R1222_U140;
  assign new_P1_R1222_U377 = ~new_P1_R1222_U200 | ~new_P1_R1222_U375;
  assign new_P1_R1222_U378 = ~new_P1_U3070 | ~new_P1_R1222_U24;
  assign new_P1_R1222_U379 = ~new_P1_U3479 | ~new_P1_R1222_U22;
  assign new_P1_R1222_U380 = ~new_P1_U3071 | ~new_P1_R1222_U20;
  assign new_P1_R1222_U381 = ~new_P1_U3476 | ~new_P1_R1222_U21;
  assign new_P1_R1222_U382 = ~new_P1_R1222_U381 | ~new_P1_R1222_U380;
  assign new_P1_R1222_U383 = ~new_P1_R1222_U351 | ~new_P1_R1222_U42;
  assign new_P1_R1222_U384 = ~new_P1_R1222_U382 | ~new_P1_R1222_U192;
  assign new_P1_R1222_U385 = ~new_P1_U3067 | ~new_P1_R1222_U36;
  assign new_P1_R1222_U386 = ~new_P1_U3473 | ~new_P1_R1222_U27;
  assign new_P1_R1222_U387 = ~new_P1_U3060 | ~new_P1_R1222_U25;
  assign new_P1_R1222_U388 = ~new_P1_U3470 | ~new_P1_R1222_U26;
  assign new_P1_R1222_U389 = ~new_P1_R1222_U388 | ~new_P1_R1222_U387;
  assign new_P1_R1222_U390 = ~new_P1_R1222_U352 | ~new_P1_R1222_U45;
  assign new_P1_R1222_U391 = ~new_P1_R1222_U389 | ~new_P1_R1222_U218;
  assign new_P1_R1222_U392 = ~new_P1_U3064 | ~new_P1_R1222_U33;
  assign new_P1_R1222_U393 = ~new_P1_U3467 | ~new_P1_R1222_U34;
  assign new_P1_R1222_U394 = ~new_P1_R1222_U393 | ~new_P1_R1222_U392;
  assign new_P1_R1222_U395 = ~new_P1_R1222_U353 | ~new_P1_R1222_U141;
  assign new_P1_R1222_U396 = ~new_P1_R1222_U227 | ~new_P1_R1222_U394;
  assign new_P1_R1222_U397 = ~new_P1_U3068 | ~new_P1_R1222_U28;
  assign new_P1_R1222_U398 = ~new_P1_U3464 | ~new_P1_R1222_U29;
  assign new_P1_R1222_U399 = ~new_P1_U3055 | ~new_P1_R1222_U143;
  assign new_P1_R1222_U400 = ~new_P1_U4028 | ~new_P1_R1222_U142;
  assign new_P1_R1222_U401 = ~new_P1_U3055 | ~new_P1_R1222_U143;
  assign new_P1_R1222_U402 = ~new_P1_U4028 | ~new_P1_R1222_U142;
  assign new_P1_R1222_U403 = ~new_P1_R1222_U402 | ~new_P1_R1222_U401;
  assign new_P1_R1222_U404 = ~new_P1_R1222_U144 | ~new_P1_R1222_U145;
  assign new_P1_R1222_U405 = ~new_P1_R1222_U302 | ~new_P1_R1222_U403;
  assign new_P1_R1222_U406 = ~new_P1_U3054 | ~new_P1_R1222_U89;
  assign new_P1_R1222_U407 = ~new_P1_U4017 | ~new_P1_R1222_U88;
  assign new_P1_R1222_U408 = ~new_P1_U3054 | ~new_P1_R1222_U89;
  assign new_P1_R1222_U409 = ~new_P1_U4017 | ~new_P1_R1222_U88;
  assign new_P1_R1222_U410 = ~new_P1_R1222_U409 | ~new_P1_R1222_U408;
  assign new_P1_R1222_U411 = ~new_P1_R1222_U146 | ~new_P1_R1222_U147;
  assign new_P1_R1222_U412 = ~new_P1_R1222_U300 | ~new_P1_R1222_U410;
  assign new_P1_R1222_U413 = ~new_P1_U3053 | ~new_P1_R1222_U47;
  assign new_P1_R1222_U414 = ~new_P1_U4018 | ~new_P1_R1222_U48;
  assign new_P1_R1222_U415 = ~new_P1_U3053 | ~new_P1_R1222_U47;
  assign new_P1_R1222_U416 = ~new_P1_U4018 | ~new_P1_R1222_U48;
  assign new_P1_R1222_U417 = ~new_P1_R1222_U416 | ~new_P1_R1222_U415;
  assign new_P1_R1222_U418 = ~new_P1_R1222_U148 | ~new_P1_R1222_U149;
  assign new_P1_R1222_U419 = ~new_P1_R1222_U297 | ~new_P1_R1222_U417;
  assign new_P1_R1222_U420 = ~new_P1_U3057 | ~new_P1_R1222_U50;
  assign new_P1_R1222_U421 = ~new_P1_U4019 | ~new_P1_R1222_U49;
  assign new_P1_R1222_U422 = ~new_P1_U3058 | ~new_P1_R1222_U51;
  assign new_P1_R1222_U423 = ~new_P1_U4020 | ~new_P1_R1222_U52;
  assign new_P1_R1222_U424 = ~new_P1_R1222_U423 | ~new_P1_R1222_U422;
  assign new_P1_R1222_U425 = ~new_P1_R1222_U354 | ~new_P1_R1222_U90;
  assign new_P1_R1222_U426 = ~new_P1_R1222_U424 | ~new_P1_R1222_U304;
  assign new_P1_R1222_U427 = ~new_P1_U3065 | ~new_P1_R1222_U53;
  assign new_P1_R1222_U428 = ~new_P1_U4021 | ~new_P1_R1222_U54;
  assign new_P1_R1222_U429 = ~new_P1_R1222_U428 | ~new_P1_R1222_U427;
  assign new_P1_R1222_U430 = ~new_P1_R1222_U355 | ~new_P1_R1222_U151;
  assign new_P1_R1222_U431 = ~new_P1_R1222_U291 | ~new_P1_R1222_U429;
  assign new_P1_R1222_U432 = ~new_P1_U3066 | ~new_P1_R1222_U85;
  assign new_P1_R1222_U433 = ~new_P1_U4022 | ~new_P1_R1222_U86;
  assign new_P1_R1222_U434 = ~new_P1_U3066 | ~new_P1_R1222_U85;
  assign new_P1_R1222_U435 = ~new_P1_U4022 | ~new_P1_R1222_U86;
  assign new_P1_R1222_U436 = ~new_P1_R1222_U435 | ~new_P1_R1222_U434;
  assign new_P1_R1222_U437 = ~new_P1_R1222_U152 | ~new_P1_R1222_U153;
  assign new_P1_R1222_U438 = ~new_P1_R1222_U287 | ~new_P1_R1222_U436;
  assign new_P1_R1222_U439 = ~new_P1_U3061 | ~new_P1_R1222_U83;
  assign new_P1_R1222_U440 = ~new_P1_U4023 | ~new_P1_R1222_U84;
  assign new_P1_R1222_U441 = ~new_P1_U3061 | ~new_P1_R1222_U83;
  assign new_P1_R1222_U442 = ~new_P1_U4023 | ~new_P1_R1222_U84;
  assign new_P1_R1222_U443 = ~new_P1_R1222_U442 | ~new_P1_R1222_U441;
  assign new_P1_R1222_U444 = ~new_P1_R1222_U154 | ~new_P1_R1222_U155;
  assign new_P1_R1222_U445 = ~new_P1_R1222_U283 | ~new_P1_R1222_U443;
  assign new_P1_R1222_U446 = ~new_P1_U3075 | ~new_P1_R1222_U55;
  assign new_P1_R1222_U447 = ~new_P1_U4024 | ~new_P1_R1222_U56;
  assign new_P1_R1222_U448 = ~new_P1_U3075 | ~new_P1_R1222_U55;
  assign new_P1_R1222_U449 = ~new_P1_U4024 | ~new_P1_R1222_U56;
  assign new_P1_R1222_U450 = ~new_P1_R1222_U449 | ~new_P1_R1222_U448;
  assign new_P1_R1222_U451 = ~new_P1_U3076 | ~new_P1_R1222_U82;
  assign new_P1_R1222_U452 = ~new_P1_U4025 | ~new_P1_R1222_U91;
  assign new_P1_R1222_U453 = ~new_P1_R1222_U179 | ~new_P1_R1222_U158;
  assign new_P1_R1222_U454 = ~new_P1_R1222_U325 | ~new_P1_R1222_U32;
  assign new_P1_R1222_U455 = ~new_P1_U3081 | ~new_P1_R1222_U79;
  assign new_P1_R1222_U456 = ~new_P1_U3514 | ~new_P1_R1222_U80;
  assign new_P1_R1222_U457 = ~new_P1_R1222_U456 | ~new_P1_R1222_U455;
  assign new_P1_R1222_U458 = ~new_P1_R1222_U356 | ~new_P1_R1222_U92;
  assign new_P1_R1222_U459 = ~new_P1_R1222_U457 | ~new_P1_R1222_U313;
  assign new_P1_R1222_U460 = ~new_P1_U3082 | ~new_P1_R1222_U76;
  assign new_P1_R1222_U461 = ~new_P1_U3512 | ~new_P1_R1222_U77;
  assign new_P1_R1222_U462 = ~new_P1_R1222_U461 | ~new_P1_R1222_U460;
  assign new_P1_R1222_U463 = ~new_P1_R1222_U357 | ~new_P1_R1222_U159;
  assign new_P1_R1222_U464 = ~new_P1_R1222_U267 | ~new_P1_R1222_U462;
  assign new_P1_R1222_U465 = ~new_P1_U3069 | ~new_P1_R1222_U61;
  assign new_P1_R1222_U466 = ~new_P1_U3509 | ~new_P1_R1222_U59;
  assign new_P1_R1222_U467 = ~new_P1_U3073 | ~new_P1_R1222_U57;
  assign new_P1_R1222_U468 = ~new_P1_U3506 | ~new_P1_R1222_U58;
  assign new_P1_R1222_U469 = ~new_P1_R1222_U468 | ~new_P1_R1222_U467;
  assign new_P1_R1222_U470 = ~new_P1_R1222_U358 | ~new_P1_R1222_U93;
  assign new_P1_R1222_U471 = ~new_P1_R1222_U469 | ~new_P1_R1222_U259;
  assign new_P1_R1222_U472 = ~new_P1_U3074 | ~new_P1_R1222_U74;
  assign new_P1_R1222_U473 = ~new_P1_U3503 | ~new_P1_R1222_U75;
  assign new_P1_R1222_U474 = ~new_P1_U3074 | ~new_P1_R1222_U74;
  assign new_P1_R1222_U475 = ~new_P1_U3503 | ~new_P1_R1222_U75;
  assign new_P1_R1222_U476 = ~new_P1_R1222_U475 | ~new_P1_R1222_U474;
  assign new_P1_R1222_U477 = ~new_P1_R1222_U160 | ~new_P1_R1222_U161;
  assign new_P1_R1222_U478 = ~new_P1_R1222_U255 | ~new_P1_R1222_U476;
  assign new_P1_R1222_U479 = ~new_P1_U3079 | ~new_P1_R1222_U72;
  assign new_P1_R1222_U480 = ~new_P1_U3500 | ~new_P1_R1222_U73;
  assign new_P1_R1222_U481 = ~new_P1_U3079 | ~new_P1_R1222_U72;
  assign new_P1_R1222_U482 = ~new_P1_U3500 | ~new_P1_R1222_U73;
  assign new_P1_R1222_U483 = ~new_P1_R1222_U482 | ~new_P1_R1222_U481;
  assign new_P1_R1222_U484 = ~new_P1_R1222_U162 | ~new_P1_R1222_U163;
  assign new_P1_R1222_U485 = ~new_P1_R1222_U251 | ~new_P1_R1222_U483;
  assign new_P1_R1222_U486 = ~new_P1_U3080 | ~new_P1_R1222_U70;
  assign new_P1_R1222_U487 = ~new_P1_U3497 | ~new_P1_R1222_U71;
  assign new_P1_R1222_U488 = ~new_P1_U3072 | ~new_P1_R1222_U65;
  assign new_P1_R1222_U489 = ~new_P1_U3494 | ~new_P1_R1222_U66;
  assign new_P1_R1222_U490 = ~new_P1_R1222_U489 | ~new_P1_R1222_U488;
  assign new_P1_R1222_U491 = ~new_P1_R1222_U359 | ~new_P1_R1222_U94;
  assign new_P1_R1222_U492 = ~new_P1_R1222_U490 | ~new_P1_R1222_U335;
  assign new_P1_R1222_U493 = ~new_P1_U3063 | ~new_P1_R1222_U67;
  assign new_P1_R1222_U494 = ~new_P1_U3491 | ~new_P1_R1222_U68;
  assign new_P1_R1222_U495 = ~new_P1_R1222_U494 | ~new_P1_R1222_U493;
  assign new_P1_R1222_U496 = ~new_P1_R1222_U360 | ~new_P1_R1222_U164;
  assign new_P1_R1222_U497 = ~new_P1_R1222_U241 | ~new_P1_R1222_U495;
  assign new_P1_R1222_U498 = ~new_P1_U3062 | ~new_P1_R1222_U63;
  assign new_P1_R1222_U499 = ~new_P1_U3488 | ~new_P1_R1222_U64;
  assign new_P1_R1222_U500 = ~new_P1_U3077 | ~new_P1_R1222_U30;
  assign new_P1_R1222_U501 = ~new_P1_U3456 | ~new_P1_R1222_U31;
  assign new_P2_ADD_1119_U4 = ~P2_REG3_REG_3_;
  assign new_P2_ADD_1119_U5 = new_P2_ADD_1119_U78 & new_P2_ADD_1119_U106;
  assign new_P2_ADD_1119_U6 = ~P2_REG3_REG_5_;
  assign new_P2_ADD_1119_U7 = ~P2_REG3_REG_4_;
  assign new_P2_ADD_1119_U8 = ~P2_REG3_REG_4_ | ~P2_REG3_REG_5_ | ~P2_REG3_REG_3_;
  assign new_P2_ADD_1119_U9 = ~P2_REG3_REG_7_;
  assign new_P2_ADD_1119_U10 = ~P2_REG3_REG_6_;
  assign new_P2_ADD_1119_U11 = ~new_P2_ADD_1119_U75 | ~new_P2_ADD_1119_U85;
  assign new_P2_ADD_1119_U12 = ~P2_REG3_REG_8_;
  assign new_P2_ADD_1119_U13 = ~P2_REG3_REG_9_;
  assign new_P2_ADD_1119_U14 = ~new_P2_ADD_1119_U76 | ~new_P2_ADD_1119_U87;
  assign new_P2_ADD_1119_U15 = ~P2_REG3_REG_11_;
  assign new_P2_ADD_1119_U16 = ~P2_REG3_REG_10_;
  assign new_P2_ADD_1119_U17 = ~new_P2_ADD_1119_U77 | ~new_P2_ADD_1119_U89;
  assign new_P2_ADD_1119_U18 = ~P2_REG3_REG_12_;
  assign new_P2_ADD_1119_U19 = ~P2_REG3_REG_12_ | ~new_P2_ADD_1119_U91;
  assign new_P2_ADD_1119_U20 = ~P2_REG3_REG_13_;
  assign new_P2_ADD_1119_U21 = ~P2_REG3_REG_13_ | ~new_P2_ADD_1119_U92;
  assign new_P2_ADD_1119_U22 = ~P2_REG3_REG_14_;
  assign new_P2_ADD_1119_U23 = ~P2_REG3_REG_14_ | ~new_P2_ADD_1119_U93;
  assign new_P2_ADD_1119_U24 = ~P2_REG3_REG_15_;
  assign new_P2_ADD_1119_U25 = ~P2_REG3_REG_15_ | ~new_P2_ADD_1119_U94;
  assign new_P2_ADD_1119_U26 = ~P2_REG3_REG_16_;
  assign new_P2_ADD_1119_U27 = ~P2_REG3_REG_16_ | ~new_P2_ADD_1119_U95;
  assign new_P2_ADD_1119_U28 = ~P2_REG3_REG_17_;
  assign new_P2_ADD_1119_U29 = ~P2_REG3_REG_17_ | ~new_P2_ADD_1119_U96;
  assign new_P2_ADD_1119_U30 = ~P2_REG3_REG_18_;
  assign new_P2_ADD_1119_U31 = ~P2_REG3_REG_18_ | ~new_P2_ADD_1119_U97;
  assign new_P2_ADD_1119_U32 = ~P2_REG3_REG_19_;
  assign new_P2_ADD_1119_U33 = ~P2_REG3_REG_19_ | ~new_P2_ADD_1119_U98;
  assign new_P2_ADD_1119_U34 = ~P2_REG3_REG_20_;
  assign new_P2_ADD_1119_U35 = ~P2_REG3_REG_20_ | ~new_P2_ADD_1119_U99;
  assign new_P2_ADD_1119_U36 = ~P2_REG3_REG_21_;
  assign new_P2_ADD_1119_U37 = ~P2_REG3_REG_21_ | ~new_P2_ADD_1119_U100;
  assign new_P2_ADD_1119_U38 = ~P2_REG3_REG_22_;
  assign new_P2_ADD_1119_U39 = ~P2_REG3_REG_22_ | ~new_P2_ADD_1119_U101;
  assign new_P2_ADD_1119_U40 = ~P2_REG3_REG_23_;
  assign new_P2_ADD_1119_U41 = ~P2_REG3_REG_23_ | ~new_P2_ADD_1119_U102;
  assign new_P2_ADD_1119_U42 = ~P2_REG3_REG_24_;
  assign new_P2_ADD_1119_U43 = ~P2_REG3_REG_24_ | ~new_P2_ADD_1119_U103;
  assign new_P2_ADD_1119_U44 = ~P2_REG3_REG_25_;
  assign new_P2_ADD_1119_U45 = ~P2_REG3_REG_25_ | ~new_P2_ADD_1119_U104;
  assign new_P2_ADD_1119_U46 = ~P2_REG3_REG_26_;
  assign new_P2_ADD_1119_U47 = ~P2_REG3_REG_26_ | ~new_P2_ADD_1119_U105;
  assign new_P2_ADD_1119_U48 = ~P2_REG3_REG_28_;
  assign new_P2_ADD_1119_U49 = ~P2_REG3_REG_27_;
  assign new_P2_ADD_1119_U50 = ~new_P2_ADD_1119_U109 | ~new_P2_ADD_1119_U108;
  assign new_P2_ADD_1119_U51 = ~new_P2_ADD_1119_U111 | ~new_P2_ADD_1119_U110;
  assign new_P2_ADD_1119_U52 = ~new_P2_ADD_1119_U113 | ~new_P2_ADD_1119_U112;
  assign new_P2_ADD_1119_U53 = ~new_P2_ADD_1119_U115 | ~new_P2_ADD_1119_U114;
  assign new_P2_ADD_1119_U54 = ~new_P2_ADD_1119_U117 | ~new_P2_ADD_1119_U116;
  assign new_P2_ADD_1119_U55 = ~new_P2_ADD_1119_U119 | ~new_P2_ADD_1119_U118;
  assign new_P2_ADD_1119_U56 = ~new_P2_ADD_1119_U121 | ~new_P2_ADD_1119_U120;
  assign new_P2_ADD_1119_U57 = ~new_P2_ADD_1119_U123 | ~new_P2_ADD_1119_U122;
  assign new_P2_ADD_1119_U58 = ~new_P2_ADD_1119_U125 | ~new_P2_ADD_1119_U124;
  assign new_P2_ADD_1119_U59 = ~new_P2_ADD_1119_U127 | ~new_P2_ADD_1119_U126;
  assign new_P2_ADD_1119_U60 = ~new_P2_ADD_1119_U129 | ~new_P2_ADD_1119_U128;
  assign new_P2_ADD_1119_U61 = ~new_P2_ADD_1119_U131 | ~new_P2_ADD_1119_U130;
  assign new_P2_ADD_1119_U62 = ~new_P2_ADD_1119_U133 | ~new_P2_ADD_1119_U132;
  assign new_P2_ADD_1119_U63 = ~new_P2_ADD_1119_U135 | ~new_P2_ADD_1119_U134;
  assign new_P2_ADD_1119_U64 = ~new_P2_ADD_1119_U137 | ~new_P2_ADD_1119_U136;
  assign new_P2_ADD_1119_U65 = ~new_P2_ADD_1119_U139 | ~new_P2_ADD_1119_U138;
  assign new_P2_ADD_1119_U66 = ~new_P2_ADD_1119_U141 | ~new_P2_ADD_1119_U140;
  assign new_P2_ADD_1119_U67 = ~new_P2_ADD_1119_U143 | ~new_P2_ADD_1119_U142;
  assign new_P2_ADD_1119_U68 = ~new_P2_ADD_1119_U145 | ~new_P2_ADD_1119_U144;
  assign new_P2_ADD_1119_U69 = ~new_P2_ADD_1119_U147 | ~new_P2_ADD_1119_U146;
  assign new_P2_ADD_1119_U70 = ~new_P2_ADD_1119_U149 | ~new_P2_ADD_1119_U148;
  assign new_P2_ADD_1119_U71 = ~new_P2_ADD_1119_U151 | ~new_P2_ADD_1119_U150;
  assign new_P2_ADD_1119_U72 = ~new_P2_ADD_1119_U153 | ~new_P2_ADD_1119_U152;
  assign new_P2_ADD_1119_U73 = ~new_P2_ADD_1119_U155 | ~new_P2_ADD_1119_U154;
  assign new_P2_ADD_1119_U74 = ~new_P2_ADD_1119_U157 | ~new_P2_ADD_1119_U156;
  assign new_P2_ADD_1119_U75 = P2_REG3_REG_7_ & P2_REG3_REG_6_;
  assign new_P2_ADD_1119_U76 = P2_REG3_REG_8_ & P2_REG3_REG_9_;
  assign new_P2_ADD_1119_U77 = P2_REG3_REG_11_ & P2_REG3_REG_10_;
  assign new_P2_ADD_1119_U78 = P2_REG3_REG_28_ & P2_REG3_REG_27_;
  assign new_P2_ADD_1119_U79 = ~P2_REG3_REG_8_ | ~new_P2_ADD_1119_U87;
  assign new_P2_ADD_1119_U80 = ~P2_REG3_REG_6_ | ~new_P2_ADD_1119_U85;
  assign new_P2_ADD_1119_U81 = ~P2_REG3_REG_4_ | ~P2_REG3_REG_3_;
  assign new_P2_ADD_1119_U82 = ~P2_REG3_REG_27_ | ~new_P2_ADD_1119_U106;
  assign new_P2_ADD_1119_U83 = ~P2_REG3_REG_10_ | ~new_P2_ADD_1119_U89;
  assign new_P2_ADD_1119_U84 = ~new_P2_ADD_1119_U81;
  assign new_P2_ADD_1119_U85 = ~new_P2_ADD_1119_U8;
  assign new_P2_ADD_1119_U86 = ~new_P2_ADD_1119_U80;
  assign new_P2_ADD_1119_U87 = ~new_P2_ADD_1119_U11;
  assign new_P2_ADD_1119_U88 = ~new_P2_ADD_1119_U79;
  assign new_P2_ADD_1119_U89 = ~new_P2_ADD_1119_U14;
  assign new_P2_ADD_1119_U90 = ~new_P2_ADD_1119_U83;
  assign new_P2_ADD_1119_U91 = ~new_P2_ADD_1119_U17;
  assign new_P2_ADD_1119_U92 = ~new_P2_ADD_1119_U19;
  assign new_P2_ADD_1119_U93 = ~new_P2_ADD_1119_U21;
  assign new_P2_ADD_1119_U94 = ~new_P2_ADD_1119_U23;
  assign new_P2_ADD_1119_U95 = ~new_P2_ADD_1119_U25;
  assign new_P2_ADD_1119_U96 = ~new_P2_ADD_1119_U27;
  assign new_P2_ADD_1119_U97 = ~new_P2_ADD_1119_U29;
  assign new_P2_ADD_1119_U98 = ~new_P2_ADD_1119_U31;
  assign new_P2_ADD_1119_U99 = ~new_P2_ADD_1119_U33;
  assign new_P2_ADD_1119_U100 = ~new_P2_ADD_1119_U35;
  assign new_P2_ADD_1119_U101 = ~new_P2_ADD_1119_U37;
  assign new_P2_ADD_1119_U102 = ~new_P2_ADD_1119_U39;
  assign new_P2_ADD_1119_U103 = ~new_P2_ADD_1119_U41;
  assign new_P2_ADD_1119_U104 = ~new_P2_ADD_1119_U43;
  assign new_P2_ADD_1119_U105 = ~new_P2_ADD_1119_U45;
  assign new_P2_ADD_1119_U106 = ~new_P2_ADD_1119_U47;
  assign new_P2_ADD_1119_U107 = ~new_P2_ADD_1119_U82;
  assign new_P2_ADD_1119_U108 = ~P2_REG3_REG_9_ | ~new_P2_ADD_1119_U79;
  assign new_P2_ADD_1119_U109 = ~new_P2_ADD_1119_U88 | ~new_P2_ADD_1119_U13;
  assign new_P2_ADD_1119_U110 = ~P2_REG3_REG_8_ | ~new_P2_ADD_1119_U11;
  assign new_P2_ADD_1119_U111 = ~new_P2_ADD_1119_U87 | ~new_P2_ADD_1119_U12;
  assign new_P2_ADD_1119_U112 = ~P2_REG3_REG_7_ | ~new_P2_ADD_1119_U80;
  assign new_P2_ADD_1119_U113 = ~new_P2_ADD_1119_U86 | ~new_P2_ADD_1119_U9;
  assign new_P2_ADD_1119_U114 = ~P2_REG3_REG_6_ | ~new_P2_ADD_1119_U8;
  assign new_P2_ADD_1119_U115 = ~new_P2_ADD_1119_U85 | ~new_P2_ADD_1119_U10;
  assign new_P2_ADD_1119_U116 = ~P2_REG3_REG_5_ | ~new_P2_ADD_1119_U81;
  assign new_P2_ADD_1119_U117 = ~new_P2_ADD_1119_U84 | ~new_P2_ADD_1119_U6;
  assign new_P2_ADD_1119_U118 = ~P2_REG3_REG_4_ | ~new_P2_ADD_1119_U4;
  assign new_P2_ADD_1119_U119 = ~P2_REG3_REG_3_ | ~new_P2_ADD_1119_U7;
  assign new_P2_ADD_1119_U120 = ~P2_REG3_REG_28_ | ~new_P2_ADD_1119_U82;
  assign new_P2_ADD_1119_U121 = ~new_P2_ADD_1119_U107 | ~new_P2_ADD_1119_U48;
  assign new_P2_ADD_1119_U122 = ~P2_REG3_REG_27_ | ~new_P2_ADD_1119_U47;
  assign new_P2_ADD_1119_U123 = ~new_P2_ADD_1119_U106 | ~new_P2_ADD_1119_U49;
  assign new_P2_ADD_1119_U124 = ~P2_REG3_REG_26_ | ~new_P2_ADD_1119_U45;
  assign new_P2_ADD_1119_U125 = ~new_P2_ADD_1119_U105 | ~new_P2_ADD_1119_U46;
  assign new_P2_ADD_1119_U126 = ~P2_REG3_REG_25_ | ~new_P2_ADD_1119_U43;
  assign new_P2_ADD_1119_U127 = ~new_P2_ADD_1119_U104 | ~new_P2_ADD_1119_U44;
  assign new_P2_ADD_1119_U128 = ~P2_REG3_REG_24_ | ~new_P2_ADD_1119_U41;
  assign new_P2_ADD_1119_U129 = ~new_P2_ADD_1119_U103 | ~new_P2_ADD_1119_U42;
  assign new_P2_ADD_1119_U130 = ~P2_REG3_REG_23_ | ~new_P2_ADD_1119_U39;
  assign new_P2_ADD_1119_U131 = ~new_P2_ADD_1119_U102 | ~new_P2_ADD_1119_U40;
  assign new_P2_ADD_1119_U132 = ~P2_REG3_REG_22_ | ~new_P2_ADD_1119_U37;
  assign new_P2_ADD_1119_U133 = ~new_P2_ADD_1119_U101 | ~new_P2_ADD_1119_U38;
  assign new_P2_ADD_1119_U134 = ~P2_REG3_REG_21_ | ~new_P2_ADD_1119_U35;
  assign new_P2_ADD_1119_U135 = ~new_P2_ADD_1119_U100 | ~new_P2_ADD_1119_U36;
  assign new_P2_ADD_1119_U136 = ~P2_REG3_REG_20_ | ~new_P2_ADD_1119_U33;
  assign new_P2_ADD_1119_U137 = ~new_P2_ADD_1119_U99 | ~new_P2_ADD_1119_U34;
  assign new_P2_ADD_1119_U138 = ~P2_REG3_REG_19_ | ~new_P2_ADD_1119_U31;
  assign new_P2_ADD_1119_U139 = ~new_P2_ADD_1119_U98 | ~new_P2_ADD_1119_U32;
  assign new_P2_ADD_1119_U140 = ~P2_REG3_REG_18_ | ~new_P2_ADD_1119_U29;
  assign new_P2_ADD_1119_U141 = ~new_P2_ADD_1119_U97 | ~new_P2_ADD_1119_U30;
  assign new_P2_ADD_1119_U142 = ~P2_REG3_REG_17_ | ~new_P2_ADD_1119_U27;
  assign new_P2_ADD_1119_U143 = ~new_P2_ADD_1119_U96 | ~new_P2_ADD_1119_U28;
  assign new_P2_ADD_1119_U144 = ~P2_REG3_REG_16_ | ~new_P2_ADD_1119_U25;
  assign new_P2_ADD_1119_U145 = ~new_P2_ADD_1119_U95 | ~new_P2_ADD_1119_U26;
  assign new_P2_ADD_1119_U146 = ~P2_REG3_REG_15_ | ~new_P2_ADD_1119_U23;
  assign new_P2_ADD_1119_U147 = ~new_P2_ADD_1119_U94 | ~new_P2_ADD_1119_U24;
  assign new_P2_ADD_1119_U148 = ~P2_REG3_REG_14_ | ~new_P2_ADD_1119_U21;
  assign new_P2_ADD_1119_U149 = ~new_P2_ADD_1119_U93 | ~new_P2_ADD_1119_U22;
  assign new_P2_ADD_1119_U150 = ~P2_REG3_REG_13_ | ~new_P2_ADD_1119_U19;
  assign new_P2_ADD_1119_U151 = ~new_P2_ADD_1119_U92 | ~new_P2_ADD_1119_U20;
  assign new_P2_ADD_1119_U152 = ~P2_REG3_REG_12_ | ~new_P2_ADD_1119_U17;
  assign new_P2_ADD_1119_U153 = ~new_P2_ADD_1119_U91 | ~new_P2_ADD_1119_U18;
  assign new_P2_ADD_1119_U154 = ~P2_REG3_REG_11_ | ~new_P2_ADD_1119_U83;
  assign new_P2_ADD_1119_U155 = ~new_P2_ADD_1119_U90 | ~new_P2_ADD_1119_U15;
  assign new_P2_ADD_1119_U156 = ~P2_REG3_REG_10_ | ~new_P2_ADD_1119_U14;
  assign new_P2_ADD_1119_U157 = ~new_P2_ADD_1119_U89 | ~new_P2_ADD_1119_U16;
  assign new_P2_SUB_1108_U6 = new_P2_SUB_1108_U172 & new_P2_SUB_1108_U40;
  assign new_P2_SUB_1108_U7 = new_P2_SUB_1108_U170 & new_P2_SUB_1108_U140;
  assign new_P2_SUB_1108_U8 = new_P2_SUB_1108_U169 & new_P2_SUB_1108_U37;
  assign new_P2_SUB_1108_U9 = new_P2_SUB_1108_U168 & new_P2_SUB_1108_U38;
  assign new_P2_SUB_1108_U10 = new_P2_SUB_1108_U166 & new_P2_SUB_1108_U143;
  assign new_P2_SUB_1108_U11 = new_P2_SUB_1108_U165 & new_P2_SUB_1108_U30;
  assign new_P2_SUB_1108_U12 = new_P2_SUB_1108_U164 & new_P2_SUB_1108_U36;
  assign new_P2_SUB_1108_U13 = new_P2_SUB_1108_U162 & new_P2_SUB_1108_U32;
  assign new_P2_SUB_1108_U14 = new_P2_SUB_1108_U160 & new_P2_SUB_1108_U33;
  assign new_P2_SUB_1108_U15 = new_P2_SUB_1108_U159 & new_P2_SUB_1108_U109;
  assign new_P2_SUB_1108_U16 = new_P2_SUB_1108_U157 & new_P2_SUB_1108_U29;
  assign new_P2_SUB_1108_U17 = new_P2_SUB_1108_U155 & new_P2_SUB_1108_U23;
  assign new_P2_SUB_1108_U18 = new_P2_SUB_1108_U138 & new_P2_SUB_1108_U128;
  assign new_P2_SUB_1108_U19 = new_P2_SUB_1108_U137 & new_P2_SUB_1108_U25;
  assign new_P2_SUB_1108_U20 = new_P2_SUB_1108_U136 & new_P2_SUB_1108_U26;
  assign new_P2_SUB_1108_U21 = new_P2_SUB_1108_U134 & new_P2_SUB_1108_U131;
  assign new_P2_SUB_1108_U22 = new_P2_SUB_1108_U133 & new_P2_SUB_1108_U24;
  assign new_P2_SUB_1108_U23 = P2_IR_REG_2_ | P2_IR_REG_1_ | P2_IR_REG_0_;
  assign new_P2_SUB_1108_U24 = ~new_P2_SUB_1108_U44 | ~new_P2_SUB_1108_U45 | ~new_P2_SUB_1108_U174;
  assign new_P2_SUB_1108_U25 = ~new_P2_SUB_1108_U46 | ~new_P2_SUB_1108_U174;
  assign new_P2_SUB_1108_U26 = ~new_P2_SUB_1108_U47 | ~new_P2_SUB_1108_U129;
  assign new_P2_SUB_1108_U27 = ~P2_IR_REG_7_;
  assign new_P2_SUB_1108_U28 = ~P2_IR_REG_3_;
  assign new_P2_SUB_1108_U29 = ~new_P2_SUB_1108_U57 | ~new_P2_SUB_1108_U52;
  assign new_P2_SUB_1108_U30 = ~new_P2_SUB_1108_U88 | ~new_P2_SUB_1108_U89 | ~new_P2_SUB_1108_U91 | ~new_P2_SUB_1108_U90;
  assign new_P2_SUB_1108_U31 = ~new_P2_SUB_1108_U92 | ~new_P2_SUB_1108_U144;
  assign new_P2_SUB_1108_U32 = ~new_P2_SUB_1108_U93 | ~new_P2_SUB_1108_U147;
  assign new_P2_SUB_1108_U33 = ~new_P2_SUB_1108_U149 | ~new_P2_SUB_1108_U34;
  assign new_P2_SUB_1108_U34 = ~P2_IR_REG_24_;
  assign new_P2_SUB_1108_U35 = ~new_P2_SUB_1108_U147 | ~new_P2_SUB_1108_U115;
  assign new_P2_SUB_1108_U36 = ~new_P2_SUB_1108_U94 | ~new_P2_SUB_1108_U144;
  assign new_P2_SUB_1108_U37 = ~new_P2_SUB_1108_U95 | ~new_P2_SUB_1108_U132;
  assign new_P2_SUB_1108_U38 = ~new_P2_SUB_1108_U96 | ~new_P2_SUB_1108_U141;
  assign new_P2_SUB_1108_U39 = ~P2_IR_REG_15_;
  assign new_P2_SUB_1108_U40 = ~new_P2_SUB_1108_U97 | ~new_P2_SUB_1108_U132;
  assign new_P2_SUB_1108_U41 = ~P2_IR_REG_11_;
  assign new_P2_SUB_1108_U42 = ~new_P2_SUB_1108_U196 | ~new_P2_SUB_1108_U195;
  assign new_P2_SUB_1108_U43 = ~new_P2_SUB_1108_U180 | ~new_P2_SUB_1108_U179;
  assign new_P2_SUB_1108_U44 = ~P2_IR_REG_6_ & ~P2_IR_REG_5_ & ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_1108_U45 = ~P2_IR_REG_7_ & ~P2_IR_REG_8_;
  assign new_P2_SUB_1108_U46 = ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_1108_U47 = ~P2_IR_REG_5_ & ~P2_IR_REG_6_;
  assign new_P2_SUB_1108_U48 = ~P2_IR_REG_13_ & ~P2_IR_REG_12_ & ~P2_IR_REG_10_ & ~P2_IR_REG_11_;
  assign new_P2_SUB_1108_U49 = ~P2_IR_REG_17_ & ~P2_IR_REG_16_ & ~P2_IR_REG_14_ & ~P2_IR_REG_15_;
  assign new_P2_SUB_1108_U50 = ~P2_IR_REG_0_ & ~P2_IR_REG_1_ & ~P2_IR_REG_18_ & ~P2_IR_REG_19_;
  assign new_P2_SUB_1108_U51 = ~P2_IR_REG_21_ & ~P2_IR_REG_22_ & ~P2_IR_REG_20_;
  assign new_P2_SUB_1108_U52 = new_P2_SUB_1108_U48 & new_P2_SUB_1108_U49 & new_P2_SUB_1108_U51 & new_P2_SUB_1108_U50;
  assign new_P2_SUB_1108_U53 = ~P2_IR_REG_26_ & ~P2_IR_REG_25_ & ~P2_IR_REG_23_ & ~P2_IR_REG_24_;
  assign new_P2_SUB_1108_U54 = ~P2_IR_REG_2_ & ~P2_IR_REG_29_ & ~P2_IR_REG_27_ & ~P2_IR_REG_28_;
  assign new_P2_SUB_1108_U55 = ~P2_IR_REG_6_ & ~P2_IR_REG_5_ & ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_1108_U56 = ~P2_IR_REG_8_ & ~P2_IR_REG_9_ & ~P2_IR_REG_7_;
  assign new_P2_SUB_1108_U57 = new_P2_SUB_1108_U53 & new_P2_SUB_1108_U54 & new_P2_SUB_1108_U56 & new_P2_SUB_1108_U55;
  assign new_P2_SUB_1108_U58 = ~P2_IR_REG_13_ & ~P2_IR_REG_12_ & ~P2_IR_REG_10_ & ~P2_IR_REG_11_;
  assign new_P2_SUB_1108_U59 = ~P2_IR_REG_17_ & ~P2_IR_REG_16_ & ~P2_IR_REG_14_ & ~P2_IR_REG_15_;
  assign new_P2_SUB_1108_U60 = ~P2_IR_REG_0_ & ~P2_IR_REG_1_ & ~P2_IR_REG_18_ & ~P2_IR_REG_19_;
  assign new_P2_SUB_1108_U61 = ~P2_IR_REG_21_ & ~P2_IR_REG_22_ & ~P2_IR_REG_20_;
  assign new_P2_SUB_1108_U62 = new_P2_SUB_1108_U58 & new_P2_SUB_1108_U59 & new_P2_SUB_1108_U61 & new_P2_SUB_1108_U60;
  assign new_P2_SUB_1108_U63 = ~P2_IR_REG_26_ & ~P2_IR_REG_25_ & ~P2_IR_REG_23_ & ~P2_IR_REG_24_;
  assign new_P2_SUB_1108_U64 = ~P2_IR_REG_28_ & ~P2_IR_REG_2_ & ~P2_IR_REG_27_;
  assign new_P2_SUB_1108_U65 = ~P2_IR_REG_6_ & ~P2_IR_REG_5_ & ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_1108_U66 = ~P2_IR_REG_8_ & ~P2_IR_REG_9_ & ~P2_IR_REG_7_;
  assign new_P2_SUB_1108_U67 = new_P2_SUB_1108_U63 & new_P2_SUB_1108_U64 & new_P2_SUB_1108_U66 & new_P2_SUB_1108_U65;
  assign new_P2_SUB_1108_U68 = ~P2_IR_REG_13_ & ~P2_IR_REG_12_ & ~P2_IR_REG_10_ & ~P2_IR_REG_11_;
  assign new_P2_SUB_1108_U69 = ~P2_IR_REG_15_ & ~P2_IR_REG_16_ & ~P2_IR_REG_14_;
  assign new_P2_SUB_1108_U70 = ~P2_IR_REG_1_ & ~P2_IR_REG_19_ & ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign new_P2_SUB_1108_U71 = ~P2_IR_REG_20_ & ~P2_IR_REG_21_ & ~P2_IR_REG_0_;
  assign new_P2_SUB_1108_U72 = new_P2_SUB_1108_U68 & new_P2_SUB_1108_U69 & new_P2_SUB_1108_U71 & new_P2_SUB_1108_U70;
  assign new_P2_SUB_1108_U73 = ~P2_IR_REG_25_ & ~P2_IR_REG_24_ & ~P2_IR_REG_22_ & ~P2_IR_REG_23_;
  assign new_P2_SUB_1108_U74 = ~P2_IR_REG_27_ & ~P2_IR_REG_2_ & ~P2_IR_REG_26_;
  assign new_P2_SUB_1108_U75 = ~P2_IR_REG_6_ & ~P2_IR_REG_5_ & ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_1108_U76 = ~P2_IR_REG_8_ & ~P2_IR_REG_9_ & ~P2_IR_REG_7_;
  assign new_P2_SUB_1108_U77 = new_P2_SUB_1108_U73 & new_P2_SUB_1108_U74 & new_P2_SUB_1108_U76 & new_P2_SUB_1108_U75;
  assign new_P2_SUB_1108_U78 = ~P2_IR_REG_13_ & ~P2_IR_REG_12_ & ~P2_IR_REG_10_ & ~P2_IR_REG_11_;
  assign new_P2_SUB_1108_U79 = ~P2_IR_REG_15_ & ~P2_IR_REG_16_ & ~P2_IR_REG_14_;
  assign new_P2_SUB_1108_U80 = ~P2_IR_REG_1_ & ~P2_IR_REG_19_ & ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign new_P2_SUB_1108_U81 = ~P2_IR_REG_20_ & ~P2_IR_REG_21_ & ~P2_IR_REG_0_;
  assign new_P2_SUB_1108_U82 = new_P2_SUB_1108_U78 & new_P2_SUB_1108_U79 & new_P2_SUB_1108_U81 & new_P2_SUB_1108_U80;
  assign new_P2_SUB_1108_U83 = ~P2_IR_REG_25_ & ~P2_IR_REG_24_ & ~P2_IR_REG_22_ & ~P2_IR_REG_23_;
  assign new_P2_SUB_1108_U84 = ~P2_IR_REG_2_ & ~P2_IR_REG_3_ & ~P2_IR_REG_26_;
  assign new_P2_SUB_1108_U85 = ~P2_IR_REG_5_ & ~P2_IR_REG_6_ & ~P2_IR_REG_4_;
  assign new_P2_SUB_1108_U86 = ~P2_IR_REG_8_ & ~P2_IR_REG_9_ & ~P2_IR_REG_7_;
  assign new_P2_SUB_1108_U87 = new_P2_SUB_1108_U83 & new_P2_SUB_1108_U84 & new_P2_SUB_1108_U86 & new_P2_SUB_1108_U85;
  assign new_P2_SUB_1108_U88 = ~P2_IR_REG_11_ & ~P2_IR_REG_10_ & ~P2_IR_REG_12_ & ~P2_IR_REG_13_ & ~P2_IR_REG_14_;
  assign new_P2_SUB_1108_U89 = ~P2_IR_REG_0_ & ~P2_IR_REG_1_ & ~P2_IR_REG_15_ & ~P2_IR_REG_16_;
  assign new_P2_SUB_1108_U90 = ~P2_IR_REG_5_ & ~P2_IR_REG_4_ & ~P2_IR_REG_2_ & ~P2_IR_REG_3_;
  assign new_P2_SUB_1108_U91 = ~P2_IR_REG_9_ & ~P2_IR_REG_8_ & ~P2_IR_REG_6_ & ~P2_IR_REG_7_;
  assign new_P2_SUB_1108_U92 = ~P2_IR_REG_20_ & ~P2_IR_REG_19_ & ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign new_P2_SUB_1108_U93 = ~P2_IR_REG_22_ & ~P2_IR_REG_23_ & ~P2_IR_REG_21_;
  assign new_P2_SUB_1108_U94 = ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign new_P2_SUB_1108_U95 = ~P2_IR_REG_9_ & ~P2_IR_REG_12_ & ~P2_IR_REG_10_ & ~P2_IR_REG_11_;
  assign new_P2_SUB_1108_U96 = ~P2_IR_REG_13_ & ~P2_IR_REG_14_;
  assign new_P2_SUB_1108_U97 = ~P2_IR_REG_10_ & ~P2_IR_REG_9_;
  assign new_P2_SUB_1108_U98 = ~P2_IR_REG_9_;
  assign new_P2_SUB_1108_U99 = new_P2_SUB_1108_U176 & new_P2_SUB_1108_U175;
  assign new_P2_SUB_1108_U100 = ~P2_IR_REG_5_;
  assign new_P2_SUB_1108_U101 = new_P2_SUB_1108_U178 & new_P2_SUB_1108_U177;
  assign new_P2_SUB_1108_U102 = ~P2_IR_REG_31_;
  assign new_P2_SUB_1108_U103 = ~P2_IR_REG_30_;
  assign new_P2_SUB_1108_U104 = new_P2_SUB_1108_U182 & new_P2_SUB_1108_U181;
  assign new_P2_SUB_1108_U105 = ~P2_IR_REG_28_;
  assign new_P2_SUB_1108_U106 = ~new_P2_SUB_1108_U77 | ~new_P2_SUB_1108_U72;
  assign new_P2_SUB_1108_U107 = new_P2_SUB_1108_U184 & new_P2_SUB_1108_U183;
  assign new_P2_SUB_1108_U108 = ~P2_IR_REG_27_;
  assign new_P2_SUB_1108_U109 = ~new_P2_SUB_1108_U87 | ~new_P2_SUB_1108_U82;
  assign new_P2_SUB_1108_U110 = new_P2_SUB_1108_U186 & new_P2_SUB_1108_U185;
  assign new_P2_SUB_1108_U111 = ~P2_IR_REG_25_;
  assign new_P2_SUB_1108_U112 = new_P2_SUB_1108_U188 & new_P2_SUB_1108_U187;
  assign new_P2_SUB_1108_U113 = ~P2_IR_REG_22_;
  assign new_P2_SUB_1108_U114 = new_P2_SUB_1108_U190 & new_P2_SUB_1108_U189;
  assign new_P2_SUB_1108_U115 = ~P2_IR_REG_21_;
  assign new_P2_SUB_1108_U116 = new_P2_SUB_1108_U192 & new_P2_SUB_1108_U191;
  assign new_P2_SUB_1108_U117 = ~P2_IR_REG_20_;
  assign new_P2_SUB_1108_U118 = ~new_P2_SUB_1108_U145 | ~new_P2_SUB_1108_U122;
  assign new_P2_SUB_1108_U119 = new_P2_SUB_1108_U194 & new_P2_SUB_1108_U193;
  assign new_P2_SUB_1108_U120 = ~P2_IR_REG_1_;
  assign new_P2_SUB_1108_U121 = ~P2_IR_REG_0_;
  assign new_P2_SUB_1108_U122 = ~P2_IR_REG_19_;
  assign new_P2_SUB_1108_U123 = new_P2_SUB_1108_U198 & new_P2_SUB_1108_U197;
  assign new_P2_SUB_1108_U124 = ~P2_IR_REG_17_;
  assign new_P2_SUB_1108_U125 = new_P2_SUB_1108_U200 & new_P2_SUB_1108_U199;
  assign new_P2_SUB_1108_U126 = ~P2_IR_REG_13_;
  assign new_P2_SUB_1108_U127 = new_P2_SUB_1108_U202 & new_P2_SUB_1108_U201;
  assign new_P2_SUB_1108_U128 = ~new_P2_SUB_1108_U174 | ~new_P2_SUB_1108_U28;
  assign new_P2_SUB_1108_U129 = ~new_P2_SUB_1108_U25;
  assign new_P2_SUB_1108_U130 = ~new_P2_SUB_1108_U26;
  assign new_P2_SUB_1108_U131 = ~new_P2_SUB_1108_U130 | ~new_P2_SUB_1108_U27;
  assign new_P2_SUB_1108_U132 = ~new_P2_SUB_1108_U24;
  assign new_P2_SUB_1108_U133 = ~P2_IR_REG_8_ | ~new_P2_SUB_1108_U131;
  assign new_P2_SUB_1108_U134 = ~P2_IR_REG_7_ | ~new_P2_SUB_1108_U26;
  assign new_P2_SUB_1108_U135 = ~new_P2_SUB_1108_U129 | ~new_P2_SUB_1108_U100;
  assign new_P2_SUB_1108_U136 = ~P2_IR_REG_6_ | ~new_P2_SUB_1108_U135;
  assign new_P2_SUB_1108_U137 = ~P2_IR_REG_4_ | ~new_P2_SUB_1108_U128;
  assign new_P2_SUB_1108_U138 = ~P2_IR_REG_3_ | ~new_P2_SUB_1108_U23;
  assign new_P2_SUB_1108_U139 = ~new_P2_SUB_1108_U40;
  assign new_P2_SUB_1108_U140 = ~new_P2_SUB_1108_U139 | ~new_P2_SUB_1108_U41;
  assign new_P2_SUB_1108_U141 = ~new_P2_SUB_1108_U37;
  assign new_P2_SUB_1108_U142 = ~new_P2_SUB_1108_U38;
  assign new_P2_SUB_1108_U143 = ~new_P2_SUB_1108_U142 | ~new_P2_SUB_1108_U39;
  assign new_P2_SUB_1108_U144 = ~new_P2_SUB_1108_U30;
  assign new_P2_SUB_1108_U145 = ~new_P2_SUB_1108_U36;
  assign new_P2_SUB_1108_U146 = ~new_P2_SUB_1108_U118;
  assign new_P2_SUB_1108_U147 = ~new_P2_SUB_1108_U31;
  assign new_P2_SUB_1108_U148 = ~new_P2_SUB_1108_U35;
  assign new_P2_SUB_1108_U149 = ~new_P2_SUB_1108_U32;
  assign new_P2_SUB_1108_U150 = ~new_P2_SUB_1108_U33;
  assign new_P2_SUB_1108_U151 = ~new_P2_SUB_1108_U109;
  assign new_P2_SUB_1108_U152 = ~new_P2_SUB_1108_U106;
  assign new_P2_SUB_1108_U153 = ~new_P2_SUB_1108_U29;
  assign new_P2_SUB_1108_U154 = P2_IR_REG_1_ | P2_IR_REG_0_;
  assign new_P2_SUB_1108_U155 = ~P2_IR_REG_2_ | ~new_P2_SUB_1108_U154;
  assign new_P2_SUB_1108_U156 = ~new_P2_SUB_1108_U67 | ~new_P2_SUB_1108_U62;
  assign new_P2_SUB_1108_U157 = ~P2_IR_REG_29_ | ~new_P2_SUB_1108_U156;
  assign new_P2_SUB_1108_U158 = ~new_P2_SUB_1108_U150 | ~new_P2_SUB_1108_U111;
  assign new_P2_SUB_1108_U159 = ~P2_IR_REG_26_ | ~new_P2_SUB_1108_U158;
  assign new_P2_SUB_1108_U160 = ~P2_IR_REG_24_ | ~new_P2_SUB_1108_U32;
  assign new_P2_SUB_1108_U161 = ~new_P2_SUB_1108_U148 | ~new_P2_SUB_1108_U113;
  assign new_P2_SUB_1108_U162 = ~P2_IR_REG_23_ | ~new_P2_SUB_1108_U161;
  assign new_P2_SUB_1108_U163 = ~new_P2_SUB_1108_U144 | ~new_P2_SUB_1108_U124;
  assign new_P2_SUB_1108_U164 = ~P2_IR_REG_18_ | ~new_P2_SUB_1108_U163;
  assign new_P2_SUB_1108_U165 = ~P2_IR_REG_16_ | ~new_P2_SUB_1108_U143;
  assign new_P2_SUB_1108_U166 = ~P2_IR_REG_15_ | ~new_P2_SUB_1108_U38;
  assign new_P2_SUB_1108_U167 = ~new_P2_SUB_1108_U141 | ~new_P2_SUB_1108_U126;
  assign new_P2_SUB_1108_U168 = ~P2_IR_REG_14_ | ~new_P2_SUB_1108_U167;
  assign new_P2_SUB_1108_U169 = ~P2_IR_REG_12_ | ~new_P2_SUB_1108_U140;
  assign new_P2_SUB_1108_U170 = ~P2_IR_REG_11_ | ~new_P2_SUB_1108_U40;
  assign new_P2_SUB_1108_U171 = ~new_P2_SUB_1108_U132 | ~new_P2_SUB_1108_U98;
  assign new_P2_SUB_1108_U172 = ~P2_IR_REG_10_ | ~new_P2_SUB_1108_U171;
  assign new_P2_SUB_1108_U173 = ~new_P2_SUB_1108_U153 | ~new_P2_SUB_1108_U103;
  assign new_P2_SUB_1108_U174 = ~new_P2_SUB_1108_U23;
  assign new_P2_SUB_1108_U175 = ~P2_IR_REG_9_ | ~new_P2_SUB_1108_U24;
  assign new_P2_SUB_1108_U176 = ~new_P2_SUB_1108_U132 | ~new_P2_SUB_1108_U98;
  assign new_P2_SUB_1108_U177 = ~P2_IR_REG_5_ | ~new_P2_SUB_1108_U25;
  assign new_P2_SUB_1108_U178 = ~new_P2_SUB_1108_U129 | ~new_P2_SUB_1108_U100;
  assign new_P2_SUB_1108_U179 = ~new_P2_SUB_1108_U173 | ~new_P2_SUB_1108_U102;
  assign new_P2_SUB_1108_U180 = ~P2_IR_REG_31_ | ~new_P2_SUB_1108_U153 | ~new_P2_SUB_1108_U103;
  assign new_P2_SUB_1108_U181 = ~P2_IR_REG_30_ | ~new_P2_SUB_1108_U29;
  assign new_P2_SUB_1108_U182 = ~new_P2_SUB_1108_U153 | ~new_P2_SUB_1108_U103;
  assign new_P2_SUB_1108_U183 = ~P2_IR_REG_28_ | ~new_P2_SUB_1108_U106;
  assign new_P2_SUB_1108_U184 = ~new_P2_SUB_1108_U152 | ~new_P2_SUB_1108_U105;
  assign new_P2_SUB_1108_U185 = ~P2_IR_REG_27_ | ~new_P2_SUB_1108_U109;
  assign new_P2_SUB_1108_U186 = ~new_P2_SUB_1108_U151 | ~new_P2_SUB_1108_U108;
  assign new_P2_SUB_1108_U187 = ~P2_IR_REG_25_ | ~new_P2_SUB_1108_U33;
  assign new_P2_SUB_1108_U188 = ~new_P2_SUB_1108_U150 | ~new_P2_SUB_1108_U111;
  assign new_P2_SUB_1108_U189 = ~P2_IR_REG_22_ | ~new_P2_SUB_1108_U35;
  assign new_P2_SUB_1108_U190 = ~new_P2_SUB_1108_U148 | ~new_P2_SUB_1108_U113;
  assign new_P2_SUB_1108_U191 = ~P2_IR_REG_21_ | ~new_P2_SUB_1108_U31;
  assign new_P2_SUB_1108_U192 = ~new_P2_SUB_1108_U147 | ~new_P2_SUB_1108_U115;
  assign new_P2_SUB_1108_U193 = ~P2_IR_REG_20_ | ~new_P2_SUB_1108_U118;
  assign new_P2_SUB_1108_U194 = ~new_P2_SUB_1108_U146 | ~new_P2_SUB_1108_U117;
  assign new_P2_SUB_1108_U195 = ~P2_IR_REG_1_ | ~new_P2_SUB_1108_U121;
  assign new_P2_SUB_1108_U196 = ~P2_IR_REG_0_ | ~new_P2_SUB_1108_U120;
  assign new_P2_SUB_1108_U197 = ~P2_IR_REG_19_ | ~new_P2_SUB_1108_U36;
  assign new_P2_SUB_1108_U198 = ~new_P2_SUB_1108_U145 | ~new_P2_SUB_1108_U122;
  assign new_P2_SUB_1108_U199 = ~P2_IR_REG_17_ | ~new_P2_SUB_1108_U30;
  assign new_P2_SUB_1108_U200 = ~new_P2_SUB_1108_U144 | ~new_P2_SUB_1108_U124;
  assign new_P2_SUB_1108_U201 = ~P2_IR_REG_13_ | ~new_P2_SUB_1108_U37;
  assign new_P2_SUB_1108_U202 = ~new_P2_SUB_1108_U141 | ~new_P2_SUB_1108_U126;
  assign new_P2_R1299_U6 = new_P2_U3061 & new_P2_R1299_U7;
  assign new_P2_R1299_U7 = ~new_P2_U3058;
  assign new_P2_R1312_U6 = new_P2_R1312_U171 & new_P2_R1312_U172 & new_P2_R1312_U170;
  assign new_P2_R1312_U7 = new_P2_R1312_U85 & new_P2_R1312_U84;
  assign new_P2_R1312_U8 = new_P2_R1312_U7 & new_P2_R1312_U173;
  assign new_P2_R1312_U9 = new_P2_R1312_U183 & new_P2_R1312_U182;
  assign new_P2_R1312_U10 = new_P2_R1312_U213 & new_P2_R1312_U212;
  assign new_P2_R1312_U11 = new_P2_R1312_U169 & new_P2_R1312_U14 & new_P2_R1312_U82;
  assign new_P2_R1312_U12 = new_P2_R1312_U154 & new_P2_R1312_U155 & new_P2_R1312_U157 & new_P2_R1312_U156;
  assign new_P2_R1312_U13 = new_P2_R1312_U173 & new_P2_R1312_U174 & new_P2_R1312_U176 & new_P2_R1312_U175;
  assign new_P2_R1312_U14 = new_P2_R1312_U164 & new_P2_R1312_U162 & new_P2_R1312_U161;
  assign new_P2_R1312_U15 = new_P2_R1312_U17 & new_P2_R1312_U165 & new_P2_R1312_U83 & new_P2_R1312_U6 & new_P2_R1312_U11;
  assign new_P2_R1312_U16 = new_P2_R1312_U165 & new_P2_R1312_U163;
  assign new_P2_R1312_U17 = new_P2_R1312_U225 & new_P2_R1312_U224;
  assign new_P2_R1312_U18 = ~new_P2_R1312_U144 | ~new_P2_R1312_U147 | ~new_P2_R1312_U150 | ~new_P2_R1312_U152 | ~new_P2_R1312_U151;
  assign new_P2_R1312_U19 = ~new_P2_U3090;
  assign new_P2_R1312_U20 = ~new_P2_U3093;
  assign new_P2_R1312_U21 = ~new_P2_U3091;
  assign new_P2_R1312_U22 = ~new_P2_U3092;
  assign new_P2_R1312_U23 = ~new_P2_U3126;
  assign new_P2_R1312_U24 = ~new_P2_U3123;
  assign new_P2_R1312_U25 = ~new_P2_U3089;
  assign new_P2_R1312_U26 = ~new_P2_U3121;
  assign new_P2_R1312_U27 = ~new_P2_U3105;
  assign new_P2_R1312_U28 = ~new_P2_U3106;
  assign new_P2_R1312_U29 = ~new_P2_U3108;
  assign new_P2_R1312_U30 = ~new_P2_U3107;
  assign new_P2_R1312_U31 = ~new_P2_U3109;
  assign new_P2_R1312_U32 = ~new_P2_U3110;
  assign new_P2_R1312_U33 = ~new_P2_U3111;
  assign new_P2_R1312_U34 = ~new_P2_U3112;
  assign new_P2_R1312_U35 = ~new_P2_U3115;
  assign new_P2_R1312_U36 = ~new_P2_U3116;
  assign new_P2_R1312_U37 = ~new_P2_U3114;
  assign new_P2_R1312_U38 = ~new_P2_U3113;
  assign new_P2_R1312_U39 = ~new_P2_U3104;
  assign new_P2_R1312_U40 = ~new_P2_U3094;
  assign new_P2_R1312_U41 = ~new_P2_U3102;
  assign new_P2_R1312_U42 = ~new_P2_U3101;
  assign new_P2_R1312_U43 = ~new_P2_U3103;
  assign new_P2_R1312_U44 = ~new_P2_U3100;
  assign new_P2_R1312_U45 = ~new_P2_U3099;
  assign new_P2_R1312_U46 = ~new_P2_U3095;
  assign new_P2_R1312_U47 = ~new_P2_U3097;
  assign new_P2_R1312_U48 = ~new_P2_U3098;
  assign new_P2_R1312_U49 = ~new_P2_U3096;
  assign new_P2_R1312_U50 = ~new_P2_U3149;
  assign new_P2_R1312_U51 = ~new_P2_U3117;
  assign new_P2_R1312_U52 = ~new_P2_U3118;
  assign new_P2_R1312_U53 = ~new_P2_U3119;
  assign new_P2_R1312_U54 = ~new_P2_U3151;
  assign new_P2_R1312_U55 = ~new_P2_U3127;
  assign new_P2_R1312_U56 = ~new_P2_U3125;
  assign new_P2_R1312_U57 = ~new_P2_U3124;
  assign new_P2_R1312_U58 = ~new_P2_U3140;
  assign new_P2_R1312_U59 = ~new_P2_U3141;
  assign new_P2_R1312_U60 = ~new_P2_U3143;
  assign new_P2_R1312_U61 = ~new_P2_U3128;
  assign new_P2_R1312_U62 = ~new_P2_U3129;
  assign new_P2_R1312_U63 = ~new_P2_U3131;
  assign new_P2_R1312_U64 = ~new_P2_U3134;
  assign new_P2_R1312_U65 = ~new_P2_U3135;
  assign new_P2_R1312_U66 = ~new_P2_U3137;
  assign new_P2_R1312_U67 = ~new_P2_U3146;
  assign new_P2_R1312_U68 = ~new_P2_U3147;
  assign new_P2_R1312_U69 = ~new_P2_U3133;
  assign new_P2_R1312_U70 = ~new_P2_U3139;
  assign new_P2_R1312_U71 = ~new_P2_U3145;
  assign new_P2_R1312_U72 = ~new_P2_U3130;
  assign new_P2_R1312_U73 = ~new_P2_U3132;
  assign new_P2_R1312_U74 = ~new_P2_U3136;
  assign new_P2_R1312_U75 = ~new_P2_U3138;
  assign new_P2_R1312_U76 = ~new_P2_U3142;
  assign new_P2_R1312_U77 = ~new_P2_U3144;
  assign new_P2_R1312_U78 = ~new_P2_U3148;
  assign new_P2_R1312_U79 = ~new_P2_U3150;
  assign new_P2_R1312_U80 = ~new_P2_U3122;
  assign new_P2_R1312_U81 = new_P2_R1312_U17 & new_P2_R1312_U166;
  assign new_P2_R1312_U82 = new_P2_R1312_U160 & new_P2_R1312_U159;
  assign new_P2_R1312_U83 = new_P2_R1312_U163 & new_P2_R1312_U158;
  assign new_P2_R1312_U84 = new_P2_R1312_U174 & new_P2_R1312_U175 & new_P2_R1312_U177 & new_P2_R1312_U176;
  assign new_P2_R1312_U85 = new_P2_R1312_U180 & new_P2_R1312_U179 & new_P2_R1312_U178;
  assign new_P2_R1312_U86 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U51;
  assign new_P2_R1312_U87 = new_P2_U3149 & new_P2_R1312_U12;
  assign new_P2_R1312_U88 = new_P2_R1312_U186 & new_P2_R1312_U173;
  assign new_P2_R1312_U89 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U88 & new_P2_R1312_U185;
  assign new_P2_R1312_U90 = new_P2_R1312_U91 & new_P2_R1312_U7 & new_P2_R1312_U187;
  assign new_P2_R1312_U91 = new_P2_R1312_U9 & new_P2_R1312_U12;
  assign new_P2_R1312_U92 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U53;
  assign new_P2_R1312_U93 = new_P2_R1312_U12 & new_P2_U3151 & new_P2_R1312_U9;
  assign new_P2_R1312_U94 = new_P2_U3127 & new_P2_R1312_U46;
  assign new_P2_R1312_U95 = new_P2_R1312_U194 & new_P2_R1312_U195;
  assign new_P2_R1312_U96 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168;
  assign new_P2_R1312_U97 = new_P2_R1312_U168 & new_P2_R1312_U173 & new_P2_R1312_U167 & new_P2_R1312_U29;
  assign new_P2_R1312_U98 = new_P2_U3140 & new_P2_R1312_U176 & new_P2_R1312_U174;
  assign new_P2_R1312_U99 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U31;
  assign new_P2_R1312_U100 = new_P2_R1312_U13 & new_P2_U3141;
  assign new_P2_R1312_U101 = new_P2_R1312_U168 & new_P2_R1312_U177 & new_P2_R1312_U167 & new_P2_R1312_U33;
  assign new_P2_R1312_U102 = new_P2_R1312_U103 & new_P2_R1312_U13;
  assign new_P2_R1312_U103 = new_P2_U3143 & new_P2_R1312_U178;
  assign new_P2_R1312_U104 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U49;
  assign new_P2_R1312_U105 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U164 & new_P2_R1312_U47;
  assign new_P2_R1312_U106 = new_P2_R1312_U168 & new_P2_R1312_U169 & new_P2_R1312_U167 & new_P2_R1312_U45;
  assign new_P2_R1312_U107 = new_P2_U3131 & new_P2_R1312_U16;
  assign new_P2_R1312_U108 = new_P2_R1312_U168 & new_P2_R1312_U171 & new_P2_R1312_U167 & new_P2_R1312_U41;
  assign new_P2_R1312_U109 = new_P2_U3134 & new_P2_R1312_U16;
  assign new_P2_R1312_U110 = new_P2_R1312_U168 & new_P2_R1312_U170 & new_P2_R1312_U167 & new_P2_R1312_U43;
  assign new_P2_R1312_U111 = new_P2_R1312_U166 & new_P2_R1312_U112 & new_P2_R1312_U17 & new_P2_R1312_U11 & new_P2_R1312_U171;
  assign new_P2_R1312_U112 = new_P2_U3135 & new_P2_R1312_U16;
  assign new_P2_R1312_U113 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U27;
  assign new_P2_R1312_U114 = new_P2_U3137 & new_P2_R1312_U168;
  assign new_P2_R1312_U115 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U157 & new_P2_R1312_U37;
  assign new_P2_R1312_U116 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U157 & new_P2_R1312_U156 & new_P2_R1312_U35;
  assign new_P2_R1312_U117 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U42;
  assign new_P2_R1312_U118 = new_P2_U3133 & new_P2_R1312_U16;
  assign new_P2_R1312_U119 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U30;
  assign new_P2_R1312_U120 = new_P2_U3139 & new_P2_R1312_U174 & new_P2_R1312_U173;
  assign new_P2_R1312_U121 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U38;
  assign new_P2_R1312_U122 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U164 & new_P2_R1312_U161 & new_P2_R1312_U48;
  assign new_P2_R1312_U123 = new_P2_R1312_U169 & new_P2_R1312_U168;
  assign new_P2_R1312_U124 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U160 & new_P2_R1312_U44;
  assign new_P2_R1312_U125 = new_P2_U3132 & new_P2_R1312_U16;
  assign new_P2_R1312_U126 = new_P2_R1312_U167 & new_P2_R1312_U39;
  assign new_P2_R1312_U127 = new_P2_R1312_U126 & new_P2_R1312_U17 & new_P2_R1312_U168;
  assign new_P2_R1312_U128 = new_P2_R1312_U6 & new_P2_U3136;
  assign new_P2_R1312_U129 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U28;
  assign new_P2_R1312_U130 = new_P2_U3138 & new_P2_R1312_U173;
  assign new_P2_R1312_U131 = new_P2_R1312_U166 & new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_R1312_U32;
  assign new_P2_R1312_U132 = new_P2_R1312_U133 & new_P2_R1312_U13;
  assign new_P2_R1312_U133 = new_P2_U3142 & new_P2_R1312_U177;
  assign new_P2_R1312_U134 = new_P2_R1312_U168 & new_P2_R1312_U177 & new_P2_R1312_U167 & new_P2_R1312_U34;
  assign new_P2_R1312_U135 = new_P2_R1312_U13 & new_P2_R1312_U136;
  assign new_P2_R1312_U136 = new_P2_U3144 & new_P2_R1312_U179 & new_P2_R1312_U178;
  assign new_P2_R1312_U137 = new_P2_R1312_U166 & new_P2_R1312_U36 & new_P2_R1312_U154 & new_P2_R1312_U157 & new_P2_R1312_U156;
  assign new_P2_R1312_U138 = new_P2_R1312_U167 & new_P2_R1312_U168 & new_P2_U3148 & new_P2_R1312_U8;
  assign new_P2_R1312_U139 = new_P2_R1312_U168 & new_P2_R1312_U221 & new_P2_R1312_U167 & new_P2_R1312_U52;
  assign new_P2_R1312_U140 = new_P2_U3150 & new_P2_R1312_U12;
  assign new_P2_R1312_U141 = new_P2_R1312_U181 & new_P2_R1312_U153;
  assign new_P2_R1312_U142 = new_P2_R1312_U192 & new_P2_R1312_U188;
  assign new_P2_R1312_U143 = new_P2_R1312_U198 & new_P2_R1312_U199 & new_P2_R1312_U197;
  assign new_P2_R1312_U144 = new_P2_R1312_U143 & new_P2_R1312_U142 & new_P2_R1312_U141;
  assign new_P2_R1312_U145 = new_P2_R1312_U203 & new_P2_R1312_U202;
  assign new_P2_R1312_U146 = new_P2_R1312_U205 & new_P2_R1312_U204;
  assign new_P2_R1312_U147 = new_P2_R1312_U206 & new_P2_R1312_U146 & new_P2_R1312_U145 & new_P2_R1312_U201 & new_P2_R1312_U200;
  assign new_P2_R1312_U148 = new_P2_R1312_U210 & new_P2_R1312_U209;
  assign new_P2_R1312_U149 = new_P2_R1312_U214 & new_P2_R1312_U215;
  assign new_P2_R1312_U150 = new_P2_R1312_U211 & new_P2_R1312_U149 & new_P2_R1312_U148 & new_P2_R1312_U208 & new_P2_R1312_U207;
  assign new_P2_R1312_U151 = new_P2_R1312_U216 & new_P2_R1312_U217 & new_P2_R1312_U219 & new_P2_R1312_U218;
  assign new_P2_R1312_U152 = new_P2_R1312_U222 & new_P2_R1312_U10 & new_P2_R1312_U220;
  assign new_P2_R1312_U153 = ~new_P2_R1312_U81 | ~new_P2_R1312_U191;
  assign new_P2_R1312_U154 = ~new_P2_U3115 | ~new_P2_R1312_U68;
  assign new_P2_R1312_U155 = ~new_P2_U3116 | ~new_P2_R1312_U78;
  assign new_P2_R1312_U156 = ~new_P2_U3114 | ~new_P2_R1312_U67;
  assign new_P2_R1312_U157 = ~new_P2_U3113 | ~new_P2_R1312_U71;
  assign new_P2_R1312_U158 = ~new_P2_U3104 | ~new_P2_R1312_U74;
  assign new_P2_R1312_U159 = ~new_P2_U3100 | ~new_P2_R1312_U73;
  assign new_P2_R1312_U160 = ~new_P2_U3099 | ~new_P2_R1312_U63;
  assign new_P2_R1312_U161 = ~new_P2_U3097 | ~new_P2_R1312_U62;
  assign new_P2_R1312_U162 = ~new_P2_U3098 | ~new_P2_R1312_U72;
  assign new_P2_R1312_U163 = ~new_P2_U3094 | ~new_P2_R1312_U23;
  assign new_P2_R1312_U164 = ~new_P2_U3096 | ~new_P2_R1312_U61;
  assign new_P2_R1312_U165 = ~new_P2_U3093 | ~new_P2_R1312_U56;
  assign new_P2_R1312_U166 = ~new_P2_U3090 | ~new_P2_R1312_U80;
  assign new_P2_R1312_U167 = ~new_P2_U3091 | ~new_P2_R1312_U24;
  assign new_P2_R1312_U168 = ~new_P2_U3092 | ~new_P2_R1312_U57;
  assign new_P2_R1312_U169 = ~new_P2_U3095 | ~new_P2_R1312_U55;
  assign new_P2_R1312_U170 = ~new_P2_U3102 | ~new_P2_R1312_U64;
  assign new_P2_R1312_U171 = ~new_P2_U3101 | ~new_P2_R1312_U69;
  assign new_P2_R1312_U172 = ~new_P2_U3103 | ~new_P2_R1312_U65;
  assign new_P2_R1312_U173 = ~new_P2_U3105 | ~new_P2_R1312_U66;
  assign new_P2_R1312_U174 = ~new_P2_U3106 | ~new_P2_R1312_U75;
  assign new_P2_R1312_U175 = ~new_P2_U3108 | ~new_P2_R1312_U58;
  assign new_P2_R1312_U176 = ~new_P2_U3107 | ~new_P2_R1312_U70;
  assign new_P2_R1312_U177 = ~new_P2_U3109 | ~new_P2_R1312_U59;
  assign new_P2_R1312_U178 = ~new_P2_U3110 | ~new_P2_R1312_U76;
  assign new_P2_R1312_U179 = ~new_P2_U3111 | ~new_P2_R1312_U60;
  assign new_P2_R1312_U180 = ~new_P2_U3112 | ~new_P2_R1312_U77;
  assign new_P2_R1312_U181 = ~new_P2_R1312_U86 | ~new_P2_R1312_U15 | ~new_P2_R1312_U8 | ~new_P2_R1312_U87;
  assign new_P2_R1312_U182 = ~new_P2_U3117 | ~new_P2_R1312_U50;
  assign new_P2_R1312_U183 = ~new_P2_U3118 | ~new_P2_R1312_U79;
  assign new_P2_R1312_U184 = ~new_P2_U3152 | ~new_P2_U3153;
  assign new_P2_R1312_U185 = ~new_P2_U3120 | ~new_P2_R1312_U184;
  assign new_P2_R1312_U186 = ~new_P2_U3119 | ~new_P2_R1312_U54;
  assign new_P2_R1312_U187 = new_P2_U3152 | new_P2_U3153;
  assign new_P2_R1312_U188 = ~new_P2_R1312_U89 | ~new_P2_R1312_U15 | ~new_P2_R1312_U90;
  assign new_P2_R1312_U189 = ~new_P2_R1312_U168 | ~new_P2_U3126 | ~new_P2_R1312_U167 | ~new_P2_R1312_U165 | ~new_P2_R1312_U40;
  assign new_P2_R1312_U190 = ~new_P2_U3123 | ~new_P2_R1312_U21;
  assign new_P2_R1312_U191 = ~new_P2_R1312_U190 | ~new_P2_R1312_U189;
  assign new_P2_R1312_U192 = ~new_P2_R1312_U92 | ~new_P2_R1312_U15 | ~new_P2_R1312_U168 | ~new_P2_R1312_U8 | ~new_P2_R1312_U93;
  assign new_P2_R1312_U193 = ~new_P2_R1312_U94 | ~new_P2_R1312_U16;
  assign new_P2_R1312_U194 = ~new_P2_U3125 | ~new_P2_R1312_U20;
  assign new_P2_R1312_U195 = ~new_P2_U3124 | ~new_P2_R1312_U22;
  assign new_P2_R1312_U196 = ~new_P2_R1312_U95 | ~new_P2_R1312_U193;
  assign new_P2_R1312_U197 = ~new_P2_R1312_U96 | ~new_P2_R1312_U17 | ~new_P2_R1312_U196;
  assign new_P2_R1312_U198 = ~new_P2_R1312_U97 | ~new_P2_R1312_U166 | ~new_P2_R1312_U98 | ~new_P2_R1312_U15;
  assign new_P2_R1312_U199 = ~new_P2_R1312_U99 | ~new_P2_R1312_U100 | ~new_P2_R1312_U15;
  assign new_P2_R1312_U200 = ~new_P2_R1312_U101 | ~new_P2_R1312_U166 | ~new_P2_R1312_U15 | ~new_P2_R1312_U102;
  assign new_P2_R1312_U201 = ~new_P2_R1312_U104 | ~new_P2_R1312_U169 | ~new_P2_R1312_U17 | ~new_P2_U3128 | ~new_P2_R1312_U16;
  assign new_P2_R1312_U202 = ~new_P2_R1312_U105 | ~new_P2_R1312_U169 | ~new_P2_R1312_U17 | ~new_P2_U3129 | ~new_P2_R1312_U16;
  assign new_P2_R1312_U203 = ~new_P2_R1312_U106 | ~new_P2_R1312_U166 | ~new_P2_R1312_U107 | ~new_P2_R1312_U17 | ~new_P2_R1312_U14;
  assign new_P2_R1312_U204 = ~new_P2_R1312_U108 | ~new_P2_R1312_U166 | ~new_P2_R1312_U109 | ~new_P2_R1312_U17 | ~new_P2_R1312_U11;
  assign new_P2_R1312_U205 = ~new_P2_R1312_U110 | ~new_P2_R1312_U111;
  assign new_P2_R1312_U206 = ~new_P2_R1312_U113 | ~new_P2_R1312_U114 | ~new_P2_R1312_U15;
  assign new_P2_R1312_U207 = ~new_P2_R1312_U115 | ~new_P2_R1312_U15 | ~new_P2_R1312_U168 | ~new_P2_U3146 | ~new_P2_R1312_U8;
  assign new_P2_R1312_U208 = ~new_P2_R1312_U116 | ~new_P2_R1312_U15 | ~new_P2_R1312_U168 | ~new_P2_U3147 | ~new_P2_R1312_U8;
  assign new_P2_R1312_U209 = ~new_P2_R1312_U117 | ~new_P2_R1312_U118 | ~new_P2_R1312_U17 | ~new_P2_R1312_U11;
  assign new_P2_R1312_U210 = ~new_P2_R1312_U119 | ~new_P2_R1312_U120 | ~new_P2_R1312_U15;
  assign new_P2_R1312_U211 = ~new_P2_R1312_U121 | ~new_P2_R1312_U15 | ~new_P2_R1312_U8 | ~new_P2_U3145;
  assign new_P2_R1312_U212 = ~new_P2_R1312_U223 | ~new_P2_R1312_U227 | ~new_P2_R1312_U226;
  assign new_P2_R1312_U213 = ~new_P2_R1312_U19 | ~new_P2_R1312_U17 | ~new_P2_U3122;
  assign new_P2_R1312_U214 = ~new_P2_R1312_U122 | ~new_P2_R1312_U123 | ~new_P2_R1312_U17 | ~new_P2_U3130 | ~new_P2_R1312_U16;
  assign new_P2_R1312_U215 = ~new_P2_R1312_U124 | ~new_P2_R1312_U125 | ~new_P2_R1312_U17 | ~new_P2_R1312_U14 | ~new_P2_R1312_U169;
  assign new_P2_R1312_U216 = ~new_P2_R1312_U127 | ~new_P2_R1312_U166 | ~new_P2_R1312_U16 | ~new_P2_R1312_U11 | ~new_P2_R1312_U128;
  assign new_P2_R1312_U217 = ~new_P2_R1312_U129 | ~new_P2_R1312_U130 | ~new_P2_R1312_U15;
  assign new_P2_R1312_U218 = ~new_P2_R1312_U131 | ~new_P2_R1312_U15 | ~new_P2_R1312_U132;
  assign new_P2_R1312_U219 = ~new_P2_R1312_U134 | ~new_P2_R1312_U166 | ~new_P2_R1312_U15 | ~new_P2_R1312_U135;
  assign new_P2_R1312_U220 = ~new_P2_R1312_U137 | ~new_P2_R1312_U15 | ~new_P2_R1312_U138;
  assign new_P2_R1312_U221 = ~new_P2_U3117 | ~new_P2_R1312_U50;
  assign new_P2_R1312_U222 = ~new_P2_R1312_U139 | ~new_P2_R1312_U166 | ~new_P2_R1312_U15 | ~new_P2_R1312_U8 | ~new_P2_R1312_U140;
  assign new_P2_R1312_U223 = ~new_P2_U3121 | ~new_P2_U3089;
  assign new_P2_R1312_U224 = ~new_P2_U3089 | ~new_P2_R1312_U26;
  assign new_P2_R1312_U225 = ~new_P2_U3121 | ~new_P2_R1312_U25;
  assign new_P2_R1312_U226 = new_P2_U3154 | new_P2_U3121;
  assign new_P2_R1312_U227 = ~new_P2_U3154 | ~new_P2_R1312_U25;
  assign new_P2_R1335_U6 = ~new_P2_U3061;
  assign new_P2_R1335_U7 = ~new_P2_U3058;
  assign new_P2_R1335_U8 = new_P2_R1335_U10 & new_P2_R1335_U9;
  assign new_P2_R1335_U9 = ~new_P2_U3058 | ~new_P2_R1335_U6;
  assign new_P2_R1335_U10 = ~new_P2_U3061 | ~new_P2_R1335_U7;
  assign new_P2_R1209_U4 = new_P2_R1209_U95 & new_P2_R1209_U94;
  assign new_P2_R1209_U5 = new_P2_R1209_U96 & new_P2_R1209_U97;
  assign new_P2_R1209_U6 = new_P2_R1209_U113 & new_P2_R1209_U112;
  assign new_P2_R1209_U7 = new_P2_R1209_U155 & new_P2_R1209_U154;
  assign new_P2_R1209_U8 = new_P2_R1209_U164 & new_P2_R1209_U163;
  assign new_P2_R1209_U9 = new_P2_R1209_U182 & new_P2_R1209_U181;
  assign new_P2_R1209_U10 = new_P2_R1209_U218 & new_P2_R1209_U215;
  assign new_P2_R1209_U11 = new_P2_R1209_U211 & new_P2_R1209_U208;
  assign new_P2_R1209_U12 = new_P2_R1209_U202 & new_P2_R1209_U199;
  assign new_P2_R1209_U13 = new_P2_R1209_U196 & new_P2_R1209_U192;
  assign new_P2_R1209_U14 = new_P2_R1209_U151 & new_P2_R1209_U148;
  assign new_P2_R1209_U15 = new_P2_R1209_U143 & new_P2_R1209_U140;
  assign new_P2_R1209_U16 = new_P2_R1209_U129 & new_P2_R1209_U126;
  assign new_P2_R1209_U17 = ~P2_REG1_REG_6_;
  assign new_P2_R1209_U18 = ~new_P2_U3446;
  assign new_P2_R1209_U19 = ~new_P2_U3449;
  assign new_P2_R1209_U20 = ~new_P2_U3446 | ~P2_REG1_REG_6_;
  assign new_P2_R1209_U21 = ~P2_REG1_REG_7_;
  assign new_P2_R1209_U22 = ~P2_REG1_REG_4_;
  assign new_P2_R1209_U23 = ~new_P2_U3440;
  assign new_P2_R1209_U24 = ~new_P2_U3443;
  assign new_P2_R1209_U25 = ~P2_REG1_REG_2_;
  assign new_P2_R1209_U26 = ~new_P2_U3434;
  assign new_P2_R1209_U27 = ~P2_REG1_REG_0_;
  assign new_P2_R1209_U28 = ~new_P2_U3425;
  assign new_P2_R1209_U29 = ~new_P2_U3425 | ~P2_REG1_REG_0_;
  assign new_P2_R1209_U30 = ~P2_REG1_REG_3_;
  assign new_P2_R1209_U31 = ~new_P2_U3437;
  assign new_P2_R1209_U32 = ~new_P2_U3440 | ~P2_REG1_REG_4_;
  assign new_P2_R1209_U33 = ~P2_REG1_REG_5_;
  assign new_P2_R1209_U34 = ~P2_REG1_REG_8_;
  assign new_P2_R1209_U35 = ~new_P2_U3452;
  assign new_P2_R1209_U36 = ~new_P2_U3455;
  assign new_P2_R1209_U37 = ~P2_REG1_REG_9_;
  assign new_P2_R1209_U38 = ~new_P2_R1209_U49 | ~new_P2_R1209_U121;
  assign new_P2_R1209_U39 = ~new_P2_R1209_U109 | ~new_P2_R1209_U110 | ~new_P2_R1209_U108;
  assign new_P2_R1209_U40 = ~new_P2_R1209_U98 | ~new_P2_R1209_U99;
  assign new_P2_R1209_U41 = ~P2_REG1_REG_1_ | ~new_P2_U3431;
  assign new_P2_R1209_U42 = ~new_P2_R1209_U135 | ~new_P2_R1209_U136 | ~new_P2_R1209_U134;
  assign new_P2_R1209_U43 = ~new_P2_R1209_U132 | ~new_P2_R1209_U131;
  assign new_P2_R1209_U44 = ~P2_REG1_REG_16_;
  assign new_P2_R1209_U45 = ~new_P2_U3476;
  assign new_P2_R1209_U46 = ~new_P2_U3479;
  assign new_P2_R1209_U47 = ~new_P2_U3476 | ~P2_REG1_REG_16_;
  assign new_P2_R1209_U48 = ~P2_REG1_REG_17_;
  assign new_P2_R1209_U49 = ~new_P2_U3452 | ~P2_REG1_REG_8_;
  assign new_P2_R1209_U50 = ~P2_REG1_REG_10_;
  assign new_P2_R1209_U51 = ~new_P2_U3458;
  assign new_P2_R1209_U52 = ~P2_REG1_REG_12_;
  assign new_P2_R1209_U53 = ~new_P2_U3464;
  assign new_P2_R1209_U54 = ~P2_REG1_REG_11_;
  assign new_P2_R1209_U55 = ~new_P2_U3461;
  assign new_P2_R1209_U56 = ~new_P2_U3461 | ~P2_REG1_REG_11_;
  assign new_P2_R1209_U57 = ~P2_REG1_REG_13_;
  assign new_P2_R1209_U58 = ~new_P2_U3467;
  assign new_P2_R1209_U59 = ~P2_REG1_REG_14_;
  assign new_P2_R1209_U60 = ~new_P2_U3470;
  assign new_P2_R1209_U61 = ~P2_REG1_REG_15_;
  assign new_P2_R1209_U62 = ~new_P2_U3473;
  assign new_P2_R1209_U63 = ~P2_REG1_REG_18_;
  assign new_P2_R1209_U64 = ~new_P2_U3482;
  assign new_P2_R1209_U65 = ~new_P2_R1209_U187 | ~new_P2_R1209_U186 | ~new_P2_R1209_U185;
  assign new_P2_R1209_U66 = ~new_P2_R1209_U179 | ~new_P2_R1209_U178;
  assign new_P2_R1209_U67 = ~new_P2_R1209_U56 | ~new_P2_R1209_U204;
  assign new_P2_R1209_U68 = ~new_P2_R1209_U259 | ~new_P2_R1209_U258;
  assign new_P2_R1209_U69 = ~new_P2_R1209_U308 | ~new_P2_R1209_U307;
  assign new_P2_R1209_U70 = ~new_P2_R1209_U231 | ~new_P2_R1209_U230;
  assign new_P2_R1209_U71 = ~new_P2_R1209_U236 | ~new_P2_R1209_U235;
  assign new_P2_R1209_U72 = ~new_P2_R1209_U243 | ~new_P2_R1209_U242;
  assign new_P2_R1209_U73 = ~new_P2_R1209_U250 | ~new_P2_R1209_U249;
  assign new_P2_R1209_U74 = ~new_P2_R1209_U255 | ~new_P2_R1209_U254;
  assign new_P2_R1209_U75 = ~new_P2_R1209_U271 | ~new_P2_R1209_U270;
  assign new_P2_R1209_U76 = ~new_P2_R1209_U278 | ~new_P2_R1209_U277;
  assign new_P2_R1209_U77 = ~new_P2_R1209_U285 | ~new_P2_R1209_U284;
  assign new_P2_R1209_U78 = ~new_P2_R1209_U292 | ~new_P2_R1209_U291;
  assign new_P2_R1209_U79 = ~new_P2_R1209_U299 | ~new_P2_R1209_U298;
  assign new_P2_R1209_U80 = ~new_P2_R1209_U304 | ~new_P2_R1209_U303;
  assign new_P2_R1209_U81 = ~new_P2_R1209_U118 | ~new_P2_R1209_U117 | ~new_P2_R1209_U116;
  assign new_P2_R1209_U82 = ~new_P2_R1209_U133 | ~new_P2_R1209_U145;
  assign new_P2_R1209_U83 = ~new_P2_R1209_U41 | ~new_P2_R1209_U152;
  assign new_P2_R1209_U84 = ~new_P2_U3424;
  assign new_P2_R1209_U85 = ~P2_REG1_REG_19_;
  assign new_P2_R1209_U86 = ~new_P2_R1209_U175 | ~new_P2_R1209_U174;
  assign new_P2_R1209_U87 = ~new_P2_R1209_U171 | ~new_P2_R1209_U170;
  assign new_P2_R1209_U88 = ~new_P2_R1209_U161 | ~new_P2_R1209_U160;
  assign new_P2_R1209_U89 = ~new_P2_R1209_U32;
  assign new_P2_R1209_U90 = ~P2_REG1_REG_9_ | ~new_P2_U3455;
  assign new_P2_R1209_U91 = ~new_P2_U3464 | ~P2_REG1_REG_12_;
  assign new_P2_R1209_U92 = ~new_P2_R1209_U56;
  assign new_P2_R1209_U93 = ~new_P2_R1209_U49;
  assign new_P2_R1209_U94 = new_P2_U3443 | P2_REG1_REG_5_;
  assign new_P2_R1209_U95 = new_P2_U3440 | P2_REG1_REG_4_;
  assign new_P2_R1209_U96 = P2_REG1_REG_3_ | new_P2_U3437;
  assign new_P2_R1209_U97 = P2_REG1_REG_2_ | new_P2_U3434;
  assign new_P2_R1209_U98 = ~new_P2_R1209_U29;
  assign new_P2_R1209_U99 = P2_REG1_REG_1_ | new_P2_U3431;
  assign new_P2_R1209_U100 = ~new_P2_R1209_U40;
  assign new_P2_R1209_U101 = ~new_P2_R1209_U41;
  assign new_P2_R1209_U102 = ~new_P2_R1209_U40 | ~new_P2_R1209_U41;
  assign new_P2_R1209_U103 = ~new_P2_R1209_U96 | ~P2_REG1_REG_2_ | ~new_P2_U3434;
  assign new_P2_R1209_U104 = ~new_P2_R1209_U5 | ~new_P2_R1209_U102;
  assign new_P2_R1209_U105 = ~new_P2_U3437 | ~P2_REG1_REG_3_;
  assign new_P2_R1209_U106 = ~new_P2_R1209_U104 | ~new_P2_R1209_U105 | ~new_P2_R1209_U103;
  assign new_P2_R1209_U107 = ~new_P2_R1209_U33 | ~new_P2_R1209_U32;
  assign new_P2_R1209_U108 = ~new_P2_U3443 | ~new_P2_R1209_U107;
  assign new_P2_R1209_U109 = ~new_P2_R1209_U4 | ~new_P2_R1209_U106;
  assign new_P2_R1209_U110 = ~P2_REG1_REG_5_ | ~new_P2_R1209_U89;
  assign new_P2_R1209_U111 = ~new_P2_R1209_U39;
  assign new_P2_R1209_U112 = new_P2_U3449 | P2_REG1_REG_7_;
  assign new_P2_R1209_U113 = new_P2_U3446 | P2_REG1_REG_6_;
  assign new_P2_R1209_U114 = ~new_P2_R1209_U20;
  assign new_P2_R1209_U115 = ~new_P2_R1209_U21 | ~new_P2_R1209_U20;
  assign new_P2_R1209_U116 = ~new_P2_U3449 | ~new_P2_R1209_U115;
  assign new_P2_R1209_U117 = ~P2_REG1_REG_7_ | ~new_P2_R1209_U114;
  assign new_P2_R1209_U118 = ~new_P2_R1209_U6 | ~new_P2_R1209_U39;
  assign new_P2_R1209_U119 = ~new_P2_R1209_U81;
  assign new_P2_R1209_U120 = P2_REG1_REG_8_ | new_P2_U3452;
  assign new_P2_R1209_U121 = ~new_P2_R1209_U120 | ~new_P2_R1209_U81;
  assign new_P2_R1209_U122 = ~new_P2_R1209_U38;
  assign new_P2_R1209_U123 = new_P2_U3455 | P2_REG1_REG_9_;
  assign new_P2_R1209_U124 = P2_REG1_REG_6_ | new_P2_U3446;
  assign new_P2_R1209_U125 = ~new_P2_R1209_U124 | ~new_P2_R1209_U39;
  assign new_P2_R1209_U126 = ~new_P2_R1209_U125 | ~new_P2_R1209_U20 | ~new_P2_R1209_U238 | ~new_P2_R1209_U237;
  assign new_P2_R1209_U127 = ~new_P2_R1209_U111 | ~new_P2_R1209_U20;
  assign new_P2_R1209_U128 = ~P2_REG1_REG_7_ | ~new_P2_U3449;
  assign new_P2_R1209_U129 = ~new_P2_R1209_U127 | ~new_P2_R1209_U128 | ~new_P2_R1209_U6;
  assign new_P2_R1209_U130 = new_P2_U3446 | P2_REG1_REG_6_;
  assign new_P2_R1209_U131 = ~new_P2_R1209_U101 | ~new_P2_R1209_U97;
  assign new_P2_R1209_U132 = ~new_P2_U3434 | ~P2_REG1_REG_2_;
  assign new_P2_R1209_U133 = ~new_P2_R1209_U43;
  assign new_P2_R1209_U134 = ~new_P2_R1209_U100 | ~new_P2_R1209_U5;
  assign new_P2_R1209_U135 = ~new_P2_R1209_U43 | ~new_P2_R1209_U96;
  assign new_P2_R1209_U136 = ~new_P2_U3437 | ~P2_REG1_REG_3_;
  assign new_P2_R1209_U137 = ~new_P2_R1209_U42;
  assign new_P2_R1209_U138 = P2_REG1_REG_4_ | new_P2_U3440;
  assign new_P2_R1209_U139 = ~new_P2_R1209_U138 | ~new_P2_R1209_U42;
  assign new_P2_R1209_U140 = ~new_P2_R1209_U139 | ~new_P2_R1209_U32 | ~new_P2_R1209_U245 | ~new_P2_R1209_U244;
  assign new_P2_R1209_U141 = ~new_P2_R1209_U137 | ~new_P2_R1209_U32;
  assign new_P2_R1209_U142 = ~P2_REG1_REG_5_ | ~new_P2_U3443;
  assign new_P2_R1209_U143 = ~new_P2_R1209_U141 | ~new_P2_R1209_U142 | ~new_P2_R1209_U4;
  assign new_P2_R1209_U144 = new_P2_U3440 | P2_REG1_REG_4_;
  assign new_P2_R1209_U145 = ~new_P2_R1209_U100 | ~new_P2_R1209_U97;
  assign new_P2_R1209_U146 = ~new_P2_R1209_U82;
  assign new_P2_R1209_U147 = ~new_P2_U3437 | ~P2_REG1_REG_3_;
  assign new_P2_R1209_U148 = ~new_P2_R1209_U40 | ~new_P2_R1209_U41 | ~new_P2_R1209_U257 | ~new_P2_R1209_U256;
  assign new_P2_R1209_U149 = ~new_P2_R1209_U41 | ~new_P2_R1209_U40;
  assign new_P2_R1209_U150 = ~new_P2_U3434 | ~P2_REG1_REG_2_;
  assign new_P2_R1209_U151 = ~new_P2_R1209_U149 | ~new_P2_R1209_U150 | ~new_P2_R1209_U97;
  assign new_P2_R1209_U152 = P2_REG1_REG_1_ | new_P2_U3431;
  assign new_P2_R1209_U153 = ~new_P2_R1209_U83;
  assign new_P2_R1209_U154 = new_P2_U3455 | P2_REG1_REG_9_;
  assign new_P2_R1209_U155 = new_P2_U3458 | P2_REG1_REG_10_;
  assign new_P2_R1209_U156 = ~new_P2_R1209_U93 | ~new_P2_R1209_U7;
  assign new_P2_R1209_U157 = ~new_P2_U3458 | ~P2_REG1_REG_10_;
  assign new_P2_R1209_U158 = ~new_P2_R1209_U156 | ~new_P2_R1209_U157 | ~new_P2_R1209_U90;
  assign new_P2_R1209_U159 = P2_REG1_REG_10_ | new_P2_U3458;
  assign new_P2_R1209_U160 = ~new_P2_R1209_U81 | ~new_P2_R1209_U120 | ~new_P2_R1209_U7;
  assign new_P2_R1209_U161 = ~new_P2_R1209_U159 | ~new_P2_R1209_U158;
  assign new_P2_R1209_U162 = ~new_P2_R1209_U88;
  assign new_P2_R1209_U163 = new_P2_U3467 | P2_REG1_REG_13_;
  assign new_P2_R1209_U164 = new_P2_U3464 | P2_REG1_REG_12_;
  assign new_P2_R1209_U165 = ~new_P2_R1209_U92 | ~new_P2_R1209_U8;
  assign new_P2_R1209_U166 = ~new_P2_U3467 | ~P2_REG1_REG_13_;
  assign new_P2_R1209_U167 = ~new_P2_R1209_U165 | ~new_P2_R1209_U166 | ~new_P2_R1209_U91;
  assign new_P2_R1209_U168 = P2_REG1_REG_11_ | new_P2_U3461;
  assign new_P2_R1209_U169 = P2_REG1_REG_13_ | new_P2_U3467;
  assign new_P2_R1209_U170 = ~new_P2_R1209_U88 | ~new_P2_R1209_U168 | ~new_P2_R1209_U8;
  assign new_P2_R1209_U171 = ~new_P2_R1209_U169 | ~new_P2_R1209_U167;
  assign new_P2_R1209_U172 = ~new_P2_R1209_U87;
  assign new_P2_R1209_U173 = P2_REG1_REG_14_ | new_P2_U3470;
  assign new_P2_R1209_U174 = ~new_P2_R1209_U173 | ~new_P2_R1209_U87;
  assign new_P2_R1209_U175 = ~new_P2_U3470 | ~P2_REG1_REG_14_;
  assign new_P2_R1209_U176 = ~new_P2_R1209_U86;
  assign new_P2_R1209_U177 = P2_REG1_REG_15_ | new_P2_U3473;
  assign new_P2_R1209_U178 = ~new_P2_R1209_U177 | ~new_P2_R1209_U86;
  assign new_P2_R1209_U179 = ~new_P2_U3473 | ~P2_REG1_REG_15_;
  assign new_P2_R1209_U180 = ~new_P2_R1209_U66;
  assign new_P2_R1209_U181 = new_P2_U3479 | P2_REG1_REG_17_;
  assign new_P2_R1209_U182 = new_P2_U3476 | P2_REG1_REG_16_;
  assign new_P2_R1209_U183 = ~new_P2_R1209_U47;
  assign new_P2_R1209_U184 = ~new_P2_R1209_U48 | ~new_P2_R1209_U47;
  assign new_P2_R1209_U185 = ~new_P2_U3479 | ~new_P2_R1209_U184;
  assign new_P2_R1209_U186 = ~P2_REG1_REG_17_ | ~new_P2_R1209_U183;
  assign new_P2_R1209_U187 = ~new_P2_R1209_U9 | ~new_P2_R1209_U66;
  assign new_P2_R1209_U188 = ~new_P2_R1209_U65;
  assign new_P2_R1209_U189 = P2_REG1_REG_18_ | new_P2_U3482;
  assign new_P2_R1209_U190 = ~new_P2_R1209_U189 | ~new_P2_R1209_U65;
  assign new_P2_R1209_U191 = ~new_P2_U3482 | ~P2_REG1_REG_18_;
  assign new_P2_R1209_U192 = ~new_P2_R1209_U190 | ~new_P2_R1209_U191 | ~new_P2_R1209_U261 | ~new_P2_R1209_U260;
  assign new_P2_R1209_U193 = ~new_P2_U3482 | ~P2_REG1_REG_18_;
  assign new_P2_R1209_U194 = ~new_P2_R1209_U188 | ~new_P2_R1209_U193;
  assign new_P2_R1209_U195 = new_P2_U3482 | P2_REG1_REG_18_;
  assign new_P2_R1209_U196 = ~new_P2_R1209_U194 | ~new_P2_R1209_U195 | ~new_P2_R1209_U264;
  assign new_P2_R1209_U197 = P2_REG1_REG_16_ | new_P2_U3476;
  assign new_P2_R1209_U198 = ~new_P2_R1209_U197 | ~new_P2_R1209_U66;
  assign new_P2_R1209_U199 = ~new_P2_R1209_U198 | ~new_P2_R1209_U47 | ~new_P2_R1209_U273 | ~new_P2_R1209_U272;
  assign new_P2_R1209_U200 = ~new_P2_R1209_U180 | ~new_P2_R1209_U47;
  assign new_P2_R1209_U201 = ~P2_REG1_REG_17_ | ~new_P2_U3479;
  assign new_P2_R1209_U202 = ~new_P2_R1209_U200 | ~new_P2_R1209_U201 | ~new_P2_R1209_U9;
  assign new_P2_R1209_U203 = new_P2_U3476 | P2_REG1_REG_16_;
  assign new_P2_R1209_U204 = ~new_P2_R1209_U168 | ~new_P2_R1209_U88;
  assign new_P2_R1209_U205 = ~new_P2_R1209_U67;
  assign new_P2_R1209_U206 = P2_REG1_REG_12_ | new_P2_U3464;
  assign new_P2_R1209_U207 = ~new_P2_R1209_U206 | ~new_P2_R1209_U67;
  assign new_P2_R1209_U208 = ~new_P2_R1209_U207 | ~new_P2_R1209_U91 | ~new_P2_R1209_U294 | ~new_P2_R1209_U293;
  assign new_P2_R1209_U209 = ~new_P2_R1209_U205 | ~new_P2_R1209_U91;
  assign new_P2_R1209_U210 = ~new_P2_U3467 | ~P2_REG1_REG_13_;
  assign new_P2_R1209_U211 = ~new_P2_R1209_U209 | ~new_P2_R1209_U210 | ~new_P2_R1209_U8;
  assign new_P2_R1209_U212 = new_P2_U3464 | P2_REG1_REG_12_;
  assign new_P2_R1209_U213 = P2_REG1_REG_9_ | new_P2_U3455;
  assign new_P2_R1209_U214 = ~new_P2_R1209_U213 | ~new_P2_R1209_U38;
  assign new_P2_R1209_U215 = ~new_P2_R1209_U214 | ~new_P2_R1209_U90 | ~new_P2_R1209_U306 | ~new_P2_R1209_U305;
  assign new_P2_R1209_U216 = ~new_P2_R1209_U122 | ~new_P2_R1209_U90;
  assign new_P2_R1209_U217 = ~new_P2_U3458 | ~P2_REG1_REG_10_;
  assign new_P2_R1209_U218 = ~new_P2_R1209_U216 | ~new_P2_R1209_U217 | ~new_P2_R1209_U7;
  assign new_P2_R1209_U219 = ~new_P2_R1209_U123 | ~new_P2_R1209_U90;
  assign new_P2_R1209_U220 = ~new_P2_R1209_U120 | ~new_P2_R1209_U49;
  assign new_P2_R1209_U221 = ~new_P2_R1209_U130 | ~new_P2_R1209_U20;
  assign new_P2_R1209_U222 = ~new_P2_R1209_U144 | ~new_P2_R1209_U32;
  assign new_P2_R1209_U223 = ~new_P2_R1209_U147 | ~new_P2_R1209_U96;
  assign new_P2_R1209_U224 = ~new_P2_R1209_U203 | ~new_P2_R1209_U47;
  assign new_P2_R1209_U225 = ~new_P2_R1209_U212 | ~new_P2_R1209_U91;
  assign new_P2_R1209_U226 = ~new_P2_R1209_U168 | ~new_P2_R1209_U56;
  assign new_P2_R1209_U227 = ~new_P2_U3455 | ~new_P2_R1209_U37;
  assign new_P2_R1209_U228 = ~P2_REG1_REG_9_ | ~new_P2_R1209_U36;
  assign new_P2_R1209_U229 = ~new_P2_R1209_U228 | ~new_P2_R1209_U227;
  assign new_P2_R1209_U230 = ~new_P2_R1209_U219 | ~new_P2_R1209_U38;
  assign new_P2_R1209_U231 = ~new_P2_R1209_U229 | ~new_P2_R1209_U122;
  assign new_P2_R1209_U232 = ~new_P2_U3452 | ~new_P2_R1209_U34;
  assign new_P2_R1209_U233 = ~P2_REG1_REG_8_ | ~new_P2_R1209_U35;
  assign new_P2_R1209_U234 = ~new_P2_R1209_U233 | ~new_P2_R1209_U232;
  assign new_P2_R1209_U235 = ~new_P2_R1209_U220 | ~new_P2_R1209_U81;
  assign new_P2_R1209_U236 = ~new_P2_R1209_U119 | ~new_P2_R1209_U234;
  assign new_P2_R1209_U237 = ~new_P2_U3449 | ~new_P2_R1209_U21;
  assign new_P2_R1209_U238 = ~P2_REG1_REG_7_ | ~new_P2_R1209_U19;
  assign new_P2_R1209_U239 = ~new_P2_U3446 | ~new_P2_R1209_U17;
  assign new_P2_R1209_U240 = ~P2_REG1_REG_6_ | ~new_P2_R1209_U18;
  assign new_P2_R1209_U241 = ~new_P2_R1209_U240 | ~new_P2_R1209_U239;
  assign new_P2_R1209_U242 = ~new_P2_R1209_U221 | ~new_P2_R1209_U39;
  assign new_P2_R1209_U243 = ~new_P2_R1209_U241 | ~new_P2_R1209_U111;
  assign new_P2_R1209_U244 = ~new_P2_U3443 | ~new_P2_R1209_U33;
  assign new_P2_R1209_U245 = ~P2_REG1_REG_5_ | ~new_P2_R1209_U24;
  assign new_P2_R1209_U246 = ~new_P2_U3440 | ~new_P2_R1209_U22;
  assign new_P2_R1209_U247 = ~P2_REG1_REG_4_ | ~new_P2_R1209_U23;
  assign new_P2_R1209_U248 = ~new_P2_R1209_U247 | ~new_P2_R1209_U246;
  assign new_P2_R1209_U249 = ~new_P2_R1209_U222 | ~new_P2_R1209_U42;
  assign new_P2_R1209_U250 = ~new_P2_R1209_U248 | ~new_P2_R1209_U137;
  assign new_P2_R1209_U251 = ~new_P2_U3437 | ~new_P2_R1209_U30;
  assign new_P2_R1209_U252 = ~P2_REG1_REG_3_ | ~new_P2_R1209_U31;
  assign new_P2_R1209_U253 = ~new_P2_R1209_U252 | ~new_P2_R1209_U251;
  assign new_P2_R1209_U254 = ~new_P2_R1209_U223 | ~new_P2_R1209_U82;
  assign new_P2_R1209_U255 = ~new_P2_R1209_U146 | ~new_P2_R1209_U253;
  assign new_P2_R1209_U256 = ~new_P2_U3434 | ~new_P2_R1209_U25;
  assign new_P2_R1209_U257 = ~P2_REG1_REG_2_ | ~new_P2_R1209_U26;
  assign new_P2_R1209_U258 = ~new_P2_R1209_U98 | ~new_P2_R1209_U83;
  assign new_P2_R1209_U259 = ~new_P2_R1209_U153 | ~new_P2_R1209_U29;
  assign new_P2_R1209_U260 = ~new_P2_U3424 | ~new_P2_R1209_U85;
  assign new_P2_R1209_U261 = ~P2_REG1_REG_19_ | ~new_P2_R1209_U84;
  assign new_P2_R1209_U262 = ~new_P2_U3424 | ~new_P2_R1209_U85;
  assign new_P2_R1209_U263 = ~P2_REG1_REG_19_ | ~new_P2_R1209_U84;
  assign new_P2_R1209_U264 = ~new_P2_R1209_U263 | ~new_P2_R1209_U262;
  assign new_P2_R1209_U265 = ~new_P2_U3482 | ~new_P2_R1209_U63;
  assign new_P2_R1209_U266 = ~P2_REG1_REG_18_ | ~new_P2_R1209_U64;
  assign new_P2_R1209_U267 = ~new_P2_U3482 | ~new_P2_R1209_U63;
  assign new_P2_R1209_U268 = ~P2_REG1_REG_18_ | ~new_P2_R1209_U64;
  assign new_P2_R1209_U269 = ~new_P2_R1209_U268 | ~new_P2_R1209_U267;
  assign new_P2_R1209_U270 = ~new_P2_R1209_U65 | ~new_P2_R1209_U266 | ~new_P2_R1209_U265;
  assign new_P2_R1209_U271 = ~new_P2_R1209_U269 | ~new_P2_R1209_U188;
  assign new_P2_R1209_U272 = ~new_P2_U3479 | ~new_P2_R1209_U48;
  assign new_P2_R1209_U273 = ~P2_REG1_REG_17_ | ~new_P2_R1209_U46;
  assign new_P2_R1209_U274 = ~new_P2_U3476 | ~new_P2_R1209_U44;
  assign new_P2_R1209_U275 = ~P2_REG1_REG_16_ | ~new_P2_R1209_U45;
  assign new_P2_R1209_U276 = ~new_P2_R1209_U275 | ~new_P2_R1209_U274;
  assign new_P2_R1209_U277 = ~new_P2_R1209_U224 | ~new_P2_R1209_U66;
  assign new_P2_R1209_U278 = ~new_P2_R1209_U276 | ~new_P2_R1209_U180;
  assign new_P2_R1209_U279 = ~new_P2_U3473 | ~new_P2_R1209_U61;
  assign new_P2_R1209_U280 = ~P2_REG1_REG_15_ | ~new_P2_R1209_U62;
  assign new_P2_R1209_U281 = ~new_P2_U3473 | ~new_P2_R1209_U61;
  assign new_P2_R1209_U282 = ~P2_REG1_REG_15_ | ~new_P2_R1209_U62;
  assign new_P2_R1209_U283 = ~new_P2_R1209_U282 | ~new_P2_R1209_U281;
  assign new_P2_R1209_U284 = ~new_P2_R1209_U86 | ~new_P2_R1209_U280 | ~new_P2_R1209_U279;
  assign new_P2_R1209_U285 = ~new_P2_R1209_U176 | ~new_P2_R1209_U283;
  assign new_P2_R1209_U286 = ~new_P2_U3470 | ~new_P2_R1209_U59;
  assign new_P2_R1209_U287 = ~P2_REG1_REG_14_ | ~new_P2_R1209_U60;
  assign new_P2_R1209_U288 = ~new_P2_U3470 | ~new_P2_R1209_U59;
  assign new_P2_R1209_U289 = ~P2_REG1_REG_14_ | ~new_P2_R1209_U60;
  assign new_P2_R1209_U290 = ~new_P2_R1209_U289 | ~new_P2_R1209_U288;
  assign new_P2_R1209_U291 = ~new_P2_R1209_U87 | ~new_P2_R1209_U287 | ~new_P2_R1209_U286;
  assign new_P2_R1209_U292 = ~new_P2_R1209_U172 | ~new_P2_R1209_U290;
  assign new_P2_R1209_U293 = ~new_P2_U3467 | ~new_P2_R1209_U57;
  assign new_P2_R1209_U294 = ~P2_REG1_REG_13_ | ~new_P2_R1209_U58;
  assign new_P2_R1209_U295 = ~new_P2_U3464 | ~new_P2_R1209_U52;
  assign new_P2_R1209_U296 = ~P2_REG1_REG_12_ | ~new_P2_R1209_U53;
  assign new_P2_R1209_U297 = ~new_P2_R1209_U296 | ~new_P2_R1209_U295;
  assign new_P2_R1209_U298 = ~new_P2_R1209_U225 | ~new_P2_R1209_U67;
  assign new_P2_R1209_U299 = ~new_P2_R1209_U297 | ~new_P2_R1209_U205;
  assign new_P2_R1209_U300 = ~new_P2_U3461 | ~new_P2_R1209_U54;
  assign new_P2_R1209_U301 = ~P2_REG1_REG_11_ | ~new_P2_R1209_U55;
  assign new_P2_R1209_U302 = ~new_P2_R1209_U301 | ~new_P2_R1209_U300;
  assign new_P2_R1209_U303 = ~new_P2_R1209_U226 | ~new_P2_R1209_U88;
  assign new_P2_R1209_U304 = ~new_P2_R1209_U162 | ~new_P2_R1209_U302;
  assign new_P2_R1209_U305 = ~new_P2_U3458 | ~new_P2_R1209_U50;
  assign new_P2_R1209_U306 = ~P2_REG1_REG_10_ | ~new_P2_R1209_U51;
  assign new_P2_R1209_U307 = ~new_P2_U3425 | ~new_P2_R1209_U27;
  assign new_P2_R1209_U308 = ~P2_REG1_REG_0_ | ~new_P2_R1209_U28;
  assign new_P2_R1170_U4 = new_P2_R1170_U95 & new_P2_R1170_U94;
  assign new_P2_R1170_U5 = new_P2_R1170_U96 & new_P2_R1170_U97;
  assign new_P2_R1170_U6 = new_P2_R1170_U113 & new_P2_R1170_U112;
  assign new_P2_R1170_U7 = new_P2_R1170_U155 & new_P2_R1170_U154;
  assign new_P2_R1170_U8 = new_P2_R1170_U164 & new_P2_R1170_U163;
  assign new_P2_R1170_U9 = new_P2_R1170_U182 & new_P2_R1170_U181;
  assign new_P2_R1170_U10 = new_P2_R1170_U218 & new_P2_R1170_U215;
  assign new_P2_R1170_U11 = new_P2_R1170_U211 & new_P2_R1170_U208;
  assign new_P2_R1170_U12 = new_P2_R1170_U202 & new_P2_R1170_U199;
  assign new_P2_R1170_U13 = new_P2_R1170_U196 & new_P2_R1170_U192;
  assign new_P2_R1170_U14 = new_P2_R1170_U151 & new_P2_R1170_U148;
  assign new_P2_R1170_U15 = new_P2_R1170_U143 & new_P2_R1170_U140;
  assign new_P2_R1170_U16 = new_P2_R1170_U129 & new_P2_R1170_U126;
  assign new_P2_R1170_U17 = ~P2_REG2_REG_6_;
  assign new_P2_R1170_U18 = ~new_P2_U3446;
  assign new_P2_R1170_U19 = ~new_P2_U3449;
  assign new_P2_R1170_U20 = ~new_P2_U3446 | ~P2_REG2_REG_6_;
  assign new_P2_R1170_U21 = ~P2_REG2_REG_7_;
  assign new_P2_R1170_U22 = ~P2_REG2_REG_4_;
  assign new_P2_R1170_U23 = ~new_P2_U3440;
  assign new_P2_R1170_U24 = ~new_P2_U3443;
  assign new_P2_R1170_U25 = ~P2_REG2_REG_2_;
  assign new_P2_R1170_U26 = ~new_P2_U3434;
  assign new_P2_R1170_U27 = ~P2_REG2_REG_0_;
  assign new_P2_R1170_U28 = ~new_P2_U3425;
  assign new_P2_R1170_U29 = ~new_P2_U3425 | ~P2_REG2_REG_0_;
  assign new_P2_R1170_U30 = ~P2_REG2_REG_3_;
  assign new_P2_R1170_U31 = ~new_P2_U3437;
  assign new_P2_R1170_U32 = ~new_P2_U3440 | ~P2_REG2_REG_4_;
  assign new_P2_R1170_U33 = ~P2_REG2_REG_5_;
  assign new_P2_R1170_U34 = ~P2_REG2_REG_8_;
  assign new_P2_R1170_U35 = ~new_P2_U3452;
  assign new_P2_R1170_U36 = ~new_P2_U3455;
  assign new_P2_R1170_U37 = ~P2_REG2_REG_9_;
  assign new_P2_R1170_U38 = ~new_P2_R1170_U49 | ~new_P2_R1170_U121;
  assign new_P2_R1170_U39 = ~new_P2_R1170_U109 | ~new_P2_R1170_U110 | ~new_P2_R1170_U108;
  assign new_P2_R1170_U40 = ~new_P2_R1170_U98 | ~new_P2_R1170_U99;
  assign new_P2_R1170_U41 = ~P2_REG2_REG_1_ | ~new_P2_U3431;
  assign new_P2_R1170_U42 = ~new_P2_R1170_U135 | ~new_P2_R1170_U136 | ~new_P2_R1170_U134;
  assign new_P2_R1170_U43 = ~new_P2_R1170_U132 | ~new_P2_R1170_U131;
  assign new_P2_R1170_U44 = ~P2_REG2_REG_16_;
  assign new_P2_R1170_U45 = ~new_P2_U3476;
  assign new_P2_R1170_U46 = ~new_P2_U3479;
  assign new_P2_R1170_U47 = ~new_P2_U3476 | ~P2_REG2_REG_16_;
  assign new_P2_R1170_U48 = ~P2_REG2_REG_17_;
  assign new_P2_R1170_U49 = ~new_P2_U3452 | ~P2_REG2_REG_8_;
  assign new_P2_R1170_U50 = ~P2_REG2_REG_10_;
  assign new_P2_R1170_U51 = ~new_P2_U3458;
  assign new_P2_R1170_U52 = ~P2_REG2_REG_12_;
  assign new_P2_R1170_U53 = ~new_P2_U3464;
  assign new_P2_R1170_U54 = ~P2_REG2_REG_11_;
  assign new_P2_R1170_U55 = ~new_P2_U3461;
  assign new_P2_R1170_U56 = ~new_P2_U3461 | ~P2_REG2_REG_11_;
  assign new_P2_R1170_U57 = ~P2_REG2_REG_13_;
  assign new_P2_R1170_U58 = ~new_P2_U3467;
  assign new_P2_R1170_U59 = ~P2_REG2_REG_14_;
  assign new_P2_R1170_U60 = ~new_P2_U3470;
  assign new_P2_R1170_U61 = ~P2_REG2_REG_15_;
  assign new_P2_R1170_U62 = ~new_P2_U3473;
  assign new_P2_R1170_U63 = ~P2_REG2_REG_18_;
  assign new_P2_R1170_U64 = ~new_P2_U3482;
  assign new_P2_R1170_U65 = ~new_P2_R1170_U187 | ~new_P2_R1170_U186 | ~new_P2_R1170_U185;
  assign new_P2_R1170_U66 = ~new_P2_R1170_U179 | ~new_P2_R1170_U178;
  assign new_P2_R1170_U67 = ~new_P2_R1170_U56 | ~new_P2_R1170_U204;
  assign new_P2_R1170_U68 = ~new_P2_R1170_U259 | ~new_P2_R1170_U258;
  assign new_P2_R1170_U69 = ~new_P2_R1170_U308 | ~new_P2_R1170_U307;
  assign new_P2_R1170_U70 = ~new_P2_R1170_U231 | ~new_P2_R1170_U230;
  assign new_P2_R1170_U71 = ~new_P2_R1170_U236 | ~new_P2_R1170_U235;
  assign new_P2_R1170_U72 = ~new_P2_R1170_U243 | ~new_P2_R1170_U242;
  assign new_P2_R1170_U73 = ~new_P2_R1170_U250 | ~new_P2_R1170_U249;
  assign new_P2_R1170_U74 = ~new_P2_R1170_U255 | ~new_P2_R1170_U254;
  assign new_P2_R1170_U75 = ~new_P2_R1170_U271 | ~new_P2_R1170_U270;
  assign new_P2_R1170_U76 = ~new_P2_R1170_U278 | ~new_P2_R1170_U277;
  assign new_P2_R1170_U77 = ~new_P2_R1170_U285 | ~new_P2_R1170_U284;
  assign new_P2_R1170_U78 = ~new_P2_R1170_U292 | ~new_P2_R1170_U291;
  assign new_P2_R1170_U79 = ~new_P2_R1170_U299 | ~new_P2_R1170_U298;
  assign new_P2_R1170_U80 = ~new_P2_R1170_U304 | ~new_P2_R1170_U303;
  assign new_P2_R1170_U81 = ~new_P2_R1170_U118 | ~new_P2_R1170_U117 | ~new_P2_R1170_U116;
  assign new_P2_R1170_U82 = ~new_P2_R1170_U133 | ~new_P2_R1170_U145;
  assign new_P2_R1170_U83 = ~new_P2_R1170_U41 | ~new_P2_R1170_U152;
  assign new_P2_R1170_U84 = ~new_P2_U3424;
  assign new_P2_R1170_U85 = ~P2_REG2_REG_19_;
  assign new_P2_R1170_U86 = ~new_P2_R1170_U175 | ~new_P2_R1170_U174;
  assign new_P2_R1170_U87 = ~new_P2_R1170_U171 | ~new_P2_R1170_U170;
  assign new_P2_R1170_U88 = ~new_P2_R1170_U161 | ~new_P2_R1170_U160;
  assign new_P2_R1170_U89 = ~new_P2_R1170_U32;
  assign new_P2_R1170_U90 = ~P2_REG2_REG_9_ | ~new_P2_U3455;
  assign new_P2_R1170_U91 = ~new_P2_U3464 | ~P2_REG2_REG_12_;
  assign new_P2_R1170_U92 = ~new_P2_R1170_U56;
  assign new_P2_R1170_U93 = ~new_P2_R1170_U49;
  assign new_P2_R1170_U94 = new_P2_U3443 | P2_REG2_REG_5_;
  assign new_P2_R1170_U95 = new_P2_U3440 | P2_REG2_REG_4_;
  assign new_P2_R1170_U96 = P2_REG2_REG_3_ | new_P2_U3437;
  assign new_P2_R1170_U97 = P2_REG2_REG_2_ | new_P2_U3434;
  assign new_P2_R1170_U98 = ~new_P2_R1170_U29;
  assign new_P2_R1170_U99 = P2_REG2_REG_1_ | new_P2_U3431;
  assign new_P2_R1170_U100 = ~new_P2_R1170_U40;
  assign new_P2_R1170_U101 = ~new_P2_R1170_U41;
  assign new_P2_R1170_U102 = ~new_P2_R1170_U40 | ~new_P2_R1170_U41;
  assign new_P2_R1170_U103 = ~new_P2_R1170_U96 | ~P2_REG2_REG_2_ | ~new_P2_U3434;
  assign new_P2_R1170_U104 = ~new_P2_R1170_U5 | ~new_P2_R1170_U102;
  assign new_P2_R1170_U105 = ~new_P2_U3437 | ~P2_REG2_REG_3_;
  assign new_P2_R1170_U106 = ~new_P2_R1170_U104 | ~new_P2_R1170_U105 | ~new_P2_R1170_U103;
  assign new_P2_R1170_U107 = ~new_P2_R1170_U33 | ~new_P2_R1170_U32;
  assign new_P2_R1170_U108 = ~new_P2_U3443 | ~new_P2_R1170_U107;
  assign new_P2_R1170_U109 = ~new_P2_R1170_U4 | ~new_P2_R1170_U106;
  assign new_P2_R1170_U110 = ~P2_REG2_REG_5_ | ~new_P2_R1170_U89;
  assign new_P2_R1170_U111 = ~new_P2_R1170_U39;
  assign new_P2_R1170_U112 = new_P2_U3449 | P2_REG2_REG_7_;
  assign new_P2_R1170_U113 = new_P2_U3446 | P2_REG2_REG_6_;
  assign new_P2_R1170_U114 = ~new_P2_R1170_U20;
  assign new_P2_R1170_U115 = ~new_P2_R1170_U21 | ~new_P2_R1170_U20;
  assign new_P2_R1170_U116 = ~new_P2_U3449 | ~new_P2_R1170_U115;
  assign new_P2_R1170_U117 = ~P2_REG2_REG_7_ | ~new_P2_R1170_U114;
  assign new_P2_R1170_U118 = ~new_P2_R1170_U6 | ~new_P2_R1170_U39;
  assign new_P2_R1170_U119 = ~new_P2_R1170_U81;
  assign new_P2_R1170_U120 = P2_REG2_REG_8_ | new_P2_U3452;
  assign new_P2_R1170_U121 = ~new_P2_R1170_U120 | ~new_P2_R1170_U81;
  assign new_P2_R1170_U122 = ~new_P2_R1170_U38;
  assign new_P2_R1170_U123 = new_P2_U3455 | P2_REG2_REG_9_;
  assign new_P2_R1170_U124 = P2_REG2_REG_6_ | new_P2_U3446;
  assign new_P2_R1170_U125 = ~new_P2_R1170_U124 | ~new_P2_R1170_U39;
  assign new_P2_R1170_U126 = ~new_P2_R1170_U125 | ~new_P2_R1170_U20 | ~new_P2_R1170_U238 | ~new_P2_R1170_U237;
  assign new_P2_R1170_U127 = ~new_P2_R1170_U111 | ~new_P2_R1170_U20;
  assign new_P2_R1170_U128 = ~P2_REG2_REG_7_ | ~new_P2_U3449;
  assign new_P2_R1170_U129 = ~new_P2_R1170_U127 | ~new_P2_R1170_U128 | ~new_P2_R1170_U6;
  assign new_P2_R1170_U130 = new_P2_U3446 | P2_REG2_REG_6_;
  assign new_P2_R1170_U131 = ~new_P2_R1170_U101 | ~new_P2_R1170_U97;
  assign new_P2_R1170_U132 = ~new_P2_U3434 | ~P2_REG2_REG_2_;
  assign new_P2_R1170_U133 = ~new_P2_R1170_U43;
  assign new_P2_R1170_U134 = ~new_P2_R1170_U100 | ~new_P2_R1170_U5;
  assign new_P2_R1170_U135 = ~new_P2_R1170_U43 | ~new_P2_R1170_U96;
  assign new_P2_R1170_U136 = ~new_P2_U3437 | ~P2_REG2_REG_3_;
  assign new_P2_R1170_U137 = ~new_P2_R1170_U42;
  assign new_P2_R1170_U138 = P2_REG2_REG_4_ | new_P2_U3440;
  assign new_P2_R1170_U139 = ~new_P2_R1170_U138 | ~new_P2_R1170_U42;
  assign new_P2_R1170_U140 = ~new_P2_R1170_U139 | ~new_P2_R1170_U32 | ~new_P2_R1170_U245 | ~new_P2_R1170_U244;
  assign new_P2_R1170_U141 = ~new_P2_R1170_U137 | ~new_P2_R1170_U32;
  assign new_P2_R1170_U142 = ~P2_REG2_REG_5_ | ~new_P2_U3443;
  assign new_P2_R1170_U143 = ~new_P2_R1170_U141 | ~new_P2_R1170_U142 | ~new_P2_R1170_U4;
  assign new_P2_R1170_U144 = new_P2_U3440 | P2_REG2_REG_4_;
  assign new_P2_R1170_U145 = ~new_P2_R1170_U100 | ~new_P2_R1170_U97;
  assign new_P2_R1170_U146 = ~new_P2_R1170_U82;
  assign new_P2_R1170_U147 = ~new_P2_U3437 | ~P2_REG2_REG_3_;
  assign new_P2_R1170_U148 = ~new_P2_R1170_U40 | ~new_P2_R1170_U41 | ~new_P2_R1170_U257 | ~new_P2_R1170_U256;
  assign new_P2_R1170_U149 = ~new_P2_R1170_U41 | ~new_P2_R1170_U40;
  assign new_P2_R1170_U150 = ~new_P2_U3434 | ~P2_REG2_REG_2_;
  assign new_P2_R1170_U151 = ~new_P2_R1170_U149 | ~new_P2_R1170_U150 | ~new_P2_R1170_U97;
  assign new_P2_R1170_U152 = P2_REG2_REG_1_ | new_P2_U3431;
  assign new_P2_R1170_U153 = ~new_P2_R1170_U83;
  assign new_P2_R1170_U154 = new_P2_U3455 | P2_REG2_REG_9_;
  assign new_P2_R1170_U155 = new_P2_U3458 | P2_REG2_REG_10_;
  assign new_P2_R1170_U156 = ~new_P2_R1170_U93 | ~new_P2_R1170_U7;
  assign new_P2_R1170_U157 = ~new_P2_U3458 | ~P2_REG2_REG_10_;
  assign new_P2_R1170_U158 = ~new_P2_R1170_U156 | ~new_P2_R1170_U157 | ~new_P2_R1170_U90;
  assign new_P2_R1170_U159 = P2_REG2_REG_10_ | new_P2_U3458;
  assign new_P2_R1170_U160 = ~new_P2_R1170_U81 | ~new_P2_R1170_U120 | ~new_P2_R1170_U7;
  assign new_P2_R1170_U161 = ~new_P2_R1170_U159 | ~new_P2_R1170_U158;
  assign new_P2_R1170_U162 = ~new_P2_R1170_U88;
  assign new_P2_R1170_U163 = new_P2_U3467 | P2_REG2_REG_13_;
  assign new_P2_R1170_U164 = new_P2_U3464 | P2_REG2_REG_12_;
  assign new_P2_R1170_U165 = ~new_P2_R1170_U92 | ~new_P2_R1170_U8;
  assign new_P2_R1170_U166 = ~new_P2_U3467 | ~P2_REG2_REG_13_;
  assign new_P2_R1170_U167 = ~new_P2_R1170_U165 | ~new_P2_R1170_U166 | ~new_P2_R1170_U91;
  assign new_P2_R1170_U168 = P2_REG2_REG_11_ | new_P2_U3461;
  assign new_P2_R1170_U169 = P2_REG2_REG_13_ | new_P2_U3467;
  assign new_P2_R1170_U170 = ~new_P2_R1170_U88 | ~new_P2_R1170_U168 | ~new_P2_R1170_U8;
  assign new_P2_R1170_U171 = ~new_P2_R1170_U169 | ~new_P2_R1170_U167;
  assign new_P2_R1170_U172 = ~new_P2_R1170_U87;
  assign new_P2_R1170_U173 = P2_REG2_REG_14_ | new_P2_U3470;
  assign new_P2_R1170_U174 = ~new_P2_R1170_U173 | ~new_P2_R1170_U87;
  assign new_P2_R1170_U175 = ~new_P2_U3470 | ~P2_REG2_REG_14_;
  assign new_P2_R1170_U176 = ~new_P2_R1170_U86;
  assign new_P2_R1170_U177 = P2_REG2_REG_15_ | new_P2_U3473;
  assign new_P2_R1170_U178 = ~new_P2_R1170_U177 | ~new_P2_R1170_U86;
  assign new_P2_R1170_U179 = ~new_P2_U3473 | ~P2_REG2_REG_15_;
  assign new_P2_R1170_U180 = ~new_P2_R1170_U66;
  assign new_P2_R1170_U181 = new_P2_U3479 | P2_REG2_REG_17_;
  assign new_P2_R1170_U182 = new_P2_U3476 | P2_REG2_REG_16_;
  assign new_P2_R1170_U183 = ~new_P2_R1170_U47;
  assign new_P2_R1170_U184 = ~new_P2_R1170_U48 | ~new_P2_R1170_U47;
  assign new_P2_R1170_U185 = ~new_P2_U3479 | ~new_P2_R1170_U184;
  assign new_P2_R1170_U186 = ~P2_REG2_REG_17_ | ~new_P2_R1170_U183;
  assign new_P2_R1170_U187 = ~new_P2_R1170_U9 | ~new_P2_R1170_U66;
  assign new_P2_R1170_U188 = ~new_P2_R1170_U65;
  assign new_P2_R1170_U189 = P2_REG2_REG_18_ | new_P2_U3482;
  assign new_P2_R1170_U190 = ~new_P2_R1170_U189 | ~new_P2_R1170_U65;
  assign new_P2_R1170_U191 = ~new_P2_U3482 | ~P2_REG2_REG_18_;
  assign new_P2_R1170_U192 = ~new_P2_R1170_U190 | ~new_P2_R1170_U191 | ~new_P2_R1170_U261 | ~new_P2_R1170_U260;
  assign new_P2_R1170_U193 = ~new_P2_U3482 | ~P2_REG2_REG_18_;
  assign new_P2_R1170_U194 = ~new_P2_R1170_U188 | ~new_P2_R1170_U193;
  assign new_P2_R1170_U195 = new_P2_U3482 | P2_REG2_REG_18_;
  assign new_P2_R1170_U196 = ~new_P2_R1170_U194 | ~new_P2_R1170_U195 | ~new_P2_R1170_U264;
  assign new_P2_R1170_U197 = P2_REG2_REG_16_ | new_P2_U3476;
  assign new_P2_R1170_U198 = ~new_P2_R1170_U197 | ~new_P2_R1170_U66;
  assign new_P2_R1170_U199 = ~new_P2_R1170_U198 | ~new_P2_R1170_U47 | ~new_P2_R1170_U273 | ~new_P2_R1170_U272;
  assign new_P2_R1170_U200 = ~new_P2_R1170_U180 | ~new_P2_R1170_U47;
  assign new_P2_R1170_U201 = ~P2_REG2_REG_17_ | ~new_P2_U3479;
  assign new_P2_R1170_U202 = ~new_P2_R1170_U200 | ~new_P2_R1170_U201 | ~new_P2_R1170_U9;
  assign new_P2_R1170_U203 = new_P2_U3476 | P2_REG2_REG_16_;
  assign new_P2_R1170_U204 = ~new_P2_R1170_U168 | ~new_P2_R1170_U88;
  assign new_P2_R1170_U205 = ~new_P2_R1170_U67;
  assign new_P2_R1170_U206 = P2_REG2_REG_12_ | new_P2_U3464;
  assign new_P2_R1170_U207 = ~new_P2_R1170_U206 | ~new_P2_R1170_U67;
  assign new_P2_R1170_U208 = ~new_P2_R1170_U207 | ~new_P2_R1170_U91 | ~new_P2_R1170_U294 | ~new_P2_R1170_U293;
  assign new_P2_R1170_U209 = ~new_P2_R1170_U205 | ~new_P2_R1170_U91;
  assign new_P2_R1170_U210 = ~new_P2_U3467 | ~P2_REG2_REG_13_;
  assign new_P2_R1170_U211 = ~new_P2_R1170_U209 | ~new_P2_R1170_U210 | ~new_P2_R1170_U8;
  assign new_P2_R1170_U212 = new_P2_U3464 | P2_REG2_REG_12_;
  assign new_P2_R1170_U213 = P2_REG2_REG_9_ | new_P2_U3455;
  assign new_P2_R1170_U214 = ~new_P2_R1170_U213 | ~new_P2_R1170_U38;
  assign new_P2_R1170_U215 = ~new_P2_R1170_U214 | ~new_P2_R1170_U90 | ~new_P2_R1170_U306 | ~new_P2_R1170_U305;
  assign new_P2_R1170_U216 = ~new_P2_R1170_U122 | ~new_P2_R1170_U90;
  assign new_P2_R1170_U217 = ~new_P2_U3458 | ~P2_REG2_REG_10_;
  assign new_P2_R1170_U218 = ~new_P2_R1170_U216 | ~new_P2_R1170_U217 | ~new_P2_R1170_U7;
  assign new_P2_R1170_U219 = ~new_P2_R1170_U123 | ~new_P2_R1170_U90;
  assign new_P2_R1170_U220 = ~new_P2_R1170_U120 | ~new_P2_R1170_U49;
  assign new_P2_R1170_U221 = ~new_P2_R1170_U130 | ~new_P2_R1170_U20;
  assign new_P2_R1170_U222 = ~new_P2_R1170_U144 | ~new_P2_R1170_U32;
  assign new_P2_R1170_U223 = ~new_P2_R1170_U147 | ~new_P2_R1170_U96;
  assign new_P2_R1170_U224 = ~new_P2_R1170_U203 | ~new_P2_R1170_U47;
  assign new_P2_R1170_U225 = ~new_P2_R1170_U212 | ~new_P2_R1170_U91;
  assign new_P2_R1170_U226 = ~new_P2_R1170_U168 | ~new_P2_R1170_U56;
  assign new_P2_R1170_U227 = ~new_P2_U3455 | ~new_P2_R1170_U37;
  assign new_P2_R1170_U228 = ~P2_REG2_REG_9_ | ~new_P2_R1170_U36;
  assign new_P2_R1170_U229 = ~new_P2_R1170_U228 | ~new_P2_R1170_U227;
  assign new_P2_R1170_U230 = ~new_P2_R1170_U219 | ~new_P2_R1170_U38;
  assign new_P2_R1170_U231 = ~new_P2_R1170_U229 | ~new_P2_R1170_U122;
  assign new_P2_R1170_U232 = ~new_P2_U3452 | ~new_P2_R1170_U34;
  assign new_P2_R1170_U233 = ~P2_REG2_REG_8_ | ~new_P2_R1170_U35;
  assign new_P2_R1170_U234 = ~new_P2_R1170_U233 | ~new_P2_R1170_U232;
  assign new_P2_R1170_U235 = ~new_P2_R1170_U220 | ~new_P2_R1170_U81;
  assign new_P2_R1170_U236 = ~new_P2_R1170_U119 | ~new_P2_R1170_U234;
  assign new_P2_R1170_U237 = ~new_P2_U3449 | ~new_P2_R1170_U21;
  assign new_P2_R1170_U238 = ~P2_REG2_REG_7_ | ~new_P2_R1170_U19;
  assign new_P2_R1170_U239 = ~new_P2_U3446 | ~new_P2_R1170_U17;
  assign new_P2_R1170_U240 = ~P2_REG2_REG_6_ | ~new_P2_R1170_U18;
  assign new_P2_R1170_U241 = ~new_P2_R1170_U240 | ~new_P2_R1170_U239;
  assign new_P2_R1170_U242 = ~new_P2_R1170_U221 | ~new_P2_R1170_U39;
  assign new_P2_R1170_U243 = ~new_P2_R1170_U241 | ~new_P2_R1170_U111;
  assign new_P2_R1170_U244 = ~new_P2_U3443 | ~new_P2_R1170_U33;
  assign new_P2_R1170_U245 = ~P2_REG2_REG_5_ | ~new_P2_R1170_U24;
  assign new_P2_R1170_U246 = ~new_P2_U3440 | ~new_P2_R1170_U22;
  assign new_P2_R1170_U247 = ~P2_REG2_REG_4_ | ~new_P2_R1170_U23;
  assign new_P2_R1170_U248 = ~new_P2_R1170_U247 | ~new_P2_R1170_U246;
  assign new_P2_R1170_U249 = ~new_P2_R1170_U222 | ~new_P2_R1170_U42;
  assign new_P2_R1170_U250 = ~new_P2_R1170_U248 | ~new_P2_R1170_U137;
  assign new_P2_R1170_U251 = ~new_P2_U3437 | ~new_P2_R1170_U30;
  assign new_P2_R1170_U252 = ~P2_REG2_REG_3_ | ~new_P2_R1170_U31;
  assign new_P2_R1170_U253 = ~new_P2_R1170_U252 | ~new_P2_R1170_U251;
  assign new_P2_R1170_U254 = ~new_P2_R1170_U223 | ~new_P2_R1170_U82;
  assign new_P2_R1170_U255 = ~new_P2_R1170_U146 | ~new_P2_R1170_U253;
  assign new_P2_R1170_U256 = ~new_P2_U3434 | ~new_P2_R1170_U25;
  assign new_P2_R1170_U257 = ~P2_REG2_REG_2_ | ~new_P2_R1170_U26;
  assign new_P2_R1170_U258 = ~new_P2_R1170_U98 | ~new_P2_R1170_U83;
  assign new_P2_R1170_U259 = ~new_P2_R1170_U153 | ~new_P2_R1170_U29;
  assign new_P2_R1170_U260 = ~new_P2_U3424 | ~new_P2_R1170_U85;
  assign new_P2_R1170_U261 = ~P2_REG2_REG_19_ | ~new_P2_R1170_U84;
  assign new_P2_R1170_U262 = ~new_P2_U3424 | ~new_P2_R1170_U85;
  assign new_P2_R1170_U263 = ~P2_REG2_REG_19_ | ~new_P2_R1170_U84;
  assign new_P2_R1170_U264 = ~new_P2_R1170_U263 | ~new_P2_R1170_U262;
  assign new_P2_R1170_U265 = ~new_P2_U3482 | ~new_P2_R1170_U63;
  assign new_P2_R1170_U266 = ~P2_REG2_REG_18_ | ~new_P2_R1170_U64;
  assign new_P2_R1170_U267 = ~new_P2_U3482 | ~new_P2_R1170_U63;
  assign new_P2_R1170_U268 = ~P2_REG2_REG_18_ | ~new_P2_R1170_U64;
  assign new_P2_R1170_U269 = ~new_P2_R1170_U268 | ~new_P2_R1170_U267;
  assign new_P2_R1170_U270 = ~new_P2_R1170_U65 | ~new_P2_R1170_U266 | ~new_P2_R1170_U265;
  assign new_P2_R1170_U271 = ~new_P2_R1170_U269 | ~new_P2_R1170_U188;
  assign new_P2_R1170_U272 = ~new_P2_U3479 | ~new_P2_R1170_U48;
  assign new_P2_R1170_U273 = ~P2_REG2_REG_17_ | ~new_P2_R1170_U46;
  assign new_P2_R1170_U274 = ~new_P2_U3476 | ~new_P2_R1170_U44;
  assign new_P2_R1170_U275 = ~P2_REG2_REG_16_ | ~new_P2_R1170_U45;
  assign new_P2_R1170_U276 = ~new_P2_R1170_U275 | ~new_P2_R1170_U274;
  assign new_P2_R1170_U277 = ~new_P2_R1170_U224 | ~new_P2_R1170_U66;
  assign new_P2_R1170_U278 = ~new_P2_R1170_U276 | ~new_P2_R1170_U180;
  assign new_P2_R1170_U279 = ~new_P2_U3473 | ~new_P2_R1170_U61;
  assign new_P2_R1170_U280 = ~P2_REG2_REG_15_ | ~new_P2_R1170_U62;
  assign new_P2_R1170_U281 = ~new_P2_U3473 | ~new_P2_R1170_U61;
  assign new_P2_R1170_U282 = ~P2_REG2_REG_15_ | ~new_P2_R1170_U62;
  assign new_P2_R1170_U283 = ~new_P2_R1170_U282 | ~new_P2_R1170_U281;
  assign new_P2_R1170_U284 = ~new_P2_R1170_U86 | ~new_P2_R1170_U280 | ~new_P2_R1170_U279;
  assign new_P2_R1170_U285 = ~new_P2_R1170_U176 | ~new_P2_R1170_U283;
  assign new_P2_R1170_U286 = ~new_P2_U3470 | ~new_P2_R1170_U59;
  assign new_P2_R1170_U287 = ~P2_REG2_REG_14_ | ~new_P2_R1170_U60;
  assign new_P2_R1170_U288 = ~new_P2_U3470 | ~new_P2_R1170_U59;
  assign new_P2_R1170_U289 = ~P2_REG2_REG_14_ | ~new_P2_R1170_U60;
  assign new_P2_R1170_U290 = ~new_P2_R1170_U289 | ~new_P2_R1170_U288;
  assign new_P2_R1170_U291 = ~new_P2_R1170_U87 | ~new_P2_R1170_U287 | ~new_P2_R1170_U286;
  assign new_P2_R1170_U292 = ~new_P2_R1170_U172 | ~new_P2_R1170_U290;
  assign new_P2_R1170_U293 = ~new_P2_U3467 | ~new_P2_R1170_U57;
  assign new_P2_R1170_U294 = ~P2_REG2_REG_13_ | ~new_P2_R1170_U58;
  assign new_P2_R1170_U295 = ~new_P2_U3464 | ~new_P2_R1170_U52;
  assign new_P2_R1170_U296 = ~P2_REG2_REG_12_ | ~new_P2_R1170_U53;
  assign new_P2_R1170_U297 = ~new_P2_R1170_U296 | ~new_P2_R1170_U295;
  assign new_P2_R1170_U298 = ~new_P2_R1170_U225 | ~new_P2_R1170_U67;
  assign new_P2_R1170_U299 = ~new_P2_R1170_U297 | ~new_P2_R1170_U205;
  assign new_P2_R1170_U300 = ~new_P2_U3461 | ~new_P2_R1170_U54;
  assign new_P2_R1170_U301 = ~P2_REG2_REG_11_ | ~new_P2_R1170_U55;
  assign new_P2_R1170_U302 = ~new_P2_R1170_U301 | ~new_P2_R1170_U300;
  assign new_P2_R1170_U303 = ~new_P2_R1170_U226 | ~new_P2_R1170_U88;
  assign new_P2_R1170_U304 = ~new_P2_R1170_U162 | ~new_P2_R1170_U302;
  assign new_P2_R1170_U305 = ~new_P2_U3458 | ~new_P2_R1170_U50;
  assign new_P2_R1170_U306 = ~P2_REG2_REG_10_ | ~new_P2_R1170_U51;
  assign new_P2_R1170_U307 = ~new_P2_U3425 | ~new_P2_R1170_U27;
  assign new_P2_R1170_U308 = ~P2_REG2_REG_0_ | ~new_P2_R1170_U28;
  assign new_P2_R1275_U6 = new_P2_R1275_U135 & new_P2_R1275_U35;
  assign new_P2_R1275_U7 = new_P2_R1275_U133 & new_P2_R1275_U36;
  assign new_P2_R1275_U8 = new_P2_R1275_U132 & new_P2_R1275_U37;
  assign new_P2_R1275_U9 = new_P2_R1275_U131 & new_P2_R1275_U38;
  assign new_P2_R1275_U10 = new_P2_R1275_U129 & new_P2_R1275_U39;
  assign new_P2_R1275_U11 = new_P2_R1275_U128 & new_P2_R1275_U40;
  assign new_P2_R1275_U12 = new_P2_R1275_U127 & new_P2_R1275_U41;
  assign new_P2_R1275_U13 = new_P2_R1275_U125 & new_P2_R1275_U42;
  assign new_P2_R1275_U14 = new_P2_R1275_U123 & new_P2_R1275_U43;
  assign new_P2_R1275_U15 = new_P2_R1275_U121 & new_P2_R1275_U44;
  assign new_P2_R1275_U16 = new_P2_R1275_U119 & new_P2_R1275_U45;
  assign new_P2_R1275_U17 = new_P2_R1275_U117 & new_P2_R1275_U46;
  assign new_P2_R1275_U18 = new_P2_R1275_U115 & new_P2_R1275_U25;
  assign new_P2_R1275_U19 = new_P2_R1275_U113 & new_P2_R1275_U67;
  assign new_P2_R1275_U20 = new_P2_R1275_U98 & new_P2_R1275_U26;
  assign new_P2_R1275_U21 = new_P2_R1275_U97 & new_P2_R1275_U27;
  assign new_P2_R1275_U22 = new_P2_R1275_U96 & new_P2_R1275_U28;
  assign new_P2_R1275_U23 = new_P2_R1275_U94 & new_P2_R1275_U29;
  assign new_P2_R1275_U24 = new_P2_R1275_U93 & new_P2_R1275_U30;
  assign new_P2_R1275_U25 = new_P2_U3435 | new_P2_U3432 | new_P2_U3427;
  assign new_P2_R1275_U26 = ~new_P2_R1275_U87 | ~new_P2_R1275_U34;
  assign new_P2_R1275_U27 = ~new_P2_R1275_U88 | ~new_P2_R1275_U33;
  assign new_P2_R1275_U28 = ~new_P2_R1275_U56 | ~new_P2_R1275_U89;
  assign new_P2_R1275_U29 = ~new_P2_R1275_U90 | ~new_P2_R1275_U32;
  assign new_P2_R1275_U30 = ~new_P2_R1275_U91 | ~new_P2_R1275_U31;
  assign new_P2_R1275_U31 = ~new_P2_U3453;
  assign new_P2_R1275_U32 = ~new_P2_U3450;
  assign new_P2_R1275_U33 = ~new_P2_U3441;
  assign new_P2_R1275_U34 = ~new_P2_U3438;
  assign new_P2_R1275_U35 = ~new_P2_R1275_U57 | ~new_P2_R1275_U92;
  assign new_P2_R1275_U36 = ~new_P2_R1275_U99 | ~new_P2_R1275_U54;
  assign new_P2_R1275_U37 = ~new_P2_R1275_U100 | ~new_P2_R1275_U53;
  assign new_P2_R1275_U38 = ~new_P2_R1275_U58 | ~new_P2_R1275_U101;
  assign new_P2_R1275_U39 = ~new_P2_R1275_U102 | ~new_P2_R1275_U52;
  assign new_P2_R1275_U40 = ~new_P2_R1275_U103 | ~new_P2_R1275_U51;
  assign new_P2_R1275_U41 = ~new_P2_R1275_U59 | ~new_P2_R1275_U104;
  assign new_P2_R1275_U42 = ~new_P2_R1275_U60 | ~new_P2_R1275_U105;
  assign new_P2_R1275_U43 = ~new_P2_R1275_U61 | ~new_P2_R1275_U106;
  assign new_P2_R1275_U44 = ~new_P2_R1275_U50 | ~new_P2_R1275_U107 | ~new_P2_R1275_U75;
  assign new_P2_R1275_U45 = ~new_P2_R1275_U49 | ~new_P2_R1275_U108 | ~new_P2_R1275_U73;
  assign new_P2_R1275_U46 = ~new_P2_R1275_U48 | ~new_P2_R1275_U109 | ~new_P2_R1275_U71;
  assign new_P2_R1275_U47 = ~new_P2_U3959;
  assign new_P2_R1275_U48 = ~new_P2_U3949;
  assign new_P2_R1275_U49 = ~new_P2_U3951;
  assign new_P2_R1275_U50 = ~new_P2_U3953;
  assign new_P2_R1275_U51 = ~new_P2_U3477;
  assign new_P2_R1275_U52 = ~new_P2_U3474;
  assign new_P2_R1275_U53 = ~new_P2_U3465;
  assign new_P2_R1275_U54 = ~new_P2_U3462;
  assign new_P2_R1275_U55 = ~new_P2_R1275_U153 | ~new_P2_R1275_U152;
  assign new_P2_R1275_U56 = ~new_P2_U3444 & ~new_P2_U3447;
  assign new_P2_R1275_U57 = ~new_P2_U3459 & ~new_P2_U3456;
  assign new_P2_R1275_U58 = ~new_P2_U3468 & ~new_P2_U3471;
  assign new_P2_R1275_U59 = ~new_P2_U3480 & ~new_P2_U3483;
  assign new_P2_R1275_U60 = ~new_P2_U3485 & ~new_P2_U3957;
  assign new_P2_R1275_U61 = ~new_P2_U3956 & ~new_P2_U3955;
  assign new_P2_R1275_U62 = ~new_P2_U3456;
  assign new_P2_R1275_U63 = new_P2_R1275_U137 & new_P2_R1275_U136;
  assign new_P2_R1275_U64 = ~new_P2_U3444;
  assign new_P2_R1275_U65 = new_P2_R1275_U139 & new_P2_R1275_U138;
  assign new_P2_R1275_U66 = ~new_P2_U3958;
  assign new_P2_R1275_U67 = ~new_P2_R1275_U47 | ~new_P2_R1275_U110 | ~new_P2_R1275_U69;
  assign new_P2_R1275_U68 = new_P2_R1275_U141 & new_P2_R1275_U140;
  assign new_P2_R1275_U69 = ~new_P2_U3960;
  assign new_P2_R1275_U70 = new_P2_R1275_U143 & new_P2_R1275_U142;
  assign new_P2_R1275_U71 = ~new_P2_U3950;
  assign new_P2_R1275_U72 = new_P2_R1275_U145 & new_P2_R1275_U144;
  assign new_P2_R1275_U73 = ~new_P2_U3952;
  assign new_P2_R1275_U74 = new_P2_R1275_U147 & new_P2_R1275_U146;
  assign new_P2_R1275_U75 = ~new_P2_U3954;
  assign new_P2_R1275_U76 = new_P2_R1275_U149 & new_P2_R1275_U148;
  assign new_P2_R1275_U77 = ~new_P2_U3956;
  assign new_P2_R1275_U78 = new_P2_R1275_U151 & new_P2_R1275_U150;
  assign new_P2_R1275_U79 = ~new_P2_U3432;
  assign new_P2_R1275_U80 = ~new_P2_U3427;
  assign new_P2_R1275_U81 = ~new_P2_U3485;
  assign new_P2_R1275_U82 = new_P2_R1275_U155 & new_P2_R1275_U154;
  assign new_P2_R1275_U83 = ~new_P2_U3480;
  assign new_P2_R1275_U84 = new_P2_R1275_U157 & new_P2_R1275_U156;
  assign new_P2_R1275_U85 = ~new_P2_U3468;
  assign new_P2_R1275_U86 = new_P2_R1275_U159 & new_P2_R1275_U158;
  assign new_P2_R1275_U87 = ~new_P2_R1275_U25;
  assign new_P2_R1275_U88 = ~new_P2_R1275_U26;
  assign new_P2_R1275_U89 = ~new_P2_R1275_U27;
  assign new_P2_R1275_U90 = ~new_P2_R1275_U28;
  assign new_P2_R1275_U91 = ~new_P2_R1275_U29;
  assign new_P2_R1275_U92 = ~new_P2_R1275_U30;
  assign new_P2_R1275_U93 = ~new_P2_U3453 | ~new_P2_R1275_U29;
  assign new_P2_R1275_U94 = ~new_P2_U3450 | ~new_P2_R1275_U28;
  assign new_P2_R1275_U95 = ~new_P2_R1275_U89 | ~new_P2_R1275_U64;
  assign new_P2_R1275_U96 = ~new_P2_U3447 | ~new_P2_R1275_U95;
  assign new_P2_R1275_U97 = ~new_P2_U3441 | ~new_P2_R1275_U26;
  assign new_P2_R1275_U98 = ~new_P2_U3438 | ~new_P2_R1275_U25;
  assign new_P2_R1275_U99 = ~new_P2_R1275_U35;
  assign new_P2_R1275_U100 = ~new_P2_R1275_U36;
  assign new_P2_R1275_U101 = ~new_P2_R1275_U37;
  assign new_P2_R1275_U102 = ~new_P2_R1275_U38;
  assign new_P2_R1275_U103 = ~new_P2_R1275_U39;
  assign new_P2_R1275_U104 = ~new_P2_R1275_U40;
  assign new_P2_R1275_U105 = ~new_P2_R1275_U41;
  assign new_P2_R1275_U106 = ~new_P2_R1275_U42;
  assign new_P2_R1275_U107 = ~new_P2_R1275_U43;
  assign new_P2_R1275_U108 = ~new_P2_R1275_U44;
  assign new_P2_R1275_U109 = ~new_P2_R1275_U45;
  assign new_P2_R1275_U110 = ~new_P2_R1275_U46;
  assign new_P2_R1275_U111 = ~new_P2_R1275_U67;
  assign new_P2_R1275_U112 = ~new_P2_R1275_U110 | ~new_P2_R1275_U69;
  assign new_P2_R1275_U113 = ~new_P2_U3959 | ~new_P2_R1275_U112;
  assign new_P2_R1275_U114 = new_P2_U3432 | new_P2_U3427;
  assign new_P2_R1275_U115 = ~new_P2_U3435 | ~new_P2_R1275_U114;
  assign new_P2_R1275_U116 = ~new_P2_R1275_U109 | ~new_P2_R1275_U71;
  assign new_P2_R1275_U117 = ~new_P2_U3949 | ~new_P2_R1275_U116;
  assign new_P2_R1275_U118 = ~new_P2_R1275_U108 | ~new_P2_R1275_U73;
  assign new_P2_R1275_U119 = ~new_P2_U3951 | ~new_P2_R1275_U118;
  assign new_P2_R1275_U120 = ~new_P2_R1275_U107 | ~new_P2_R1275_U75;
  assign new_P2_R1275_U121 = ~new_P2_U3953 | ~new_P2_R1275_U120;
  assign new_P2_R1275_U122 = ~new_P2_R1275_U106 | ~new_P2_R1275_U77;
  assign new_P2_R1275_U123 = ~new_P2_U3955 | ~new_P2_R1275_U122;
  assign new_P2_R1275_U124 = ~new_P2_R1275_U105 | ~new_P2_R1275_U81;
  assign new_P2_R1275_U125 = ~new_P2_U3957 | ~new_P2_R1275_U124;
  assign new_P2_R1275_U126 = ~new_P2_R1275_U104 | ~new_P2_R1275_U83;
  assign new_P2_R1275_U127 = ~new_P2_U3483 | ~new_P2_R1275_U126;
  assign new_P2_R1275_U128 = ~new_P2_U3477 | ~new_P2_R1275_U39;
  assign new_P2_R1275_U129 = ~new_P2_U3474 | ~new_P2_R1275_U38;
  assign new_P2_R1275_U130 = ~new_P2_R1275_U101 | ~new_P2_R1275_U85;
  assign new_P2_R1275_U131 = ~new_P2_U3471 | ~new_P2_R1275_U130;
  assign new_P2_R1275_U132 = ~new_P2_U3465 | ~new_P2_R1275_U36;
  assign new_P2_R1275_U133 = ~new_P2_U3462 | ~new_P2_R1275_U35;
  assign new_P2_R1275_U134 = ~new_P2_R1275_U92 | ~new_P2_R1275_U62;
  assign new_P2_R1275_U135 = ~new_P2_U3459 | ~new_P2_R1275_U134;
  assign new_P2_R1275_U136 = ~new_P2_U3456 | ~new_P2_R1275_U30;
  assign new_P2_R1275_U137 = ~new_P2_R1275_U92 | ~new_P2_R1275_U62;
  assign new_P2_R1275_U138 = ~new_P2_U3444 | ~new_P2_R1275_U27;
  assign new_P2_R1275_U139 = ~new_P2_R1275_U89 | ~new_P2_R1275_U64;
  assign new_P2_R1275_U140 = ~new_P2_U3958 | ~new_P2_R1275_U67;
  assign new_P2_R1275_U141 = ~new_P2_R1275_U111 | ~new_P2_R1275_U66;
  assign new_P2_R1275_U142 = ~new_P2_U3960 | ~new_P2_R1275_U46;
  assign new_P2_R1275_U143 = ~new_P2_R1275_U110 | ~new_P2_R1275_U69;
  assign new_P2_R1275_U144 = ~new_P2_U3950 | ~new_P2_R1275_U45;
  assign new_P2_R1275_U145 = ~new_P2_R1275_U109 | ~new_P2_R1275_U71;
  assign new_P2_R1275_U146 = ~new_P2_U3952 | ~new_P2_R1275_U44;
  assign new_P2_R1275_U147 = ~new_P2_R1275_U108 | ~new_P2_R1275_U73;
  assign new_P2_R1275_U148 = ~new_P2_U3954 | ~new_P2_R1275_U43;
  assign new_P2_R1275_U149 = ~new_P2_R1275_U107 | ~new_P2_R1275_U75;
  assign new_P2_R1275_U150 = ~new_P2_U3956 | ~new_P2_R1275_U42;
  assign new_P2_R1275_U151 = ~new_P2_R1275_U106 | ~new_P2_R1275_U77;
  assign new_P2_R1275_U152 = ~new_P2_U3432 | ~new_P2_R1275_U80;
  assign new_P2_R1275_U153 = ~new_P2_U3427 | ~new_P2_R1275_U79;
  assign new_P2_R1275_U154 = ~new_P2_U3485 | ~new_P2_R1275_U41;
  assign new_P2_R1275_U155 = ~new_P2_R1275_U105 | ~new_P2_R1275_U81;
  assign new_P2_R1275_U156 = ~new_P2_U3480 | ~new_P2_R1275_U40;
  assign new_P2_R1275_U157 = ~new_P2_R1275_U104 | ~new_P2_R1275_U83;
  assign new_P2_R1275_U158 = ~new_P2_U3468 | ~new_P2_R1275_U37;
  assign new_P2_R1275_U159 = ~new_P2_R1275_U101 | ~new_P2_R1275_U85;
  assign new_P2_R1179_U6 = new_P2_R1179_U202 & new_P2_R1179_U201;
  assign new_P2_R1179_U7 = new_P2_R1179_U241 & new_P2_R1179_U240;
  assign new_P2_R1179_U8 = new_P2_R1179_U181 & new_P2_R1179_U256;
  assign new_P2_R1179_U9 = new_P2_R1179_U258 & new_P2_R1179_U257;
  assign new_P2_R1179_U10 = new_P2_R1179_U182 & new_P2_R1179_U282;
  assign new_P2_R1179_U11 = new_P2_R1179_U284 & new_P2_R1179_U283;
  assign new_P2_R1179_U12 = ~new_P2_R1179_U344 | ~new_P2_R1179_U347;
  assign new_P2_R1179_U13 = ~new_P2_R1179_U333 | ~new_P2_R1179_U336;
  assign new_P2_R1179_U14 = ~new_P2_R1179_U322 | ~new_P2_R1179_U325;
  assign new_P2_R1179_U15 = ~new_P2_R1179_U314 | ~new_P2_R1179_U316;
  assign new_P2_R1179_U16 = ~new_P2_R1179_U352 | ~new_P2_R1179_U312;
  assign new_P2_R1179_U17 = ~new_P2_R1179_U235 | ~new_P2_R1179_U237;
  assign new_P2_R1179_U18 = ~new_P2_R1179_U227 | ~new_P2_R1179_U230;
  assign new_P2_R1179_U19 = ~new_P2_R1179_U219 | ~new_P2_R1179_U221;
  assign new_P2_R1179_U20 = ~new_P2_R1179_U166 | ~new_P2_R1179_U350;
  assign new_P2_R1179_U21 = ~new_P2_U3450;
  assign new_P2_R1179_U22 = ~new_P2_U3444;
  assign new_P2_R1179_U23 = ~new_P2_U3435;
  assign new_P2_R1179_U24 = ~new_P2_U3427;
  assign new_P2_R1179_U25 = ~new_P2_U3080;
  assign new_P2_R1179_U26 = ~new_P2_U3438;
  assign new_P2_R1179_U27 = ~new_P2_U3070;
  assign new_P2_R1179_U28 = ~new_P2_U3070 | ~new_P2_R1179_U23;
  assign new_P2_R1179_U29 = ~new_P2_U3066;
  assign new_P2_R1179_U30 = ~new_P2_U3447;
  assign new_P2_R1179_U31 = ~new_P2_U3441;
  assign new_P2_R1179_U32 = ~new_P2_U3073;
  assign new_P2_R1179_U33 = ~new_P2_U3069;
  assign new_P2_R1179_U34 = ~new_P2_U3062;
  assign new_P2_R1179_U35 = ~new_P2_U3062 | ~new_P2_R1179_U31;
  assign new_P2_R1179_U36 = ~new_P2_U3453;
  assign new_P2_R1179_U37 = ~new_P2_U3072;
  assign new_P2_R1179_U38 = ~new_P2_U3072 | ~new_P2_R1179_U21;
  assign new_P2_R1179_U39 = ~new_P2_U3086;
  assign new_P2_R1179_U40 = ~new_P2_U3456;
  assign new_P2_R1179_U41 = ~new_P2_U3085;
  assign new_P2_R1179_U42 = ~new_P2_R1179_U208 | ~new_P2_R1179_U207;
  assign new_P2_R1179_U43 = ~new_P2_R1179_U35 | ~new_P2_R1179_U223;
  assign new_P2_R1179_U44 = ~new_P2_R1179_U351 | ~new_P2_R1179_U192 | ~new_P2_R1179_U176;
  assign new_P2_R1179_U45 = ~new_P2_U3951;
  assign new_P2_R1179_U46 = ~new_P2_U3459;
  assign new_P2_R1179_U47 = ~new_P2_U3462;
  assign new_P2_R1179_U48 = ~new_P2_U3065;
  assign new_P2_R1179_U49 = ~new_P2_U3064;
  assign new_P2_R1179_U50 = ~new_P2_U3085 | ~new_P2_R1179_U40;
  assign new_P2_R1179_U51 = ~new_P2_U3465;
  assign new_P2_R1179_U52 = ~new_P2_U3074;
  assign new_P2_R1179_U53 = ~new_P2_U3468;
  assign new_P2_R1179_U54 = ~new_P2_U3082;
  assign new_P2_R1179_U55 = ~new_P2_U3477;
  assign new_P2_R1179_U56 = ~new_P2_U3474;
  assign new_P2_R1179_U57 = ~new_P2_U3471;
  assign new_P2_R1179_U58 = ~new_P2_U3075;
  assign new_P2_R1179_U59 = ~new_P2_U3076;
  assign new_P2_R1179_U60 = ~new_P2_U3081;
  assign new_P2_R1179_U61 = ~new_P2_U3081 | ~new_P2_R1179_U57;
  assign new_P2_R1179_U62 = ~new_P2_U3480;
  assign new_P2_R1179_U63 = ~new_P2_U3071;
  assign new_P2_R1179_U64 = ~new_P2_R1179_U268 | ~new_P2_R1179_U267;
  assign new_P2_R1179_U65 = ~new_P2_U3084;
  assign new_P2_R1179_U66 = ~new_P2_U3485;
  assign new_P2_R1179_U67 = ~new_P2_U3083;
  assign new_P2_R1179_U68 = ~new_P2_U3957;
  assign new_P2_R1179_U69 = ~new_P2_U3078;
  assign new_P2_R1179_U70 = ~new_P2_U3954;
  assign new_P2_R1179_U71 = ~new_P2_U3955;
  assign new_P2_R1179_U72 = ~new_P2_U3956;
  assign new_P2_R1179_U73 = ~new_P2_U3068;
  assign new_P2_R1179_U74 = ~new_P2_U3063;
  assign new_P2_R1179_U75 = ~new_P2_U3077;
  assign new_P2_R1179_U76 = ~new_P2_U3077 | ~new_P2_R1179_U72;
  assign new_P2_R1179_U77 = ~new_P2_U3953;
  assign new_P2_R1179_U78 = ~new_P2_U3067;
  assign new_P2_R1179_U79 = ~new_P2_U3952;
  assign new_P2_R1179_U80 = ~new_P2_U3060;
  assign new_P2_R1179_U81 = ~new_P2_U3950;
  assign new_P2_R1179_U82 = ~new_P2_U3059;
  assign new_P2_R1179_U83 = ~new_P2_U3059 | ~new_P2_R1179_U45;
  assign new_P2_R1179_U84 = ~new_P2_U3055;
  assign new_P2_R1179_U85 = ~new_P2_U3949;
  assign new_P2_R1179_U86 = ~new_P2_U3056;
  assign new_P2_R1179_U87 = ~new_P2_R1179_U128 | ~new_P2_R1179_U301;
  assign new_P2_R1179_U88 = ~new_P2_R1179_U298 | ~new_P2_R1179_U297;
  assign new_P2_R1179_U89 = ~new_P2_R1179_U76 | ~new_P2_R1179_U318;
  assign new_P2_R1179_U90 = ~new_P2_R1179_U61 | ~new_P2_R1179_U329;
  assign new_P2_R1179_U91 = ~new_P2_R1179_U50 | ~new_P2_R1179_U340;
  assign new_P2_R1179_U92 = ~new_P2_U3079;
  assign new_P2_R1179_U93 = ~new_P2_R1179_U395 | ~new_P2_R1179_U394;
  assign new_P2_R1179_U94 = ~new_P2_R1179_U409 | ~new_P2_R1179_U408;
  assign new_P2_R1179_U95 = ~new_P2_R1179_U414 | ~new_P2_R1179_U413;
  assign new_P2_R1179_U96 = ~new_P2_R1179_U430 | ~new_P2_R1179_U429;
  assign new_P2_R1179_U97 = ~new_P2_R1179_U435 | ~new_P2_R1179_U434;
  assign new_P2_R1179_U98 = ~new_P2_R1179_U440 | ~new_P2_R1179_U439;
  assign new_P2_R1179_U99 = ~new_P2_R1179_U445 | ~new_P2_R1179_U444;
  assign new_P2_R1179_U100 = ~new_P2_R1179_U450 | ~new_P2_R1179_U449;
  assign new_P2_R1179_U101 = ~new_P2_R1179_U466 | ~new_P2_R1179_U465;
  assign new_P2_R1179_U102 = ~new_P2_R1179_U471 | ~new_P2_R1179_U470;
  assign new_P2_R1179_U103 = ~new_P2_R1179_U356 | ~new_P2_R1179_U355;
  assign new_P2_R1179_U104 = ~new_P2_R1179_U365 | ~new_P2_R1179_U364;
  assign new_P2_R1179_U105 = ~new_P2_R1179_U372 | ~new_P2_R1179_U371;
  assign new_P2_R1179_U106 = ~new_P2_R1179_U376 | ~new_P2_R1179_U375;
  assign new_P2_R1179_U107 = ~new_P2_R1179_U385 | ~new_P2_R1179_U384;
  assign new_P2_R1179_U108 = ~new_P2_R1179_U404 | ~new_P2_R1179_U403;
  assign new_P2_R1179_U109 = ~new_P2_R1179_U421 | ~new_P2_R1179_U420;
  assign new_P2_R1179_U110 = ~new_P2_R1179_U425 | ~new_P2_R1179_U424;
  assign new_P2_R1179_U111 = ~new_P2_R1179_U457 | ~new_P2_R1179_U456;
  assign new_P2_R1179_U112 = ~new_P2_R1179_U461 | ~new_P2_R1179_U460;
  assign new_P2_R1179_U113 = ~new_P2_R1179_U478 | ~new_P2_R1179_U477;
  assign new_P2_R1179_U114 = new_P2_R1179_U194 & new_P2_R1179_U184;
  assign new_P2_R1179_U115 = new_P2_R1179_U197 & new_P2_R1179_U198;
  assign new_P2_R1179_U116 = new_P2_R1179_U185 & new_P2_R1179_U205 & new_P2_R1179_U200;
  assign new_P2_R1179_U117 = new_P2_R1179_U210 & new_P2_R1179_U186;
  assign new_P2_R1179_U118 = new_P2_R1179_U213 & new_P2_R1179_U214;
  assign new_P2_R1179_U119 = new_P2_R1179_U38 & new_P2_R1179_U358 & new_P2_R1179_U357;
  assign new_P2_R1179_U120 = new_P2_R1179_U361 & new_P2_R1179_U186;
  assign new_P2_R1179_U121 = new_P2_R1179_U229 & new_P2_R1179_U6;
  assign new_P2_R1179_U122 = new_P2_R1179_U368 & new_P2_R1179_U185;
  assign new_P2_R1179_U123 = new_P2_R1179_U28 & new_P2_R1179_U378 & new_P2_R1179_U377;
  assign new_P2_R1179_U124 = new_P2_R1179_U381 & new_P2_R1179_U184;
  assign new_P2_R1179_U125 = new_P2_R1179_U180 & new_P2_R1179_U239 & new_P2_R1179_U216;
  assign new_P2_R1179_U126 = new_P2_R1179_U261 & new_P2_R1179_U8;
  assign new_P2_R1179_U127 = new_P2_R1179_U287 & new_P2_R1179_U10;
  assign new_P2_R1179_U128 = new_P2_R1179_U303 & new_P2_R1179_U304;
  assign new_P2_R1179_U129 = new_P2_R1179_U311 & new_P2_R1179_U387 & new_P2_R1179_U386;
  assign new_P2_R1179_U130 = new_P2_R1179_U308 & new_P2_R1179_U390;
  assign new_P2_R1179_U131 = ~new_P2_R1179_U392 | ~new_P2_R1179_U391;
  assign new_P2_R1179_U132 = new_P2_R1179_U83 & new_P2_R1179_U397 & new_P2_R1179_U396;
  assign new_P2_R1179_U133 = new_P2_R1179_U400 & new_P2_R1179_U183;
  assign new_P2_R1179_U134 = ~new_P2_R1179_U406 | ~new_P2_R1179_U405;
  assign new_P2_R1179_U135 = ~new_P2_R1179_U411 | ~new_P2_R1179_U410;
  assign new_P2_R1179_U136 = new_P2_R1179_U324 & new_P2_R1179_U11;
  assign new_P2_R1179_U137 = new_P2_R1179_U417 & new_P2_R1179_U182;
  assign new_P2_R1179_U138 = ~new_P2_R1179_U427 | ~new_P2_R1179_U426;
  assign new_P2_R1179_U139 = ~new_P2_R1179_U432 | ~new_P2_R1179_U431;
  assign new_P2_R1179_U140 = ~new_P2_R1179_U437 | ~new_P2_R1179_U436;
  assign new_P2_R1179_U141 = ~new_P2_R1179_U442 | ~new_P2_R1179_U441;
  assign new_P2_R1179_U142 = ~new_P2_R1179_U447 | ~new_P2_R1179_U446;
  assign new_P2_R1179_U143 = new_P2_R1179_U335 & new_P2_R1179_U9;
  assign new_P2_R1179_U144 = new_P2_R1179_U453 & new_P2_R1179_U181;
  assign new_P2_R1179_U145 = ~new_P2_R1179_U463 | ~new_P2_R1179_U462;
  assign new_P2_R1179_U146 = ~new_P2_R1179_U468 | ~new_P2_R1179_U467;
  assign new_P2_R1179_U147 = new_P2_R1179_U346 & new_P2_R1179_U7;
  assign new_P2_R1179_U148 = new_P2_R1179_U474 & new_P2_R1179_U180;
  assign new_P2_R1179_U149 = new_P2_R1179_U354 & new_P2_R1179_U353;
  assign new_P2_R1179_U150 = ~new_P2_R1179_U118 | ~new_P2_R1179_U211;
  assign new_P2_R1179_U151 = new_P2_R1179_U363 & new_P2_R1179_U362;
  assign new_P2_R1179_U152 = new_P2_R1179_U370 & new_P2_R1179_U369;
  assign new_P2_R1179_U153 = new_P2_R1179_U374 & new_P2_R1179_U373;
  assign new_P2_R1179_U154 = ~new_P2_R1179_U115 | ~new_P2_R1179_U195;
  assign new_P2_R1179_U155 = new_P2_R1179_U383 & new_P2_R1179_U382;
  assign new_P2_R1179_U156 = ~new_P2_U3960;
  assign new_P2_R1179_U157 = ~new_P2_U3057;
  assign new_P2_R1179_U158 = new_P2_R1179_U402 & new_P2_R1179_U401;
  assign new_P2_R1179_U159 = ~new_P2_R1179_U294 | ~new_P2_R1179_U293;
  assign new_P2_R1179_U160 = ~new_P2_R1179_U290 | ~new_P2_R1179_U289;
  assign new_P2_R1179_U161 = new_P2_R1179_U419 & new_P2_R1179_U418;
  assign new_P2_R1179_U162 = new_P2_R1179_U423 & new_P2_R1179_U422;
  assign new_P2_R1179_U163 = ~new_P2_R1179_U280 | ~new_P2_R1179_U279;
  assign new_P2_R1179_U164 = ~new_P2_R1179_U276 | ~new_P2_R1179_U275;
  assign new_P2_R1179_U165 = ~new_P2_U3432;
  assign new_P2_R1179_U166 = ~new_P2_U3427 | ~new_P2_R1179_U92;
  assign new_P2_R1179_U167 = ~new_P2_R1179_U272 | ~new_P2_R1179_U271;
  assign new_P2_R1179_U168 = ~new_P2_U3483;
  assign new_P2_R1179_U169 = ~new_P2_R1179_U264 | ~new_P2_R1179_U263;
  assign new_P2_R1179_U170 = new_P2_R1179_U455 & new_P2_R1179_U454;
  assign new_P2_R1179_U171 = new_P2_R1179_U459 & new_P2_R1179_U458;
  assign new_P2_R1179_U172 = ~new_P2_R1179_U254 | ~new_P2_R1179_U253;
  assign new_P2_R1179_U173 = ~new_P2_R1179_U250 | ~new_P2_R1179_U249;
  assign new_P2_R1179_U174 = ~new_P2_R1179_U246 | ~new_P2_R1179_U245;
  assign new_P2_R1179_U175 = new_P2_R1179_U476 & new_P2_R1179_U475;
  assign new_P2_R1179_U176 = ~new_P2_R1179_U166 | ~new_P2_R1179_U165;
  assign new_P2_R1179_U177 = ~new_P2_R1179_U83;
  assign new_P2_R1179_U178 = ~new_P2_R1179_U28;
  assign new_P2_R1179_U179 = ~new_P2_R1179_U38;
  assign new_P2_R1179_U180 = ~new_P2_U3459 | ~new_P2_R1179_U49;
  assign new_P2_R1179_U181 = ~new_P2_U3474 | ~new_P2_R1179_U59;
  assign new_P2_R1179_U182 = ~new_P2_U3955 | ~new_P2_R1179_U74;
  assign new_P2_R1179_U183 = ~new_P2_U3951 | ~new_P2_R1179_U82;
  assign new_P2_R1179_U184 = ~new_P2_U3435 | ~new_P2_R1179_U27;
  assign new_P2_R1179_U185 = ~new_P2_U3444 | ~new_P2_R1179_U33;
  assign new_P2_R1179_U186 = ~new_P2_U3450 | ~new_P2_R1179_U37;
  assign new_P2_R1179_U187 = ~new_P2_R1179_U61;
  assign new_P2_R1179_U188 = ~new_P2_R1179_U76;
  assign new_P2_R1179_U189 = ~new_P2_R1179_U35;
  assign new_P2_R1179_U190 = ~new_P2_R1179_U50;
  assign new_P2_R1179_U191 = ~new_P2_R1179_U166;
  assign new_P2_R1179_U192 = ~new_P2_U3080 | ~new_P2_R1179_U166;
  assign new_P2_R1179_U193 = ~new_P2_R1179_U44;
  assign new_P2_R1179_U194 = ~new_P2_U3438 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U195 = ~new_P2_R1179_U114 | ~new_P2_R1179_U44;
  assign new_P2_R1179_U196 = ~new_P2_R1179_U29 | ~new_P2_R1179_U28;
  assign new_P2_R1179_U197 = ~new_P2_R1179_U196 | ~new_P2_R1179_U26;
  assign new_P2_R1179_U198 = ~new_P2_U3066 | ~new_P2_R1179_U178;
  assign new_P2_R1179_U199 = ~new_P2_R1179_U154;
  assign new_P2_R1179_U200 = ~new_P2_U3447 | ~new_P2_R1179_U32;
  assign new_P2_R1179_U201 = ~new_P2_U3073 | ~new_P2_R1179_U30;
  assign new_P2_R1179_U202 = ~new_P2_U3069 | ~new_P2_R1179_U22;
  assign new_P2_R1179_U203 = ~new_P2_R1179_U189 | ~new_P2_R1179_U185;
  assign new_P2_R1179_U204 = ~new_P2_R1179_U6 | ~new_P2_R1179_U203;
  assign new_P2_R1179_U205 = ~new_P2_U3441 | ~new_P2_R1179_U34;
  assign new_P2_R1179_U206 = ~new_P2_U3447 | ~new_P2_R1179_U32;
  assign new_P2_R1179_U207 = ~new_P2_R1179_U154 | ~new_P2_R1179_U116;
  assign new_P2_R1179_U208 = ~new_P2_R1179_U206 | ~new_P2_R1179_U204;
  assign new_P2_R1179_U209 = ~new_P2_R1179_U42;
  assign new_P2_R1179_U210 = ~new_P2_U3453 | ~new_P2_R1179_U39;
  assign new_P2_R1179_U211 = ~new_P2_R1179_U117 | ~new_P2_R1179_U42;
  assign new_P2_R1179_U212 = ~new_P2_R1179_U39 | ~new_P2_R1179_U38;
  assign new_P2_R1179_U213 = ~new_P2_R1179_U212 | ~new_P2_R1179_U36;
  assign new_P2_R1179_U214 = ~new_P2_U3086 | ~new_P2_R1179_U179;
  assign new_P2_R1179_U215 = ~new_P2_R1179_U150;
  assign new_P2_R1179_U216 = ~new_P2_U3456 | ~new_P2_R1179_U41;
  assign new_P2_R1179_U217 = ~new_P2_R1179_U216 | ~new_P2_R1179_U50;
  assign new_P2_R1179_U218 = ~new_P2_R1179_U209 | ~new_P2_R1179_U38;
  assign new_P2_R1179_U219 = ~new_P2_R1179_U120 | ~new_P2_R1179_U218;
  assign new_P2_R1179_U220 = ~new_P2_R1179_U42 | ~new_P2_R1179_U186;
  assign new_P2_R1179_U221 = ~new_P2_R1179_U119 | ~new_P2_R1179_U220;
  assign new_P2_R1179_U222 = ~new_P2_R1179_U38 | ~new_P2_R1179_U186;
  assign new_P2_R1179_U223 = ~new_P2_R1179_U205 | ~new_P2_R1179_U154;
  assign new_P2_R1179_U224 = ~new_P2_R1179_U43;
  assign new_P2_R1179_U225 = ~new_P2_U3069 | ~new_P2_R1179_U22;
  assign new_P2_R1179_U226 = ~new_P2_R1179_U224 | ~new_P2_R1179_U225;
  assign new_P2_R1179_U227 = ~new_P2_R1179_U122 | ~new_P2_R1179_U226;
  assign new_P2_R1179_U228 = ~new_P2_R1179_U43 | ~new_P2_R1179_U185;
  assign new_P2_R1179_U229 = ~new_P2_U3447 | ~new_P2_R1179_U32;
  assign new_P2_R1179_U230 = ~new_P2_R1179_U121 | ~new_P2_R1179_U228;
  assign new_P2_R1179_U231 = ~new_P2_U3069 | ~new_P2_R1179_U22;
  assign new_P2_R1179_U232 = ~new_P2_R1179_U185 | ~new_P2_R1179_U231;
  assign new_P2_R1179_U233 = ~new_P2_R1179_U205 | ~new_P2_R1179_U35;
  assign new_P2_R1179_U234 = ~new_P2_R1179_U193 | ~new_P2_R1179_U28;
  assign new_P2_R1179_U235 = ~new_P2_R1179_U124 | ~new_P2_R1179_U234;
  assign new_P2_R1179_U236 = ~new_P2_R1179_U44 | ~new_P2_R1179_U184;
  assign new_P2_R1179_U237 = ~new_P2_R1179_U123 | ~new_P2_R1179_U236;
  assign new_P2_R1179_U238 = ~new_P2_R1179_U28 | ~new_P2_R1179_U184;
  assign new_P2_R1179_U239 = ~new_P2_U3462 | ~new_P2_R1179_U48;
  assign new_P2_R1179_U240 = ~new_P2_U3065 | ~new_P2_R1179_U47;
  assign new_P2_R1179_U241 = ~new_P2_U3064 | ~new_P2_R1179_U46;
  assign new_P2_R1179_U242 = ~new_P2_R1179_U190 | ~new_P2_R1179_U180;
  assign new_P2_R1179_U243 = ~new_P2_R1179_U7 | ~new_P2_R1179_U242;
  assign new_P2_R1179_U244 = ~new_P2_U3462 | ~new_P2_R1179_U48;
  assign new_P2_R1179_U245 = ~new_P2_R1179_U150 | ~new_P2_R1179_U125;
  assign new_P2_R1179_U246 = ~new_P2_R1179_U244 | ~new_P2_R1179_U243;
  assign new_P2_R1179_U247 = ~new_P2_R1179_U174;
  assign new_P2_R1179_U248 = ~new_P2_U3465 | ~new_P2_R1179_U52;
  assign new_P2_R1179_U249 = ~new_P2_R1179_U248 | ~new_P2_R1179_U174;
  assign new_P2_R1179_U250 = ~new_P2_U3074 | ~new_P2_R1179_U51;
  assign new_P2_R1179_U251 = ~new_P2_R1179_U173;
  assign new_P2_R1179_U252 = ~new_P2_U3468 | ~new_P2_R1179_U54;
  assign new_P2_R1179_U253 = ~new_P2_R1179_U252 | ~new_P2_R1179_U173;
  assign new_P2_R1179_U254 = ~new_P2_U3082 | ~new_P2_R1179_U53;
  assign new_P2_R1179_U255 = ~new_P2_R1179_U172;
  assign new_P2_R1179_U256 = ~new_P2_U3477 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U257 = ~new_P2_U3075 | ~new_P2_R1179_U55;
  assign new_P2_R1179_U258 = ~new_P2_U3076 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U259 = ~new_P2_R1179_U187 | ~new_P2_R1179_U8;
  assign new_P2_R1179_U260 = ~new_P2_R1179_U9 | ~new_P2_R1179_U259;
  assign new_P2_R1179_U261 = ~new_P2_U3471 | ~new_P2_R1179_U60;
  assign new_P2_R1179_U262 = ~new_P2_U3477 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U263 = ~new_P2_R1179_U126 | ~new_P2_R1179_U172;
  assign new_P2_R1179_U264 = ~new_P2_R1179_U262 | ~new_P2_R1179_U260;
  assign new_P2_R1179_U265 = ~new_P2_R1179_U169;
  assign new_P2_R1179_U266 = ~new_P2_U3480 | ~new_P2_R1179_U63;
  assign new_P2_R1179_U267 = ~new_P2_R1179_U266 | ~new_P2_R1179_U169;
  assign new_P2_R1179_U268 = ~new_P2_U3071 | ~new_P2_R1179_U62;
  assign new_P2_R1179_U269 = ~new_P2_R1179_U64;
  assign new_P2_R1179_U270 = ~new_P2_R1179_U269 | ~new_P2_R1179_U65;
  assign new_P2_R1179_U271 = ~new_P2_R1179_U270 | ~new_P2_R1179_U168;
  assign new_P2_R1179_U272 = ~new_P2_U3084 | ~new_P2_R1179_U64;
  assign new_P2_R1179_U273 = ~new_P2_R1179_U167;
  assign new_P2_R1179_U274 = ~new_P2_U3485 | ~new_P2_R1179_U67;
  assign new_P2_R1179_U275 = ~new_P2_R1179_U274 | ~new_P2_R1179_U167;
  assign new_P2_R1179_U276 = ~new_P2_U3083 | ~new_P2_R1179_U66;
  assign new_P2_R1179_U277 = ~new_P2_R1179_U164;
  assign new_P2_R1179_U278 = ~new_P2_U3957 | ~new_P2_R1179_U69;
  assign new_P2_R1179_U279 = ~new_P2_R1179_U278 | ~new_P2_R1179_U164;
  assign new_P2_R1179_U280 = ~new_P2_U3078 | ~new_P2_R1179_U68;
  assign new_P2_R1179_U281 = ~new_P2_R1179_U163;
  assign new_P2_R1179_U282 = ~new_P2_U3954 | ~new_P2_R1179_U73;
  assign new_P2_R1179_U283 = ~new_P2_U3068 | ~new_P2_R1179_U70;
  assign new_P2_R1179_U284 = ~new_P2_U3063 | ~new_P2_R1179_U71;
  assign new_P2_R1179_U285 = ~new_P2_R1179_U188 | ~new_P2_R1179_U10;
  assign new_P2_R1179_U286 = ~new_P2_R1179_U11 | ~new_P2_R1179_U285;
  assign new_P2_R1179_U287 = ~new_P2_U3956 | ~new_P2_R1179_U75;
  assign new_P2_R1179_U288 = ~new_P2_U3954 | ~new_P2_R1179_U73;
  assign new_P2_R1179_U289 = ~new_P2_R1179_U127 | ~new_P2_R1179_U163;
  assign new_P2_R1179_U290 = ~new_P2_R1179_U288 | ~new_P2_R1179_U286;
  assign new_P2_R1179_U291 = ~new_P2_R1179_U160;
  assign new_P2_R1179_U292 = ~new_P2_U3953 | ~new_P2_R1179_U78;
  assign new_P2_R1179_U293 = ~new_P2_R1179_U292 | ~new_P2_R1179_U160;
  assign new_P2_R1179_U294 = ~new_P2_U3067 | ~new_P2_R1179_U77;
  assign new_P2_R1179_U295 = ~new_P2_R1179_U159;
  assign new_P2_R1179_U296 = ~new_P2_U3952 | ~new_P2_R1179_U80;
  assign new_P2_R1179_U297 = ~new_P2_R1179_U296 | ~new_P2_R1179_U159;
  assign new_P2_R1179_U298 = ~new_P2_U3060 | ~new_P2_R1179_U79;
  assign new_P2_R1179_U299 = ~new_P2_R1179_U88;
  assign new_P2_R1179_U300 = ~new_P2_U3950 | ~new_P2_R1179_U84;
  assign new_P2_R1179_U301 = ~new_P2_R1179_U300 | ~new_P2_R1179_U88 | ~new_P2_R1179_U183;
  assign new_P2_R1179_U302 = ~new_P2_R1179_U84 | ~new_P2_R1179_U83;
  assign new_P2_R1179_U303 = ~new_P2_R1179_U302 | ~new_P2_R1179_U81;
  assign new_P2_R1179_U304 = ~new_P2_U3055 | ~new_P2_R1179_U177;
  assign new_P2_R1179_U305 = ~new_P2_R1179_U87;
  assign new_P2_R1179_U306 = ~new_P2_U3056 | ~new_P2_R1179_U85;
  assign new_P2_R1179_U307 = ~new_P2_R1179_U305 | ~new_P2_R1179_U306;
  assign new_P2_R1179_U308 = ~new_P2_U3949 | ~new_P2_R1179_U86;
  assign new_P2_R1179_U309 = ~new_P2_U3949 | ~new_P2_R1179_U86;
  assign new_P2_R1179_U310 = ~new_P2_R1179_U309 | ~new_P2_R1179_U87;
  assign new_P2_R1179_U311 = ~new_P2_U3056 | ~new_P2_R1179_U85;
  assign new_P2_R1179_U312 = ~new_P2_R1179_U129 | ~new_P2_R1179_U310;
  assign new_P2_R1179_U313 = ~new_P2_R1179_U299 | ~new_P2_R1179_U83;
  assign new_P2_R1179_U314 = ~new_P2_R1179_U133 | ~new_P2_R1179_U313;
  assign new_P2_R1179_U315 = ~new_P2_R1179_U88 | ~new_P2_R1179_U183;
  assign new_P2_R1179_U316 = ~new_P2_R1179_U132 | ~new_P2_R1179_U315;
  assign new_P2_R1179_U317 = ~new_P2_R1179_U83 | ~new_P2_R1179_U183;
  assign new_P2_R1179_U318 = ~new_P2_R1179_U287 | ~new_P2_R1179_U163;
  assign new_P2_R1179_U319 = ~new_P2_R1179_U89;
  assign new_P2_R1179_U320 = ~new_P2_U3063 | ~new_P2_R1179_U71;
  assign new_P2_R1179_U321 = ~new_P2_R1179_U319 | ~new_P2_R1179_U320;
  assign new_P2_R1179_U322 = ~new_P2_R1179_U137 | ~new_P2_R1179_U321;
  assign new_P2_R1179_U323 = ~new_P2_R1179_U89 | ~new_P2_R1179_U182;
  assign new_P2_R1179_U324 = ~new_P2_U3954 | ~new_P2_R1179_U73;
  assign new_P2_R1179_U325 = ~new_P2_R1179_U136 | ~new_P2_R1179_U323;
  assign new_P2_R1179_U326 = ~new_P2_U3063 | ~new_P2_R1179_U71;
  assign new_P2_R1179_U327 = ~new_P2_R1179_U182 | ~new_P2_R1179_U326;
  assign new_P2_R1179_U328 = ~new_P2_R1179_U287 | ~new_P2_R1179_U76;
  assign new_P2_R1179_U329 = ~new_P2_R1179_U261 | ~new_P2_R1179_U172;
  assign new_P2_R1179_U330 = ~new_P2_R1179_U90;
  assign new_P2_R1179_U331 = ~new_P2_U3076 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U332 = ~new_P2_R1179_U330 | ~new_P2_R1179_U331;
  assign new_P2_R1179_U333 = ~new_P2_R1179_U144 | ~new_P2_R1179_U332;
  assign new_P2_R1179_U334 = ~new_P2_R1179_U90 | ~new_P2_R1179_U181;
  assign new_P2_R1179_U335 = ~new_P2_U3477 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U336 = ~new_P2_R1179_U143 | ~new_P2_R1179_U334;
  assign new_P2_R1179_U337 = ~new_P2_U3076 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U338 = ~new_P2_R1179_U181 | ~new_P2_R1179_U337;
  assign new_P2_R1179_U339 = ~new_P2_R1179_U261 | ~new_P2_R1179_U61;
  assign new_P2_R1179_U340 = ~new_P2_R1179_U216 | ~new_P2_R1179_U150;
  assign new_P2_R1179_U341 = ~new_P2_R1179_U91;
  assign new_P2_R1179_U342 = ~new_P2_U3064 | ~new_P2_R1179_U46;
  assign new_P2_R1179_U343 = ~new_P2_R1179_U341 | ~new_P2_R1179_U342;
  assign new_P2_R1179_U344 = ~new_P2_R1179_U148 | ~new_P2_R1179_U343;
  assign new_P2_R1179_U345 = ~new_P2_R1179_U91 | ~new_P2_R1179_U180;
  assign new_P2_R1179_U346 = ~new_P2_U3462 | ~new_P2_R1179_U48;
  assign new_P2_R1179_U347 = ~new_P2_R1179_U147 | ~new_P2_R1179_U345;
  assign new_P2_R1179_U348 = ~new_P2_U3064 | ~new_P2_R1179_U46;
  assign new_P2_R1179_U349 = ~new_P2_R1179_U180 | ~new_P2_R1179_U348;
  assign new_P2_R1179_U350 = ~new_P2_U3079 | ~new_P2_R1179_U24;
  assign new_P2_R1179_U351 = ~new_P2_U3080 | ~new_P2_R1179_U165;
  assign new_P2_R1179_U352 = ~new_P2_R1179_U130 | ~new_P2_R1179_U307;
  assign new_P2_R1179_U353 = ~new_P2_U3456 | ~new_P2_R1179_U41;
  assign new_P2_R1179_U354 = ~new_P2_U3085 | ~new_P2_R1179_U40;
  assign new_P2_R1179_U355 = ~new_P2_R1179_U217 | ~new_P2_R1179_U150;
  assign new_P2_R1179_U356 = ~new_P2_R1179_U215 | ~new_P2_R1179_U149;
  assign new_P2_R1179_U357 = ~new_P2_U3453 | ~new_P2_R1179_U39;
  assign new_P2_R1179_U358 = ~new_P2_U3086 | ~new_P2_R1179_U36;
  assign new_P2_R1179_U359 = ~new_P2_U3453 | ~new_P2_R1179_U39;
  assign new_P2_R1179_U360 = ~new_P2_U3086 | ~new_P2_R1179_U36;
  assign new_P2_R1179_U361 = ~new_P2_R1179_U360 | ~new_P2_R1179_U359;
  assign new_P2_R1179_U362 = ~new_P2_U3450 | ~new_P2_R1179_U37;
  assign new_P2_R1179_U363 = ~new_P2_U3072 | ~new_P2_R1179_U21;
  assign new_P2_R1179_U364 = ~new_P2_R1179_U222 | ~new_P2_R1179_U42;
  assign new_P2_R1179_U365 = ~new_P2_R1179_U151 | ~new_P2_R1179_U209;
  assign new_P2_R1179_U366 = ~new_P2_U3447 | ~new_P2_R1179_U32;
  assign new_P2_R1179_U367 = ~new_P2_U3073 | ~new_P2_R1179_U30;
  assign new_P2_R1179_U368 = ~new_P2_R1179_U367 | ~new_P2_R1179_U366;
  assign new_P2_R1179_U369 = ~new_P2_U3444 | ~new_P2_R1179_U33;
  assign new_P2_R1179_U370 = ~new_P2_U3069 | ~new_P2_R1179_U22;
  assign new_P2_R1179_U371 = ~new_P2_R1179_U232 | ~new_P2_R1179_U43;
  assign new_P2_R1179_U372 = ~new_P2_R1179_U152 | ~new_P2_R1179_U224;
  assign new_P2_R1179_U373 = ~new_P2_U3441 | ~new_P2_R1179_U34;
  assign new_P2_R1179_U374 = ~new_P2_U3062 | ~new_P2_R1179_U31;
  assign new_P2_R1179_U375 = ~new_P2_R1179_U233 | ~new_P2_R1179_U154;
  assign new_P2_R1179_U376 = ~new_P2_R1179_U199 | ~new_P2_R1179_U153;
  assign new_P2_R1179_U377 = ~new_P2_U3438 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U378 = ~new_P2_U3066 | ~new_P2_R1179_U26;
  assign new_P2_R1179_U379 = ~new_P2_U3438 | ~new_P2_R1179_U29;
  assign new_P2_R1179_U380 = ~new_P2_U3066 | ~new_P2_R1179_U26;
  assign new_P2_R1179_U381 = ~new_P2_R1179_U380 | ~new_P2_R1179_U379;
  assign new_P2_R1179_U382 = ~new_P2_U3435 | ~new_P2_R1179_U27;
  assign new_P2_R1179_U383 = ~new_P2_U3070 | ~new_P2_R1179_U23;
  assign new_P2_R1179_U384 = ~new_P2_R1179_U238 | ~new_P2_R1179_U44;
  assign new_P2_R1179_U385 = ~new_P2_R1179_U155 | ~new_P2_R1179_U193;
  assign new_P2_R1179_U386 = ~new_P2_U3960 | ~new_P2_R1179_U157;
  assign new_P2_R1179_U387 = ~new_P2_U3057 | ~new_P2_R1179_U156;
  assign new_P2_R1179_U388 = ~new_P2_U3960 | ~new_P2_R1179_U157;
  assign new_P2_R1179_U389 = ~new_P2_U3057 | ~new_P2_R1179_U156;
  assign new_P2_R1179_U390 = ~new_P2_R1179_U389 | ~new_P2_R1179_U388;
  assign new_P2_R1179_U391 = ~new_P2_U3949 | ~new_P2_R1179_U86;
  assign new_P2_R1179_U392 = ~new_P2_U3056 | ~new_P2_R1179_U85;
  assign new_P2_R1179_U393 = ~new_P2_R1179_U131;
  assign new_P2_R1179_U394 = ~new_P2_R1179_U393 | ~new_P2_R1179_U305;
  assign new_P2_R1179_U395 = ~new_P2_R1179_U131 | ~new_P2_R1179_U87;
  assign new_P2_R1179_U396 = ~new_P2_U3950 | ~new_P2_R1179_U84;
  assign new_P2_R1179_U397 = ~new_P2_U3055 | ~new_P2_R1179_U81;
  assign new_P2_R1179_U398 = ~new_P2_U3950 | ~new_P2_R1179_U84;
  assign new_P2_R1179_U399 = ~new_P2_U3055 | ~new_P2_R1179_U81;
  assign new_P2_R1179_U400 = ~new_P2_R1179_U399 | ~new_P2_R1179_U398;
  assign new_P2_R1179_U401 = ~new_P2_U3951 | ~new_P2_R1179_U82;
  assign new_P2_R1179_U402 = ~new_P2_U3059 | ~new_P2_R1179_U45;
  assign new_P2_R1179_U403 = ~new_P2_R1179_U317 | ~new_P2_R1179_U88;
  assign new_P2_R1179_U404 = ~new_P2_R1179_U158 | ~new_P2_R1179_U299;
  assign new_P2_R1179_U405 = ~new_P2_U3952 | ~new_P2_R1179_U80;
  assign new_P2_R1179_U406 = ~new_P2_U3060 | ~new_P2_R1179_U79;
  assign new_P2_R1179_U407 = ~new_P2_R1179_U134;
  assign new_P2_R1179_U408 = ~new_P2_R1179_U295 | ~new_P2_R1179_U407;
  assign new_P2_R1179_U409 = ~new_P2_R1179_U134 | ~new_P2_R1179_U159;
  assign new_P2_R1179_U410 = ~new_P2_U3953 | ~new_P2_R1179_U78;
  assign new_P2_R1179_U411 = ~new_P2_U3067 | ~new_P2_R1179_U77;
  assign new_P2_R1179_U412 = ~new_P2_R1179_U135;
  assign new_P2_R1179_U413 = ~new_P2_R1179_U291 | ~new_P2_R1179_U412;
  assign new_P2_R1179_U414 = ~new_P2_R1179_U135 | ~new_P2_R1179_U160;
  assign new_P2_R1179_U415 = ~new_P2_U3954 | ~new_P2_R1179_U73;
  assign new_P2_R1179_U416 = ~new_P2_U3068 | ~new_P2_R1179_U70;
  assign new_P2_R1179_U417 = ~new_P2_R1179_U416 | ~new_P2_R1179_U415;
  assign new_P2_R1179_U418 = ~new_P2_U3955 | ~new_P2_R1179_U74;
  assign new_P2_R1179_U419 = ~new_P2_U3063 | ~new_P2_R1179_U71;
  assign new_P2_R1179_U420 = ~new_P2_R1179_U327 | ~new_P2_R1179_U89;
  assign new_P2_R1179_U421 = ~new_P2_R1179_U161 | ~new_P2_R1179_U319;
  assign new_P2_R1179_U422 = ~new_P2_U3956 | ~new_P2_R1179_U75;
  assign new_P2_R1179_U423 = ~new_P2_U3077 | ~new_P2_R1179_U72;
  assign new_P2_R1179_U424 = ~new_P2_R1179_U328 | ~new_P2_R1179_U163;
  assign new_P2_R1179_U425 = ~new_P2_R1179_U281 | ~new_P2_R1179_U162;
  assign new_P2_R1179_U426 = ~new_P2_U3957 | ~new_P2_R1179_U69;
  assign new_P2_R1179_U427 = ~new_P2_U3078 | ~new_P2_R1179_U68;
  assign new_P2_R1179_U428 = ~new_P2_R1179_U138;
  assign new_P2_R1179_U429 = ~new_P2_R1179_U277 | ~new_P2_R1179_U428;
  assign new_P2_R1179_U430 = ~new_P2_R1179_U138 | ~new_P2_R1179_U164;
  assign new_P2_R1179_U431 = ~new_P2_U3432 | ~new_P2_R1179_U25;
  assign new_P2_R1179_U432 = ~new_P2_U3080 | ~new_P2_R1179_U165;
  assign new_P2_R1179_U433 = ~new_P2_R1179_U139;
  assign new_P2_R1179_U434 = ~new_P2_R1179_U191 | ~new_P2_R1179_U433;
  assign new_P2_R1179_U435 = ~new_P2_R1179_U139 | ~new_P2_R1179_U166;
  assign new_P2_R1179_U436 = ~new_P2_U3485 | ~new_P2_R1179_U67;
  assign new_P2_R1179_U437 = ~new_P2_U3083 | ~new_P2_R1179_U66;
  assign new_P2_R1179_U438 = ~new_P2_R1179_U140;
  assign new_P2_R1179_U439 = ~new_P2_R1179_U273 | ~new_P2_R1179_U438;
  assign new_P2_R1179_U440 = ~new_P2_R1179_U140 | ~new_P2_R1179_U167;
  assign new_P2_R1179_U441 = ~new_P2_U3483 | ~new_P2_R1179_U65;
  assign new_P2_R1179_U442 = ~new_P2_U3084 | ~new_P2_R1179_U168;
  assign new_P2_R1179_U443 = ~new_P2_R1179_U141;
  assign new_P2_R1179_U444 = ~new_P2_R1179_U443 | ~new_P2_R1179_U269;
  assign new_P2_R1179_U445 = ~new_P2_R1179_U141 | ~new_P2_R1179_U64;
  assign new_P2_R1179_U446 = ~new_P2_U3480 | ~new_P2_R1179_U63;
  assign new_P2_R1179_U447 = ~new_P2_U3071 | ~new_P2_R1179_U62;
  assign new_P2_R1179_U448 = ~new_P2_R1179_U142;
  assign new_P2_R1179_U449 = ~new_P2_R1179_U265 | ~new_P2_R1179_U448;
  assign new_P2_R1179_U450 = ~new_P2_R1179_U142 | ~new_P2_R1179_U169;
  assign new_P2_R1179_U451 = ~new_P2_U3477 | ~new_P2_R1179_U58;
  assign new_P2_R1179_U452 = ~new_P2_U3075 | ~new_P2_R1179_U55;
  assign new_P2_R1179_U453 = ~new_P2_R1179_U452 | ~new_P2_R1179_U451;
  assign new_P2_R1179_U454 = ~new_P2_U3474 | ~new_P2_R1179_U59;
  assign new_P2_R1179_U455 = ~new_P2_U3076 | ~new_P2_R1179_U56;
  assign new_P2_R1179_U456 = ~new_P2_R1179_U338 | ~new_P2_R1179_U90;
  assign new_P2_R1179_U457 = ~new_P2_R1179_U170 | ~new_P2_R1179_U330;
  assign new_P2_R1179_U458 = ~new_P2_U3471 | ~new_P2_R1179_U60;
  assign new_P2_R1179_U459 = ~new_P2_U3081 | ~new_P2_R1179_U57;
  assign new_P2_R1179_U460 = ~new_P2_R1179_U339 | ~new_P2_R1179_U172;
  assign new_P2_R1179_U461 = ~new_P2_R1179_U255 | ~new_P2_R1179_U171;
  assign new_P2_R1179_U462 = ~new_P2_U3468 | ~new_P2_R1179_U54;
  assign new_P2_R1179_U463 = ~new_P2_U3082 | ~new_P2_R1179_U53;
  assign new_P2_R1179_U464 = ~new_P2_R1179_U145;
  assign new_P2_R1179_U465 = ~new_P2_R1179_U251 | ~new_P2_R1179_U464;
  assign new_P2_R1179_U466 = ~new_P2_R1179_U145 | ~new_P2_R1179_U173;
  assign new_P2_R1179_U467 = ~new_P2_U3465 | ~new_P2_R1179_U52;
  assign new_P2_R1179_U468 = ~new_P2_U3074 | ~new_P2_R1179_U51;
  assign new_P2_R1179_U469 = ~new_P2_R1179_U146;
  assign new_P2_R1179_U470 = ~new_P2_R1179_U247 | ~new_P2_R1179_U469;
  assign new_P2_R1179_U471 = ~new_P2_R1179_U146 | ~new_P2_R1179_U174;
  assign new_P2_R1179_U472 = ~new_P2_U3462 | ~new_P2_R1179_U48;
  assign new_P2_R1179_U473 = ~new_P2_U3065 | ~new_P2_R1179_U47;
  assign new_P2_R1179_U474 = ~new_P2_R1179_U473 | ~new_P2_R1179_U472;
  assign new_P2_R1179_U475 = ~new_P2_U3459 | ~new_P2_R1179_U49;
  assign new_P2_R1179_U476 = ~new_P2_U3064 | ~new_P2_R1179_U46;
  assign new_P2_R1179_U477 = ~new_P2_R1179_U349 | ~new_P2_R1179_U91;
  assign new_P2_R1179_U478 = ~new_P2_R1179_U175 | ~new_P2_R1179_U341;
  assign new_P2_R1215_U4 = new_P2_R1215_U179 & new_P2_R1215_U178;
  assign new_P2_R1215_U5 = new_P2_R1215_U180 & new_P2_R1215_U181;
  assign new_P2_R1215_U6 = new_P2_R1215_U197 & new_P2_R1215_U196;
  assign new_P2_R1215_U7 = new_P2_R1215_U237 & new_P2_R1215_U236;
  assign new_P2_R1215_U8 = new_P2_R1215_U246 & new_P2_R1215_U245;
  assign new_P2_R1215_U9 = new_P2_R1215_U264 & new_P2_R1215_U263;
  assign new_P2_R1215_U10 = new_P2_R1215_U272 & new_P2_R1215_U271;
  assign new_P2_R1215_U11 = new_P2_R1215_U351 & new_P2_R1215_U348;
  assign new_P2_R1215_U12 = new_P2_R1215_U344 & new_P2_R1215_U341;
  assign new_P2_R1215_U13 = new_P2_R1215_U335 & new_P2_R1215_U332;
  assign new_P2_R1215_U14 = new_P2_R1215_U326 & new_P2_R1215_U323;
  assign new_P2_R1215_U15 = new_P2_R1215_U320 & new_P2_R1215_U318;
  assign new_P2_R1215_U16 = new_P2_R1215_U313 & new_P2_R1215_U310;
  assign new_P2_R1215_U17 = new_P2_R1215_U235 & new_P2_R1215_U232;
  assign new_P2_R1215_U18 = new_P2_R1215_U227 & new_P2_R1215_U224;
  assign new_P2_R1215_U19 = new_P2_R1215_U213 & new_P2_R1215_U210;
  assign new_P2_R1215_U20 = ~new_P2_U3447;
  assign new_P2_R1215_U21 = ~new_P2_U3073;
  assign new_P2_R1215_U22 = ~new_P2_U3072;
  assign new_P2_R1215_U23 = ~new_P2_U3073 | ~new_P2_U3447;
  assign new_P2_R1215_U24 = ~new_P2_U3450;
  assign new_P2_R1215_U25 = ~new_P2_U3441;
  assign new_P2_R1215_U26 = ~new_P2_U3062;
  assign new_P2_R1215_U27 = ~new_P2_U3069;
  assign new_P2_R1215_U28 = ~new_P2_U3435;
  assign new_P2_R1215_U29 = ~new_P2_U3070;
  assign new_P2_R1215_U30 = ~new_P2_U3427;
  assign new_P2_R1215_U31 = ~new_P2_U3079;
  assign new_P2_R1215_U32 = ~new_P2_U3079 | ~new_P2_U3427;
  assign new_P2_R1215_U33 = ~new_P2_U3438;
  assign new_P2_R1215_U34 = ~new_P2_U3066;
  assign new_P2_R1215_U35 = ~new_P2_U3062 | ~new_P2_U3441;
  assign new_P2_R1215_U36 = ~new_P2_U3444;
  assign new_P2_R1215_U37 = ~new_P2_U3453;
  assign new_P2_R1215_U38 = ~new_P2_U3086;
  assign new_P2_R1215_U39 = ~new_P2_U3085;
  assign new_P2_R1215_U40 = ~new_P2_U3456;
  assign new_P2_R1215_U41 = ~new_P2_R1215_U62 | ~new_P2_R1215_U205;
  assign new_P2_R1215_U42 = ~new_P2_R1215_U118 | ~new_P2_R1215_U193;
  assign new_P2_R1215_U43 = ~new_P2_R1215_U182 | ~new_P2_R1215_U183;
  assign new_P2_R1215_U44 = ~new_P2_U3432 | ~new_P2_U3080;
  assign new_P2_R1215_U45 = ~new_P2_R1215_U122 | ~new_P2_R1215_U219;
  assign new_P2_R1215_U46 = ~new_P2_R1215_U216 | ~new_P2_R1215_U215;
  assign new_P2_R1215_U47 = ~new_P2_U3950;
  assign new_P2_R1215_U48 = ~new_P2_U3055;
  assign new_P2_R1215_U49 = ~new_P2_U3059;
  assign new_P2_R1215_U50 = ~new_P2_U3951;
  assign new_P2_R1215_U51 = ~new_P2_U3952;
  assign new_P2_R1215_U52 = ~new_P2_U3060;
  assign new_P2_R1215_U53 = ~new_P2_U3953;
  assign new_P2_R1215_U54 = ~new_P2_U3067;
  assign new_P2_R1215_U55 = ~new_P2_U3956;
  assign new_P2_R1215_U56 = ~new_P2_U3077;
  assign new_P2_R1215_U57 = ~new_P2_U3477;
  assign new_P2_R1215_U58 = ~new_P2_U3075;
  assign new_P2_R1215_U59 = ~new_P2_U3071;
  assign new_P2_R1215_U60 = ~new_P2_U3075 | ~new_P2_U3477;
  assign new_P2_R1215_U61 = ~new_P2_U3480;
  assign new_P2_R1215_U62 = ~new_P2_U3086 | ~new_P2_U3453;
  assign new_P2_R1215_U63 = ~new_P2_U3459;
  assign new_P2_R1215_U64 = ~new_P2_U3064;
  assign new_P2_R1215_U65 = ~new_P2_U3465;
  assign new_P2_R1215_U66 = ~new_P2_U3074;
  assign new_P2_R1215_U67 = ~new_P2_U3462;
  assign new_P2_R1215_U68 = ~new_P2_U3065;
  assign new_P2_R1215_U69 = ~new_P2_U3065 | ~new_P2_U3462;
  assign new_P2_R1215_U70 = ~new_P2_U3468;
  assign new_P2_R1215_U71 = ~new_P2_U3082;
  assign new_P2_R1215_U72 = ~new_P2_U3471;
  assign new_P2_R1215_U73 = ~new_P2_U3081;
  assign new_P2_R1215_U74 = ~new_P2_U3474;
  assign new_P2_R1215_U75 = ~new_P2_U3076;
  assign new_P2_R1215_U76 = ~new_P2_U3483;
  assign new_P2_R1215_U77 = ~new_P2_U3084;
  assign new_P2_R1215_U78 = ~new_P2_U3084 | ~new_P2_U3483;
  assign new_P2_R1215_U79 = ~new_P2_U3485;
  assign new_P2_R1215_U80 = ~new_P2_U3083;
  assign new_P2_R1215_U81 = ~new_P2_U3083 | ~new_P2_U3485;
  assign new_P2_R1215_U82 = ~new_P2_U3957;
  assign new_P2_R1215_U83 = ~new_P2_U3955;
  assign new_P2_R1215_U84 = ~new_P2_U3063;
  assign new_P2_R1215_U85 = ~new_P2_U3954;
  assign new_P2_R1215_U86 = ~new_P2_U3068;
  assign new_P2_R1215_U87 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1215_U88 = ~new_P2_U3056;
  assign new_P2_R1215_U89 = ~new_P2_U3949;
  assign new_P2_R1215_U90 = ~new_P2_R1215_U306 | ~new_P2_R1215_U176;
  assign new_P2_R1215_U91 = ~new_P2_U3078;
  assign new_P2_R1215_U92 = ~new_P2_R1215_U78 | ~new_P2_R1215_U315;
  assign new_P2_R1215_U93 = ~new_P2_R1215_U261 | ~new_P2_R1215_U260;
  assign new_P2_R1215_U94 = ~new_P2_R1215_U69 | ~new_P2_R1215_U337;
  assign new_P2_R1215_U95 = ~new_P2_R1215_U457 | ~new_P2_R1215_U456;
  assign new_P2_R1215_U96 = ~new_P2_R1215_U504 | ~new_P2_R1215_U503;
  assign new_P2_R1215_U97 = ~new_P2_R1215_U375 | ~new_P2_R1215_U374;
  assign new_P2_R1215_U98 = ~new_P2_R1215_U380 | ~new_P2_R1215_U379;
  assign new_P2_R1215_U99 = ~new_P2_R1215_U387 | ~new_P2_R1215_U386;
  assign new_P2_R1215_U100 = ~new_P2_R1215_U394 | ~new_P2_R1215_U393;
  assign new_P2_R1215_U101 = ~new_P2_R1215_U399 | ~new_P2_R1215_U398;
  assign new_P2_R1215_U102 = ~new_P2_R1215_U408 | ~new_P2_R1215_U407;
  assign new_P2_R1215_U103 = ~new_P2_R1215_U415 | ~new_P2_R1215_U414;
  assign new_P2_R1215_U104 = ~new_P2_R1215_U422 | ~new_P2_R1215_U421;
  assign new_P2_R1215_U105 = ~new_P2_R1215_U429 | ~new_P2_R1215_U428;
  assign new_P2_R1215_U106 = ~new_P2_R1215_U434 | ~new_P2_R1215_U433;
  assign new_P2_R1215_U107 = ~new_P2_R1215_U441 | ~new_P2_R1215_U440;
  assign new_P2_R1215_U108 = ~new_P2_R1215_U448 | ~new_P2_R1215_U447;
  assign new_P2_R1215_U109 = ~new_P2_R1215_U462 | ~new_P2_R1215_U461;
  assign new_P2_R1215_U110 = ~new_P2_R1215_U467 | ~new_P2_R1215_U466;
  assign new_P2_R1215_U111 = ~new_P2_R1215_U474 | ~new_P2_R1215_U473;
  assign new_P2_R1215_U112 = ~new_P2_R1215_U481 | ~new_P2_R1215_U480;
  assign new_P2_R1215_U113 = ~new_P2_R1215_U488 | ~new_P2_R1215_U487;
  assign new_P2_R1215_U114 = ~new_P2_R1215_U495 | ~new_P2_R1215_U494;
  assign new_P2_R1215_U115 = ~new_P2_R1215_U500 | ~new_P2_R1215_U499;
  assign new_P2_R1215_U116 = new_P2_U3435 & new_P2_U3070;
  assign new_P2_R1215_U117 = new_P2_R1215_U189 & new_P2_R1215_U187;
  assign new_P2_R1215_U118 = new_P2_R1215_U194 & new_P2_R1215_U192;
  assign new_P2_R1215_U119 = new_P2_R1215_U201 & new_P2_R1215_U200;
  assign new_P2_R1215_U120 = new_P2_R1215_U23 & new_P2_R1215_U382 & new_P2_R1215_U381;
  assign new_P2_R1215_U121 = new_P2_R1215_U212 & new_P2_R1215_U6;
  assign new_P2_R1215_U122 = new_P2_R1215_U220 & new_P2_R1215_U218;
  assign new_P2_R1215_U123 = new_P2_R1215_U35 & new_P2_R1215_U389 & new_P2_R1215_U388;
  assign new_P2_R1215_U124 = new_P2_R1215_U226 & new_P2_R1215_U4;
  assign new_P2_R1215_U125 = new_P2_R1215_U234 & new_P2_R1215_U181;
  assign new_P2_R1215_U126 = new_P2_R1215_U204 & new_P2_R1215_U7;
  assign new_P2_R1215_U127 = new_P2_R1215_U239 & new_P2_R1215_U171;
  assign new_P2_R1215_U128 = new_P2_R1215_U250 & new_P2_R1215_U8;
  assign new_P2_R1215_U129 = new_P2_R1215_U248 & new_P2_R1215_U172;
  assign new_P2_R1215_U130 = new_P2_R1215_U268 & new_P2_R1215_U267;
  assign new_P2_R1215_U131 = new_P2_R1215_U10 & new_P2_R1215_U282;
  assign new_P2_R1215_U132 = new_P2_R1215_U285 & new_P2_R1215_U280;
  assign new_P2_R1215_U133 = new_P2_R1215_U301 & new_P2_R1215_U298;
  assign new_P2_R1215_U134 = new_P2_R1215_U368 & new_P2_R1215_U302;
  assign new_P2_R1215_U135 = new_P2_R1215_U160 & new_P2_R1215_U278;
  assign new_P2_R1215_U136 = new_P2_R1215_U81 & new_P2_R1215_U455 & new_P2_R1215_U454;
  assign new_P2_R1215_U137 = new_P2_R1215_U325 & new_P2_R1215_U10;
  assign new_P2_R1215_U138 = new_P2_R1215_U60 & new_P2_R1215_U469 & new_P2_R1215_U468;
  assign new_P2_R1215_U139 = new_P2_R1215_U334 & new_P2_R1215_U9;
  assign new_P2_R1215_U140 = new_P2_R1215_U172 & new_P2_R1215_U490 & new_P2_R1215_U489;
  assign new_P2_R1215_U141 = new_P2_R1215_U343 & new_P2_R1215_U8;
  assign new_P2_R1215_U142 = new_P2_R1215_U171 & new_P2_R1215_U502 & new_P2_R1215_U501;
  assign new_P2_R1215_U143 = new_P2_R1215_U350 & new_P2_R1215_U7;
  assign new_P2_R1215_U144 = ~new_P2_R1215_U119 | ~new_P2_R1215_U202;
  assign new_P2_R1215_U145 = ~new_P2_R1215_U217 | ~new_P2_R1215_U229;
  assign new_P2_R1215_U146 = ~new_P2_U3057;
  assign new_P2_R1215_U147 = ~new_P2_U3960;
  assign new_P2_R1215_U148 = new_P2_R1215_U403 & new_P2_R1215_U402;
  assign new_P2_R1215_U149 = ~new_P2_R1215_U364 | ~new_P2_R1215_U304 | ~new_P2_R1215_U169;
  assign new_P2_R1215_U150 = new_P2_R1215_U410 & new_P2_R1215_U409;
  assign new_P2_R1215_U151 = ~new_P2_R1215_U134 | ~new_P2_R1215_U370 | ~new_P2_R1215_U369;
  assign new_P2_R1215_U152 = new_P2_R1215_U417 & new_P2_R1215_U416;
  assign new_P2_R1215_U153 = ~new_P2_R1215_U87 | ~new_P2_R1215_U365 | ~new_P2_R1215_U299;
  assign new_P2_R1215_U154 = new_P2_R1215_U424 & new_P2_R1215_U423;
  assign new_P2_R1215_U155 = ~new_P2_R1215_U293 | ~new_P2_R1215_U292;
  assign new_P2_R1215_U156 = new_P2_R1215_U436 & new_P2_R1215_U435;
  assign new_P2_R1215_U157 = ~new_P2_R1215_U289 | ~new_P2_R1215_U288;
  assign new_P2_R1215_U158 = new_P2_R1215_U443 & new_P2_R1215_U442;
  assign new_P2_R1215_U159 = ~new_P2_R1215_U132 | ~new_P2_R1215_U284;
  assign new_P2_R1215_U160 = new_P2_R1215_U450 & new_P2_R1215_U449;
  assign new_P2_R1215_U161 = ~new_P2_R1215_U44 | ~new_P2_R1215_U327;
  assign new_P2_R1215_U162 = ~new_P2_R1215_U130 | ~new_P2_R1215_U269;
  assign new_P2_R1215_U163 = new_P2_R1215_U476 & new_P2_R1215_U475;
  assign new_P2_R1215_U164 = ~new_P2_R1215_U257 | ~new_P2_R1215_U256;
  assign new_P2_R1215_U165 = new_P2_R1215_U483 & new_P2_R1215_U482;
  assign new_P2_R1215_U166 = ~new_P2_R1215_U253 | ~new_P2_R1215_U252;
  assign new_P2_R1215_U167 = ~new_P2_R1215_U243 | ~new_P2_R1215_U242;
  assign new_P2_R1215_U168 = ~new_P2_R1215_U367 | ~new_P2_R1215_U366;
  assign new_P2_R1215_U169 = ~new_P2_U3056 | ~new_P2_R1215_U151;
  assign new_P2_R1215_U170 = ~new_P2_R1215_U35;
  assign new_P2_R1215_U171 = ~new_P2_U3456 | ~new_P2_U3085;
  assign new_P2_R1215_U172 = ~new_P2_U3074 | ~new_P2_U3465;
  assign new_P2_R1215_U173 = ~new_P2_U3060 | ~new_P2_U3952;
  assign new_P2_R1215_U174 = ~new_P2_R1215_U69;
  assign new_P2_R1215_U175 = ~new_P2_R1215_U78;
  assign new_P2_R1215_U176 = ~new_P2_U3067 | ~new_P2_U3953;
  assign new_P2_R1215_U177 = ~new_P2_R1215_U62;
  assign new_P2_R1215_U178 = new_P2_U3069 | new_P2_U3444;
  assign new_P2_R1215_U179 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1215_U180 = new_P2_U3438 | new_P2_U3066;
  assign new_P2_R1215_U181 = new_P2_U3435 | new_P2_U3070;
  assign new_P2_R1215_U182 = ~new_P2_R1215_U32;
  assign new_P2_R1215_U183 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1215_U184 = ~new_P2_R1215_U43;
  assign new_P2_R1215_U185 = ~new_P2_R1215_U44;
  assign new_P2_R1215_U186 = ~new_P2_R1215_U43 | ~new_P2_R1215_U44;
  assign new_P2_R1215_U187 = ~new_P2_R1215_U116 | ~new_P2_R1215_U180;
  assign new_P2_R1215_U188 = ~new_P2_R1215_U5 | ~new_P2_R1215_U186;
  assign new_P2_R1215_U189 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1215_U190 = ~new_P2_R1215_U117 | ~new_P2_R1215_U188;
  assign new_P2_R1215_U191 = ~new_P2_R1215_U36 | ~new_P2_R1215_U35;
  assign new_P2_R1215_U192 = ~new_P2_U3069 | ~new_P2_R1215_U191;
  assign new_P2_R1215_U193 = ~new_P2_R1215_U4 | ~new_P2_R1215_U190;
  assign new_P2_R1215_U194 = ~new_P2_U3444 | ~new_P2_R1215_U170;
  assign new_P2_R1215_U195 = ~new_P2_R1215_U42;
  assign new_P2_R1215_U196 = new_P2_U3072 | new_P2_U3450;
  assign new_P2_R1215_U197 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1215_U198 = ~new_P2_R1215_U23;
  assign new_P2_R1215_U199 = ~new_P2_R1215_U24 | ~new_P2_R1215_U23;
  assign new_P2_R1215_U200 = ~new_P2_U3072 | ~new_P2_R1215_U199;
  assign new_P2_R1215_U201 = ~new_P2_U3450 | ~new_P2_R1215_U198;
  assign new_P2_R1215_U202 = ~new_P2_R1215_U6 | ~new_P2_R1215_U42;
  assign new_P2_R1215_U203 = ~new_P2_R1215_U144;
  assign new_P2_R1215_U204 = new_P2_U3453 | new_P2_U3086;
  assign new_P2_R1215_U205 = ~new_P2_R1215_U204 | ~new_P2_R1215_U144;
  assign new_P2_R1215_U206 = ~new_P2_R1215_U41;
  assign new_P2_R1215_U207 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1215_U208 = new_P2_U3447 | new_P2_U3073;
  assign new_P2_R1215_U209 = ~new_P2_R1215_U208 | ~new_P2_R1215_U42;
  assign new_P2_R1215_U210 = ~new_P2_R1215_U120 | ~new_P2_R1215_U209;
  assign new_P2_R1215_U211 = ~new_P2_R1215_U195 | ~new_P2_R1215_U23;
  assign new_P2_R1215_U212 = ~new_P2_U3450 | ~new_P2_U3072;
  assign new_P2_R1215_U213 = ~new_P2_R1215_U121 | ~new_P2_R1215_U211;
  assign new_P2_R1215_U214 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1215_U215 = ~new_P2_R1215_U185 | ~new_P2_R1215_U181;
  assign new_P2_R1215_U216 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1215_U217 = ~new_P2_R1215_U46;
  assign new_P2_R1215_U218 = ~new_P2_R1215_U184 | ~new_P2_R1215_U5;
  assign new_P2_R1215_U219 = ~new_P2_R1215_U46 | ~new_P2_R1215_U180;
  assign new_P2_R1215_U220 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1215_U221 = ~new_P2_R1215_U45;
  assign new_P2_R1215_U222 = new_P2_U3441 | new_P2_U3062;
  assign new_P2_R1215_U223 = ~new_P2_R1215_U222 | ~new_P2_R1215_U45;
  assign new_P2_R1215_U224 = ~new_P2_R1215_U123 | ~new_P2_R1215_U223;
  assign new_P2_R1215_U225 = ~new_P2_R1215_U221 | ~new_P2_R1215_U35;
  assign new_P2_R1215_U226 = ~new_P2_U3444 | ~new_P2_U3069;
  assign new_P2_R1215_U227 = ~new_P2_R1215_U124 | ~new_P2_R1215_U225;
  assign new_P2_R1215_U228 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1215_U229 = ~new_P2_R1215_U184 | ~new_P2_R1215_U181;
  assign new_P2_R1215_U230 = ~new_P2_R1215_U145;
  assign new_P2_R1215_U231 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1215_U232 = ~new_P2_R1215_U43 | ~new_P2_R1215_U44 | ~new_P2_R1215_U401 | ~new_P2_R1215_U400;
  assign new_P2_R1215_U233 = ~new_P2_R1215_U44 | ~new_P2_R1215_U43;
  assign new_P2_R1215_U234 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1215_U235 = ~new_P2_R1215_U125 | ~new_P2_R1215_U233;
  assign new_P2_R1215_U236 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1215_U237 = new_P2_U3064 | new_P2_U3459;
  assign new_P2_R1215_U238 = ~new_P2_R1215_U177 | ~new_P2_R1215_U7;
  assign new_P2_R1215_U239 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1215_U240 = ~new_P2_R1215_U127 | ~new_P2_R1215_U238;
  assign new_P2_R1215_U241 = new_P2_U3459 | new_P2_U3064;
  assign new_P2_R1215_U242 = ~new_P2_R1215_U126 | ~new_P2_R1215_U144;
  assign new_P2_R1215_U243 = ~new_P2_R1215_U241 | ~new_P2_R1215_U240;
  assign new_P2_R1215_U244 = ~new_P2_R1215_U167;
  assign new_P2_R1215_U245 = new_P2_U3082 | new_P2_U3468;
  assign new_P2_R1215_U246 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1215_U247 = ~new_P2_R1215_U174 | ~new_P2_R1215_U8;
  assign new_P2_R1215_U248 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1215_U249 = ~new_P2_R1215_U129 | ~new_P2_R1215_U247;
  assign new_P2_R1215_U250 = new_P2_U3462 | new_P2_U3065;
  assign new_P2_R1215_U251 = new_P2_U3468 | new_P2_U3082;
  assign new_P2_R1215_U252 = ~new_P2_R1215_U128 | ~new_P2_R1215_U167;
  assign new_P2_R1215_U253 = ~new_P2_R1215_U251 | ~new_P2_R1215_U249;
  assign new_P2_R1215_U254 = ~new_P2_R1215_U166;
  assign new_P2_R1215_U255 = new_P2_U3471 | new_P2_U3081;
  assign new_P2_R1215_U256 = ~new_P2_R1215_U255 | ~new_P2_R1215_U166;
  assign new_P2_R1215_U257 = ~new_P2_U3081 | ~new_P2_U3471;
  assign new_P2_R1215_U258 = ~new_P2_R1215_U164;
  assign new_P2_R1215_U259 = new_P2_U3474 | new_P2_U3076;
  assign new_P2_R1215_U260 = ~new_P2_R1215_U259 | ~new_P2_R1215_U164;
  assign new_P2_R1215_U261 = ~new_P2_U3076 | ~new_P2_U3474;
  assign new_P2_R1215_U262 = ~new_P2_R1215_U93;
  assign new_P2_R1215_U263 = new_P2_U3071 | new_P2_U3480;
  assign new_P2_R1215_U264 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1215_U265 = ~new_P2_R1215_U60;
  assign new_P2_R1215_U266 = ~new_P2_R1215_U61 | ~new_P2_R1215_U60;
  assign new_P2_R1215_U267 = ~new_P2_U3071 | ~new_P2_R1215_U266;
  assign new_P2_R1215_U268 = ~new_P2_U3480 | ~new_P2_R1215_U265;
  assign new_P2_R1215_U269 = ~new_P2_R1215_U9 | ~new_P2_R1215_U93;
  assign new_P2_R1215_U270 = ~new_P2_R1215_U162;
  assign new_P2_R1215_U271 = new_P2_U3078 | new_P2_U3957;
  assign new_P2_R1215_U272 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1215_U273 = new_P2_U3077 | new_P2_U3956;
  assign new_P2_R1215_U274 = ~new_P2_R1215_U81;
  assign new_P2_R1215_U275 = ~new_P2_U3957 | ~new_P2_R1215_U274;
  assign new_P2_R1215_U276 = ~new_P2_R1215_U275 | ~new_P2_R1215_U91;
  assign new_P2_R1215_U277 = ~new_P2_R1215_U81 | ~new_P2_R1215_U82;
  assign new_P2_R1215_U278 = ~new_P2_R1215_U277 | ~new_P2_R1215_U276;
  assign new_P2_R1215_U279 = ~new_P2_R1215_U175 | ~new_P2_R1215_U10;
  assign new_P2_R1215_U280 = ~new_P2_U3077 | ~new_P2_U3956;
  assign new_P2_R1215_U281 = ~new_P2_R1215_U278 | ~new_P2_R1215_U279;
  assign new_P2_R1215_U282 = new_P2_U3483 | new_P2_U3084;
  assign new_P2_R1215_U283 = new_P2_U3956 | new_P2_U3077;
  assign new_P2_R1215_U284 = ~new_P2_R1215_U131 | ~new_P2_R1215_U273 | ~new_P2_R1215_U162;
  assign new_P2_R1215_U285 = ~new_P2_R1215_U283 | ~new_P2_R1215_U281;
  assign new_P2_R1215_U286 = ~new_P2_R1215_U159;
  assign new_P2_R1215_U287 = new_P2_U3955 | new_P2_U3063;
  assign new_P2_R1215_U288 = ~new_P2_R1215_U287 | ~new_P2_R1215_U159;
  assign new_P2_R1215_U289 = ~new_P2_U3063 | ~new_P2_U3955;
  assign new_P2_R1215_U290 = ~new_P2_R1215_U157;
  assign new_P2_R1215_U291 = new_P2_U3954 | new_P2_U3068;
  assign new_P2_R1215_U292 = ~new_P2_R1215_U291 | ~new_P2_R1215_U157;
  assign new_P2_R1215_U293 = ~new_P2_U3068 | ~new_P2_U3954;
  assign new_P2_R1215_U294 = ~new_P2_R1215_U155;
  assign new_P2_R1215_U295 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1215_U296 = ~new_P2_R1215_U176 | ~new_P2_R1215_U173;
  assign new_P2_R1215_U297 = ~new_P2_R1215_U87;
  assign new_P2_R1215_U298 = new_P2_U3953 | new_P2_U3067;
  assign new_P2_R1215_U299 = ~new_P2_R1215_U168 | ~new_P2_R1215_U155 | ~new_P2_R1215_U298;
  assign new_P2_R1215_U300 = ~new_P2_R1215_U153;
  assign new_P2_R1215_U301 = new_P2_U3950 | new_P2_U3055;
  assign new_P2_R1215_U302 = ~new_P2_U3055 | ~new_P2_U3950;
  assign new_P2_R1215_U303 = ~new_P2_R1215_U151;
  assign new_P2_R1215_U304 = ~new_P2_U3949 | ~new_P2_R1215_U151;
  assign new_P2_R1215_U305 = ~new_P2_R1215_U149;
  assign new_P2_R1215_U306 = ~new_P2_R1215_U298 | ~new_P2_R1215_U155;
  assign new_P2_R1215_U307 = ~new_P2_R1215_U90;
  assign new_P2_R1215_U308 = new_P2_U3952 | new_P2_U3060;
  assign new_P2_R1215_U309 = ~new_P2_R1215_U308 | ~new_P2_R1215_U90;
  assign new_P2_R1215_U310 = ~new_P2_R1215_U154 | ~new_P2_R1215_U309 | ~new_P2_R1215_U173;
  assign new_P2_R1215_U311 = ~new_P2_R1215_U307 | ~new_P2_R1215_U173;
  assign new_P2_R1215_U312 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1215_U313 = ~new_P2_R1215_U168 | ~new_P2_R1215_U311 | ~new_P2_R1215_U312;
  assign new_P2_R1215_U314 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1215_U315 = ~new_P2_R1215_U282 | ~new_P2_R1215_U162;
  assign new_P2_R1215_U316 = ~new_P2_R1215_U92;
  assign new_P2_R1215_U317 = ~new_P2_R1215_U10 | ~new_P2_R1215_U92;
  assign new_P2_R1215_U318 = ~new_P2_R1215_U135 | ~new_P2_R1215_U317;
  assign new_P2_R1215_U319 = ~new_P2_R1215_U317 | ~new_P2_R1215_U278;
  assign new_P2_R1215_U320 = ~new_P2_R1215_U453 | ~new_P2_R1215_U319;
  assign new_P2_R1215_U321 = new_P2_U3485 | new_P2_U3083;
  assign new_P2_R1215_U322 = ~new_P2_R1215_U321 | ~new_P2_R1215_U92;
  assign new_P2_R1215_U323 = ~new_P2_R1215_U136 | ~new_P2_R1215_U322;
  assign new_P2_R1215_U324 = ~new_P2_R1215_U316 | ~new_P2_R1215_U81;
  assign new_P2_R1215_U325 = ~new_P2_U3078 | ~new_P2_U3957;
  assign new_P2_R1215_U326 = ~new_P2_R1215_U137 | ~new_P2_R1215_U324;
  assign new_P2_R1215_U327 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1215_U328 = ~new_P2_R1215_U161;
  assign new_P2_R1215_U329 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1215_U330 = new_P2_U3477 | new_P2_U3075;
  assign new_P2_R1215_U331 = ~new_P2_R1215_U330 | ~new_P2_R1215_U93;
  assign new_P2_R1215_U332 = ~new_P2_R1215_U138 | ~new_P2_R1215_U331;
  assign new_P2_R1215_U333 = ~new_P2_R1215_U262 | ~new_P2_R1215_U60;
  assign new_P2_R1215_U334 = ~new_P2_U3480 | ~new_P2_U3071;
  assign new_P2_R1215_U335 = ~new_P2_R1215_U139 | ~new_P2_R1215_U333;
  assign new_P2_R1215_U336 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1215_U337 = ~new_P2_R1215_U250 | ~new_P2_R1215_U167;
  assign new_P2_R1215_U338 = ~new_P2_R1215_U94;
  assign new_P2_R1215_U339 = new_P2_U3465 | new_P2_U3074;
  assign new_P2_R1215_U340 = ~new_P2_R1215_U339 | ~new_P2_R1215_U94;
  assign new_P2_R1215_U341 = ~new_P2_R1215_U140 | ~new_P2_R1215_U340;
  assign new_P2_R1215_U342 = ~new_P2_R1215_U338 | ~new_P2_R1215_U172;
  assign new_P2_R1215_U343 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1215_U344 = ~new_P2_R1215_U141 | ~new_P2_R1215_U342;
  assign new_P2_R1215_U345 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1215_U346 = new_P2_U3456 | new_P2_U3085;
  assign new_P2_R1215_U347 = ~new_P2_R1215_U346 | ~new_P2_R1215_U41;
  assign new_P2_R1215_U348 = ~new_P2_R1215_U142 | ~new_P2_R1215_U347;
  assign new_P2_R1215_U349 = ~new_P2_R1215_U206 | ~new_P2_R1215_U171;
  assign new_P2_R1215_U350 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1215_U351 = ~new_P2_R1215_U143 | ~new_P2_R1215_U349;
  assign new_P2_R1215_U352 = ~new_P2_R1215_U207 | ~new_P2_R1215_U171;
  assign new_P2_R1215_U353 = ~new_P2_R1215_U204 | ~new_P2_R1215_U62;
  assign new_P2_R1215_U354 = ~new_P2_R1215_U214 | ~new_P2_R1215_U23;
  assign new_P2_R1215_U355 = ~new_P2_R1215_U228 | ~new_P2_R1215_U35;
  assign new_P2_R1215_U356 = ~new_P2_R1215_U231 | ~new_P2_R1215_U180;
  assign new_P2_R1215_U357 = ~new_P2_R1215_U314 | ~new_P2_R1215_U173;
  assign new_P2_R1215_U358 = ~new_P2_R1215_U298 | ~new_P2_R1215_U176;
  assign new_P2_R1215_U359 = ~new_P2_R1215_U329 | ~new_P2_R1215_U81;
  assign new_P2_R1215_U360 = ~new_P2_R1215_U282 | ~new_P2_R1215_U78;
  assign new_P2_R1215_U361 = ~new_P2_R1215_U336 | ~new_P2_R1215_U60;
  assign new_P2_R1215_U362 = ~new_P2_R1215_U345 | ~new_P2_R1215_U172;
  assign new_P2_R1215_U363 = ~new_P2_R1215_U250 | ~new_P2_R1215_U69;
  assign new_P2_R1215_U364 = ~new_P2_U3949 | ~new_P2_U3056;
  assign new_P2_R1215_U365 = ~new_P2_R1215_U296 | ~new_P2_R1215_U168;
  assign new_P2_R1215_U366 = ~new_P2_U3059 | ~new_P2_R1215_U295;
  assign new_P2_R1215_U367 = ~new_P2_U3951 | ~new_P2_R1215_U295;
  assign new_P2_R1215_U368 = ~new_P2_R1215_U301 | ~new_P2_R1215_U296 | ~new_P2_R1215_U168;
  assign new_P2_R1215_U369 = ~new_P2_R1215_U133 | ~new_P2_R1215_U155 | ~new_P2_R1215_U168;
  assign new_P2_R1215_U370 = ~new_P2_R1215_U297 | ~new_P2_R1215_U301;
  assign new_P2_R1215_U371 = ~new_P2_U3085 | ~new_P2_R1215_U40;
  assign new_P2_R1215_U372 = ~new_P2_U3456 | ~new_P2_R1215_U39;
  assign new_P2_R1215_U373 = ~new_P2_R1215_U372 | ~new_P2_R1215_U371;
  assign new_P2_R1215_U374 = ~new_P2_R1215_U352 | ~new_P2_R1215_U41;
  assign new_P2_R1215_U375 = ~new_P2_R1215_U373 | ~new_P2_R1215_U206;
  assign new_P2_R1215_U376 = ~new_P2_U3086 | ~new_P2_R1215_U37;
  assign new_P2_R1215_U377 = ~new_P2_U3453 | ~new_P2_R1215_U38;
  assign new_P2_R1215_U378 = ~new_P2_R1215_U377 | ~new_P2_R1215_U376;
  assign new_P2_R1215_U379 = ~new_P2_R1215_U353 | ~new_P2_R1215_U144;
  assign new_P2_R1215_U380 = ~new_P2_R1215_U203 | ~new_P2_R1215_U378;
  assign new_P2_R1215_U381 = ~new_P2_U3072 | ~new_P2_R1215_U24;
  assign new_P2_R1215_U382 = ~new_P2_U3450 | ~new_P2_R1215_U22;
  assign new_P2_R1215_U383 = ~new_P2_U3073 | ~new_P2_R1215_U20;
  assign new_P2_R1215_U384 = ~new_P2_U3447 | ~new_P2_R1215_U21;
  assign new_P2_R1215_U385 = ~new_P2_R1215_U384 | ~new_P2_R1215_U383;
  assign new_P2_R1215_U386 = ~new_P2_R1215_U354 | ~new_P2_R1215_U42;
  assign new_P2_R1215_U387 = ~new_P2_R1215_U385 | ~new_P2_R1215_U195;
  assign new_P2_R1215_U388 = ~new_P2_U3069 | ~new_P2_R1215_U36;
  assign new_P2_R1215_U389 = ~new_P2_U3444 | ~new_P2_R1215_U27;
  assign new_P2_R1215_U390 = ~new_P2_U3062 | ~new_P2_R1215_U25;
  assign new_P2_R1215_U391 = ~new_P2_U3441 | ~new_P2_R1215_U26;
  assign new_P2_R1215_U392 = ~new_P2_R1215_U391 | ~new_P2_R1215_U390;
  assign new_P2_R1215_U393 = ~new_P2_R1215_U355 | ~new_P2_R1215_U45;
  assign new_P2_R1215_U394 = ~new_P2_R1215_U392 | ~new_P2_R1215_U221;
  assign new_P2_R1215_U395 = ~new_P2_U3066 | ~new_P2_R1215_U33;
  assign new_P2_R1215_U396 = ~new_P2_U3438 | ~new_P2_R1215_U34;
  assign new_P2_R1215_U397 = ~new_P2_R1215_U396 | ~new_P2_R1215_U395;
  assign new_P2_R1215_U398 = ~new_P2_R1215_U356 | ~new_P2_R1215_U145;
  assign new_P2_R1215_U399 = ~new_P2_R1215_U230 | ~new_P2_R1215_U397;
  assign new_P2_R1215_U400 = ~new_P2_U3070 | ~new_P2_R1215_U28;
  assign new_P2_R1215_U401 = ~new_P2_U3435 | ~new_P2_R1215_U29;
  assign new_P2_R1215_U402 = ~new_P2_U3057 | ~new_P2_R1215_U147;
  assign new_P2_R1215_U403 = ~new_P2_U3960 | ~new_P2_R1215_U146;
  assign new_P2_R1215_U404 = ~new_P2_U3057 | ~new_P2_R1215_U147;
  assign new_P2_R1215_U405 = ~new_P2_U3960 | ~new_P2_R1215_U146;
  assign new_P2_R1215_U406 = ~new_P2_R1215_U405 | ~new_P2_R1215_U404;
  assign new_P2_R1215_U407 = ~new_P2_R1215_U148 | ~new_P2_R1215_U149;
  assign new_P2_R1215_U408 = ~new_P2_R1215_U305 | ~new_P2_R1215_U406;
  assign new_P2_R1215_U409 = ~new_P2_U3056 | ~new_P2_R1215_U89;
  assign new_P2_R1215_U410 = ~new_P2_U3949 | ~new_P2_R1215_U88;
  assign new_P2_R1215_U411 = ~new_P2_U3056 | ~new_P2_R1215_U89;
  assign new_P2_R1215_U412 = ~new_P2_U3949 | ~new_P2_R1215_U88;
  assign new_P2_R1215_U413 = ~new_P2_R1215_U412 | ~new_P2_R1215_U411;
  assign new_P2_R1215_U414 = ~new_P2_R1215_U150 | ~new_P2_R1215_U151;
  assign new_P2_R1215_U415 = ~new_P2_R1215_U303 | ~new_P2_R1215_U413;
  assign new_P2_R1215_U416 = ~new_P2_U3055 | ~new_P2_R1215_U47;
  assign new_P2_R1215_U417 = ~new_P2_U3950 | ~new_P2_R1215_U48;
  assign new_P2_R1215_U418 = ~new_P2_U3055 | ~new_P2_R1215_U47;
  assign new_P2_R1215_U419 = ~new_P2_U3950 | ~new_P2_R1215_U48;
  assign new_P2_R1215_U420 = ~new_P2_R1215_U419 | ~new_P2_R1215_U418;
  assign new_P2_R1215_U421 = ~new_P2_R1215_U152 | ~new_P2_R1215_U153;
  assign new_P2_R1215_U422 = ~new_P2_R1215_U300 | ~new_P2_R1215_U420;
  assign new_P2_R1215_U423 = ~new_P2_U3059 | ~new_P2_R1215_U50;
  assign new_P2_R1215_U424 = ~new_P2_U3951 | ~new_P2_R1215_U49;
  assign new_P2_R1215_U425 = ~new_P2_U3060 | ~new_P2_R1215_U51;
  assign new_P2_R1215_U426 = ~new_P2_U3952 | ~new_P2_R1215_U52;
  assign new_P2_R1215_U427 = ~new_P2_R1215_U426 | ~new_P2_R1215_U425;
  assign new_P2_R1215_U428 = ~new_P2_R1215_U357 | ~new_P2_R1215_U90;
  assign new_P2_R1215_U429 = ~new_P2_R1215_U427 | ~new_P2_R1215_U307;
  assign new_P2_R1215_U430 = ~new_P2_U3067 | ~new_P2_R1215_U53;
  assign new_P2_R1215_U431 = ~new_P2_U3953 | ~new_P2_R1215_U54;
  assign new_P2_R1215_U432 = ~new_P2_R1215_U431 | ~new_P2_R1215_U430;
  assign new_P2_R1215_U433 = ~new_P2_R1215_U358 | ~new_P2_R1215_U155;
  assign new_P2_R1215_U434 = ~new_P2_R1215_U294 | ~new_P2_R1215_U432;
  assign new_P2_R1215_U435 = ~new_P2_U3068 | ~new_P2_R1215_U85;
  assign new_P2_R1215_U436 = ~new_P2_U3954 | ~new_P2_R1215_U86;
  assign new_P2_R1215_U437 = ~new_P2_U3068 | ~new_P2_R1215_U85;
  assign new_P2_R1215_U438 = ~new_P2_U3954 | ~new_P2_R1215_U86;
  assign new_P2_R1215_U439 = ~new_P2_R1215_U438 | ~new_P2_R1215_U437;
  assign new_P2_R1215_U440 = ~new_P2_R1215_U156 | ~new_P2_R1215_U157;
  assign new_P2_R1215_U441 = ~new_P2_R1215_U290 | ~new_P2_R1215_U439;
  assign new_P2_R1215_U442 = ~new_P2_U3063 | ~new_P2_R1215_U83;
  assign new_P2_R1215_U443 = ~new_P2_U3955 | ~new_P2_R1215_U84;
  assign new_P2_R1215_U444 = ~new_P2_U3063 | ~new_P2_R1215_U83;
  assign new_P2_R1215_U445 = ~new_P2_U3955 | ~new_P2_R1215_U84;
  assign new_P2_R1215_U446 = ~new_P2_R1215_U445 | ~new_P2_R1215_U444;
  assign new_P2_R1215_U447 = ~new_P2_R1215_U158 | ~new_P2_R1215_U159;
  assign new_P2_R1215_U448 = ~new_P2_R1215_U286 | ~new_P2_R1215_U446;
  assign new_P2_R1215_U449 = ~new_P2_U3077 | ~new_P2_R1215_U55;
  assign new_P2_R1215_U450 = ~new_P2_U3956 | ~new_P2_R1215_U56;
  assign new_P2_R1215_U451 = ~new_P2_U3077 | ~new_P2_R1215_U55;
  assign new_P2_R1215_U452 = ~new_P2_U3956 | ~new_P2_R1215_U56;
  assign new_P2_R1215_U453 = ~new_P2_R1215_U452 | ~new_P2_R1215_U451;
  assign new_P2_R1215_U454 = ~new_P2_U3078 | ~new_P2_R1215_U82;
  assign new_P2_R1215_U455 = ~new_P2_U3957 | ~new_P2_R1215_U91;
  assign new_P2_R1215_U456 = ~new_P2_R1215_U182 | ~new_P2_R1215_U161;
  assign new_P2_R1215_U457 = ~new_P2_R1215_U328 | ~new_P2_R1215_U32;
  assign new_P2_R1215_U458 = ~new_P2_U3083 | ~new_P2_R1215_U79;
  assign new_P2_R1215_U459 = ~new_P2_U3485 | ~new_P2_R1215_U80;
  assign new_P2_R1215_U460 = ~new_P2_R1215_U459 | ~new_P2_R1215_U458;
  assign new_P2_R1215_U461 = ~new_P2_R1215_U359 | ~new_P2_R1215_U92;
  assign new_P2_R1215_U462 = ~new_P2_R1215_U460 | ~new_P2_R1215_U316;
  assign new_P2_R1215_U463 = ~new_P2_U3084 | ~new_P2_R1215_U76;
  assign new_P2_R1215_U464 = ~new_P2_U3483 | ~new_P2_R1215_U77;
  assign new_P2_R1215_U465 = ~new_P2_R1215_U464 | ~new_P2_R1215_U463;
  assign new_P2_R1215_U466 = ~new_P2_R1215_U360 | ~new_P2_R1215_U162;
  assign new_P2_R1215_U467 = ~new_P2_R1215_U270 | ~new_P2_R1215_U465;
  assign new_P2_R1215_U468 = ~new_P2_U3071 | ~new_P2_R1215_U61;
  assign new_P2_R1215_U469 = ~new_P2_U3480 | ~new_P2_R1215_U59;
  assign new_P2_R1215_U470 = ~new_P2_U3075 | ~new_P2_R1215_U57;
  assign new_P2_R1215_U471 = ~new_P2_U3477 | ~new_P2_R1215_U58;
  assign new_P2_R1215_U472 = ~new_P2_R1215_U471 | ~new_P2_R1215_U470;
  assign new_P2_R1215_U473 = ~new_P2_R1215_U361 | ~new_P2_R1215_U93;
  assign new_P2_R1215_U474 = ~new_P2_R1215_U472 | ~new_P2_R1215_U262;
  assign new_P2_R1215_U475 = ~new_P2_U3076 | ~new_P2_R1215_U74;
  assign new_P2_R1215_U476 = ~new_P2_U3474 | ~new_P2_R1215_U75;
  assign new_P2_R1215_U477 = ~new_P2_U3076 | ~new_P2_R1215_U74;
  assign new_P2_R1215_U478 = ~new_P2_U3474 | ~new_P2_R1215_U75;
  assign new_P2_R1215_U479 = ~new_P2_R1215_U478 | ~new_P2_R1215_U477;
  assign new_P2_R1215_U480 = ~new_P2_R1215_U163 | ~new_P2_R1215_U164;
  assign new_P2_R1215_U481 = ~new_P2_R1215_U258 | ~new_P2_R1215_U479;
  assign new_P2_R1215_U482 = ~new_P2_U3081 | ~new_P2_R1215_U72;
  assign new_P2_R1215_U483 = ~new_P2_U3471 | ~new_P2_R1215_U73;
  assign new_P2_R1215_U484 = ~new_P2_U3081 | ~new_P2_R1215_U72;
  assign new_P2_R1215_U485 = ~new_P2_U3471 | ~new_P2_R1215_U73;
  assign new_P2_R1215_U486 = ~new_P2_R1215_U485 | ~new_P2_R1215_U484;
  assign new_P2_R1215_U487 = ~new_P2_R1215_U165 | ~new_P2_R1215_U166;
  assign new_P2_R1215_U488 = ~new_P2_R1215_U254 | ~new_P2_R1215_U486;
  assign new_P2_R1215_U489 = ~new_P2_U3082 | ~new_P2_R1215_U70;
  assign new_P2_R1215_U490 = ~new_P2_U3468 | ~new_P2_R1215_U71;
  assign new_P2_R1215_U491 = ~new_P2_U3074 | ~new_P2_R1215_U65;
  assign new_P2_R1215_U492 = ~new_P2_U3465 | ~new_P2_R1215_U66;
  assign new_P2_R1215_U493 = ~new_P2_R1215_U492 | ~new_P2_R1215_U491;
  assign new_P2_R1215_U494 = ~new_P2_R1215_U362 | ~new_P2_R1215_U94;
  assign new_P2_R1215_U495 = ~new_P2_R1215_U493 | ~new_P2_R1215_U338;
  assign new_P2_R1215_U496 = ~new_P2_U3065 | ~new_P2_R1215_U67;
  assign new_P2_R1215_U497 = ~new_P2_U3462 | ~new_P2_R1215_U68;
  assign new_P2_R1215_U498 = ~new_P2_R1215_U497 | ~new_P2_R1215_U496;
  assign new_P2_R1215_U499 = ~new_P2_R1215_U363 | ~new_P2_R1215_U167;
  assign new_P2_R1215_U500 = ~new_P2_R1215_U244 | ~new_P2_R1215_U498;
  assign new_P2_R1215_U501 = ~new_P2_U3064 | ~new_P2_R1215_U63;
  assign new_P2_R1215_U502 = ~new_P2_U3459 | ~new_P2_R1215_U64;
  assign new_P2_R1215_U503 = ~new_P2_U3079 | ~new_P2_R1215_U30;
  assign new_P2_R1215_U504 = ~new_P2_U3427 | ~new_P2_R1215_U31;
  assign new_P2_R1164_U4 = new_P2_R1164_U179 & new_P2_R1164_U178;
  assign new_P2_R1164_U5 = new_P2_R1164_U197 & new_P2_R1164_U196;
  assign new_P2_R1164_U6 = new_P2_R1164_U237 & new_P2_R1164_U236;
  assign new_P2_R1164_U7 = new_P2_R1164_U246 & new_P2_R1164_U245;
  assign new_P2_R1164_U8 = new_P2_R1164_U264 & new_P2_R1164_U263;
  assign new_P2_R1164_U9 = new_P2_R1164_U272 & new_P2_R1164_U271;
  assign new_P2_R1164_U10 = new_P2_R1164_U351 & new_P2_R1164_U348;
  assign new_P2_R1164_U11 = new_P2_R1164_U344 & new_P2_R1164_U341;
  assign new_P2_R1164_U12 = new_P2_R1164_U335 & new_P2_R1164_U332;
  assign new_P2_R1164_U13 = new_P2_R1164_U326 & new_P2_R1164_U323;
  assign new_P2_R1164_U14 = new_P2_R1164_U320 & new_P2_R1164_U318;
  assign new_P2_R1164_U15 = new_P2_R1164_U313 & new_P2_R1164_U310;
  assign new_P2_R1164_U16 = new_P2_R1164_U235 & new_P2_R1164_U232;
  assign new_P2_R1164_U17 = new_P2_R1164_U227 & new_P2_R1164_U224;
  assign new_P2_R1164_U18 = new_P2_R1164_U213 & new_P2_R1164_U210;
  assign new_P2_R1164_U19 = ~new_P2_U3447;
  assign new_P2_R1164_U20 = ~new_P2_U3073;
  assign new_P2_R1164_U21 = ~new_P2_U3072;
  assign new_P2_R1164_U22 = ~new_P2_U3073 | ~new_P2_U3447;
  assign new_P2_R1164_U23 = ~new_P2_U3450;
  assign new_P2_R1164_U24 = ~new_P2_U3441;
  assign new_P2_R1164_U25 = ~new_P2_U3062;
  assign new_P2_R1164_U26 = ~new_P2_U3069;
  assign new_P2_R1164_U27 = ~new_P2_U3435;
  assign new_P2_R1164_U28 = ~new_P2_U3070;
  assign new_P2_R1164_U29 = ~new_P2_U3427;
  assign new_P2_R1164_U30 = ~new_P2_U3079;
  assign new_P2_R1164_U31 = ~new_P2_U3079 | ~new_P2_U3427;
  assign new_P2_R1164_U32 = ~new_P2_U3438;
  assign new_P2_R1164_U33 = ~new_P2_U3066;
  assign new_P2_R1164_U34 = ~new_P2_U3062 | ~new_P2_U3441;
  assign new_P2_R1164_U35 = ~new_P2_U3444;
  assign new_P2_R1164_U36 = ~new_P2_U3453;
  assign new_P2_R1164_U37 = ~new_P2_U3086;
  assign new_P2_R1164_U38 = ~new_P2_U3085;
  assign new_P2_R1164_U39 = ~new_P2_U3456;
  assign new_P2_R1164_U40 = ~new_P2_R1164_U61 | ~new_P2_R1164_U205;
  assign new_P2_R1164_U41 = ~new_P2_R1164_U117 | ~new_P2_R1164_U193;
  assign new_P2_R1164_U42 = ~new_P2_R1164_U182 | ~new_P2_R1164_U183;
  assign new_P2_R1164_U43 = ~new_P2_U3432 | ~new_P2_U3080;
  assign new_P2_R1164_U44 = ~new_P2_R1164_U122 | ~new_P2_R1164_U219;
  assign new_P2_R1164_U45 = ~new_P2_R1164_U216 | ~new_P2_R1164_U215;
  assign new_P2_R1164_U46 = ~new_P2_U3950;
  assign new_P2_R1164_U47 = ~new_P2_U3055;
  assign new_P2_R1164_U48 = ~new_P2_U3059;
  assign new_P2_R1164_U49 = ~new_P2_U3951;
  assign new_P2_R1164_U50 = ~new_P2_U3952;
  assign new_P2_R1164_U51 = ~new_P2_U3060;
  assign new_P2_R1164_U52 = ~new_P2_U3953;
  assign new_P2_R1164_U53 = ~new_P2_U3067;
  assign new_P2_R1164_U54 = ~new_P2_U3956;
  assign new_P2_R1164_U55 = ~new_P2_U3077;
  assign new_P2_R1164_U56 = ~new_P2_U3477;
  assign new_P2_R1164_U57 = ~new_P2_U3075;
  assign new_P2_R1164_U58 = ~new_P2_U3071;
  assign new_P2_R1164_U59 = ~new_P2_U3075 | ~new_P2_U3477;
  assign new_P2_R1164_U60 = ~new_P2_U3480;
  assign new_P2_R1164_U61 = ~new_P2_U3086 | ~new_P2_U3453;
  assign new_P2_R1164_U62 = ~new_P2_U3459;
  assign new_P2_R1164_U63 = ~new_P2_U3064;
  assign new_P2_R1164_U64 = ~new_P2_U3465;
  assign new_P2_R1164_U65 = ~new_P2_U3074;
  assign new_P2_R1164_U66 = ~new_P2_U3462;
  assign new_P2_R1164_U67 = ~new_P2_U3065;
  assign new_P2_R1164_U68 = ~new_P2_U3065 | ~new_P2_U3462;
  assign new_P2_R1164_U69 = ~new_P2_U3468;
  assign new_P2_R1164_U70 = ~new_P2_U3082;
  assign new_P2_R1164_U71 = ~new_P2_U3471;
  assign new_P2_R1164_U72 = ~new_P2_U3081;
  assign new_P2_R1164_U73 = ~new_P2_U3474;
  assign new_P2_R1164_U74 = ~new_P2_U3076;
  assign new_P2_R1164_U75 = ~new_P2_U3483;
  assign new_P2_R1164_U76 = ~new_P2_U3084;
  assign new_P2_R1164_U77 = ~new_P2_U3084 | ~new_P2_U3483;
  assign new_P2_R1164_U78 = ~new_P2_U3485;
  assign new_P2_R1164_U79 = ~new_P2_U3083;
  assign new_P2_R1164_U80 = ~new_P2_U3083 | ~new_P2_U3485;
  assign new_P2_R1164_U81 = ~new_P2_U3957;
  assign new_P2_R1164_U82 = ~new_P2_U3955;
  assign new_P2_R1164_U83 = ~new_P2_U3063;
  assign new_P2_R1164_U84 = ~new_P2_U3954;
  assign new_P2_R1164_U85 = ~new_P2_U3068;
  assign new_P2_R1164_U86 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1164_U87 = ~new_P2_U3056;
  assign new_P2_R1164_U88 = ~new_P2_U3949;
  assign new_P2_R1164_U89 = ~new_P2_R1164_U306 | ~new_P2_R1164_U176;
  assign new_P2_R1164_U90 = ~new_P2_U3078;
  assign new_P2_R1164_U91 = ~new_P2_R1164_U77 | ~new_P2_R1164_U315;
  assign new_P2_R1164_U92 = ~new_P2_R1164_U261 | ~new_P2_R1164_U260;
  assign new_P2_R1164_U93 = ~new_P2_R1164_U68 | ~new_P2_R1164_U337;
  assign new_P2_R1164_U94 = ~new_P2_R1164_U457 | ~new_P2_R1164_U456;
  assign new_P2_R1164_U95 = ~new_P2_R1164_U504 | ~new_P2_R1164_U503;
  assign new_P2_R1164_U96 = ~new_P2_R1164_U375 | ~new_P2_R1164_U374;
  assign new_P2_R1164_U97 = ~new_P2_R1164_U380 | ~new_P2_R1164_U379;
  assign new_P2_R1164_U98 = ~new_P2_R1164_U387 | ~new_P2_R1164_U386;
  assign new_P2_R1164_U99 = ~new_P2_R1164_U394 | ~new_P2_R1164_U393;
  assign new_P2_R1164_U100 = ~new_P2_R1164_U399 | ~new_P2_R1164_U398;
  assign new_P2_R1164_U101 = ~new_P2_R1164_U408 | ~new_P2_R1164_U407;
  assign new_P2_R1164_U102 = ~new_P2_R1164_U415 | ~new_P2_R1164_U414;
  assign new_P2_R1164_U103 = ~new_P2_R1164_U422 | ~new_P2_R1164_U421;
  assign new_P2_R1164_U104 = ~new_P2_R1164_U429 | ~new_P2_R1164_U428;
  assign new_P2_R1164_U105 = ~new_P2_R1164_U434 | ~new_P2_R1164_U433;
  assign new_P2_R1164_U106 = ~new_P2_R1164_U441 | ~new_P2_R1164_U440;
  assign new_P2_R1164_U107 = ~new_P2_R1164_U448 | ~new_P2_R1164_U447;
  assign new_P2_R1164_U108 = ~new_P2_R1164_U462 | ~new_P2_R1164_U461;
  assign new_P2_R1164_U109 = ~new_P2_R1164_U467 | ~new_P2_R1164_U466;
  assign new_P2_R1164_U110 = ~new_P2_R1164_U474 | ~new_P2_R1164_U473;
  assign new_P2_R1164_U111 = ~new_P2_R1164_U481 | ~new_P2_R1164_U480;
  assign new_P2_R1164_U112 = ~new_P2_R1164_U488 | ~new_P2_R1164_U487;
  assign new_P2_R1164_U113 = ~new_P2_R1164_U495 | ~new_P2_R1164_U494;
  assign new_P2_R1164_U114 = ~new_P2_R1164_U500 | ~new_P2_R1164_U499;
  assign new_P2_R1164_U115 = new_P2_R1164_U189 & new_P2_R1164_U187;
  assign new_P2_R1164_U116 = new_P2_R1164_U4 & new_P2_R1164_U180;
  assign new_P2_R1164_U117 = new_P2_R1164_U194 & new_P2_R1164_U192;
  assign new_P2_R1164_U118 = new_P2_R1164_U201 & new_P2_R1164_U200;
  assign new_P2_R1164_U119 = new_P2_R1164_U22 & new_P2_R1164_U382 & new_P2_R1164_U381;
  assign new_P2_R1164_U120 = new_P2_R1164_U212 & new_P2_R1164_U5;
  assign new_P2_R1164_U121 = new_P2_R1164_U181 & new_P2_R1164_U180;
  assign new_P2_R1164_U122 = new_P2_R1164_U220 & new_P2_R1164_U218;
  assign new_P2_R1164_U123 = new_P2_R1164_U34 & new_P2_R1164_U389 & new_P2_R1164_U388;
  assign new_P2_R1164_U124 = new_P2_R1164_U226 & new_P2_R1164_U4;
  assign new_P2_R1164_U125 = new_P2_R1164_U234 & new_P2_R1164_U181;
  assign new_P2_R1164_U126 = new_P2_R1164_U204 & new_P2_R1164_U6;
  assign new_P2_R1164_U127 = new_P2_R1164_U239 & new_P2_R1164_U171;
  assign new_P2_R1164_U128 = new_P2_R1164_U250 & new_P2_R1164_U7;
  assign new_P2_R1164_U129 = new_P2_R1164_U248 & new_P2_R1164_U172;
  assign new_P2_R1164_U130 = new_P2_R1164_U268 & new_P2_R1164_U267;
  assign new_P2_R1164_U131 = new_P2_R1164_U9 & new_P2_R1164_U282;
  assign new_P2_R1164_U132 = new_P2_R1164_U285 & new_P2_R1164_U280;
  assign new_P2_R1164_U133 = new_P2_R1164_U301 & new_P2_R1164_U298;
  assign new_P2_R1164_U134 = new_P2_R1164_U368 & new_P2_R1164_U302;
  assign new_P2_R1164_U135 = new_P2_R1164_U160 & new_P2_R1164_U278;
  assign new_P2_R1164_U136 = new_P2_R1164_U80 & new_P2_R1164_U455 & new_P2_R1164_U454;
  assign new_P2_R1164_U137 = new_P2_R1164_U325 & new_P2_R1164_U9;
  assign new_P2_R1164_U138 = new_P2_R1164_U59 & new_P2_R1164_U469 & new_P2_R1164_U468;
  assign new_P2_R1164_U139 = new_P2_R1164_U334 & new_P2_R1164_U8;
  assign new_P2_R1164_U140 = new_P2_R1164_U172 & new_P2_R1164_U490 & new_P2_R1164_U489;
  assign new_P2_R1164_U141 = new_P2_R1164_U343 & new_P2_R1164_U7;
  assign new_P2_R1164_U142 = new_P2_R1164_U171 & new_P2_R1164_U502 & new_P2_R1164_U501;
  assign new_P2_R1164_U143 = new_P2_R1164_U350 & new_P2_R1164_U6;
  assign new_P2_R1164_U144 = ~new_P2_R1164_U118 | ~new_P2_R1164_U202;
  assign new_P2_R1164_U145 = ~new_P2_R1164_U217 | ~new_P2_R1164_U229;
  assign new_P2_R1164_U146 = ~new_P2_U3057;
  assign new_P2_R1164_U147 = ~new_P2_U3960;
  assign new_P2_R1164_U148 = new_P2_R1164_U403 & new_P2_R1164_U402;
  assign new_P2_R1164_U149 = ~new_P2_R1164_U364 | ~new_P2_R1164_U304 | ~new_P2_R1164_U169;
  assign new_P2_R1164_U150 = new_P2_R1164_U410 & new_P2_R1164_U409;
  assign new_P2_R1164_U151 = ~new_P2_R1164_U134 | ~new_P2_R1164_U370 | ~new_P2_R1164_U369;
  assign new_P2_R1164_U152 = new_P2_R1164_U417 & new_P2_R1164_U416;
  assign new_P2_R1164_U153 = ~new_P2_R1164_U86 | ~new_P2_R1164_U365 | ~new_P2_R1164_U299;
  assign new_P2_R1164_U154 = new_P2_R1164_U424 & new_P2_R1164_U423;
  assign new_P2_R1164_U155 = ~new_P2_R1164_U293 | ~new_P2_R1164_U292;
  assign new_P2_R1164_U156 = new_P2_R1164_U436 & new_P2_R1164_U435;
  assign new_P2_R1164_U157 = ~new_P2_R1164_U289 | ~new_P2_R1164_U288;
  assign new_P2_R1164_U158 = new_P2_R1164_U443 & new_P2_R1164_U442;
  assign new_P2_R1164_U159 = ~new_P2_R1164_U132 | ~new_P2_R1164_U284;
  assign new_P2_R1164_U160 = new_P2_R1164_U450 & new_P2_R1164_U449;
  assign new_P2_R1164_U161 = ~new_P2_R1164_U43 | ~new_P2_R1164_U327;
  assign new_P2_R1164_U162 = ~new_P2_R1164_U130 | ~new_P2_R1164_U269;
  assign new_P2_R1164_U163 = new_P2_R1164_U476 & new_P2_R1164_U475;
  assign new_P2_R1164_U164 = ~new_P2_R1164_U257 | ~new_P2_R1164_U256;
  assign new_P2_R1164_U165 = new_P2_R1164_U483 & new_P2_R1164_U482;
  assign new_P2_R1164_U166 = ~new_P2_R1164_U253 | ~new_P2_R1164_U252;
  assign new_P2_R1164_U167 = ~new_P2_R1164_U243 | ~new_P2_R1164_U242;
  assign new_P2_R1164_U168 = ~new_P2_R1164_U367 | ~new_P2_R1164_U366;
  assign new_P2_R1164_U169 = ~new_P2_U3056 | ~new_P2_R1164_U151;
  assign new_P2_R1164_U170 = ~new_P2_R1164_U34;
  assign new_P2_R1164_U171 = ~new_P2_U3456 | ~new_P2_U3085;
  assign new_P2_R1164_U172 = ~new_P2_U3074 | ~new_P2_U3465;
  assign new_P2_R1164_U173 = ~new_P2_U3060 | ~new_P2_U3952;
  assign new_P2_R1164_U174 = ~new_P2_R1164_U68;
  assign new_P2_R1164_U175 = ~new_P2_R1164_U77;
  assign new_P2_R1164_U176 = ~new_P2_U3067 | ~new_P2_U3953;
  assign new_P2_R1164_U177 = ~new_P2_R1164_U61;
  assign new_P2_R1164_U178 = new_P2_U3069 | new_P2_U3444;
  assign new_P2_R1164_U179 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1164_U180 = new_P2_U3438 | new_P2_U3066;
  assign new_P2_R1164_U181 = new_P2_U3435 | new_P2_U3070;
  assign new_P2_R1164_U182 = ~new_P2_R1164_U31;
  assign new_P2_R1164_U183 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1164_U184 = ~new_P2_R1164_U42;
  assign new_P2_R1164_U185 = ~new_P2_R1164_U43;
  assign new_P2_R1164_U186 = ~new_P2_R1164_U42 | ~new_P2_R1164_U43;
  assign new_P2_R1164_U187 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1164_U188 = ~new_P2_R1164_U186 | ~new_P2_R1164_U181;
  assign new_P2_R1164_U189 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1164_U190 = ~new_P2_R1164_U115 | ~new_P2_R1164_U188;
  assign new_P2_R1164_U191 = ~new_P2_R1164_U35 | ~new_P2_R1164_U34;
  assign new_P2_R1164_U192 = ~new_P2_U3069 | ~new_P2_R1164_U191;
  assign new_P2_R1164_U193 = ~new_P2_R1164_U116 | ~new_P2_R1164_U190;
  assign new_P2_R1164_U194 = ~new_P2_U3444 | ~new_P2_R1164_U170;
  assign new_P2_R1164_U195 = ~new_P2_R1164_U41;
  assign new_P2_R1164_U196 = new_P2_U3072 | new_P2_U3450;
  assign new_P2_R1164_U197 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1164_U198 = ~new_P2_R1164_U22;
  assign new_P2_R1164_U199 = ~new_P2_R1164_U23 | ~new_P2_R1164_U22;
  assign new_P2_R1164_U200 = ~new_P2_U3072 | ~new_P2_R1164_U199;
  assign new_P2_R1164_U201 = ~new_P2_U3450 | ~new_P2_R1164_U198;
  assign new_P2_R1164_U202 = ~new_P2_R1164_U5 | ~new_P2_R1164_U41;
  assign new_P2_R1164_U203 = ~new_P2_R1164_U144;
  assign new_P2_R1164_U204 = new_P2_U3453 | new_P2_U3086;
  assign new_P2_R1164_U205 = ~new_P2_R1164_U204 | ~new_P2_R1164_U144;
  assign new_P2_R1164_U206 = ~new_P2_R1164_U40;
  assign new_P2_R1164_U207 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1164_U208 = new_P2_U3447 | new_P2_U3073;
  assign new_P2_R1164_U209 = ~new_P2_R1164_U208 | ~new_P2_R1164_U41;
  assign new_P2_R1164_U210 = ~new_P2_R1164_U119 | ~new_P2_R1164_U209;
  assign new_P2_R1164_U211 = ~new_P2_R1164_U195 | ~new_P2_R1164_U22;
  assign new_P2_R1164_U212 = ~new_P2_U3450 | ~new_P2_U3072;
  assign new_P2_R1164_U213 = ~new_P2_R1164_U120 | ~new_P2_R1164_U211;
  assign new_P2_R1164_U214 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1164_U215 = ~new_P2_R1164_U185 | ~new_P2_R1164_U181;
  assign new_P2_R1164_U216 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1164_U217 = ~new_P2_R1164_U45;
  assign new_P2_R1164_U218 = ~new_P2_R1164_U121 | ~new_P2_R1164_U184;
  assign new_P2_R1164_U219 = ~new_P2_R1164_U45 | ~new_P2_R1164_U180;
  assign new_P2_R1164_U220 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1164_U221 = ~new_P2_R1164_U44;
  assign new_P2_R1164_U222 = new_P2_U3441 | new_P2_U3062;
  assign new_P2_R1164_U223 = ~new_P2_R1164_U222 | ~new_P2_R1164_U44;
  assign new_P2_R1164_U224 = ~new_P2_R1164_U123 | ~new_P2_R1164_U223;
  assign new_P2_R1164_U225 = ~new_P2_R1164_U221 | ~new_P2_R1164_U34;
  assign new_P2_R1164_U226 = ~new_P2_U3444 | ~new_P2_U3069;
  assign new_P2_R1164_U227 = ~new_P2_R1164_U124 | ~new_P2_R1164_U225;
  assign new_P2_R1164_U228 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1164_U229 = ~new_P2_R1164_U184 | ~new_P2_R1164_U181;
  assign new_P2_R1164_U230 = ~new_P2_R1164_U145;
  assign new_P2_R1164_U231 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1164_U232 = ~new_P2_R1164_U42 | ~new_P2_R1164_U43 | ~new_P2_R1164_U401 | ~new_P2_R1164_U400;
  assign new_P2_R1164_U233 = ~new_P2_R1164_U43 | ~new_P2_R1164_U42;
  assign new_P2_R1164_U234 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1164_U235 = ~new_P2_R1164_U125 | ~new_P2_R1164_U233;
  assign new_P2_R1164_U236 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1164_U237 = new_P2_U3064 | new_P2_U3459;
  assign new_P2_R1164_U238 = ~new_P2_R1164_U177 | ~new_P2_R1164_U6;
  assign new_P2_R1164_U239 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1164_U240 = ~new_P2_R1164_U127 | ~new_P2_R1164_U238;
  assign new_P2_R1164_U241 = new_P2_U3459 | new_P2_U3064;
  assign new_P2_R1164_U242 = ~new_P2_R1164_U126 | ~new_P2_R1164_U144;
  assign new_P2_R1164_U243 = ~new_P2_R1164_U241 | ~new_P2_R1164_U240;
  assign new_P2_R1164_U244 = ~new_P2_R1164_U167;
  assign new_P2_R1164_U245 = new_P2_U3082 | new_P2_U3468;
  assign new_P2_R1164_U246 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1164_U247 = ~new_P2_R1164_U174 | ~new_P2_R1164_U7;
  assign new_P2_R1164_U248 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1164_U249 = ~new_P2_R1164_U129 | ~new_P2_R1164_U247;
  assign new_P2_R1164_U250 = new_P2_U3462 | new_P2_U3065;
  assign new_P2_R1164_U251 = new_P2_U3468 | new_P2_U3082;
  assign new_P2_R1164_U252 = ~new_P2_R1164_U128 | ~new_P2_R1164_U167;
  assign new_P2_R1164_U253 = ~new_P2_R1164_U251 | ~new_P2_R1164_U249;
  assign new_P2_R1164_U254 = ~new_P2_R1164_U166;
  assign new_P2_R1164_U255 = new_P2_U3471 | new_P2_U3081;
  assign new_P2_R1164_U256 = ~new_P2_R1164_U255 | ~new_P2_R1164_U166;
  assign new_P2_R1164_U257 = ~new_P2_U3081 | ~new_P2_U3471;
  assign new_P2_R1164_U258 = ~new_P2_R1164_U164;
  assign new_P2_R1164_U259 = new_P2_U3474 | new_P2_U3076;
  assign new_P2_R1164_U260 = ~new_P2_R1164_U259 | ~new_P2_R1164_U164;
  assign new_P2_R1164_U261 = ~new_P2_U3076 | ~new_P2_U3474;
  assign new_P2_R1164_U262 = ~new_P2_R1164_U92;
  assign new_P2_R1164_U263 = new_P2_U3071 | new_P2_U3480;
  assign new_P2_R1164_U264 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1164_U265 = ~new_P2_R1164_U59;
  assign new_P2_R1164_U266 = ~new_P2_R1164_U60 | ~new_P2_R1164_U59;
  assign new_P2_R1164_U267 = ~new_P2_U3071 | ~new_P2_R1164_U266;
  assign new_P2_R1164_U268 = ~new_P2_U3480 | ~new_P2_R1164_U265;
  assign new_P2_R1164_U269 = ~new_P2_R1164_U8 | ~new_P2_R1164_U92;
  assign new_P2_R1164_U270 = ~new_P2_R1164_U162;
  assign new_P2_R1164_U271 = new_P2_U3078 | new_P2_U3957;
  assign new_P2_R1164_U272 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1164_U273 = new_P2_U3077 | new_P2_U3956;
  assign new_P2_R1164_U274 = ~new_P2_R1164_U80;
  assign new_P2_R1164_U275 = ~new_P2_U3957 | ~new_P2_R1164_U274;
  assign new_P2_R1164_U276 = ~new_P2_R1164_U275 | ~new_P2_R1164_U90;
  assign new_P2_R1164_U277 = ~new_P2_R1164_U80 | ~new_P2_R1164_U81;
  assign new_P2_R1164_U278 = ~new_P2_R1164_U277 | ~new_P2_R1164_U276;
  assign new_P2_R1164_U279 = ~new_P2_R1164_U175 | ~new_P2_R1164_U9;
  assign new_P2_R1164_U280 = ~new_P2_U3077 | ~new_P2_U3956;
  assign new_P2_R1164_U281 = ~new_P2_R1164_U278 | ~new_P2_R1164_U279;
  assign new_P2_R1164_U282 = new_P2_U3483 | new_P2_U3084;
  assign new_P2_R1164_U283 = new_P2_U3956 | new_P2_U3077;
  assign new_P2_R1164_U284 = ~new_P2_R1164_U131 | ~new_P2_R1164_U273 | ~new_P2_R1164_U162;
  assign new_P2_R1164_U285 = ~new_P2_R1164_U283 | ~new_P2_R1164_U281;
  assign new_P2_R1164_U286 = ~new_P2_R1164_U159;
  assign new_P2_R1164_U287 = new_P2_U3955 | new_P2_U3063;
  assign new_P2_R1164_U288 = ~new_P2_R1164_U287 | ~new_P2_R1164_U159;
  assign new_P2_R1164_U289 = ~new_P2_U3063 | ~new_P2_U3955;
  assign new_P2_R1164_U290 = ~new_P2_R1164_U157;
  assign new_P2_R1164_U291 = new_P2_U3954 | new_P2_U3068;
  assign new_P2_R1164_U292 = ~new_P2_R1164_U291 | ~new_P2_R1164_U157;
  assign new_P2_R1164_U293 = ~new_P2_U3068 | ~new_P2_U3954;
  assign new_P2_R1164_U294 = ~new_P2_R1164_U155;
  assign new_P2_R1164_U295 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1164_U296 = ~new_P2_R1164_U176 | ~new_P2_R1164_U173;
  assign new_P2_R1164_U297 = ~new_P2_R1164_U86;
  assign new_P2_R1164_U298 = new_P2_U3953 | new_P2_U3067;
  assign new_P2_R1164_U299 = ~new_P2_R1164_U168 | ~new_P2_R1164_U155 | ~new_P2_R1164_U298;
  assign new_P2_R1164_U300 = ~new_P2_R1164_U153;
  assign new_P2_R1164_U301 = new_P2_U3950 | new_P2_U3055;
  assign new_P2_R1164_U302 = ~new_P2_U3055 | ~new_P2_U3950;
  assign new_P2_R1164_U303 = ~new_P2_R1164_U151;
  assign new_P2_R1164_U304 = ~new_P2_U3949 | ~new_P2_R1164_U151;
  assign new_P2_R1164_U305 = ~new_P2_R1164_U149;
  assign new_P2_R1164_U306 = ~new_P2_R1164_U298 | ~new_P2_R1164_U155;
  assign new_P2_R1164_U307 = ~new_P2_R1164_U89;
  assign new_P2_R1164_U308 = new_P2_U3952 | new_P2_U3060;
  assign new_P2_R1164_U309 = ~new_P2_R1164_U308 | ~new_P2_R1164_U89;
  assign new_P2_R1164_U310 = ~new_P2_R1164_U154 | ~new_P2_R1164_U309 | ~new_P2_R1164_U173;
  assign new_P2_R1164_U311 = ~new_P2_R1164_U307 | ~new_P2_R1164_U173;
  assign new_P2_R1164_U312 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1164_U313 = ~new_P2_R1164_U168 | ~new_P2_R1164_U311 | ~new_P2_R1164_U312;
  assign new_P2_R1164_U314 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1164_U315 = ~new_P2_R1164_U282 | ~new_P2_R1164_U162;
  assign new_P2_R1164_U316 = ~new_P2_R1164_U91;
  assign new_P2_R1164_U317 = ~new_P2_R1164_U9 | ~new_P2_R1164_U91;
  assign new_P2_R1164_U318 = ~new_P2_R1164_U135 | ~new_P2_R1164_U317;
  assign new_P2_R1164_U319 = ~new_P2_R1164_U317 | ~new_P2_R1164_U278;
  assign new_P2_R1164_U320 = ~new_P2_R1164_U453 | ~new_P2_R1164_U319;
  assign new_P2_R1164_U321 = new_P2_U3485 | new_P2_U3083;
  assign new_P2_R1164_U322 = ~new_P2_R1164_U321 | ~new_P2_R1164_U91;
  assign new_P2_R1164_U323 = ~new_P2_R1164_U136 | ~new_P2_R1164_U322;
  assign new_P2_R1164_U324 = ~new_P2_R1164_U316 | ~new_P2_R1164_U80;
  assign new_P2_R1164_U325 = ~new_P2_U3078 | ~new_P2_U3957;
  assign new_P2_R1164_U326 = ~new_P2_R1164_U137 | ~new_P2_R1164_U324;
  assign new_P2_R1164_U327 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1164_U328 = ~new_P2_R1164_U161;
  assign new_P2_R1164_U329 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1164_U330 = new_P2_U3477 | new_P2_U3075;
  assign new_P2_R1164_U331 = ~new_P2_R1164_U330 | ~new_P2_R1164_U92;
  assign new_P2_R1164_U332 = ~new_P2_R1164_U138 | ~new_P2_R1164_U331;
  assign new_P2_R1164_U333 = ~new_P2_R1164_U262 | ~new_P2_R1164_U59;
  assign new_P2_R1164_U334 = ~new_P2_U3480 | ~new_P2_U3071;
  assign new_P2_R1164_U335 = ~new_P2_R1164_U139 | ~new_P2_R1164_U333;
  assign new_P2_R1164_U336 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1164_U337 = ~new_P2_R1164_U250 | ~new_P2_R1164_U167;
  assign new_P2_R1164_U338 = ~new_P2_R1164_U93;
  assign new_P2_R1164_U339 = new_P2_U3465 | new_P2_U3074;
  assign new_P2_R1164_U340 = ~new_P2_R1164_U339 | ~new_P2_R1164_U93;
  assign new_P2_R1164_U341 = ~new_P2_R1164_U140 | ~new_P2_R1164_U340;
  assign new_P2_R1164_U342 = ~new_P2_R1164_U338 | ~new_P2_R1164_U172;
  assign new_P2_R1164_U343 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1164_U344 = ~new_P2_R1164_U141 | ~new_P2_R1164_U342;
  assign new_P2_R1164_U345 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1164_U346 = new_P2_U3456 | new_P2_U3085;
  assign new_P2_R1164_U347 = ~new_P2_R1164_U346 | ~new_P2_R1164_U40;
  assign new_P2_R1164_U348 = ~new_P2_R1164_U142 | ~new_P2_R1164_U347;
  assign new_P2_R1164_U349 = ~new_P2_R1164_U206 | ~new_P2_R1164_U171;
  assign new_P2_R1164_U350 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1164_U351 = ~new_P2_R1164_U143 | ~new_P2_R1164_U349;
  assign new_P2_R1164_U352 = ~new_P2_R1164_U207 | ~new_P2_R1164_U171;
  assign new_P2_R1164_U353 = ~new_P2_R1164_U204 | ~new_P2_R1164_U61;
  assign new_P2_R1164_U354 = ~new_P2_R1164_U214 | ~new_P2_R1164_U22;
  assign new_P2_R1164_U355 = ~new_P2_R1164_U228 | ~new_P2_R1164_U34;
  assign new_P2_R1164_U356 = ~new_P2_R1164_U231 | ~new_P2_R1164_U180;
  assign new_P2_R1164_U357 = ~new_P2_R1164_U314 | ~new_P2_R1164_U173;
  assign new_P2_R1164_U358 = ~new_P2_R1164_U298 | ~new_P2_R1164_U176;
  assign new_P2_R1164_U359 = ~new_P2_R1164_U329 | ~new_P2_R1164_U80;
  assign new_P2_R1164_U360 = ~new_P2_R1164_U282 | ~new_P2_R1164_U77;
  assign new_P2_R1164_U361 = ~new_P2_R1164_U336 | ~new_P2_R1164_U59;
  assign new_P2_R1164_U362 = ~new_P2_R1164_U345 | ~new_P2_R1164_U172;
  assign new_P2_R1164_U363 = ~new_P2_R1164_U250 | ~new_P2_R1164_U68;
  assign new_P2_R1164_U364 = ~new_P2_U3949 | ~new_P2_U3056;
  assign new_P2_R1164_U365 = ~new_P2_R1164_U296 | ~new_P2_R1164_U168;
  assign new_P2_R1164_U366 = ~new_P2_U3059 | ~new_P2_R1164_U295;
  assign new_P2_R1164_U367 = ~new_P2_U3951 | ~new_P2_R1164_U295;
  assign new_P2_R1164_U368 = ~new_P2_R1164_U301 | ~new_P2_R1164_U296 | ~new_P2_R1164_U168;
  assign new_P2_R1164_U369 = ~new_P2_R1164_U133 | ~new_P2_R1164_U155 | ~new_P2_R1164_U168;
  assign new_P2_R1164_U370 = ~new_P2_R1164_U297 | ~new_P2_R1164_U301;
  assign new_P2_R1164_U371 = ~new_P2_U3085 | ~new_P2_R1164_U39;
  assign new_P2_R1164_U372 = ~new_P2_U3456 | ~new_P2_R1164_U38;
  assign new_P2_R1164_U373 = ~new_P2_R1164_U372 | ~new_P2_R1164_U371;
  assign new_P2_R1164_U374 = ~new_P2_R1164_U352 | ~new_P2_R1164_U40;
  assign new_P2_R1164_U375 = ~new_P2_R1164_U373 | ~new_P2_R1164_U206;
  assign new_P2_R1164_U376 = ~new_P2_U3086 | ~new_P2_R1164_U36;
  assign new_P2_R1164_U377 = ~new_P2_U3453 | ~new_P2_R1164_U37;
  assign new_P2_R1164_U378 = ~new_P2_R1164_U377 | ~new_P2_R1164_U376;
  assign new_P2_R1164_U379 = ~new_P2_R1164_U353 | ~new_P2_R1164_U144;
  assign new_P2_R1164_U380 = ~new_P2_R1164_U203 | ~new_P2_R1164_U378;
  assign new_P2_R1164_U381 = ~new_P2_U3072 | ~new_P2_R1164_U23;
  assign new_P2_R1164_U382 = ~new_P2_U3450 | ~new_P2_R1164_U21;
  assign new_P2_R1164_U383 = ~new_P2_U3073 | ~new_P2_R1164_U19;
  assign new_P2_R1164_U384 = ~new_P2_U3447 | ~new_P2_R1164_U20;
  assign new_P2_R1164_U385 = ~new_P2_R1164_U384 | ~new_P2_R1164_U383;
  assign new_P2_R1164_U386 = ~new_P2_R1164_U354 | ~new_P2_R1164_U41;
  assign new_P2_R1164_U387 = ~new_P2_R1164_U385 | ~new_P2_R1164_U195;
  assign new_P2_R1164_U388 = ~new_P2_U3069 | ~new_P2_R1164_U35;
  assign new_P2_R1164_U389 = ~new_P2_U3444 | ~new_P2_R1164_U26;
  assign new_P2_R1164_U390 = ~new_P2_U3062 | ~new_P2_R1164_U24;
  assign new_P2_R1164_U391 = ~new_P2_U3441 | ~new_P2_R1164_U25;
  assign new_P2_R1164_U392 = ~new_P2_R1164_U391 | ~new_P2_R1164_U390;
  assign new_P2_R1164_U393 = ~new_P2_R1164_U355 | ~new_P2_R1164_U44;
  assign new_P2_R1164_U394 = ~new_P2_R1164_U392 | ~new_P2_R1164_U221;
  assign new_P2_R1164_U395 = ~new_P2_U3066 | ~new_P2_R1164_U32;
  assign new_P2_R1164_U396 = ~new_P2_U3438 | ~new_P2_R1164_U33;
  assign new_P2_R1164_U397 = ~new_P2_R1164_U396 | ~new_P2_R1164_U395;
  assign new_P2_R1164_U398 = ~new_P2_R1164_U356 | ~new_P2_R1164_U145;
  assign new_P2_R1164_U399 = ~new_P2_R1164_U230 | ~new_P2_R1164_U397;
  assign new_P2_R1164_U400 = ~new_P2_U3070 | ~new_P2_R1164_U27;
  assign new_P2_R1164_U401 = ~new_P2_U3435 | ~new_P2_R1164_U28;
  assign new_P2_R1164_U402 = ~new_P2_U3057 | ~new_P2_R1164_U147;
  assign new_P2_R1164_U403 = ~new_P2_U3960 | ~new_P2_R1164_U146;
  assign new_P2_R1164_U404 = ~new_P2_U3057 | ~new_P2_R1164_U147;
  assign new_P2_R1164_U405 = ~new_P2_U3960 | ~new_P2_R1164_U146;
  assign new_P2_R1164_U406 = ~new_P2_R1164_U405 | ~new_P2_R1164_U404;
  assign new_P2_R1164_U407 = ~new_P2_R1164_U148 | ~new_P2_R1164_U149;
  assign new_P2_R1164_U408 = ~new_P2_R1164_U305 | ~new_P2_R1164_U406;
  assign new_P2_R1164_U409 = ~new_P2_U3056 | ~new_P2_R1164_U88;
  assign new_P2_R1164_U410 = ~new_P2_U3949 | ~new_P2_R1164_U87;
  assign new_P2_R1164_U411 = ~new_P2_U3056 | ~new_P2_R1164_U88;
  assign new_P2_R1164_U412 = ~new_P2_U3949 | ~new_P2_R1164_U87;
  assign new_P2_R1164_U413 = ~new_P2_R1164_U412 | ~new_P2_R1164_U411;
  assign new_P2_R1164_U414 = ~new_P2_R1164_U150 | ~new_P2_R1164_U151;
  assign new_P2_R1164_U415 = ~new_P2_R1164_U303 | ~new_P2_R1164_U413;
  assign new_P2_R1164_U416 = ~new_P2_U3055 | ~new_P2_R1164_U46;
  assign new_P2_R1164_U417 = ~new_P2_U3950 | ~new_P2_R1164_U47;
  assign new_P2_R1164_U418 = ~new_P2_U3055 | ~new_P2_R1164_U46;
  assign new_P2_R1164_U419 = ~new_P2_U3950 | ~new_P2_R1164_U47;
  assign new_P2_R1164_U420 = ~new_P2_R1164_U419 | ~new_P2_R1164_U418;
  assign new_P2_R1164_U421 = ~new_P2_R1164_U152 | ~new_P2_R1164_U153;
  assign new_P2_R1164_U422 = ~new_P2_R1164_U300 | ~new_P2_R1164_U420;
  assign new_P2_R1164_U423 = ~new_P2_U3059 | ~new_P2_R1164_U49;
  assign new_P2_R1164_U424 = ~new_P2_U3951 | ~new_P2_R1164_U48;
  assign new_P2_R1164_U425 = ~new_P2_U3060 | ~new_P2_R1164_U50;
  assign new_P2_R1164_U426 = ~new_P2_U3952 | ~new_P2_R1164_U51;
  assign new_P2_R1164_U427 = ~new_P2_R1164_U426 | ~new_P2_R1164_U425;
  assign new_P2_R1164_U428 = ~new_P2_R1164_U357 | ~new_P2_R1164_U89;
  assign new_P2_R1164_U429 = ~new_P2_R1164_U427 | ~new_P2_R1164_U307;
  assign new_P2_R1164_U430 = ~new_P2_U3067 | ~new_P2_R1164_U52;
  assign new_P2_R1164_U431 = ~new_P2_U3953 | ~new_P2_R1164_U53;
  assign new_P2_R1164_U432 = ~new_P2_R1164_U431 | ~new_P2_R1164_U430;
  assign new_P2_R1164_U433 = ~new_P2_R1164_U358 | ~new_P2_R1164_U155;
  assign new_P2_R1164_U434 = ~new_P2_R1164_U294 | ~new_P2_R1164_U432;
  assign new_P2_R1164_U435 = ~new_P2_U3068 | ~new_P2_R1164_U84;
  assign new_P2_R1164_U436 = ~new_P2_U3954 | ~new_P2_R1164_U85;
  assign new_P2_R1164_U437 = ~new_P2_U3068 | ~new_P2_R1164_U84;
  assign new_P2_R1164_U438 = ~new_P2_U3954 | ~new_P2_R1164_U85;
  assign new_P2_R1164_U439 = ~new_P2_R1164_U438 | ~new_P2_R1164_U437;
  assign new_P2_R1164_U440 = ~new_P2_R1164_U156 | ~new_P2_R1164_U157;
  assign new_P2_R1164_U441 = ~new_P2_R1164_U290 | ~new_P2_R1164_U439;
  assign new_P2_R1164_U442 = ~new_P2_U3063 | ~new_P2_R1164_U82;
  assign new_P2_R1164_U443 = ~new_P2_U3955 | ~new_P2_R1164_U83;
  assign new_P2_R1164_U444 = ~new_P2_U3063 | ~new_P2_R1164_U82;
  assign new_P2_R1164_U445 = ~new_P2_U3955 | ~new_P2_R1164_U83;
  assign new_P2_R1164_U446 = ~new_P2_R1164_U445 | ~new_P2_R1164_U444;
  assign new_P2_R1164_U447 = ~new_P2_R1164_U158 | ~new_P2_R1164_U159;
  assign new_P2_R1164_U448 = ~new_P2_R1164_U286 | ~new_P2_R1164_U446;
  assign new_P2_R1164_U449 = ~new_P2_U3077 | ~new_P2_R1164_U54;
  assign new_P2_R1164_U450 = ~new_P2_U3956 | ~new_P2_R1164_U55;
  assign new_P2_R1164_U451 = ~new_P2_U3077 | ~new_P2_R1164_U54;
  assign new_P2_R1164_U452 = ~new_P2_U3956 | ~new_P2_R1164_U55;
  assign new_P2_R1164_U453 = ~new_P2_R1164_U452 | ~new_P2_R1164_U451;
  assign new_P2_R1164_U454 = ~new_P2_U3078 | ~new_P2_R1164_U81;
  assign new_P2_R1164_U455 = ~new_P2_U3957 | ~new_P2_R1164_U90;
  assign new_P2_R1164_U456 = ~new_P2_R1164_U182 | ~new_P2_R1164_U161;
  assign new_P2_R1164_U457 = ~new_P2_R1164_U328 | ~new_P2_R1164_U31;
  assign new_P2_R1164_U458 = ~new_P2_U3083 | ~new_P2_R1164_U78;
  assign new_P2_R1164_U459 = ~new_P2_U3485 | ~new_P2_R1164_U79;
  assign new_P2_R1164_U460 = ~new_P2_R1164_U459 | ~new_P2_R1164_U458;
  assign new_P2_R1164_U461 = ~new_P2_R1164_U359 | ~new_P2_R1164_U91;
  assign new_P2_R1164_U462 = ~new_P2_R1164_U460 | ~new_P2_R1164_U316;
  assign new_P2_R1164_U463 = ~new_P2_U3084 | ~new_P2_R1164_U75;
  assign new_P2_R1164_U464 = ~new_P2_U3483 | ~new_P2_R1164_U76;
  assign new_P2_R1164_U465 = ~new_P2_R1164_U464 | ~new_P2_R1164_U463;
  assign new_P2_R1164_U466 = ~new_P2_R1164_U360 | ~new_P2_R1164_U162;
  assign new_P2_R1164_U467 = ~new_P2_R1164_U270 | ~new_P2_R1164_U465;
  assign new_P2_R1164_U468 = ~new_P2_U3071 | ~new_P2_R1164_U60;
  assign new_P2_R1164_U469 = ~new_P2_U3480 | ~new_P2_R1164_U58;
  assign new_P2_R1164_U470 = ~new_P2_U3075 | ~new_P2_R1164_U56;
  assign new_P2_R1164_U471 = ~new_P2_U3477 | ~new_P2_R1164_U57;
  assign new_P2_R1164_U472 = ~new_P2_R1164_U471 | ~new_P2_R1164_U470;
  assign new_P2_R1164_U473 = ~new_P2_R1164_U361 | ~new_P2_R1164_U92;
  assign new_P2_R1164_U474 = ~new_P2_R1164_U472 | ~new_P2_R1164_U262;
  assign new_P2_R1164_U475 = ~new_P2_U3076 | ~new_P2_R1164_U73;
  assign new_P2_R1164_U476 = ~new_P2_U3474 | ~new_P2_R1164_U74;
  assign new_P2_R1164_U477 = ~new_P2_U3076 | ~new_P2_R1164_U73;
  assign new_P2_R1164_U478 = ~new_P2_U3474 | ~new_P2_R1164_U74;
  assign new_P2_R1164_U479 = ~new_P2_R1164_U478 | ~new_P2_R1164_U477;
  assign new_P2_R1164_U480 = ~new_P2_R1164_U163 | ~new_P2_R1164_U164;
  assign new_P2_R1164_U481 = ~new_P2_R1164_U258 | ~new_P2_R1164_U479;
  assign new_P2_R1164_U482 = ~new_P2_U3081 | ~new_P2_R1164_U71;
  assign new_P2_R1164_U483 = ~new_P2_U3471 | ~new_P2_R1164_U72;
  assign new_P2_R1164_U484 = ~new_P2_U3081 | ~new_P2_R1164_U71;
  assign new_P2_R1164_U485 = ~new_P2_U3471 | ~new_P2_R1164_U72;
  assign new_P2_R1164_U486 = ~new_P2_R1164_U485 | ~new_P2_R1164_U484;
  assign new_P2_R1164_U487 = ~new_P2_R1164_U165 | ~new_P2_R1164_U166;
  assign new_P2_R1164_U488 = ~new_P2_R1164_U254 | ~new_P2_R1164_U486;
  assign new_P2_R1164_U489 = ~new_P2_U3082 | ~new_P2_R1164_U69;
  assign new_P2_R1164_U490 = ~new_P2_U3468 | ~new_P2_R1164_U70;
  assign new_P2_R1164_U491 = ~new_P2_U3074 | ~new_P2_R1164_U64;
  assign new_P2_R1164_U492 = ~new_P2_U3465 | ~new_P2_R1164_U65;
  assign new_P2_R1164_U493 = ~new_P2_R1164_U492 | ~new_P2_R1164_U491;
  assign new_P2_R1164_U494 = ~new_P2_R1164_U362 | ~new_P2_R1164_U93;
  assign new_P2_R1164_U495 = ~new_P2_R1164_U493 | ~new_P2_R1164_U338;
  assign new_P2_R1164_U496 = ~new_P2_U3065 | ~new_P2_R1164_U66;
  assign new_P2_R1164_U497 = ~new_P2_U3462 | ~new_P2_R1164_U67;
  assign new_P2_R1164_U498 = ~new_P2_R1164_U497 | ~new_P2_R1164_U496;
  assign new_P2_R1164_U499 = ~new_P2_R1164_U363 | ~new_P2_R1164_U167;
  assign new_P2_R1164_U500 = ~new_P2_R1164_U244 | ~new_P2_R1164_U498;
  assign new_P2_R1164_U501 = ~new_P2_U3064 | ~new_P2_R1164_U62;
  assign new_P2_R1164_U502 = ~new_P2_U3459 | ~new_P2_R1164_U63;
  assign new_P2_R1164_U503 = ~new_P2_U3079 | ~new_P2_R1164_U29;
  assign new_P2_R1164_U504 = ~new_P2_U3427 | ~new_P2_R1164_U30;
  assign new_P2_R1233_U4 = new_P2_R1233_U179 & new_P2_R1233_U178;
  assign new_P2_R1233_U5 = new_P2_R1233_U197 & new_P2_R1233_U196;
  assign new_P2_R1233_U6 = new_P2_R1233_U237 & new_P2_R1233_U236;
  assign new_P2_R1233_U7 = new_P2_R1233_U246 & new_P2_R1233_U245;
  assign new_P2_R1233_U8 = new_P2_R1233_U264 & new_P2_R1233_U263;
  assign new_P2_R1233_U9 = new_P2_R1233_U272 & new_P2_R1233_U271;
  assign new_P2_R1233_U10 = new_P2_R1233_U351 & new_P2_R1233_U348;
  assign new_P2_R1233_U11 = new_P2_R1233_U344 & new_P2_R1233_U341;
  assign new_P2_R1233_U12 = new_P2_R1233_U335 & new_P2_R1233_U332;
  assign new_P2_R1233_U13 = new_P2_R1233_U326 & new_P2_R1233_U323;
  assign new_P2_R1233_U14 = new_P2_R1233_U320 & new_P2_R1233_U318;
  assign new_P2_R1233_U15 = new_P2_R1233_U313 & new_P2_R1233_U310;
  assign new_P2_R1233_U16 = new_P2_R1233_U235 & new_P2_R1233_U232;
  assign new_P2_R1233_U17 = new_P2_R1233_U227 & new_P2_R1233_U224;
  assign new_P2_R1233_U18 = new_P2_R1233_U213 & new_P2_R1233_U210;
  assign new_P2_R1233_U19 = ~new_P2_U3447;
  assign new_P2_R1233_U20 = ~new_P2_U3073;
  assign new_P2_R1233_U21 = ~new_P2_U3072;
  assign new_P2_R1233_U22 = ~new_P2_U3073 | ~new_P2_U3447;
  assign new_P2_R1233_U23 = ~new_P2_U3450;
  assign new_P2_R1233_U24 = ~new_P2_U3441;
  assign new_P2_R1233_U25 = ~new_P2_U3062;
  assign new_P2_R1233_U26 = ~new_P2_U3069;
  assign new_P2_R1233_U27 = ~new_P2_U3435;
  assign new_P2_R1233_U28 = ~new_P2_U3070;
  assign new_P2_R1233_U29 = ~new_P2_U3427;
  assign new_P2_R1233_U30 = ~new_P2_U3079;
  assign new_P2_R1233_U31 = ~new_P2_U3079 | ~new_P2_U3427;
  assign new_P2_R1233_U32 = ~new_P2_U3438;
  assign new_P2_R1233_U33 = ~new_P2_U3066;
  assign new_P2_R1233_U34 = ~new_P2_U3062 | ~new_P2_U3441;
  assign new_P2_R1233_U35 = ~new_P2_U3444;
  assign new_P2_R1233_U36 = ~new_P2_U3453;
  assign new_P2_R1233_U37 = ~new_P2_U3086;
  assign new_P2_R1233_U38 = ~new_P2_U3085;
  assign new_P2_R1233_U39 = ~new_P2_U3456;
  assign new_P2_R1233_U40 = ~new_P2_R1233_U61 | ~new_P2_R1233_U205;
  assign new_P2_R1233_U41 = ~new_P2_R1233_U117 | ~new_P2_R1233_U193;
  assign new_P2_R1233_U42 = ~new_P2_R1233_U182 | ~new_P2_R1233_U183;
  assign new_P2_R1233_U43 = ~new_P2_U3432 | ~new_P2_U3080;
  assign new_P2_R1233_U44 = ~new_P2_R1233_U122 | ~new_P2_R1233_U219;
  assign new_P2_R1233_U45 = ~new_P2_R1233_U216 | ~new_P2_R1233_U215;
  assign new_P2_R1233_U46 = ~new_P2_U3950;
  assign new_P2_R1233_U47 = ~new_P2_U3055;
  assign new_P2_R1233_U48 = ~new_P2_U3059;
  assign new_P2_R1233_U49 = ~new_P2_U3951;
  assign new_P2_R1233_U50 = ~new_P2_U3952;
  assign new_P2_R1233_U51 = ~new_P2_U3060;
  assign new_P2_R1233_U52 = ~new_P2_U3953;
  assign new_P2_R1233_U53 = ~new_P2_U3067;
  assign new_P2_R1233_U54 = ~new_P2_U3956;
  assign new_P2_R1233_U55 = ~new_P2_U3077;
  assign new_P2_R1233_U56 = ~new_P2_U3477;
  assign new_P2_R1233_U57 = ~new_P2_U3075;
  assign new_P2_R1233_U58 = ~new_P2_U3071;
  assign new_P2_R1233_U59 = ~new_P2_U3075 | ~new_P2_U3477;
  assign new_P2_R1233_U60 = ~new_P2_U3480;
  assign new_P2_R1233_U61 = ~new_P2_U3086 | ~new_P2_U3453;
  assign new_P2_R1233_U62 = ~new_P2_U3459;
  assign new_P2_R1233_U63 = ~new_P2_U3064;
  assign new_P2_R1233_U64 = ~new_P2_U3465;
  assign new_P2_R1233_U65 = ~new_P2_U3074;
  assign new_P2_R1233_U66 = ~new_P2_U3462;
  assign new_P2_R1233_U67 = ~new_P2_U3065;
  assign new_P2_R1233_U68 = ~new_P2_U3065 | ~new_P2_U3462;
  assign new_P2_R1233_U69 = ~new_P2_U3468;
  assign new_P2_R1233_U70 = ~new_P2_U3082;
  assign new_P2_R1233_U71 = ~new_P2_U3471;
  assign new_P2_R1233_U72 = ~new_P2_U3081;
  assign new_P2_R1233_U73 = ~new_P2_U3474;
  assign new_P2_R1233_U74 = ~new_P2_U3076;
  assign new_P2_R1233_U75 = ~new_P2_U3483;
  assign new_P2_R1233_U76 = ~new_P2_U3084;
  assign new_P2_R1233_U77 = ~new_P2_U3084 | ~new_P2_U3483;
  assign new_P2_R1233_U78 = ~new_P2_U3485;
  assign new_P2_R1233_U79 = ~new_P2_U3083;
  assign new_P2_R1233_U80 = ~new_P2_U3083 | ~new_P2_U3485;
  assign new_P2_R1233_U81 = ~new_P2_U3957;
  assign new_P2_R1233_U82 = ~new_P2_U3955;
  assign new_P2_R1233_U83 = ~new_P2_U3063;
  assign new_P2_R1233_U84 = ~new_P2_U3954;
  assign new_P2_R1233_U85 = ~new_P2_U3068;
  assign new_P2_R1233_U86 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1233_U87 = ~new_P2_U3056;
  assign new_P2_R1233_U88 = ~new_P2_U3949;
  assign new_P2_R1233_U89 = ~new_P2_R1233_U306 | ~new_P2_R1233_U176;
  assign new_P2_R1233_U90 = ~new_P2_U3078;
  assign new_P2_R1233_U91 = ~new_P2_R1233_U77 | ~new_P2_R1233_U315;
  assign new_P2_R1233_U92 = ~new_P2_R1233_U261 | ~new_P2_R1233_U260;
  assign new_P2_R1233_U93 = ~new_P2_R1233_U68 | ~new_P2_R1233_U337;
  assign new_P2_R1233_U94 = ~new_P2_R1233_U457 | ~new_P2_R1233_U456;
  assign new_P2_R1233_U95 = ~new_P2_R1233_U504 | ~new_P2_R1233_U503;
  assign new_P2_R1233_U96 = ~new_P2_R1233_U375 | ~new_P2_R1233_U374;
  assign new_P2_R1233_U97 = ~new_P2_R1233_U380 | ~new_P2_R1233_U379;
  assign new_P2_R1233_U98 = ~new_P2_R1233_U387 | ~new_P2_R1233_U386;
  assign new_P2_R1233_U99 = ~new_P2_R1233_U394 | ~new_P2_R1233_U393;
  assign new_P2_R1233_U100 = ~new_P2_R1233_U399 | ~new_P2_R1233_U398;
  assign new_P2_R1233_U101 = ~new_P2_R1233_U408 | ~new_P2_R1233_U407;
  assign new_P2_R1233_U102 = ~new_P2_R1233_U415 | ~new_P2_R1233_U414;
  assign new_P2_R1233_U103 = ~new_P2_R1233_U422 | ~new_P2_R1233_U421;
  assign new_P2_R1233_U104 = ~new_P2_R1233_U429 | ~new_P2_R1233_U428;
  assign new_P2_R1233_U105 = ~new_P2_R1233_U434 | ~new_P2_R1233_U433;
  assign new_P2_R1233_U106 = ~new_P2_R1233_U441 | ~new_P2_R1233_U440;
  assign new_P2_R1233_U107 = ~new_P2_R1233_U448 | ~new_P2_R1233_U447;
  assign new_P2_R1233_U108 = ~new_P2_R1233_U462 | ~new_P2_R1233_U461;
  assign new_P2_R1233_U109 = ~new_P2_R1233_U467 | ~new_P2_R1233_U466;
  assign new_P2_R1233_U110 = ~new_P2_R1233_U474 | ~new_P2_R1233_U473;
  assign new_P2_R1233_U111 = ~new_P2_R1233_U481 | ~new_P2_R1233_U480;
  assign new_P2_R1233_U112 = ~new_P2_R1233_U488 | ~new_P2_R1233_U487;
  assign new_P2_R1233_U113 = ~new_P2_R1233_U495 | ~new_P2_R1233_U494;
  assign new_P2_R1233_U114 = ~new_P2_R1233_U500 | ~new_P2_R1233_U499;
  assign new_P2_R1233_U115 = new_P2_R1233_U189 & new_P2_R1233_U187;
  assign new_P2_R1233_U116 = new_P2_R1233_U4 & new_P2_R1233_U180;
  assign new_P2_R1233_U117 = new_P2_R1233_U194 & new_P2_R1233_U192;
  assign new_P2_R1233_U118 = new_P2_R1233_U201 & new_P2_R1233_U200;
  assign new_P2_R1233_U119 = new_P2_R1233_U22 & new_P2_R1233_U382 & new_P2_R1233_U381;
  assign new_P2_R1233_U120 = new_P2_R1233_U212 & new_P2_R1233_U5;
  assign new_P2_R1233_U121 = new_P2_R1233_U181 & new_P2_R1233_U180;
  assign new_P2_R1233_U122 = new_P2_R1233_U220 & new_P2_R1233_U218;
  assign new_P2_R1233_U123 = new_P2_R1233_U34 & new_P2_R1233_U389 & new_P2_R1233_U388;
  assign new_P2_R1233_U124 = new_P2_R1233_U226 & new_P2_R1233_U4;
  assign new_P2_R1233_U125 = new_P2_R1233_U234 & new_P2_R1233_U181;
  assign new_P2_R1233_U126 = new_P2_R1233_U204 & new_P2_R1233_U6;
  assign new_P2_R1233_U127 = new_P2_R1233_U239 & new_P2_R1233_U171;
  assign new_P2_R1233_U128 = new_P2_R1233_U250 & new_P2_R1233_U7;
  assign new_P2_R1233_U129 = new_P2_R1233_U248 & new_P2_R1233_U172;
  assign new_P2_R1233_U130 = new_P2_R1233_U268 & new_P2_R1233_U267;
  assign new_P2_R1233_U131 = new_P2_R1233_U9 & new_P2_R1233_U282;
  assign new_P2_R1233_U132 = new_P2_R1233_U285 & new_P2_R1233_U280;
  assign new_P2_R1233_U133 = new_P2_R1233_U301 & new_P2_R1233_U298;
  assign new_P2_R1233_U134 = new_P2_R1233_U368 & new_P2_R1233_U302;
  assign new_P2_R1233_U135 = new_P2_R1233_U160 & new_P2_R1233_U278;
  assign new_P2_R1233_U136 = new_P2_R1233_U80 & new_P2_R1233_U455 & new_P2_R1233_U454;
  assign new_P2_R1233_U137 = new_P2_R1233_U325 & new_P2_R1233_U9;
  assign new_P2_R1233_U138 = new_P2_R1233_U59 & new_P2_R1233_U469 & new_P2_R1233_U468;
  assign new_P2_R1233_U139 = new_P2_R1233_U334 & new_P2_R1233_U8;
  assign new_P2_R1233_U140 = new_P2_R1233_U172 & new_P2_R1233_U490 & new_P2_R1233_U489;
  assign new_P2_R1233_U141 = new_P2_R1233_U343 & new_P2_R1233_U7;
  assign new_P2_R1233_U142 = new_P2_R1233_U171 & new_P2_R1233_U502 & new_P2_R1233_U501;
  assign new_P2_R1233_U143 = new_P2_R1233_U350 & new_P2_R1233_U6;
  assign new_P2_R1233_U144 = ~new_P2_R1233_U118 | ~new_P2_R1233_U202;
  assign new_P2_R1233_U145 = ~new_P2_R1233_U217 | ~new_P2_R1233_U229;
  assign new_P2_R1233_U146 = ~new_P2_U3057;
  assign new_P2_R1233_U147 = ~new_P2_U3960;
  assign new_P2_R1233_U148 = new_P2_R1233_U403 & new_P2_R1233_U402;
  assign new_P2_R1233_U149 = ~new_P2_R1233_U364 | ~new_P2_R1233_U304 | ~new_P2_R1233_U169;
  assign new_P2_R1233_U150 = new_P2_R1233_U410 & new_P2_R1233_U409;
  assign new_P2_R1233_U151 = ~new_P2_R1233_U134 | ~new_P2_R1233_U370 | ~new_P2_R1233_U369;
  assign new_P2_R1233_U152 = new_P2_R1233_U417 & new_P2_R1233_U416;
  assign new_P2_R1233_U153 = ~new_P2_R1233_U86 | ~new_P2_R1233_U365 | ~new_P2_R1233_U299;
  assign new_P2_R1233_U154 = new_P2_R1233_U424 & new_P2_R1233_U423;
  assign new_P2_R1233_U155 = ~new_P2_R1233_U293 | ~new_P2_R1233_U292;
  assign new_P2_R1233_U156 = new_P2_R1233_U436 & new_P2_R1233_U435;
  assign new_P2_R1233_U157 = ~new_P2_R1233_U289 | ~new_P2_R1233_U288;
  assign new_P2_R1233_U158 = new_P2_R1233_U443 & new_P2_R1233_U442;
  assign new_P2_R1233_U159 = ~new_P2_R1233_U132 | ~new_P2_R1233_U284;
  assign new_P2_R1233_U160 = new_P2_R1233_U450 & new_P2_R1233_U449;
  assign new_P2_R1233_U161 = ~new_P2_R1233_U43 | ~new_P2_R1233_U327;
  assign new_P2_R1233_U162 = ~new_P2_R1233_U130 | ~new_P2_R1233_U269;
  assign new_P2_R1233_U163 = new_P2_R1233_U476 & new_P2_R1233_U475;
  assign new_P2_R1233_U164 = ~new_P2_R1233_U257 | ~new_P2_R1233_U256;
  assign new_P2_R1233_U165 = new_P2_R1233_U483 & new_P2_R1233_U482;
  assign new_P2_R1233_U166 = ~new_P2_R1233_U253 | ~new_P2_R1233_U252;
  assign new_P2_R1233_U167 = ~new_P2_R1233_U243 | ~new_P2_R1233_U242;
  assign new_P2_R1233_U168 = ~new_P2_R1233_U367 | ~new_P2_R1233_U366;
  assign new_P2_R1233_U169 = ~new_P2_U3056 | ~new_P2_R1233_U151;
  assign new_P2_R1233_U170 = ~new_P2_R1233_U34;
  assign new_P2_R1233_U171 = ~new_P2_U3456 | ~new_P2_U3085;
  assign new_P2_R1233_U172 = ~new_P2_U3074 | ~new_P2_U3465;
  assign new_P2_R1233_U173 = ~new_P2_U3060 | ~new_P2_U3952;
  assign new_P2_R1233_U174 = ~new_P2_R1233_U68;
  assign new_P2_R1233_U175 = ~new_P2_R1233_U77;
  assign new_P2_R1233_U176 = ~new_P2_U3067 | ~new_P2_U3953;
  assign new_P2_R1233_U177 = ~new_P2_R1233_U61;
  assign new_P2_R1233_U178 = new_P2_U3069 | new_P2_U3444;
  assign new_P2_R1233_U179 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1233_U180 = new_P2_U3438 | new_P2_U3066;
  assign new_P2_R1233_U181 = new_P2_U3435 | new_P2_U3070;
  assign new_P2_R1233_U182 = ~new_P2_R1233_U31;
  assign new_P2_R1233_U183 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1233_U184 = ~new_P2_R1233_U42;
  assign new_P2_R1233_U185 = ~new_P2_R1233_U43;
  assign new_P2_R1233_U186 = ~new_P2_R1233_U42 | ~new_P2_R1233_U43;
  assign new_P2_R1233_U187 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1233_U188 = ~new_P2_R1233_U186 | ~new_P2_R1233_U181;
  assign new_P2_R1233_U189 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1233_U190 = ~new_P2_R1233_U115 | ~new_P2_R1233_U188;
  assign new_P2_R1233_U191 = ~new_P2_R1233_U35 | ~new_P2_R1233_U34;
  assign new_P2_R1233_U192 = ~new_P2_U3069 | ~new_P2_R1233_U191;
  assign new_P2_R1233_U193 = ~new_P2_R1233_U116 | ~new_P2_R1233_U190;
  assign new_P2_R1233_U194 = ~new_P2_U3444 | ~new_P2_R1233_U170;
  assign new_P2_R1233_U195 = ~new_P2_R1233_U41;
  assign new_P2_R1233_U196 = new_P2_U3072 | new_P2_U3450;
  assign new_P2_R1233_U197 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1233_U198 = ~new_P2_R1233_U22;
  assign new_P2_R1233_U199 = ~new_P2_R1233_U23 | ~new_P2_R1233_U22;
  assign new_P2_R1233_U200 = ~new_P2_U3072 | ~new_P2_R1233_U199;
  assign new_P2_R1233_U201 = ~new_P2_U3450 | ~new_P2_R1233_U198;
  assign new_P2_R1233_U202 = ~new_P2_R1233_U5 | ~new_P2_R1233_U41;
  assign new_P2_R1233_U203 = ~new_P2_R1233_U144;
  assign new_P2_R1233_U204 = new_P2_U3453 | new_P2_U3086;
  assign new_P2_R1233_U205 = ~new_P2_R1233_U204 | ~new_P2_R1233_U144;
  assign new_P2_R1233_U206 = ~new_P2_R1233_U40;
  assign new_P2_R1233_U207 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1233_U208 = new_P2_U3447 | new_P2_U3073;
  assign new_P2_R1233_U209 = ~new_P2_R1233_U208 | ~new_P2_R1233_U41;
  assign new_P2_R1233_U210 = ~new_P2_R1233_U119 | ~new_P2_R1233_U209;
  assign new_P2_R1233_U211 = ~new_P2_R1233_U195 | ~new_P2_R1233_U22;
  assign new_P2_R1233_U212 = ~new_P2_U3450 | ~new_P2_U3072;
  assign new_P2_R1233_U213 = ~new_P2_R1233_U120 | ~new_P2_R1233_U211;
  assign new_P2_R1233_U214 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1233_U215 = ~new_P2_R1233_U185 | ~new_P2_R1233_U181;
  assign new_P2_R1233_U216 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1233_U217 = ~new_P2_R1233_U45;
  assign new_P2_R1233_U218 = ~new_P2_R1233_U121 | ~new_P2_R1233_U184;
  assign new_P2_R1233_U219 = ~new_P2_R1233_U45 | ~new_P2_R1233_U180;
  assign new_P2_R1233_U220 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1233_U221 = ~new_P2_R1233_U44;
  assign new_P2_R1233_U222 = new_P2_U3441 | new_P2_U3062;
  assign new_P2_R1233_U223 = ~new_P2_R1233_U222 | ~new_P2_R1233_U44;
  assign new_P2_R1233_U224 = ~new_P2_R1233_U123 | ~new_P2_R1233_U223;
  assign new_P2_R1233_U225 = ~new_P2_R1233_U221 | ~new_P2_R1233_U34;
  assign new_P2_R1233_U226 = ~new_P2_U3444 | ~new_P2_U3069;
  assign new_P2_R1233_U227 = ~new_P2_R1233_U124 | ~new_P2_R1233_U225;
  assign new_P2_R1233_U228 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1233_U229 = ~new_P2_R1233_U184 | ~new_P2_R1233_U181;
  assign new_P2_R1233_U230 = ~new_P2_R1233_U145;
  assign new_P2_R1233_U231 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1233_U232 = ~new_P2_R1233_U42 | ~new_P2_R1233_U43 | ~new_P2_R1233_U401 | ~new_P2_R1233_U400;
  assign new_P2_R1233_U233 = ~new_P2_R1233_U43 | ~new_P2_R1233_U42;
  assign new_P2_R1233_U234 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1233_U235 = ~new_P2_R1233_U125 | ~new_P2_R1233_U233;
  assign new_P2_R1233_U236 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1233_U237 = new_P2_U3064 | new_P2_U3459;
  assign new_P2_R1233_U238 = ~new_P2_R1233_U177 | ~new_P2_R1233_U6;
  assign new_P2_R1233_U239 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1233_U240 = ~new_P2_R1233_U127 | ~new_P2_R1233_U238;
  assign new_P2_R1233_U241 = new_P2_U3459 | new_P2_U3064;
  assign new_P2_R1233_U242 = ~new_P2_R1233_U126 | ~new_P2_R1233_U144;
  assign new_P2_R1233_U243 = ~new_P2_R1233_U241 | ~new_P2_R1233_U240;
  assign new_P2_R1233_U244 = ~new_P2_R1233_U167;
  assign new_P2_R1233_U245 = new_P2_U3082 | new_P2_U3468;
  assign new_P2_R1233_U246 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1233_U247 = ~new_P2_R1233_U174 | ~new_P2_R1233_U7;
  assign new_P2_R1233_U248 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1233_U249 = ~new_P2_R1233_U129 | ~new_P2_R1233_U247;
  assign new_P2_R1233_U250 = new_P2_U3462 | new_P2_U3065;
  assign new_P2_R1233_U251 = new_P2_U3468 | new_P2_U3082;
  assign new_P2_R1233_U252 = ~new_P2_R1233_U128 | ~new_P2_R1233_U167;
  assign new_P2_R1233_U253 = ~new_P2_R1233_U251 | ~new_P2_R1233_U249;
  assign new_P2_R1233_U254 = ~new_P2_R1233_U166;
  assign new_P2_R1233_U255 = new_P2_U3471 | new_P2_U3081;
  assign new_P2_R1233_U256 = ~new_P2_R1233_U255 | ~new_P2_R1233_U166;
  assign new_P2_R1233_U257 = ~new_P2_U3081 | ~new_P2_U3471;
  assign new_P2_R1233_U258 = ~new_P2_R1233_U164;
  assign new_P2_R1233_U259 = new_P2_U3474 | new_P2_U3076;
  assign new_P2_R1233_U260 = ~new_P2_R1233_U259 | ~new_P2_R1233_U164;
  assign new_P2_R1233_U261 = ~new_P2_U3076 | ~new_P2_U3474;
  assign new_P2_R1233_U262 = ~new_P2_R1233_U92;
  assign new_P2_R1233_U263 = new_P2_U3071 | new_P2_U3480;
  assign new_P2_R1233_U264 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1233_U265 = ~new_P2_R1233_U59;
  assign new_P2_R1233_U266 = ~new_P2_R1233_U60 | ~new_P2_R1233_U59;
  assign new_P2_R1233_U267 = ~new_P2_U3071 | ~new_P2_R1233_U266;
  assign new_P2_R1233_U268 = ~new_P2_U3480 | ~new_P2_R1233_U265;
  assign new_P2_R1233_U269 = ~new_P2_R1233_U8 | ~new_P2_R1233_U92;
  assign new_P2_R1233_U270 = ~new_P2_R1233_U162;
  assign new_P2_R1233_U271 = new_P2_U3078 | new_P2_U3957;
  assign new_P2_R1233_U272 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1233_U273 = new_P2_U3077 | new_P2_U3956;
  assign new_P2_R1233_U274 = ~new_P2_R1233_U80;
  assign new_P2_R1233_U275 = ~new_P2_U3957 | ~new_P2_R1233_U274;
  assign new_P2_R1233_U276 = ~new_P2_R1233_U275 | ~new_P2_R1233_U90;
  assign new_P2_R1233_U277 = ~new_P2_R1233_U80 | ~new_P2_R1233_U81;
  assign new_P2_R1233_U278 = ~new_P2_R1233_U277 | ~new_P2_R1233_U276;
  assign new_P2_R1233_U279 = ~new_P2_R1233_U175 | ~new_P2_R1233_U9;
  assign new_P2_R1233_U280 = ~new_P2_U3077 | ~new_P2_U3956;
  assign new_P2_R1233_U281 = ~new_P2_R1233_U278 | ~new_P2_R1233_U279;
  assign new_P2_R1233_U282 = new_P2_U3483 | new_P2_U3084;
  assign new_P2_R1233_U283 = new_P2_U3956 | new_P2_U3077;
  assign new_P2_R1233_U284 = ~new_P2_R1233_U131 | ~new_P2_R1233_U273 | ~new_P2_R1233_U162;
  assign new_P2_R1233_U285 = ~new_P2_R1233_U283 | ~new_P2_R1233_U281;
  assign new_P2_R1233_U286 = ~new_P2_R1233_U159;
  assign new_P2_R1233_U287 = new_P2_U3955 | new_P2_U3063;
  assign new_P2_R1233_U288 = ~new_P2_R1233_U287 | ~new_P2_R1233_U159;
  assign new_P2_R1233_U289 = ~new_P2_U3063 | ~new_P2_U3955;
  assign new_P2_R1233_U290 = ~new_P2_R1233_U157;
  assign new_P2_R1233_U291 = new_P2_U3954 | new_P2_U3068;
  assign new_P2_R1233_U292 = ~new_P2_R1233_U291 | ~new_P2_R1233_U157;
  assign new_P2_R1233_U293 = ~new_P2_U3068 | ~new_P2_U3954;
  assign new_P2_R1233_U294 = ~new_P2_R1233_U155;
  assign new_P2_R1233_U295 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1233_U296 = ~new_P2_R1233_U176 | ~new_P2_R1233_U173;
  assign new_P2_R1233_U297 = ~new_P2_R1233_U86;
  assign new_P2_R1233_U298 = new_P2_U3953 | new_P2_U3067;
  assign new_P2_R1233_U299 = ~new_P2_R1233_U168 | ~new_P2_R1233_U155 | ~new_P2_R1233_U298;
  assign new_P2_R1233_U300 = ~new_P2_R1233_U153;
  assign new_P2_R1233_U301 = new_P2_U3950 | new_P2_U3055;
  assign new_P2_R1233_U302 = ~new_P2_U3055 | ~new_P2_U3950;
  assign new_P2_R1233_U303 = ~new_P2_R1233_U151;
  assign new_P2_R1233_U304 = ~new_P2_U3949 | ~new_P2_R1233_U151;
  assign new_P2_R1233_U305 = ~new_P2_R1233_U149;
  assign new_P2_R1233_U306 = ~new_P2_R1233_U298 | ~new_P2_R1233_U155;
  assign new_P2_R1233_U307 = ~new_P2_R1233_U89;
  assign new_P2_R1233_U308 = new_P2_U3952 | new_P2_U3060;
  assign new_P2_R1233_U309 = ~new_P2_R1233_U308 | ~new_P2_R1233_U89;
  assign new_P2_R1233_U310 = ~new_P2_R1233_U154 | ~new_P2_R1233_U309 | ~new_P2_R1233_U173;
  assign new_P2_R1233_U311 = ~new_P2_R1233_U307 | ~new_P2_R1233_U173;
  assign new_P2_R1233_U312 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1233_U313 = ~new_P2_R1233_U168 | ~new_P2_R1233_U311 | ~new_P2_R1233_U312;
  assign new_P2_R1233_U314 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1233_U315 = ~new_P2_R1233_U282 | ~new_P2_R1233_U162;
  assign new_P2_R1233_U316 = ~new_P2_R1233_U91;
  assign new_P2_R1233_U317 = ~new_P2_R1233_U9 | ~new_P2_R1233_U91;
  assign new_P2_R1233_U318 = ~new_P2_R1233_U135 | ~new_P2_R1233_U317;
  assign new_P2_R1233_U319 = ~new_P2_R1233_U317 | ~new_P2_R1233_U278;
  assign new_P2_R1233_U320 = ~new_P2_R1233_U453 | ~new_P2_R1233_U319;
  assign new_P2_R1233_U321 = new_P2_U3485 | new_P2_U3083;
  assign new_P2_R1233_U322 = ~new_P2_R1233_U321 | ~new_P2_R1233_U91;
  assign new_P2_R1233_U323 = ~new_P2_R1233_U136 | ~new_P2_R1233_U322;
  assign new_P2_R1233_U324 = ~new_P2_R1233_U316 | ~new_P2_R1233_U80;
  assign new_P2_R1233_U325 = ~new_P2_U3078 | ~new_P2_U3957;
  assign new_P2_R1233_U326 = ~new_P2_R1233_U137 | ~new_P2_R1233_U324;
  assign new_P2_R1233_U327 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1233_U328 = ~new_P2_R1233_U161;
  assign new_P2_R1233_U329 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1233_U330 = new_P2_U3477 | new_P2_U3075;
  assign new_P2_R1233_U331 = ~new_P2_R1233_U330 | ~new_P2_R1233_U92;
  assign new_P2_R1233_U332 = ~new_P2_R1233_U138 | ~new_P2_R1233_U331;
  assign new_P2_R1233_U333 = ~new_P2_R1233_U262 | ~new_P2_R1233_U59;
  assign new_P2_R1233_U334 = ~new_P2_U3480 | ~new_P2_U3071;
  assign new_P2_R1233_U335 = ~new_P2_R1233_U139 | ~new_P2_R1233_U333;
  assign new_P2_R1233_U336 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1233_U337 = ~new_P2_R1233_U250 | ~new_P2_R1233_U167;
  assign new_P2_R1233_U338 = ~new_P2_R1233_U93;
  assign new_P2_R1233_U339 = new_P2_U3465 | new_P2_U3074;
  assign new_P2_R1233_U340 = ~new_P2_R1233_U339 | ~new_P2_R1233_U93;
  assign new_P2_R1233_U341 = ~new_P2_R1233_U140 | ~new_P2_R1233_U340;
  assign new_P2_R1233_U342 = ~new_P2_R1233_U338 | ~new_P2_R1233_U172;
  assign new_P2_R1233_U343 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1233_U344 = ~new_P2_R1233_U141 | ~new_P2_R1233_U342;
  assign new_P2_R1233_U345 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1233_U346 = new_P2_U3456 | new_P2_U3085;
  assign new_P2_R1233_U347 = ~new_P2_R1233_U346 | ~new_P2_R1233_U40;
  assign new_P2_R1233_U348 = ~new_P2_R1233_U142 | ~new_P2_R1233_U347;
  assign new_P2_R1233_U349 = ~new_P2_R1233_U206 | ~new_P2_R1233_U171;
  assign new_P2_R1233_U350 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1233_U351 = ~new_P2_R1233_U143 | ~new_P2_R1233_U349;
  assign new_P2_R1233_U352 = ~new_P2_R1233_U207 | ~new_P2_R1233_U171;
  assign new_P2_R1233_U353 = ~new_P2_R1233_U204 | ~new_P2_R1233_U61;
  assign new_P2_R1233_U354 = ~new_P2_R1233_U214 | ~new_P2_R1233_U22;
  assign new_P2_R1233_U355 = ~new_P2_R1233_U228 | ~new_P2_R1233_U34;
  assign new_P2_R1233_U356 = ~new_P2_R1233_U231 | ~new_P2_R1233_U180;
  assign new_P2_R1233_U357 = ~new_P2_R1233_U314 | ~new_P2_R1233_U173;
  assign new_P2_R1233_U358 = ~new_P2_R1233_U298 | ~new_P2_R1233_U176;
  assign new_P2_R1233_U359 = ~new_P2_R1233_U329 | ~new_P2_R1233_U80;
  assign new_P2_R1233_U360 = ~new_P2_R1233_U282 | ~new_P2_R1233_U77;
  assign new_P2_R1233_U361 = ~new_P2_R1233_U336 | ~new_P2_R1233_U59;
  assign new_P2_R1233_U362 = ~new_P2_R1233_U345 | ~new_P2_R1233_U172;
  assign new_P2_R1233_U363 = ~new_P2_R1233_U250 | ~new_P2_R1233_U68;
  assign new_P2_R1233_U364 = ~new_P2_U3949 | ~new_P2_U3056;
  assign new_P2_R1233_U365 = ~new_P2_R1233_U296 | ~new_P2_R1233_U168;
  assign new_P2_R1233_U366 = ~new_P2_U3059 | ~new_P2_R1233_U295;
  assign new_P2_R1233_U367 = ~new_P2_U3951 | ~new_P2_R1233_U295;
  assign new_P2_R1233_U368 = ~new_P2_R1233_U301 | ~new_P2_R1233_U296 | ~new_P2_R1233_U168;
  assign new_P2_R1233_U369 = ~new_P2_R1233_U133 | ~new_P2_R1233_U155 | ~new_P2_R1233_U168;
  assign new_P2_R1233_U370 = ~new_P2_R1233_U297 | ~new_P2_R1233_U301;
  assign new_P2_R1233_U371 = ~new_P2_U3085 | ~new_P2_R1233_U39;
  assign new_P2_R1233_U372 = ~new_P2_U3456 | ~new_P2_R1233_U38;
  assign new_P2_R1233_U373 = ~new_P2_R1233_U372 | ~new_P2_R1233_U371;
  assign new_P2_R1233_U374 = ~new_P2_R1233_U352 | ~new_P2_R1233_U40;
  assign new_P2_R1233_U375 = ~new_P2_R1233_U373 | ~new_P2_R1233_U206;
  assign new_P2_R1233_U376 = ~new_P2_U3086 | ~new_P2_R1233_U36;
  assign new_P2_R1233_U377 = ~new_P2_U3453 | ~new_P2_R1233_U37;
  assign new_P2_R1233_U378 = ~new_P2_R1233_U377 | ~new_P2_R1233_U376;
  assign new_P2_R1233_U379 = ~new_P2_R1233_U353 | ~new_P2_R1233_U144;
  assign new_P2_R1233_U380 = ~new_P2_R1233_U203 | ~new_P2_R1233_U378;
  assign new_P2_R1233_U381 = ~new_P2_U3072 | ~new_P2_R1233_U23;
  assign new_P2_R1233_U382 = ~new_P2_U3450 | ~new_P2_R1233_U21;
  assign new_P2_R1233_U383 = ~new_P2_U3073 | ~new_P2_R1233_U19;
  assign new_P2_R1233_U384 = ~new_P2_U3447 | ~new_P2_R1233_U20;
  assign new_P2_R1233_U385 = ~new_P2_R1233_U384 | ~new_P2_R1233_U383;
  assign new_P2_R1233_U386 = ~new_P2_R1233_U354 | ~new_P2_R1233_U41;
  assign new_P2_R1233_U387 = ~new_P2_R1233_U385 | ~new_P2_R1233_U195;
  assign new_P2_R1233_U388 = ~new_P2_U3069 | ~new_P2_R1233_U35;
  assign new_P2_R1233_U389 = ~new_P2_U3444 | ~new_P2_R1233_U26;
  assign new_P2_R1233_U390 = ~new_P2_U3062 | ~new_P2_R1233_U24;
  assign new_P2_R1233_U391 = ~new_P2_U3441 | ~new_P2_R1233_U25;
  assign new_P2_R1233_U392 = ~new_P2_R1233_U391 | ~new_P2_R1233_U390;
  assign new_P2_R1233_U393 = ~new_P2_R1233_U355 | ~new_P2_R1233_U44;
  assign new_P2_R1233_U394 = ~new_P2_R1233_U392 | ~new_P2_R1233_U221;
  assign new_P2_R1233_U395 = ~new_P2_U3066 | ~new_P2_R1233_U32;
  assign new_P2_R1233_U396 = ~new_P2_U3438 | ~new_P2_R1233_U33;
  assign new_P2_R1233_U397 = ~new_P2_R1233_U396 | ~new_P2_R1233_U395;
  assign new_P2_R1233_U398 = ~new_P2_R1233_U356 | ~new_P2_R1233_U145;
  assign new_P2_R1233_U399 = ~new_P2_R1233_U230 | ~new_P2_R1233_U397;
  assign new_P2_R1233_U400 = ~new_P2_U3070 | ~new_P2_R1233_U27;
  assign new_P2_R1233_U401 = ~new_P2_U3435 | ~new_P2_R1233_U28;
  assign new_P2_R1233_U402 = ~new_P2_U3057 | ~new_P2_R1233_U147;
  assign new_P2_R1233_U403 = ~new_P2_U3960 | ~new_P2_R1233_U146;
  assign new_P2_R1233_U404 = ~new_P2_U3057 | ~new_P2_R1233_U147;
  assign new_P2_R1233_U405 = ~new_P2_U3960 | ~new_P2_R1233_U146;
  assign new_P2_R1233_U406 = ~new_P2_R1233_U405 | ~new_P2_R1233_U404;
  assign new_P2_R1233_U407 = ~new_P2_R1233_U148 | ~new_P2_R1233_U149;
  assign new_P2_R1233_U408 = ~new_P2_R1233_U305 | ~new_P2_R1233_U406;
  assign new_P2_R1233_U409 = ~new_P2_U3056 | ~new_P2_R1233_U88;
  assign new_P2_R1233_U410 = ~new_P2_U3949 | ~new_P2_R1233_U87;
  assign new_P2_R1233_U411 = ~new_P2_U3056 | ~new_P2_R1233_U88;
  assign new_P2_R1233_U412 = ~new_P2_U3949 | ~new_P2_R1233_U87;
  assign new_P2_R1233_U413 = ~new_P2_R1233_U412 | ~new_P2_R1233_U411;
  assign new_P2_R1233_U414 = ~new_P2_R1233_U150 | ~new_P2_R1233_U151;
  assign new_P2_R1233_U415 = ~new_P2_R1233_U303 | ~new_P2_R1233_U413;
  assign new_P2_R1233_U416 = ~new_P2_U3055 | ~new_P2_R1233_U46;
  assign new_P2_R1233_U417 = ~new_P2_U3950 | ~new_P2_R1233_U47;
  assign new_P2_R1233_U418 = ~new_P2_U3055 | ~new_P2_R1233_U46;
  assign new_P2_R1233_U419 = ~new_P2_U3950 | ~new_P2_R1233_U47;
  assign new_P2_R1233_U420 = ~new_P2_R1233_U419 | ~new_P2_R1233_U418;
  assign new_P2_R1233_U421 = ~new_P2_R1233_U152 | ~new_P2_R1233_U153;
  assign new_P2_R1233_U422 = ~new_P2_R1233_U300 | ~new_P2_R1233_U420;
  assign new_P2_R1233_U423 = ~new_P2_U3059 | ~new_P2_R1233_U49;
  assign new_P2_R1233_U424 = ~new_P2_U3951 | ~new_P2_R1233_U48;
  assign new_P2_R1233_U425 = ~new_P2_U3060 | ~new_P2_R1233_U50;
  assign new_P2_R1233_U426 = ~new_P2_U3952 | ~new_P2_R1233_U51;
  assign new_P2_R1233_U427 = ~new_P2_R1233_U426 | ~new_P2_R1233_U425;
  assign new_P2_R1233_U428 = ~new_P2_R1233_U357 | ~new_P2_R1233_U89;
  assign new_P2_R1233_U429 = ~new_P2_R1233_U427 | ~new_P2_R1233_U307;
  assign new_P2_R1233_U430 = ~new_P2_U3067 | ~new_P2_R1233_U52;
  assign new_P2_R1233_U431 = ~new_P2_U3953 | ~new_P2_R1233_U53;
  assign new_P2_R1233_U432 = ~new_P2_R1233_U431 | ~new_P2_R1233_U430;
  assign new_P2_R1233_U433 = ~new_P2_R1233_U358 | ~new_P2_R1233_U155;
  assign new_P2_R1233_U434 = ~new_P2_R1233_U294 | ~new_P2_R1233_U432;
  assign new_P2_R1233_U435 = ~new_P2_U3068 | ~new_P2_R1233_U84;
  assign new_P2_R1233_U436 = ~new_P2_U3954 | ~new_P2_R1233_U85;
  assign new_P2_R1233_U437 = ~new_P2_U3068 | ~new_P2_R1233_U84;
  assign new_P2_R1233_U438 = ~new_P2_U3954 | ~new_P2_R1233_U85;
  assign new_P2_R1233_U439 = ~new_P2_R1233_U438 | ~new_P2_R1233_U437;
  assign new_P2_R1233_U440 = ~new_P2_R1233_U156 | ~new_P2_R1233_U157;
  assign new_P2_R1233_U441 = ~new_P2_R1233_U290 | ~new_P2_R1233_U439;
  assign new_P2_R1233_U442 = ~new_P2_U3063 | ~new_P2_R1233_U82;
  assign new_P2_R1233_U443 = ~new_P2_U3955 | ~new_P2_R1233_U83;
  assign new_P2_R1233_U444 = ~new_P2_U3063 | ~new_P2_R1233_U82;
  assign new_P2_R1233_U445 = ~new_P2_U3955 | ~new_P2_R1233_U83;
  assign new_P2_R1233_U446 = ~new_P2_R1233_U445 | ~new_P2_R1233_U444;
  assign new_P2_R1233_U447 = ~new_P2_R1233_U158 | ~new_P2_R1233_U159;
  assign new_P2_R1233_U448 = ~new_P2_R1233_U286 | ~new_P2_R1233_U446;
  assign new_P2_R1233_U449 = ~new_P2_U3077 | ~new_P2_R1233_U54;
  assign new_P2_R1233_U450 = ~new_P2_U3956 | ~new_P2_R1233_U55;
  assign new_P2_R1233_U451 = ~new_P2_U3077 | ~new_P2_R1233_U54;
  assign new_P2_R1233_U452 = ~new_P2_U3956 | ~new_P2_R1233_U55;
  assign new_P2_R1233_U453 = ~new_P2_R1233_U452 | ~new_P2_R1233_U451;
  assign new_P2_R1233_U454 = ~new_P2_U3078 | ~new_P2_R1233_U81;
  assign new_P2_R1233_U455 = ~new_P2_U3957 | ~new_P2_R1233_U90;
  assign new_P2_R1233_U456 = ~new_P2_R1233_U182 | ~new_P2_R1233_U161;
  assign new_P2_R1233_U457 = ~new_P2_R1233_U328 | ~new_P2_R1233_U31;
  assign new_P2_R1233_U458 = ~new_P2_U3083 | ~new_P2_R1233_U78;
  assign new_P2_R1233_U459 = ~new_P2_U3485 | ~new_P2_R1233_U79;
  assign new_P2_R1233_U460 = ~new_P2_R1233_U459 | ~new_P2_R1233_U458;
  assign new_P2_R1233_U461 = ~new_P2_R1233_U359 | ~new_P2_R1233_U91;
  assign new_P2_R1233_U462 = ~new_P2_R1233_U460 | ~new_P2_R1233_U316;
  assign new_P2_R1233_U463 = ~new_P2_U3084 | ~new_P2_R1233_U75;
  assign new_P2_R1233_U464 = ~new_P2_U3483 | ~new_P2_R1233_U76;
  assign new_P2_R1233_U465 = ~new_P2_R1233_U464 | ~new_P2_R1233_U463;
  assign new_P2_R1233_U466 = ~new_P2_R1233_U360 | ~new_P2_R1233_U162;
  assign new_P2_R1233_U467 = ~new_P2_R1233_U270 | ~new_P2_R1233_U465;
  assign new_P2_R1233_U468 = ~new_P2_U3071 | ~new_P2_R1233_U60;
  assign new_P2_R1233_U469 = ~new_P2_U3480 | ~new_P2_R1233_U58;
  assign new_P2_R1233_U470 = ~new_P2_U3075 | ~new_P2_R1233_U56;
  assign new_P2_R1233_U471 = ~new_P2_U3477 | ~new_P2_R1233_U57;
  assign new_P2_R1233_U472 = ~new_P2_R1233_U471 | ~new_P2_R1233_U470;
  assign new_P2_R1233_U473 = ~new_P2_R1233_U361 | ~new_P2_R1233_U92;
  assign new_P2_R1233_U474 = ~new_P2_R1233_U472 | ~new_P2_R1233_U262;
  assign new_P2_R1233_U475 = ~new_P2_U3076 | ~new_P2_R1233_U73;
  assign new_P2_R1233_U476 = ~new_P2_U3474 | ~new_P2_R1233_U74;
  assign new_P2_R1233_U477 = ~new_P2_U3076 | ~new_P2_R1233_U73;
  assign new_P2_R1233_U478 = ~new_P2_U3474 | ~new_P2_R1233_U74;
  assign new_P2_R1233_U479 = ~new_P2_R1233_U478 | ~new_P2_R1233_U477;
  assign new_P2_R1233_U480 = ~new_P2_R1233_U163 | ~new_P2_R1233_U164;
  assign new_P2_R1233_U481 = ~new_P2_R1233_U258 | ~new_P2_R1233_U479;
  assign new_P2_R1233_U482 = ~new_P2_U3081 | ~new_P2_R1233_U71;
  assign new_P2_R1233_U483 = ~new_P2_U3471 | ~new_P2_R1233_U72;
  assign new_P2_R1233_U484 = ~new_P2_U3081 | ~new_P2_R1233_U71;
  assign new_P2_R1233_U485 = ~new_P2_U3471 | ~new_P2_R1233_U72;
  assign new_P2_R1233_U486 = ~new_P2_R1233_U485 | ~new_P2_R1233_U484;
  assign new_P2_R1233_U487 = ~new_P2_R1233_U165 | ~new_P2_R1233_U166;
  assign new_P2_R1233_U488 = ~new_P2_R1233_U254 | ~new_P2_R1233_U486;
  assign new_P2_R1233_U489 = ~new_P2_U3082 | ~new_P2_R1233_U69;
  assign new_P2_R1233_U490 = ~new_P2_U3468 | ~new_P2_R1233_U70;
  assign new_P2_R1233_U491 = ~new_P2_U3074 | ~new_P2_R1233_U64;
  assign new_P2_R1233_U492 = ~new_P2_U3465 | ~new_P2_R1233_U65;
  assign new_P2_R1233_U493 = ~new_P2_R1233_U492 | ~new_P2_R1233_U491;
  assign new_P2_R1233_U494 = ~new_P2_R1233_U362 | ~new_P2_R1233_U93;
  assign new_P2_R1233_U495 = ~new_P2_R1233_U493 | ~new_P2_R1233_U338;
  assign new_P2_R1233_U496 = ~new_P2_U3065 | ~new_P2_R1233_U66;
  assign new_P2_R1233_U497 = ~new_P2_U3462 | ~new_P2_R1233_U67;
  assign new_P2_R1233_U498 = ~new_P2_R1233_U497 | ~new_P2_R1233_U496;
  assign new_P2_R1233_U499 = ~new_P2_R1233_U363 | ~new_P2_R1233_U167;
  assign new_P2_R1233_U500 = ~new_P2_R1233_U244 | ~new_P2_R1233_U498;
  assign new_P2_R1233_U501 = ~new_P2_U3064 | ~new_P2_R1233_U62;
  assign new_P2_R1233_U502 = ~new_P2_U3459 | ~new_P2_R1233_U63;
  assign new_P2_R1233_U503 = ~new_P2_U3079 | ~new_P2_R1233_U29;
  assign new_P2_R1233_U504 = ~new_P2_U3427 | ~new_P2_R1233_U30;
  assign new_P2_R1176_U4 = new_P2_R1176_U221 & new_P2_R1176_U220;
  assign new_P2_R1176_U5 = new_P2_R1176_U234 & new_P2_R1176_U233;
  assign new_P2_R1176_U6 = new_P2_R1176_U264 & new_P2_R1176_U263;
  assign new_P2_R1176_U7 = new_P2_R1176_U280 & new_P2_R1176_U279;
  assign new_P2_R1176_U8 = new_P2_R1176_U292 & new_P2_R1176_U291;
  assign new_P2_R1176_U9 = new_P2_R1176_U6 & new_P2_R1176_U268;
  assign new_P2_R1176_U10 = new_P2_R1176_U5 & new_P2_R1176_U229;
  assign new_P2_R1176_U11 = new_P2_R1176_U9 & new_P2_R1176_U259;
  assign new_P2_R1176_U12 = new_P2_R1176_U528 & new_P2_R1176_U527;
  assign new_P2_R1176_U13 = new_P2_R1176_U351 & new_P2_R1176_U348;
  assign new_P2_R1176_U14 = new_P2_R1176_U342 & new_P2_R1176_U339;
  assign new_P2_R1176_U15 = new_P2_R1176_U335 & new_P2_R1176_U332;
  assign new_P2_R1176_U16 = new_P2_R1176_U385 & new_P2_R1176_U326 & new_P2_R1176_U323;
  assign new_P2_R1176_U17 = new_P2_R1176_U255 & new_P2_R1176_U252;
  assign new_P2_R1176_U18 = new_P2_R1176_U248 & new_P2_R1176_U245;
  assign new_P2_R1176_U19 = ~new_P2_U3184;
  assign new_P2_R1176_U20 = ~new_P2_U3175;
  assign new_P2_R1176_U21 = ~new_P2_U3181;
  assign new_P2_R1176_U22 = ~new_P2_U3181 | ~new_P2_R1176_U66;
  assign new_P2_R1176_U23 = ~new_P2_U3180;
  assign new_P2_R1176_U24 = ~new_P2_U3182;
  assign new_P2_R1176_U25 = ~new_P2_U3183;
  assign new_P2_R1176_U26 = ~new_P2_U3184 | ~new_P2_R1176_U69;
  assign new_P2_R1176_U27 = ~new_P2_U3179;
  assign new_P2_R1176_U28 = ~new_P2_U3177;
  assign new_P2_R1176_U29 = ~new_P2_U3177 | ~new_P2_R1176_U73;
  assign new_P2_R1176_U30 = ~new_P2_U3176;
  assign new_P2_R1176_U31 = ~new_P2_U3178;
  assign new_P2_R1176_U32 = ~new_P2_U3178 | ~new_P2_R1176_U71;
  assign new_P2_R1176_U33 = ~new_P2_U3174;
  assign new_P2_R1176_U34 = ~new_P2_R1176_U369 | ~new_P2_R1176_U238 | ~new_P2_R1176_U237;
  assign new_P2_R1176_U35 = ~new_P2_R1176_U32 | ~new_P2_R1176_U230;
  assign new_P2_R1176_U36 = ~new_P2_R1176_U365 | ~new_P2_R1176_U366 | ~new_P2_R1176_U218;
  assign new_P2_R1176_U37 = ~new_P2_U3156;
  assign new_P2_R1176_U38 = ~new_P2_U3158;
  assign new_P2_R1176_U39 = ~new_P2_U3159;
  assign new_P2_R1176_U40 = ~new_P2_U3157;
  assign new_P2_R1176_U41 = ~new_P2_U3167;
  assign new_P2_R1176_U42 = ~new_P2_U3167 | ~new_P2_R1176_U78;
  assign new_P2_R1176_U43 = ~new_P2_U3166;
  assign new_P2_R1176_U44 = ~new_P2_U3169;
  assign new_P2_R1176_U45 = ~new_P2_U3171;
  assign new_P2_R1176_U46 = ~new_P2_U3172;
  assign new_P2_R1176_U47 = ~new_P2_U3172 | ~new_P2_R1176_U82;
  assign new_P2_R1176_U48 = ~new_P2_U3170;
  assign new_P2_R1176_U49 = ~new_P2_U3173;
  assign new_P2_R1176_U50 = ~new_P2_U3173 | ~new_P2_R1176_U81;
  assign new_P2_R1176_U51 = ~new_P2_U3168;
  assign new_P2_R1176_U52 = ~new_P2_U3165;
  assign new_P2_R1176_U53 = ~new_P2_U3163;
  assign new_P2_R1176_U54 = ~new_P2_U3164;
  assign new_P2_R1176_U55 = ~new_P2_U3164 | ~new_P2_R1176_U87;
  assign new_P2_R1176_U56 = ~new_P2_U3162;
  assign new_P2_R1176_U57 = ~new_P2_U3161;
  assign new_P2_R1176_U58 = ~new_P2_U3160;
  assign new_P2_R1176_U59 = ~new_P2_R1176_U212 | ~new_P2_R1176_U321;
  assign new_P2_R1176_U60 = ~new_P2_R1176_U55 | ~new_P2_R1176_U328;
  assign new_P2_R1176_U61 = ~new_P2_R1176_U277 | ~new_P2_R1176_U276;
  assign new_P2_R1176_U62 = ~new_P2_R1176_U374 | ~new_P2_R1176_U270;
  assign new_P2_R1176_U63 = ~new_P2_R1176_U47 | ~new_P2_R1176_U344;
  assign new_P2_R1176_U64 = ~new_P2_R1176_U387 | ~new_P2_R1176_U386;
  assign new_P2_R1176_U65 = ~new_P2_R1176_U419 | ~new_P2_R1176_U418;
  assign new_P2_R1176_U66 = ~new_P2_R1176_U407 | ~new_P2_R1176_U406;
  assign new_P2_R1176_U67 = ~new_P2_R1176_U404 | ~new_P2_R1176_U403;
  assign new_P2_R1176_U68 = ~new_P2_R1176_U398 | ~new_P2_R1176_U397;
  assign new_P2_R1176_U69 = ~new_P2_R1176_U401 | ~new_P2_R1176_U400;
  assign new_P2_R1176_U70 = ~new_P2_R1176_U395 | ~new_P2_R1176_U394;
  assign new_P2_R1176_U71 = ~new_P2_R1176_U410 | ~new_P2_R1176_U409;
  assign new_P2_R1176_U72 = ~new_P2_R1176_U413 | ~new_P2_R1176_U412;
  assign new_P2_R1176_U73 = ~new_P2_R1176_U416 | ~new_P2_R1176_U415;
  assign new_P2_R1176_U74 = ~new_P2_R1176_U459 | ~new_P2_R1176_U458;
  assign new_P2_R1176_U75 = ~new_P2_R1176_U507 | ~new_P2_R1176_U506;
  assign new_P2_R1176_U76 = ~new_P2_R1176_U510 | ~new_P2_R1176_U509;
  assign new_P2_R1176_U77 = ~new_P2_R1176_U462 | ~new_P2_R1176_U461;
  assign new_P2_R1176_U78 = ~new_P2_R1176_U486 | ~new_P2_R1176_U485;
  assign new_P2_R1176_U79 = ~new_P2_R1176_U483 | ~new_P2_R1176_U482;
  assign new_P2_R1176_U80 = ~new_P2_R1176_U477 | ~new_P2_R1176_U476;
  assign new_P2_R1176_U81 = ~new_P2_R1176_U465 | ~new_P2_R1176_U464;
  assign new_P2_R1176_U82 = ~new_P2_R1176_U468 | ~new_P2_R1176_U467;
  assign new_P2_R1176_U83 = ~new_P2_R1176_U471 | ~new_P2_R1176_U470;
  assign new_P2_R1176_U84 = ~new_P2_R1176_U474 | ~new_P2_R1176_U473;
  assign new_P2_R1176_U85 = ~new_P2_R1176_U480 | ~new_P2_R1176_U479;
  assign new_P2_R1176_U86 = ~new_P2_R1176_U489 | ~new_P2_R1176_U488;
  assign new_P2_R1176_U87 = ~new_P2_R1176_U498 | ~new_P2_R1176_U497;
  assign new_P2_R1176_U88 = ~new_P2_R1176_U492 | ~new_P2_R1176_U491;
  assign new_P2_R1176_U89 = ~new_P2_R1176_U495 | ~new_P2_R1176_U494;
  assign new_P2_R1176_U90 = ~new_P2_R1176_U501 | ~new_P2_R1176_U500;
  assign new_P2_R1176_U91 = ~new_P2_R1176_U504 | ~new_P2_R1176_U503;
  assign new_P2_R1176_U92 = ~new_P2_R1176_U516 | ~new_P2_R1176_U515;
  assign new_P2_R1176_U93 = ~new_P2_R1176_U623 | ~new_P2_R1176_U622;
  assign new_P2_R1176_U94 = ~new_P2_R1176_U422 | ~new_P2_R1176_U421;
  assign new_P2_R1176_U95 = ~new_P2_R1176_U429 | ~new_P2_R1176_U428;
  assign new_P2_R1176_U96 = ~new_P2_R1176_U436 | ~new_P2_R1176_U435;
  assign new_P2_R1176_U97 = ~new_P2_R1176_U443 | ~new_P2_R1176_U442;
  assign new_P2_R1176_U98 = ~new_P2_R1176_U450 | ~new_P2_R1176_U449;
  assign new_P2_R1176_U99 = ~new_P2_R1176_U457 | ~new_P2_R1176_U456;
  assign new_P2_R1176_U100 = ~new_P2_R1176_U519 | ~new_P2_R1176_U518;
  assign new_P2_R1176_U101 = ~new_P2_R1176_U526 | ~new_P2_R1176_U525;
  assign new_P2_R1176_U102 = ~new_P2_R1176_U533 | ~new_P2_R1176_U532;
  assign new_P2_R1176_U103 = ~new_P2_R1176_U538 | ~new_P2_R1176_U537;
  assign new_P2_R1176_U104 = ~new_P2_R1176_U545 | ~new_P2_R1176_U544;
  assign new_P2_R1176_U105 = ~new_P2_R1176_U552 | ~new_P2_R1176_U551;
  assign new_P2_R1176_U106 = ~new_P2_R1176_U559 | ~new_P2_R1176_U558;
  assign new_P2_R1176_U107 = ~new_P2_R1176_U566 | ~new_P2_R1176_U565;
  assign new_P2_R1176_U108 = ~new_P2_R1176_U571 | ~new_P2_R1176_U570;
  assign new_P2_R1176_U109 = ~new_P2_R1176_U578 | ~new_P2_R1176_U577;
  assign new_P2_R1176_U110 = ~new_P2_R1176_U585 | ~new_P2_R1176_U584;
  assign new_P2_R1176_U111 = ~new_P2_R1176_U592 | ~new_P2_R1176_U591;
  assign new_P2_R1176_U112 = ~new_P2_R1176_U599 | ~new_P2_R1176_U598;
  assign new_P2_R1176_U113 = ~new_P2_R1176_U606 | ~new_P2_R1176_U605;
  assign new_P2_R1176_U114 = ~new_P2_R1176_U611 | ~new_P2_R1176_U610;
  assign new_P2_R1176_U115 = ~new_P2_R1176_U618 | ~new_P2_R1176_U617;
  assign new_P2_R1176_U116 = new_P2_R1176_U224 & new_P2_R1176_U223;
  assign new_P2_R1176_U117 = new_P2_R1176_U240 & new_P2_R1176_U10;
  assign new_P2_R1176_U118 = new_P2_R1176_U372 & new_P2_R1176_U241;
  assign new_P2_R1176_U119 = new_P2_R1176_U29 & new_P2_R1176_U431 & new_P2_R1176_U430;
  assign new_P2_R1176_U120 = new_P2_R1176_U247 & new_P2_R1176_U5;
  assign new_P2_R1176_U121 = new_P2_R1176_U22 & new_P2_R1176_U452 & new_P2_R1176_U451;
  assign new_P2_R1176_U122 = new_P2_R1176_U254 & new_P2_R1176_U4;
  assign new_P2_R1176_U123 = new_P2_R1176_U272 & new_P2_R1176_U11;
  assign new_P2_R1176_U124 = new_P2_R1176_U266 & new_P2_R1176_U207;
  assign new_P2_R1176_U125 = new_P2_R1176_U380 & new_P2_R1176_U273;
  assign new_P2_R1176_U126 = new_P2_R1176_U284 & new_P2_R1176_U283;
  assign new_P2_R1176_U127 = new_P2_R1176_U296 & new_P2_R1176_U8;
  assign new_P2_R1176_U128 = new_P2_R1176_U294 & new_P2_R1176_U208;
  assign new_P2_R1176_U129 = new_P2_R1176_U312 & new_P2_R1176_U203;
  assign new_P2_R1176_U130 = new_P2_R1176_U383 & new_P2_R1176_U318;
  assign new_P2_R1176_U131 = new_P2_R1176_U320 & new_P2_R1176_U310;
  assign new_P2_R1176_U132 = new_P2_R1176_U320 & new_P2_R1176_U312;
  assign new_P2_R1176_U133 = new_P2_R1176_U381 & new_P2_R1176_U319;
  assign new_P2_R1176_U134 = ~new_P2_R1176_U513 | ~new_P2_R1176_U512;
  assign new_P2_R1176_U135 = new_P2_R1176_U508 & new_P2_R1176_U38;
  assign new_P2_R1176_U136 = new_P2_R1176_U212 & new_P2_R1176_U209;
  assign new_P2_R1176_U137 = new_P2_R1176_U325 & new_P2_R1176_U203;
  assign new_P2_R1176_U138 = new_P2_R1176_U12 & new_P2_R1176_U209;
  assign new_P2_R1176_U139 = new_P2_R1176_U208 & new_P2_R1176_U554 & new_P2_R1176_U553;
  assign new_P2_R1176_U140 = new_P2_R1176_U334 & new_P2_R1176_U8;
  assign new_P2_R1176_U141 = new_P2_R1176_U42 & new_P2_R1176_U580 & new_P2_R1176_U579;
  assign new_P2_R1176_U142 = new_P2_R1176_U341 & new_P2_R1176_U7;
  assign new_P2_R1176_U143 = new_P2_R1176_U207 & new_P2_R1176_U601 & new_P2_R1176_U600;
  assign new_P2_R1176_U144 = new_P2_R1176_U350 & new_P2_R1176_U6;
  assign new_P2_R1176_U145 = ~new_P2_R1176_U620 | ~new_P2_R1176_U619;
  assign new_P2_R1176_U146 = ~new_P2_U3456;
  assign new_P2_R1176_U147 = new_P2_R1176_U390 & new_P2_R1176_U389;
  assign new_P2_R1176_U148 = ~new_P2_U3441;
  assign new_P2_R1176_U149 = ~new_P2_U3432;
  assign new_P2_R1176_U150 = ~new_P2_U3427;
  assign new_P2_R1176_U151 = ~new_P2_U3438;
  assign new_P2_R1176_U152 = ~new_P2_U3435;
  assign new_P2_R1176_U153 = ~new_P2_U3444;
  assign new_P2_R1176_U154 = ~new_P2_U3450;
  assign new_P2_R1176_U155 = ~new_P2_U3447;
  assign new_P2_R1176_U156 = ~new_P2_U3453;
  assign new_P2_R1176_U157 = ~new_P2_R1176_U118 | ~new_P2_R1176_U371;
  assign new_P2_R1176_U158 = new_P2_R1176_U424 & new_P2_R1176_U423;
  assign new_P2_R1176_U159 = ~new_P2_R1176_U370 | ~new_P2_R1176_U368;
  assign new_P2_R1176_U160 = new_P2_R1176_U438 & new_P2_R1176_U437;
  assign new_P2_R1176_U161 = ~new_P2_R1176_U362 | ~new_P2_R1176_U227 | ~new_P2_R1176_U205;
  assign new_P2_R1176_U162 = new_P2_R1176_U445 & new_P2_R1176_U444;
  assign new_P2_R1176_U163 = ~new_P2_R1176_U116 | ~new_P2_R1176_U225;
  assign new_P2_R1176_U164 = ~new_P2_U3950;
  assign new_P2_R1176_U165 = ~new_P2_U3951;
  assign new_P2_R1176_U166 = ~new_P2_U3459;
  assign new_P2_R1176_U167 = ~new_P2_U3462;
  assign new_P2_R1176_U168 = ~new_P2_U3468;
  assign new_P2_R1176_U169 = ~new_P2_U3465;
  assign new_P2_R1176_U170 = ~new_P2_U3471;
  assign new_P2_R1176_U171 = ~new_P2_U3474;
  assign new_P2_R1176_U172 = ~new_P2_U3480;
  assign new_P2_R1176_U173 = ~new_P2_U3477;
  assign new_P2_R1176_U174 = ~new_P2_U3483;
  assign new_P2_R1176_U175 = ~new_P2_U3956;
  assign new_P2_R1176_U176 = ~new_P2_U3957;
  assign new_P2_R1176_U177 = ~new_P2_U3485;
  assign new_P2_R1176_U178 = ~new_P2_U3955;
  assign new_P2_R1176_U179 = ~new_P2_U3954;
  assign new_P2_R1176_U180 = ~new_P2_U3952;
  assign new_P2_R1176_U181 = ~new_P2_U3953;
  assign new_P2_R1176_U182 = ~new_P2_U3949;
  assign new_P2_R1176_U183 = ~new_P2_U3155;
  assign new_P2_R1176_U184 = new_P2_R1176_U521 & new_P2_R1176_U520;
  assign new_P2_R1176_U185 = ~new_P2_R1176_U315 | ~new_P2_R1176_U314;
  assign new_P2_R1176_U186 = ~new_P2_R1176_U307 | ~new_P2_R1176_U306;
  assign new_P2_R1176_U187 = new_P2_R1176_U540 & new_P2_R1176_U539;
  assign new_P2_R1176_U188 = ~new_P2_R1176_U303 | ~new_P2_R1176_U302;
  assign new_P2_R1176_U189 = new_P2_R1176_U547 & new_P2_R1176_U546;
  assign new_P2_R1176_U190 = ~new_P2_R1176_U299 | ~new_P2_R1176_U298;
  assign new_P2_R1176_U191 = new_P2_R1176_U561 & new_P2_R1176_U560;
  assign new_P2_R1176_U192 = ~new_P2_R1176_U26 | ~new_P2_R1176_U214;
  assign new_P2_R1176_U193 = ~new_P2_R1176_U289 | ~new_P2_R1176_U288;
  assign new_P2_R1176_U194 = new_P2_R1176_U573 & new_P2_R1176_U572;
  assign new_P2_R1176_U195 = ~new_P2_R1176_U126 | ~new_P2_R1176_U285;
  assign new_P2_R1176_U196 = new_P2_R1176_U587 & new_P2_R1176_U586;
  assign new_P2_R1176_U197 = ~new_P2_R1176_U125 | ~new_P2_R1176_U379;
  assign new_P2_R1176_U198 = new_P2_R1176_U594 & new_P2_R1176_U593;
  assign new_P2_R1176_U199 = ~new_P2_R1176_U378 | ~new_P2_R1176_U373;
  assign new_P2_R1176_U200 = ~new_P2_R1176_U50 | ~new_P2_R1176_U260;
  assign new_P2_R1176_U201 = new_P2_R1176_U613 & new_P2_R1176_U612;
  assign new_P2_R1176_U202 = ~new_P2_R1176_U363 | ~new_P2_R1176_U257 | ~new_P2_R1176_U204;
  assign new_P2_R1176_U203 = ~new_P2_R1176_U377 | ~new_P2_R1176_U376;
  assign new_P2_R1176_U204 = ~new_P2_R1176_U64 | ~new_P2_R1176_U157;
  assign new_P2_R1176_U205 = ~new_P2_R1176_U70 | ~new_P2_R1176_U163;
  assign new_P2_R1176_U206 = ~new_P2_R1176_U22;
  assign new_P2_R1176_U207 = ~new_P2_U3171 | ~new_P2_R1176_U84;
  assign new_P2_R1176_U208 = ~new_P2_U3163 | ~new_P2_R1176_U89;
  assign new_P2_R1176_U209 = ~new_P2_U3158 | ~new_P2_R1176_U75;
  assign new_P2_R1176_U210 = ~new_P2_R1176_U47;
  assign new_P2_R1176_U211 = ~new_P2_R1176_U55;
  assign new_P2_R1176_U212 = ~new_P2_U3159 | ~new_P2_R1176_U76;
  assign new_P2_R1176_U213 = ~new_P2_R1176_U402 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U214 = ~new_P2_U3183 | ~new_P2_R1176_U213;
  assign new_P2_R1176_U215 = ~new_P2_R1176_U26;
  assign new_P2_R1176_U216 = ~new_P2_R1176_U192;
  assign new_P2_R1176_U217 = ~new_P2_R1176_U399 | ~new_P2_R1176_U24;
  assign new_P2_R1176_U218 = ~new_P2_U3182 | ~new_P2_R1176_U68;
  assign new_P2_R1176_U219 = ~new_P2_R1176_U36;
  assign new_P2_R1176_U220 = ~new_P2_R1176_U405 | ~new_P2_R1176_U23;
  assign new_P2_R1176_U221 = ~new_P2_R1176_U408 | ~new_P2_R1176_U21;
  assign new_P2_R1176_U222 = ~new_P2_R1176_U23 | ~new_P2_R1176_U22;
  assign new_P2_R1176_U223 = ~new_P2_R1176_U67 | ~new_P2_R1176_U222;
  assign new_P2_R1176_U224 = ~new_P2_U3180 | ~new_P2_R1176_U206;
  assign new_P2_R1176_U225 = ~new_P2_R1176_U4 | ~new_P2_R1176_U36;
  assign new_P2_R1176_U226 = ~new_P2_R1176_U163;
  assign new_P2_R1176_U227 = ~new_P2_U3179 | ~new_P2_R1176_U163;
  assign new_P2_R1176_U228 = ~new_P2_R1176_U161;
  assign new_P2_R1176_U229 = ~new_P2_R1176_U411 | ~new_P2_R1176_U31;
  assign new_P2_R1176_U230 = ~new_P2_R1176_U229 | ~new_P2_R1176_U161;
  assign new_P2_R1176_U231 = ~new_P2_R1176_U32;
  assign new_P2_R1176_U232 = ~new_P2_R1176_U35;
  assign new_P2_R1176_U233 = ~new_P2_R1176_U414 | ~new_P2_R1176_U30;
  assign new_P2_R1176_U234 = ~new_P2_R1176_U417 | ~new_P2_R1176_U28;
  assign new_P2_R1176_U235 = ~new_P2_R1176_U29;
  assign new_P2_R1176_U236 = ~new_P2_R1176_U30 | ~new_P2_R1176_U29;
  assign new_P2_R1176_U237 = ~new_P2_R1176_U72 | ~new_P2_R1176_U236;
  assign new_P2_R1176_U238 = ~new_P2_U3176 | ~new_P2_R1176_U235;
  assign new_P2_R1176_U239 = ~new_P2_R1176_U159;
  assign new_P2_R1176_U240 = ~new_P2_R1176_U420 | ~new_P2_R1176_U20;
  assign new_P2_R1176_U241 = ~new_P2_U3175 | ~new_P2_R1176_U65;
  assign new_P2_R1176_U242 = ~new_P2_R1176_U157;
  assign new_P2_R1176_U243 = ~new_P2_R1176_U417 | ~new_P2_R1176_U28;
  assign new_P2_R1176_U244 = ~new_P2_R1176_U243 | ~new_P2_R1176_U35;
  assign new_P2_R1176_U245 = ~new_P2_R1176_U119 | ~new_P2_R1176_U244;
  assign new_P2_R1176_U246 = ~new_P2_R1176_U232 | ~new_P2_R1176_U29;
  assign new_P2_R1176_U247 = ~new_P2_U3176 | ~new_P2_R1176_U72;
  assign new_P2_R1176_U248 = ~new_P2_R1176_U120 | ~new_P2_R1176_U246;
  assign new_P2_R1176_U249 = ~new_P2_R1176_U417 | ~new_P2_R1176_U28;
  assign new_P2_R1176_U250 = ~new_P2_R1176_U408 | ~new_P2_R1176_U21;
  assign new_P2_R1176_U251 = ~new_P2_R1176_U250 | ~new_P2_R1176_U36;
  assign new_P2_R1176_U252 = ~new_P2_R1176_U121 | ~new_P2_R1176_U251;
  assign new_P2_R1176_U253 = ~new_P2_R1176_U219 | ~new_P2_R1176_U22;
  assign new_P2_R1176_U254 = ~new_P2_U3180 | ~new_P2_R1176_U67;
  assign new_P2_R1176_U255 = ~new_P2_R1176_U122 | ~new_P2_R1176_U253;
  assign new_P2_R1176_U256 = ~new_P2_R1176_U408 | ~new_P2_R1176_U21;
  assign new_P2_R1176_U257 = ~new_P2_U3174 | ~new_P2_R1176_U157;
  assign new_P2_R1176_U258 = ~new_P2_R1176_U202;
  assign new_P2_R1176_U259 = ~new_P2_R1176_U466 | ~new_P2_R1176_U49;
  assign new_P2_R1176_U260 = ~new_P2_R1176_U259 | ~new_P2_R1176_U202;
  assign new_P2_R1176_U261 = ~new_P2_R1176_U50;
  assign new_P2_R1176_U262 = ~new_P2_R1176_U200;
  assign new_P2_R1176_U263 = ~new_P2_R1176_U472 | ~new_P2_R1176_U48;
  assign new_P2_R1176_U264 = ~new_P2_R1176_U475 | ~new_P2_R1176_U45;
  assign new_P2_R1176_U265 = ~new_P2_R1176_U210 | ~new_P2_R1176_U6;
  assign new_P2_R1176_U266 = ~new_P2_U3170 | ~new_P2_R1176_U83;
  assign new_P2_R1176_U267 = ~new_P2_R1176_U124 | ~new_P2_R1176_U265;
  assign new_P2_R1176_U268 = ~new_P2_R1176_U469 | ~new_P2_R1176_U46;
  assign new_P2_R1176_U269 = ~new_P2_R1176_U472 | ~new_P2_R1176_U48;
  assign new_P2_R1176_U270 = ~new_P2_R1176_U269 | ~new_P2_R1176_U267;
  assign new_P2_R1176_U271 = ~new_P2_R1176_U199;
  assign new_P2_R1176_U272 = ~new_P2_R1176_U478 | ~new_P2_R1176_U44;
  assign new_P2_R1176_U273 = ~new_P2_U3169 | ~new_P2_R1176_U80;
  assign new_P2_R1176_U274 = ~new_P2_R1176_U197;
  assign new_P2_R1176_U275 = ~new_P2_R1176_U481 | ~new_P2_R1176_U51;
  assign new_P2_R1176_U276 = ~new_P2_R1176_U275 | ~new_P2_R1176_U197;
  assign new_P2_R1176_U277 = ~new_P2_U3168 | ~new_P2_R1176_U85;
  assign new_P2_R1176_U278 = ~new_P2_R1176_U61;
  assign new_P2_R1176_U279 = ~new_P2_R1176_U484 | ~new_P2_R1176_U43;
  assign new_P2_R1176_U280 = ~new_P2_R1176_U487 | ~new_P2_R1176_U41;
  assign new_P2_R1176_U281 = ~new_P2_R1176_U42;
  assign new_P2_R1176_U282 = ~new_P2_R1176_U43 | ~new_P2_R1176_U42;
  assign new_P2_R1176_U283 = ~new_P2_R1176_U79 | ~new_P2_R1176_U282;
  assign new_P2_R1176_U284 = ~new_P2_U3166 | ~new_P2_R1176_U281;
  assign new_P2_R1176_U285 = ~new_P2_R1176_U7 | ~new_P2_R1176_U61;
  assign new_P2_R1176_U286 = ~new_P2_R1176_U195;
  assign new_P2_R1176_U287 = ~new_P2_R1176_U490 | ~new_P2_R1176_U52;
  assign new_P2_R1176_U288 = ~new_P2_R1176_U287 | ~new_P2_R1176_U195;
  assign new_P2_R1176_U289 = ~new_P2_U3165 | ~new_P2_R1176_U86;
  assign new_P2_R1176_U290 = ~new_P2_R1176_U193;
  assign new_P2_R1176_U291 = ~new_P2_R1176_U493 | ~new_P2_R1176_U56;
  assign new_P2_R1176_U292 = ~new_P2_R1176_U496 | ~new_P2_R1176_U53;
  assign new_P2_R1176_U293 = ~new_P2_R1176_U211 | ~new_P2_R1176_U8;
  assign new_P2_R1176_U294 = ~new_P2_U3162 | ~new_P2_R1176_U88;
  assign new_P2_R1176_U295 = ~new_P2_R1176_U128 | ~new_P2_R1176_U293;
  assign new_P2_R1176_U296 = ~new_P2_R1176_U499 | ~new_P2_R1176_U54;
  assign new_P2_R1176_U297 = ~new_P2_R1176_U493 | ~new_P2_R1176_U56;
  assign new_P2_R1176_U298 = ~new_P2_R1176_U127 | ~new_P2_R1176_U193;
  assign new_P2_R1176_U299 = ~new_P2_R1176_U297 | ~new_P2_R1176_U295;
  assign new_P2_R1176_U300 = ~new_P2_R1176_U190;
  assign new_P2_R1176_U301 = ~new_P2_R1176_U502 | ~new_P2_R1176_U57;
  assign new_P2_R1176_U302 = ~new_P2_R1176_U301 | ~new_P2_R1176_U190;
  assign new_P2_R1176_U303 = ~new_P2_U3161 | ~new_P2_R1176_U90;
  assign new_P2_R1176_U304 = ~new_P2_R1176_U188;
  assign new_P2_R1176_U305 = ~new_P2_R1176_U505 | ~new_P2_R1176_U58;
  assign new_P2_R1176_U306 = ~new_P2_R1176_U305 | ~new_P2_R1176_U188;
  assign new_P2_R1176_U307 = ~new_P2_U3160 | ~new_P2_R1176_U91;
  assign new_P2_R1176_U308 = ~new_P2_R1176_U186;
  assign new_P2_R1176_U309 = ~new_P2_R1176_U508 | ~new_P2_R1176_U38;
  assign new_P2_R1176_U310 = ~new_P2_R1176_U311 | ~new_P2_R1176_U212 | ~new_P2_R1176_U209;
  assign new_P2_R1176_U311 = ~new_P2_U3157 | ~new_P2_R1176_U77;
  assign new_P2_R1176_U312 = ~new_P2_R1176_U511 | ~new_P2_R1176_U39;
  assign new_P2_R1176_U313 = ~new_P2_R1176_U463 | ~new_P2_R1176_U40;
  assign new_P2_R1176_U314 = ~new_P2_R1176_U129 | ~new_P2_R1176_U186;
  assign new_P2_R1176_U315 = ~new_P2_R1176_U375 | ~new_P2_R1176_U310;
  assign new_P2_R1176_U316 = ~new_P2_R1176_U185;
  assign new_P2_R1176_U317 = ~new_P2_R1176_U460 | ~new_P2_R1176_U37;
  assign new_P2_R1176_U318 = ~new_P2_U3156 | ~new_P2_R1176_U74;
  assign new_P2_R1176_U319 = ~new_P2_U3156 | ~new_P2_R1176_U74;
  assign new_P2_R1176_U320 = ~new_P2_R1176_U460 | ~new_P2_R1176_U37;
  assign new_P2_R1176_U321 = ~new_P2_R1176_U312 | ~new_P2_R1176_U186;
  assign new_P2_R1176_U322 = ~new_P2_R1176_U59;
  assign new_P2_R1176_U323 = ~new_P2_R1176_U135 | ~new_P2_R1176_U12;
  assign new_P2_R1176_U324 = ~new_P2_R1176_U136 | ~new_P2_R1176_U321;
  assign new_P2_R1176_U325 = ~new_P2_U3157 | ~new_P2_R1176_U77;
  assign new_P2_R1176_U326 = ~new_P2_R1176_U137 | ~new_P2_R1176_U324;
  assign new_P2_R1176_U327 = ~new_P2_R1176_U508 | ~new_P2_R1176_U38;
  assign new_P2_R1176_U328 = ~new_P2_R1176_U296 | ~new_P2_R1176_U193;
  assign new_P2_R1176_U329 = ~new_P2_R1176_U60;
  assign new_P2_R1176_U330 = ~new_P2_R1176_U496 | ~new_P2_R1176_U53;
  assign new_P2_R1176_U331 = ~new_P2_R1176_U330 | ~new_P2_R1176_U60;
  assign new_P2_R1176_U332 = ~new_P2_R1176_U139 | ~new_P2_R1176_U331;
  assign new_P2_R1176_U333 = ~new_P2_R1176_U329 | ~new_P2_R1176_U208;
  assign new_P2_R1176_U334 = ~new_P2_U3162 | ~new_P2_R1176_U88;
  assign new_P2_R1176_U335 = ~new_P2_R1176_U140 | ~new_P2_R1176_U333;
  assign new_P2_R1176_U336 = ~new_P2_R1176_U496 | ~new_P2_R1176_U53;
  assign new_P2_R1176_U337 = ~new_P2_R1176_U487 | ~new_P2_R1176_U41;
  assign new_P2_R1176_U338 = ~new_P2_R1176_U337 | ~new_P2_R1176_U61;
  assign new_P2_R1176_U339 = ~new_P2_R1176_U141 | ~new_P2_R1176_U338;
  assign new_P2_R1176_U340 = ~new_P2_R1176_U278 | ~new_P2_R1176_U42;
  assign new_P2_R1176_U341 = ~new_P2_U3166 | ~new_P2_R1176_U79;
  assign new_P2_R1176_U342 = ~new_P2_R1176_U142 | ~new_P2_R1176_U340;
  assign new_P2_R1176_U343 = ~new_P2_R1176_U487 | ~new_P2_R1176_U41;
  assign new_P2_R1176_U344 = ~new_P2_R1176_U268 | ~new_P2_R1176_U200;
  assign new_P2_R1176_U345 = ~new_P2_R1176_U63;
  assign new_P2_R1176_U346 = ~new_P2_R1176_U475 | ~new_P2_R1176_U45;
  assign new_P2_R1176_U347 = ~new_P2_R1176_U346 | ~new_P2_R1176_U63;
  assign new_P2_R1176_U348 = ~new_P2_R1176_U143 | ~new_P2_R1176_U347;
  assign new_P2_R1176_U349 = ~new_P2_R1176_U345 | ~new_P2_R1176_U207;
  assign new_P2_R1176_U350 = ~new_P2_U3170 | ~new_P2_R1176_U83;
  assign new_P2_R1176_U351 = ~new_P2_R1176_U144 | ~new_P2_R1176_U349;
  assign new_P2_R1176_U352 = ~new_P2_R1176_U475 | ~new_P2_R1176_U45;
  assign new_P2_R1176_U353 = ~new_P2_R1176_U249 | ~new_P2_R1176_U29;
  assign new_P2_R1176_U354 = ~new_P2_R1176_U256 | ~new_P2_R1176_U22;
  assign new_P2_R1176_U355 = ~new_P2_R1176_U327 | ~new_P2_R1176_U209;
  assign new_P2_R1176_U356 = ~new_P2_R1176_U312 | ~new_P2_R1176_U212;
  assign new_P2_R1176_U357 = ~new_P2_R1176_U336 | ~new_P2_R1176_U208;
  assign new_P2_R1176_U358 = ~new_P2_R1176_U296 | ~new_P2_R1176_U55;
  assign new_P2_R1176_U359 = ~new_P2_R1176_U343 | ~new_P2_R1176_U42;
  assign new_P2_R1176_U360 = ~new_P2_R1176_U352 | ~new_P2_R1176_U207;
  assign new_P2_R1176_U361 = ~new_P2_R1176_U268 | ~new_P2_R1176_U47;
  assign new_P2_R1176_U362 = ~new_P2_U3179 | ~new_P2_R1176_U70;
  assign new_P2_R1176_U363 = ~new_P2_U3174 | ~new_P2_R1176_U64;
  assign new_P2_R1176_U364 = ~new_P2_R1176_U130 | ~new_P2_R1176_U314 | ~new_P2_R1176_U311;
  assign new_P2_R1176_U365 = ~new_P2_R1176_U367 | ~new_P2_U3183 | ~new_P2_R1176_U213;
  assign new_P2_R1176_U366 = ~new_P2_R1176_U215 | ~new_P2_R1176_U217;
  assign new_P2_R1176_U367 = ~new_P2_R1176_U399 | ~new_P2_R1176_U24;
  assign new_P2_R1176_U368 = ~new_P2_R1176_U10 | ~new_P2_R1176_U161;
  assign new_P2_R1176_U369 = ~new_P2_R1176_U231 | ~new_P2_R1176_U5;
  assign new_P2_R1176_U370 = ~new_P2_R1176_U34;
  assign new_P2_R1176_U371 = ~new_P2_R1176_U117 | ~new_P2_R1176_U161;
  assign new_P2_R1176_U372 = ~new_P2_R1176_U34 | ~new_P2_R1176_U240;
  assign new_P2_R1176_U373 = ~new_P2_R1176_U11 | ~new_P2_R1176_U202;
  assign new_P2_R1176_U374 = ~new_P2_R1176_U261 | ~new_P2_R1176_U9;
  assign new_P2_R1176_U375 = ~new_P2_R1176_U377 | ~new_P2_R1176_U376 | ~new_P2_R1176_U311;
  assign new_P2_R1176_U376 = ~new_P2_R1176_U77 | ~new_P2_R1176_U309;
  assign new_P2_R1176_U377 = ~new_P2_U3157 | ~new_P2_R1176_U309;
  assign new_P2_R1176_U378 = ~new_P2_R1176_U62;
  assign new_P2_R1176_U379 = ~new_P2_R1176_U123 | ~new_P2_R1176_U202;
  assign new_P2_R1176_U380 = ~new_P2_R1176_U62 | ~new_P2_R1176_U272;
  assign new_P2_R1176_U381 = ~new_P2_R1176_U131 | ~new_P2_R1176_U375;
  assign new_P2_R1176_U382 = ~new_P2_R1176_U132 | ~new_P2_R1176_U186 | ~new_P2_R1176_U203;
  assign new_P2_R1176_U383 = ~new_P2_R1176_U313 | ~new_P2_R1176_U384 | ~new_P2_R1176_U309;
  assign new_P2_R1176_U384 = ~new_P2_R1176_U212 | ~new_P2_R1176_U209;
  assign new_P2_R1176_U385 = ~new_P2_R1176_U138 | ~new_P2_R1176_U322;
  assign new_P2_R1176_U386 = ~new_P2_U3184 | ~new_P2_R1176_U146;
  assign new_P2_R1176_U387 = ~new_P2_U3456 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U388 = ~new_P2_R1176_U64;
  assign new_P2_R1176_U389 = ~new_P2_R1176_U388 | ~new_P2_U3174;
  assign new_P2_R1176_U390 = ~new_P2_R1176_U64 | ~new_P2_R1176_U33;
  assign new_P2_R1176_U391 = ~new_P2_R1176_U388 | ~new_P2_U3174;
  assign new_P2_R1176_U392 = ~new_P2_R1176_U64 | ~new_P2_R1176_U33;
  assign new_P2_R1176_U393 = ~new_P2_R1176_U392 | ~new_P2_R1176_U391;
  assign new_P2_R1176_U394 = ~new_P2_U3184 | ~new_P2_R1176_U148;
  assign new_P2_R1176_U395 = ~new_P2_U3441 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U396 = ~new_P2_R1176_U70;
  assign new_P2_R1176_U397 = ~new_P2_U3184 | ~new_P2_R1176_U149;
  assign new_P2_R1176_U398 = ~new_P2_U3432 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U399 = ~new_P2_R1176_U68;
  assign new_P2_R1176_U400 = ~new_P2_U3184 | ~new_P2_R1176_U150;
  assign new_P2_R1176_U401 = ~new_P2_U3427 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U402 = ~new_P2_R1176_U69;
  assign new_P2_R1176_U403 = ~new_P2_U3184 | ~new_P2_R1176_U151;
  assign new_P2_R1176_U404 = ~new_P2_U3438 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U405 = ~new_P2_R1176_U67;
  assign new_P2_R1176_U406 = ~new_P2_U3184 | ~new_P2_R1176_U152;
  assign new_P2_R1176_U407 = ~new_P2_U3435 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U408 = ~new_P2_R1176_U66;
  assign new_P2_R1176_U409 = ~new_P2_U3184 | ~new_P2_R1176_U153;
  assign new_P2_R1176_U410 = ~new_P2_U3444 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U411 = ~new_P2_R1176_U71;
  assign new_P2_R1176_U412 = ~new_P2_U3184 | ~new_P2_R1176_U154;
  assign new_P2_R1176_U413 = ~new_P2_U3450 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U414 = ~new_P2_R1176_U72;
  assign new_P2_R1176_U415 = ~new_P2_U3184 | ~new_P2_R1176_U155;
  assign new_P2_R1176_U416 = ~new_P2_U3447 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U417 = ~new_P2_R1176_U73;
  assign new_P2_R1176_U418 = ~new_P2_U3184 | ~new_P2_R1176_U156;
  assign new_P2_R1176_U419 = ~new_P2_U3453 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U420 = ~new_P2_R1176_U65;
  assign new_P2_R1176_U421 = ~new_P2_R1176_U147 | ~new_P2_R1176_U157;
  assign new_P2_R1176_U422 = ~new_P2_R1176_U242 | ~new_P2_R1176_U393;
  assign new_P2_R1176_U423 = ~new_P2_R1176_U420 | ~new_P2_U3175;
  assign new_P2_R1176_U424 = ~new_P2_R1176_U65 | ~new_P2_R1176_U20;
  assign new_P2_R1176_U425 = ~new_P2_R1176_U420 | ~new_P2_U3175;
  assign new_P2_R1176_U426 = ~new_P2_R1176_U65 | ~new_P2_R1176_U20;
  assign new_P2_R1176_U427 = ~new_P2_R1176_U426 | ~new_P2_R1176_U425;
  assign new_P2_R1176_U428 = ~new_P2_R1176_U158 | ~new_P2_R1176_U159;
  assign new_P2_R1176_U429 = ~new_P2_R1176_U239 | ~new_P2_R1176_U427;
  assign new_P2_R1176_U430 = ~new_P2_R1176_U414 | ~new_P2_U3176;
  assign new_P2_R1176_U431 = ~new_P2_R1176_U72 | ~new_P2_R1176_U30;
  assign new_P2_R1176_U432 = ~new_P2_R1176_U417 | ~new_P2_U3177;
  assign new_P2_R1176_U433 = ~new_P2_R1176_U73 | ~new_P2_R1176_U28;
  assign new_P2_R1176_U434 = ~new_P2_R1176_U433 | ~new_P2_R1176_U432;
  assign new_P2_R1176_U435 = ~new_P2_R1176_U353 | ~new_P2_R1176_U35;
  assign new_P2_R1176_U436 = ~new_P2_R1176_U434 | ~new_P2_R1176_U232;
  assign new_P2_R1176_U437 = ~new_P2_R1176_U411 | ~new_P2_U3178;
  assign new_P2_R1176_U438 = ~new_P2_R1176_U71 | ~new_P2_R1176_U31;
  assign new_P2_R1176_U439 = ~new_P2_R1176_U411 | ~new_P2_U3178;
  assign new_P2_R1176_U440 = ~new_P2_R1176_U71 | ~new_P2_R1176_U31;
  assign new_P2_R1176_U441 = ~new_P2_R1176_U440 | ~new_P2_R1176_U439;
  assign new_P2_R1176_U442 = ~new_P2_R1176_U160 | ~new_P2_R1176_U161;
  assign new_P2_R1176_U443 = ~new_P2_R1176_U228 | ~new_P2_R1176_U441;
  assign new_P2_R1176_U444 = ~new_P2_R1176_U396 | ~new_P2_U3179;
  assign new_P2_R1176_U445 = ~new_P2_R1176_U70 | ~new_P2_R1176_U27;
  assign new_P2_R1176_U446 = ~new_P2_R1176_U396 | ~new_P2_U3179;
  assign new_P2_R1176_U447 = ~new_P2_R1176_U70 | ~new_P2_R1176_U27;
  assign new_P2_R1176_U448 = ~new_P2_R1176_U447 | ~new_P2_R1176_U446;
  assign new_P2_R1176_U449 = ~new_P2_R1176_U162 | ~new_P2_R1176_U163;
  assign new_P2_R1176_U450 = ~new_P2_R1176_U226 | ~new_P2_R1176_U448;
  assign new_P2_R1176_U451 = ~new_P2_R1176_U405 | ~new_P2_U3180;
  assign new_P2_R1176_U452 = ~new_P2_R1176_U67 | ~new_P2_R1176_U23;
  assign new_P2_R1176_U453 = ~new_P2_R1176_U408 | ~new_P2_U3181;
  assign new_P2_R1176_U454 = ~new_P2_R1176_U66 | ~new_P2_R1176_U21;
  assign new_P2_R1176_U455 = ~new_P2_R1176_U454 | ~new_P2_R1176_U453;
  assign new_P2_R1176_U456 = ~new_P2_R1176_U354 | ~new_P2_R1176_U36;
  assign new_P2_R1176_U457 = ~new_P2_R1176_U455 | ~new_P2_R1176_U219;
  assign new_P2_R1176_U458 = ~new_P2_U3184 | ~new_P2_R1176_U164;
  assign new_P2_R1176_U459 = ~new_P2_U3950 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U460 = ~new_P2_R1176_U74;
  assign new_P2_R1176_U461 = ~new_P2_U3184 | ~new_P2_R1176_U165;
  assign new_P2_R1176_U462 = ~new_P2_U3951 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U463 = ~new_P2_R1176_U77;
  assign new_P2_R1176_U464 = ~new_P2_U3184 | ~new_P2_R1176_U166;
  assign new_P2_R1176_U465 = ~new_P2_U3459 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U466 = ~new_P2_R1176_U81;
  assign new_P2_R1176_U467 = ~new_P2_U3184 | ~new_P2_R1176_U167;
  assign new_P2_R1176_U468 = ~new_P2_U3462 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U469 = ~new_P2_R1176_U82;
  assign new_P2_R1176_U470 = ~new_P2_U3184 | ~new_P2_R1176_U168;
  assign new_P2_R1176_U471 = ~new_P2_U3468 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U472 = ~new_P2_R1176_U83;
  assign new_P2_R1176_U473 = ~new_P2_U3184 | ~new_P2_R1176_U169;
  assign new_P2_R1176_U474 = ~new_P2_U3465 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U475 = ~new_P2_R1176_U84;
  assign new_P2_R1176_U476 = ~new_P2_U3184 | ~new_P2_R1176_U170;
  assign new_P2_R1176_U477 = ~new_P2_U3471 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U478 = ~new_P2_R1176_U80;
  assign new_P2_R1176_U479 = ~new_P2_U3184 | ~new_P2_R1176_U171;
  assign new_P2_R1176_U480 = ~new_P2_U3474 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U481 = ~new_P2_R1176_U85;
  assign new_P2_R1176_U482 = ~new_P2_U3184 | ~new_P2_R1176_U172;
  assign new_P2_R1176_U483 = ~new_P2_U3480 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U484 = ~new_P2_R1176_U79;
  assign new_P2_R1176_U485 = ~new_P2_U3184 | ~new_P2_R1176_U173;
  assign new_P2_R1176_U486 = ~new_P2_U3477 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U487 = ~new_P2_R1176_U78;
  assign new_P2_R1176_U488 = ~new_P2_U3184 | ~new_P2_R1176_U174;
  assign new_P2_R1176_U489 = ~new_P2_U3483 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U490 = ~new_P2_R1176_U86;
  assign new_P2_R1176_U491 = ~new_P2_U3184 | ~new_P2_R1176_U175;
  assign new_P2_R1176_U492 = ~new_P2_U3956 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U493 = ~new_P2_R1176_U88;
  assign new_P2_R1176_U494 = ~new_P2_U3184 | ~new_P2_R1176_U176;
  assign new_P2_R1176_U495 = ~new_P2_U3957 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U496 = ~new_P2_R1176_U89;
  assign new_P2_R1176_U497 = ~new_P2_U3184 | ~new_P2_R1176_U177;
  assign new_P2_R1176_U498 = ~new_P2_U3485 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U499 = ~new_P2_R1176_U87;
  assign new_P2_R1176_U500 = ~new_P2_U3184 | ~new_P2_R1176_U178;
  assign new_P2_R1176_U501 = ~new_P2_U3955 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U502 = ~new_P2_R1176_U90;
  assign new_P2_R1176_U503 = ~new_P2_U3184 | ~new_P2_R1176_U179;
  assign new_P2_R1176_U504 = ~new_P2_U3954 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U505 = ~new_P2_R1176_U91;
  assign new_P2_R1176_U506 = ~new_P2_U3184 | ~new_P2_R1176_U180;
  assign new_P2_R1176_U507 = ~new_P2_U3952 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U508 = ~new_P2_R1176_U75;
  assign new_P2_R1176_U509 = ~new_P2_U3184 | ~new_P2_R1176_U181;
  assign new_P2_R1176_U510 = ~new_P2_U3953 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U511 = ~new_P2_R1176_U76;
  assign new_P2_R1176_U512 = ~new_P2_U3184 | ~new_P2_R1176_U182;
  assign new_P2_R1176_U513 = ~new_P2_U3949 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U514 = ~new_P2_R1176_U134;
  assign new_P2_R1176_U515 = ~new_P2_U3155 | ~new_P2_R1176_U514;
  assign new_P2_R1176_U516 = ~new_P2_R1176_U134 | ~new_P2_R1176_U183;
  assign new_P2_R1176_U517 = ~new_P2_R1176_U92;
  assign new_P2_R1176_U518 = ~new_P2_R1176_U517 | ~new_P2_R1176_U364 | ~new_P2_R1176_U317;
  assign new_P2_R1176_U519 = ~new_P2_R1176_U92 | ~new_P2_R1176_U133 | ~new_P2_R1176_U382;
  assign new_P2_R1176_U520 = ~new_P2_R1176_U460 | ~new_P2_U3156;
  assign new_P2_R1176_U521 = ~new_P2_R1176_U74 | ~new_P2_R1176_U37;
  assign new_P2_R1176_U522 = ~new_P2_R1176_U460 | ~new_P2_U3156;
  assign new_P2_R1176_U523 = ~new_P2_R1176_U74 | ~new_P2_R1176_U37;
  assign new_P2_R1176_U524 = ~new_P2_R1176_U523 | ~new_P2_R1176_U522;
  assign new_P2_R1176_U525 = ~new_P2_R1176_U184 | ~new_P2_R1176_U185;
  assign new_P2_R1176_U526 = ~new_P2_R1176_U316 | ~new_P2_R1176_U524;
  assign new_P2_R1176_U527 = ~new_P2_R1176_U463 | ~new_P2_U3157;
  assign new_P2_R1176_U528 = ~new_P2_R1176_U77 | ~new_P2_R1176_U40;
  assign new_P2_R1176_U529 = ~new_P2_R1176_U508 | ~new_P2_U3158;
  assign new_P2_R1176_U530 = ~new_P2_R1176_U75 | ~new_P2_R1176_U38;
  assign new_P2_R1176_U531 = ~new_P2_R1176_U530 | ~new_P2_R1176_U529;
  assign new_P2_R1176_U532 = ~new_P2_R1176_U355 | ~new_P2_R1176_U59;
  assign new_P2_R1176_U533 = ~new_P2_R1176_U531 | ~new_P2_R1176_U322;
  assign new_P2_R1176_U534 = ~new_P2_R1176_U511 | ~new_P2_U3159;
  assign new_P2_R1176_U535 = ~new_P2_R1176_U76 | ~new_P2_R1176_U39;
  assign new_P2_R1176_U536 = ~new_P2_R1176_U535 | ~new_P2_R1176_U534;
  assign new_P2_R1176_U537 = ~new_P2_R1176_U356 | ~new_P2_R1176_U186;
  assign new_P2_R1176_U538 = ~new_P2_R1176_U308 | ~new_P2_R1176_U536;
  assign new_P2_R1176_U539 = ~new_P2_R1176_U505 | ~new_P2_U3160;
  assign new_P2_R1176_U540 = ~new_P2_R1176_U91 | ~new_P2_R1176_U58;
  assign new_P2_R1176_U541 = ~new_P2_R1176_U505 | ~new_P2_U3160;
  assign new_P2_R1176_U542 = ~new_P2_R1176_U91 | ~new_P2_R1176_U58;
  assign new_P2_R1176_U543 = ~new_P2_R1176_U542 | ~new_P2_R1176_U541;
  assign new_P2_R1176_U544 = ~new_P2_R1176_U187 | ~new_P2_R1176_U188;
  assign new_P2_R1176_U545 = ~new_P2_R1176_U304 | ~new_P2_R1176_U543;
  assign new_P2_R1176_U546 = ~new_P2_R1176_U502 | ~new_P2_U3161;
  assign new_P2_R1176_U547 = ~new_P2_R1176_U90 | ~new_P2_R1176_U57;
  assign new_P2_R1176_U548 = ~new_P2_R1176_U502 | ~new_P2_U3161;
  assign new_P2_R1176_U549 = ~new_P2_R1176_U90 | ~new_P2_R1176_U57;
  assign new_P2_R1176_U550 = ~new_P2_R1176_U549 | ~new_P2_R1176_U548;
  assign new_P2_R1176_U551 = ~new_P2_R1176_U189 | ~new_P2_R1176_U190;
  assign new_P2_R1176_U552 = ~new_P2_R1176_U300 | ~new_P2_R1176_U550;
  assign new_P2_R1176_U553 = ~new_P2_R1176_U493 | ~new_P2_U3162;
  assign new_P2_R1176_U554 = ~new_P2_R1176_U88 | ~new_P2_R1176_U56;
  assign new_P2_R1176_U555 = ~new_P2_R1176_U496 | ~new_P2_U3163;
  assign new_P2_R1176_U556 = ~new_P2_R1176_U89 | ~new_P2_R1176_U53;
  assign new_P2_R1176_U557 = ~new_P2_R1176_U556 | ~new_P2_R1176_U555;
  assign new_P2_R1176_U558 = ~new_P2_R1176_U357 | ~new_P2_R1176_U60;
  assign new_P2_R1176_U559 = ~new_P2_R1176_U557 | ~new_P2_R1176_U329;
  assign new_P2_R1176_U560 = ~new_P2_R1176_U399 | ~new_P2_U3182;
  assign new_P2_R1176_U561 = ~new_P2_R1176_U68 | ~new_P2_R1176_U24;
  assign new_P2_R1176_U562 = ~new_P2_R1176_U399 | ~new_P2_U3182;
  assign new_P2_R1176_U563 = ~new_P2_R1176_U68 | ~new_P2_R1176_U24;
  assign new_P2_R1176_U564 = ~new_P2_R1176_U563 | ~new_P2_R1176_U562;
  assign new_P2_R1176_U565 = ~new_P2_R1176_U191 | ~new_P2_R1176_U192;
  assign new_P2_R1176_U566 = ~new_P2_R1176_U216 | ~new_P2_R1176_U564;
  assign new_P2_R1176_U567 = ~new_P2_R1176_U499 | ~new_P2_U3164;
  assign new_P2_R1176_U568 = ~new_P2_R1176_U87 | ~new_P2_R1176_U54;
  assign new_P2_R1176_U569 = ~new_P2_R1176_U568 | ~new_P2_R1176_U567;
  assign new_P2_R1176_U570 = ~new_P2_R1176_U358 | ~new_P2_R1176_U193;
  assign new_P2_R1176_U571 = ~new_P2_R1176_U290 | ~new_P2_R1176_U569;
  assign new_P2_R1176_U572 = ~new_P2_R1176_U490 | ~new_P2_U3165;
  assign new_P2_R1176_U573 = ~new_P2_R1176_U86 | ~new_P2_R1176_U52;
  assign new_P2_R1176_U574 = ~new_P2_R1176_U490 | ~new_P2_U3165;
  assign new_P2_R1176_U575 = ~new_P2_R1176_U86 | ~new_P2_R1176_U52;
  assign new_P2_R1176_U576 = ~new_P2_R1176_U575 | ~new_P2_R1176_U574;
  assign new_P2_R1176_U577 = ~new_P2_R1176_U194 | ~new_P2_R1176_U195;
  assign new_P2_R1176_U578 = ~new_P2_R1176_U286 | ~new_P2_R1176_U576;
  assign new_P2_R1176_U579 = ~new_P2_R1176_U484 | ~new_P2_U3166;
  assign new_P2_R1176_U580 = ~new_P2_R1176_U79 | ~new_P2_R1176_U43;
  assign new_P2_R1176_U581 = ~new_P2_R1176_U487 | ~new_P2_U3167;
  assign new_P2_R1176_U582 = ~new_P2_R1176_U78 | ~new_P2_R1176_U41;
  assign new_P2_R1176_U583 = ~new_P2_R1176_U582 | ~new_P2_R1176_U581;
  assign new_P2_R1176_U584 = ~new_P2_R1176_U359 | ~new_P2_R1176_U61;
  assign new_P2_R1176_U585 = ~new_P2_R1176_U583 | ~new_P2_R1176_U278;
  assign new_P2_R1176_U586 = ~new_P2_R1176_U481 | ~new_P2_U3168;
  assign new_P2_R1176_U587 = ~new_P2_R1176_U85 | ~new_P2_R1176_U51;
  assign new_P2_R1176_U588 = ~new_P2_R1176_U481 | ~new_P2_U3168;
  assign new_P2_R1176_U589 = ~new_P2_R1176_U85 | ~new_P2_R1176_U51;
  assign new_P2_R1176_U590 = ~new_P2_R1176_U589 | ~new_P2_R1176_U588;
  assign new_P2_R1176_U591 = ~new_P2_R1176_U196 | ~new_P2_R1176_U197;
  assign new_P2_R1176_U592 = ~new_P2_R1176_U274 | ~new_P2_R1176_U590;
  assign new_P2_R1176_U593 = ~new_P2_R1176_U478 | ~new_P2_U3169;
  assign new_P2_R1176_U594 = ~new_P2_R1176_U80 | ~new_P2_R1176_U44;
  assign new_P2_R1176_U595 = ~new_P2_R1176_U478 | ~new_P2_U3169;
  assign new_P2_R1176_U596 = ~new_P2_R1176_U80 | ~new_P2_R1176_U44;
  assign new_P2_R1176_U597 = ~new_P2_R1176_U596 | ~new_P2_R1176_U595;
  assign new_P2_R1176_U598 = ~new_P2_R1176_U198 | ~new_P2_R1176_U199;
  assign new_P2_R1176_U599 = ~new_P2_R1176_U271 | ~new_P2_R1176_U597;
  assign new_P2_R1176_U600 = ~new_P2_R1176_U472 | ~new_P2_U3170;
  assign new_P2_R1176_U601 = ~new_P2_R1176_U83 | ~new_P2_R1176_U48;
  assign new_P2_R1176_U602 = ~new_P2_R1176_U475 | ~new_P2_U3171;
  assign new_P2_R1176_U603 = ~new_P2_R1176_U84 | ~new_P2_R1176_U45;
  assign new_P2_R1176_U604 = ~new_P2_R1176_U603 | ~new_P2_R1176_U602;
  assign new_P2_R1176_U605 = ~new_P2_R1176_U360 | ~new_P2_R1176_U63;
  assign new_P2_R1176_U606 = ~new_P2_R1176_U604 | ~new_P2_R1176_U345;
  assign new_P2_R1176_U607 = ~new_P2_R1176_U469 | ~new_P2_U3172;
  assign new_P2_R1176_U608 = ~new_P2_R1176_U82 | ~new_P2_R1176_U46;
  assign new_P2_R1176_U609 = ~new_P2_R1176_U608 | ~new_P2_R1176_U607;
  assign new_P2_R1176_U610 = ~new_P2_R1176_U361 | ~new_P2_R1176_U200;
  assign new_P2_R1176_U611 = ~new_P2_R1176_U262 | ~new_P2_R1176_U609;
  assign new_P2_R1176_U612 = ~new_P2_R1176_U466 | ~new_P2_U3173;
  assign new_P2_R1176_U613 = ~new_P2_R1176_U81 | ~new_P2_R1176_U49;
  assign new_P2_R1176_U614 = ~new_P2_R1176_U466 | ~new_P2_U3173;
  assign new_P2_R1176_U615 = ~new_P2_R1176_U81 | ~new_P2_R1176_U49;
  assign new_P2_R1176_U616 = ~new_P2_R1176_U615 | ~new_P2_R1176_U614;
  assign new_P2_R1176_U617 = ~new_P2_R1176_U201 | ~new_P2_R1176_U202;
  assign new_P2_R1176_U618 = ~new_P2_R1176_U258 | ~new_P2_R1176_U616;
  assign new_P2_R1176_U619 = ~new_P2_R1176_U69 | ~new_P2_R1176_U19;
  assign new_P2_R1176_U620 = ~new_P2_R1176_U402 | ~new_P2_U3184;
  assign new_P2_R1176_U621 = ~new_P2_R1176_U145;
  assign new_P2_R1176_U622 = ~new_P2_R1176_U621 | ~new_P2_U3183;
  assign new_P2_R1176_U623 = ~new_P2_R1176_U145 | ~new_P2_R1176_U25;
  assign new_P2_R1131_U4 = new_P2_R1131_U179 & new_P2_R1131_U178;
  assign new_P2_R1131_U5 = new_P2_R1131_U197 & new_P2_R1131_U196;
  assign new_P2_R1131_U6 = new_P2_R1131_U237 & new_P2_R1131_U236;
  assign new_P2_R1131_U7 = new_P2_R1131_U246 & new_P2_R1131_U245;
  assign new_P2_R1131_U8 = new_P2_R1131_U264 & new_P2_R1131_U263;
  assign new_P2_R1131_U9 = new_P2_R1131_U272 & new_P2_R1131_U271;
  assign new_P2_R1131_U10 = new_P2_R1131_U351 & new_P2_R1131_U348;
  assign new_P2_R1131_U11 = new_P2_R1131_U344 & new_P2_R1131_U341;
  assign new_P2_R1131_U12 = new_P2_R1131_U335 & new_P2_R1131_U332;
  assign new_P2_R1131_U13 = new_P2_R1131_U326 & new_P2_R1131_U323;
  assign new_P2_R1131_U14 = new_P2_R1131_U320 & new_P2_R1131_U318;
  assign new_P2_R1131_U15 = new_P2_R1131_U313 & new_P2_R1131_U310;
  assign new_P2_R1131_U16 = new_P2_R1131_U235 & new_P2_R1131_U232;
  assign new_P2_R1131_U17 = new_P2_R1131_U227 & new_P2_R1131_U224;
  assign new_P2_R1131_U18 = new_P2_R1131_U213 & new_P2_R1131_U210;
  assign new_P2_R1131_U19 = ~new_P2_U3447;
  assign new_P2_R1131_U20 = ~new_P2_U3073;
  assign new_P2_R1131_U21 = ~new_P2_U3072;
  assign new_P2_R1131_U22 = ~new_P2_U3073 | ~new_P2_U3447;
  assign new_P2_R1131_U23 = ~new_P2_U3450;
  assign new_P2_R1131_U24 = ~new_P2_U3441;
  assign new_P2_R1131_U25 = ~new_P2_U3062;
  assign new_P2_R1131_U26 = ~new_P2_U3069;
  assign new_P2_R1131_U27 = ~new_P2_U3435;
  assign new_P2_R1131_U28 = ~new_P2_U3070;
  assign new_P2_R1131_U29 = ~new_P2_U3427;
  assign new_P2_R1131_U30 = ~new_P2_U3079;
  assign new_P2_R1131_U31 = ~new_P2_U3079 | ~new_P2_U3427;
  assign new_P2_R1131_U32 = ~new_P2_U3438;
  assign new_P2_R1131_U33 = ~new_P2_U3066;
  assign new_P2_R1131_U34 = ~new_P2_U3062 | ~new_P2_U3441;
  assign new_P2_R1131_U35 = ~new_P2_U3444;
  assign new_P2_R1131_U36 = ~new_P2_U3453;
  assign new_P2_R1131_U37 = ~new_P2_U3086;
  assign new_P2_R1131_U38 = ~new_P2_U3085;
  assign new_P2_R1131_U39 = ~new_P2_U3456;
  assign new_P2_R1131_U40 = ~new_P2_R1131_U61 | ~new_P2_R1131_U205;
  assign new_P2_R1131_U41 = ~new_P2_R1131_U117 | ~new_P2_R1131_U193;
  assign new_P2_R1131_U42 = ~new_P2_R1131_U182 | ~new_P2_R1131_U183;
  assign new_P2_R1131_U43 = ~new_P2_U3432 | ~new_P2_U3080;
  assign new_P2_R1131_U44 = ~new_P2_R1131_U122 | ~new_P2_R1131_U219;
  assign new_P2_R1131_U45 = ~new_P2_R1131_U216 | ~new_P2_R1131_U215;
  assign new_P2_R1131_U46 = ~new_P2_U3950;
  assign new_P2_R1131_U47 = ~new_P2_U3055;
  assign new_P2_R1131_U48 = ~new_P2_U3059;
  assign new_P2_R1131_U49 = ~new_P2_U3951;
  assign new_P2_R1131_U50 = ~new_P2_U3952;
  assign new_P2_R1131_U51 = ~new_P2_U3060;
  assign new_P2_R1131_U52 = ~new_P2_U3953;
  assign new_P2_R1131_U53 = ~new_P2_U3067;
  assign new_P2_R1131_U54 = ~new_P2_U3956;
  assign new_P2_R1131_U55 = ~new_P2_U3077;
  assign new_P2_R1131_U56 = ~new_P2_U3477;
  assign new_P2_R1131_U57 = ~new_P2_U3075;
  assign new_P2_R1131_U58 = ~new_P2_U3071;
  assign new_P2_R1131_U59 = ~new_P2_U3075 | ~new_P2_U3477;
  assign new_P2_R1131_U60 = ~new_P2_U3480;
  assign new_P2_R1131_U61 = ~new_P2_U3086 | ~new_P2_U3453;
  assign new_P2_R1131_U62 = ~new_P2_U3459;
  assign new_P2_R1131_U63 = ~new_P2_U3064;
  assign new_P2_R1131_U64 = ~new_P2_U3465;
  assign new_P2_R1131_U65 = ~new_P2_U3074;
  assign new_P2_R1131_U66 = ~new_P2_U3462;
  assign new_P2_R1131_U67 = ~new_P2_U3065;
  assign new_P2_R1131_U68 = ~new_P2_U3065 | ~new_P2_U3462;
  assign new_P2_R1131_U69 = ~new_P2_U3468;
  assign new_P2_R1131_U70 = ~new_P2_U3082;
  assign new_P2_R1131_U71 = ~new_P2_U3471;
  assign new_P2_R1131_U72 = ~new_P2_U3081;
  assign new_P2_R1131_U73 = ~new_P2_U3474;
  assign new_P2_R1131_U74 = ~new_P2_U3076;
  assign new_P2_R1131_U75 = ~new_P2_U3483;
  assign new_P2_R1131_U76 = ~new_P2_U3084;
  assign new_P2_R1131_U77 = ~new_P2_U3084 | ~new_P2_U3483;
  assign new_P2_R1131_U78 = ~new_P2_U3485;
  assign new_P2_R1131_U79 = ~new_P2_U3083;
  assign new_P2_R1131_U80 = ~new_P2_U3083 | ~new_P2_U3485;
  assign new_P2_R1131_U81 = ~new_P2_U3957;
  assign new_P2_R1131_U82 = ~new_P2_U3955;
  assign new_P2_R1131_U83 = ~new_P2_U3063;
  assign new_P2_R1131_U84 = ~new_P2_U3954;
  assign new_P2_R1131_U85 = ~new_P2_U3068;
  assign new_P2_R1131_U86 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1131_U87 = ~new_P2_U3056;
  assign new_P2_R1131_U88 = ~new_P2_U3949;
  assign new_P2_R1131_U89 = ~new_P2_R1131_U306 | ~new_P2_R1131_U176;
  assign new_P2_R1131_U90 = ~new_P2_U3078;
  assign new_P2_R1131_U91 = ~new_P2_R1131_U77 | ~new_P2_R1131_U315;
  assign new_P2_R1131_U92 = ~new_P2_R1131_U261 | ~new_P2_R1131_U260;
  assign new_P2_R1131_U93 = ~new_P2_R1131_U68 | ~new_P2_R1131_U337;
  assign new_P2_R1131_U94 = ~new_P2_R1131_U457 | ~new_P2_R1131_U456;
  assign new_P2_R1131_U95 = ~new_P2_R1131_U504 | ~new_P2_R1131_U503;
  assign new_P2_R1131_U96 = ~new_P2_R1131_U375 | ~new_P2_R1131_U374;
  assign new_P2_R1131_U97 = ~new_P2_R1131_U380 | ~new_P2_R1131_U379;
  assign new_P2_R1131_U98 = ~new_P2_R1131_U387 | ~new_P2_R1131_U386;
  assign new_P2_R1131_U99 = ~new_P2_R1131_U394 | ~new_P2_R1131_U393;
  assign new_P2_R1131_U100 = ~new_P2_R1131_U399 | ~new_P2_R1131_U398;
  assign new_P2_R1131_U101 = ~new_P2_R1131_U408 | ~new_P2_R1131_U407;
  assign new_P2_R1131_U102 = ~new_P2_R1131_U415 | ~new_P2_R1131_U414;
  assign new_P2_R1131_U103 = ~new_P2_R1131_U422 | ~new_P2_R1131_U421;
  assign new_P2_R1131_U104 = ~new_P2_R1131_U429 | ~new_P2_R1131_U428;
  assign new_P2_R1131_U105 = ~new_P2_R1131_U434 | ~new_P2_R1131_U433;
  assign new_P2_R1131_U106 = ~new_P2_R1131_U441 | ~new_P2_R1131_U440;
  assign new_P2_R1131_U107 = ~new_P2_R1131_U448 | ~new_P2_R1131_U447;
  assign new_P2_R1131_U108 = ~new_P2_R1131_U462 | ~new_P2_R1131_U461;
  assign new_P2_R1131_U109 = ~new_P2_R1131_U467 | ~new_P2_R1131_U466;
  assign new_P2_R1131_U110 = ~new_P2_R1131_U474 | ~new_P2_R1131_U473;
  assign new_P2_R1131_U111 = ~new_P2_R1131_U481 | ~new_P2_R1131_U480;
  assign new_P2_R1131_U112 = ~new_P2_R1131_U488 | ~new_P2_R1131_U487;
  assign new_P2_R1131_U113 = ~new_P2_R1131_U495 | ~new_P2_R1131_U494;
  assign new_P2_R1131_U114 = ~new_P2_R1131_U500 | ~new_P2_R1131_U499;
  assign new_P2_R1131_U115 = new_P2_R1131_U189 & new_P2_R1131_U187;
  assign new_P2_R1131_U116 = new_P2_R1131_U4 & new_P2_R1131_U180;
  assign new_P2_R1131_U117 = new_P2_R1131_U194 & new_P2_R1131_U192;
  assign new_P2_R1131_U118 = new_P2_R1131_U201 & new_P2_R1131_U200;
  assign new_P2_R1131_U119 = new_P2_R1131_U22 & new_P2_R1131_U382 & new_P2_R1131_U381;
  assign new_P2_R1131_U120 = new_P2_R1131_U212 & new_P2_R1131_U5;
  assign new_P2_R1131_U121 = new_P2_R1131_U181 & new_P2_R1131_U180;
  assign new_P2_R1131_U122 = new_P2_R1131_U220 & new_P2_R1131_U218;
  assign new_P2_R1131_U123 = new_P2_R1131_U34 & new_P2_R1131_U389 & new_P2_R1131_U388;
  assign new_P2_R1131_U124 = new_P2_R1131_U226 & new_P2_R1131_U4;
  assign new_P2_R1131_U125 = new_P2_R1131_U234 & new_P2_R1131_U181;
  assign new_P2_R1131_U126 = new_P2_R1131_U204 & new_P2_R1131_U6;
  assign new_P2_R1131_U127 = new_P2_R1131_U239 & new_P2_R1131_U171;
  assign new_P2_R1131_U128 = new_P2_R1131_U250 & new_P2_R1131_U7;
  assign new_P2_R1131_U129 = new_P2_R1131_U248 & new_P2_R1131_U172;
  assign new_P2_R1131_U130 = new_P2_R1131_U268 & new_P2_R1131_U267;
  assign new_P2_R1131_U131 = new_P2_R1131_U9 & new_P2_R1131_U282;
  assign new_P2_R1131_U132 = new_P2_R1131_U285 & new_P2_R1131_U280;
  assign new_P2_R1131_U133 = new_P2_R1131_U301 & new_P2_R1131_U298;
  assign new_P2_R1131_U134 = new_P2_R1131_U368 & new_P2_R1131_U302;
  assign new_P2_R1131_U135 = new_P2_R1131_U160 & new_P2_R1131_U278;
  assign new_P2_R1131_U136 = new_P2_R1131_U80 & new_P2_R1131_U455 & new_P2_R1131_U454;
  assign new_P2_R1131_U137 = new_P2_R1131_U325 & new_P2_R1131_U9;
  assign new_P2_R1131_U138 = new_P2_R1131_U59 & new_P2_R1131_U469 & new_P2_R1131_U468;
  assign new_P2_R1131_U139 = new_P2_R1131_U334 & new_P2_R1131_U8;
  assign new_P2_R1131_U140 = new_P2_R1131_U172 & new_P2_R1131_U490 & new_P2_R1131_U489;
  assign new_P2_R1131_U141 = new_P2_R1131_U343 & new_P2_R1131_U7;
  assign new_P2_R1131_U142 = new_P2_R1131_U171 & new_P2_R1131_U502 & new_P2_R1131_U501;
  assign new_P2_R1131_U143 = new_P2_R1131_U350 & new_P2_R1131_U6;
  assign new_P2_R1131_U144 = ~new_P2_R1131_U118 | ~new_P2_R1131_U202;
  assign new_P2_R1131_U145 = ~new_P2_R1131_U217 | ~new_P2_R1131_U229;
  assign new_P2_R1131_U146 = ~new_P2_U3057;
  assign new_P2_R1131_U147 = ~new_P2_U3960;
  assign new_P2_R1131_U148 = new_P2_R1131_U403 & new_P2_R1131_U402;
  assign new_P2_R1131_U149 = ~new_P2_R1131_U364 | ~new_P2_R1131_U304 | ~new_P2_R1131_U169;
  assign new_P2_R1131_U150 = new_P2_R1131_U410 & new_P2_R1131_U409;
  assign new_P2_R1131_U151 = ~new_P2_R1131_U134 | ~new_P2_R1131_U370 | ~new_P2_R1131_U369;
  assign new_P2_R1131_U152 = new_P2_R1131_U417 & new_P2_R1131_U416;
  assign new_P2_R1131_U153 = ~new_P2_R1131_U86 | ~new_P2_R1131_U365 | ~new_P2_R1131_U299;
  assign new_P2_R1131_U154 = new_P2_R1131_U424 & new_P2_R1131_U423;
  assign new_P2_R1131_U155 = ~new_P2_R1131_U293 | ~new_P2_R1131_U292;
  assign new_P2_R1131_U156 = new_P2_R1131_U436 & new_P2_R1131_U435;
  assign new_P2_R1131_U157 = ~new_P2_R1131_U289 | ~new_P2_R1131_U288;
  assign new_P2_R1131_U158 = new_P2_R1131_U443 & new_P2_R1131_U442;
  assign new_P2_R1131_U159 = ~new_P2_R1131_U132 | ~new_P2_R1131_U284;
  assign new_P2_R1131_U160 = new_P2_R1131_U450 & new_P2_R1131_U449;
  assign new_P2_R1131_U161 = ~new_P2_R1131_U43 | ~new_P2_R1131_U327;
  assign new_P2_R1131_U162 = ~new_P2_R1131_U130 | ~new_P2_R1131_U269;
  assign new_P2_R1131_U163 = new_P2_R1131_U476 & new_P2_R1131_U475;
  assign new_P2_R1131_U164 = ~new_P2_R1131_U257 | ~new_P2_R1131_U256;
  assign new_P2_R1131_U165 = new_P2_R1131_U483 & new_P2_R1131_U482;
  assign new_P2_R1131_U166 = ~new_P2_R1131_U253 | ~new_P2_R1131_U252;
  assign new_P2_R1131_U167 = ~new_P2_R1131_U243 | ~new_P2_R1131_U242;
  assign new_P2_R1131_U168 = ~new_P2_R1131_U367 | ~new_P2_R1131_U366;
  assign new_P2_R1131_U169 = ~new_P2_U3056 | ~new_P2_R1131_U151;
  assign new_P2_R1131_U170 = ~new_P2_R1131_U34;
  assign new_P2_R1131_U171 = ~new_P2_U3456 | ~new_P2_U3085;
  assign new_P2_R1131_U172 = ~new_P2_U3074 | ~new_P2_U3465;
  assign new_P2_R1131_U173 = ~new_P2_U3060 | ~new_P2_U3952;
  assign new_P2_R1131_U174 = ~new_P2_R1131_U68;
  assign new_P2_R1131_U175 = ~new_P2_R1131_U77;
  assign new_P2_R1131_U176 = ~new_P2_U3067 | ~new_P2_U3953;
  assign new_P2_R1131_U177 = ~new_P2_R1131_U61;
  assign new_P2_R1131_U178 = new_P2_U3069 | new_P2_U3444;
  assign new_P2_R1131_U179 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1131_U180 = new_P2_U3438 | new_P2_U3066;
  assign new_P2_R1131_U181 = new_P2_U3435 | new_P2_U3070;
  assign new_P2_R1131_U182 = ~new_P2_R1131_U31;
  assign new_P2_R1131_U183 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1131_U184 = ~new_P2_R1131_U42;
  assign new_P2_R1131_U185 = ~new_P2_R1131_U43;
  assign new_P2_R1131_U186 = ~new_P2_R1131_U42 | ~new_P2_R1131_U43;
  assign new_P2_R1131_U187 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1131_U188 = ~new_P2_R1131_U186 | ~new_P2_R1131_U181;
  assign new_P2_R1131_U189 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1131_U190 = ~new_P2_R1131_U115 | ~new_P2_R1131_U188;
  assign new_P2_R1131_U191 = ~new_P2_R1131_U35 | ~new_P2_R1131_U34;
  assign new_P2_R1131_U192 = ~new_P2_U3069 | ~new_P2_R1131_U191;
  assign new_P2_R1131_U193 = ~new_P2_R1131_U116 | ~new_P2_R1131_U190;
  assign new_P2_R1131_U194 = ~new_P2_U3444 | ~new_P2_R1131_U170;
  assign new_P2_R1131_U195 = ~new_P2_R1131_U41;
  assign new_P2_R1131_U196 = new_P2_U3072 | new_P2_U3450;
  assign new_P2_R1131_U197 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1131_U198 = ~new_P2_R1131_U22;
  assign new_P2_R1131_U199 = ~new_P2_R1131_U23 | ~new_P2_R1131_U22;
  assign new_P2_R1131_U200 = ~new_P2_U3072 | ~new_P2_R1131_U199;
  assign new_P2_R1131_U201 = ~new_P2_U3450 | ~new_P2_R1131_U198;
  assign new_P2_R1131_U202 = ~new_P2_R1131_U5 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U203 = ~new_P2_R1131_U144;
  assign new_P2_R1131_U204 = new_P2_U3453 | new_P2_U3086;
  assign new_P2_R1131_U205 = ~new_P2_R1131_U204 | ~new_P2_R1131_U144;
  assign new_P2_R1131_U206 = ~new_P2_R1131_U40;
  assign new_P2_R1131_U207 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1131_U208 = new_P2_U3447 | new_P2_U3073;
  assign new_P2_R1131_U209 = ~new_P2_R1131_U208 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U210 = ~new_P2_R1131_U119 | ~new_P2_R1131_U209;
  assign new_P2_R1131_U211 = ~new_P2_R1131_U195 | ~new_P2_R1131_U22;
  assign new_P2_R1131_U212 = ~new_P2_U3450 | ~new_P2_U3072;
  assign new_P2_R1131_U213 = ~new_P2_R1131_U120 | ~new_P2_R1131_U211;
  assign new_P2_R1131_U214 = new_P2_U3073 | new_P2_U3447;
  assign new_P2_R1131_U215 = ~new_P2_R1131_U185 | ~new_P2_R1131_U181;
  assign new_P2_R1131_U216 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1131_U217 = ~new_P2_R1131_U45;
  assign new_P2_R1131_U218 = ~new_P2_R1131_U121 | ~new_P2_R1131_U184;
  assign new_P2_R1131_U219 = ~new_P2_R1131_U45 | ~new_P2_R1131_U180;
  assign new_P2_R1131_U220 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1131_U221 = ~new_P2_R1131_U44;
  assign new_P2_R1131_U222 = new_P2_U3441 | new_P2_U3062;
  assign new_P2_R1131_U223 = ~new_P2_R1131_U222 | ~new_P2_R1131_U44;
  assign new_P2_R1131_U224 = ~new_P2_R1131_U123 | ~new_P2_R1131_U223;
  assign new_P2_R1131_U225 = ~new_P2_R1131_U221 | ~new_P2_R1131_U34;
  assign new_P2_R1131_U226 = ~new_P2_U3444 | ~new_P2_U3069;
  assign new_P2_R1131_U227 = ~new_P2_R1131_U124 | ~new_P2_R1131_U225;
  assign new_P2_R1131_U228 = new_P2_U3062 | new_P2_U3441;
  assign new_P2_R1131_U229 = ~new_P2_R1131_U184 | ~new_P2_R1131_U181;
  assign new_P2_R1131_U230 = ~new_P2_R1131_U145;
  assign new_P2_R1131_U231 = ~new_P2_U3066 | ~new_P2_U3438;
  assign new_P2_R1131_U232 = ~new_P2_R1131_U42 | ~new_P2_R1131_U43 | ~new_P2_R1131_U401 | ~new_P2_R1131_U400;
  assign new_P2_R1131_U233 = ~new_P2_R1131_U43 | ~new_P2_R1131_U42;
  assign new_P2_R1131_U234 = ~new_P2_U3070 | ~new_P2_U3435;
  assign new_P2_R1131_U235 = ~new_P2_R1131_U125 | ~new_P2_R1131_U233;
  assign new_P2_R1131_U236 = new_P2_U3085 | new_P2_U3456;
  assign new_P2_R1131_U237 = new_P2_U3064 | new_P2_U3459;
  assign new_P2_R1131_U238 = ~new_P2_R1131_U177 | ~new_P2_R1131_U6;
  assign new_P2_R1131_U239 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1131_U240 = ~new_P2_R1131_U127 | ~new_P2_R1131_U238;
  assign new_P2_R1131_U241 = new_P2_U3459 | new_P2_U3064;
  assign new_P2_R1131_U242 = ~new_P2_R1131_U126 | ~new_P2_R1131_U144;
  assign new_P2_R1131_U243 = ~new_P2_R1131_U241 | ~new_P2_R1131_U240;
  assign new_P2_R1131_U244 = ~new_P2_R1131_U167;
  assign new_P2_R1131_U245 = new_P2_U3082 | new_P2_U3468;
  assign new_P2_R1131_U246 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1131_U247 = ~new_P2_R1131_U174 | ~new_P2_R1131_U7;
  assign new_P2_R1131_U248 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1131_U249 = ~new_P2_R1131_U129 | ~new_P2_R1131_U247;
  assign new_P2_R1131_U250 = new_P2_U3462 | new_P2_U3065;
  assign new_P2_R1131_U251 = new_P2_U3468 | new_P2_U3082;
  assign new_P2_R1131_U252 = ~new_P2_R1131_U128 | ~new_P2_R1131_U167;
  assign new_P2_R1131_U253 = ~new_P2_R1131_U251 | ~new_P2_R1131_U249;
  assign new_P2_R1131_U254 = ~new_P2_R1131_U166;
  assign new_P2_R1131_U255 = new_P2_U3471 | new_P2_U3081;
  assign new_P2_R1131_U256 = ~new_P2_R1131_U255 | ~new_P2_R1131_U166;
  assign new_P2_R1131_U257 = ~new_P2_U3081 | ~new_P2_U3471;
  assign new_P2_R1131_U258 = ~new_P2_R1131_U164;
  assign new_P2_R1131_U259 = new_P2_U3474 | new_P2_U3076;
  assign new_P2_R1131_U260 = ~new_P2_R1131_U259 | ~new_P2_R1131_U164;
  assign new_P2_R1131_U261 = ~new_P2_U3076 | ~new_P2_U3474;
  assign new_P2_R1131_U262 = ~new_P2_R1131_U92;
  assign new_P2_R1131_U263 = new_P2_U3071 | new_P2_U3480;
  assign new_P2_R1131_U264 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1131_U265 = ~new_P2_R1131_U59;
  assign new_P2_R1131_U266 = ~new_P2_R1131_U60 | ~new_P2_R1131_U59;
  assign new_P2_R1131_U267 = ~new_P2_U3071 | ~new_P2_R1131_U266;
  assign new_P2_R1131_U268 = ~new_P2_U3480 | ~new_P2_R1131_U265;
  assign new_P2_R1131_U269 = ~new_P2_R1131_U8 | ~new_P2_R1131_U92;
  assign new_P2_R1131_U270 = ~new_P2_R1131_U162;
  assign new_P2_R1131_U271 = new_P2_U3078 | new_P2_U3957;
  assign new_P2_R1131_U272 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1131_U273 = new_P2_U3077 | new_P2_U3956;
  assign new_P2_R1131_U274 = ~new_P2_R1131_U80;
  assign new_P2_R1131_U275 = ~new_P2_U3957 | ~new_P2_R1131_U274;
  assign new_P2_R1131_U276 = ~new_P2_R1131_U275 | ~new_P2_R1131_U90;
  assign new_P2_R1131_U277 = ~new_P2_R1131_U80 | ~new_P2_R1131_U81;
  assign new_P2_R1131_U278 = ~new_P2_R1131_U277 | ~new_P2_R1131_U276;
  assign new_P2_R1131_U279 = ~new_P2_R1131_U175 | ~new_P2_R1131_U9;
  assign new_P2_R1131_U280 = ~new_P2_U3077 | ~new_P2_U3956;
  assign new_P2_R1131_U281 = ~new_P2_R1131_U278 | ~new_P2_R1131_U279;
  assign new_P2_R1131_U282 = new_P2_U3483 | new_P2_U3084;
  assign new_P2_R1131_U283 = new_P2_U3956 | new_P2_U3077;
  assign new_P2_R1131_U284 = ~new_P2_R1131_U131 | ~new_P2_R1131_U273 | ~new_P2_R1131_U162;
  assign new_P2_R1131_U285 = ~new_P2_R1131_U283 | ~new_P2_R1131_U281;
  assign new_P2_R1131_U286 = ~new_P2_R1131_U159;
  assign new_P2_R1131_U287 = new_P2_U3955 | new_P2_U3063;
  assign new_P2_R1131_U288 = ~new_P2_R1131_U287 | ~new_P2_R1131_U159;
  assign new_P2_R1131_U289 = ~new_P2_U3063 | ~new_P2_U3955;
  assign new_P2_R1131_U290 = ~new_P2_R1131_U157;
  assign new_P2_R1131_U291 = new_P2_U3954 | new_P2_U3068;
  assign new_P2_R1131_U292 = ~new_P2_R1131_U291 | ~new_P2_R1131_U157;
  assign new_P2_R1131_U293 = ~new_P2_U3068 | ~new_P2_U3954;
  assign new_P2_R1131_U294 = ~new_P2_R1131_U155;
  assign new_P2_R1131_U295 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1131_U296 = ~new_P2_R1131_U176 | ~new_P2_R1131_U173;
  assign new_P2_R1131_U297 = ~new_P2_R1131_U86;
  assign new_P2_R1131_U298 = new_P2_U3953 | new_P2_U3067;
  assign new_P2_R1131_U299 = ~new_P2_R1131_U168 | ~new_P2_R1131_U155 | ~new_P2_R1131_U298;
  assign new_P2_R1131_U300 = ~new_P2_R1131_U153;
  assign new_P2_R1131_U301 = new_P2_U3950 | new_P2_U3055;
  assign new_P2_R1131_U302 = ~new_P2_U3055 | ~new_P2_U3950;
  assign new_P2_R1131_U303 = ~new_P2_R1131_U151;
  assign new_P2_R1131_U304 = ~new_P2_U3949 | ~new_P2_R1131_U151;
  assign new_P2_R1131_U305 = ~new_P2_R1131_U149;
  assign new_P2_R1131_U306 = ~new_P2_R1131_U298 | ~new_P2_R1131_U155;
  assign new_P2_R1131_U307 = ~new_P2_R1131_U89;
  assign new_P2_R1131_U308 = new_P2_U3952 | new_P2_U3060;
  assign new_P2_R1131_U309 = ~new_P2_R1131_U308 | ~new_P2_R1131_U89;
  assign new_P2_R1131_U310 = ~new_P2_R1131_U154 | ~new_P2_R1131_U309 | ~new_P2_R1131_U173;
  assign new_P2_R1131_U311 = ~new_P2_R1131_U307 | ~new_P2_R1131_U173;
  assign new_P2_R1131_U312 = ~new_P2_U3951 | ~new_P2_U3059;
  assign new_P2_R1131_U313 = ~new_P2_R1131_U168 | ~new_P2_R1131_U311 | ~new_P2_R1131_U312;
  assign new_P2_R1131_U314 = new_P2_U3060 | new_P2_U3952;
  assign new_P2_R1131_U315 = ~new_P2_R1131_U282 | ~new_P2_R1131_U162;
  assign new_P2_R1131_U316 = ~new_P2_R1131_U91;
  assign new_P2_R1131_U317 = ~new_P2_R1131_U9 | ~new_P2_R1131_U91;
  assign new_P2_R1131_U318 = ~new_P2_R1131_U135 | ~new_P2_R1131_U317;
  assign new_P2_R1131_U319 = ~new_P2_R1131_U317 | ~new_P2_R1131_U278;
  assign new_P2_R1131_U320 = ~new_P2_R1131_U453 | ~new_P2_R1131_U319;
  assign new_P2_R1131_U321 = new_P2_U3485 | new_P2_U3083;
  assign new_P2_R1131_U322 = ~new_P2_R1131_U321 | ~new_P2_R1131_U91;
  assign new_P2_R1131_U323 = ~new_P2_R1131_U136 | ~new_P2_R1131_U322;
  assign new_P2_R1131_U324 = ~new_P2_R1131_U316 | ~new_P2_R1131_U80;
  assign new_P2_R1131_U325 = ~new_P2_U3078 | ~new_P2_U3957;
  assign new_P2_R1131_U326 = ~new_P2_R1131_U137 | ~new_P2_R1131_U324;
  assign new_P2_R1131_U327 = new_P2_U3432 | new_P2_U3080;
  assign new_P2_R1131_U328 = ~new_P2_R1131_U161;
  assign new_P2_R1131_U329 = new_P2_U3083 | new_P2_U3485;
  assign new_P2_R1131_U330 = new_P2_U3477 | new_P2_U3075;
  assign new_P2_R1131_U331 = ~new_P2_R1131_U330 | ~new_P2_R1131_U92;
  assign new_P2_R1131_U332 = ~new_P2_R1131_U138 | ~new_P2_R1131_U331;
  assign new_P2_R1131_U333 = ~new_P2_R1131_U262 | ~new_P2_R1131_U59;
  assign new_P2_R1131_U334 = ~new_P2_U3480 | ~new_P2_U3071;
  assign new_P2_R1131_U335 = ~new_P2_R1131_U139 | ~new_P2_R1131_U333;
  assign new_P2_R1131_U336 = new_P2_U3075 | new_P2_U3477;
  assign new_P2_R1131_U337 = ~new_P2_R1131_U250 | ~new_P2_R1131_U167;
  assign new_P2_R1131_U338 = ~new_P2_R1131_U93;
  assign new_P2_R1131_U339 = new_P2_U3465 | new_P2_U3074;
  assign new_P2_R1131_U340 = ~new_P2_R1131_U339 | ~new_P2_R1131_U93;
  assign new_P2_R1131_U341 = ~new_P2_R1131_U140 | ~new_P2_R1131_U340;
  assign new_P2_R1131_U342 = ~new_P2_R1131_U338 | ~new_P2_R1131_U172;
  assign new_P2_R1131_U343 = ~new_P2_U3082 | ~new_P2_U3468;
  assign new_P2_R1131_U344 = ~new_P2_R1131_U141 | ~new_P2_R1131_U342;
  assign new_P2_R1131_U345 = new_P2_U3074 | new_P2_U3465;
  assign new_P2_R1131_U346 = new_P2_U3456 | new_P2_U3085;
  assign new_P2_R1131_U347 = ~new_P2_R1131_U346 | ~new_P2_R1131_U40;
  assign new_P2_R1131_U348 = ~new_P2_R1131_U142 | ~new_P2_R1131_U347;
  assign new_P2_R1131_U349 = ~new_P2_R1131_U206 | ~new_P2_R1131_U171;
  assign new_P2_R1131_U350 = ~new_P2_U3064 | ~new_P2_U3459;
  assign new_P2_R1131_U351 = ~new_P2_R1131_U143 | ~new_P2_R1131_U349;
  assign new_P2_R1131_U352 = ~new_P2_R1131_U207 | ~new_P2_R1131_U171;
  assign new_P2_R1131_U353 = ~new_P2_R1131_U204 | ~new_P2_R1131_U61;
  assign new_P2_R1131_U354 = ~new_P2_R1131_U214 | ~new_P2_R1131_U22;
  assign new_P2_R1131_U355 = ~new_P2_R1131_U228 | ~new_P2_R1131_U34;
  assign new_P2_R1131_U356 = ~new_P2_R1131_U231 | ~new_P2_R1131_U180;
  assign new_P2_R1131_U357 = ~new_P2_R1131_U314 | ~new_P2_R1131_U173;
  assign new_P2_R1131_U358 = ~new_P2_R1131_U298 | ~new_P2_R1131_U176;
  assign new_P2_R1131_U359 = ~new_P2_R1131_U329 | ~new_P2_R1131_U80;
  assign new_P2_R1131_U360 = ~new_P2_R1131_U282 | ~new_P2_R1131_U77;
  assign new_P2_R1131_U361 = ~new_P2_R1131_U336 | ~new_P2_R1131_U59;
  assign new_P2_R1131_U362 = ~new_P2_R1131_U345 | ~new_P2_R1131_U172;
  assign new_P2_R1131_U363 = ~new_P2_R1131_U250 | ~new_P2_R1131_U68;
  assign new_P2_R1131_U364 = ~new_P2_U3949 | ~new_P2_U3056;
  assign new_P2_R1131_U365 = ~new_P2_R1131_U296 | ~new_P2_R1131_U168;
  assign new_P2_R1131_U366 = ~new_P2_U3059 | ~new_P2_R1131_U295;
  assign new_P2_R1131_U367 = ~new_P2_U3951 | ~new_P2_R1131_U295;
  assign new_P2_R1131_U368 = ~new_P2_R1131_U301 | ~new_P2_R1131_U296 | ~new_P2_R1131_U168;
  assign new_P2_R1131_U369 = ~new_P2_R1131_U133 | ~new_P2_R1131_U155 | ~new_P2_R1131_U168;
  assign new_P2_R1131_U370 = ~new_P2_R1131_U297 | ~new_P2_R1131_U301;
  assign new_P2_R1131_U371 = ~new_P2_U3085 | ~new_P2_R1131_U39;
  assign new_P2_R1131_U372 = ~new_P2_U3456 | ~new_P2_R1131_U38;
  assign new_P2_R1131_U373 = ~new_P2_R1131_U372 | ~new_P2_R1131_U371;
  assign new_P2_R1131_U374 = ~new_P2_R1131_U352 | ~new_P2_R1131_U40;
  assign new_P2_R1131_U375 = ~new_P2_R1131_U373 | ~new_P2_R1131_U206;
  assign new_P2_R1131_U376 = ~new_P2_U3086 | ~new_P2_R1131_U36;
  assign new_P2_R1131_U377 = ~new_P2_U3453 | ~new_P2_R1131_U37;
  assign new_P2_R1131_U378 = ~new_P2_R1131_U377 | ~new_P2_R1131_U376;
  assign new_P2_R1131_U379 = ~new_P2_R1131_U353 | ~new_P2_R1131_U144;
  assign new_P2_R1131_U380 = ~new_P2_R1131_U203 | ~new_P2_R1131_U378;
  assign new_P2_R1131_U381 = ~new_P2_U3072 | ~new_P2_R1131_U23;
  assign new_P2_R1131_U382 = ~new_P2_U3450 | ~new_P2_R1131_U21;
  assign new_P2_R1131_U383 = ~new_P2_U3073 | ~new_P2_R1131_U19;
  assign new_P2_R1131_U384 = ~new_P2_U3447 | ~new_P2_R1131_U20;
  assign new_P2_R1131_U385 = ~new_P2_R1131_U384 | ~new_P2_R1131_U383;
  assign new_P2_R1131_U386 = ~new_P2_R1131_U354 | ~new_P2_R1131_U41;
  assign new_P2_R1131_U387 = ~new_P2_R1131_U385 | ~new_P2_R1131_U195;
  assign new_P2_R1131_U388 = ~new_P2_U3069 | ~new_P2_R1131_U35;
  assign new_P2_R1131_U389 = ~new_P2_U3444 | ~new_P2_R1131_U26;
  assign new_P2_R1131_U390 = ~new_P2_U3062 | ~new_P2_R1131_U24;
  assign new_P2_R1131_U391 = ~new_P2_U3441 | ~new_P2_R1131_U25;
  assign new_P2_R1131_U392 = ~new_P2_R1131_U391 | ~new_P2_R1131_U390;
  assign new_P2_R1131_U393 = ~new_P2_R1131_U355 | ~new_P2_R1131_U44;
  assign new_P2_R1131_U394 = ~new_P2_R1131_U392 | ~new_P2_R1131_U221;
  assign new_P2_R1131_U395 = ~new_P2_U3066 | ~new_P2_R1131_U32;
  assign new_P2_R1131_U396 = ~new_P2_U3438 | ~new_P2_R1131_U33;
  assign new_P2_R1131_U397 = ~new_P2_R1131_U396 | ~new_P2_R1131_U395;
  assign new_P2_R1131_U398 = ~new_P2_R1131_U356 | ~new_P2_R1131_U145;
  assign new_P2_R1131_U399 = ~new_P2_R1131_U230 | ~new_P2_R1131_U397;
  assign new_P2_R1131_U400 = ~new_P2_U3070 | ~new_P2_R1131_U27;
  assign new_P2_R1131_U401 = ~new_P2_U3435 | ~new_P2_R1131_U28;
  assign new_P2_R1131_U402 = ~new_P2_U3057 | ~new_P2_R1131_U147;
  assign new_P2_R1131_U403 = ~new_P2_U3960 | ~new_P2_R1131_U146;
  assign new_P2_R1131_U404 = ~new_P2_U3057 | ~new_P2_R1131_U147;
  assign new_P2_R1131_U405 = ~new_P2_U3960 | ~new_P2_R1131_U146;
  assign new_P2_R1131_U406 = ~new_P2_R1131_U405 | ~new_P2_R1131_U404;
  assign new_P2_R1131_U407 = ~new_P2_R1131_U148 | ~new_P2_R1131_U149;
  assign new_P2_R1131_U408 = ~new_P2_R1131_U305 | ~new_P2_R1131_U406;
  assign new_P2_R1131_U409 = ~new_P2_U3056 | ~new_P2_R1131_U88;
  assign new_P2_R1131_U410 = ~new_P2_U3949 | ~new_P2_R1131_U87;
  assign new_P2_R1131_U411 = ~new_P2_U3056 | ~new_P2_R1131_U88;
  assign new_P2_R1131_U412 = ~new_P2_U3949 | ~new_P2_R1131_U87;
  assign new_P2_R1131_U413 = ~new_P2_R1131_U412 | ~new_P2_R1131_U411;
  assign new_P2_R1131_U414 = ~new_P2_R1131_U150 | ~new_P2_R1131_U151;
  assign new_P2_R1131_U415 = ~new_P2_R1131_U303 | ~new_P2_R1131_U413;
  assign new_P2_R1131_U416 = ~new_P2_U3055 | ~new_P2_R1131_U46;
  assign new_P2_R1131_U417 = ~new_P2_U3950 | ~new_P2_R1131_U47;
  assign new_P2_R1131_U418 = ~new_P2_U3055 | ~new_P2_R1131_U46;
  assign new_P2_R1131_U419 = ~new_P2_U3950 | ~new_P2_R1131_U47;
  assign new_P2_R1131_U420 = ~new_P2_R1131_U419 | ~new_P2_R1131_U418;
  assign new_P2_R1131_U421 = ~new_P2_R1131_U152 | ~new_P2_R1131_U153;
  assign new_P2_R1131_U422 = ~new_P2_R1131_U300 | ~new_P2_R1131_U420;
  assign new_P2_R1131_U423 = ~new_P2_U3059 | ~new_P2_R1131_U49;
  assign new_P2_R1131_U424 = ~new_P2_U3951 | ~new_P2_R1131_U48;
  assign new_P2_R1131_U425 = ~new_P2_U3060 | ~new_P2_R1131_U50;
  assign new_P2_R1131_U426 = ~new_P2_U3952 | ~new_P2_R1131_U51;
  assign new_P2_R1131_U427 = ~new_P2_R1131_U426 | ~new_P2_R1131_U425;
  assign new_P2_R1131_U428 = ~new_P2_R1131_U357 | ~new_P2_R1131_U89;
  assign new_P2_R1131_U429 = ~new_P2_R1131_U427 | ~new_P2_R1131_U307;
  assign new_P2_R1131_U430 = ~new_P2_U3067 | ~new_P2_R1131_U52;
  assign new_P2_R1131_U431 = ~new_P2_U3953 | ~new_P2_R1131_U53;
  assign new_P2_R1131_U432 = ~new_P2_R1131_U431 | ~new_P2_R1131_U430;
  assign new_P2_R1131_U433 = ~new_P2_R1131_U358 | ~new_P2_R1131_U155;
  assign new_P2_R1131_U434 = ~new_P2_R1131_U294 | ~new_P2_R1131_U432;
  assign new_P2_R1131_U435 = ~new_P2_U3068 | ~new_P2_R1131_U84;
  assign new_P2_R1131_U436 = ~new_P2_U3954 | ~new_P2_R1131_U85;
  assign new_P2_R1131_U437 = ~new_P2_U3068 | ~new_P2_R1131_U84;
  assign new_P2_R1131_U438 = ~new_P2_U3954 | ~new_P2_R1131_U85;
  assign new_P2_R1131_U439 = ~new_P2_R1131_U438 | ~new_P2_R1131_U437;
  assign new_P2_R1131_U440 = ~new_P2_R1131_U156 | ~new_P2_R1131_U157;
  assign new_P2_R1131_U441 = ~new_P2_R1131_U290 | ~new_P2_R1131_U439;
  assign new_P2_R1131_U442 = ~new_P2_U3063 | ~new_P2_R1131_U82;
  assign new_P2_R1131_U443 = ~new_P2_U3955 | ~new_P2_R1131_U83;
  assign new_P2_R1131_U444 = ~new_P2_U3063 | ~new_P2_R1131_U82;
  assign new_P2_R1131_U445 = ~new_P2_U3955 | ~new_P2_R1131_U83;
  assign new_P2_R1131_U446 = ~new_P2_R1131_U445 | ~new_P2_R1131_U444;
  assign new_P2_R1131_U447 = ~new_P2_R1131_U158 | ~new_P2_R1131_U159;
  assign new_P2_R1131_U448 = ~new_P2_R1131_U286 | ~new_P2_R1131_U446;
  assign new_P2_R1131_U449 = ~new_P2_U3077 | ~new_P2_R1131_U54;
  assign new_P2_R1131_U450 = ~new_P2_U3956 | ~new_P2_R1131_U55;
  assign new_P2_R1131_U451 = ~new_P2_U3077 | ~new_P2_R1131_U54;
  assign new_P2_R1131_U452 = ~new_P2_U3956 | ~new_P2_R1131_U55;
  assign new_P2_R1131_U453 = ~new_P2_R1131_U452 | ~new_P2_R1131_U451;
  assign new_P2_R1131_U454 = ~new_P2_U3078 | ~new_P2_R1131_U81;
  assign new_P2_R1131_U455 = ~new_P2_U3957 | ~new_P2_R1131_U90;
  assign new_P2_R1131_U456 = ~new_P2_R1131_U182 | ~new_P2_R1131_U161;
  assign new_P2_R1131_U457 = ~new_P2_R1131_U328 | ~new_P2_R1131_U31;
  assign new_P2_R1131_U458 = ~new_P2_U3083 | ~new_P2_R1131_U78;
  assign new_P2_R1131_U459 = ~new_P2_U3485 | ~new_P2_R1131_U79;
  assign new_P2_R1131_U460 = ~new_P2_R1131_U459 | ~new_P2_R1131_U458;
  assign new_P2_R1131_U461 = ~new_P2_R1131_U359 | ~new_P2_R1131_U91;
  assign new_P2_R1131_U462 = ~new_P2_R1131_U460 | ~new_P2_R1131_U316;
  assign new_P2_R1131_U463 = ~new_P2_U3084 | ~new_P2_R1131_U75;
  assign new_P2_R1131_U464 = ~new_P2_U3483 | ~new_P2_R1131_U76;
  assign new_P2_R1131_U465 = ~new_P2_R1131_U464 | ~new_P2_R1131_U463;
  assign new_P2_R1131_U466 = ~new_P2_R1131_U360 | ~new_P2_R1131_U162;
  assign new_P2_R1131_U467 = ~new_P2_R1131_U270 | ~new_P2_R1131_U465;
  assign new_P2_R1131_U468 = ~new_P2_U3071 | ~new_P2_R1131_U60;
  assign new_P2_R1131_U469 = ~new_P2_U3480 | ~new_P2_R1131_U58;
  assign new_P2_R1131_U470 = ~new_P2_U3075 | ~new_P2_R1131_U56;
  assign new_P2_R1131_U471 = ~new_P2_U3477 | ~new_P2_R1131_U57;
  assign new_P2_R1131_U472 = ~new_P2_R1131_U471 | ~new_P2_R1131_U470;
  assign new_P2_R1131_U473 = ~new_P2_R1131_U361 | ~new_P2_R1131_U92;
  assign new_P2_R1131_U474 = ~new_P2_R1131_U472 | ~new_P2_R1131_U262;
  assign new_P2_R1131_U475 = ~new_P2_U3076 | ~new_P2_R1131_U73;
  assign new_P2_R1131_U476 = ~new_P2_U3474 | ~new_P2_R1131_U74;
  assign new_P2_R1131_U477 = ~new_P2_U3076 | ~new_P2_R1131_U73;
  assign new_P2_R1131_U478 = ~new_P2_U3474 | ~new_P2_R1131_U74;
  assign new_P2_R1131_U479 = ~new_P2_R1131_U478 | ~new_P2_R1131_U477;
  assign new_P2_R1131_U480 = ~new_P2_R1131_U163 | ~new_P2_R1131_U164;
  assign new_P2_R1131_U481 = ~new_P2_R1131_U258 | ~new_P2_R1131_U479;
  assign new_P2_R1131_U482 = ~new_P2_U3081 | ~new_P2_R1131_U71;
  assign new_P2_R1131_U483 = ~new_P2_U3471 | ~new_P2_R1131_U72;
  assign new_P2_R1131_U484 = ~new_P2_U3081 | ~new_P2_R1131_U71;
  assign new_P2_R1131_U485 = ~new_P2_U3471 | ~new_P2_R1131_U72;
  assign new_P2_R1131_U486 = ~new_P2_R1131_U485 | ~new_P2_R1131_U484;
  assign new_P2_R1131_U487 = ~new_P2_R1131_U165 | ~new_P2_R1131_U166;
  assign new_P2_R1131_U488 = ~new_P2_R1131_U254 | ~new_P2_R1131_U486;
  assign new_P2_R1131_U489 = ~new_P2_U3082 | ~new_P2_R1131_U69;
  assign new_P2_R1131_U490 = ~new_P2_U3468 | ~new_P2_R1131_U70;
  assign new_P2_R1131_U491 = ~new_P2_U3074 | ~new_P2_R1131_U64;
  assign new_P2_R1131_U492 = ~new_P2_U3465 | ~new_P2_R1131_U65;
  assign new_P2_R1131_U493 = ~new_P2_R1131_U492 | ~new_P2_R1131_U491;
  assign new_P2_R1131_U494 = ~new_P2_R1131_U362 | ~new_P2_R1131_U93;
  assign new_P2_R1131_U495 = ~new_P2_R1131_U493 | ~new_P2_R1131_U338;
  assign new_P2_R1131_U496 = ~new_P2_U3065 | ~new_P2_R1131_U66;
  assign new_P2_R1131_U497 = ~new_P2_U3462 | ~new_P2_R1131_U67;
  assign new_P2_R1131_U498 = ~new_P2_R1131_U497 | ~new_P2_R1131_U496;
  assign new_P2_R1131_U499 = ~new_P2_R1131_U363 | ~new_P2_R1131_U167;
  assign new_P2_R1131_U500 = ~new_P2_R1131_U244 | ~new_P2_R1131_U498;
  assign new_P2_R1131_U501 = ~new_P2_U3064 | ~new_P2_R1131_U62;
  assign new_P2_R1131_U502 = ~new_P2_U3459 | ~new_P2_R1131_U63;
  assign new_P2_R1131_U503 = ~new_P2_U3079 | ~new_P2_R1131_U29;
  assign new_P2_R1131_U504 = ~new_P2_U3427 | ~new_P2_R1131_U30;
  assign new_P2_R1146_U6 = new_P2_R1146_U202 & new_P2_R1146_U201;
  assign new_P2_R1146_U7 = new_P2_R1146_U241 & new_P2_R1146_U240;
  assign new_P2_R1146_U8 = new_P2_R1146_U181 & new_P2_R1146_U256;
  assign new_P2_R1146_U9 = new_P2_R1146_U258 & new_P2_R1146_U257;
  assign new_P2_R1146_U10 = new_P2_R1146_U182 & new_P2_R1146_U282;
  assign new_P2_R1146_U11 = new_P2_R1146_U284 & new_P2_R1146_U283;
  assign new_P2_R1146_U12 = ~new_P2_R1146_U344 | ~new_P2_R1146_U347;
  assign new_P2_R1146_U13 = ~new_P2_R1146_U333 | ~new_P2_R1146_U336;
  assign new_P2_R1146_U14 = ~new_P2_R1146_U322 | ~new_P2_R1146_U325;
  assign new_P2_R1146_U15 = ~new_P2_R1146_U314 | ~new_P2_R1146_U316;
  assign new_P2_R1146_U16 = ~new_P2_R1146_U352 | ~new_P2_R1146_U312;
  assign new_P2_R1146_U17 = ~new_P2_R1146_U235 | ~new_P2_R1146_U237;
  assign new_P2_R1146_U18 = ~new_P2_R1146_U227 | ~new_P2_R1146_U230;
  assign new_P2_R1146_U19 = ~new_P2_R1146_U219 | ~new_P2_R1146_U221;
  assign new_P2_R1146_U20 = ~new_P2_R1146_U166 | ~new_P2_R1146_U350;
  assign new_P2_R1146_U21 = ~new_P2_U3450;
  assign new_P2_R1146_U22 = ~new_P2_U3444;
  assign new_P2_R1146_U23 = ~new_P2_U3435;
  assign new_P2_R1146_U24 = ~new_P2_U3427;
  assign new_P2_R1146_U25 = ~new_P2_U3080;
  assign new_P2_R1146_U26 = ~new_P2_U3438;
  assign new_P2_R1146_U27 = ~new_P2_U3070;
  assign new_P2_R1146_U28 = ~new_P2_U3070 | ~new_P2_R1146_U23;
  assign new_P2_R1146_U29 = ~new_P2_U3066;
  assign new_P2_R1146_U30 = ~new_P2_U3447;
  assign new_P2_R1146_U31 = ~new_P2_U3441;
  assign new_P2_R1146_U32 = ~new_P2_U3073;
  assign new_P2_R1146_U33 = ~new_P2_U3069;
  assign new_P2_R1146_U34 = ~new_P2_U3062;
  assign new_P2_R1146_U35 = ~new_P2_U3062 | ~new_P2_R1146_U31;
  assign new_P2_R1146_U36 = ~new_P2_U3453;
  assign new_P2_R1146_U37 = ~new_P2_U3072;
  assign new_P2_R1146_U38 = ~new_P2_U3072 | ~new_P2_R1146_U21;
  assign new_P2_R1146_U39 = ~new_P2_U3086;
  assign new_P2_R1146_U40 = ~new_P2_U3456;
  assign new_P2_R1146_U41 = ~new_P2_U3085;
  assign new_P2_R1146_U42 = ~new_P2_R1146_U208 | ~new_P2_R1146_U207;
  assign new_P2_R1146_U43 = ~new_P2_R1146_U35 | ~new_P2_R1146_U223;
  assign new_P2_R1146_U44 = ~new_P2_R1146_U351 | ~new_P2_R1146_U192 | ~new_P2_R1146_U176;
  assign new_P2_R1146_U45 = ~new_P2_U3951;
  assign new_P2_R1146_U46 = ~new_P2_U3459;
  assign new_P2_R1146_U47 = ~new_P2_U3462;
  assign new_P2_R1146_U48 = ~new_P2_U3065;
  assign new_P2_R1146_U49 = ~new_P2_U3064;
  assign new_P2_R1146_U50 = ~new_P2_U3085 | ~new_P2_R1146_U40;
  assign new_P2_R1146_U51 = ~new_P2_U3465;
  assign new_P2_R1146_U52 = ~new_P2_U3074;
  assign new_P2_R1146_U53 = ~new_P2_U3468;
  assign new_P2_R1146_U54 = ~new_P2_U3082;
  assign new_P2_R1146_U55 = ~new_P2_U3477;
  assign new_P2_R1146_U56 = ~new_P2_U3474;
  assign new_P2_R1146_U57 = ~new_P2_U3471;
  assign new_P2_R1146_U58 = ~new_P2_U3075;
  assign new_P2_R1146_U59 = ~new_P2_U3076;
  assign new_P2_R1146_U60 = ~new_P2_U3081;
  assign new_P2_R1146_U61 = ~new_P2_U3081 | ~new_P2_R1146_U57;
  assign new_P2_R1146_U62 = ~new_P2_U3480;
  assign new_P2_R1146_U63 = ~new_P2_U3071;
  assign new_P2_R1146_U64 = ~new_P2_R1146_U268 | ~new_P2_R1146_U267;
  assign new_P2_R1146_U65 = ~new_P2_U3084;
  assign new_P2_R1146_U66 = ~new_P2_U3485;
  assign new_P2_R1146_U67 = ~new_P2_U3083;
  assign new_P2_R1146_U68 = ~new_P2_U3957;
  assign new_P2_R1146_U69 = ~new_P2_U3078;
  assign new_P2_R1146_U70 = ~new_P2_U3954;
  assign new_P2_R1146_U71 = ~new_P2_U3955;
  assign new_P2_R1146_U72 = ~new_P2_U3956;
  assign new_P2_R1146_U73 = ~new_P2_U3068;
  assign new_P2_R1146_U74 = ~new_P2_U3063;
  assign new_P2_R1146_U75 = ~new_P2_U3077;
  assign new_P2_R1146_U76 = ~new_P2_U3077 | ~new_P2_R1146_U72;
  assign new_P2_R1146_U77 = ~new_P2_U3953;
  assign new_P2_R1146_U78 = ~new_P2_U3067;
  assign new_P2_R1146_U79 = ~new_P2_U3952;
  assign new_P2_R1146_U80 = ~new_P2_U3060;
  assign new_P2_R1146_U81 = ~new_P2_U3950;
  assign new_P2_R1146_U82 = ~new_P2_U3059;
  assign new_P2_R1146_U83 = ~new_P2_U3059 | ~new_P2_R1146_U45;
  assign new_P2_R1146_U84 = ~new_P2_U3055;
  assign new_P2_R1146_U85 = ~new_P2_U3949;
  assign new_P2_R1146_U86 = ~new_P2_U3056;
  assign new_P2_R1146_U87 = ~new_P2_R1146_U128 | ~new_P2_R1146_U301;
  assign new_P2_R1146_U88 = ~new_P2_R1146_U298 | ~new_P2_R1146_U297;
  assign new_P2_R1146_U89 = ~new_P2_R1146_U76 | ~new_P2_R1146_U318;
  assign new_P2_R1146_U90 = ~new_P2_R1146_U61 | ~new_P2_R1146_U329;
  assign new_P2_R1146_U91 = ~new_P2_R1146_U50 | ~new_P2_R1146_U340;
  assign new_P2_R1146_U92 = ~new_P2_U3079;
  assign new_P2_R1146_U93 = ~new_P2_R1146_U395 | ~new_P2_R1146_U394;
  assign new_P2_R1146_U94 = ~new_P2_R1146_U409 | ~new_P2_R1146_U408;
  assign new_P2_R1146_U95 = ~new_P2_R1146_U414 | ~new_P2_R1146_U413;
  assign new_P2_R1146_U96 = ~new_P2_R1146_U430 | ~new_P2_R1146_U429;
  assign new_P2_R1146_U97 = ~new_P2_R1146_U435 | ~new_P2_R1146_U434;
  assign new_P2_R1146_U98 = ~new_P2_R1146_U440 | ~new_P2_R1146_U439;
  assign new_P2_R1146_U99 = ~new_P2_R1146_U445 | ~new_P2_R1146_U444;
  assign new_P2_R1146_U100 = ~new_P2_R1146_U450 | ~new_P2_R1146_U449;
  assign new_P2_R1146_U101 = ~new_P2_R1146_U466 | ~new_P2_R1146_U465;
  assign new_P2_R1146_U102 = ~new_P2_R1146_U471 | ~new_P2_R1146_U470;
  assign new_P2_R1146_U103 = ~new_P2_R1146_U356 | ~new_P2_R1146_U355;
  assign new_P2_R1146_U104 = ~new_P2_R1146_U365 | ~new_P2_R1146_U364;
  assign new_P2_R1146_U105 = ~new_P2_R1146_U372 | ~new_P2_R1146_U371;
  assign new_P2_R1146_U106 = ~new_P2_R1146_U376 | ~new_P2_R1146_U375;
  assign new_P2_R1146_U107 = ~new_P2_R1146_U385 | ~new_P2_R1146_U384;
  assign new_P2_R1146_U108 = ~new_P2_R1146_U404 | ~new_P2_R1146_U403;
  assign new_P2_R1146_U109 = ~new_P2_R1146_U421 | ~new_P2_R1146_U420;
  assign new_P2_R1146_U110 = ~new_P2_R1146_U425 | ~new_P2_R1146_U424;
  assign new_P2_R1146_U111 = ~new_P2_R1146_U457 | ~new_P2_R1146_U456;
  assign new_P2_R1146_U112 = ~new_P2_R1146_U461 | ~new_P2_R1146_U460;
  assign new_P2_R1146_U113 = ~new_P2_R1146_U478 | ~new_P2_R1146_U477;
  assign new_P2_R1146_U114 = new_P2_R1146_U194 & new_P2_R1146_U184;
  assign new_P2_R1146_U115 = new_P2_R1146_U197 & new_P2_R1146_U198;
  assign new_P2_R1146_U116 = new_P2_R1146_U185 & new_P2_R1146_U205 & new_P2_R1146_U200;
  assign new_P2_R1146_U117 = new_P2_R1146_U210 & new_P2_R1146_U186;
  assign new_P2_R1146_U118 = new_P2_R1146_U213 & new_P2_R1146_U214;
  assign new_P2_R1146_U119 = new_P2_R1146_U38 & new_P2_R1146_U358 & new_P2_R1146_U357;
  assign new_P2_R1146_U120 = new_P2_R1146_U361 & new_P2_R1146_U186;
  assign new_P2_R1146_U121 = new_P2_R1146_U229 & new_P2_R1146_U6;
  assign new_P2_R1146_U122 = new_P2_R1146_U368 & new_P2_R1146_U185;
  assign new_P2_R1146_U123 = new_P2_R1146_U28 & new_P2_R1146_U378 & new_P2_R1146_U377;
  assign new_P2_R1146_U124 = new_P2_R1146_U381 & new_P2_R1146_U184;
  assign new_P2_R1146_U125 = new_P2_R1146_U180 & new_P2_R1146_U239 & new_P2_R1146_U216;
  assign new_P2_R1146_U126 = new_P2_R1146_U261 & new_P2_R1146_U8;
  assign new_P2_R1146_U127 = new_P2_R1146_U287 & new_P2_R1146_U10;
  assign new_P2_R1146_U128 = new_P2_R1146_U303 & new_P2_R1146_U304;
  assign new_P2_R1146_U129 = new_P2_R1146_U311 & new_P2_R1146_U387 & new_P2_R1146_U386;
  assign new_P2_R1146_U130 = new_P2_R1146_U308 & new_P2_R1146_U390;
  assign new_P2_R1146_U131 = ~new_P2_R1146_U392 | ~new_P2_R1146_U391;
  assign new_P2_R1146_U132 = new_P2_R1146_U83 & new_P2_R1146_U397 & new_P2_R1146_U396;
  assign new_P2_R1146_U133 = new_P2_R1146_U400 & new_P2_R1146_U183;
  assign new_P2_R1146_U134 = ~new_P2_R1146_U406 | ~new_P2_R1146_U405;
  assign new_P2_R1146_U135 = ~new_P2_R1146_U411 | ~new_P2_R1146_U410;
  assign new_P2_R1146_U136 = new_P2_R1146_U324 & new_P2_R1146_U11;
  assign new_P2_R1146_U137 = new_P2_R1146_U417 & new_P2_R1146_U182;
  assign new_P2_R1146_U138 = ~new_P2_R1146_U427 | ~new_P2_R1146_U426;
  assign new_P2_R1146_U139 = ~new_P2_R1146_U432 | ~new_P2_R1146_U431;
  assign new_P2_R1146_U140 = ~new_P2_R1146_U437 | ~new_P2_R1146_U436;
  assign new_P2_R1146_U141 = ~new_P2_R1146_U442 | ~new_P2_R1146_U441;
  assign new_P2_R1146_U142 = ~new_P2_R1146_U447 | ~new_P2_R1146_U446;
  assign new_P2_R1146_U143 = new_P2_R1146_U335 & new_P2_R1146_U9;
  assign new_P2_R1146_U144 = new_P2_R1146_U453 & new_P2_R1146_U181;
  assign new_P2_R1146_U145 = ~new_P2_R1146_U463 | ~new_P2_R1146_U462;
  assign new_P2_R1146_U146 = ~new_P2_R1146_U468 | ~new_P2_R1146_U467;
  assign new_P2_R1146_U147 = new_P2_R1146_U346 & new_P2_R1146_U7;
  assign new_P2_R1146_U148 = new_P2_R1146_U474 & new_P2_R1146_U180;
  assign new_P2_R1146_U149 = new_P2_R1146_U354 & new_P2_R1146_U353;
  assign new_P2_R1146_U150 = ~new_P2_R1146_U118 | ~new_P2_R1146_U211;
  assign new_P2_R1146_U151 = new_P2_R1146_U363 & new_P2_R1146_U362;
  assign new_P2_R1146_U152 = new_P2_R1146_U370 & new_P2_R1146_U369;
  assign new_P2_R1146_U153 = new_P2_R1146_U374 & new_P2_R1146_U373;
  assign new_P2_R1146_U154 = ~new_P2_R1146_U115 | ~new_P2_R1146_U195;
  assign new_P2_R1146_U155 = new_P2_R1146_U383 & new_P2_R1146_U382;
  assign new_P2_R1146_U156 = ~new_P2_U3960;
  assign new_P2_R1146_U157 = ~new_P2_U3057;
  assign new_P2_R1146_U158 = new_P2_R1146_U402 & new_P2_R1146_U401;
  assign new_P2_R1146_U159 = ~new_P2_R1146_U294 | ~new_P2_R1146_U293;
  assign new_P2_R1146_U160 = ~new_P2_R1146_U290 | ~new_P2_R1146_U289;
  assign new_P2_R1146_U161 = new_P2_R1146_U419 & new_P2_R1146_U418;
  assign new_P2_R1146_U162 = new_P2_R1146_U423 & new_P2_R1146_U422;
  assign new_P2_R1146_U163 = ~new_P2_R1146_U280 | ~new_P2_R1146_U279;
  assign new_P2_R1146_U164 = ~new_P2_R1146_U276 | ~new_P2_R1146_U275;
  assign new_P2_R1146_U165 = ~new_P2_U3432;
  assign new_P2_R1146_U166 = ~new_P2_U3427 | ~new_P2_R1146_U92;
  assign new_P2_R1146_U167 = ~new_P2_R1146_U272 | ~new_P2_R1146_U271;
  assign new_P2_R1146_U168 = ~new_P2_U3483;
  assign new_P2_R1146_U169 = ~new_P2_R1146_U264 | ~new_P2_R1146_U263;
  assign new_P2_R1146_U170 = new_P2_R1146_U455 & new_P2_R1146_U454;
  assign new_P2_R1146_U171 = new_P2_R1146_U459 & new_P2_R1146_U458;
  assign new_P2_R1146_U172 = ~new_P2_R1146_U254 | ~new_P2_R1146_U253;
  assign new_P2_R1146_U173 = ~new_P2_R1146_U250 | ~new_P2_R1146_U249;
  assign new_P2_R1146_U174 = ~new_P2_R1146_U246 | ~new_P2_R1146_U245;
  assign new_P2_R1146_U175 = new_P2_R1146_U476 & new_P2_R1146_U475;
  assign new_P2_R1146_U176 = ~new_P2_R1146_U166 | ~new_P2_R1146_U165;
  assign new_P2_R1146_U177 = ~new_P2_R1146_U83;
  assign new_P2_R1146_U178 = ~new_P2_R1146_U28;
  assign new_P2_R1146_U179 = ~new_P2_R1146_U38;
  assign new_P2_R1146_U180 = ~new_P2_U3459 | ~new_P2_R1146_U49;
  assign new_P2_R1146_U181 = ~new_P2_U3474 | ~new_P2_R1146_U59;
  assign new_P2_R1146_U182 = ~new_P2_U3955 | ~new_P2_R1146_U74;
  assign new_P2_R1146_U183 = ~new_P2_U3951 | ~new_P2_R1146_U82;
  assign new_P2_R1146_U184 = ~new_P2_U3435 | ~new_P2_R1146_U27;
  assign new_P2_R1146_U185 = ~new_P2_U3444 | ~new_P2_R1146_U33;
  assign new_P2_R1146_U186 = ~new_P2_U3450 | ~new_P2_R1146_U37;
  assign new_P2_R1146_U187 = ~new_P2_R1146_U61;
  assign new_P2_R1146_U188 = ~new_P2_R1146_U76;
  assign new_P2_R1146_U189 = ~new_P2_R1146_U35;
  assign new_P2_R1146_U190 = ~new_P2_R1146_U50;
  assign new_P2_R1146_U191 = ~new_P2_R1146_U166;
  assign new_P2_R1146_U192 = ~new_P2_U3080 | ~new_P2_R1146_U166;
  assign new_P2_R1146_U193 = ~new_P2_R1146_U44;
  assign new_P2_R1146_U194 = ~new_P2_U3438 | ~new_P2_R1146_U29;
  assign new_P2_R1146_U195 = ~new_P2_R1146_U114 | ~new_P2_R1146_U44;
  assign new_P2_R1146_U196 = ~new_P2_R1146_U29 | ~new_P2_R1146_U28;
  assign new_P2_R1146_U197 = ~new_P2_R1146_U196 | ~new_P2_R1146_U26;
  assign new_P2_R1146_U198 = ~new_P2_U3066 | ~new_P2_R1146_U178;
  assign new_P2_R1146_U199 = ~new_P2_R1146_U154;
  assign new_P2_R1146_U200 = ~new_P2_U3447 | ~new_P2_R1146_U32;
  assign new_P2_R1146_U201 = ~new_P2_U3073 | ~new_P2_R1146_U30;
  assign new_P2_R1146_U202 = ~new_P2_U3069 | ~new_P2_R1146_U22;
  assign new_P2_R1146_U203 = ~new_P2_R1146_U189 | ~new_P2_R1146_U185;
  assign new_P2_R1146_U204 = ~new_P2_R1146_U6 | ~new_P2_R1146_U203;
  assign new_P2_R1146_U205 = ~new_P2_U3441 | ~new_P2_R1146_U34;
  assign new_P2_R1146_U206 = ~new_P2_U3447 | ~new_P2_R1146_U32;
  assign new_P2_R1146_U207 = ~new_P2_R1146_U154 | ~new_P2_R1146_U116;
  assign new_P2_R1146_U208 = ~new_P2_R1146_U206 | ~new_P2_R1146_U204;
  assign new_P2_R1146_U209 = ~new_P2_R1146_U42;
  assign new_P2_R1146_U210 = ~new_P2_U3453 | ~new_P2_R1146_U39;
  assign new_P2_R1146_U211 = ~new_P2_R1146_U117 | ~new_P2_R1146_U42;
  assign new_P2_R1146_U212 = ~new_P2_R1146_U39 | ~new_P2_R1146_U38;
  assign new_P2_R1146_U213 = ~new_P2_R1146_U212 | ~new_P2_R1146_U36;
  assign new_P2_R1146_U214 = ~new_P2_U3086 | ~new_P2_R1146_U179;
  assign new_P2_R1146_U215 = ~new_P2_R1146_U150;
  assign new_P2_R1146_U216 = ~new_P2_U3456 | ~new_P2_R1146_U41;
  assign new_P2_R1146_U217 = ~new_P2_R1146_U216 | ~new_P2_R1146_U50;
  assign new_P2_R1146_U218 = ~new_P2_R1146_U209 | ~new_P2_R1146_U38;
  assign new_P2_R1146_U219 = ~new_P2_R1146_U120 | ~new_P2_R1146_U218;
  assign new_P2_R1146_U220 = ~new_P2_R1146_U42 | ~new_P2_R1146_U186;
  assign new_P2_R1146_U221 = ~new_P2_R1146_U119 | ~new_P2_R1146_U220;
  assign new_P2_R1146_U222 = ~new_P2_R1146_U38 | ~new_P2_R1146_U186;
  assign new_P2_R1146_U223 = ~new_P2_R1146_U205 | ~new_P2_R1146_U154;
  assign new_P2_R1146_U224 = ~new_P2_R1146_U43;
  assign new_P2_R1146_U225 = ~new_P2_U3069 | ~new_P2_R1146_U22;
  assign new_P2_R1146_U226 = ~new_P2_R1146_U224 | ~new_P2_R1146_U225;
  assign new_P2_R1146_U227 = ~new_P2_R1146_U122 | ~new_P2_R1146_U226;
  assign new_P2_R1146_U228 = ~new_P2_R1146_U43 | ~new_P2_R1146_U185;
  assign new_P2_R1146_U229 = ~new_P2_U3447 | ~new_P2_R1146_U32;
  assign new_P2_R1146_U230 = ~new_P2_R1146_U121 | ~new_P2_R1146_U228;
  assign new_P2_R1146_U231 = ~new_P2_U3069 | ~new_P2_R1146_U22;
  assign new_P2_R1146_U232 = ~new_P2_R1146_U185 | ~new_P2_R1146_U231;
  assign new_P2_R1146_U233 = ~new_P2_R1146_U205 | ~new_P2_R1146_U35;
  assign new_P2_R1146_U234 = ~new_P2_R1146_U193 | ~new_P2_R1146_U28;
  assign new_P2_R1146_U235 = ~new_P2_R1146_U124 | ~new_P2_R1146_U234;
  assign new_P2_R1146_U236 = ~new_P2_R1146_U44 | ~new_P2_R1146_U184;
  assign new_P2_R1146_U237 = ~new_P2_R1146_U123 | ~new_P2_R1146_U236;
  assign new_P2_R1146_U238 = ~new_P2_R1146_U28 | ~new_P2_R1146_U184;
  assign new_P2_R1146_U239 = ~new_P2_U3462 | ~new_P2_R1146_U48;
  assign new_P2_R1146_U240 = ~new_P2_U3065 | ~new_P2_R1146_U47;
  assign new_P2_R1146_U241 = ~new_P2_U3064 | ~new_P2_R1146_U46;
  assign new_P2_R1146_U242 = ~new_P2_R1146_U190 | ~new_P2_R1146_U180;
  assign new_P2_R1146_U243 = ~new_P2_R1146_U7 | ~new_P2_R1146_U242;
  assign new_P2_R1146_U244 = ~new_P2_U3462 | ~new_P2_R1146_U48;
  assign new_P2_R1146_U245 = ~new_P2_R1146_U150 | ~new_P2_R1146_U125;
  assign new_P2_R1146_U246 = ~new_P2_R1146_U244 | ~new_P2_R1146_U243;
  assign new_P2_R1146_U247 = ~new_P2_R1146_U174;
  assign new_P2_R1146_U248 = ~new_P2_U3465 | ~new_P2_R1146_U52;
  assign new_P2_R1146_U249 = ~new_P2_R1146_U248 | ~new_P2_R1146_U174;
  assign new_P2_R1146_U250 = ~new_P2_U3074 | ~new_P2_R1146_U51;
  assign new_P2_R1146_U251 = ~new_P2_R1146_U173;
  assign new_P2_R1146_U252 = ~new_P2_U3468 | ~new_P2_R1146_U54;
  assign new_P2_R1146_U253 = ~new_P2_R1146_U252 | ~new_P2_R1146_U173;
  assign new_P2_R1146_U254 = ~new_P2_U3082 | ~new_P2_R1146_U53;
  assign new_P2_R1146_U255 = ~new_P2_R1146_U172;
  assign new_P2_R1146_U256 = ~new_P2_U3477 | ~new_P2_R1146_U58;
  assign new_P2_R1146_U257 = ~new_P2_U3075 | ~new_P2_R1146_U55;
  assign new_P2_R1146_U258 = ~new_P2_U3076 | ~new_P2_R1146_U56;
  assign new_P2_R1146_U259 = ~new_P2_R1146_U187 | ~new_P2_R1146_U8;
  assign new_P2_R1146_U260 = ~new_P2_R1146_U9 | ~new_P2_R1146_U259;
  assign new_P2_R1146_U261 = ~new_P2_U3471 | ~new_P2_R1146_U60;
  assign new_P2_R1146_U262 = ~new_P2_U3477 | ~new_P2_R1146_U58;
  assign new_P2_R1146_U263 = ~new_P2_R1146_U126 | ~new_P2_R1146_U172;
  assign new_P2_R1146_U264 = ~new_P2_R1146_U262 | ~new_P2_R1146_U260;
  assign new_P2_R1146_U265 = ~new_P2_R1146_U169;
  assign new_P2_R1146_U266 = ~new_P2_U3480 | ~new_P2_R1146_U63;
  assign new_P2_R1146_U267 = ~new_P2_R1146_U266 | ~new_P2_R1146_U169;
  assign new_P2_R1146_U268 = ~new_P2_U3071 | ~new_P2_R1146_U62;
  assign new_P2_R1146_U269 = ~new_P2_R1146_U64;
  assign new_P2_R1146_U270 = ~new_P2_R1146_U269 | ~new_P2_R1146_U65;
  assign new_P2_R1146_U271 = ~new_P2_R1146_U270 | ~new_P2_R1146_U168;
  assign new_P2_R1146_U272 = ~new_P2_U3084 | ~new_P2_R1146_U64;
  assign new_P2_R1146_U273 = ~new_P2_R1146_U167;
  assign new_P2_R1146_U274 = ~new_P2_U3485 | ~new_P2_R1146_U67;
  assign new_P2_R1146_U275 = ~new_P2_R1146_U274 | ~new_P2_R1146_U167;
  assign new_P2_R1146_U276 = ~new_P2_U3083 | ~new_P2_R1146_U66;
  assign new_P2_R1146_U277 = ~new_P2_R1146_U164;
  assign new_P2_R1146_U278 = ~new_P2_U3957 | ~new_P2_R1146_U69;
  assign new_P2_R1146_U279 = ~new_P2_R1146_U278 | ~new_P2_R1146_U164;
  assign new_P2_R1146_U280 = ~new_P2_U3078 | ~new_P2_R1146_U68;
  assign new_P2_R1146_U281 = ~new_P2_R1146_U163;
  assign new_P2_R1146_U282 = ~new_P2_U3954 | ~new_P2_R1146_U73;
  assign new_P2_R1146_U283 = ~new_P2_U3068 | ~new_P2_R1146_U70;
  assign new_P2_R1146_U284 = ~new_P2_U3063 | ~new_P2_R1146_U71;
  assign new_P2_R1146_U285 = ~new_P2_R1146_U188 | ~new_P2_R1146_U10;
  assign new_P2_R1146_U286 = ~new_P2_R1146_U11 | ~new_P2_R1146_U285;
  assign new_P2_R1146_U287 = ~new_P2_U3956 | ~new_P2_R1146_U75;
  assign new_P2_R1146_U288 = ~new_P2_U3954 | ~new_P2_R1146_U73;
  assign new_P2_R1146_U289 = ~new_P2_R1146_U127 | ~new_P2_R1146_U163;
  assign new_P2_R1146_U290 = ~new_P2_R1146_U288 | ~new_P2_R1146_U286;
  assign new_P2_R1146_U291 = ~new_P2_R1146_U160;
  assign new_P2_R1146_U292 = ~new_P2_U3953 | ~new_P2_R1146_U78;
  assign new_P2_R1146_U293 = ~new_P2_R1146_U292 | ~new_P2_R1146_U160;
  assign new_P2_R1146_U294 = ~new_P2_U3067 | ~new_P2_R1146_U77;
  assign new_P2_R1146_U295 = ~new_P2_R1146_U159;
  assign new_P2_R1146_U296 = ~new_P2_U3952 | ~new_P2_R1146_U80;
  assign new_P2_R1146_U297 = ~new_P2_R1146_U296 | ~new_P2_R1146_U159;
  assign new_P2_R1146_U298 = ~new_P2_U3060 | ~new_P2_R1146_U79;
  assign new_P2_R1146_U299 = ~new_P2_R1146_U88;
  assign new_P2_R1146_U300 = ~new_P2_U3950 | ~new_P2_R1146_U84;
  assign new_P2_R1146_U301 = ~new_P2_R1146_U300 | ~new_P2_R1146_U88 | ~new_P2_R1146_U183;
  assign new_P2_R1146_U302 = ~new_P2_R1146_U84 | ~new_P2_R1146_U83;
  assign new_P2_R1146_U303 = ~new_P2_R1146_U302 | ~new_P2_R1146_U81;
  assign new_P2_R1146_U304 = ~new_P2_U3055 | ~new_P2_R1146_U177;
  assign new_P2_R1146_U305 = ~new_P2_R1146_U87;
  assign new_P2_R1146_U306 = ~new_P2_U3056 | ~new_P2_R1146_U85;
  assign new_P2_R1146_U307 = ~new_P2_R1146_U305 | ~new_P2_R1146_U306;
  assign new_P2_R1146_U308 = ~new_P2_U3949 | ~new_P2_R1146_U86;
  assign new_P2_R1146_U309 = ~new_P2_U3949 | ~new_P2_R1146_U86;
  assign new_P2_R1146_U310 = ~new_P2_R1146_U309 | ~new_P2_R1146_U87;
  assign new_P2_R1146_U311 = ~new_P2_U3056 | ~new_P2_R1146_U85;
  assign new_P2_R1146_U312 = ~new_P2_R1146_U129 | ~new_P2_R1146_U310;
  assign new_P2_R1146_U313 = ~new_P2_R1146_U299 | ~new_P2_R1146_U83;
  assign new_P2_R1146_U314 = ~new_P2_R1146_U133 | ~new_P2_R1146_U313;
  assign new_P2_R1146_U315 = ~new_P2_R1146_U88 | ~new_P2_R1146_U183;
  assign new_P2_R1146_U316 = ~new_P2_R1146_U132 | ~new_P2_R1146_U315;
  assign new_P2_R1146_U317 = ~new_P2_R1146_U83 | ~new_P2_R1146_U183;
  assign new_P2_R1146_U318 = ~new_P2_R1146_U287 | ~new_P2_R1146_U163;
  assign new_P2_R1146_U319 = ~new_P2_R1146_U89;
  assign new_P2_R1146_U320 = ~new_P2_U3063 | ~new_P2_R1146_U71;
  assign new_P2_R1146_U321 = ~new_P2_R1146_U319 | ~new_P2_R1146_U320;
  assign new_P2_R1146_U322 = ~new_P2_R1146_U137 | ~new_P2_R1146_U321;
  assign new_P2_R1146_U323 = ~new_P2_R1146_U89 | ~new_P2_R1146_U182;
  assign new_P2_R1146_U324 = ~new_P2_U3954 | ~new_P2_R1146_U73;
  assign new_P2_R1146_U325 = ~new_P2_R1146_U136 | ~new_P2_R1146_U323;
  assign new_P2_R1146_U326 = ~new_P2_U3063 | ~new_P2_R1146_U71;
  assign new_P2_R1146_U327 = ~new_P2_R1146_U182 | ~new_P2_R1146_U326;
  assign new_P2_R1146_U328 = ~new_P2_R1146_U287 | ~new_P2_R1146_U76;
  assign new_P2_R1146_U329 = ~new_P2_R1146_U261 | ~new_P2_R1146_U172;
  assign new_P2_R1146_U330 = ~new_P2_R1146_U90;
  assign new_P2_R1146_U331 = ~new_P2_U3076 | ~new_P2_R1146_U56;
  assign new_P2_R1146_U332 = ~new_P2_R1146_U330 | ~new_P2_R1146_U331;
  assign new_P2_R1146_U333 = ~new_P2_R1146_U144 | ~new_P2_R1146_U332;
  assign new_P2_R1146_U334 = ~new_P2_R1146_U90 | ~new_P2_R1146_U181;
  assign new_P2_R1146_U335 = ~new_P2_U3477 | ~new_P2_R1146_U58;
  assign new_P2_R1146_U336 = ~new_P2_R1146_U143 | ~new_P2_R1146_U334;
  assign new_P2_R1146_U337 = ~new_P2_U3076 | ~new_P2_R1146_U56;
  assign new_P2_R1146_U338 = ~new_P2_R1146_U181 | ~new_P2_R1146_U337;
  assign new_P2_R1146_U339 = ~new_P2_R1146_U261 | ~new_P2_R1146_U61;
  assign new_P2_R1146_U340 = ~new_P2_R1146_U216 | ~new_P2_R1146_U150;
  assign new_P2_R1146_U341 = ~new_P2_R1146_U91;
  assign new_P2_R1146_U342 = ~new_P2_U3064 | ~new_P2_R1146_U46;
  assign new_P2_R1146_U343 = ~new_P2_R1146_U341 | ~new_P2_R1146_U342;
  assign new_P2_R1146_U344 = ~new_P2_R1146_U148 | ~new_P2_R1146_U343;
  assign new_P2_R1146_U345 = ~new_P2_R1146_U91 | ~new_P2_R1146_U180;
  assign new_P2_R1146_U346 = ~new_P2_U3462 | ~new_P2_R1146_U48;
  assign new_P2_R1146_U347 = ~new_P2_R1146_U147 | ~new_P2_R1146_U345;
  assign new_P2_R1146_U348 = ~new_P2_U3064 | ~new_P2_R1146_U46;
  assign new_P2_R1146_U349 = ~new_P2_R1146_U180 | ~new_P2_R1146_U348;
  assign new_P2_R1146_U350 = ~new_P2_U3079 | ~new_P2_R1146_U24;
  assign new_P2_R1146_U351 = ~new_P2_U3080 | ~new_P2_R1146_U165;
  assign new_P2_R1146_U352 = ~new_P2_R1146_U130 | ~new_P2_R1146_U307;
  assign new_P2_R1146_U353 = ~new_P2_U3456 | ~new_P2_R1146_U41;
  assign new_P2_R1146_U354 = ~new_P2_U3085 | ~new_P2_R1146_U40;
  assign new_P2_R1146_U355 = ~new_P2_R1146_U217 | ~new_P2_R1146_U150;
  assign new_P2_R1146_U356 = ~new_P2_R1146_U215 | ~new_P2_R1146_U149;
  assign new_P2_R1146_U357 = ~new_P2_U3453 | ~new_P2_R1146_U39;
  assign new_P2_R1146_U358 = ~new_P2_U3086 | ~new_P2_R1146_U36;
  assign new_P2_R1146_U359 = ~new_P2_U3453 | ~new_P2_R1146_U39;
  assign new_P2_R1146_U360 = ~new_P2_U3086 | ~new_P2_R1146_U36;
  assign new_P2_R1146_U361 = ~new_P2_R1146_U360 | ~new_P2_R1146_U359;
  assign new_P2_R1146_U362 = ~new_P2_U3450 | ~new_P2_R1146_U37;
  assign new_P2_R1146_U363 = ~new_P2_U3072 | ~new_P2_R1146_U21;
  assign new_P2_R1146_U364 = ~new_P2_R1146_U222 | ~new_P2_R1146_U42;
  assign new_P2_R1146_U365 = ~new_P2_R1146_U151 | ~new_P2_R1146_U209;
  assign new_P2_R1146_U366 = ~new_P2_U3447 | ~new_P2_R1146_U32;
  assign new_P2_R1146_U367 = ~new_P2_U3073 | ~new_P2_R1146_U30;
  assign new_P2_R1146_U368 = ~new_P2_R1146_U367 | ~new_P2_R1146_U366;
  assign new_P2_R1146_U369 = ~new_P2_U3444 | ~new_P2_R1146_U33;
  assign new_P2_R1146_U370 = ~new_P2_U3069 | ~new_P2_R1146_U22;
  assign new_P2_R1146_U371 = ~new_P2_R1146_U232 | ~new_P2_R1146_U43;
  assign new_P2_R1146_U372 = ~new_P2_R1146_U152 | ~new_P2_R1146_U224;
  assign new_P2_R1146_U373 = ~new_P2_U3441 | ~new_P2_R1146_U34;
  assign new_P2_R1146_U374 = ~new_P2_U3062 | ~new_P2_R1146_U31;
  assign new_P2_R1146_U375 = ~new_P2_R1146_U233 | ~new_P2_R1146_U154;
  assign new_P2_R1146_U376 = ~new_P2_R1146_U199 | ~new_P2_R1146_U153;
  assign new_P2_R1146_U377 = ~new_P2_U3438 | ~new_P2_R1146_U29;
  assign new_P2_R1146_U378 = ~new_P2_U3066 | ~new_P2_R1146_U26;
  assign new_P2_R1146_U379 = ~new_P2_U3438 | ~new_P2_R1146_U29;
  assign new_P2_R1146_U380 = ~new_P2_U3066 | ~new_P2_R1146_U26;
  assign new_P2_R1146_U381 = ~new_P2_R1146_U380 | ~new_P2_R1146_U379;
  assign new_P2_R1146_U382 = ~new_P2_U3435 | ~new_P2_R1146_U27;
  assign new_P2_R1146_U383 = ~new_P2_U3070 | ~new_P2_R1146_U23;
  assign new_P2_R1146_U384 = ~new_P2_R1146_U238 | ~new_P2_R1146_U44;
  assign new_P2_R1146_U385 = ~new_P2_R1146_U155 | ~new_P2_R1146_U193;
  assign new_P2_R1146_U386 = ~new_P2_U3960 | ~new_P2_R1146_U157;
  assign new_P2_R1146_U387 = ~new_P2_U3057 | ~new_P2_R1146_U156;
  assign new_P2_R1146_U388 = ~new_P2_U3960 | ~new_P2_R1146_U157;
  assign new_P2_R1146_U389 = ~new_P2_U3057 | ~new_P2_R1146_U156;
  assign new_P2_R1146_U390 = ~new_P2_R1146_U389 | ~new_P2_R1146_U388;
  assign new_P2_R1146_U391 = ~new_P2_U3949 | ~new_P2_R1146_U86;
  assign new_P2_R1146_U392 = ~new_P2_U3056 | ~new_P2_R1146_U85;
  assign new_P2_R1146_U393 = ~new_P2_R1146_U131;
  assign new_P2_R1146_U394 = ~new_P2_R1146_U393 | ~new_P2_R1146_U305;
  assign new_P2_R1146_U395 = ~new_P2_R1146_U131 | ~new_P2_R1146_U87;
  assign new_P2_R1146_U396 = ~new_P2_U3950 | ~new_P2_R1146_U84;
  assign new_P2_R1146_U397 = ~new_P2_U3055 | ~new_P2_R1146_U81;
  assign new_P2_R1146_U398 = ~new_P2_U3950 | ~new_P2_R1146_U84;
  assign new_P2_R1146_U399 = ~new_P2_U3055 | ~new_P2_R1146_U81;
  assign new_P2_R1146_U400 = ~new_P2_R1146_U399 | ~new_P2_R1146_U398;
  assign new_P2_R1146_U401 = ~new_P2_U3951 | ~new_P2_R1146_U82;
  assign new_P2_R1146_U402 = ~new_P2_U3059 | ~new_P2_R1146_U45;
  assign new_P2_R1146_U403 = ~new_P2_R1146_U317 | ~new_P2_R1146_U88;
  assign new_P2_R1146_U404 = ~new_P2_R1146_U158 | ~new_P2_R1146_U299;
  assign new_P2_R1146_U405 = ~new_P2_U3952 | ~new_P2_R1146_U80;
  assign new_P2_R1146_U406 = ~new_P2_U3060 | ~new_P2_R1146_U79;
  assign new_P2_R1146_U407 = ~new_P2_R1146_U134;
  assign new_P2_R1146_U408 = ~new_P2_R1146_U295 | ~new_P2_R1146_U407;
  assign new_P2_R1146_U409 = ~new_P2_R1146_U134 | ~new_P2_R1146_U159;
  assign new_P2_R1146_U410 = ~new_P2_U3953 | ~new_P2_R1146_U78;
  assign new_P2_R1146_U411 = ~new_P2_U3067 | ~new_P2_R1146_U77;
  assign new_P2_R1146_U412 = ~new_P2_R1146_U135;
  assign new_P2_R1146_U413 = ~new_P2_R1146_U291 | ~new_P2_R1146_U412;
  assign new_P2_R1146_U414 = ~new_P2_R1146_U135 | ~new_P2_R1146_U160;
  assign new_P2_R1146_U415 = ~new_P2_U3954 | ~new_P2_R1146_U73;
  assign new_P2_R1146_U416 = ~new_P2_U3068 | ~new_P2_R1146_U70;
  assign new_P2_R1146_U417 = ~new_P2_R1146_U416 | ~new_P2_R1146_U415;
  assign new_P2_R1146_U418 = ~new_P2_U3955 | ~new_P2_R1146_U74;
  assign new_P2_R1146_U419 = ~new_P2_U3063 | ~new_P2_R1146_U71;
  assign new_P2_R1146_U420 = ~new_P2_R1146_U327 | ~new_P2_R1146_U89;
  assign new_P2_R1146_U421 = ~new_P2_R1146_U161 | ~new_P2_R1146_U319;
  assign new_P2_R1146_U422 = ~new_P2_U3956 | ~new_P2_R1146_U75;
  assign new_P2_R1146_U423 = ~new_P2_U3077 | ~new_P2_R1146_U72;
  assign new_P2_R1146_U424 = ~new_P2_R1146_U328 | ~new_P2_R1146_U163;
  assign new_P2_R1146_U425 = ~new_P2_R1146_U281 | ~new_P2_R1146_U162;
  assign new_P2_R1146_U426 = ~new_P2_U3957 | ~new_P2_R1146_U69;
  assign new_P2_R1146_U427 = ~new_P2_U3078 | ~new_P2_R1146_U68;
  assign new_P2_R1146_U428 = ~new_P2_R1146_U138;
  assign new_P2_R1146_U429 = ~new_P2_R1146_U277 | ~new_P2_R1146_U428;
  assign new_P2_R1146_U430 = ~new_P2_R1146_U138 | ~new_P2_R1146_U164;
  assign new_P2_R1146_U431 = ~new_P2_U3432 | ~new_P2_R1146_U25;
  assign new_P2_R1146_U432 = ~new_P2_U3080 | ~new_P2_R1146_U165;
  assign new_P2_R1146_U433 = ~new_P2_R1146_U139;
  assign new_P2_R1146_U434 = ~new_P2_R1146_U191 | ~new_P2_R1146_U433;
  assign new_P2_R1146_U435 = ~new_P2_R1146_U139 | ~new_P2_R1146_U166;
  assign new_P2_R1146_U436 = ~new_P2_U3485 | ~new_P2_R1146_U67;
  assign new_P2_R1146_U437 = ~new_P2_U3083 | ~new_P2_R1146_U66;
  assign new_P2_R1146_U438 = ~new_P2_R1146_U140;
  assign new_P2_R1146_U439 = ~new_P2_R1146_U273 | ~new_P2_R1146_U438;
  assign new_P2_R1146_U440 = ~new_P2_R1146_U140 | ~new_P2_R1146_U167;
  assign new_P2_R1146_U441 = ~new_P2_U3483 | ~new_P2_R1146_U65;
  assign new_P2_R1146_U442 = ~new_P2_U3084 | ~new_P2_R1146_U168;
  assign new_P2_R1146_U443 = ~new_P2_R1146_U141;
  assign new_P2_R1146_U444 = ~new_P2_R1146_U443 | ~new_P2_R1146_U269;
  assign new_P2_R1146_U445 = ~new_P2_R1146_U141 | ~new_P2_R1146_U64;
  assign new_P2_R1146_U446 = ~new_P2_U3480 | ~new_P2_R1146_U63;
  assign new_P2_R1146_U447 = ~new_P2_U3071 | ~new_P2_R1146_U62;
  assign new_P2_R1146_U448 = ~new_P2_R1146_U142;
  assign new_P2_R1146_U449 = ~new_P2_R1146_U265 | ~new_P2_R1146_U448;
  assign new_P2_R1146_U450 = ~new_P2_R1146_U142 | ~new_P2_R1146_U169;
  assign new_P2_R1146_U451 = ~new_P2_U3477 | ~new_P2_R1146_U58;
  assign new_P2_R1146_U452 = ~new_P2_U3075 | ~new_P2_R1146_U55;
  assign new_P2_R1146_U453 = ~new_P2_R1146_U452 | ~new_P2_R1146_U451;
  assign new_P2_R1146_U454 = ~new_P2_U3474 | ~new_P2_R1146_U59;
  assign new_P2_R1146_U455 = ~new_P2_U3076 | ~new_P2_R1146_U56;
  assign new_P2_R1146_U456 = ~new_P2_R1146_U338 | ~new_P2_R1146_U90;
  assign new_P2_R1146_U457 = ~new_P2_R1146_U170 | ~new_P2_R1146_U330;
  assign new_P2_R1146_U458 = ~new_P2_U3471 | ~new_P2_R1146_U60;
  assign new_P2_R1146_U459 = ~new_P2_U3081 | ~new_P2_R1146_U57;
  assign new_P2_R1146_U460 = ~new_P2_R1146_U339 | ~new_P2_R1146_U172;
  assign new_P2_R1146_U461 = ~new_P2_R1146_U255 | ~new_P2_R1146_U171;
  assign new_P2_R1146_U462 = ~new_P2_U3468 | ~new_P2_R1146_U54;
  assign new_P2_R1146_U463 = ~new_P2_U3082 | ~new_P2_R1146_U53;
  assign new_P2_R1146_U464 = ~new_P2_R1146_U145;
  assign new_P2_R1146_U465 = ~new_P2_R1146_U251 | ~new_P2_R1146_U464;
  assign new_P2_R1146_U466 = ~new_P2_R1146_U145 | ~new_P2_R1146_U173;
  assign new_P2_R1146_U467 = ~new_P2_U3465 | ~new_P2_R1146_U52;
  assign new_P2_R1146_U468 = ~new_P2_U3074 | ~new_P2_R1146_U51;
  assign new_P2_R1146_U469 = ~new_P2_R1146_U146;
  assign new_P2_R1146_U470 = ~new_P2_R1146_U247 | ~new_P2_R1146_U469;
  assign new_P2_R1146_U471 = ~new_P2_R1146_U146 | ~new_P2_R1146_U174;
  assign new_P2_R1146_U472 = ~new_P2_U3462 | ~new_P2_R1146_U48;
  assign new_P2_R1146_U473 = ~new_P2_U3065 | ~new_P2_R1146_U47;
  assign new_P2_R1146_U474 = ~new_P2_R1146_U473 | ~new_P2_R1146_U472;
  assign new_P2_R1146_U475 = ~new_P2_U3459 | ~new_P2_R1146_U49;
  assign new_P2_R1146_U476 = ~new_P2_U3064 | ~new_P2_R1146_U46;
  assign new_P2_R1146_U477 = ~new_P2_R1146_U349 | ~new_P2_R1146_U91;
  assign new_P2_R1146_U478 = ~new_P2_R1146_U175 | ~new_P2_R1146_U341;
  assign new_P2_R1203_U6 = new_P2_R1203_U202 & new_P2_R1203_U201;
  assign new_P2_R1203_U7 = new_P2_R1203_U241 & new_P2_R1203_U240;
  assign new_P2_R1203_U8 = new_P2_R1203_U181 & new_P2_R1203_U256;
  assign new_P2_R1203_U9 = new_P2_R1203_U258 & new_P2_R1203_U257;
  assign new_P2_R1203_U10 = new_P2_R1203_U182 & new_P2_R1203_U282;
  assign new_P2_R1203_U11 = new_P2_R1203_U284 & new_P2_R1203_U283;
  assign new_P2_R1203_U12 = ~new_P2_R1203_U344 | ~new_P2_R1203_U347;
  assign new_P2_R1203_U13 = ~new_P2_R1203_U333 | ~new_P2_R1203_U336;
  assign new_P2_R1203_U14 = ~new_P2_R1203_U322 | ~new_P2_R1203_U325;
  assign new_P2_R1203_U15 = ~new_P2_R1203_U314 | ~new_P2_R1203_U316;
  assign new_P2_R1203_U16 = ~new_P2_R1203_U352 | ~new_P2_R1203_U312;
  assign new_P2_R1203_U17 = ~new_P2_R1203_U235 | ~new_P2_R1203_U237;
  assign new_P2_R1203_U18 = ~new_P2_R1203_U227 | ~new_P2_R1203_U230;
  assign new_P2_R1203_U19 = ~new_P2_R1203_U219 | ~new_P2_R1203_U221;
  assign new_P2_R1203_U20 = ~new_P2_R1203_U166 | ~new_P2_R1203_U350;
  assign new_P2_R1203_U21 = ~new_P2_U3450;
  assign new_P2_R1203_U22 = ~new_P2_U3444;
  assign new_P2_R1203_U23 = ~new_P2_U3435;
  assign new_P2_R1203_U24 = ~new_P2_U3427;
  assign new_P2_R1203_U25 = ~new_P2_U3080;
  assign new_P2_R1203_U26 = ~new_P2_U3438;
  assign new_P2_R1203_U27 = ~new_P2_U3070;
  assign new_P2_R1203_U28 = ~new_P2_U3070 | ~new_P2_R1203_U23;
  assign new_P2_R1203_U29 = ~new_P2_U3066;
  assign new_P2_R1203_U30 = ~new_P2_U3447;
  assign new_P2_R1203_U31 = ~new_P2_U3441;
  assign new_P2_R1203_U32 = ~new_P2_U3073;
  assign new_P2_R1203_U33 = ~new_P2_U3069;
  assign new_P2_R1203_U34 = ~new_P2_U3062;
  assign new_P2_R1203_U35 = ~new_P2_U3062 | ~new_P2_R1203_U31;
  assign new_P2_R1203_U36 = ~new_P2_U3453;
  assign new_P2_R1203_U37 = ~new_P2_U3072;
  assign new_P2_R1203_U38 = ~new_P2_U3072 | ~new_P2_R1203_U21;
  assign new_P2_R1203_U39 = ~new_P2_U3086;
  assign new_P2_R1203_U40 = ~new_P2_U3456;
  assign new_P2_R1203_U41 = ~new_P2_U3085;
  assign new_P2_R1203_U42 = ~new_P2_R1203_U208 | ~new_P2_R1203_U207;
  assign new_P2_R1203_U43 = ~new_P2_R1203_U35 | ~new_P2_R1203_U223;
  assign new_P2_R1203_U44 = ~new_P2_R1203_U351 | ~new_P2_R1203_U192 | ~new_P2_R1203_U176;
  assign new_P2_R1203_U45 = ~new_P2_U3951;
  assign new_P2_R1203_U46 = ~new_P2_U3459;
  assign new_P2_R1203_U47 = ~new_P2_U3462;
  assign new_P2_R1203_U48 = ~new_P2_U3065;
  assign new_P2_R1203_U49 = ~new_P2_U3064;
  assign new_P2_R1203_U50 = ~new_P2_U3085 | ~new_P2_R1203_U40;
  assign new_P2_R1203_U51 = ~new_P2_U3465;
  assign new_P2_R1203_U52 = ~new_P2_U3074;
  assign new_P2_R1203_U53 = ~new_P2_U3468;
  assign new_P2_R1203_U54 = ~new_P2_U3082;
  assign new_P2_R1203_U55 = ~new_P2_U3477;
  assign new_P2_R1203_U56 = ~new_P2_U3474;
  assign new_P2_R1203_U57 = ~new_P2_U3471;
  assign new_P2_R1203_U58 = ~new_P2_U3075;
  assign new_P2_R1203_U59 = ~new_P2_U3076;
  assign new_P2_R1203_U60 = ~new_P2_U3081;
  assign new_P2_R1203_U61 = ~new_P2_U3081 | ~new_P2_R1203_U57;
  assign new_P2_R1203_U62 = ~new_P2_U3480;
  assign new_P2_R1203_U63 = ~new_P2_U3071;
  assign new_P2_R1203_U64 = ~new_P2_R1203_U268 | ~new_P2_R1203_U267;
  assign new_P2_R1203_U65 = ~new_P2_U3084;
  assign new_P2_R1203_U66 = ~new_P2_U3485;
  assign new_P2_R1203_U67 = ~new_P2_U3083;
  assign new_P2_R1203_U68 = ~new_P2_U3957;
  assign new_P2_R1203_U69 = ~new_P2_U3078;
  assign new_P2_R1203_U70 = ~new_P2_U3954;
  assign new_P2_R1203_U71 = ~new_P2_U3955;
  assign new_P2_R1203_U72 = ~new_P2_U3956;
  assign new_P2_R1203_U73 = ~new_P2_U3068;
  assign new_P2_R1203_U74 = ~new_P2_U3063;
  assign new_P2_R1203_U75 = ~new_P2_U3077;
  assign new_P2_R1203_U76 = ~new_P2_U3077 | ~new_P2_R1203_U72;
  assign new_P2_R1203_U77 = ~new_P2_U3953;
  assign new_P2_R1203_U78 = ~new_P2_U3067;
  assign new_P2_R1203_U79 = ~new_P2_U3952;
  assign new_P2_R1203_U80 = ~new_P2_U3060;
  assign new_P2_R1203_U81 = ~new_P2_U3950;
  assign new_P2_R1203_U82 = ~new_P2_U3059;
  assign new_P2_R1203_U83 = ~new_P2_U3059 | ~new_P2_R1203_U45;
  assign new_P2_R1203_U84 = ~new_P2_U3055;
  assign new_P2_R1203_U85 = ~new_P2_U3949;
  assign new_P2_R1203_U86 = ~new_P2_U3056;
  assign new_P2_R1203_U87 = ~new_P2_R1203_U128 | ~new_P2_R1203_U301;
  assign new_P2_R1203_U88 = ~new_P2_R1203_U298 | ~new_P2_R1203_U297;
  assign new_P2_R1203_U89 = ~new_P2_R1203_U76 | ~new_P2_R1203_U318;
  assign new_P2_R1203_U90 = ~new_P2_R1203_U61 | ~new_P2_R1203_U329;
  assign new_P2_R1203_U91 = ~new_P2_R1203_U50 | ~new_P2_R1203_U340;
  assign new_P2_R1203_U92 = ~new_P2_U3079;
  assign new_P2_R1203_U93 = ~new_P2_R1203_U395 | ~new_P2_R1203_U394;
  assign new_P2_R1203_U94 = ~new_P2_R1203_U409 | ~new_P2_R1203_U408;
  assign new_P2_R1203_U95 = ~new_P2_R1203_U414 | ~new_P2_R1203_U413;
  assign new_P2_R1203_U96 = ~new_P2_R1203_U430 | ~new_P2_R1203_U429;
  assign new_P2_R1203_U97 = ~new_P2_R1203_U435 | ~new_P2_R1203_U434;
  assign new_P2_R1203_U98 = ~new_P2_R1203_U440 | ~new_P2_R1203_U439;
  assign new_P2_R1203_U99 = ~new_P2_R1203_U445 | ~new_P2_R1203_U444;
  assign new_P2_R1203_U100 = ~new_P2_R1203_U450 | ~new_P2_R1203_U449;
  assign new_P2_R1203_U101 = ~new_P2_R1203_U466 | ~new_P2_R1203_U465;
  assign new_P2_R1203_U102 = ~new_P2_R1203_U471 | ~new_P2_R1203_U470;
  assign new_P2_R1203_U103 = ~new_P2_R1203_U356 | ~new_P2_R1203_U355;
  assign new_P2_R1203_U104 = ~new_P2_R1203_U365 | ~new_P2_R1203_U364;
  assign new_P2_R1203_U105 = ~new_P2_R1203_U372 | ~new_P2_R1203_U371;
  assign new_P2_R1203_U106 = ~new_P2_R1203_U376 | ~new_P2_R1203_U375;
  assign new_P2_R1203_U107 = ~new_P2_R1203_U385 | ~new_P2_R1203_U384;
  assign new_P2_R1203_U108 = ~new_P2_R1203_U404 | ~new_P2_R1203_U403;
  assign new_P2_R1203_U109 = ~new_P2_R1203_U421 | ~new_P2_R1203_U420;
  assign new_P2_R1203_U110 = ~new_P2_R1203_U425 | ~new_P2_R1203_U424;
  assign new_P2_R1203_U111 = ~new_P2_R1203_U457 | ~new_P2_R1203_U456;
  assign new_P2_R1203_U112 = ~new_P2_R1203_U461 | ~new_P2_R1203_U460;
  assign new_P2_R1203_U113 = ~new_P2_R1203_U478 | ~new_P2_R1203_U477;
  assign new_P2_R1203_U114 = new_P2_R1203_U194 & new_P2_R1203_U184;
  assign new_P2_R1203_U115 = new_P2_R1203_U197 & new_P2_R1203_U198;
  assign new_P2_R1203_U116 = new_P2_R1203_U185 & new_P2_R1203_U205 & new_P2_R1203_U200;
  assign new_P2_R1203_U117 = new_P2_R1203_U210 & new_P2_R1203_U186;
  assign new_P2_R1203_U118 = new_P2_R1203_U213 & new_P2_R1203_U214;
  assign new_P2_R1203_U119 = new_P2_R1203_U38 & new_P2_R1203_U358 & new_P2_R1203_U357;
  assign new_P2_R1203_U120 = new_P2_R1203_U361 & new_P2_R1203_U186;
  assign new_P2_R1203_U121 = new_P2_R1203_U229 & new_P2_R1203_U6;
  assign new_P2_R1203_U122 = new_P2_R1203_U368 & new_P2_R1203_U185;
  assign new_P2_R1203_U123 = new_P2_R1203_U28 & new_P2_R1203_U378 & new_P2_R1203_U377;
  assign new_P2_R1203_U124 = new_P2_R1203_U381 & new_P2_R1203_U184;
  assign new_P2_R1203_U125 = new_P2_R1203_U180 & new_P2_R1203_U239 & new_P2_R1203_U216;
  assign new_P2_R1203_U126 = new_P2_R1203_U261 & new_P2_R1203_U8;
  assign new_P2_R1203_U127 = new_P2_R1203_U287 & new_P2_R1203_U10;
  assign new_P2_R1203_U128 = new_P2_R1203_U303 & new_P2_R1203_U304;
  assign new_P2_R1203_U129 = new_P2_R1203_U311 & new_P2_R1203_U387 & new_P2_R1203_U386;
  assign new_P2_R1203_U130 = new_P2_R1203_U308 & new_P2_R1203_U390;
  assign new_P2_R1203_U131 = ~new_P2_R1203_U392 | ~new_P2_R1203_U391;
  assign new_P2_R1203_U132 = new_P2_R1203_U83 & new_P2_R1203_U397 & new_P2_R1203_U396;
  assign new_P2_R1203_U133 = new_P2_R1203_U400 & new_P2_R1203_U183;
  assign new_P2_R1203_U134 = ~new_P2_R1203_U406 | ~new_P2_R1203_U405;
  assign new_P2_R1203_U135 = ~new_P2_R1203_U411 | ~new_P2_R1203_U410;
  assign new_P2_R1203_U136 = new_P2_R1203_U324 & new_P2_R1203_U11;
  assign new_P2_R1203_U137 = new_P2_R1203_U417 & new_P2_R1203_U182;
  assign new_P2_R1203_U138 = ~new_P2_R1203_U427 | ~new_P2_R1203_U426;
  assign new_P2_R1203_U139 = ~new_P2_R1203_U432 | ~new_P2_R1203_U431;
  assign new_P2_R1203_U140 = ~new_P2_R1203_U437 | ~new_P2_R1203_U436;
  assign new_P2_R1203_U141 = ~new_P2_R1203_U442 | ~new_P2_R1203_U441;
  assign new_P2_R1203_U142 = ~new_P2_R1203_U447 | ~new_P2_R1203_U446;
  assign new_P2_R1203_U143 = new_P2_R1203_U335 & new_P2_R1203_U9;
  assign new_P2_R1203_U144 = new_P2_R1203_U453 & new_P2_R1203_U181;
  assign new_P2_R1203_U145 = ~new_P2_R1203_U463 | ~new_P2_R1203_U462;
  assign new_P2_R1203_U146 = ~new_P2_R1203_U468 | ~new_P2_R1203_U467;
  assign new_P2_R1203_U147 = new_P2_R1203_U346 & new_P2_R1203_U7;
  assign new_P2_R1203_U148 = new_P2_R1203_U474 & new_P2_R1203_U180;
  assign new_P2_R1203_U149 = new_P2_R1203_U354 & new_P2_R1203_U353;
  assign new_P2_R1203_U150 = ~new_P2_R1203_U118 | ~new_P2_R1203_U211;
  assign new_P2_R1203_U151 = new_P2_R1203_U363 & new_P2_R1203_U362;
  assign new_P2_R1203_U152 = new_P2_R1203_U370 & new_P2_R1203_U369;
  assign new_P2_R1203_U153 = new_P2_R1203_U374 & new_P2_R1203_U373;
  assign new_P2_R1203_U154 = ~new_P2_R1203_U115 | ~new_P2_R1203_U195;
  assign new_P2_R1203_U155 = new_P2_R1203_U383 & new_P2_R1203_U382;
  assign new_P2_R1203_U156 = ~new_P2_U3960;
  assign new_P2_R1203_U157 = ~new_P2_U3057;
  assign new_P2_R1203_U158 = new_P2_R1203_U402 & new_P2_R1203_U401;
  assign new_P2_R1203_U159 = ~new_P2_R1203_U294 | ~new_P2_R1203_U293;
  assign new_P2_R1203_U160 = ~new_P2_R1203_U290 | ~new_P2_R1203_U289;
  assign new_P2_R1203_U161 = new_P2_R1203_U419 & new_P2_R1203_U418;
  assign new_P2_R1203_U162 = new_P2_R1203_U423 & new_P2_R1203_U422;
  assign new_P2_R1203_U163 = ~new_P2_R1203_U280 | ~new_P2_R1203_U279;
  assign new_P2_R1203_U164 = ~new_P2_R1203_U276 | ~new_P2_R1203_U275;
  assign new_P2_R1203_U165 = ~new_P2_U3432;
  assign new_P2_R1203_U166 = ~new_P2_U3427 | ~new_P2_R1203_U92;
  assign new_P2_R1203_U167 = ~new_P2_R1203_U272 | ~new_P2_R1203_U271;
  assign new_P2_R1203_U168 = ~new_P2_U3483;
  assign new_P2_R1203_U169 = ~new_P2_R1203_U264 | ~new_P2_R1203_U263;
  assign new_P2_R1203_U170 = new_P2_R1203_U455 & new_P2_R1203_U454;
  assign new_P2_R1203_U171 = new_P2_R1203_U459 & new_P2_R1203_U458;
  assign new_P2_R1203_U172 = ~new_P2_R1203_U254 | ~new_P2_R1203_U253;
  assign new_P2_R1203_U173 = ~new_P2_R1203_U250 | ~new_P2_R1203_U249;
  assign new_P2_R1203_U174 = ~new_P2_R1203_U246 | ~new_P2_R1203_U245;
  assign new_P2_R1203_U175 = new_P2_R1203_U476 & new_P2_R1203_U475;
  assign new_P2_R1203_U176 = ~new_P2_R1203_U166 | ~new_P2_R1203_U165;
  assign new_P2_R1203_U177 = ~new_P2_R1203_U83;
  assign new_P2_R1203_U178 = ~new_P2_R1203_U28;
  assign new_P2_R1203_U179 = ~new_P2_R1203_U38;
  assign new_P2_R1203_U180 = ~new_P2_U3459 | ~new_P2_R1203_U49;
  assign new_P2_R1203_U181 = ~new_P2_U3474 | ~new_P2_R1203_U59;
  assign new_P2_R1203_U182 = ~new_P2_U3955 | ~new_P2_R1203_U74;
  assign new_P2_R1203_U183 = ~new_P2_U3951 | ~new_P2_R1203_U82;
  assign new_P2_R1203_U184 = ~new_P2_U3435 | ~new_P2_R1203_U27;
  assign new_P2_R1203_U185 = ~new_P2_U3444 | ~new_P2_R1203_U33;
  assign new_P2_R1203_U186 = ~new_P2_U3450 | ~new_P2_R1203_U37;
  assign new_P2_R1203_U187 = ~new_P2_R1203_U61;
  assign new_P2_R1203_U188 = ~new_P2_R1203_U76;
  assign new_P2_R1203_U189 = ~new_P2_R1203_U35;
  assign new_P2_R1203_U190 = ~new_P2_R1203_U50;
  assign new_P2_R1203_U191 = ~new_P2_R1203_U166;
  assign new_P2_R1203_U192 = ~new_P2_U3080 | ~new_P2_R1203_U166;
  assign new_P2_R1203_U193 = ~new_P2_R1203_U44;
  assign new_P2_R1203_U194 = ~new_P2_U3438 | ~new_P2_R1203_U29;
  assign new_P2_R1203_U195 = ~new_P2_R1203_U114 | ~new_P2_R1203_U44;
  assign new_P2_R1203_U196 = ~new_P2_R1203_U29 | ~new_P2_R1203_U28;
  assign new_P2_R1203_U197 = ~new_P2_R1203_U196 | ~new_P2_R1203_U26;
  assign new_P2_R1203_U198 = ~new_P2_U3066 | ~new_P2_R1203_U178;
  assign new_P2_R1203_U199 = ~new_P2_R1203_U154;
  assign new_P2_R1203_U200 = ~new_P2_U3447 | ~new_P2_R1203_U32;
  assign new_P2_R1203_U201 = ~new_P2_U3073 | ~new_P2_R1203_U30;
  assign new_P2_R1203_U202 = ~new_P2_U3069 | ~new_P2_R1203_U22;
  assign new_P2_R1203_U203 = ~new_P2_R1203_U189 | ~new_P2_R1203_U185;
  assign new_P2_R1203_U204 = ~new_P2_R1203_U6 | ~new_P2_R1203_U203;
  assign new_P2_R1203_U205 = ~new_P2_U3441 | ~new_P2_R1203_U34;
  assign new_P2_R1203_U206 = ~new_P2_U3447 | ~new_P2_R1203_U32;
  assign new_P2_R1203_U207 = ~new_P2_R1203_U154 | ~new_P2_R1203_U116;
  assign new_P2_R1203_U208 = ~new_P2_R1203_U206 | ~new_P2_R1203_U204;
  assign new_P2_R1203_U209 = ~new_P2_R1203_U42;
  assign new_P2_R1203_U210 = ~new_P2_U3453 | ~new_P2_R1203_U39;
  assign new_P2_R1203_U211 = ~new_P2_R1203_U117 | ~new_P2_R1203_U42;
  assign new_P2_R1203_U212 = ~new_P2_R1203_U39 | ~new_P2_R1203_U38;
  assign new_P2_R1203_U213 = ~new_P2_R1203_U212 | ~new_P2_R1203_U36;
  assign new_P2_R1203_U214 = ~new_P2_U3086 | ~new_P2_R1203_U179;
  assign new_P2_R1203_U215 = ~new_P2_R1203_U150;
  assign new_P2_R1203_U216 = ~new_P2_U3456 | ~new_P2_R1203_U41;
  assign new_P2_R1203_U217 = ~new_P2_R1203_U216 | ~new_P2_R1203_U50;
  assign new_P2_R1203_U218 = ~new_P2_R1203_U209 | ~new_P2_R1203_U38;
  assign new_P2_R1203_U219 = ~new_P2_R1203_U120 | ~new_P2_R1203_U218;
  assign new_P2_R1203_U220 = ~new_P2_R1203_U42 | ~new_P2_R1203_U186;
  assign new_P2_R1203_U221 = ~new_P2_R1203_U119 | ~new_P2_R1203_U220;
  assign new_P2_R1203_U222 = ~new_P2_R1203_U38 | ~new_P2_R1203_U186;
  assign new_P2_R1203_U223 = ~new_P2_R1203_U205 | ~new_P2_R1203_U154;
  assign new_P2_R1203_U224 = ~new_P2_R1203_U43;
  assign new_P2_R1203_U225 = ~new_P2_U3069 | ~new_P2_R1203_U22;
  assign new_P2_R1203_U226 = ~new_P2_R1203_U224 | ~new_P2_R1203_U225;
  assign new_P2_R1203_U227 = ~new_P2_R1203_U122 | ~new_P2_R1203_U226;
  assign new_P2_R1203_U228 = ~new_P2_R1203_U43 | ~new_P2_R1203_U185;
  assign new_P2_R1203_U229 = ~new_P2_U3447 | ~new_P2_R1203_U32;
  assign new_P2_R1203_U230 = ~new_P2_R1203_U121 | ~new_P2_R1203_U228;
  assign new_P2_R1203_U231 = ~new_P2_U3069 | ~new_P2_R1203_U22;
  assign new_P2_R1203_U232 = ~new_P2_R1203_U185 | ~new_P2_R1203_U231;
  assign new_P2_R1203_U233 = ~new_P2_R1203_U205 | ~new_P2_R1203_U35;
  assign new_P2_R1203_U234 = ~new_P2_R1203_U193 | ~new_P2_R1203_U28;
  assign new_P2_R1203_U235 = ~new_P2_R1203_U124 | ~new_P2_R1203_U234;
  assign new_P2_R1203_U236 = ~new_P2_R1203_U44 | ~new_P2_R1203_U184;
  assign new_P2_R1203_U237 = ~new_P2_R1203_U123 | ~new_P2_R1203_U236;
  assign new_P2_R1203_U238 = ~new_P2_R1203_U28 | ~new_P2_R1203_U184;
  assign new_P2_R1203_U239 = ~new_P2_U3462 | ~new_P2_R1203_U48;
  assign new_P2_R1203_U240 = ~new_P2_U3065 | ~new_P2_R1203_U47;
  assign new_P2_R1203_U241 = ~new_P2_U3064 | ~new_P2_R1203_U46;
  assign new_P2_R1203_U242 = ~new_P2_R1203_U190 | ~new_P2_R1203_U180;
  assign new_P2_R1203_U243 = ~new_P2_R1203_U7 | ~new_P2_R1203_U242;
  assign new_P2_R1203_U244 = ~new_P2_U3462 | ~new_P2_R1203_U48;
  assign new_P2_R1203_U245 = ~new_P2_R1203_U150 | ~new_P2_R1203_U125;
  assign new_P2_R1203_U246 = ~new_P2_R1203_U244 | ~new_P2_R1203_U243;
  assign new_P2_R1203_U247 = ~new_P2_R1203_U174;
  assign new_P2_R1203_U248 = ~new_P2_U3465 | ~new_P2_R1203_U52;
  assign new_P2_R1203_U249 = ~new_P2_R1203_U248 | ~new_P2_R1203_U174;
  assign new_P2_R1203_U250 = ~new_P2_U3074 | ~new_P2_R1203_U51;
  assign new_P2_R1203_U251 = ~new_P2_R1203_U173;
  assign new_P2_R1203_U252 = ~new_P2_U3468 | ~new_P2_R1203_U54;
  assign new_P2_R1203_U253 = ~new_P2_R1203_U252 | ~new_P2_R1203_U173;
  assign new_P2_R1203_U254 = ~new_P2_U3082 | ~new_P2_R1203_U53;
  assign new_P2_R1203_U255 = ~new_P2_R1203_U172;
  assign new_P2_R1203_U256 = ~new_P2_U3477 | ~new_P2_R1203_U58;
  assign new_P2_R1203_U257 = ~new_P2_U3075 | ~new_P2_R1203_U55;
  assign new_P2_R1203_U258 = ~new_P2_U3076 | ~new_P2_R1203_U56;
  assign new_P2_R1203_U259 = ~new_P2_R1203_U187 | ~new_P2_R1203_U8;
  assign new_P2_R1203_U260 = ~new_P2_R1203_U9 | ~new_P2_R1203_U259;
  assign new_P2_R1203_U261 = ~new_P2_U3471 | ~new_P2_R1203_U60;
  assign new_P2_R1203_U262 = ~new_P2_U3477 | ~new_P2_R1203_U58;
  assign new_P2_R1203_U263 = ~new_P2_R1203_U126 | ~new_P2_R1203_U172;
  assign new_P2_R1203_U264 = ~new_P2_R1203_U262 | ~new_P2_R1203_U260;
  assign new_P2_R1203_U265 = ~new_P2_R1203_U169;
  assign new_P2_R1203_U266 = ~new_P2_U3480 | ~new_P2_R1203_U63;
  assign new_P2_R1203_U267 = ~new_P2_R1203_U266 | ~new_P2_R1203_U169;
  assign new_P2_R1203_U268 = ~new_P2_U3071 | ~new_P2_R1203_U62;
  assign new_P2_R1203_U269 = ~new_P2_R1203_U64;
  assign new_P2_R1203_U270 = ~new_P2_R1203_U269 | ~new_P2_R1203_U65;
  assign new_P2_R1203_U271 = ~new_P2_R1203_U270 | ~new_P2_R1203_U168;
  assign new_P2_R1203_U272 = ~new_P2_U3084 | ~new_P2_R1203_U64;
  assign new_P2_R1203_U273 = ~new_P2_R1203_U167;
  assign new_P2_R1203_U274 = ~new_P2_U3485 | ~new_P2_R1203_U67;
  assign new_P2_R1203_U275 = ~new_P2_R1203_U274 | ~new_P2_R1203_U167;
  assign new_P2_R1203_U276 = ~new_P2_U3083 | ~new_P2_R1203_U66;
  assign new_P2_R1203_U277 = ~new_P2_R1203_U164;
  assign new_P2_R1203_U278 = ~new_P2_U3957 | ~new_P2_R1203_U69;
  assign new_P2_R1203_U279 = ~new_P2_R1203_U278 | ~new_P2_R1203_U164;
  assign new_P2_R1203_U280 = ~new_P2_U3078 | ~new_P2_R1203_U68;
  assign new_P2_R1203_U281 = ~new_P2_R1203_U163;
  assign new_P2_R1203_U282 = ~new_P2_U3954 | ~new_P2_R1203_U73;
  assign new_P2_R1203_U283 = ~new_P2_U3068 | ~new_P2_R1203_U70;
  assign new_P2_R1203_U284 = ~new_P2_U3063 | ~new_P2_R1203_U71;
  assign new_P2_R1203_U285 = ~new_P2_R1203_U188 | ~new_P2_R1203_U10;
  assign new_P2_R1203_U286 = ~new_P2_R1203_U11 | ~new_P2_R1203_U285;
  assign new_P2_R1203_U287 = ~new_P2_U3956 | ~new_P2_R1203_U75;
  assign new_P2_R1203_U288 = ~new_P2_U3954 | ~new_P2_R1203_U73;
  assign new_P2_R1203_U289 = ~new_P2_R1203_U127 | ~new_P2_R1203_U163;
  assign new_P2_R1203_U290 = ~new_P2_R1203_U288 | ~new_P2_R1203_U286;
  assign new_P2_R1203_U291 = ~new_P2_R1203_U160;
  assign new_P2_R1203_U292 = ~new_P2_U3953 | ~new_P2_R1203_U78;
  assign new_P2_R1203_U293 = ~new_P2_R1203_U292 | ~new_P2_R1203_U160;
  assign new_P2_R1203_U294 = ~new_P2_U3067 | ~new_P2_R1203_U77;
  assign new_P2_R1203_U295 = ~new_P2_R1203_U159;
  assign new_P2_R1203_U296 = ~new_P2_U3952 | ~new_P2_R1203_U80;
  assign new_P2_R1203_U297 = ~new_P2_R1203_U296 | ~new_P2_R1203_U159;
  assign new_P2_R1203_U298 = ~new_P2_U3060 | ~new_P2_R1203_U79;
  assign new_P2_R1203_U299 = ~new_P2_R1203_U88;
  assign new_P2_R1203_U300 = ~new_P2_U3950 | ~new_P2_R1203_U84;
  assign new_P2_R1203_U301 = ~new_P2_R1203_U300 | ~new_P2_R1203_U88 | ~new_P2_R1203_U183;
  assign new_P2_R1203_U302 = ~new_P2_R1203_U84 | ~new_P2_R1203_U83;
  assign new_P2_R1203_U303 = ~new_P2_R1203_U302 | ~new_P2_R1203_U81;
  assign new_P2_R1203_U304 = ~new_P2_U3055 | ~new_P2_R1203_U177;
  assign new_P2_R1203_U305 = ~new_P2_R1203_U87;
  assign new_P2_R1203_U306 = ~new_P2_U3056 | ~new_P2_R1203_U85;
  assign new_P2_R1203_U307 = ~new_P2_R1203_U305 | ~new_P2_R1203_U306;
  assign new_P2_R1203_U308 = ~new_P2_U3949 | ~new_P2_R1203_U86;
  assign new_P2_R1203_U309 = ~new_P2_U3949 | ~new_P2_R1203_U86;
  assign new_P2_R1203_U310 = ~new_P2_R1203_U309 | ~new_P2_R1203_U87;
  assign new_P2_R1203_U311 = ~new_P2_U3056 | ~new_P2_R1203_U85;
  assign new_P2_R1203_U312 = ~new_P2_R1203_U129 | ~new_P2_R1203_U310;
  assign new_P2_R1203_U313 = ~new_P2_R1203_U299 | ~new_P2_R1203_U83;
  assign new_P2_R1203_U314 = ~new_P2_R1203_U133 | ~new_P2_R1203_U313;
  assign new_P2_R1203_U315 = ~new_P2_R1203_U88 | ~new_P2_R1203_U183;
  assign new_P2_R1203_U316 = ~new_P2_R1203_U132 | ~new_P2_R1203_U315;
  assign new_P2_R1203_U317 = ~new_P2_R1203_U83 | ~new_P2_R1203_U183;
  assign new_P2_R1203_U318 = ~new_P2_R1203_U287 | ~new_P2_R1203_U163;
  assign new_P2_R1203_U319 = ~new_P2_R1203_U89;
  assign new_P2_R1203_U320 = ~new_P2_U3063 | ~new_P2_R1203_U71;
  assign new_P2_R1203_U321 = ~new_P2_R1203_U319 | ~new_P2_R1203_U320;
  assign new_P2_R1203_U322 = ~new_P2_R1203_U137 | ~new_P2_R1203_U321;
  assign new_P2_R1203_U323 = ~new_P2_R1203_U89 | ~new_P2_R1203_U182;
  assign new_P2_R1203_U324 = ~new_P2_U3954 | ~new_P2_R1203_U73;
  assign new_P2_R1203_U325 = ~new_P2_R1203_U136 | ~new_P2_R1203_U323;
  assign new_P2_R1203_U326 = ~new_P2_U3063 | ~new_P2_R1203_U71;
  assign new_P2_R1203_U327 = ~new_P2_R1203_U182 | ~new_P2_R1203_U326;
  assign new_P2_R1203_U328 = ~new_P2_R1203_U287 | ~new_P2_R1203_U76;
  assign new_P2_R1203_U329 = ~new_P2_R1203_U261 | ~new_P2_R1203_U172;
  assign new_P2_R1203_U330 = ~new_P2_R1203_U90;
  assign new_P2_R1203_U331 = ~new_P2_U3076 | ~new_P2_R1203_U56;
  assign new_P2_R1203_U332 = ~new_P2_R1203_U330 | ~new_P2_R1203_U331;
  assign new_P2_R1203_U333 = ~new_P2_R1203_U144 | ~new_P2_R1203_U332;
  assign new_P2_R1203_U334 = ~new_P2_R1203_U90 | ~new_P2_R1203_U181;
  assign new_P2_R1203_U335 = ~new_P2_U3477 | ~new_P2_R1203_U58;
  assign new_P2_R1203_U336 = ~new_P2_R1203_U143 | ~new_P2_R1203_U334;
  assign new_P2_R1203_U337 = ~new_P2_U3076 | ~new_P2_R1203_U56;
  assign new_P2_R1203_U338 = ~new_P2_R1203_U181 | ~new_P2_R1203_U337;
  assign new_P2_R1203_U339 = ~new_P2_R1203_U261 | ~new_P2_R1203_U61;
  assign new_P2_R1203_U340 = ~new_P2_R1203_U216 | ~new_P2_R1203_U150;
  assign new_P2_R1203_U341 = ~new_P2_R1203_U91;
  assign new_P2_R1203_U342 = ~new_P2_U3064 | ~new_P2_R1203_U46;
  assign new_P2_R1203_U343 = ~new_P2_R1203_U341 | ~new_P2_R1203_U342;
  assign new_P2_R1203_U344 = ~new_P2_R1203_U148 | ~new_P2_R1203_U343;
  assign new_P2_R1203_U345 = ~new_P2_R1203_U91 | ~new_P2_R1203_U180;
  assign new_P2_R1203_U346 = ~new_P2_U3462 | ~new_P2_R1203_U48;
  assign new_P2_R1203_U347 = ~new_P2_R1203_U147 | ~new_P2_R1203_U345;
  assign new_P2_R1203_U348 = ~new_P2_U3064 | ~new_P2_R1203_U46;
  assign new_P2_R1203_U349 = ~new_P2_R1203_U180 | ~new_P2_R1203_U348;
  assign new_P2_R1203_U350 = ~new_P2_U3079 | ~new_P2_R1203_U24;
  assign new_P2_R1203_U351 = ~new_P2_U3080 | ~new_P2_R1203_U165;
  assign new_P2_R1203_U352 = ~new_P2_R1203_U130 | ~new_P2_R1203_U307;
  assign new_P2_R1203_U353 = ~new_P2_U3456 | ~new_P2_R1203_U41;
  assign new_P2_R1203_U354 = ~new_P2_U3085 | ~new_P2_R1203_U40;
  assign new_P2_R1203_U355 = ~new_P2_R1203_U217 | ~new_P2_R1203_U150;
  assign new_P2_R1203_U356 = ~new_P2_R1203_U215 | ~new_P2_R1203_U149;
  assign new_P2_R1203_U357 = ~new_P2_U3453 | ~new_P2_R1203_U39;
  assign new_P2_R1203_U358 = ~new_P2_U3086 | ~new_P2_R1203_U36;
  assign new_P2_R1203_U359 = ~new_P2_U3453 | ~new_P2_R1203_U39;
  assign new_P2_R1203_U360 = ~new_P2_U3086 | ~new_P2_R1203_U36;
  assign new_P2_R1203_U361 = ~new_P2_R1203_U360 | ~new_P2_R1203_U359;
  assign new_P2_R1203_U362 = ~new_P2_U3450 | ~new_P2_R1203_U37;
  assign new_P2_R1203_U363 = ~new_P2_U3072 | ~new_P2_R1203_U21;
  assign new_P2_R1203_U364 = ~new_P2_R1203_U222 | ~new_P2_R1203_U42;
  assign new_P2_R1203_U365 = ~new_P2_R1203_U151 | ~new_P2_R1203_U209;
  assign new_P2_R1203_U366 = ~new_P2_U3447 | ~new_P2_R1203_U32;
  assign new_P2_R1203_U367 = ~new_P2_U3073 | ~new_P2_R1203_U30;
  assign new_P2_R1203_U368 = ~new_P2_R1203_U367 | ~new_P2_R1203_U366;
  assign new_P2_R1203_U369 = ~new_P2_U3444 | ~new_P2_R1203_U33;
  assign new_P2_R1203_U370 = ~new_P2_U3069 | ~new_P2_R1203_U22;
  assign new_P2_R1203_U371 = ~new_P2_R1203_U232 | ~new_P2_R1203_U43;
  assign new_P2_R1203_U372 = ~new_P2_R1203_U152 | ~new_P2_R1203_U224;
  assign new_P2_R1203_U373 = ~new_P2_U3441 | ~new_P2_R1203_U34;
  assign new_P2_R1203_U374 = ~new_P2_U3062 | ~new_P2_R1203_U31;
  assign new_P2_R1203_U375 = ~new_P2_R1203_U233 | ~new_P2_R1203_U154;
  assign new_P2_R1203_U376 = ~new_P2_R1203_U199 | ~new_P2_R1203_U153;
  assign new_P2_R1203_U377 = ~new_P2_U3438 | ~new_P2_R1203_U29;
  assign new_P2_R1203_U378 = ~new_P2_U3066 | ~new_P2_R1203_U26;
  assign new_P2_R1203_U379 = ~new_P2_U3438 | ~new_P2_R1203_U29;
  assign new_P2_R1203_U380 = ~new_P2_U3066 | ~new_P2_R1203_U26;
  assign new_P2_R1203_U381 = ~new_P2_R1203_U380 | ~new_P2_R1203_U379;
  assign new_P2_R1203_U382 = ~new_P2_U3435 | ~new_P2_R1203_U27;
  assign new_P2_R1203_U383 = ~new_P2_U3070 | ~new_P2_R1203_U23;
  assign new_P2_R1203_U384 = ~new_P2_R1203_U238 | ~new_P2_R1203_U44;
  assign new_P2_R1203_U385 = ~new_P2_R1203_U155 | ~new_P2_R1203_U193;
  assign new_P2_R1203_U386 = ~new_P2_U3960 | ~new_P2_R1203_U157;
  assign new_P2_R1203_U387 = ~new_P2_U3057 | ~new_P2_R1203_U156;
  assign new_P2_R1203_U388 = ~new_P2_U3960 | ~new_P2_R1203_U157;
  assign new_P2_R1203_U389 = ~new_P2_U3057 | ~new_P2_R1203_U156;
  assign new_P2_R1203_U390 = ~new_P2_R1203_U389 | ~new_P2_R1203_U388;
  assign new_P2_R1203_U391 = ~new_P2_U3949 | ~new_P2_R1203_U86;
  assign new_P2_R1203_U392 = ~new_P2_U3056 | ~new_P2_R1203_U85;
  assign new_P2_R1203_U393 = ~new_P2_R1203_U131;
  assign new_P2_R1203_U394 = ~new_P2_R1203_U393 | ~new_P2_R1203_U305;
  assign new_P2_R1203_U395 = ~new_P2_R1203_U131 | ~new_P2_R1203_U87;
  assign new_P2_R1203_U396 = ~new_P2_U3950 | ~new_P2_R1203_U84;
  assign new_P2_R1203_U397 = ~new_P2_U3055 | ~new_P2_R1203_U81;
  assign new_P2_R1203_U398 = ~new_P2_U3950 | ~new_P2_R1203_U84;
  assign new_P2_R1203_U399 = ~new_P2_U3055 | ~new_P2_R1203_U81;
  assign new_P2_R1203_U400 = ~new_P2_R1203_U399 | ~new_P2_R1203_U398;
  assign new_P2_R1203_U401 = ~new_P2_U3951 | ~new_P2_R1203_U82;
  assign new_P2_R1203_U402 = ~new_P2_U3059 | ~new_P2_R1203_U45;
  assign new_P2_R1203_U403 = ~new_P2_R1203_U317 | ~new_P2_R1203_U88;
  assign new_P2_R1203_U404 = ~new_P2_R1203_U158 | ~new_P2_R1203_U299;
  assign new_P2_R1203_U405 = ~new_P2_U3952 | ~new_P2_R1203_U80;
  assign new_P2_R1203_U406 = ~new_P2_U3060 | ~new_P2_R1203_U79;
  assign new_P2_R1203_U407 = ~new_P2_R1203_U134;
  assign new_P2_R1203_U408 = ~new_P2_R1203_U295 | ~new_P2_R1203_U407;
  assign new_P2_R1203_U409 = ~new_P2_R1203_U134 | ~new_P2_R1203_U159;
  assign new_P2_R1203_U410 = ~new_P2_U3953 | ~new_P2_R1203_U78;
  assign new_P2_R1203_U411 = ~new_P2_U3067 | ~new_P2_R1203_U77;
  assign new_P2_R1203_U412 = ~new_P2_R1203_U135;
  assign new_P2_R1203_U413 = ~new_P2_R1203_U291 | ~new_P2_R1203_U412;
  assign new_P2_R1203_U414 = ~new_P2_R1203_U135 | ~new_P2_R1203_U160;
  assign new_P2_R1203_U415 = ~new_P2_U3954 | ~new_P2_R1203_U73;
  assign new_P2_R1203_U416 = ~new_P2_U3068 | ~new_P2_R1203_U70;
  assign new_P2_R1203_U417 = ~new_P2_R1203_U416 | ~new_P2_R1203_U415;
  assign new_P2_R1203_U418 = ~new_P2_U3955 | ~new_P2_R1203_U74;
  assign new_P2_R1203_U419 = ~new_P2_U3063 | ~new_P2_R1203_U71;
  assign new_P2_R1203_U420 = ~new_P2_R1203_U327 | ~new_P2_R1203_U89;
  assign new_P2_R1203_U421 = ~new_P2_R1203_U161 | ~new_P2_R1203_U319;
  assign new_P2_R1203_U422 = ~new_P2_U3956 | ~new_P2_R1203_U75;
  assign new_P2_R1203_U423 = ~new_P2_U3077 | ~new_P2_R1203_U72;
  assign new_P2_R1203_U424 = ~new_P2_R1203_U328 | ~new_P2_R1203_U163;
  assign new_P2_R1203_U425 = ~new_P2_R1203_U281 | ~new_P2_R1203_U162;
  assign new_P2_R1203_U426 = ~new_P2_U3957 | ~new_P2_R1203_U69;
  assign new_P2_R1203_U427 = ~new_P2_U3078 | ~new_P2_R1203_U68;
  assign new_P2_R1203_U428 = ~new_P2_R1203_U138;
  assign new_P2_R1203_U429 = ~new_P2_R1203_U277 | ~new_P2_R1203_U428;
  assign new_P2_R1203_U430 = ~new_P2_R1203_U138 | ~new_P2_R1203_U164;
  assign new_P2_R1203_U431 = ~new_P2_U3432 | ~new_P2_R1203_U25;
  assign new_P2_R1203_U432 = ~new_P2_U3080 | ~new_P2_R1203_U165;
  assign new_P2_R1203_U433 = ~new_P2_R1203_U139;
  assign new_P2_R1203_U434 = ~new_P2_R1203_U191 | ~new_P2_R1203_U433;
  assign new_P2_R1203_U435 = ~new_P2_R1203_U139 | ~new_P2_R1203_U166;
  assign new_P2_R1203_U436 = ~new_P2_U3485 | ~new_P2_R1203_U67;
  assign new_P2_R1203_U437 = ~new_P2_U3083 | ~new_P2_R1203_U66;
  assign new_P2_R1203_U438 = ~new_P2_R1203_U140;
  assign new_P2_R1203_U439 = ~new_P2_R1203_U273 | ~new_P2_R1203_U438;
  assign new_P2_R1203_U440 = ~new_P2_R1203_U140 | ~new_P2_R1203_U167;
  assign new_P2_R1203_U441 = ~new_P2_U3483 | ~new_P2_R1203_U65;
  assign new_P2_R1203_U442 = ~new_P2_U3084 | ~new_P2_R1203_U168;
  assign new_P2_R1203_U443 = ~new_P2_R1203_U141;
  assign new_P2_R1203_U444 = ~new_P2_R1203_U443 | ~new_P2_R1203_U269;
  assign new_P2_R1203_U445 = ~new_P2_R1203_U141 | ~new_P2_R1203_U64;
  assign new_P2_R1203_U446 = ~new_P2_U3480 | ~new_P2_R1203_U63;
  assign new_P2_R1203_U447 = ~new_P2_U3071 | ~new_P2_R1203_U62;
  assign new_P2_R1203_U448 = ~new_P2_R1203_U142;
  assign new_P2_R1203_U449 = ~new_P2_R1203_U265 | ~new_P2_R1203_U448;
  assign new_P2_R1203_U450 = ~new_P2_R1203_U142 | ~new_P2_R1203_U169;
  assign new_P2_R1203_U451 = ~new_P2_U3477 | ~new_P2_R1203_U58;
  assign new_P2_R1203_U452 = ~new_P2_U3075 | ~new_P2_R1203_U55;
  assign new_P2_R1203_U453 = ~new_P2_R1203_U452 | ~new_P2_R1203_U451;
  assign new_P2_R1203_U454 = ~new_P2_U3474 | ~new_P2_R1203_U59;
  assign new_P2_R1203_U455 = ~new_P2_U3076 | ~new_P2_R1203_U56;
  assign new_P2_R1203_U456 = ~new_P2_R1203_U338 | ~new_P2_R1203_U90;
  assign new_P2_R1203_U457 = ~new_P2_R1203_U170 | ~new_P2_R1203_U330;
  assign new_P2_R1203_U458 = ~new_P2_U3471 | ~new_P2_R1203_U60;
  assign new_P2_R1203_U459 = ~new_P2_U3081 | ~new_P2_R1203_U57;
  assign new_P2_R1203_U460 = ~new_P2_R1203_U339 | ~new_P2_R1203_U172;
  assign new_P2_R1203_U461 = ~new_P2_R1203_U255 | ~new_P2_R1203_U171;
  assign new_P2_R1203_U462 = ~new_P2_U3468 | ~new_P2_R1203_U54;
  assign new_P2_R1203_U463 = ~new_P2_U3082 | ~new_P2_R1203_U53;
  assign new_P2_R1203_U464 = ~new_P2_R1203_U145;
  assign new_P2_R1203_U465 = ~new_P2_R1203_U251 | ~new_P2_R1203_U464;
  assign new_P2_R1203_U466 = ~new_P2_R1203_U145 | ~new_P2_R1203_U173;
  assign new_P2_R1203_U467 = ~new_P2_U3465 | ~new_P2_R1203_U52;
  assign new_P2_R1203_U468 = ~new_P2_U3074 | ~new_P2_R1203_U51;
  assign new_P2_R1203_U469 = ~new_P2_R1203_U146;
  assign new_P2_R1203_U470 = ~new_P2_R1203_U247 | ~new_P2_R1203_U469;
  assign new_P2_R1203_U471 = ~new_P2_R1203_U146 | ~new_P2_R1203_U174;
  assign new_P2_R1203_U472 = ~new_P2_U3462 | ~new_P2_R1203_U48;
  assign new_P2_R1203_U473 = ~new_P2_U3065 | ~new_P2_R1203_U47;
  assign new_P2_R1203_U474 = ~new_P2_R1203_U473 | ~new_P2_R1203_U472;
  assign new_P2_R1203_U475 = ~new_P2_U3459 | ~new_P2_R1203_U49;
  assign new_P2_R1203_U476 = ~new_P2_U3064 | ~new_P2_R1203_U46;
  assign new_P2_R1203_U477 = ~new_P2_R1203_U349 | ~new_P2_R1203_U91;
  assign new_P2_R1203_U478 = ~new_P2_R1203_U175 | ~new_P2_R1203_U341;
  assign new_P2_R1113_U6 = new_P2_R1113_U202 & new_P2_R1113_U201;
  assign new_P2_R1113_U7 = new_P2_R1113_U241 & new_P2_R1113_U240;
  assign new_P2_R1113_U8 = new_P2_R1113_U181 & new_P2_R1113_U256;
  assign new_P2_R1113_U9 = new_P2_R1113_U258 & new_P2_R1113_U257;
  assign new_P2_R1113_U10 = new_P2_R1113_U182 & new_P2_R1113_U282;
  assign new_P2_R1113_U11 = new_P2_R1113_U284 & new_P2_R1113_U283;
  assign new_P2_R1113_U12 = ~new_P2_R1113_U344 | ~new_P2_R1113_U347;
  assign new_P2_R1113_U13 = ~new_P2_R1113_U333 | ~new_P2_R1113_U336;
  assign new_P2_R1113_U14 = ~new_P2_R1113_U322 | ~new_P2_R1113_U325;
  assign new_P2_R1113_U15 = ~new_P2_R1113_U314 | ~new_P2_R1113_U316;
  assign new_P2_R1113_U16 = ~new_P2_R1113_U352 | ~new_P2_R1113_U312;
  assign new_P2_R1113_U17 = ~new_P2_R1113_U235 | ~new_P2_R1113_U237;
  assign new_P2_R1113_U18 = ~new_P2_R1113_U227 | ~new_P2_R1113_U230;
  assign new_P2_R1113_U19 = ~new_P2_R1113_U219 | ~new_P2_R1113_U221;
  assign new_P2_R1113_U20 = ~new_P2_R1113_U166 | ~new_P2_R1113_U350;
  assign new_P2_R1113_U21 = ~new_P2_U3450;
  assign new_P2_R1113_U22 = ~new_P2_U3444;
  assign new_P2_R1113_U23 = ~new_P2_U3435;
  assign new_P2_R1113_U24 = ~new_P2_U3427;
  assign new_P2_R1113_U25 = ~new_P2_U3080;
  assign new_P2_R1113_U26 = ~new_P2_U3438;
  assign new_P2_R1113_U27 = ~new_P2_U3070;
  assign new_P2_R1113_U28 = ~new_P2_U3070 | ~new_P2_R1113_U23;
  assign new_P2_R1113_U29 = ~new_P2_U3066;
  assign new_P2_R1113_U30 = ~new_P2_U3447;
  assign new_P2_R1113_U31 = ~new_P2_U3441;
  assign new_P2_R1113_U32 = ~new_P2_U3073;
  assign new_P2_R1113_U33 = ~new_P2_U3069;
  assign new_P2_R1113_U34 = ~new_P2_U3062;
  assign new_P2_R1113_U35 = ~new_P2_U3062 | ~new_P2_R1113_U31;
  assign new_P2_R1113_U36 = ~new_P2_U3453;
  assign new_P2_R1113_U37 = ~new_P2_U3072;
  assign new_P2_R1113_U38 = ~new_P2_U3072 | ~new_P2_R1113_U21;
  assign new_P2_R1113_U39 = ~new_P2_U3086;
  assign new_P2_R1113_U40 = ~new_P2_U3456;
  assign new_P2_R1113_U41 = ~new_P2_U3085;
  assign new_P2_R1113_U42 = ~new_P2_R1113_U208 | ~new_P2_R1113_U207;
  assign new_P2_R1113_U43 = ~new_P2_R1113_U35 | ~new_P2_R1113_U223;
  assign new_P2_R1113_U44 = ~new_P2_R1113_U351 | ~new_P2_R1113_U192 | ~new_P2_R1113_U176;
  assign new_P2_R1113_U45 = ~new_P2_U3951;
  assign new_P2_R1113_U46 = ~new_P2_U3459;
  assign new_P2_R1113_U47 = ~new_P2_U3462;
  assign new_P2_R1113_U48 = ~new_P2_U3065;
  assign new_P2_R1113_U49 = ~new_P2_U3064;
  assign new_P2_R1113_U50 = ~new_P2_U3085 | ~new_P2_R1113_U40;
  assign new_P2_R1113_U51 = ~new_P2_U3465;
  assign new_P2_R1113_U52 = ~new_P2_U3074;
  assign new_P2_R1113_U53 = ~new_P2_U3468;
  assign new_P2_R1113_U54 = ~new_P2_U3082;
  assign new_P2_R1113_U55 = ~new_P2_U3477;
  assign new_P2_R1113_U56 = ~new_P2_U3474;
  assign new_P2_R1113_U57 = ~new_P2_U3471;
  assign new_P2_R1113_U58 = ~new_P2_U3075;
  assign new_P2_R1113_U59 = ~new_P2_U3076;
  assign new_P2_R1113_U60 = ~new_P2_U3081;
  assign new_P2_R1113_U61 = ~new_P2_U3081 | ~new_P2_R1113_U57;
  assign new_P2_R1113_U62 = ~new_P2_U3480;
  assign new_P2_R1113_U63 = ~new_P2_U3071;
  assign new_P2_R1113_U64 = ~new_P2_R1113_U268 | ~new_P2_R1113_U267;
  assign new_P2_R1113_U65 = ~new_P2_U3084;
  assign new_P2_R1113_U66 = ~new_P2_U3485;
  assign new_P2_R1113_U67 = ~new_P2_U3083;
  assign new_P2_R1113_U68 = ~new_P2_U3957;
  assign new_P2_R1113_U69 = ~new_P2_U3078;
  assign new_P2_R1113_U70 = ~new_P2_U3954;
  assign new_P2_R1113_U71 = ~new_P2_U3955;
  assign new_P2_R1113_U72 = ~new_P2_U3956;
  assign new_P2_R1113_U73 = ~new_P2_U3068;
  assign new_P2_R1113_U74 = ~new_P2_U3063;
  assign new_P2_R1113_U75 = ~new_P2_U3077;
  assign new_P2_R1113_U76 = ~new_P2_U3077 | ~new_P2_R1113_U72;
  assign new_P2_R1113_U77 = ~new_P2_U3953;
  assign new_P2_R1113_U78 = ~new_P2_U3067;
  assign new_P2_R1113_U79 = ~new_P2_U3952;
  assign new_P2_R1113_U80 = ~new_P2_U3060;
  assign new_P2_R1113_U81 = ~new_P2_U3950;
  assign new_P2_R1113_U82 = ~new_P2_U3059;
  assign new_P2_R1113_U83 = ~new_P2_U3059 | ~new_P2_R1113_U45;
  assign new_P2_R1113_U84 = ~new_P2_U3055;
  assign new_P2_R1113_U85 = ~new_P2_U3949;
  assign new_P2_R1113_U86 = ~new_P2_U3056;
  assign new_P2_R1113_U87 = ~new_P2_R1113_U128 | ~new_P2_R1113_U301;
  assign new_P2_R1113_U88 = ~new_P2_R1113_U298 | ~new_P2_R1113_U297;
  assign new_P2_R1113_U89 = ~new_P2_R1113_U76 | ~new_P2_R1113_U318;
  assign new_P2_R1113_U90 = ~new_P2_R1113_U61 | ~new_P2_R1113_U329;
  assign new_P2_R1113_U91 = ~new_P2_R1113_U50 | ~new_P2_R1113_U340;
  assign new_P2_R1113_U92 = ~new_P2_U3079;
  assign new_P2_R1113_U93 = ~new_P2_R1113_U395 | ~new_P2_R1113_U394;
  assign new_P2_R1113_U94 = ~new_P2_R1113_U409 | ~new_P2_R1113_U408;
  assign new_P2_R1113_U95 = ~new_P2_R1113_U414 | ~new_P2_R1113_U413;
  assign new_P2_R1113_U96 = ~new_P2_R1113_U430 | ~new_P2_R1113_U429;
  assign new_P2_R1113_U97 = ~new_P2_R1113_U435 | ~new_P2_R1113_U434;
  assign new_P2_R1113_U98 = ~new_P2_R1113_U440 | ~new_P2_R1113_U439;
  assign new_P2_R1113_U99 = ~new_P2_R1113_U445 | ~new_P2_R1113_U444;
  assign new_P2_R1113_U100 = ~new_P2_R1113_U450 | ~new_P2_R1113_U449;
  assign new_P2_R1113_U101 = ~new_P2_R1113_U466 | ~new_P2_R1113_U465;
  assign new_P2_R1113_U102 = ~new_P2_R1113_U471 | ~new_P2_R1113_U470;
  assign new_P2_R1113_U103 = ~new_P2_R1113_U356 | ~new_P2_R1113_U355;
  assign new_P2_R1113_U104 = ~new_P2_R1113_U365 | ~new_P2_R1113_U364;
  assign new_P2_R1113_U105 = ~new_P2_R1113_U372 | ~new_P2_R1113_U371;
  assign new_P2_R1113_U106 = ~new_P2_R1113_U376 | ~new_P2_R1113_U375;
  assign new_P2_R1113_U107 = ~new_P2_R1113_U385 | ~new_P2_R1113_U384;
  assign new_P2_R1113_U108 = ~new_P2_R1113_U404 | ~new_P2_R1113_U403;
  assign new_P2_R1113_U109 = ~new_P2_R1113_U421 | ~new_P2_R1113_U420;
  assign new_P2_R1113_U110 = ~new_P2_R1113_U425 | ~new_P2_R1113_U424;
  assign new_P2_R1113_U111 = ~new_P2_R1113_U457 | ~new_P2_R1113_U456;
  assign new_P2_R1113_U112 = ~new_P2_R1113_U461 | ~new_P2_R1113_U460;
  assign new_P2_R1113_U113 = ~new_P2_R1113_U478 | ~new_P2_R1113_U477;
  assign new_P2_R1113_U114 = new_P2_R1113_U194 & new_P2_R1113_U184;
  assign new_P2_R1113_U115 = new_P2_R1113_U197 & new_P2_R1113_U198;
  assign new_P2_R1113_U116 = new_P2_R1113_U185 & new_P2_R1113_U205 & new_P2_R1113_U200;
  assign new_P2_R1113_U117 = new_P2_R1113_U210 & new_P2_R1113_U186;
  assign new_P2_R1113_U118 = new_P2_R1113_U213 & new_P2_R1113_U214;
  assign new_P2_R1113_U119 = new_P2_R1113_U38 & new_P2_R1113_U358 & new_P2_R1113_U357;
  assign new_P2_R1113_U120 = new_P2_R1113_U361 & new_P2_R1113_U186;
  assign new_P2_R1113_U121 = new_P2_R1113_U229 & new_P2_R1113_U6;
  assign new_P2_R1113_U122 = new_P2_R1113_U368 & new_P2_R1113_U185;
  assign new_P2_R1113_U123 = new_P2_R1113_U28 & new_P2_R1113_U378 & new_P2_R1113_U377;
  assign new_P2_R1113_U124 = new_P2_R1113_U381 & new_P2_R1113_U184;
  assign new_P2_R1113_U125 = new_P2_R1113_U180 & new_P2_R1113_U239 & new_P2_R1113_U216;
  assign new_P2_R1113_U126 = new_P2_R1113_U261 & new_P2_R1113_U8;
  assign new_P2_R1113_U127 = new_P2_R1113_U287 & new_P2_R1113_U10;
  assign new_P2_R1113_U128 = new_P2_R1113_U303 & new_P2_R1113_U304;
  assign new_P2_R1113_U129 = new_P2_R1113_U311 & new_P2_R1113_U387 & new_P2_R1113_U386;
  assign new_P2_R1113_U130 = new_P2_R1113_U308 & new_P2_R1113_U390;
  assign new_P2_R1113_U131 = ~new_P2_R1113_U392 | ~new_P2_R1113_U391;
  assign new_P2_R1113_U132 = new_P2_R1113_U83 & new_P2_R1113_U397 & new_P2_R1113_U396;
  assign new_P2_R1113_U133 = new_P2_R1113_U400 & new_P2_R1113_U183;
  assign new_P2_R1113_U134 = ~new_P2_R1113_U406 | ~new_P2_R1113_U405;
  assign new_P2_R1113_U135 = ~new_P2_R1113_U411 | ~new_P2_R1113_U410;
  assign new_P2_R1113_U136 = new_P2_R1113_U324 & new_P2_R1113_U11;
  assign new_P2_R1113_U137 = new_P2_R1113_U417 & new_P2_R1113_U182;
  assign new_P2_R1113_U138 = ~new_P2_R1113_U427 | ~new_P2_R1113_U426;
  assign new_P2_R1113_U139 = ~new_P2_R1113_U432 | ~new_P2_R1113_U431;
  assign new_P2_R1113_U140 = ~new_P2_R1113_U437 | ~new_P2_R1113_U436;
  assign new_P2_R1113_U141 = ~new_P2_R1113_U442 | ~new_P2_R1113_U441;
  assign new_P2_R1113_U142 = ~new_P2_R1113_U447 | ~new_P2_R1113_U446;
  assign new_P2_R1113_U143 = new_P2_R1113_U335 & new_P2_R1113_U9;
  assign new_P2_R1113_U144 = new_P2_R1113_U453 & new_P2_R1113_U181;
  assign new_P2_R1113_U145 = ~new_P2_R1113_U463 | ~new_P2_R1113_U462;
  assign new_P2_R1113_U146 = ~new_P2_R1113_U468 | ~new_P2_R1113_U467;
  assign new_P2_R1113_U147 = new_P2_R1113_U346 & new_P2_R1113_U7;
  assign new_P2_R1113_U148 = new_P2_R1113_U474 & new_P2_R1113_U180;
  assign new_P2_R1113_U149 = new_P2_R1113_U354 & new_P2_R1113_U353;
  assign new_P2_R1113_U150 = ~new_P2_R1113_U118 | ~new_P2_R1113_U211;
  assign new_P2_R1113_U151 = new_P2_R1113_U363 & new_P2_R1113_U362;
  assign new_P2_R1113_U152 = new_P2_R1113_U370 & new_P2_R1113_U369;
  assign new_P2_R1113_U153 = new_P2_R1113_U374 & new_P2_R1113_U373;
  assign new_P2_R1113_U154 = ~new_P2_R1113_U115 | ~new_P2_R1113_U195;
  assign new_P2_R1113_U155 = new_P2_R1113_U383 & new_P2_R1113_U382;
  assign new_P2_R1113_U156 = ~new_P2_U3960;
  assign new_P2_R1113_U157 = ~new_P2_U3057;
  assign new_P2_R1113_U158 = new_P2_R1113_U402 & new_P2_R1113_U401;
  assign new_P2_R1113_U159 = ~new_P2_R1113_U294 | ~new_P2_R1113_U293;
  assign new_P2_R1113_U160 = ~new_P2_R1113_U290 | ~new_P2_R1113_U289;
  assign new_P2_R1113_U161 = new_P2_R1113_U419 & new_P2_R1113_U418;
  assign new_P2_R1113_U162 = new_P2_R1113_U423 & new_P2_R1113_U422;
  assign new_P2_R1113_U163 = ~new_P2_R1113_U280 | ~new_P2_R1113_U279;
  assign new_P2_R1113_U164 = ~new_P2_R1113_U276 | ~new_P2_R1113_U275;
  assign new_P2_R1113_U165 = ~new_P2_U3432;
  assign new_P2_R1113_U166 = ~new_P2_U3427 | ~new_P2_R1113_U92;
  assign new_P2_R1113_U167 = ~new_P2_R1113_U272 | ~new_P2_R1113_U271;
  assign new_P2_R1113_U168 = ~new_P2_U3483;
  assign new_P2_R1113_U169 = ~new_P2_R1113_U264 | ~new_P2_R1113_U263;
  assign new_P2_R1113_U170 = new_P2_R1113_U455 & new_P2_R1113_U454;
  assign new_P2_R1113_U171 = new_P2_R1113_U459 & new_P2_R1113_U458;
  assign new_P2_R1113_U172 = ~new_P2_R1113_U254 | ~new_P2_R1113_U253;
  assign new_P2_R1113_U173 = ~new_P2_R1113_U250 | ~new_P2_R1113_U249;
  assign new_P2_R1113_U174 = ~new_P2_R1113_U246 | ~new_P2_R1113_U245;
  assign new_P2_R1113_U175 = new_P2_R1113_U476 & new_P2_R1113_U475;
  assign new_P2_R1113_U176 = ~new_P2_R1113_U166 | ~new_P2_R1113_U165;
  assign new_P2_R1113_U177 = ~new_P2_R1113_U83;
  assign new_P2_R1113_U178 = ~new_P2_R1113_U28;
  assign new_P2_R1113_U179 = ~new_P2_R1113_U38;
  assign new_P2_R1113_U180 = ~new_P2_U3459 | ~new_P2_R1113_U49;
  assign new_P2_R1113_U181 = ~new_P2_U3474 | ~new_P2_R1113_U59;
  assign new_P2_R1113_U182 = ~new_P2_U3955 | ~new_P2_R1113_U74;
  assign new_P2_R1113_U183 = ~new_P2_U3951 | ~new_P2_R1113_U82;
  assign new_P2_R1113_U184 = ~new_P2_U3435 | ~new_P2_R1113_U27;
  assign new_P2_R1113_U185 = ~new_P2_U3444 | ~new_P2_R1113_U33;
  assign new_P2_R1113_U186 = ~new_P2_U3450 | ~new_P2_R1113_U37;
  assign new_P2_R1113_U187 = ~new_P2_R1113_U61;
  assign new_P2_R1113_U188 = ~new_P2_R1113_U76;
  assign new_P2_R1113_U189 = ~new_P2_R1113_U35;
  assign new_P2_R1113_U190 = ~new_P2_R1113_U50;
  assign new_P2_R1113_U191 = ~new_P2_R1113_U166;
  assign new_P2_R1113_U192 = ~new_P2_U3080 | ~new_P2_R1113_U166;
  assign new_P2_R1113_U193 = ~new_P2_R1113_U44;
  assign new_P2_R1113_U194 = ~new_P2_U3438 | ~new_P2_R1113_U29;
  assign new_P2_R1113_U195 = ~new_P2_R1113_U114 | ~new_P2_R1113_U44;
  assign new_P2_R1113_U196 = ~new_P2_R1113_U29 | ~new_P2_R1113_U28;
  assign new_P2_R1113_U197 = ~new_P2_R1113_U196 | ~new_P2_R1113_U26;
  assign new_P2_R1113_U198 = ~new_P2_U3066 | ~new_P2_R1113_U178;
  assign new_P2_R1113_U199 = ~new_P2_R1113_U154;
  assign new_P2_R1113_U200 = ~new_P2_U3447 | ~new_P2_R1113_U32;
  assign new_P2_R1113_U201 = ~new_P2_U3073 | ~new_P2_R1113_U30;
  assign new_P2_R1113_U202 = ~new_P2_U3069 | ~new_P2_R1113_U22;
  assign new_P2_R1113_U203 = ~new_P2_R1113_U189 | ~new_P2_R1113_U185;
  assign new_P2_R1113_U204 = ~new_P2_R1113_U6 | ~new_P2_R1113_U203;
  assign new_P2_R1113_U205 = ~new_P2_U3441 | ~new_P2_R1113_U34;
  assign new_P2_R1113_U206 = ~new_P2_U3447 | ~new_P2_R1113_U32;
  assign new_P2_R1113_U207 = ~new_P2_R1113_U154 | ~new_P2_R1113_U116;
  assign new_P2_R1113_U208 = ~new_P2_R1113_U206 | ~new_P2_R1113_U204;
  assign new_P2_R1113_U209 = ~new_P2_R1113_U42;
  assign new_P2_R1113_U210 = ~new_P2_U3453 | ~new_P2_R1113_U39;
  assign new_P2_R1113_U211 = ~new_P2_R1113_U117 | ~new_P2_R1113_U42;
  assign new_P2_R1113_U212 = ~new_P2_R1113_U39 | ~new_P2_R1113_U38;
  assign new_P2_R1113_U213 = ~new_P2_R1113_U212 | ~new_P2_R1113_U36;
  assign new_P2_R1113_U214 = ~new_P2_U3086 | ~new_P2_R1113_U179;
  assign new_P2_R1113_U215 = ~new_P2_R1113_U150;
  assign new_P2_R1113_U216 = ~new_P2_U3456 | ~new_P2_R1113_U41;
  assign new_P2_R1113_U217 = ~new_P2_R1113_U216 | ~new_P2_R1113_U50;
  assign new_P2_R1113_U218 = ~new_P2_R1113_U209 | ~new_P2_R1113_U38;
  assign new_P2_R1113_U219 = ~new_P2_R1113_U120 | ~new_P2_R1113_U218;
  assign new_P2_R1113_U220 = ~new_P2_R1113_U42 | ~new_P2_R1113_U186;
  assign new_P2_R1113_U221 = ~new_P2_R1113_U119 | ~new_P2_R1113_U220;
  assign new_P2_R1113_U222 = ~new_P2_R1113_U38 | ~new_P2_R1113_U186;
  assign new_P2_R1113_U223 = ~new_P2_R1113_U205 | ~new_P2_R1113_U154;
  assign new_P2_R1113_U224 = ~new_P2_R1113_U43;
  assign new_P2_R1113_U225 = ~new_P2_U3069 | ~new_P2_R1113_U22;
  assign new_P2_R1113_U226 = ~new_P2_R1113_U224 | ~new_P2_R1113_U225;
  assign new_P2_R1113_U227 = ~new_P2_R1113_U122 | ~new_P2_R1113_U226;
  assign new_P2_R1113_U228 = ~new_P2_R1113_U43 | ~new_P2_R1113_U185;
  assign new_P2_R1113_U229 = ~new_P2_U3447 | ~new_P2_R1113_U32;
  assign new_P2_R1113_U230 = ~new_P2_R1113_U121 | ~new_P2_R1113_U228;
  assign new_P2_R1113_U231 = ~new_P2_U3069 | ~new_P2_R1113_U22;
  assign new_P2_R1113_U232 = ~new_P2_R1113_U185 | ~new_P2_R1113_U231;
  assign new_P2_R1113_U233 = ~new_P2_R1113_U205 | ~new_P2_R1113_U35;
  assign new_P2_R1113_U234 = ~new_P2_R1113_U193 | ~new_P2_R1113_U28;
  assign new_P2_R1113_U235 = ~new_P2_R1113_U124 | ~new_P2_R1113_U234;
  assign new_P2_R1113_U236 = ~new_P2_R1113_U44 | ~new_P2_R1113_U184;
  assign new_P2_R1113_U237 = ~new_P2_R1113_U123 | ~new_P2_R1113_U236;
  assign new_P2_R1113_U238 = ~new_P2_R1113_U28 | ~new_P2_R1113_U184;
  assign new_P2_R1113_U239 = ~new_P2_U3462 | ~new_P2_R1113_U48;
  assign new_P2_R1113_U240 = ~new_P2_U3065 | ~new_P2_R1113_U47;
  assign new_P2_R1113_U241 = ~new_P2_U3064 | ~new_P2_R1113_U46;
  assign new_P2_R1113_U242 = ~new_P2_R1113_U190 | ~new_P2_R1113_U180;
  assign new_P2_R1113_U243 = ~new_P2_R1113_U7 | ~new_P2_R1113_U242;
  assign new_P2_R1113_U244 = ~new_P2_U3462 | ~new_P2_R1113_U48;
  assign new_P2_R1113_U245 = ~new_P2_R1113_U150 | ~new_P2_R1113_U125;
  assign new_P2_R1113_U246 = ~new_P2_R1113_U244 | ~new_P2_R1113_U243;
  assign new_P2_R1113_U247 = ~new_P2_R1113_U174;
  assign new_P2_R1113_U248 = ~new_P2_U3465 | ~new_P2_R1113_U52;
  assign new_P2_R1113_U249 = ~new_P2_R1113_U248 | ~new_P2_R1113_U174;
  assign new_P2_R1113_U250 = ~new_P2_U3074 | ~new_P2_R1113_U51;
  assign new_P2_R1113_U251 = ~new_P2_R1113_U173;
  assign new_P2_R1113_U252 = ~new_P2_U3468 | ~new_P2_R1113_U54;
  assign new_P2_R1113_U253 = ~new_P2_R1113_U252 | ~new_P2_R1113_U173;
  assign new_P2_R1113_U254 = ~new_P2_U3082 | ~new_P2_R1113_U53;
  assign new_P2_R1113_U255 = ~new_P2_R1113_U172;
  assign new_P2_R1113_U256 = ~new_P2_U3477 | ~new_P2_R1113_U58;
  assign new_P2_R1113_U257 = ~new_P2_U3075 | ~new_P2_R1113_U55;
  assign new_P2_R1113_U258 = ~new_P2_U3076 | ~new_P2_R1113_U56;
  assign new_P2_R1113_U259 = ~new_P2_R1113_U187 | ~new_P2_R1113_U8;
  assign new_P2_R1113_U260 = ~new_P2_R1113_U9 | ~new_P2_R1113_U259;
  assign new_P2_R1113_U261 = ~new_P2_U3471 | ~new_P2_R1113_U60;
  assign new_P2_R1113_U262 = ~new_P2_U3477 | ~new_P2_R1113_U58;
  assign new_P2_R1113_U263 = ~new_P2_R1113_U126 | ~new_P2_R1113_U172;
  assign new_P2_R1113_U264 = ~new_P2_R1113_U262 | ~new_P2_R1113_U260;
  assign new_P2_R1113_U265 = ~new_P2_R1113_U169;
  assign new_P2_R1113_U266 = ~new_P2_U3480 | ~new_P2_R1113_U63;
  assign new_P2_R1113_U267 = ~new_P2_R1113_U266 | ~new_P2_R1113_U169;
  assign new_P2_R1113_U268 = ~new_P2_U3071 | ~new_P2_R1113_U62;
  assign new_P2_R1113_U269 = ~new_P2_R1113_U64;
  assign new_P2_R1113_U270 = ~new_P2_R1113_U269 | ~new_P2_R1113_U65;
  assign new_P2_R1113_U271 = ~new_P2_R1113_U270 | ~new_P2_R1113_U168;
  assign new_P2_R1113_U272 = ~new_P2_U3084 | ~new_P2_R1113_U64;
  assign new_P2_R1113_U273 = ~new_P2_R1113_U167;
  assign new_P2_R1113_U274 = ~new_P2_U3485 | ~new_P2_R1113_U67;
  assign new_P2_R1113_U275 = ~new_P2_R1113_U274 | ~new_P2_R1113_U167;
  assign new_P2_R1113_U276 = ~new_P2_U3083 | ~new_P2_R1113_U66;
  assign new_P2_R1113_U277 = ~new_P2_R1113_U164;
  assign new_P2_R1113_U278 = ~new_P2_U3957 | ~new_P2_R1113_U69;
  assign new_P2_R1113_U279 = ~new_P2_R1113_U278 | ~new_P2_R1113_U164;
  assign new_P2_R1113_U280 = ~new_P2_U3078 | ~new_P2_R1113_U68;
  assign new_P2_R1113_U281 = ~new_P2_R1113_U163;
  assign new_P2_R1113_U282 = ~new_P2_U3954 | ~new_P2_R1113_U73;
  assign new_P2_R1113_U283 = ~new_P2_U3068 | ~new_P2_R1113_U70;
  assign new_P2_R1113_U284 = ~new_P2_U3063 | ~new_P2_R1113_U71;
  assign new_P2_R1113_U285 = ~new_P2_R1113_U188 | ~new_P2_R1113_U10;
  assign new_P2_R1113_U286 = ~new_P2_R1113_U11 | ~new_P2_R1113_U285;
  assign new_P2_R1113_U287 = ~new_P2_U3956 | ~new_P2_R1113_U75;
  assign new_P2_R1113_U288 = ~new_P2_U3954 | ~new_P2_R1113_U73;
  assign new_P2_R1113_U289 = ~new_P2_R1113_U127 | ~new_P2_R1113_U163;
  assign new_P2_R1113_U290 = ~new_P2_R1113_U288 | ~new_P2_R1113_U286;
  assign new_P2_R1113_U291 = ~new_P2_R1113_U160;
  assign new_P2_R1113_U292 = ~new_P2_U3953 | ~new_P2_R1113_U78;
  assign new_P2_R1113_U293 = ~new_P2_R1113_U292 | ~new_P2_R1113_U160;
  assign new_P2_R1113_U294 = ~new_P2_U3067 | ~new_P2_R1113_U77;
  assign new_P2_R1113_U295 = ~new_P2_R1113_U159;
  assign new_P2_R1113_U296 = ~new_P2_U3952 | ~new_P2_R1113_U80;
  assign new_P2_R1113_U297 = ~new_P2_R1113_U296 | ~new_P2_R1113_U159;
  assign new_P2_R1113_U298 = ~new_P2_U3060 | ~new_P2_R1113_U79;
  assign new_P2_R1113_U299 = ~new_P2_R1113_U88;
  assign new_P2_R1113_U300 = ~new_P2_U3950 | ~new_P2_R1113_U84;
  assign new_P2_R1113_U301 = ~new_P2_R1113_U300 | ~new_P2_R1113_U88 | ~new_P2_R1113_U183;
  assign new_P2_R1113_U302 = ~new_P2_R1113_U84 | ~new_P2_R1113_U83;
  assign new_P2_R1113_U303 = ~new_P2_R1113_U302 | ~new_P2_R1113_U81;
  assign new_P2_R1113_U304 = ~new_P2_U3055 | ~new_P2_R1113_U177;
  assign new_P2_R1113_U305 = ~new_P2_R1113_U87;
  assign new_P2_R1113_U306 = ~new_P2_U3056 | ~new_P2_R1113_U85;
  assign new_P2_R1113_U307 = ~new_P2_R1113_U305 | ~new_P2_R1113_U306;
  assign new_P2_R1113_U308 = ~new_P2_U3949 | ~new_P2_R1113_U86;
  assign new_P2_R1113_U309 = ~new_P2_U3949 | ~new_P2_R1113_U86;
  assign new_P2_R1113_U310 = ~new_P2_R1113_U309 | ~new_P2_R1113_U87;
  assign new_P2_R1113_U311 = ~new_P2_U3056 | ~new_P2_R1113_U85;
  assign new_P2_R1113_U312 = ~new_P2_R1113_U129 | ~new_P2_R1113_U310;
  assign new_P2_R1113_U313 = ~new_P2_R1113_U299 | ~new_P2_R1113_U83;
  assign new_P2_R1113_U314 = ~new_P2_R1113_U133 | ~new_P2_R1113_U313;
  assign new_P2_R1113_U315 = ~new_P2_R1113_U88 | ~new_P2_R1113_U183;
  assign new_P2_R1113_U316 = ~new_P2_R1113_U132 | ~new_P2_R1113_U315;
  assign new_P2_R1113_U317 = ~new_P2_R1113_U83 | ~new_P2_R1113_U183;
  assign new_P2_R1113_U318 = ~new_P2_R1113_U287 | ~new_P2_R1113_U163;
  assign new_P2_R1113_U319 = ~new_P2_R1113_U89;
  assign new_P2_R1113_U320 = ~new_P2_U3063 | ~new_P2_R1113_U71;
  assign new_P2_R1113_U321 = ~new_P2_R1113_U319 | ~new_P2_R1113_U320;
  assign new_P2_R1113_U322 = ~new_P2_R1113_U137 | ~new_P2_R1113_U321;
  assign new_P2_R1113_U323 = ~new_P2_R1113_U89 | ~new_P2_R1113_U182;
  assign new_P2_R1113_U324 = ~new_P2_U3954 | ~new_P2_R1113_U73;
  assign new_P2_R1113_U325 = ~new_P2_R1113_U136 | ~new_P2_R1113_U323;
  assign new_P2_R1113_U326 = ~new_P2_U3063 | ~new_P2_R1113_U71;
  assign new_P2_R1113_U327 = ~new_P2_R1113_U182 | ~new_P2_R1113_U326;
  assign new_P2_R1113_U328 = ~new_P2_R1113_U287 | ~new_P2_R1113_U76;
  assign new_P2_R1113_U329 = ~new_P2_R1113_U261 | ~new_P2_R1113_U172;
  assign new_P2_R1113_U330 = ~new_P2_R1113_U90;
  assign new_P2_R1113_U331 = ~new_P2_U3076 | ~new_P2_R1113_U56;
  assign new_P2_R1113_U332 = ~new_P2_R1113_U330 | ~new_P2_R1113_U331;
  assign new_P2_R1113_U333 = ~new_P2_R1113_U144 | ~new_P2_R1113_U332;
  assign new_P2_R1113_U334 = ~new_P2_R1113_U90 | ~new_P2_R1113_U181;
  assign new_P2_R1113_U335 = ~new_P2_U3477 | ~new_P2_R1113_U58;
  assign new_P2_R1113_U336 = ~new_P2_R1113_U143 | ~new_P2_R1113_U334;
  assign new_P2_R1113_U337 = ~new_P2_U3076 | ~new_P2_R1113_U56;
  assign new_P2_R1113_U338 = ~new_P2_R1113_U181 | ~new_P2_R1113_U337;
  assign new_P2_R1113_U339 = ~new_P2_R1113_U261 | ~new_P2_R1113_U61;
  assign new_P2_R1113_U340 = ~new_P2_R1113_U216 | ~new_P2_R1113_U150;
  assign new_P2_R1113_U341 = ~new_P2_R1113_U91;
  assign new_P2_R1113_U342 = ~new_P2_U3064 | ~new_P2_R1113_U46;
  assign new_P2_R1113_U343 = ~new_P2_R1113_U341 | ~new_P2_R1113_U342;
  assign new_P2_R1113_U344 = ~new_P2_R1113_U148 | ~new_P2_R1113_U343;
  assign new_P2_R1113_U345 = ~new_P2_R1113_U91 | ~new_P2_R1113_U180;
  assign new_P2_R1113_U346 = ~new_P2_U3462 | ~new_P2_R1113_U48;
  assign new_P2_R1113_U347 = ~new_P2_R1113_U147 | ~new_P2_R1113_U345;
  assign new_P2_R1113_U348 = ~new_P2_U3064 | ~new_P2_R1113_U46;
  assign new_P2_R1113_U349 = ~new_P2_R1113_U180 | ~new_P2_R1113_U348;
  assign new_P2_R1113_U350 = ~new_P2_U3079 | ~new_P2_R1113_U24;
  assign new_P2_R1113_U351 = ~new_P2_U3080 | ~new_P2_R1113_U165;
  assign new_P2_R1113_U352 = ~new_P2_R1113_U130 | ~new_P2_R1113_U307;
  assign new_P2_R1113_U353 = ~new_P2_U3456 | ~new_P2_R1113_U41;
  assign new_P2_R1113_U354 = ~new_P2_U3085 | ~new_P2_R1113_U40;
  assign new_P2_R1113_U355 = ~new_P2_R1113_U217 | ~new_P2_R1113_U150;
  assign new_P2_R1113_U356 = ~new_P2_R1113_U215 | ~new_P2_R1113_U149;
  assign new_P2_R1113_U357 = ~new_P2_U3453 | ~new_P2_R1113_U39;
  assign new_P2_R1113_U358 = ~new_P2_U3086 | ~new_P2_R1113_U36;
  assign new_P2_R1113_U359 = ~new_P2_U3453 | ~new_P2_R1113_U39;
  assign new_P2_R1113_U360 = ~new_P2_U3086 | ~new_P2_R1113_U36;
  assign new_P2_R1113_U361 = ~new_P2_R1113_U360 | ~new_P2_R1113_U359;
  assign new_P2_R1113_U362 = ~new_P2_U3450 | ~new_P2_R1113_U37;
  assign new_P2_R1113_U363 = ~new_P2_U3072 | ~new_P2_R1113_U21;
  assign new_P2_R1113_U364 = ~new_P2_R1113_U222 | ~new_P2_R1113_U42;
  assign new_P2_R1113_U365 = ~new_P2_R1113_U151 | ~new_P2_R1113_U209;
  assign new_P2_R1113_U366 = ~new_P2_U3447 | ~new_P2_R1113_U32;
  assign new_P2_R1113_U367 = ~new_P2_U3073 | ~new_P2_R1113_U30;
  assign new_P2_R1113_U368 = ~new_P2_R1113_U367 | ~new_P2_R1113_U366;
  assign new_P2_R1113_U369 = ~new_P2_U3444 | ~new_P2_R1113_U33;
  assign new_P2_R1113_U370 = ~new_P2_U3069 | ~new_P2_R1113_U22;
  assign new_P2_R1113_U371 = ~new_P2_R1113_U232 | ~new_P2_R1113_U43;
  assign new_P2_R1113_U372 = ~new_P2_R1113_U152 | ~new_P2_R1113_U224;
  assign new_P2_R1113_U373 = ~new_P2_U3441 | ~new_P2_R1113_U34;
  assign new_P2_R1113_U374 = ~new_P2_U3062 | ~new_P2_R1113_U31;
  assign new_P2_R1113_U375 = ~new_P2_R1113_U233 | ~new_P2_R1113_U154;
  assign new_P2_R1113_U376 = ~new_P2_R1113_U199 | ~new_P2_R1113_U153;
  assign new_P2_R1113_U377 = ~new_P2_U3438 | ~new_P2_R1113_U29;
  assign new_P2_R1113_U378 = ~new_P2_U3066 | ~new_P2_R1113_U26;
  assign new_P2_R1113_U379 = ~new_P2_U3438 | ~new_P2_R1113_U29;
  assign new_P2_R1113_U380 = ~new_P2_U3066 | ~new_P2_R1113_U26;
  assign new_P2_R1113_U381 = ~new_P2_R1113_U380 | ~new_P2_R1113_U379;
  assign new_P2_R1113_U382 = ~new_P2_U3435 | ~new_P2_R1113_U27;
  assign new_P2_R1113_U383 = ~new_P2_U3070 | ~new_P2_R1113_U23;
  assign new_P2_R1113_U384 = ~new_P2_R1113_U238 | ~new_P2_R1113_U44;
  assign new_P2_R1113_U385 = ~new_P2_R1113_U155 | ~new_P2_R1113_U193;
  assign new_P2_R1113_U386 = ~new_P2_U3960 | ~new_P2_R1113_U157;
  assign new_P2_R1113_U387 = ~new_P2_U3057 | ~new_P2_R1113_U156;
  assign new_P2_R1113_U388 = ~new_P2_U3960 | ~new_P2_R1113_U157;
  assign new_P2_R1113_U389 = ~new_P2_U3057 | ~new_P2_R1113_U156;
  assign new_P2_R1113_U390 = ~new_P2_R1113_U389 | ~new_P2_R1113_U388;
  assign new_P2_R1113_U391 = ~new_P2_U3949 | ~new_P2_R1113_U86;
  assign new_P2_R1113_U392 = ~new_P2_U3056 | ~new_P2_R1113_U85;
  assign new_P2_R1113_U393 = ~new_P2_R1113_U131;
  assign new_P2_R1113_U394 = ~new_P2_R1113_U393 | ~new_P2_R1113_U305;
  assign new_P2_R1113_U395 = ~new_P2_R1113_U131 | ~new_P2_R1113_U87;
  assign new_P2_R1113_U396 = ~new_P2_U3950 | ~new_P2_R1113_U84;
  assign new_P2_R1113_U397 = ~new_P2_U3055 | ~new_P2_R1113_U81;
  assign new_P2_R1113_U398 = ~new_P2_U3950 | ~new_P2_R1113_U84;
  assign new_P2_R1113_U399 = ~new_P2_U3055 | ~new_P2_R1113_U81;
  assign new_P2_R1113_U400 = ~new_P2_R1113_U399 | ~new_P2_R1113_U398;
  assign new_P2_R1113_U401 = ~new_P2_U3951 | ~new_P2_R1113_U82;
  assign new_P2_R1113_U402 = ~new_P2_U3059 | ~new_P2_R1113_U45;
  assign new_P2_R1113_U403 = ~new_P2_R1113_U317 | ~new_P2_R1113_U88;
  assign new_P2_R1113_U404 = ~new_P2_R1113_U158 | ~new_P2_R1113_U299;
  assign new_P2_R1113_U405 = ~new_P2_U3952 | ~new_P2_R1113_U80;
  assign new_P2_R1113_U406 = ~new_P2_U3060 | ~new_P2_R1113_U79;
  assign new_P2_R1113_U407 = ~new_P2_R1113_U134;
  assign new_P2_R1113_U408 = ~new_P2_R1113_U295 | ~new_P2_R1113_U407;
  assign new_P2_R1113_U409 = ~new_P2_R1113_U134 | ~new_P2_R1113_U159;
  assign new_P2_R1113_U410 = ~new_P2_U3953 | ~new_P2_R1113_U78;
  assign new_P2_R1113_U411 = ~new_P2_U3067 | ~new_P2_R1113_U77;
  assign new_P2_R1113_U412 = ~new_P2_R1113_U135;
  assign new_P2_R1113_U413 = ~new_P2_R1113_U291 | ~new_P2_R1113_U412;
  assign new_P2_R1113_U414 = ~new_P2_R1113_U135 | ~new_P2_R1113_U160;
  assign new_P2_R1113_U415 = ~new_P2_U3954 | ~new_P2_R1113_U73;
  assign new_P2_R1113_U416 = ~new_P2_U3068 | ~new_P2_R1113_U70;
  assign new_P2_R1113_U417 = ~new_P2_R1113_U416 | ~new_P2_R1113_U415;
  assign new_P2_R1113_U418 = ~new_P2_U3955 | ~new_P2_R1113_U74;
  assign new_P2_R1113_U419 = ~new_P2_U3063 | ~new_P2_R1113_U71;
  assign new_P2_R1113_U420 = ~new_P2_R1113_U327 | ~new_P2_R1113_U89;
  assign new_P2_R1113_U421 = ~new_P2_R1113_U161 | ~new_P2_R1113_U319;
  assign new_P2_R1113_U422 = ~new_P2_U3956 | ~new_P2_R1113_U75;
  assign new_P2_R1113_U423 = ~new_P2_U3077 | ~new_P2_R1113_U72;
  assign new_P2_R1113_U424 = ~new_P2_R1113_U328 | ~new_P2_R1113_U163;
  assign new_P2_R1113_U425 = ~new_P2_R1113_U281 | ~new_P2_R1113_U162;
  assign new_P2_R1113_U426 = ~new_P2_U3957 | ~new_P2_R1113_U69;
  assign new_P2_R1113_U427 = ~new_P2_U3078 | ~new_P2_R1113_U68;
  assign new_P2_R1113_U428 = ~new_P2_R1113_U138;
  assign new_P2_R1113_U429 = ~new_P2_R1113_U277 | ~new_P2_R1113_U428;
  assign new_P2_R1113_U430 = ~new_P2_R1113_U138 | ~new_P2_R1113_U164;
  assign new_P2_R1113_U431 = ~new_P2_U3432 | ~new_P2_R1113_U25;
  assign new_P2_R1113_U432 = ~new_P2_U3080 | ~new_P2_R1113_U165;
  assign new_P2_R1113_U433 = ~new_P2_R1113_U139;
  assign new_P2_R1113_U434 = ~new_P2_R1113_U191 | ~new_P2_R1113_U433;
  assign new_P2_R1113_U435 = ~new_P2_R1113_U139 | ~new_P2_R1113_U166;
  assign new_P2_R1113_U436 = ~new_P2_U3485 | ~new_P2_R1113_U67;
  assign new_P2_R1113_U437 = ~new_P2_U3083 | ~new_P2_R1113_U66;
  assign new_P2_R1113_U438 = ~new_P2_R1113_U140;
  assign new_P2_R1113_U439 = ~new_P2_R1113_U273 | ~new_P2_R1113_U438;
  assign new_P2_R1113_U440 = ~new_P2_R1113_U140 | ~new_P2_R1113_U167;
  assign new_P2_R1113_U441 = ~new_P2_U3483 | ~new_P2_R1113_U65;
  assign new_P2_R1113_U442 = ~new_P2_U3084 | ~new_P2_R1113_U168;
  assign new_P2_R1113_U443 = ~new_P2_R1113_U141;
  assign new_P2_R1113_U444 = ~new_P2_R1113_U443 | ~new_P2_R1113_U269;
  assign new_P2_R1113_U445 = ~new_P2_R1113_U141 | ~new_P2_R1113_U64;
  assign new_P2_R1113_U446 = ~new_P2_U3480 | ~new_P2_R1113_U63;
  assign new_P2_R1113_U447 = ~new_P2_U3071 | ~new_P2_R1113_U62;
  assign new_P2_R1113_U448 = ~new_P2_R1113_U142;
  assign new_P2_R1113_U449 = ~new_P2_R1113_U265 | ~new_P2_R1113_U448;
  assign new_P2_R1113_U450 = ~new_P2_R1113_U142 | ~new_P2_R1113_U169;
  assign new_P2_R1113_U451 = ~new_P2_U3477 | ~new_P2_R1113_U58;
  assign new_P2_R1113_U452 = ~new_P2_U3075 | ~new_P2_R1113_U55;
  assign new_P2_R1113_U453 = ~new_P2_R1113_U452 | ~new_P2_R1113_U451;
  assign new_P2_R1113_U454 = ~new_P2_U3474 | ~new_P2_R1113_U59;
  assign new_P2_R1113_U455 = ~new_P2_U3076 | ~new_P2_R1113_U56;
  assign new_P2_R1113_U456 = ~new_P2_R1113_U338 | ~new_P2_R1113_U90;
  assign new_P2_R1113_U457 = ~new_P2_R1113_U170 | ~new_P2_R1113_U330;
  assign new_P2_R1113_U458 = ~new_P2_U3471 | ~new_P2_R1113_U60;
  assign new_P2_R1113_U459 = ~new_P2_U3081 | ~new_P2_R1113_U57;
  assign new_P2_R1113_U460 = ~new_P2_R1113_U339 | ~new_P2_R1113_U172;
  assign new_P2_R1113_U461 = ~new_P2_R1113_U255 | ~new_P2_R1113_U171;
  assign new_P2_R1113_U462 = ~new_P2_U3468 | ~new_P2_R1113_U54;
  assign new_P2_R1113_U463 = ~new_P2_U3082 | ~new_P2_R1113_U53;
  assign new_P2_R1113_U464 = ~new_P2_R1113_U145;
  assign new_P2_R1113_U465 = ~new_P2_R1113_U251 | ~new_P2_R1113_U464;
  assign new_P2_R1113_U466 = ~new_P2_R1113_U145 | ~new_P2_R1113_U173;
  assign new_P2_R1113_U467 = ~new_P2_U3465 | ~new_P2_R1113_U52;
  assign new_P2_R1113_U468 = ~new_P2_U3074 | ~new_P2_R1113_U51;
  assign new_P2_R1113_U469 = ~new_P2_R1113_U146;
  assign new_P2_R1113_U470 = ~new_P2_R1113_U247 | ~new_P2_R1113_U469;
  assign new_P2_R1113_U471 = ~new_P2_R1113_U146 | ~new_P2_R1113_U174;
  assign new_P2_R1113_U472 = ~new_P2_U3462 | ~new_P2_R1113_U48;
  assign new_P2_R1113_U473 = ~new_P2_U3065 | ~new_P2_R1113_U47;
  assign new_P2_R1113_U474 = ~new_P2_R1113_U473 | ~new_P2_R1113_U472;
  assign new_P2_R1113_U475 = ~new_P2_U3459 | ~new_P2_R1113_U49;
  assign new_P2_R1113_U476 = ~new_P2_U3064 | ~new_P2_R1113_U46;
  assign new_P2_R1113_U477 = ~new_P2_R1113_U349 | ~new_P2_R1113_U91;
  assign new_P2_R1113_U478 = ~new_P2_R1113_U175 | ~new_P2_R1113_U341;
  assign new_P3_SUB_598_U6 = ~P3_IR_REG_18_ & ~P3_IR_REG_17_ & ~P3_IR_REG_19_ & ~P3_IR_REG_20_;
  assign new_P3_SUB_598_U7 = new_P3_SUB_598_U136 & new_P3_SUB_598_U49;
  assign new_P3_SUB_598_U8 = new_P3_SUB_598_U134 & new_P3_SUB_598_U102;
  assign new_P3_SUB_598_U9 = new_P3_SUB_598_U133 & new_P3_SUB_598_U46;
  assign new_P3_SUB_598_U10 = new_P3_SUB_598_U132 & new_P3_SUB_598_U47;
  assign new_P3_SUB_598_U11 = new_P3_SUB_598_U130 & new_P3_SUB_598_U105;
  assign new_P3_SUB_598_U12 = new_P3_SUB_598_U129 & new_P3_SUB_598_U34;
  assign new_P3_SUB_598_U13 = new_P3_SUB_598_U128 & new_P3_SUB_598_U44;
  assign new_P3_SUB_598_U14 = new_P3_SUB_598_U126 & new_P3_SUB_598_U108;
  assign new_P3_SUB_598_U15 = new_P3_SUB_598_U125 & new_P3_SUB_598_U40;
  assign new_P3_SUB_598_U16 = new_P3_SUB_598_U124 & new_P3_SUB_598_U41;
  assign new_P3_SUB_598_U17 = new_P3_SUB_598_U122 & new_P3_SUB_598_U111;
  assign new_P3_SUB_598_U18 = new_P3_SUB_598_U121 & new_P3_SUB_598_U35;
  assign new_P3_SUB_598_U19 = new_P3_SUB_598_U120 & new_P3_SUB_598_U78;
  assign new_P3_SUB_598_U20 = new_P3_SUB_598_U65 & new_P3_SUB_598_U139;
  assign new_P3_SUB_598_U21 = new_P3_SUB_598_U118 & new_P3_SUB_598_U37;
  assign new_P3_SUB_598_U22 = new_P3_SUB_598_U117 & new_P3_SUB_598_U28;
  assign new_P3_SUB_598_U23 = new_P3_SUB_598_U100 & new_P3_SUB_598_U90;
  assign new_P3_SUB_598_U24 = new_P3_SUB_598_U99 & new_P3_SUB_598_U30;
  assign new_P3_SUB_598_U25 = new_P3_SUB_598_U98 & new_P3_SUB_598_U31;
  assign new_P3_SUB_598_U26 = new_P3_SUB_598_U96 & new_P3_SUB_598_U93;
  assign new_P3_SUB_598_U27 = new_P3_SUB_598_U95 & new_P3_SUB_598_U29;
  assign new_P3_SUB_598_U28 = P3_IR_REG_2_ | P3_IR_REG_1_ | P3_IR_REG_0_;
  assign new_P3_SUB_598_U29 = ~new_P3_SUB_598_U53 | ~new_P3_SUB_598_U54 | ~new_P3_SUB_598_U140;
  assign new_P3_SUB_598_U30 = ~new_P3_SUB_598_U55 | ~new_P3_SUB_598_U140;
  assign new_P3_SUB_598_U31 = ~new_P3_SUB_598_U56 | ~new_P3_SUB_598_U91;
  assign new_P3_SUB_598_U32 = ~P3_IR_REG_7_;
  assign new_P3_SUB_598_U33 = ~P3_IR_REG_3_;
  assign new_P3_SUB_598_U34 = ~new_P3_SUB_598_U57 | ~new_P3_SUB_598_U58 | ~new_P3_SUB_598_U60 | ~new_P3_SUB_598_U59;
  assign new_P3_SUB_598_U35 = ~new_P3_SUB_598_U62 | ~new_P3_SUB_598_U106;
  assign new_P3_SUB_598_U36 = ~new_P3_SUB_598_U63 | ~new_P3_SUB_598_U112;
  assign new_P3_SUB_598_U37 = ~new_P3_SUB_598_U114 | ~new_P3_SUB_598_U38;
  assign new_P3_SUB_598_U38 = ~P3_IR_REG_29_;
  assign new_P3_SUB_598_U39 = ~P3_IR_REG_27_;
  assign new_P3_SUB_598_U40 = ~new_P3_SUB_598_U106 | ~new_P3_SUB_598_U6;
  assign new_P3_SUB_598_U41 = ~new_P3_SUB_598_U66 | ~new_P3_SUB_598_U109;
  assign new_P3_SUB_598_U42 = ~P3_IR_REG_24_;
  assign new_P3_SUB_598_U43 = ~P3_IR_REG_23_;
  assign new_P3_SUB_598_U44 = ~new_P3_SUB_598_U67 | ~new_P3_SUB_598_U106;
  assign new_P3_SUB_598_U45 = ~P3_IR_REG_19_;
  assign new_P3_SUB_598_U46 = ~new_P3_SUB_598_U68 | ~new_P3_SUB_598_U94;
  assign new_P3_SUB_598_U47 = ~new_P3_SUB_598_U69 | ~new_P3_SUB_598_U103;
  assign new_P3_SUB_598_U48 = ~P3_IR_REG_15_;
  assign new_P3_SUB_598_U49 = ~new_P3_SUB_598_U70 | ~new_P3_SUB_598_U94;
  assign new_P3_SUB_598_U50 = ~P3_IR_REG_11_;
  assign new_P3_SUB_598_U51 = ~new_P3_SUB_598_U156 | ~new_P3_SUB_598_U155;
  assign new_P3_SUB_598_U52 = ~new_P3_SUB_598_U146 | ~new_P3_SUB_598_U145;
  assign new_P3_SUB_598_U53 = ~P3_IR_REG_6_ & ~P3_IR_REG_5_ & ~P3_IR_REG_3_ & ~P3_IR_REG_4_;
  assign new_P3_SUB_598_U54 = ~P3_IR_REG_7_ & ~P3_IR_REG_8_;
  assign new_P3_SUB_598_U55 = ~P3_IR_REG_3_ & ~P3_IR_REG_4_;
  assign new_P3_SUB_598_U56 = ~P3_IR_REG_5_ & ~P3_IR_REG_6_;
  assign new_P3_SUB_598_U57 = ~P3_IR_REG_11_ & ~P3_IR_REG_10_ & ~P3_IR_REG_12_ & ~P3_IR_REG_13_ & ~P3_IR_REG_14_;
  assign new_P3_SUB_598_U58 = ~P3_IR_REG_0_ & ~P3_IR_REG_1_ & ~P3_IR_REG_15_ & ~P3_IR_REG_16_;
  assign new_P3_SUB_598_U59 = ~P3_IR_REG_5_ & ~P3_IR_REG_4_ & ~P3_IR_REG_2_ & ~P3_IR_REG_3_;
  assign new_P3_SUB_598_U60 = ~P3_IR_REG_9_ & ~P3_IR_REG_8_ & ~P3_IR_REG_6_ & ~P3_IR_REG_7_;
  assign new_P3_SUB_598_U61 = ~P3_IR_REG_22_ & ~P3_IR_REG_23_ & ~P3_IR_REG_21_;
  assign new_P3_SUB_598_U62 = new_P3_SUB_598_U61 & new_P3_SUB_598_U6 & new_P3_SUB_598_U42;
  assign new_P3_SUB_598_U63 = ~P3_IR_REG_28_ & ~P3_IR_REG_27_ & ~P3_IR_REG_25_ & ~P3_IR_REG_26_;
  assign new_P3_SUB_598_U64 = ~P3_IR_REG_25_ & ~P3_IR_REG_26_;
  assign new_P3_SUB_598_U65 = new_P3_SUB_598_U138 & new_P3_SUB_598_U36;
  assign new_P3_SUB_598_U66 = ~P3_IR_REG_21_ & ~P3_IR_REG_22_;
  assign new_P3_SUB_598_U67 = ~P3_IR_REG_17_ & ~P3_IR_REG_18_;
  assign new_P3_SUB_598_U68 = ~P3_IR_REG_9_ & ~P3_IR_REG_12_ & ~P3_IR_REG_10_ & ~P3_IR_REG_11_;
  assign new_P3_SUB_598_U69 = ~P3_IR_REG_13_ & ~P3_IR_REG_14_;
  assign new_P3_SUB_598_U70 = ~P3_IR_REG_10_ & ~P3_IR_REG_9_;
  assign new_P3_SUB_598_U71 = ~P3_IR_REG_9_;
  assign new_P3_SUB_598_U72 = new_P3_SUB_598_U142 & new_P3_SUB_598_U141;
  assign new_P3_SUB_598_U73 = ~P3_IR_REG_5_;
  assign new_P3_SUB_598_U74 = new_P3_SUB_598_U144 & new_P3_SUB_598_U143;
  assign new_P3_SUB_598_U75 = ~P3_IR_REG_31_;
  assign new_P3_SUB_598_U76 = ~P3_IR_REG_30_;
  assign new_P3_SUB_598_U77 = new_P3_SUB_598_U148 & new_P3_SUB_598_U147;
  assign new_P3_SUB_598_U78 = ~new_P3_SUB_598_U64 | ~new_P3_SUB_598_U112;
  assign new_P3_SUB_598_U79 = new_P3_SUB_598_U150 & new_P3_SUB_598_U149;
  assign new_P3_SUB_598_U80 = ~P3_IR_REG_25_;
  assign new_P3_SUB_598_U81 = new_P3_SUB_598_U152 & new_P3_SUB_598_U151;
  assign new_P3_SUB_598_U82 = ~P3_IR_REG_21_;
  assign new_P3_SUB_598_U83 = new_P3_SUB_598_U154 & new_P3_SUB_598_U153;
  assign new_P3_SUB_598_U84 = ~P3_IR_REG_1_;
  assign new_P3_SUB_598_U85 = ~P3_IR_REG_0_;
  assign new_P3_SUB_598_U86 = ~P3_IR_REG_17_;
  assign new_P3_SUB_598_U87 = new_P3_SUB_598_U158 & new_P3_SUB_598_U157;
  assign new_P3_SUB_598_U88 = ~P3_IR_REG_13_;
  assign new_P3_SUB_598_U89 = new_P3_SUB_598_U160 & new_P3_SUB_598_U159;
  assign new_P3_SUB_598_U90 = ~new_P3_SUB_598_U140 | ~new_P3_SUB_598_U33;
  assign new_P3_SUB_598_U91 = ~new_P3_SUB_598_U30;
  assign new_P3_SUB_598_U92 = ~new_P3_SUB_598_U31;
  assign new_P3_SUB_598_U93 = ~new_P3_SUB_598_U92 | ~new_P3_SUB_598_U32;
  assign new_P3_SUB_598_U94 = ~new_P3_SUB_598_U29;
  assign new_P3_SUB_598_U95 = ~P3_IR_REG_8_ | ~new_P3_SUB_598_U93;
  assign new_P3_SUB_598_U96 = ~P3_IR_REG_7_ | ~new_P3_SUB_598_U31;
  assign new_P3_SUB_598_U97 = ~new_P3_SUB_598_U91 | ~new_P3_SUB_598_U73;
  assign new_P3_SUB_598_U98 = ~P3_IR_REG_6_ | ~new_P3_SUB_598_U97;
  assign new_P3_SUB_598_U99 = ~P3_IR_REG_4_ | ~new_P3_SUB_598_U90;
  assign new_P3_SUB_598_U100 = ~P3_IR_REG_3_ | ~new_P3_SUB_598_U28;
  assign new_P3_SUB_598_U101 = ~new_P3_SUB_598_U49;
  assign new_P3_SUB_598_U102 = ~new_P3_SUB_598_U101 | ~new_P3_SUB_598_U50;
  assign new_P3_SUB_598_U103 = ~new_P3_SUB_598_U46;
  assign new_P3_SUB_598_U104 = ~new_P3_SUB_598_U47;
  assign new_P3_SUB_598_U105 = ~new_P3_SUB_598_U104 | ~new_P3_SUB_598_U48;
  assign new_P3_SUB_598_U106 = ~new_P3_SUB_598_U34;
  assign new_P3_SUB_598_U107 = ~new_P3_SUB_598_U44;
  assign new_P3_SUB_598_U108 = ~new_P3_SUB_598_U107 | ~new_P3_SUB_598_U45;
  assign new_P3_SUB_598_U109 = ~new_P3_SUB_598_U40;
  assign new_P3_SUB_598_U110 = ~new_P3_SUB_598_U41;
  assign new_P3_SUB_598_U111 = ~new_P3_SUB_598_U110 | ~new_P3_SUB_598_U43;
  assign new_P3_SUB_598_U112 = ~new_P3_SUB_598_U35;
  assign new_P3_SUB_598_U113 = ~new_P3_SUB_598_U78;
  assign new_P3_SUB_598_U114 = ~new_P3_SUB_598_U36;
  assign new_P3_SUB_598_U115 = ~new_P3_SUB_598_U37;
  assign new_P3_SUB_598_U116 = P3_IR_REG_1_ | P3_IR_REG_0_;
  assign new_P3_SUB_598_U117 = ~P3_IR_REG_2_ | ~new_P3_SUB_598_U116;
  assign new_P3_SUB_598_U118 = ~P3_IR_REG_29_ | ~new_P3_SUB_598_U36;
  assign new_P3_SUB_598_U119 = ~new_P3_SUB_598_U112 | ~new_P3_SUB_598_U80;
  assign new_P3_SUB_598_U120 = ~P3_IR_REG_26_ | ~new_P3_SUB_598_U119;
  assign new_P3_SUB_598_U121 = ~P3_IR_REG_24_ | ~new_P3_SUB_598_U111;
  assign new_P3_SUB_598_U122 = ~P3_IR_REG_23_ | ~new_P3_SUB_598_U41;
  assign new_P3_SUB_598_U123 = ~new_P3_SUB_598_U109 | ~new_P3_SUB_598_U82;
  assign new_P3_SUB_598_U124 = ~P3_IR_REG_22_ | ~new_P3_SUB_598_U123;
  assign new_P3_SUB_598_U125 = ~P3_IR_REG_20_ | ~new_P3_SUB_598_U108;
  assign new_P3_SUB_598_U126 = ~P3_IR_REG_19_ | ~new_P3_SUB_598_U44;
  assign new_P3_SUB_598_U127 = ~new_P3_SUB_598_U106 | ~new_P3_SUB_598_U86;
  assign new_P3_SUB_598_U128 = ~P3_IR_REG_18_ | ~new_P3_SUB_598_U127;
  assign new_P3_SUB_598_U129 = ~P3_IR_REG_16_ | ~new_P3_SUB_598_U105;
  assign new_P3_SUB_598_U130 = ~P3_IR_REG_15_ | ~new_P3_SUB_598_U47;
  assign new_P3_SUB_598_U131 = ~new_P3_SUB_598_U103 | ~new_P3_SUB_598_U88;
  assign new_P3_SUB_598_U132 = ~P3_IR_REG_14_ | ~new_P3_SUB_598_U131;
  assign new_P3_SUB_598_U133 = ~P3_IR_REG_12_ | ~new_P3_SUB_598_U102;
  assign new_P3_SUB_598_U134 = ~P3_IR_REG_11_ | ~new_P3_SUB_598_U49;
  assign new_P3_SUB_598_U135 = ~new_P3_SUB_598_U94 | ~new_P3_SUB_598_U71;
  assign new_P3_SUB_598_U136 = ~P3_IR_REG_10_ | ~new_P3_SUB_598_U135;
  assign new_P3_SUB_598_U137 = ~new_P3_SUB_598_U115 | ~new_P3_SUB_598_U76;
  assign new_P3_SUB_598_U138 = ~P3_IR_REG_27_ | ~P3_IR_REG_28_;
  assign new_P3_SUB_598_U139 = ~P3_IR_REG_28_ | ~new_P3_SUB_598_U78;
  assign new_P3_SUB_598_U140 = ~new_P3_SUB_598_U28;
  assign new_P3_SUB_598_U141 = ~P3_IR_REG_9_ | ~new_P3_SUB_598_U29;
  assign new_P3_SUB_598_U142 = ~new_P3_SUB_598_U94 | ~new_P3_SUB_598_U71;
  assign new_P3_SUB_598_U143 = ~P3_IR_REG_5_ | ~new_P3_SUB_598_U30;
  assign new_P3_SUB_598_U144 = ~new_P3_SUB_598_U91 | ~new_P3_SUB_598_U73;
  assign new_P3_SUB_598_U145 = ~new_P3_SUB_598_U137 | ~new_P3_SUB_598_U75;
  assign new_P3_SUB_598_U146 = ~P3_IR_REG_31_ | ~new_P3_SUB_598_U115 | ~new_P3_SUB_598_U76;
  assign new_P3_SUB_598_U147 = ~P3_IR_REG_30_ | ~new_P3_SUB_598_U37;
  assign new_P3_SUB_598_U148 = ~new_P3_SUB_598_U115 | ~new_P3_SUB_598_U76;
  assign new_P3_SUB_598_U149 = ~P3_IR_REG_27_ | ~new_P3_SUB_598_U78;
  assign new_P3_SUB_598_U150 = ~new_P3_SUB_598_U113 | ~new_P3_SUB_598_U39;
  assign new_P3_SUB_598_U151 = ~P3_IR_REG_25_ | ~new_P3_SUB_598_U35;
  assign new_P3_SUB_598_U152 = ~new_P3_SUB_598_U112 | ~new_P3_SUB_598_U80;
  assign new_P3_SUB_598_U153 = ~P3_IR_REG_21_ | ~new_P3_SUB_598_U40;
  assign new_P3_SUB_598_U154 = ~new_P3_SUB_598_U109 | ~new_P3_SUB_598_U82;
  assign new_P3_SUB_598_U155 = ~P3_IR_REG_1_ | ~new_P3_SUB_598_U85;
  assign new_P3_SUB_598_U156 = ~P3_IR_REG_0_ | ~new_P3_SUB_598_U84;
  assign new_P3_SUB_598_U157 = ~P3_IR_REG_17_ | ~new_P3_SUB_598_U34;
  assign new_P3_SUB_598_U158 = ~new_P3_SUB_598_U106 | ~new_P3_SUB_598_U86;
  assign new_P3_SUB_598_U159 = ~P3_IR_REG_13_ | ~new_P3_SUB_598_U46;
  assign new_P3_SUB_598_U160 = ~new_P3_SUB_598_U103 | ~new_P3_SUB_598_U88;
  assign new_P3_R693_U6 = new_P3_R693_U113 & new_P3_R693_U114;
  assign new_P3_R693_U7 = new_P3_R693_U115 & new_P3_R693_U116;
  assign new_P3_R693_U8 = new_P3_R693_U7 & new_P3_R693_U120 & new_P3_R693_U80 & new_P3_R693_U118;
  assign new_P3_R693_U9 = new_P3_R693_U126 & new_P3_R693_U125;
  assign new_P3_R693_U10 = new_P3_R693_U130 & new_P3_R693_U131;
  assign new_P3_R693_U11 = new_P3_R693_U84 & new_P3_R693_U10;
  assign new_P3_R693_U12 = new_P3_R693_U142 & new_P3_R693_U141;
  assign new_P3_R693_U13 = new_P3_R693_U177 & new_P3_R693_U178 & new_P3_R693_U179;
  assign new_P3_R693_U14 = new_P3_R693_U109 & new_P3_R693_U108 & new_P3_R693_U189 & new_P3_R693_U188;
  assign new_P3_R693_U15 = ~new_P3_U3529;
  assign new_P3_R693_U16 = ~new_P3_U3537;
  assign new_P3_R693_U17 = ~new_P3_U3536;
  assign new_P3_R693_U18 = ~new_P3_U3905;
  assign new_P3_R693_U19 = ~new_P3_U3540;
  assign new_P3_R693_U20 = ~new_P3_U3906;
  assign new_P3_R693_U21 = ~new_P3_U3541;
  assign new_P3_R693_U22 = ~new_P3_U3543;
  assign new_P3_R693_U23 = ~new_P3_U3443;
  assign new_P3_R693_U24 = ~new_P3_U3544;
  assign new_P3_R693_U25 = ~new_P3_U3440;
  assign new_P3_R693_U26 = ~new_P3_U3445;
  assign new_P3_R693_U27 = ~new_P3_U3907;
  assign new_P3_R693_U28 = ~new_P3_U3545;
  assign new_P3_R693_U29 = ~new_P3_U3546;
  assign new_P3_R693_U30 = ~new_P3_U3437;
  assign new_P3_R693_U31 = ~new_P3_U3434;
  assign new_P3_R693_U32 = ~new_P3_U3526;
  assign new_P3_R693_U33 = ~new_P3_U3525;
  assign new_P3_R693_U34 = ~new_P3_U3404;
  assign new_P3_R693_U35 = ~new_P3_U3407;
  assign new_P3_R693_U36 = ~new_P3_U3416;
  assign new_P3_R693_U37 = ~new_P3_U3419;
  assign new_P3_R693_U38 = ~new_P3_U3410;
  assign new_P3_R693_U39 = ~new_P3_U3413;
  assign new_P3_R693_U40 = ~new_P3_U3398;
  assign new_P3_R693_U41 = ~new_P3_U3401;
  assign new_P3_R693_U42 = ~new_P3_U3553;
  assign new_P3_R693_U43 = ~new_P3_U3395;
  assign new_P3_R693_U44 = ~new_P3_U3392;
  assign new_P3_R693_U45 = ~new_P3_U3550;
  assign new_P3_R693_U46 = ~new_P3_U3549;
  assign new_P3_R693_U47 = ~new_P3_U3542;
  assign new_P3_R693_U48 = ~new_P3_U3531;
  assign new_P3_R693_U49 = ~new_P3_U3528;
  assign new_P3_R693_U50 = ~new_P3_U3527;
  assign new_P3_R693_U51 = ~new_P3_U3523;
  assign new_P3_R693_U52 = ~new_P3_U3524;
  assign new_P3_R693_U53 = ~new_P3_U3552;
  assign new_P3_R693_U54 = ~new_P3_U3551;
  assign new_P3_R693_U55 = ~new_P3_U3425;
  assign new_P3_R693_U56 = ~new_P3_U3422;
  assign new_P3_R693_U57 = ~new_P3_U3431;
  assign new_P3_R693_U58 = ~new_P3_U3428;
  assign new_P3_R693_U59 = ~new_P3_U3548;
  assign new_P3_R693_U60 = ~new_P3_U3547;
  assign new_P3_R693_U61 = ~new_P3_U3539;
  assign new_P3_R693_U62 = ~new_P3_U3538;
  assign new_P3_R693_U63 = ~new_P3_U3908;
  assign new_P3_R693_U64 = ~new_P3_U3900;
  assign new_P3_R693_U65 = ~new_P3_U3899;
  assign new_P3_R693_U66 = ~new_P3_U3904;
  assign new_P3_R693_U67 = ~new_P3_U3903;
  assign new_P3_R693_U68 = ~new_P3_U3902;
  assign new_P3_R693_U69 = ~new_P3_U3901;
  assign new_P3_R693_U70 = ~new_P3_U3533;
  assign new_P3_R693_U71 = ~new_P3_U3534;
  assign new_P3_R693_U72 = ~new_P3_U3872;
  assign new_P3_R693_U73 = ~new_P3_U3532;
  assign new_P3_R693_U74 = ~new_P3_U3535;
  assign new_P3_R693_U75 = new_P3_U3540 & new_P3_R693_U20;
  assign new_P3_R693_U76 = new_P3_U3541 & new_P3_R693_U27;
  assign new_P3_R693_U77 = new_P3_R693_U168 & new_P3_R693_U167;
  assign new_P3_R693_U78 = new_P3_U3443 & new_P3_R693_U24;
  assign new_P3_R693_U79 = new_P3_U3440 & new_P3_R693_U28;
  assign new_P3_R693_U80 = new_P3_R693_U119 & new_P3_R693_U117;
  assign new_P3_R693_U81 = new_P3_U3404 & new_P3_R693_U50;
  assign new_P3_R693_U82 = new_P3_U3407 & new_P3_R693_U32;
  assign new_P3_R693_U83 = new_P3_U3387 & new_P3_R693_U111;
  assign new_P3_R693_U84 = new_P3_R693_U133 & new_P3_R693_U132;
  assign new_P3_R693_U85 = new_P3_R693_U129 & new_P3_R693_U86;
  assign new_P3_R693_U86 = new_P3_R693_U135 & new_P3_R693_U134;
  assign new_P3_R693_U87 = new_P3_R693_U138 & new_P3_R693_U137;
  assign new_P3_R693_U88 = new_P3_R693_U135 & new_P3_R693_U134;
  assign new_P3_R693_U89 = new_P3_R693_U9 & new_P3_R693_U148;
  assign new_P3_R693_U90 = new_P3_R693_U11 & new_P3_R693_U129 & new_P3_R693_U127;
  assign new_P3_R693_U91 = new_P3_U3523 & new_P3_R693_U36;
  assign new_P3_R693_U92 = new_P3_U3524 & new_P3_R693_U39;
  assign new_P3_R693_U93 = new_P3_R693_U95 & new_P3_R693_U152 & new_P3_R693_U151;
  assign new_P3_R693_U94 = new_P3_R693_U154 & new_P3_R693_U153;
  assign new_P3_R693_U95 = new_P3_R693_U94 & new_P3_R693_U12;
  assign new_P3_R693_U96 = new_P3_U3425 & new_P3_R693_U45;
  assign new_P3_R693_U97 = new_P3_U3422 & new_P3_R693_U54;
  assign new_P3_R693_U98 = new_P3_R693_U157 & new_P3_R693_U100;
  assign new_P3_R693_U99 = new_P3_R693_U98 & new_P3_R693_U158;
  assign new_P3_R693_U100 = new_P3_R693_U160 & new_P3_R693_U159;
  assign new_P3_R693_U101 = new_P3_R693_U123 & new_P3_R693_U122 & new_P3_R693_U171 & new_P3_R693_U170;
  assign new_P3_R693_U102 = new_P3_R693_U175 & new_P3_R693_U174;
  assign new_P3_R693_U103 = new_P3_R693_U187 & new_P3_R693_U186;
  assign new_P3_R693_U104 = new_P3_R693_U103 & new_P3_R693_U13;
  assign new_P3_R693_U105 = new_P3_R693_U106 & new_P3_R693_U190;
  assign new_P3_R693_U106 = new_P3_U3533 & new_P3_R693_U65;
  assign new_P3_R693_U107 = new_P3_U3532 & new_P3_R693_U63;
  assign new_P3_R693_U108 = new_P3_R693_U192 & new_P3_R693_U191;
  assign new_P3_R693_U109 = new_P3_R693_U195 & new_P3_R693_U194 & new_P3_R693_U193;
  assign new_P3_R693_U110 = ~new_P3_U3873;
  assign new_P3_R693_U111 = ~new_P3_U3554;
  assign new_P3_R693_U112 = ~new_P3_R693_U181 | ~new_P3_R693_U196;
  assign new_P3_R693_U113 = ~new_P3_U3543 | ~new_P3_R693_U26;
  assign new_P3_R693_U114 = ~new_P3_U3544 | ~new_P3_R693_U23;
  assign new_P3_R693_U115 = ~new_P3_U3905 | ~new_P3_R693_U61;
  assign new_P3_R693_U116 = ~new_P3_U3906 | ~new_P3_R693_U19;
  assign new_P3_R693_U117 = ~new_P3_R693_U78 | ~new_P3_R693_U113;
  assign new_P3_R693_U118 = ~new_P3_R693_U79 | ~new_P3_R693_U6;
  assign new_P3_R693_U119 = ~new_P3_U3445 | ~new_P3_R693_U22;
  assign new_P3_R693_U120 = ~new_P3_U3907 | ~new_P3_R693_U21;
  assign new_P3_R693_U121 = ~new_P3_U3437 | ~new_P3_R693_U29;
  assign new_P3_R693_U122 = ~new_P3_U3537 | ~new_P3_R693_U67;
  assign new_P3_R693_U123 = ~new_P3_U3536 | ~new_P3_R693_U68;
  assign new_P3_R693_U124 = ~new_P3_U3434 | ~new_P3_R693_U60;
  assign new_P3_R693_U125 = ~new_P3_U3526 | ~new_P3_R693_U35;
  assign new_P3_R693_U126 = ~new_P3_U3525 | ~new_P3_R693_U38;
  assign new_P3_R693_U127 = ~new_P3_R693_U81 | ~new_P3_R693_U9;
  assign new_P3_R693_U128 = ~new_P3_U3525 | ~new_P3_R693_U38;
  assign new_P3_R693_U129 = ~new_P3_R693_U82 | ~new_P3_R693_U128;
  assign new_P3_R693_U130 = ~new_P3_U3419 | ~new_P3_R693_U53;
  assign new_P3_R693_U131 = ~new_P3_U3416 | ~new_P3_R693_U51;
  assign new_P3_R693_U132 = ~new_P3_U3410 | ~new_P3_R693_U33;
  assign new_P3_R693_U133 = ~new_P3_U3413 | ~new_P3_R693_U52;
  assign new_P3_R693_U134 = ~new_P3_U3398 | ~new_P3_R693_U48;
  assign new_P3_R693_U135 = ~new_P3_U3401 | ~new_P3_R693_U49;
  assign new_P3_R693_U136 = ~new_P3_U3553 | ~new_P3_R693_U44;
  assign new_P3_R693_U137 = ~new_P3_R693_U83 | ~new_P3_R693_U136;
  assign new_P3_R693_U138 = ~new_P3_U3395 | ~new_P3_R693_U47;
  assign new_P3_R693_U139 = ~new_P3_U3392 | ~new_P3_R693_U42;
  assign new_P3_R693_U140 = ~new_P3_R693_U85 | ~new_P3_R693_U127 | ~new_P3_R693_U87 | ~new_P3_R693_U11 | ~new_P3_R693_U139;
  assign new_P3_R693_U141 = ~new_P3_U3550 | ~new_P3_R693_U55;
  assign new_P3_R693_U142 = ~new_P3_U3549 | ~new_P3_R693_U58;
  assign new_P3_R693_U143 = ~new_P3_U3542 | ~new_P3_R693_U43;
  assign new_P3_R693_U144 = ~new_P3_U3531 | ~new_P3_R693_U40;
  assign new_P3_R693_U145 = ~new_P3_R693_U144 | ~new_P3_R693_U143;
  assign new_P3_R693_U146 = ~new_P3_R693_U88 | ~new_P3_R693_U145;
  assign new_P3_R693_U147 = ~new_P3_U3528 | ~new_P3_R693_U41;
  assign new_P3_R693_U148 = ~new_P3_U3527 | ~new_P3_R693_U34;
  assign new_P3_R693_U149 = ~new_P3_R693_U89 | ~new_P3_R693_U147 | ~new_P3_R693_U146;
  assign new_P3_R693_U150 = ~new_P3_R693_U90 | ~new_P3_R693_U149;
  assign new_P3_R693_U151 = ~new_P3_R693_U91 | ~new_P3_R693_U130;
  assign new_P3_R693_U152 = ~new_P3_R693_U92 | ~new_P3_R693_U10;
  assign new_P3_R693_U153 = ~new_P3_U3552 | ~new_P3_R693_U37;
  assign new_P3_R693_U154 = ~new_P3_U3551 | ~new_P3_R693_U56;
  assign new_P3_R693_U155 = ~new_P3_R693_U93 | ~new_P3_R693_U150 | ~new_P3_R693_U140;
  assign new_P3_R693_U156 = ~new_P3_U3549 | ~new_P3_R693_U58;
  assign new_P3_R693_U157 = ~new_P3_R693_U96 | ~new_P3_R693_U156;
  assign new_P3_R693_U158 = ~new_P3_R693_U97 | ~new_P3_R693_U12;
  assign new_P3_R693_U159 = ~new_P3_U3431 | ~new_P3_R693_U59;
  assign new_P3_R693_U160 = ~new_P3_U3428 | ~new_P3_R693_U46;
  assign new_P3_R693_U161 = ~new_P3_R693_U155 | ~new_P3_R693_U99;
  assign new_P3_R693_U162 = ~new_P3_U3548 | ~new_P3_R693_U57;
  assign new_P3_R693_U163 = ~new_P3_R693_U162 | ~new_P3_R693_U161;
  assign new_P3_R693_U164 = ~new_P3_R693_U163 | ~new_P3_R693_U124;
  assign new_P3_R693_U165 = ~new_P3_U3547 | ~new_P3_R693_U31;
  assign new_P3_R693_U166 = ~new_P3_R693_U165 | ~new_P3_R693_U164;
  assign new_P3_R693_U167 = ~new_P3_U3545 | ~new_P3_R693_U25;
  assign new_P3_R693_U168 = ~new_P3_U3546 | ~new_P3_R693_U30;
  assign new_P3_R693_U169 = ~new_P3_R693_U77 | ~new_P3_R693_U6;
  assign new_P3_R693_U170 = ~new_P3_R693_U75 | ~new_P3_R693_U115;
  assign new_P3_R693_U171 = ~new_P3_R693_U76 | ~new_P3_R693_U7;
  assign new_P3_R693_U172 = ~new_P3_R693_U8 | ~new_P3_R693_U169;
  assign new_P3_R693_U173 = ~new_P3_R693_U8 | ~new_P3_R693_U166 | ~new_P3_R693_U121;
  assign new_P3_R693_U174 = ~new_P3_U3539 | ~new_P3_R693_U18;
  assign new_P3_R693_U175 = ~new_P3_U3538 | ~new_P3_R693_U66;
  assign new_P3_R693_U176 = ~new_P3_R693_U101 | ~new_P3_R693_U102 | ~new_P3_R693_U173 | ~new_P3_R693_U172;
  assign new_P3_R693_U177 = ~new_P3_U3908 | ~new_P3_R693_U73;
  assign new_P3_R693_U178 = ~new_P3_U3900 | ~new_P3_R693_U71;
  assign new_P3_R693_U179 = ~new_P3_U3899 | ~new_P3_R693_U70;
  assign new_P3_R693_U180 = ~new_P3_U3529 | ~new_P3_R693_U72;
  assign new_P3_R693_U181 = ~new_P3_R693_U180 | ~new_P3_R693_U110;
  assign new_P3_R693_U182 = ~new_P3_U3904 | ~new_P3_R693_U62;
  assign new_P3_R693_U183 = ~new_P3_U3903 | ~new_P3_R693_U16;
  assign new_P3_R693_U184 = ~new_P3_R693_U183 | ~new_P3_R693_U182;
  assign new_P3_R693_U185 = ~new_P3_R693_U123 | ~new_P3_R693_U184 | ~new_P3_R693_U122;
  assign new_P3_R693_U186 = ~new_P3_U3902 | ~new_P3_R693_U17;
  assign new_P3_R693_U187 = ~new_P3_U3901 | ~new_P3_R693_U74;
  assign new_P3_R693_U188 = ~new_P3_R693_U104 | ~new_P3_R693_U112 | ~new_P3_R693_U176 | ~new_P3_R693_U185;
  assign new_P3_R693_U189 = ~new_P3_R693_U110 | ~new_P3_R693_U180 | ~new_P3_U3530;
  assign new_P3_R693_U190 = ~new_P3_U3908 | ~new_P3_R693_U73;
  assign new_P3_R693_U191 = ~new_P3_R693_U112 | ~new_P3_R693_U105;
  assign new_P3_R693_U192 = ~new_P3_R693_U64 | ~new_P3_R693_U112 | ~new_P3_U3534 | ~new_P3_R693_U13;
  assign new_P3_R693_U193 = ~new_P3_U3872 | ~new_P3_R693_U15;
  assign new_P3_R693_U194 = ~new_P3_R693_U107 | ~new_P3_R693_U112;
  assign new_P3_R693_U195 = ~new_P3_R693_U69 | ~new_P3_R693_U112 | ~new_P3_U3535 | ~new_P3_R693_U13;
  assign new_P3_R693_U196 = ~new_P3_U3530 | ~new_P3_R693_U180;
  assign new_P3_SUB_609_U6 = ~new_P3_SUB_609_U40 | ~new_P3_SUB_609_U98;
  assign new_P3_SUB_609_U7 = ~new_P3_SUB_609_U79 | ~new_P3_SUB_609_U105;
  assign new_P3_SUB_609_U8 = ~new_P3_SUB_609_U65 | ~new_P3_SUB_609_U113;
  assign new_P3_SUB_609_U9 = ~new_P3_SUB_609_U34 | ~new_P3_SUB_609_U110;
  assign new_P3_SUB_609_U10 = ~new_P3_SUB_609_U87 | ~new_P3_SUB_609_U97;
  assign new_P3_SUB_609_U11 = ~new_P3_SUB_609_U81 | ~new_P3_SUB_609_U103;
  assign new_P3_SUB_609_U12 = ~new_P3_SUB_609_U67 | ~new_P3_SUB_609_U70;
  assign new_P3_SUB_609_U13 = ~new_P3_SUB_609_U73 | ~new_P3_SUB_609_U111;
  assign new_P3_SUB_609_U14 = ~new_P3_SUB_609_U33 | ~new_P3_SUB_609_U69;
  assign new_P3_SUB_609_U15 = ~new_P3_SUB_609_U38 | ~new_P3_SUB_609_U102;
  assign new_P3_SUB_609_U16 = ~new_P3_SUB_609_U41 | ~new_P3_SUB_609_U96;
  assign new_P3_SUB_609_U17 = ~new_P3_SUB_609_U85 | ~new_P3_SUB_609_U99;
  assign new_P3_SUB_609_U18 = ~new_P3_SUB_609_U31 | ~new_P3_SUB_609_U71;
  assign new_P3_SUB_609_U19 = ~new_P3_SUB_609_U37 | ~new_P3_SUB_609_U104;
  assign new_P3_SUB_609_U20 = ~new_P3_SUB_609_U83 | ~new_P3_SUB_609_U101;
  assign new_P3_SUB_609_U21 = ~new_P3_SUB_609_U36 | ~new_P3_SUB_609_U106;
  assign new_P3_SUB_609_U22 = ~new_P3_SUB_609_U42 | ~new_P3_SUB_609_U94;
  assign new_P3_SUB_609_U23 = ~new_P3_SUB_609_U75 | ~new_P3_SUB_609_U109;
  assign new_P3_SUB_609_U24 = ~new_P3_SUB_609_U35 | ~new_P3_SUB_609_U108;
  assign new_P3_SUB_609_U25 = ~P3_REG3_REG_3_;
  assign new_P3_SUB_609_U26 = ~new_P3_SUB_609_U89 | ~new_P3_SUB_609_U95;
  assign new_P3_SUB_609_U27 = ~new_P3_SUB_609_U39 | ~new_P3_SUB_609_U100;
  assign new_P3_SUB_609_U28 = ~new_P3_SUB_609_U91 | ~new_P3_SUB_609_U93;
  assign new_P3_SUB_609_U29 = ~new_P3_SUB_609_U64 | ~new_P3_SUB_609_U72;
  assign new_P3_SUB_609_U30 = ~new_P3_SUB_609_U77 | ~new_P3_SUB_609_U107;
  assign new_P3_SUB_609_U31 = P3_REG3_REG_7_ | P3_REG3_REG_6_ | P3_REG3_REG_5_ | P3_REG3_REG_4_ | P3_REG3_REG_3_;
  assign new_P3_SUB_609_U32 = ~P3_REG3_REG_8_;
  assign new_P3_SUB_609_U33 = ~new_P3_SUB_609_U54 | ~new_P3_SUB_609_U66;
  assign new_P3_SUB_609_U34 = ~new_P3_SUB_609_U55 | ~new_P3_SUB_609_U68;
  assign new_P3_SUB_609_U35 = ~new_P3_SUB_609_U56 | ~new_P3_SUB_609_U74;
  assign new_P3_SUB_609_U36 = ~new_P3_SUB_609_U57 | ~new_P3_SUB_609_U76;
  assign new_P3_SUB_609_U37 = ~new_P3_SUB_609_U58 | ~new_P3_SUB_609_U78;
  assign new_P3_SUB_609_U38 = ~new_P3_SUB_609_U59 | ~new_P3_SUB_609_U80;
  assign new_P3_SUB_609_U39 = ~new_P3_SUB_609_U60 | ~new_P3_SUB_609_U82;
  assign new_P3_SUB_609_U40 = ~new_P3_SUB_609_U61 | ~new_P3_SUB_609_U84;
  assign new_P3_SUB_609_U41 = ~new_P3_SUB_609_U62 | ~new_P3_SUB_609_U86;
  assign new_P3_SUB_609_U42 = ~new_P3_SUB_609_U63 | ~new_P3_SUB_609_U88;
  assign new_P3_SUB_609_U43 = ~P3_REG3_REG_28_;
  assign new_P3_SUB_609_U44 = ~P3_REG3_REG_26_;
  assign new_P3_SUB_609_U45 = ~P3_REG3_REG_24_;
  assign new_P3_SUB_609_U46 = ~P3_REG3_REG_22_;
  assign new_P3_SUB_609_U47 = ~P3_REG3_REG_20_;
  assign new_P3_SUB_609_U48 = ~P3_REG3_REG_18_;
  assign new_P3_SUB_609_U49 = ~P3_REG3_REG_16_;
  assign new_P3_SUB_609_U50 = ~P3_REG3_REG_14_;
  assign new_P3_SUB_609_U51 = ~P3_REG3_REG_12_;
  assign new_P3_SUB_609_U52 = ~P3_REG3_REG_10_;
  assign new_P3_SUB_609_U53 = ~new_P3_SUB_609_U115 | ~new_P3_SUB_609_U114;
  assign new_P3_SUB_609_U54 = ~P3_REG3_REG_8_ & ~P3_REG3_REG_9_;
  assign new_P3_SUB_609_U55 = ~P3_REG3_REG_10_ & ~P3_REG3_REG_11_;
  assign new_P3_SUB_609_U56 = ~P3_REG3_REG_12_ & ~P3_REG3_REG_13_;
  assign new_P3_SUB_609_U57 = ~P3_REG3_REG_14_ & ~P3_REG3_REG_15_;
  assign new_P3_SUB_609_U58 = ~P3_REG3_REG_16_ & ~P3_REG3_REG_17_;
  assign new_P3_SUB_609_U59 = ~P3_REG3_REG_18_ & ~P3_REG3_REG_19_;
  assign new_P3_SUB_609_U60 = ~P3_REG3_REG_20_ & ~P3_REG3_REG_21_;
  assign new_P3_SUB_609_U61 = ~P3_REG3_REG_22_ & ~P3_REG3_REG_23_;
  assign new_P3_SUB_609_U62 = ~P3_REG3_REG_24_ & ~P3_REG3_REG_25_;
  assign new_P3_SUB_609_U63 = ~P3_REG3_REG_26_ & ~P3_REG3_REG_27_;
  assign new_P3_SUB_609_U64 = P3_REG3_REG_3_ | P3_REG3_REG_4_;
  assign new_P3_SUB_609_U65 = P3_REG3_REG_3_ | P3_REG3_REG_4_ | P3_REG3_REG_5_ | P3_REG3_REG_6_;
  assign new_P3_SUB_609_U66 = ~new_P3_SUB_609_U31;
  assign new_P3_SUB_609_U67 = ~new_P3_SUB_609_U66 | ~new_P3_SUB_609_U32;
  assign new_P3_SUB_609_U68 = ~new_P3_SUB_609_U33;
  assign new_P3_SUB_609_U69 = ~P3_REG3_REG_9_ | ~new_P3_SUB_609_U67;
  assign new_P3_SUB_609_U70 = ~P3_REG3_REG_8_ | ~new_P3_SUB_609_U31;
  assign new_P3_SUB_609_U71 = ~P3_REG3_REG_7_ | ~new_P3_SUB_609_U65;
  assign new_P3_SUB_609_U72 = ~P3_REG3_REG_4_ | ~P3_REG3_REG_3_;
  assign new_P3_SUB_609_U73 = ~new_P3_SUB_609_U68 | ~new_P3_SUB_609_U52;
  assign new_P3_SUB_609_U74 = ~new_P3_SUB_609_U34;
  assign new_P3_SUB_609_U75 = ~new_P3_SUB_609_U74 | ~new_P3_SUB_609_U51;
  assign new_P3_SUB_609_U76 = ~new_P3_SUB_609_U35;
  assign new_P3_SUB_609_U77 = ~new_P3_SUB_609_U76 | ~new_P3_SUB_609_U50;
  assign new_P3_SUB_609_U78 = ~new_P3_SUB_609_U36;
  assign new_P3_SUB_609_U79 = ~new_P3_SUB_609_U78 | ~new_P3_SUB_609_U49;
  assign new_P3_SUB_609_U80 = ~new_P3_SUB_609_U37;
  assign new_P3_SUB_609_U81 = ~new_P3_SUB_609_U80 | ~new_P3_SUB_609_U48;
  assign new_P3_SUB_609_U82 = ~new_P3_SUB_609_U38;
  assign new_P3_SUB_609_U83 = ~new_P3_SUB_609_U82 | ~new_P3_SUB_609_U47;
  assign new_P3_SUB_609_U84 = ~new_P3_SUB_609_U39;
  assign new_P3_SUB_609_U85 = ~new_P3_SUB_609_U84 | ~new_P3_SUB_609_U46;
  assign new_P3_SUB_609_U86 = ~new_P3_SUB_609_U40;
  assign new_P3_SUB_609_U87 = ~new_P3_SUB_609_U86 | ~new_P3_SUB_609_U45;
  assign new_P3_SUB_609_U88 = ~new_P3_SUB_609_U41;
  assign new_P3_SUB_609_U89 = ~new_P3_SUB_609_U88 | ~new_P3_SUB_609_U44;
  assign new_P3_SUB_609_U90 = ~new_P3_SUB_609_U42;
  assign new_P3_SUB_609_U91 = ~new_P3_SUB_609_U90 | ~new_P3_SUB_609_U43;
  assign new_P3_SUB_609_U92 = ~new_P3_SUB_609_U91;
  assign new_P3_SUB_609_U93 = ~P3_REG3_REG_28_ | ~new_P3_SUB_609_U42;
  assign new_P3_SUB_609_U94 = ~P3_REG3_REG_27_ | ~new_P3_SUB_609_U89;
  assign new_P3_SUB_609_U95 = ~P3_REG3_REG_26_ | ~new_P3_SUB_609_U41;
  assign new_P3_SUB_609_U96 = ~P3_REG3_REG_25_ | ~new_P3_SUB_609_U87;
  assign new_P3_SUB_609_U97 = ~P3_REG3_REG_24_ | ~new_P3_SUB_609_U40;
  assign new_P3_SUB_609_U98 = ~P3_REG3_REG_23_ | ~new_P3_SUB_609_U85;
  assign new_P3_SUB_609_U99 = ~P3_REG3_REG_22_ | ~new_P3_SUB_609_U39;
  assign new_P3_SUB_609_U100 = ~P3_REG3_REG_21_ | ~new_P3_SUB_609_U83;
  assign new_P3_SUB_609_U101 = ~P3_REG3_REG_20_ | ~new_P3_SUB_609_U38;
  assign new_P3_SUB_609_U102 = ~P3_REG3_REG_19_ | ~new_P3_SUB_609_U81;
  assign new_P3_SUB_609_U103 = ~P3_REG3_REG_18_ | ~new_P3_SUB_609_U37;
  assign new_P3_SUB_609_U104 = ~P3_REG3_REG_17_ | ~new_P3_SUB_609_U79;
  assign new_P3_SUB_609_U105 = ~P3_REG3_REG_16_ | ~new_P3_SUB_609_U36;
  assign new_P3_SUB_609_U106 = ~P3_REG3_REG_15_ | ~new_P3_SUB_609_U77;
  assign new_P3_SUB_609_U107 = ~P3_REG3_REG_14_ | ~new_P3_SUB_609_U35;
  assign new_P3_SUB_609_U108 = ~P3_REG3_REG_13_ | ~new_P3_SUB_609_U75;
  assign new_P3_SUB_609_U109 = ~P3_REG3_REG_12_ | ~new_P3_SUB_609_U34;
  assign new_P3_SUB_609_U110 = ~P3_REG3_REG_11_ | ~new_P3_SUB_609_U73;
  assign new_P3_SUB_609_U111 = ~P3_REG3_REG_10_ | ~new_P3_SUB_609_U33;
  assign new_P3_SUB_609_U112 = P3_REG3_REG_5_ | P3_REG3_REG_4_ | P3_REG3_REG_3_;
  assign new_P3_SUB_609_U113 = ~P3_REG3_REG_6_ | ~new_P3_SUB_609_U112;
  assign new_P3_SUB_609_U114 = ~P3_REG3_REG_5_ | ~new_P3_SUB_609_U64;
  assign new_P3_SUB_609_U115 = P3_REG3_REG_5_ | P3_REG3_REG_4_ | P3_REG3_REG_3_;
  assign new_P3_R1095_U6 = new_P3_R1095_U210 & new_P3_R1095_U209;
  assign new_P3_R1095_U7 = new_P3_R1095_U189 & new_P3_R1095_U245;
  assign new_P3_R1095_U8 = new_P3_R1095_U247 & new_P3_R1095_U246;
  assign new_P3_R1095_U9 = new_P3_R1095_U190 & new_P3_R1095_U262;
  assign new_P3_R1095_U10 = new_P3_R1095_U264 & new_P3_R1095_U263;
  assign new_P3_R1095_U11 = new_P3_R1095_U191 & new_P3_R1095_U286;
  assign new_P3_R1095_U12 = new_P3_R1095_U288 & new_P3_R1095_U287;
  assign new_P3_R1095_U13 = new_P3_R1095_U213 & new_P3_R1095_U208 & new_P3_R1095_U194;
  assign new_P3_R1095_U14 = new_P3_R1095_U218 & new_P3_R1095_U195;
  assign new_P3_R1095_U15 = new_P3_R1095_U392 & new_P3_R1095_U391;
  assign new_P3_R1095_U16 = ~new_P3_R1095_U342 | ~new_P3_R1095_U345;
  assign new_P3_R1095_U17 = ~new_P3_R1095_U331 | ~new_P3_R1095_U334;
  assign new_P3_R1095_U18 = ~new_P3_R1095_U320 | ~new_P3_R1095_U323;
  assign new_P3_R1095_U19 = ~new_P3_R1095_U312 | ~new_P3_R1095_U314;
  assign new_P3_R1095_U20 = ~new_P3_R1095_U351 | ~new_P3_R1095_U162 | ~new_P3_R1095_U183;
  assign new_P3_R1095_U21 = ~new_P3_R1095_U241 | ~new_P3_R1095_U243;
  assign new_P3_R1095_U22 = ~new_P3_R1095_U233 | ~new_P3_R1095_U236;
  assign new_P3_R1095_U23 = ~new_P3_R1095_U225 | ~new_P3_R1095_U227;
  assign new_P3_R1095_U24 = ~new_P3_R1095_U172 | ~new_P3_R1095_U348;
  assign new_P3_R1095_U25 = ~new_P3_U3069;
  assign new_P3_R1095_U26 = ~new_P3_U3069 | ~new_P3_R1095_U39;
  assign new_P3_R1095_U27 = ~new_P3_U3083;
  assign new_P3_R1095_U28 = ~new_P3_U3413;
  assign new_P3_R1095_U29 = ~new_P3_U3395;
  assign new_P3_R1095_U30 = ~new_P3_U3387;
  assign new_P3_R1095_U31 = ~new_P3_U3077;
  assign new_P3_R1095_U32 = ~new_P3_U3398;
  assign new_P3_R1095_U33 = ~new_P3_U3067;
  assign new_P3_R1095_U34 = ~new_P3_U3067 | ~new_P3_R1095_U29;
  assign new_P3_R1095_U35 = ~new_P3_U3063;
  assign new_P3_R1095_U36 = ~new_P3_U3404;
  assign new_P3_R1095_U37 = ~new_P3_U3407;
  assign new_P3_R1095_U38 = ~new_P3_U3401;
  assign new_P3_R1095_U39 = ~new_P3_U3410;
  assign new_P3_R1095_U40 = ~new_P3_U3070;
  assign new_P3_R1095_U41 = ~new_P3_U3066;
  assign new_P3_R1095_U42 = ~new_P3_U3059;
  assign new_P3_R1095_U43 = ~new_P3_U3059 | ~new_P3_R1095_U38;
  assign new_P3_R1095_U44 = ~new_P3_R1095_U214 | ~new_P3_R1095_U212;
  assign new_P3_R1095_U45 = ~new_P3_U3416;
  assign new_P3_R1095_U46 = ~new_P3_U3082;
  assign new_P3_R1095_U47 = ~new_P3_R1095_U44 | ~new_P3_R1095_U215;
  assign new_P3_R1095_U48 = ~new_P3_R1095_U43 | ~new_P3_R1095_U229;
  assign new_P3_R1095_U49 = ~new_P3_R1095_U349 | ~new_P3_R1095_U201 | ~new_P3_R1095_U185;
  assign new_P3_R1095_U50 = ~new_P3_U3901;
  assign new_P3_R1095_U51 = ~new_P3_U3422;
  assign new_P3_R1095_U52 = ~new_P3_U3419;
  assign new_P3_R1095_U53 = ~new_P3_U3062;
  assign new_P3_R1095_U54 = ~new_P3_U3061;
  assign new_P3_R1095_U55 = ~new_P3_U3082 | ~new_P3_R1095_U45;
  assign new_P3_R1095_U56 = ~new_P3_U3425;
  assign new_P3_R1095_U57 = ~new_P3_U3071;
  assign new_P3_R1095_U58 = ~new_P3_U3428;
  assign new_P3_R1095_U59 = ~new_P3_U3079;
  assign new_P3_R1095_U60 = ~new_P3_U3437;
  assign new_P3_R1095_U61 = ~new_P3_U3434;
  assign new_P3_R1095_U62 = ~new_P3_U3431;
  assign new_P3_R1095_U63 = ~new_P3_U3072;
  assign new_P3_R1095_U64 = ~new_P3_U3073;
  assign new_P3_R1095_U65 = ~new_P3_U3078;
  assign new_P3_R1095_U66 = ~new_P3_U3078 | ~new_P3_R1095_U62;
  assign new_P3_R1095_U67 = ~new_P3_U3440;
  assign new_P3_R1095_U68 = ~new_P3_U3068;
  assign new_P3_R1095_U69 = ~new_P3_U3081;
  assign new_P3_R1095_U70 = ~new_P3_U3445;
  assign new_P3_R1095_U71 = ~new_P3_U3080;
  assign new_P3_R1095_U72 = ~new_P3_U3907;
  assign new_P3_R1095_U73 = ~new_P3_U3075;
  assign new_P3_R1095_U74 = ~new_P3_U3904;
  assign new_P3_R1095_U75 = ~new_P3_U3905;
  assign new_P3_R1095_U76 = ~new_P3_U3906;
  assign new_P3_R1095_U77 = ~new_P3_U3065;
  assign new_P3_R1095_U78 = ~new_P3_U3060;
  assign new_P3_R1095_U79 = ~new_P3_U3074;
  assign new_P3_R1095_U80 = ~new_P3_U3074 | ~new_P3_R1095_U76;
  assign new_P3_R1095_U81 = ~new_P3_U3903;
  assign new_P3_R1095_U82 = ~new_P3_U3064;
  assign new_P3_R1095_U83 = ~new_P3_U3902;
  assign new_P3_R1095_U84 = ~new_P3_U3057;
  assign new_P3_R1095_U85 = ~new_P3_U3900;
  assign new_P3_R1095_U86 = ~new_P3_U3056;
  assign new_P3_R1095_U87 = ~new_P3_U3056 | ~new_P3_R1095_U50;
  assign new_P3_R1095_U88 = ~new_P3_U3052;
  assign new_P3_R1095_U89 = ~new_P3_U3899;
  assign new_P3_R1095_U90 = ~new_P3_U3053;
  assign new_P3_R1095_U91 = ~new_P3_R1095_U302 | ~new_P3_R1095_U301;
  assign new_P3_R1095_U92 = ~new_P3_R1095_U80 | ~new_P3_R1095_U316;
  assign new_P3_R1095_U93 = ~new_P3_R1095_U66 | ~new_P3_R1095_U327;
  assign new_P3_R1095_U94 = ~new_P3_R1095_U55 | ~new_P3_R1095_U338;
  assign new_P3_R1095_U95 = ~new_P3_U3076;
  assign new_P3_R1095_U96 = ~new_P3_R1095_U402 | ~new_P3_R1095_U401;
  assign new_P3_R1095_U97 = ~new_P3_R1095_U416 | ~new_P3_R1095_U415;
  assign new_P3_R1095_U98 = ~new_P3_R1095_U421 | ~new_P3_R1095_U420;
  assign new_P3_R1095_U99 = ~new_P3_R1095_U437 | ~new_P3_R1095_U436;
  assign new_P3_R1095_U100 = ~new_P3_R1095_U442 | ~new_P3_R1095_U441;
  assign new_P3_R1095_U101 = ~new_P3_R1095_U447 | ~new_P3_R1095_U446;
  assign new_P3_R1095_U102 = ~new_P3_R1095_U452 | ~new_P3_R1095_U451;
  assign new_P3_R1095_U103 = ~new_P3_R1095_U457 | ~new_P3_R1095_U456;
  assign new_P3_R1095_U104 = ~new_P3_R1095_U473 | ~new_P3_R1095_U472;
  assign new_P3_R1095_U105 = ~new_P3_R1095_U478 | ~new_P3_R1095_U477;
  assign new_P3_R1095_U106 = ~new_P3_R1095_U361 | ~new_P3_R1095_U360;
  assign new_P3_R1095_U107 = ~new_P3_R1095_U370 | ~new_P3_R1095_U369;
  assign new_P3_R1095_U108 = ~new_P3_R1095_U377 | ~new_P3_R1095_U376;
  assign new_P3_R1095_U109 = ~new_P3_R1095_U381 | ~new_P3_R1095_U380;
  assign new_P3_R1095_U110 = ~new_P3_R1095_U390 | ~new_P3_R1095_U389;
  assign new_P3_R1095_U111 = ~new_P3_R1095_U411 | ~new_P3_R1095_U410;
  assign new_P3_R1095_U112 = ~new_P3_R1095_U428 | ~new_P3_R1095_U427;
  assign new_P3_R1095_U113 = ~new_P3_R1095_U432 | ~new_P3_R1095_U431;
  assign new_P3_R1095_U114 = ~new_P3_R1095_U464 | ~new_P3_R1095_U463;
  assign new_P3_R1095_U115 = ~new_P3_R1095_U468 | ~new_P3_R1095_U467;
  assign new_P3_R1095_U116 = ~new_P3_R1095_U485 | ~new_P3_R1095_U484;
  assign new_P3_R1095_U117 = new_P3_R1095_U352 & new_P3_R1095_U193;
  assign new_P3_R1095_U118 = new_P3_R1095_U205 & new_P3_R1095_U206;
  assign new_P3_R1095_U119 = new_P3_R1095_U14 & new_P3_R1095_U13;
  assign new_P3_R1095_U120 = new_P3_R1095_U357 & new_P3_R1095_U354;
  assign new_P3_R1095_U121 = new_P3_R1095_U26 & new_P3_R1095_U363 & new_P3_R1095_U362;
  assign new_P3_R1095_U122 = new_P3_R1095_U366 & new_P3_R1095_U195;
  assign new_P3_R1095_U123 = new_P3_R1095_U235 & new_P3_R1095_U6;
  assign new_P3_R1095_U124 = new_P3_R1095_U373 & new_P3_R1095_U194;
  assign new_P3_R1095_U125 = new_P3_R1095_U34 & new_P3_R1095_U383 & new_P3_R1095_U382;
  assign new_P3_R1095_U126 = new_P3_R1095_U386 & new_P3_R1095_U193;
  assign new_P3_R1095_U127 = new_P3_R1095_U222 & new_P3_R1095_U7;
  assign new_P3_R1095_U128 = new_P3_R1095_U267 & new_P3_R1095_U9;
  assign new_P3_R1095_U129 = new_P3_R1095_U291 & new_P3_R1095_U11;
  assign new_P3_R1095_U130 = new_P3_R1095_U355 & new_P3_R1095_U192;
  assign new_P3_R1095_U131 = new_P3_R1095_U306 & new_P3_R1095_U307;
  assign new_P3_R1095_U132 = new_P3_R1095_U309 & new_P3_R1095_U395;
  assign new_P3_R1095_U133 = new_P3_R1095_U306 & new_P3_R1095_U307;
  assign new_P3_R1095_U134 = new_P3_R1095_U15 & new_P3_R1095_U310;
  assign new_P3_R1095_U135 = ~new_P3_R1095_U399 | ~new_P3_R1095_U398;
  assign new_P3_R1095_U136 = new_P3_R1095_U87 & new_P3_R1095_U404 & new_P3_R1095_U403;
  assign new_P3_R1095_U137 = new_P3_R1095_U407 & new_P3_R1095_U192;
  assign new_P3_R1095_U138 = ~new_P3_R1095_U413 | ~new_P3_R1095_U412;
  assign new_P3_R1095_U139 = ~new_P3_R1095_U418 | ~new_P3_R1095_U417;
  assign new_P3_R1095_U140 = new_P3_R1095_U322 & new_P3_R1095_U12;
  assign new_P3_R1095_U141 = new_P3_R1095_U424 & new_P3_R1095_U191;
  assign new_P3_R1095_U142 = ~new_P3_R1095_U434 | ~new_P3_R1095_U433;
  assign new_P3_R1095_U143 = ~new_P3_R1095_U439 | ~new_P3_R1095_U438;
  assign new_P3_R1095_U144 = ~new_P3_R1095_U444 | ~new_P3_R1095_U443;
  assign new_P3_R1095_U145 = ~new_P3_R1095_U449 | ~new_P3_R1095_U448;
  assign new_P3_R1095_U146 = ~new_P3_R1095_U454 | ~new_P3_R1095_U453;
  assign new_P3_R1095_U147 = new_P3_R1095_U333 & new_P3_R1095_U10;
  assign new_P3_R1095_U148 = new_P3_R1095_U460 & new_P3_R1095_U190;
  assign new_P3_R1095_U149 = ~new_P3_R1095_U470 | ~new_P3_R1095_U469;
  assign new_P3_R1095_U150 = ~new_P3_R1095_U475 | ~new_P3_R1095_U474;
  assign new_P3_R1095_U151 = new_P3_R1095_U344 & new_P3_R1095_U8;
  assign new_P3_R1095_U152 = new_P3_R1095_U481 & new_P3_R1095_U189;
  assign new_P3_R1095_U153 = new_P3_R1095_U359 & new_P3_R1095_U358;
  assign new_P3_R1095_U154 = ~new_P3_R1095_U120 | ~new_P3_R1095_U356;
  assign new_P3_R1095_U155 = new_P3_R1095_U368 & new_P3_R1095_U367;
  assign new_P3_R1095_U156 = new_P3_R1095_U375 & new_P3_R1095_U374;
  assign new_P3_R1095_U157 = new_P3_R1095_U379 & new_P3_R1095_U378;
  assign new_P3_R1095_U158 = ~new_P3_R1095_U118 | ~new_P3_R1095_U203;
  assign new_P3_R1095_U159 = new_P3_R1095_U388 & new_P3_R1095_U387;
  assign new_P3_R1095_U160 = ~new_P3_U3908;
  assign new_P3_R1095_U161 = ~new_P3_U3054;
  assign new_P3_R1095_U162 = new_P3_R1095_U397 & new_P3_R1095_U396;
  assign new_P3_R1095_U163 = ~new_P3_R1095_U131 | ~new_P3_R1095_U304;
  assign new_P3_R1095_U164 = new_P3_R1095_U409 & new_P3_R1095_U408;
  assign new_P3_R1095_U165 = ~new_P3_R1095_U298 | ~new_P3_R1095_U297;
  assign new_P3_R1095_U166 = ~new_P3_R1095_U294 | ~new_P3_R1095_U293;
  assign new_P3_R1095_U167 = new_P3_R1095_U426 & new_P3_R1095_U425;
  assign new_P3_R1095_U168 = new_P3_R1095_U430 & new_P3_R1095_U429;
  assign new_P3_R1095_U169 = ~new_P3_R1095_U284 | ~new_P3_R1095_U283;
  assign new_P3_R1095_U170 = ~new_P3_R1095_U280 | ~new_P3_R1095_U279;
  assign new_P3_R1095_U171 = ~new_P3_U3392;
  assign new_P3_R1095_U172 = ~new_P3_U3387 | ~new_P3_R1095_U95;
  assign new_P3_R1095_U173 = ~new_P3_R1095_U350 | ~new_P3_R1095_U276 | ~new_P3_R1095_U184;
  assign new_P3_R1095_U174 = ~new_P3_U3443;
  assign new_P3_R1095_U175 = ~new_P3_R1095_U274 | ~new_P3_R1095_U273;
  assign new_P3_R1095_U176 = ~new_P3_R1095_U270 | ~new_P3_R1095_U269;
  assign new_P3_R1095_U177 = new_P3_R1095_U462 & new_P3_R1095_U461;
  assign new_P3_R1095_U178 = new_P3_R1095_U466 & new_P3_R1095_U465;
  assign new_P3_R1095_U179 = ~new_P3_R1095_U260 | ~new_P3_R1095_U259;
  assign new_P3_R1095_U180 = ~new_P3_R1095_U256 | ~new_P3_R1095_U255;
  assign new_P3_R1095_U181 = ~new_P3_R1095_U252 | ~new_P3_R1095_U251;
  assign new_P3_R1095_U182 = new_P3_R1095_U483 & new_P3_R1095_U482;
  assign new_P3_R1095_U183 = ~new_P3_R1095_U132 | ~new_P3_R1095_U163;
  assign new_P3_R1095_U184 = ~new_P3_R1095_U175 | ~new_P3_R1095_U174;
  assign new_P3_R1095_U185 = ~new_P3_R1095_U172 | ~new_P3_R1095_U171;
  assign new_P3_R1095_U186 = ~new_P3_R1095_U87;
  assign new_P3_R1095_U187 = ~new_P3_R1095_U34;
  assign new_P3_R1095_U188 = ~new_P3_R1095_U26;
  assign new_P3_R1095_U189 = ~new_P3_U3419 | ~new_P3_R1095_U54;
  assign new_P3_R1095_U190 = ~new_P3_U3434 | ~new_P3_R1095_U64;
  assign new_P3_R1095_U191 = ~new_P3_U3905 | ~new_P3_R1095_U78;
  assign new_P3_R1095_U192 = ~new_P3_U3901 | ~new_P3_R1095_U86;
  assign new_P3_R1095_U193 = ~new_P3_U3395 | ~new_P3_R1095_U33;
  assign new_P3_R1095_U194 = ~new_P3_U3404 | ~new_P3_R1095_U41;
  assign new_P3_R1095_U195 = ~new_P3_U3410 | ~new_P3_R1095_U25;
  assign new_P3_R1095_U196 = ~new_P3_R1095_U66;
  assign new_P3_R1095_U197 = ~new_P3_R1095_U80;
  assign new_P3_R1095_U198 = ~new_P3_R1095_U43;
  assign new_P3_R1095_U199 = ~new_P3_R1095_U55;
  assign new_P3_R1095_U200 = ~new_P3_R1095_U172;
  assign new_P3_R1095_U201 = ~new_P3_U3077 | ~new_P3_R1095_U172;
  assign new_P3_R1095_U202 = ~new_P3_R1095_U49;
  assign new_P3_R1095_U203 = ~new_P3_R1095_U117 | ~new_P3_R1095_U49;
  assign new_P3_R1095_U204 = ~new_P3_R1095_U35 | ~new_P3_R1095_U34;
  assign new_P3_R1095_U205 = ~new_P3_R1095_U204 | ~new_P3_R1095_U32;
  assign new_P3_R1095_U206 = ~new_P3_U3063 | ~new_P3_R1095_U187;
  assign new_P3_R1095_U207 = ~new_P3_R1095_U158;
  assign new_P3_R1095_U208 = ~new_P3_U3407 | ~new_P3_R1095_U40;
  assign new_P3_R1095_U209 = ~new_P3_U3070 | ~new_P3_R1095_U37;
  assign new_P3_R1095_U210 = ~new_P3_U3066 | ~new_P3_R1095_U36;
  assign new_P3_R1095_U211 = ~new_P3_R1095_U198 | ~new_P3_R1095_U194;
  assign new_P3_R1095_U212 = ~new_P3_R1095_U6 | ~new_P3_R1095_U211;
  assign new_P3_R1095_U213 = ~new_P3_U3401 | ~new_P3_R1095_U42;
  assign new_P3_R1095_U214 = ~new_P3_U3407 | ~new_P3_R1095_U40;
  assign new_P3_R1095_U215 = ~new_P3_R1095_U13 | ~new_P3_R1095_U158;
  assign new_P3_R1095_U216 = ~new_P3_R1095_U44;
  assign new_P3_R1095_U217 = ~new_P3_R1095_U47;
  assign new_P3_R1095_U218 = ~new_P3_U3413 | ~new_P3_R1095_U27;
  assign new_P3_R1095_U219 = ~new_P3_R1095_U27 | ~new_P3_R1095_U26;
  assign new_P3_R1095_U220 = ~new_P3_U3083 | ~new_P3_R1095_U188;
  assign new_P3_R1095_U221 = ~new_P3_R1095_U154;
  assign new_P3_R1095_U222 = ~new_P3_U3416 | ~new_P3_R1095_U46;
  assign new_P3_R1095_U223 = ~new_P3_R1095_U222 | ~new_P3_R1095_U55;
  assign new_P3_R1095_U224 = ~new_P3_R1095_U217 | ~new_P3_R1095_U26;
  assign new_P3_R1095_U225 = ~new_P3_R1095_U122 | ~new_P3_R1095_U224;
  assign new_P3_R1095_U226 = ~new_P3_R1095_U47 | ~new_P3_R1095_U195;
  assign new_P3_R1095_U227 = ~new_P3_R1095_U121 | ~new_P3_R1095_U226;
  assign new_P3_R1095_U228 = ~new_P3_R1095_U26 | ~new_P3_R1095_U195;
  assign new_P3_R1095_U229 = ~new_P3_R1095_U213 | ~new_P3_R1095_U158;
  assign new_P3_R1095_U230 = ~new_P3_R1095_U48;
  assign new_P3_R1095_U231 = ~new_P3_U3066 | ~new_P3_R1095_U36;
  assign new_P3_R1095_U232 = ~new_P3_R1095_U230 | ~new_P3_R1095_U231;
  assign new_P3_R1095_U233 = ~new_P3_R1095_U124 | ~new_P3_R1095_U232;
  assign new_P3_R1095_U234 = ~new_P3_R1095_U48 | ~new_P3_R1095_U194;
  assign new_P3_R1095_U235 = ~new_P3_U3407 | ~new_P3_R1095_U40;
  assign new_P3_R1095_U236 = ~new_P3_R1095_U123 | ~new_P3_R1095_U234;
  assign new_P3_R1095_U237 = ~new_P3_U3066 | ~new_P3_R1095_U36;
  assign new_P3_R1095_U238 = ~new_P3_R1095_U194 | ~new_P3_R1095_U237;
  assign new_P3_R1095_U239 = ~new_P3_R1095_U213 | ~new_P3_R1095_U43;
  assign new_P3_R1095_U240 = ~new_P3_R1095_U202 | ~new_P3_R1095_U34;
  assign new_P3_R1095_U241 = ~new_P3_R1095_U126 | ~new_P3_R1095_U240;
  assign new_P3_R1095_U242 = ~new_P3_R1095_U49 | ~new_P3_R1095_U193;
  assign new_P3_R1095_U243 = ~new_P3_R1095_U125 | ~new_P3_R1095_U242;
  assign new_P3_R1095_U244 = ~new_P3_R1095_U193 | ~new_P3_R1095_U34;
  assign new_P3_R1095_U245 = ~new_P3_U3422 | ~new_P3_R1095_U53;
  assign new_P3_R1095_U246 = ~new_P3_U3062 | ~new_P3_R1095_U51;
  assign new_P3_R1095_U247 = ~new_P3_U3061 | ~new_P3_R1095_U52;
  assign new_P3_R1095_U248 = ~new_P3_R1095_U199 | ~new_P3_R1095_U7;
  assign new_P3_R1095_U249 = ~new_P3_R1095_U8 | ~new_P3_R1095_U248;
  assign new_P3_R1095_U250 = ~new_P3_U3422 | ~new_P3_R1095_U53;
  assign new_P3_R1095_U251 = ~new_P3_R1095_U127 | ~new_P3_R1095_U154;
  assign new_P3_R1095_U252 = ~new_P3_R1095_U250 | ~new_P3_R1095_U249;
  assign new_P3_R1095_U253 = ~new_P3_R1095_U181;
  assign new_P3_R1095_U254 = ~new_P3_U3425 | ~new_P3_R1095_U57;
  assign new_P3_R1095_U255 = ~new_P3_R1095_U254 | ~new_P3_R1095_U181;
  assign new_P3_R1095_U256 = ~new_P3_U3071 | ~new_P3_R1095_U56;
  assign new_P3_R1095_U257 = ~new_P3_R1095_U180;
  assign new_P3_R1095_U258 = ~new_P3_U3428 | ~new_P3_R1095_U59;
  assign new_P3_R1095_U259 = ~new_P3_R1095_U258 | ~new_P3_R1095_U180;
  assign new_P3_R1095_U260 = ~new_P3_U3079 | ~new_P3_R1095_U58;
  assign new_P3_R1095_U261 = ~new_P3_R1095_U179;
  assign new_P3_R1095_U262 = ~new_P3_U3437 | ~new_P3_R1095_U63;
  assign new_P3_R1095_U263 = ~new_P3_U3072 | ~new_P3_R1095_U60;
  assign new_P3_R1095_U264 = ~new_P3_U3073 | ~new_P3_R1095_U61;
  assign new_P3_R1095_U265 = ~new_P3_R1095_U196 | ~new_P3_R1095_U9;
  assign new_P3_R1095_U266 = ~new_P3_R1095_U10 | ~new_P3_R1095_U265;
  assign new_P3_R1095_U267 = ~new_P3_U3431 | ~new_P3_R1095_U65;
  assign new_P3_R1095_U268 = ~new_P3_U3437 | ~new_P3_R1095_U63;
  assign new_P3_R1095_U269 = ~new_P3_R1095_U128 | ~new_P3_R1095_U179;
  assign new_P3_R1095_U270 = ~new_P3_R1095_U268 | ~new_P3_R1095_U266;
  assign new_P3_R1095_U271 = ~new_P3_R1095_U176;
  assign new_P3_R1095_U272 = ~new_P3_U3440 | ~new_P3_R1095_U68;
  assign new_P3_R1095_U273 = ~new_P3_R1095_U272 | ~new_P3_R1095_U176;
  assign new_P3_R1095_U274 = ~new_P3_U3068 | ~new_P3_R1095_U67;
  assign new_P3_R1095_U275 = ~new_P3_R1095_U175;
  assign new_P3_R1095_U276 = ~new_P3_U3081 | ~new_P3_R1095_U175;
  assign new_P3_R1095_U277 = ~new_P3_R1095_U173;
  assign new_P3_R1095_U278 = ~new_P3_U3445 | ~new_P3_R1095_U71;
  assign new_P3_R1095_U279 = ~new_P3_R1095_U278 | ~new_P3_R1095_U173;
  assign new_P3_R1095_U280 = ~new_P3_U3080 | ~new_P3_R1095_U70;
  assign new_P3_R1095_U281 = ~new_P3_R1095_U170;
  assign new_P3_R1095_U282 = ~new_P3_U3907 | ~new_P3_R1095_U73;
  assign new_P3_R1095_U283 = ~new_P3_R1095_U282 | ~new_P3_R1095_U170;
  assign new_P3_R1095_U284 = ~new_P3_U3075 | ~new_P3_R1095_U72;
  assign new_P3_R1095_U285 = ~new_P3_R1095_U169;
  assign new_P3_R1095_U286 = ~new_P3_U3904 | ~new_P3_R1095_U77;
  assign new_P3_R1095_U287 = ~new_P3_U3065 | ~new_P3_R1095_U74;
  assign new_P3_R1095_U288 = ~new_P3_U3060 | ~new_P3_R1095_U75;
  assign new_P3_R1095_U289 = ~new_P3_R1095_U197 | ~new_P3_R1095_U11;
  assign new_P3_R1095_U290 = ~new_P3_R1095_U12 | ~new_P3_R1095_U289;
  assign new_P3_R1095_U291 = ~new_P3_U3906 | ~new_P3_R1095_U79;
  assign new_P3_R1095_U292 = ~new_P3_U3904 | ~new_P3_R1095_U77;
  assign new_P3_R1095_U293 = ~new_P3_R1095_U129 | ~new_P3_R1095_U169;
  assign new_P3_R1095_U294 = ~new_P3_R1095_U292 | ~new_P3_R1095_U290;
  assign new_P3_R1095_U295 = ~new_P3_R1095_U166;
  assign new_P3_R1095_U296 = ~new_P3_U3903 | ~new_P3_R1095_U82;
  assign new_P3_R1095_U297 = ~new_P3_R1095_U296 | ~new_P3_R1095_U166;
  assign new_P3_R1095_U298 = ~new_P3_U3064 | ~new_P3_R1095_U81;
  assign new_P3_R1095_U299 = ~new_P3_R1095_U165;
  assign new_P3_R1095_U300 = ~new_P3_U3902 | ~new_P3_R1095_U84;
  assign new_P3_R1095_U301 = ~new_P3_R1095_U300 | ~new_P3_R1095_U165;
  assign new_P3_R1095_U302 = ~new_P3_U3057 | ~new_P3_R1095_U83;
  assign new_P3_R1095_U303 = ~new_P3_R1095_U91;
  assign new_P3_R1095_U304 = ~new_P3_R1095_U130 | ~new_P3_R1095_U91;
  assign new_P3_R1095_U305 = ~new_P3_R1095_U88 | ~new_P3_R1095_U87;
  assign new_P3_R1095_U306 = ~new_P3_R1095_U305 | ~new_P3_R1095_U85;
  assign new_P3_R1095_U307 = ~new_P3_U3052 | ~new_P3_R1095_U186;
  assign new_P3_R1095_U308 = ~new_P3_R1095_U163;
  assign new_P3_R1095_U309 = ~new_P3_U3899 | ~new_P3_R1095_U90;
  assign new_P3_R1095_U310 = ~new_P3_U3053 | ~new_P3_R1095_U89;
  assign new_P3_R1095_U311 = ~new_P3_R1095_U303 | ~new_P3_R1095_U87;
  assign new_P3_R1095_U312 = ~new_P3_R1095_U137 | ~new_P3_R1095_U311;
  assign new_P3_R1095_U313 = ~new_P3_R1095_U91 | ~new_P3_R1095_U192;
  assign new_P3_R1095_U314 = ~new_P3_R1095_U136 | ~new_P3_R1095_U313;
  assign new_P3_R1095_U315 = ~new_P3_R1095_U192 | ~new_P3_R1095_U87;
  assign new_P3_R1095_U316 = ~new_P3_R1095_U291 | ~new_P3_R1095_U169;
  assign new_P3_R1095_U317 = ~new_P3_R1095_U92;
  assign new_P3_R1095_U318 = ~new_P3_U3060 | ~new_P3_R1095_U75;
  assign new_P3_R1095_U319 = ~new_P3_R1095_U317 | ~new_P3_R1095_U318;
  assign new_P3_R1095_U320 = ~new_P3_R1095_U141 | ~new_P3_R1095_U319;
  assign new_P3_R1095_U321 = ~new_P3_R1095_U92 | ~new_P3_R1095_U191;
  assign new_P3_R1095_U322 = ~new_P3_U3904 | ~new_P3_R1095_U77;
  assign new_P3_R1095_U323 = ~new_P3_R1095_U140 | ~new_P3_R1095_U321;
  assign new_P3_R1095_U324 = ~new_P3_U3060 | ~new_P3_R1095_U75;
  assign new_P3_R1095_U325 = ~new_P3_R1095_U191 | ~new_P3_R1095_U324;
  assign new_P3_R1095_U326 = ~new_P3_R1095_U291 | ~new_P3_R1095_U80;
  assign new_P3_R1095_U327 = ~new_P3_R1095_U267 | ~new_P3_R1095_U179;
  assign new_P3_R1095_U328 = ~new_P3_R1095_U93;
  assign new_P3_R1095_U329 = ~new_P3_U3073 | ~new_P3_R1095_U61;
  assign new_P3_R1095_U330 = ~new_P3_R1095_U328 | ~new_P3_R1095_U329;
  assign new_P3_R1095_U331 = ~new_P3_R1095_U148 | ~new_P3_R1095_U330;
  assign new_P3_R1095_U332 = ~new_P3_R1095_U93 | ~new_P3_R1095_U190;
  assign new_P3_R1095_U333 = ~new_P3_U3437 | ~new_P3_R1095_U63;
  assign new_P3_R1095_U334 = ~new_P3_R1095_U147 | ~new_P3_R1095_U332;
  assign new_P3_R1095_U335 = ~new_P3_U3073 | ~new_P3_R1095_U61;
  assign new_P3_R1095_U336 = ~new_P3_R1095_U190 | ~new_P3_R1095_U335;
  assign new_P3_R1095_U337 = ~new_P3_R1095_U267 | ~new_P3_R1095_U66;
  assign new_P3_R1095_U338 = ~new_P3_R1095_U222 | ~new_P3_R1095_U154;
  assign new_P3_R1095_U339 = ~new_P3_R1095_U94;
  assign new_P3_R1095_U340 = ~new_P3_U3061 | ~new_P3_R1095_U52;
  assign new_P3_R1095_U341 = ~new_P3_R1095_U339 | ~new_P3_R1095_U340;
  assign new_P3_R1095_U342 = ~new_P3_R1095_U152 | ~new_P3_R1095_U341;
  assign new_P3_R1095_U343 = ~new_P3_R1095_U94 | ~new_P3_R1095_U189;
  assign new_P3_R1095_U344 = ~new_P3_U3422 | ~new_P3_R1095_U53;
  assign new_P3_R1095_U345 = ~new_P3_R1095_U151 | ~new_P3_R1095_U343;
  assign new_P3_R1095_U346 = ~new_P3_U3061 | ~new_P3_R1095_U52;
  assign new_P3_R1095_U347 = ~new_P3_R1095_U189 | ~new_P3_R1095_U346;
  assign new_P3_R1095_U348 = ~new_P3_U3076 | ~new_P3_R1095_U30;
  assign new_P3_R1095_U349 = ~new_P3_U3077 | ~new_P3_R1095_U171;
  assign new_P3_R1095_U350 = ~new_P3_U3081 | ~new_P3_R1095_U174;
  assign new_P3_R1095_U351 = ~new_P3_R1095_U134 | ~new_P3_R1095_U133 | ~new_P3_R1095_U304;
  assign new_P3_R1095_U352 = ~new_P3_U3398 | ~new_P3_R1095_U35;
  assign new_P3_R1095_U353 = ~new_P3_U3413 | ~new_P3_R1095_U220;
  assign new_P3_R1095_U354 = ~new_P3_R1095_U353 | ~new_P3_R1095_U219;
  assign new_P3_R1095_U355 = ~new_P3_U3900 | ~new_P3_R1095_U88;
  assign new_P3_R1095_U356 = ~new_P3_R1095_U119 | ~new_P3_R1095_U158;
  assign new_P3_R1095_U357 = ~new_P3_R1095_U216 | ~new_P3_R1095_U14;
  assign new_P3_R1095_U358 = ~new_P3_U3416 | ~new_P3_R1095_U46;
  assign new_P3_R1095_U359 = ~new_P3_U3082 | ~new_P3_R1095_U45;
  assign new_P3_R1095_U360 = ~new_P3_R1095_U223 | ~new_P3_R1095_U154;
  assign new_P3_R1095_U361 = ~new_P3_R1095_U221 | ~new_P3_R1095_U153;
  assign new_P3_R1095_U362 = ~new_P3_U3413 | ~new_P3_R1095_U27;
  assign new_P3_R1095_U363 = ~new_P3_U3083 | ~new_P3_R1095_U28;
  assign new_P3_R1095_U364 = ~new_P3_U3413 | ~new_P3_R1095_U27;
  assign new_P3_R1095_U365 = ~new_P3_U3083 | ~new_P3_R1095_U28;
  assign new_P3_R1095_U366 = ~new_P3_R1095_U365 | ~new_P3_R1095_U364;
  assign new_P3_R1095_U367 = ~new_P3_U3410 | ~new_P3_R1095_U25;
  assign new_P3_R1095_U368 = ~new_P3_U3069 | ~new_P3_R1095_U39;
  assign new_P3_R1095_U369 = ~new_P3_R1095_U228 | ~new_P3_R1095_U47;
  assign new_P3_R1095_U370 = ~new_P3_R1095_U155 | ~new_P3_R1095_U217;
  assign new_P3_R1095_U371 = ~new_P3_U3407 | ~new_P3_R1095_U40;
  assign new_P3_R1095_U372 = ~new_P3_U3070 | ~new_P3_R1095_U37;
  assign new_P3_R1095_U373 = ~new_P3_R1095_U372 | ~new_P3_R1095_U371;
  assign new_P3_R1095_U374 = ~new_P3_U3404 | ~new_P3_R1095_U41;
  assign new_P3_R1095_U375 = ~new_P3_U3066 | ~new_P3_R1095_U36;
  assign new_P3_R1095_U376 = ~new_P3_R1095_U238 | ~new_P3_R1095_U48;
  assign new_P3_R1095_U377 = ~new_P3_R1095_U156 | ~new_P3_R1095_U230;
  assign new_P3_R1095_U378 = ~new_P3_U3401 | ~new_P3_R1095_U42;
  assign new_P3_R1095_U379 = ~new_P3_U3059 | ~new_P3_R1095_U38;
  assign new_P3_R1095_U380 = ~new_P3_R1095_U239 | ~new_P3_R1095_U158;
  assign new_P3_R1095_U381 = ~new_P3_R1095_U207 | ~new_P3_R1095_U157;
  assign new_P3_R1095_U382 = ~new_P3_U3398 | ~new_P3_R1095_U35;
  assign new_P3_R1095_U383 = ~new_P3_U3063 | ~new_P3_R1095_U32;
  assign new_P3_R1095_U384 = ~new_P3_U3398 | ~new_P3_R1095_U35;
  assign new_P3_R1095_U385 = ~new_P3_U3063 | ~new_P3_R1095_U32;
  assign new_P3_R1095_U386 = ~new_P3_R1095_U385 | ~new_P3_R1095_U384;
  assign new_P3_R1095_U387 = ~new_P3_U3395 | ~new_P3_R1095_U33;
  assign new_P3_R1095_U388 = ~new_P3_U3067 | ~new_P3_R1095_U29;
  assign new_P3_R1095_U389 = ~new_P3_R1095_U244 | ~new_P3_R1095_U49;
  assign new_P3_R1095_U390 = ~new_P3_R1095_U159 | ~new_P3_R1095_U202;
  assign new_P3_R1095_U391 = ~new_P3_U3908 | ~new_P3_R1095_U161;
  assign new_P3_R1095_U392 = ~new_P3_U3054 | ~new_P3_R1095_U160;
  assign new_P3_R1095_U393 = ~new_P3_U3908 | ~new_P3_R1095_U161;
  assign new_P3_R1095_U394 = ~new_P3_U3054 | ~new_P3_R1095_U160;
  assign new_P3_R1095_U395 = ~new_P3_R1095_U394 | ~new_P3_R1095_U393;
  assign new_P3_R1095_U396 = ~new_P3_R1095_U89 | ~new_P3_U3053 | ~new_P3_R1095_U395;
  assign new_P3_R1095_U397 = ~new_P3_U3899 | ~new_P3_R1095_U15 | ~new_P3_R1095_U90;
  assign new_P3_R1095_U398 = ~new_P3_U3899 | ~new_P3_R1095_U90;
  assign new_P3_R1095_U399 = ~new_P3_U3053 | ~new_P3_R1095_U89;
  assign new_P3_R1095_U400 = ~new_P3_R1095_U135;
  assign new_P3_R1095_U401 = ~new_P3_R1095_U308 | ~new_P3_R1095_U400;
  assign new_P3_R1095_U402 = ~new_P3_R1095_U135 | ~new_P3_R1095_U163;
  assign new_P3_R1095_U403 = ~new_P3_U3900 | ~new_P3_R1095_U88;
  assign new_P3_R1095_U404 = ~new_P3_U3052 | ~new_P3_R1095_U85;
  assign new_P3_R1095_U405 = ~new_P3_U3900 | ~new_P3_R1095_U88;
  assign new_P3_R1095_U406 = ~new_P3_U3052 | ~new_P3_R1095_U85;
  assign new_P3_R1095_U407 = ~new_P3_R1095_U406 | ~new_P3_R1095_U405;
  assign new_P3_R1095_U408 = ~new_P3_U3901 | ~new_P3_R1095_U86;
  assign new_P3_R1095_U409 = ~new_P3_U3056 | ~new_P3_R1095_U50;
  assign new_P3_R1095_U410 = ~new_P3_R1095_U315 | ~new_P3_R1095_U91;
  assign new_P3_R1095_U411 = ~new_P3_R1095_U164 | ~new_P3_R1095_U303;
  assign new_P3_R1095_U412 = ~new_P3_U3902 | ~new_P3_R1095_U84;
  assign new_P3_R1095_U413 = ~new_P3_U3057 | ~new_P3_R1095_U83;
  assign new_P3_R1095_U414 = ~new_P3_R1095_U138;
  assign new_P3_R1095_U415 = ~new_P3_R1095_U299 | ~new_P3_R1095_U414;
  assign new_P3_R1095_U416 = ~new_P3_R1095_U138 | ~new_P3_R1095_U165;
  assign new_P3_R1095_U417 = ~new_P3_U3903 | ~new_P3_R1095_U82;
  assign new_P3_R1095_U418 = ~new_P3_U3064 | ~new_P3_R1095_U81;
  assign new_P3_R1095_U419 = ~new_P3_R1095_U139;
  assign new_P3_R1095_U420 = ~new_P3_R1095_U295 | ~new_P3_R1095_U419;
  assign new_P3_R1095_U421 = ~new_P3_R1095_U139 | ~new_P3_R1095_U166;
  assign new_P3_R1095_U422 = ~new_P3_U3904 | ~new_P3_R1095_U77;
  assign new_P3_R1095_U423 = ~new_P3_U3065 | ~new_P3_R1095_U74;
  assign new_P3_R1095_U424 = ~new_P3_R1095_U423 | ~new_P3_R1095_U422;
  assign new_P3_R1095_U425 = ~new_P3_U3905 | ~new_P3_R1095_U78;
  assign new_P3_R1095_U426 = ~new_P3_U3060 | ~new_P3_R1095_U75;
  assign new_P3_R1095_U427 = ~new_P3_R1095_U325 | ~new_P3_R1095_U92;
  assign new_P3_R1095_U428 = ~new_P3_R1095_U167 | ~new_P3_R1095_U317;
  assign new_P3_R1095_U429 = ~new_P3_U3906 | ~new_P3_R1095_U79;
  assign new_P3_R1095_U430 = ~new_P3_U3074 | ~new_P3_R1095_U76;
  assign new_P3_R1095_U431 = ~new_P3_R1095_U326 | ~new_P3_R1095_U169;
  assign new_P3_R1095_U432 = ~new_P3_R1095_U285 | ~new_P3_R1095_U168;
  assign new_P3_R1095_U433 = ~new_P3_U3907 | ~new_P3_R1095_U73;
  assign new_P3_R1095_U434 = ~new_P3_U3075 | ~new_P3_R1095_U72;
  assign new_P3_R1095_U435 = ~new_P3_R1095_U142;
  assign new_P3_R1095_U436 = ~new_P3_R1095_U281 | ~new_P3_R1095_U435;
  assign new_P3_R1095_U437 = ~new_P3_R1095_U142 | ~new_P3_R1095_U170;
  assign new_P3_R1095_U438 = ~new_P3_U3392 | ~new_P3_R1095_U31;
  assign new_P3_R1095_U439 = ~new_P3_U3077 | ~new_P3_R1095_U171;
  assign new_P3_R1095_U440 = ~new_P3_R1095_U143;
  assign new_P3_R1095_U441 = ~new_P3_R1095_U200 | ~new_P3_R1095_U440;
  assign new_P3_R1095_U442 = ~new_P3_R1095_U143 | ~new_P3_R1095_U172;
  assign new_P3_R1095_U443 = ~new_P3_U3445 | ~new_P3_R1095_U71;
  assign new_P3_R1095_U444 = ~new_P3_U3080 | ~new_P3_R1095_U70;
  assign new_P3_R1095_U445 = ~new_P3_R1095_U144;
  assign new_P3_R1095_U446 = ~new_P3_R1095_U277 | ~new_P3_R1095_U445;
  assign new_P3_R1095_U447 = ~new_P3_R1095_U144 | ~new_P3_R1095_U173;
  assign new_P3_R1095_U448 = ~new_P3_U3443 | ~new_P3_R1095_U69;
  assign new_P3_R1095_U449 = ~new_P3_U3081 | ~new_P3_R1095_U174;
  assign new_P3_R1095_U450 = ~new_P3_R1095_U145;
  assign new_P3_R1095_U451 = ~new_P3_R1095_U275 | ~new_P3_R1095_U450;
  assign new_P3_R1095_U452 = ~new_P3_R1095_U145 | ~new_P3_R1095_U175;
  assign new_P3_R1095_U453 = ~new_P3_U3440 | ~new_P3_R1095_U68;
  assign new_P3_R1095_U454 = ~new_P3_U3068 | ~new_P3_R1095_U67;
  assign new_P3_R1095_U455 = ~new_P3_R1095_U146;
  assign new_P3_R1095_U456 = ~new_P3_R1095_U271 | ~new_P3_R1095_U455;
  assign new_P3_R1095_U457 = ~new_P3_R1095_U146 | ~new_P3_R1095_U176;
  assign new_P3_R1095_U458 = ~new_P3_U3437 | ~new_P3_R1095_U63;
  assign new_P3_R1095_U459 = ~new_P3_U3072 | ~new_P3_R1095_U60;
  assign new_P3_R1095_U460 = ~new_P3_R1095_U459 | ~new_P3_R1095_U458;
  assign new_P3_R1095_U461 = ~new_P3_U3434 | ~new_P3_R1095_U64;
  assign new_P3_R1095_U462 = ~new_P3_U3073 | ~new_P3_R1095_U61;
  assign new_P3_R1095_U463 = ~new_P3_R1095_U336 | ~new_P3_R1095_U93;
  assign new_P3_R1095_U464 = ~new_P3_R1095_U177 | ~new_P3_R1095_U328;
  assign new_P3_R1095_U465 = ~new_P3_U3431 | ~new_P3_R1095_U65;
  assign new_P3_R1095_U466 = ~new_P3_U3078 | ~new_P3_R1095_U62;
  assign new_P3_R1095_U467 = ~new_P3_R1095_U337 | ~new_P3_R1095_U179;
  assign new_P3_R1095_U468 = ~new_P3_R1095_U261 | ~new_P3_R1095_U178;
  assign new_P3_R1095_U469 = ~new_P3_U3428 | ~new_P3_R1095_U59;
  assign new_P3_R1095_U470 = ~new_P3_U3079 | ~new_P3_R1095_U58;
  assign new_P3_R1095_U471 = ~new_P3_R1095_U149;
  assign new_P3_R1095_U472 = ~new_P3_R1095_U257 | ~new_P3_R1095_U471;
  assign new_P3_R1095_U473 = ~new_P3_R1095_U149 | ~new_P3_R1095_U180;
  assign new_P3_R1095_U474 = ~new_P3_U3425 | ~new_P3_R1095_U57;
  assign new_P3_R1095_U475 = ~new_P3_U3071 | ~new_P3_R1095_U56;
  assign new_P3_R1095_U476 = ~new_P3_R1095_U150;
  assign new_P3_R1095_U477 = ~new_P3_R1095_U253 | ~new_P3_R1095_U476;
  assign new_P3_R1095_U478 = ~new_P3_R1095_U150 | ~new_P3_R1095_U181;
  assign new_P3_R1095_U479 = ~new_P3_U3422 | ~new_P3_R1095_U53;
  assign new_P3_R1095_U480 = ~new_P3_U3062 | ~new_P3_R1095_U51;
  assign new_P3_R1095_U481 = ~new_P3_R1095_U480 | ~new_P3_R1095_U479;
  assign new_P3_R1095_U482 = ~new_P3_U3419 | ~new_P3_R1095_U54;
  assign new_P3_R1095_U483 = ~new_P3_U3061 | ~new_P3_R1095_U52;
  assign new_P3_R1095_U484 = ~new_P3_R1095_U347 | ~new_P3_R1095_U94;
  assign new_P3_R1095_U485 = ~new_P3_R1095_U182 | ~new_P3_R1095_U339;
  assign new_P3_R1212_U6 = ~new_P3_R1212_U176 | ~new_P3_R1212_U180;
  assign new_P3_R1212_U7 = ~new_P3_R1212_U9 | ~new_P3_R1212_U181;
  assign new_P3_R1212_U8 = ~P3_REG2_REG_0_;
  assign new_P3_R1212_U9 = ~P3_REG2_REG_0_ | ~new_P3_R1212_U48;
  assign new_P3_R1212_U10 = ~P3_REG2_REG_1_;
  assign new_P3_R1212_U11 = ~new_P3_U3391;
  assign new_P3_R1212_U12 = ~P3_REG2_REG_2_;
  assign new_P3_R1212_U13 = ~new_P3_U3394;
  assign new_P3_R1212_U14 = ~P3_REG2_REG_3_;
  assign new_P3_R1212_U15 = ~new_P3_U3397;
  assign new_P3_R1212_U16 = ~P3_REG2_REG_4_;
  assign new_P3_R1212_U17 = ~new_P3_U3400;
  assign new_P3_R1212_U18 = ~P3_REG2_REG_5_;
  assign new_P3_R1212_U19 = ~new_P3_U3403;
  assign new_P3_R1212_U20 = ~P3_REG2_REG_6_;
  assign new_P3_R1212_U21 = ~new_P3_U3406;
  assign new_P3_R1212_U22 = ~P3_REG2_REG_7_;
  assign new_P3_R1212_U23 = ~new_P3_U3409;
  assign new_P3_R1212_U24 = ~P3_REG2_REG_8_;
  assign new_P3_R1212_U25 = ~new_P3_U3412;
  assign new_P3_R1212_U26 = ~P3_REG2_REG_9_;
  assign new_P3_R1212_U27 = ~new_P3_U3415;
  assign new_P3_R1212_U28 = ~P3_REG2_REG_10_;
  assign new_P3_R1212_U29 = ~new_P3_U3418;
  assign new_P3_R1212_U30 = ~P3_REG2_REG_11_;
  assign new_P3_R1212_U31 = ~new_P3_U3421;
  assign new_P3_R1212_U32 = ~P3_REG2_REG_12_;
  assign new_P3_R1212_U33 = ~new_P3_U3424;
  assign new_P3_R1212_U34 = ~P3_REG2_REG_13_;
  assign new_P3_R1212_U35 = ~new_P3_U3427;
  assign new_P3_R1212_U36 = ~P3_REG2_REG_14_;
  assign new_P3_R1212_U37 = ~new_P3_U3430;
  assign new_P3_R1212_U38 = ~new_P3_R1212_U159 | ~new_P3_R1212_U158;
  assign new_P3_R1212_U39 = ~P3_REG2_REG_15_;
  assign new_P3_R1212_U40 = ~new_P3_U3433;
  assign new_P3_R1212_U41 = ~P3_REG2_REG_16_;
  assign new_P3_R1212_U42 = ~new_P3_U3436;
  assign new_P3_R1212_U43 = ~P3_REG2_REG_17_;
  assign new_P3_R1212_U44 = ~new_P3_U3439;
  assign new_P3_R1212_U45 = ~P3_REG2_REG_18_;
  assign new_P3_R1212_U46 = ~new_P3_U3442;
  assign new_P3_R1212_U47 = ~new_P3_R1212_U171 | ~new_P3_R1212_U170;
  assign new_P3_R1212_U48 = ~new_P3_U3386;
  assign new_P3_R1212_U49 = ~new_P3_R1212_U186 | ~new_P3_R1212_U185;
  assign new_P3_R1212_U50 = ~new_P3_R1212_U191 | ~new_P3_R1212_U190;
  assign new_P3_R1212_U51 = ~new_P3_R1212_U196 | ~new_P3_R1212_U195;
  assign new_P3_R1212_U52 = ~new_P3_R1212_U201 | ~new_P3_R1212_U200;
  assign new_P3_R1212_U53 = ~new_P3_R1212_U206 | ~new_P3_R1212_U205;
  assign new_P3_R1212_U54 = ~new_P3_R1212_U211 | ~new_P3_R1212_U210;
  assign new_P3_R1212_U55 = ~new_P3_R1212_U216 | ~new_P3_R1212_U215;
  assign new_P3_R1212_U56 = ~new_P3_R1212_U221 | ~new_P3_R1212_U220;
  assign new_P3_R1212_U57 = ~new_P3_R1212_U226 | ~new_P3_R1212_U225;
  assign new_P3_R1212_U58 = ~new_P3_R1212_U236 | ~new_P3_R1212_U235;
  assign new_P3_R1212_U59 = ~new_P3_R1212_U241 | ~new_P3_R1212_U240;
  assign new_P3_R1212_U60 = ~new_P3_R1212_U246 | ~new_P3_R1212_U245;
  assign new_P3_R1212_U61 = ~new_P3_R1212_U251 | ~new_P3_R1212_U250;
  assign new_P3_R1212_U62 = ~new_P3_R1212_U256 | ~new_P3_R1212_U255;
  assign new_P3_R1212_U63 = ~new_P3_R1212_U261 | ~new_P3_R1212_U260;
  assign new_P3_R1212_U64 = ~new_P3_R1212_U266 | ~new_P3_R1212_U265;
  assign new_P3_R1212_U65 = ~new_P3_R1212_U271 | ~new_P3_R1212_U270;
  assign new_P3_R1212_U66 = ~new_P3_R1212_U276 | ~new_P3_R1212_U275;
  assign new_P3_R1212_U67 = ~new_P3_R1212_U183 | ~new_P3_R1212_U182;
  assign new_P3_R1212_U68 = ~new_P3_R1212_U188 | ~new_P3_R1212_U187;
  assign new_P3_R1212_U69 = ~new_P3_R1212_U193 | ~new_P3_R1212_U192;
  assign new_P3_R1212_U70 = ~new_P3_R1212_U198 | ~new_P3_R1212_U197;
  assign new_P3_R1212_U71 = ~new_P3_R1212_U203 | ~new_P3_R1212_U202;
  assign new_P3_R1212_U72 = ~new_P3_R1212_U208 | ~new_P3_R1212_U207;
  assign new_P3_R1212_U73 = ~new_P3_R1212_U213 | ~new_P3_R1212_U212;
  assign new_P3_R1212_U74 = ~new_P3_R1212_U218 | ~new_P3_R1212_U217;
  assign new_P3_R1212_U75 = ~new_P3_R1212_U223 | ~new_P3_R1212_U222;
  assign new_P3_R1212_U76 = new_P3_R1212_U179 & new_P3_R1212_U228 & new_P3_R1212_U227;
  assign new_P3_R1212_U77 = new_P3_R1212_U175 & new_P3_R1212_U231;
  assign new_P3_R1212_U78 = ~new_P3_R1212_U233 | ~new_P3_R1212_U232;
  assign new_P3_R1212_U79 = ~new_P3_R1212_U238 | ~new_P3_R1212_U237;
  assign new_P3_R1212_U80 = ~new_P3_R1212_U243 | ~new_P3_R1212_U242;
  assign new_P3_R1212_U81 = ~new_P3_R1212_U248 | ~new_P3_R1212_U247;
  assign new_P3_R1212_U82 = ~new_P3_R1212_U253 | ~new_P3_R1212_U252;
  assign new_P3_R1212_U83 = ~new_P3_R1212_U258 | ~new_P3_R1212_U257;
  assign new_P3_R1212_U84 = ~new_P3_R1212_U263 | ~new_P3_R1212_U262;
  assign new_P3_R1212_U85 = ~new_P3_R1212_U268 | ~new_P3_R1212_U267;
  assign new_P3_R1212_U86 = ~new_P3_R1212_U273 | ~new_P3_R1212_U272;
  assign new_P3_R1212_U87 = ~new_P3_R1212_U135 | ~new_P3_R1212_U134;
  assign new_P3_R1212_U88 = ~new_P3_R1212_U131 | ~new_P3_R1212_U130;
  assign new_P3_R1212_U89 = ~new_P3_R1212_U127 | ~new_P3_R1212_U126;
  assign new_P3_R1212_U90 = ~new_P3_R1212_U123 | ~new_P3_R1212_U122;
  assign new_P3_R1212_U91 = ~new_P3_R1212_U119 | ~new_P3_R1212_U118;
  assign new_P3_R1212_U92 = ~new_P3_R1212_U115 | ~new_P3_R1212_U114;
  assign new_P3_R1212_U93 = ~new_P3_R1212_U111 | ~new_P3_R1212_U110;
  assign new_P3_R1212_U94 = ~new_P3_R1212_U107 | ~new_P3_R1212_U106;
  assign new_P3_R1212_U95 = ~P3_REG2_REG_19_;
  assign new_P3_R1212_U96 = ~new_P3_U3379;
  assign new_P3_R1212_U97 = ~new_P3_R1212_U167 | ~new_P3_R1212_U166;
  assign new_P3_R1212_U98 = ~new_P3_R1212_U163 | ~new_P3_R1212_U162;
  assign new_P3_R1212_U99 = ~new_P3_R1212_U155 | ~new_P3_R1212_U154;
  assign new_P3_R1212_U100 = ~new_P3_R1212_U151 | ~new_P3_R1212_U150;
  assign new_P3_R1212_U101 = ~new_P3_R1212_U147 | ~new_P3_R1212_U146;
  assign new_P3_R1212_U102 = ~new_P3_R1212_U143 | ~new_P3_R1212_U142;
  assign new_P3_R1212_U103 = ~new_P3_R1212_U139 | ~new_P3_R1212_U138;
  assign new_P3_R1212_U104 = ~new_P3_R1212_U9;
  assign new_P3_R1212_U105 = ~P3_REG2_REG_1_ | ~new_P3_R1212_U104;
  assign new_P3_R1212_U106 = ~new_P3_U3391 | ~new_P3_R1212_U105;
  assign new_P3_R1212_U107 = ~new_P3_R1212_U9 | ~new_P3_R1212_U10;
  assign new_P3_R1212_U108 = ~new_P3_R1212_U94;
  assign new_P3_R1212_U109 = ~P3_REG2_REG_2_ | ~new_P3_R1212_U13;
  assign new_P3_R1212_U110 = ~new_P3_R1212_U109 | ~new_P3_R1212_U94;
  assign new_P3_R1212_U111 = ~new_P3_U3394 | ~new_P3_R1212_U12;
  assign new_P3_R1212_U112 = ~new_P3_R1212_U93;
  assign new_P3_R1212_U113 = ~P3_REG2_REG_3_ | ~new_P3_R1212_U15;
  assign new_P3_R1212_U114 = ~new_P3_R1212_U113 | ~new_P3_R1212_U93;
  assign new_P3_R1212_U115 = ~new_P3_U3397 | ~new_P3_R1212_U14;
  assign new_P3_R1212_U116 = ~new_P3_R1212_U92;
  assign new_P3_R1212_U117 = ~P3_REG2_REG_4_ | ~new_P3_R1212_U17;
  assign new_P3_R1212_U118 = ~new_P3_R1212_U117 | ~new_P3_R1212_U92;
  assign new_P3_R1212_U119 = ~new_P3_U3400 | ~new_P3_R1212_U16;
  assign new_P3_R1212_U120 = ~new_P3_R1212_U91;
  assign new_P3_R1212_U121 = ~P3_REG2_REG_5_ | ~new_P3_R1212_U19;
  assign new_P3_R1212_U122 = ~new_P3_R1212_U121 | ~new_P3_R1212_U91;
  assign new_P3_R1212_U123 = ~new_P3_U3403 | ~new_P3_R1212_U18;
  assign new_P3_R1212_U124 = ~new_P3_R1212_U90;
  assign new_P3_R1212_U125 = ~P3_REG2_REG_6_ | ~new_P3_R1212_U21;
  assign new_P3_R1212_U126 = ~new_P3_R1212_U125 | ~new_P3_R1212_U90;
  assign new_P3_R1212_U127 = ~new_P3_U3406 | ~new_P3_R1212_U20;
  assign new_P3_R1212_U128 = ~new_P3_R1212_U89;
  assign new_P3_R1212_U129 = ~P3_REG2_REG_7_ | ~new_P3_R1212_U23;
  assign new_P3_R1212_U130 = ~new_P3_R1212_U129 | ~new_P3_R1212_U89;
  assign new_P3_R1212_U131 = ~new_P3_U3409 | ~new_P3_R1212_U22;
  assign new_P3_R1212_U132 = ~new_P3_R1212_U88;
  assign new_P3_R1212_U133 = ~P3_REG2_REG_8_ | ~new_P3_R1212_U25;
  assign new_P3_R1212_U134 = ~new_P3_R1212_U133 | ~new_P3_R1212_U88;
  assign new_P3_R1212_U135 = ~new_P3_U3412 | ~new_P3_R1212_U24;
  assign new_P3_R1212_U136 = ~new_P3_R1212_U87;
  assign new_P3_R1212_U137 = ~P3_REG2_REG_9_ | ~new_P3_R1212_U27;
  assign new_P3_R1212_U138 = ~new_P3_R1212_U137 | ~new_P3_R1212_U87;
  assign new_P3_R1212_U139 = ~new_P3_U3415 | ~new_P3_R1212_U26;
  assign new_P3_R1212_U140 = ~new_P3_R1212_U103;
  assign new_P3_R1212_U141 = ~P3_REG2_REG_10_ | ~new_P3_R1212_U29;
  assign new_P3_R1212_U142 = ~new_P3_R1212_U141 | ~new_P3_R1212_U103;
  assign new_P3_R1212_U143 = ~new_P3_U3418 | ~new_P3_R1212_U28;
  assign new_P3_R1212_U144 = ~new_P3_R1212_U102;
  assign new_P3_R1212_U145 = ~P3_REG2_REG_11_ | ~new_P3_R1212_U31;
  assign new_P3_R1212_U146 = ~new_P3_R1212_U145 | ~new_P3_R1212_U102;
  assign new_P3_R1212_U147 = ~new_P3_U3421 | ~new_P3_R1212_U30;
  assign new_P3_R1212_U148 = ~new_P3_R1212_U101;
  assign new_P3_R1212_U149 = ~P3_REG2_REG_12_ | ~new_P3_R1212_U33;
  assign new_P3_R1212_U150 = ~new_P3_R1212_U149 | ~new_P3_R1212_U101;
  assign new_P3_R1212_U151 = ~new_P3_U3424 | ~new_P3_R1212_U32;
  assign new_P3_R1212_U152 = ~new_P3_R1212_U100;
  assign new_P3_R1212_U153 = ~P3_REG2_REG_13_ | ~new_P3_R1212_U35;
  assign new_P3_R1212_U154 = ~new_P3_R1212_U153 | ~new_P3_R1212_U100;
  assign new_P3_R1212_U155 = ~new_P3_U3427 | ~new_P3_R1212_U34;
  assign new_P3_R1212_U156 = ~new_P3_R1212_U99;
  assign new_P3_R1212_U157 = ~P3_REG2_REG_14_ | ~new_P3_R1212_U37;
  assign new_P3_R1212_U158 = ~new_P3_R1212_U157 | ~new_P3_R1212_U99;
  assign new_P3_R1212_U159 = ~new_P3_U3430 | ~new_P3_R1212_U36;
  assign new_P3_R1212_U160 = ~new_P3_R1212_U38;
  assign new_P3_R1212_U161 = ~P3_REG2_REG_15_ | ~new_P3_R1212_U160;
  assign new_P3_R1212_U162 = ~new_P3_U3433 | ~new_P3_R1212_U161;
  assign new_P3_R1212_U163 = ~new_P3_R1212_U38 | ~new_P3_R1212_U39;
  assign new_P3_R1212_U164 = ~new_P3_R1212_U98;
  assign new_P3_R1212_U165 = ~P3_REG2_REG_16_ | ~new_P3_R1212_U42;
  assign new_P3_R1212_U166 = ~new_P3_R1212_U165 | ~new_P3_R1212_U98;
  assign new_P3_R1212_U167 = ~new_P3_U3436 | ~new_P3_R1212_U41;
  assign new_P3_R1212_U168 = ~new_P3_R1212_U97;
  assign new_P3_R1212_U169 = ~P3_REG2_REG_17_ | ~new_P3_R1212_U44;
  assign new_P3_R1212_U170 = ~new_P3_R1212_U169 | ~new_P3_R1212_U97;
  assign new_P3_R1212_U171 = ~new_P3_U3439 | ~new_P3_R1212_U43;
  assign new_P3_R1212_U172 = ~new_P3_R1212_U47;
  assign new_P3_R1212_U173 = ~new_P3_U3442 | ~new_P3_R1212_U45;
  assign new_P3_R1212_U174 = ~new_P3_R1212_U172 | ~new_P3_R1212_U173;
  assign new_P3_R1212_U175 = ~P3_REG2_REG_18_ | ~new_P3_R1212_U46;
  assign new_P3_R1212_U176 = ~new_P3_R1212_U77 | ~new_P3_R1212_U174;
  assign new_P3_R1212_U177 = ~P3_REG2_REG_18_ | ~new_P3_R1212_U46;
  assign new_P3_R1212_U178 = ~new_P3_R1212_U177 | ~new_P3_R1212_U47;
  assign new_P3_R1212_U179 = ~new_P3_U3442 | ~new_P3_R1212_U45;
  assign new_P3_R1212_U180 = ~new_P3_R1212_U76 | ~new_P3_R1212_U178;
  assign new_P3_R1212_U181 = ~new_P3_U3386 | ~new_P3_R1212_U8;
  assign new_P3_R1212_U182 = ~P3_REG2_REG_9_ | ~new_P3_R1212_U27;
  assign new_P3_R1212_U183 = ~new_P3_U3415 | ~new_P3_R1212_U26;
  assign new_P3_R1212_U184 = ~new_P3_R1212_U67;
  assign new_P3_R1212_U185 = ~new_P3_R1212_U136 | ~new_P3_R1212_U184;
  assign new_P3_R1212_U186 = ~new_P3_R1212_U67 | ~new_P3_R1212_U87;
  assign new_P3_R1212_U187 = ~P3_REG2_REG_8_ | ~new_P3_R1212_U25;
  assign new_P3_R1212_U188 = ~new_P3_U3412 | ~new_P3_R1212_U24;
  assign new_P3_R1212_U189 = ~new_P3_R1212_U68;
  assign new_P3_R1212_U190 = ~new_P3_R1212_U132 | ~new_P3_R1212_U189;
  assign new_P3_R1212_U191 = ~new_P3_R1212_U68 | ~new_P3_R1212_U88;
  assign new_P3_R1212_U192 = ~P3_REG2_REG_7_ | ~new_P3_R1212_U23;
  assign new_P3_R1212_U193 = ~new_P3_U3409 | ~new_P3_R1212_U22;
  assign new_P3_R1212_U194 = ~new_P3_R1212_U69;
  assign new_P3_R1212_U195 = ~new_P3_R1212_U128 | ~new_P3_R1212_U194;
  assign new_P3_R1212_U196 = ~new_P3_R1212_U69 | ~new_P3_R1212_U89;
  assign new_P3_R1212_U197 = ~P3_REG2_REG_6_ | ~new_P3_R1212_U21;
  assign new_P3_R1212_U198 = ~new_P3_U3406 | ~new_P3_R1212_U20;
  assign new_P3_R1212_U199 = ~new_P3_R1212_U70;
  assign new_P3_R1212_U200 = ~new_P3_R1212_U124 | ~new_P3_R1212_U199;
  assign new_P3_R1212_U201 = ~new_P3_R1212_U70 | ~new_P3_R1212_U90;
  assign new_P3_R1212_U202 = ~P3_REG2_REG_5_ | ~new_P3_R1212_U19;
  assign new_P3_R1212_U203 = ~new_P3_U3403 | ~new_P3_R1212_U18;
  assign new_P3_R1212_U204 = ~new_P3_R1212_U71;
  assign new_P3_R1212_U205 = ~new_P3_R1212_U120 | ~new_P3_R1212_U204;
  assign new_P3_R1212_U206 = ~new_P3_R1212_U71 | ~new_P3_R1212_U91;
  assign new_P3_R1212_U207 = ~P3_REG2_REG_4_ | ~new_P3_R1212_U17;
  assign new_P3_R1212_U208 = ~new_P3_U3400 | ~new_P3_R1212_U16;
  assign new_P3_R1212_U209 = ~new_P3_R1212_U72;
  assign new_P3_R1212_U210 = ~new_P3_R1212_U116 | ~new_P3_R1212_U209;
  assign new_P3_R1212_U211 = ~new_P3_R1212_U72 | ~new_P3_R1212_U92;
  assign new_P3_R1212_U212 = ~P3_REG2_REG_3_ | ~new_P3_R1212_U15;
  assign new_P3_R1212_U213 = ~new_P3_U3397 | ~new_P3_R1212_U14;
  assign new_P3_R1212_U214 = ~new_P3_R1212_U73;
  assign new_P3_R1212_U215 = ~new_P3_R1212_U112 | ~new_P3_R1212_U214;
  assign new_P3_R1212_U216 = ~new_P3_R1212_U73 | ~new_P3_R1212_U93;
  assign new_P3_R1212_U217 = ~P3_REG2_REG_2_ | ~new_P3_R1212_U13;
  assign new_P3_R1212_U218 = ~new_P3_U3394 | ~new_P3_R1212_U12;
  assign new_P3_R1212_U219 = ~new_P3_R1212_U74;
  assign new_P3_R1212_U220 = ~new_P3_R1212_U108 | ~new_P3_R1212_U219;
  assign new_P3_R1212_U221 = ~new_P3_R1212_U74 | ~new_P3_R1212_U94;
  assign new_P3_R1212_U222 = ~new_P3_R1212_U104 | ~new_P3_R1212_U10;
  assign new_P3_R1212_U223 = ~P3_REG2_REG_1_ | ~new_P3_R1212_U9;
  assign new_P3_R1212_U224 = ~new_P3_R1212_U75;
  assign new_P3_R1212_U225 = ~new_P3_R1212_U224 | ~new_P3_U3391;
  assign new_P3_R1212_U226 = ~new_P3_R1212_U75 | ~new_P3_R1212_U11;
  assign new_P3_R1212_U227 = ~P3_REG2_REG_19_ | ~new_P3_R1212_U96;
  assign new_P3_R1212_U228 = ~new_P3_U3379 | ~new_P3_R1212_U95;
  assign new_P3_R1212_U229 = ~P3_REG2_REG_19_ | ~new_P3_R1212_U96;
  assign new_P3_R1212_U230 = ~new_P3_U3379 | ~new_P3_R1212_U95;
  assign new_P3_R1212_U231 = ~new_P3_R1212_U230 | ~new_P3_R1212_U229;
  assign new_P3_R1212_U232 = ~P3_REG2_REG_18_ | ~new_P3_R1212_U46;
  assign new_P3_R1212_U233 = ~new_P3_U3442 | ~new_P3_R1212_U45;
  assign new_P3_R1212_U234 = ~new_P3_R1212_U78;
  assign new_P3_R1212_U235 = ~new_P3_R1212_U234 | ~new_P3_R1212_U172;
  assign new_P3_R1212_U236 = ~new_P3_R1212_U78 | ~new_P3_R1212_U47;
  assign new_P3_R1212_U237 = ~P3_REG2_REG_17_ | ~new_P3_R1212_U44;
  assign new_P3_R1212_U238 = ~new_P3_U3439 | ~new_P3_R1212_U43;
  assign new_P3_R1212_U239 = ~new_P3_R1212_U79;
  assign new_P3_R1212_U240 = ~new_P3_R1212_U168 | ~new_P3_R1212_U239;
  assign new_P3_R1212_U241 = ~new_P3_R1212_U79 | ~new_P3_R1212_U97;
  assign new_P3_R1212_U242 = ~P3_REG2_REG_16_ | ~new_P3_R1212_U42;
  assign new_P3_R1212_U243 = ~new_P3_U3436 | ~new_P3_R1212_U41;
  assign new_P3_R1212_U244 = ~new_P3_R1212_U80;
  assign new_P3_R1212_U245 = ~new_P3_R1212_U164 | ~new_P3_R1212_U244;
  assign new_P3_R1212_U246 = ~new_P3_R1212_U80 | ~new_P3_R1212_U98;
  assign new_P3_R1212_U247 = ~new_P3_U3433 | ~new_P3_R1212_U39;
  assign new_P3_R1212_U248 = ~P3_REG2_REG_15_ | ~new_P3_R1212_U40;
  assign new_P3_R1212_U249 = ~new_P3_R1212_U81;
  assign new_P3_R1212_U250 = ~new_P3_R1212_U249 | ~new_P3_R1212_U160;
  assign new_P3_R1212_U251 = ~new_P3_R1212_U81 | ~new_P3_R1212_U38;
  assign new_P3_R1212_U252 = ~P3_REG2_REG_14_ | ~new_P3_R1212_U37;
  assign new_P3_R1212_U253 = ~new_P3_U3430 | ~new_P3_R1212_U36;
  assign new_P3_R1212_U254 = ~new_P3_R1212_U82;
  assign new_P3_R1212_U255 = ~new_P3_R1212_U156 | ~new_P3_R1212_U254;
  assign new_P3_R1212_U256 = ~new_P3_R1212_U82 | ~new_P3_R1212_U99;
  assign new_P3_R1212_U257 = ~P3_REG2_REG_13_ | ~new_P3_R1212_U35;
  assign new_P3_R1212_U258 = ~new_P3_U3427 | ~new_P3_R1212_U34;
  assign new_P3_R1212_U259 = ~new_P3_R1212_U83;
  assign new_P3_R1212_U260 = ~new_P3_R1212_U152 | ~new_P3_R1212_U259;
  assign new_P3_R1212_U261 = ~new_P3_R1212_U83 | ~new_P3_R1212_U100;
  assign new_P3_R1212_U262 = ~P3_REG2_REG_12_ | ~new_P3_R1212_U33;
  assign new_P3_R1212_U263 = ~new_P3_U3424 | ~new_P3_R1212_U32;
  assign new_P3_R1212_U264 = ~new_P3_R1212_U84;
  assign new_P3_R1212_U265 = ~new_P3_R1212_U148 | ~new_P3_R1212_U264;
  assign new_P3_R1212_U266 = ~new_P3_R1212_U84 | ~new_P3_R1212_U101;
  assign new_P3_R1212_U267 = ~P3_REG2_REG_11_ | ~new_P3_R1212_U31;
  assign new_P3_R1212_U268 = ~new_P3_U3421 | ~new_P3_R1212_U30;
  assign new_P3_R1212_U269 = ~new_P3_R1212_U85;
  assign new_P3_R1212_U270 = ~new_P3_R1212_U144 | ~new_P3_R1212_U269;
  assign new_P3_R1212_U271 = ~new_P3_R1212_U85 | ~new_P3_R1212_U102;
  assign new_P3_R1212_U272 = ~P3_REG2_REG_10_ | ~new_P3_R1212_U29;
  assign new_P3_R1212_U273 = ~new_P3_U3418 | ~new_P3_R1212_U28;
  assign new_P3_R1212_U274 = ~new_P3_R1212_U86;
  assign new_P3_R1212_U275 = ~new_P3_R1212_U140 | ~new_P3_R1212_U274;
  assign new_P3_R1212_U276 = ~new_P3_R1212_U86 | ~new_P3_R1212_U103;
  assign new_P3_R1209_U6 = ~new_P3_R1209_U176 | ~new_P3_R1209_U180;
  assign new_P3_R1209_U7 = ~new_P3_R1209_U9 | ~new_P3_R1209_U181;
  assign new_P3_R1209_U8 = ~P3_REG1_REG_0_;
  assign new_P3_R1209_U9 = ~P3_REG1_REG_0_ | ~new_P3_R1209_U48;
  assign new_P3_R1209_U10 = ~P3_REG1_REG_1_;
  assign new_P3_R1209_U11 = ~new_P3_U3391;
  assign new_P3_R1209_U12 = ~P3_REG1_REG_2_;
  assign new_P3_R1209_U13 = ~new_P3_U3394;
  assign new_P3_R1209_U14 = ~P3_REG1_REG_3_;
  assign new_P3_R1209_U15 = ~new_P3_U3397;
  assign new_P3_R1209_U16 = ~P3_REG1_REG_4_;
  assign new_P3_R1209_U17 = ~new_P3_U3400;
  assign new_P3_R1209_U18 = ~P3_REG1_REG_5_;
  assign new_P3_R1209_U19 = ~new_P3_U3403;
  assign new_P3_R1209_U20 = ~P3_REG1_REG_6_;
  assign new_P3_R1209_U21 = ~new_P3_U3406;
  assign new_P3_R1209_U22 = ~P3_REG1_REG_7_;
  assign new_P3_R1209_U23 = ~new_P3_U3409;
  assign new_P3_R1209_U24 = ~P3_REG1_REG_8_;
  assign new_P3_R1209_U25 = ~new_P3_U3412;
  assign new_P3_R1209_U26 = ~P3_REG1_REG_9_;
  assign new_P3_R1209_U27 = ~new_P3_U3415;
  assign new_P3_R1209_U28 = ~P3_REG1_REG_10_;
  assign new_P3_R1209_U29 = ~new_P3_U3418;
  assign new_P3_R1209_U30 = ~P3_REG1_REG_11_;
  assign new_P3_R1209_U31 = ~new_P3_U3421;
  assign new_P3_R1209_U32 = ~P3_REG1_REG_12_;
  assign new_P3_R1209_U33 = ~new_P3_U3424;
  assign new_P3_R1209_U34 = ~P3_REG1_REG_13_;
  assign new_P3_R1209_U35 = ~new_P3_U3427;
  assign new_P3_R1209_U36 = ~P3_REG1_REG_14_;
  assign new_P3_R1209_U37 = ~new_P3_U3430;
  assign new_P3_R1209_U38 = ~new_P3_R1209_U159 | ~new_P3_R1209_U158;
  assign new_P3_R1209_U39 = ~P3_REG1_REG_15_;
  assign new_P3_R1209_U40 = ~new_P3_U3433;
  assign new_P3_R1209_U41 = ~P3_REG1_REG_16_;
  assign new_P3_R1209_U42 = ~new_P3_U3436;
  assign new_P3_R1209_U43 = ~P3_REG1_REG_17_;
  assign new_P3_R1209_U44 = ~new_P3_U3439;
  assign new_P3_R1209_U45 = ~P3_REG1_REG_18_;
  assign new_P3_R1209_U46 = ~new_P3_U3442;
  assign new_P3_R1209_U47 = ~new_P3_R1209_U171 | ~new_P3_R1209_U170;
  assign new_P3_R1209_U48 = ~new_P3_U3386;
  assign new_P3_R1209_U49 = ~new_P3_R1209_U186 | ~new_P3_R1209_U185;
  assign new_P3_R1209_U50 = ~new_P3_R1209_U191 | ~new_P3_R1209_U190;
  assign new_P3_R1209_U51 = ~new_P3_R1209_U196 | ~new_P3_R1209_U195;
  assign new_P3_R1209_U52 = ~new_P3_R1209_U201 | ~new_P3_R1209_U200;
  assign new_P3_R1209_U53 = ~new_P3_R1209_U206 | ~new_P3_R1209_U205;
  assign new_P3_R1209_U54 = ~new_P3_R1209_U211 | ~new_P3_R1209_U210;
  assign new_P3_R1209_U55 = ~new_P3_R1209_U216 | ~new_P3_R1209_U215;
  assign new_P3_R1209_U56 = ~new_P3_R1209_U221 | ~new_P3_R1209_U220;
  assign new_P3_R1209_U57 = ~new_P3_R1209_U226 | ~new_P3_R1209_U225;
  assign new_P3_R1209_U58 = ~new_P3_R1209_U236 | ~new_P3_R1209_U235;
  assign new_P3_R1209_U59 = ~new_P3_R1209_U241 | ~new_P3_R1209_U240;
  assign new_P3_R1209_U60 = ~new_P3_R1209_U246 | ~new_P3_R1209_U245;
  assign new_P3_R1209_U61 = ~new_P3_R1209_U251 | ~new_P3_R1209_U250;
  assign new_P3_R1209_U62 = ~new_P3_R1209_U256 | ~new_P3_R1209_U255;
  assign new_P3_R1209_U63 = ~new_P3_R1209_U261 | ~new_P3_R1209_U260;
  assign new_P3_R1209_U64 = ~new_P3_R1209_U266 | ~new_P3_R1209_U265;
  assign new_P3_R1209_U65 = ~new_P3_R1209_U271 | ~new_P3_R1209_U270;
  assign new_P3_R1209_U66 = ~new_P3_R1209_U276 | ~new_P3_R1209_U275;
  assign new_P3_R1209_U67 = ~new_P3_R1209_U183 | ~new_P3_R1209_U182;
  assign new_P3_R1209_U68 = ~new_P3_R1209_U188 | ~new_P3_R1209_U187;
  assign new_P3_R1209_U69 = ~new_P3_R1209_U193 | ~new_P3_R1209_U192;
  assign new_P3_R1209_U70 = ~new_P3_R1209_U198 | ~new_P3_R1209_U197;
  assign new_P3_R1209_U71 = ~new_P3_R1209_U203 | ~new_P3_R1209_U202;
  assign new_P3_R1209_U72 = ~new_P3_R1209_U208 | ~new_P3_R1209_U207;
  assign new_P3_R1209_U73 = ~new_P3_R1209_U213 | ~new_P3_R1209_U212;
  assign new_P3_R1209_U74 = ~new_P3_R1209_U218 | ~new_P3_R1209_U217;
  assign new_P3_R1209_U75 = ~new_P3_R1209_U223 | ~new_P3_R1209_U222;
  assign new_P3_R1209_U76 = new_P3_R1209_U179 & new_P3_R1209_U228 & new_P3_R1209_U227;
  assign new_P3_R1209_U77 = new_P3_R1209_U175 & new_P3_R1209_U231;
  assign new_P3_R1209_U78 = ~new_P3_R1209_U233 | ~new_P3_R1209_U232;
  assign new_P3_R1209_U79 = ~new_P3_R1209_U238 | ~new_P3_R1209_U237;
  assign new_P3_R1209_U80 = ~new_P3_R1209_U243 | ~new_P3_R1209_U242;
  assign new_P3_R1209_U81 = ~new_P3_R1209_U248 | ~new_P3_R1209_U247;
  assign new_P3_R1209_U82 = ~new_P3_R1209_U253 | ~new_P3_R1209_U252;
  assign new_P3_R1209_U83 = ~new_P3_R1209_U258 | ~new_P3_R1209_U257;
  assign new_P3_R1209_U84 = ~new_P3_R1209_U263 | ~new_P3_R1209_U262;
  assign new_P3_R1209_U85 = ~new_P3_R1209_U268 | ~new_P3_R1209_U267;
  assign new_P3_R1209_U86 = ~new_P3_R1209_U273 | ~new_P3_R1209_U272;
  assign new_P3_R1209_U87 = ~new_P3_R1209_U135 | ~new_P3_R1209_U134;
  assign new_P3_R1209_U88 = ~new_P3_R1209_U131 | ~new_P3_R1209_U130;
  assign new_P3_R1209_U89 = ~new_P3_R1209_U127 | ~new_P3_R1209_U126;
  assign new_P3_R1209_U90 = ~new_P3_R1209_U123 | ~new_P3_R1209_U122;
  assign new_P3_R1209_U91 = ~new_P3_R1209_U119 | ~new_P3_R1209_U118;
  assign new_P3_R1209_U92 = ~new_P3_R1209_U115 | ~new_P3_R1209_U114;
  assign new_P3_R1209_U93 = ~new_P3_R1209_U111 | ~new_P3_R1209_U110;
  assign new_P3_R1209_U94 = ~new_P3_R1209_U107 | ~new_P3_R1209_U106;
  assign new_P3_R1209_U95 = ~P3_REG1_REG_19_;
  assign new_P3_R1209_U96 = ~new_P3_U3379;
  assign new_P3_R1209_U97 = ~new_P3_R1209_U167 | ~new_P3_R1209_U166;
  assign new_P3_R1209_U98 = ~new_P3_R1209_U163 | ~new_P3_R1209_U162;
  assign new_P3_R1209_U99 = ~new_P3_R1209_U155 | ~new_P3_R1209_U154;
  assign new_P3_R1209_U100 = ~new_P3_R1209_U151 | ~new_P3_R1209_U150;
  assign new_P3_R1209_U101 = ~new_P3_R1209_U147 | ~new_P3_R1209_U146;
  assign new_P3_R1209_U102 = ~new_P3_R1209_U143 | ~new_P3_R1209_U142;
  assign new_P3_R1209_U103 = ~new_P3_R1209_U139 | ~new_P3_R1209_U138;
  assign new_P3_R1209_U104 = ~new_P3_R1209_U9;
  assign new_P3_R1209_U105 = ~P3_REG1_REG_1_ | ~new_P3_R1209_U104;
  assign new_P3_R1209_U106 = ~new_P3_U3391 | ~new_P3_R1209_U105;
  assign new_P3_R1209_U107 = ~new_P3_R1209_U9 | ~new_P3_R1209_U10;
  assign new_P3_R1209_U108 = ~new_P3_R1209_U94;
  assign new_P3_R1209_U109 = ~P3_REG1_REG_2_ | ~new_P3_R1209_U13;
  assign new_P3_R1209_U110 = ~new_P3_R1209_U109 | ~new_P3_R1209_U94;
  assign new_P3_R1209_U111 = ~new_P3_U3394 | ~new_P3_R1209_U12;
  assign new_P3_R1209_U112 = ~new_P3_R1209_U93;
  assign new_P3_R1209_U113 = ~P3_REG1_REG_3_ | ~new_P3_R1209_U15;
  assign new_P3_R1209_U114 = ~new_P3_R1209_U113 | ~new_P3_R1209_U93;
  assign new_P3_R1209_U115 = ~new_P3_U3397 | ~new_P3_R1209_U14;
  assign new_P3_R1209_U116 = ~new_P3_R1209_U92;
  assign new_P3_R1209_U117 = ~P3_REG1_REG_4_ | ~new_P3_R1209_U17;
  assign new_P3_R1209_U118 = ~new_P3_R1209_U117 | ~new_P3_R1209_U92;
  assign new_P3_R1209_U119 = ~new_P3_U3400 | ~new_P3_R1209_U16;
  assign new_P3_R1209_U120 = ~new_P3_R1209_U91;
  assign new_P3_R1209_U121 = ~P3_REG1_REG_5_ | ~new_P3_R1209_U19;
  assign new_P3_R1209_U122 = ~new_P3_R1209_U121 | ~new_P3_R1209_U91;
  assign new_P3_R1209_U123 = ~new_P3_U3403 | ~new_P3_R1209_U18;
  assign new_P3_R1209_U124 = ~new_P3_R1209_U90;
  assign new_P3_R1209_U125 = ~P3_REG1_REG_6_ | ~new_P3_R1209_U21;
  assign new_P3_R1209_U126 = ~new_P3_R1209_U125 | ~new_P3_R1209_U90;
  assign new_P3_R1209_U127 = ~new_P3_U3406 | ~new_P3_R1209_U20;
  assign new_P3_R1209_U128 = ~new_P3_R1209_U89;
  assign new_P3_R1209_U129 = ~P3_REG1_REG_7_ | ~new_P3_R1209_U23;
  assign new_P3_R1209_U130 = ~new_P3_R1209_U129 | ~new_P3_R1209_U89;
  assign new_P3_R1209_U131 = ~new_P3_U3409 | ~new_P3_R1209_U22;
  assign new_P3_R1209_U132 = ~new_P3_R1209_U88;
  assign new_P3_R1209_U133 = ~P3_REG1_REG_8_ | ~new_P3_R1209_U25;
  assign new_P3_R1209_U134 = ~new_P3_R1209_U133 | ~new_P3_R1209_U88;
  assign new_P3_R1209_U135 = ~new_P3_U3412 | ~new_P3_R1209_U24;
  assign new_P3_R1209_U136 = ~new_P3_R1209_U87;
  assign new_P3_R1209_U137 = ~P3_REG1_REG_9_ | ~new_P3_R1209_U27;
  assign new_P3_R1209_U138 = ~new_P3_R1209_U137 | ~new_P3_R1209_U87;
  assign new_P3_R1209_U139 = ~new_P3_U3415 | ~new_P3_R1209_U26;
  assign new_P3_R1209_U140 = ~new_P3_R1209_U103;
  assign new_P3_R1209_U141 = ~P3_REG1_REG_10_ | ~new_P3_R1209_U29;
  assign new_P3_R1209_U142 = ~new_P3_R1209_U141 | ~new_P3_R1209_U103;
  assign new_P3_R1209_U143 = ~new_P3_U3418 | ~new_P3_R1209_U28;
  assign new_P3_R1209_U144 = ~new_P3_R1209_U102;
  assign new_P3_R1209_U145 = ~P3_REG1_REG_11_ | ~new_P3_R1209_U31;
  assign new_P3_R1209_U146 = ~new_P3_R1209_U145 | ~new_P3_R1209_U102;
  assign new_P3_R1209_U147 = ~new_P3_U3421 | ~new_P3_R1209_U30;
  assign new_P3_R1209_U148 = ~new_P3_R1209_U101;
  assign new_P3_R1209_U149 = ~P3_REG1_REG_12_ | ~new_P3_R1209_U33;
  assign new_P3_R1209_U150 = ~new_P3_R1209_U149 | ~new_P3_R1209_U101;
  assign new_P3_R1209_U151 = ~new_P3_U3424 | ~new_P3_R1209_U32;
  assign new_P3_R1209_U152 = ~new_P3_R1209_U100;
  assign new_P3_R1209_U153 = ~P3_REG1_REG_13_ | ~new_P3_R1209_U35;
  assign new_P3_R1209_U154 = ~new_P3_R1209_U153 | ~new_P3_R1209_U100;
  assign new_P3_R1209_U155 = ~new_P3_U3427 | ~new_P3_R1209_U34;
  assign new_P3_R1209_U156 = ~new_P3_R1209_U99;
  assign new_P3_R1209_U157 = ~P3_REG1_REG_14_ | ~new_P3_R1209_U37;
  assign new_P3_R1209_U158 = ~new_P3_R1209_U157 | ~new_P3_R1209_U99;
  assign new_P3_R1209_U159 = ~new_P3_U3430 | ~new_P3_R1209_U36;
  assign new_P3_R1209_U160 = ~new_P3_R1209_U38;
  assign new_P3_R1209_U161 = ~P3_REG1_REG_15_ | ~new_P3_R1209_U160;
  assign new_P3_R1209_U162 = ~new_P3_U3433 | ~new_P3_R1209_U161;
  assign new_P3_R1209_U163 = ~new_P3_R1209_U38 | ~new_P3_R1209_U39;
  assign new_P3_R1209_U164 = ~new_P3_R1209_U98;
  assign new_P3_R1209_U165 = ~P3_REG1_REG_16_ | ~new_P3_R1209_U42;
  assign new_P3_R1209_U166 = ~new_P3_R1209_U165 | ~new_P3_R1209_U98;
  assign new_P3_R1209_U167 = ~new_P3_U3436 | ~new_P3_R1209_U41;
  assign new_P3_R1209_U168 = ~new_P3_R1209_U97;
  assign new_P3_R1209_U169 = ~P3_REG1_REG_17_ | ~new_P3_R1209_U44;
  assign new_P3_R1209_U170 = ~new_P3_R1209_U169 | ~new_P3_R1209_U97;
  assign new_P3_R1209_U171 = ~new_P3_U3439 | ~new_P3_R1209_U43;
  assign new_P3_R1209_U172 = ~new_P3_R1209_U47;
  assign new_P3_R1209_U173 = ~new_P3_U3442 | ~new_P3_R1209_U45;
  assign new_P3_R1209_U174 = ~new_P3_R1209_U172 | ~new_P3_R1209_U173;
  assign new_P3_R1209_U175 = ~P3_REG1_REG_18_ | ~new_P3_R1209_U46;
  assign new_P3_R1209_U176 = ~new_P3_R1209_U77 | ~new_P3_R1209_U174;
  assign new_P3_R1209_U177 = ~P3_REG1_REG_18_ | ~new_P3_R1209_U46;
  assign new_P3_R1209_U178 = ~new_P3_R1209_U177 | ~new_P3_R1209_U47;
  assign new_P3_R1209_U179 = ~new_P3_U3442 | ~new_P3_R1209_U45;
  assign new_P3_R1209_U180 = ~new_P3_R1209_U76 | ~new_P3_R1209_U178;
  assign new_P3_R1209_U181 = ~new_P3_U3386 | ~new_P3_R1209_U8;
  assign new_P3_R1209_U182 = ~P3_REG1_REG_9_ | ~new_P3_R1209_U27;
  assign new_P3_R1209_U183 = ~new_P3_U3415 | ~new_P3_R1209_U26;
  assign new_P3_R1209_U184 = ~new_P3_R1209_U67;
  assign new_P3_R1209_U185 = ~new_P3_R1209_U136 | ~new_P3_R1209_U184;
  assign new_P3_R1209_U186 = ~new_P3_R1209_U67 | ~new_P3_R1209_U87;
  assign new_P3_R1209_U187 = ~P3_REG1_REG_8_ | ~new_P3_R1209_U25;
  assign new_P3_R1209_U188 = ~new_P3_U3412 | ~new_P3_R1209_U24;
  assign new_P3_R1209_U189 = ~new_P3_R1209_U68;
  assign new_P3_R1209_U190 = ~new_P3_R1209_U132 | ~new_P3_R1209_U189;
  assign new_P3_R1209_U191 = ~new_P3_R1209_U68 | ~new_P3_R1209_U88;
  assign new_P3_R1209_U192 = ~P3_REG1_REG_7_ | ~new_P3_R1209_U23;
  assign new_P3_R1209_U193 = ~new_P3_U3409 | ~new_P3_R1209_U22;
  assign new_P3_R1209_U194 = ~new_P3_R1209_U69;
  assign new_P3_R1209_U195 = ~new_P3_R1209_U128 | ~new_P3_R1209_U194;
  assign new_P3_R1209_U196 = ~new_P3_R1209_U69 | ~new_P3_R1209_U89;
  assign new_P3_R1209_U197 = ~P3_REG1_REG_6_ | ~new_P3_R1209_U21;
  assign new_P3_R1209_U198 = ~new_P3_U3406 | ~new_P3_R1209_U20;
  assign new_P3_R1209_U199 = ~new_P3_R1209_U70;
  assign new_P3_R1209_U200 = ~new_P3_R1209_U124 | ~new_P3_R1209_U199;
  assign new_P3_R1209_U201 = ~new_P3_R1209_U70 | ~new_P3_R1209_U90;
  assign new_P3_R1209_U202 = ~P3_REG1_REG_5_ | ~new_P3_R1209_U19;
  assign new_P3_R1209_U203 = ~new_P3_U3403 | ~new_P3_R1209_U18;
  assign new_P3_R1209_U204 = ~new_P3_R1209_U71;
  assign new_P3_R1209_U205 = ~new_P3_R1209_U120 | ~new_P3_R1209_U204;
  assign new_P3_R1209_U206 = ~new_P3_R1209_U71 | ~new_P3_R1209_U91;
  assign new_P3_R1209_U207 = ~P3_REG1_REG_4_ | ~new_P3_R1209_U17;
  assign new_P3_R1209_U208 = ~new_P3_U3400 | ~new_P3_R1209_U16;
  assign new_P3_R1209_U209 = ~new_P3_R1209_U72;
  assign new_P3_R1209_U210 = ~new_P3_R1209_U116 | ~new_P3_R1209_U209;
  assign new_P3_R1209_U211 = ~new_P3_R1209_U72 | ~new_P3_R1209_U92;
  assign new_P3_R1209_U212 = ~P3_REG1_REG_3_ | ~new_P3_R1209_U15;
  assign new_P3_R1209_U213 = ~new_P3_U3397 | ~new_P3_R1209_U14;
  assign new_P3_R1209_U214 = ~new_P3_R1209_U73;
  assign new_P3_R1209_U215 = ~new_P3_R1209_U112 | ~new_P3_R1209_U214;
  assign new_P3_R1209_U216 = ~new_P3_R1209_U73 | ~new_P3_R1209_U93;
  assign new_P3_R1209_U217 = ~P3_REG1_REG_2_ | ~new_P3_R1209_U13;
  assign new_P3_R1209_U218 = ~new_P3_U3394 | ~new_P3_R1209_U12;
  assign new_P3_R1209_U219 = ~new_P3_R1209_U74;
  assign new_P3_R1209_U220 = ~new_P3_R1209_U108 | ~new_P3_R1209_U219;
  assign new_P3_R1209_U221 = ~new_P3_R1209_U74 | ~new_P3_R1209_U94;
  assign new_P3_R1209_U222 = ~new_P3_R1209_U104 | ~new_P3_R1209_U10;
  assign new_P3_R1209_U223 = ~P3_REG1_REG_1_ | ~new_P3_R1209_U9;
  assign new_P3_R1209_U224 = ~new_P3_R1209_U75;
  assign new_P3_R1209_U225 = ~new_P3_R1209_U224 | ~new_P3_U3391;
  assign new_P3_R1209_U226 = ~new_P3_R1209_U75 | ~new_P3_R1209_U11;
  assign new_P3_R1209_U227 = ~P3_REG1_REG_19_ | ~new_P3_R1209_U96;
  assign new_P3_R1209_U228 = ~new_P3_U3379 | ~new_P3_R1209_U95;
  assign new_P3_R1209_U229 = ~P3_REG1_REG_19_ | ~new_P3_R1209_U96;
  assign new_P3_R1209_U230 = ~new_P3_U3379 | ~new_P3_R1209_U95;
  assign new_P3_R1209_U231 = ~new_P3_R1209_U230 | ~new_P3_R1209_U229;
  assign new_P3_R1209_U232 = ~P3_REG1_REG_18_ | ~new_P3_R1209_U46;
  assign new_P3_R1209_U233 = ~new_P3_U3442 | ~new_P3_R1209_U45;
  assign new_P3_R1209_U234 = ~new_P3_R1209_U78;
  assign new_P3_R1209_U235 = ~new_P3_R1209_U234 | ~new_P3_R1209_U172;
  assign new_P3_R1209_U236 = ~new_P3_R1209_U78 | ~new_P3_R1209_U47;
  assign new_P3_R1209_U237 = ~P3_REG1_REG_17_ | ~new_P3_R1209_U44;
  assign new_P3_R1209_U238 = ~new_P3_U3439 | ~new_P3_R1209_U43;
  assign new_P3_R1209_U239 = ~new_P3_R1209_U79;
  assign new_P3_R1209_U240 = ~new_P3_R1209_U168 | ~new_P3_R1209_U239;
  assign new_P3_R1209_U241 = ~new_P3_R1209_U79 | ~new_P3_R1209_U97;
  assign new_P3_R1209_U242 = ~P3_REG1_REG_16_ | ~new_P3_R1209_U42;
  assign new_P3_R1209_U243 = ~new_P3_U3436 | ~new_P3_R1209_U41;
  assign new_P3_R1209_U244 = ~new_P3_R1209_U80;
  assign new_P3_R1209_U245 = ~new_P3_R1209_U164 | ~new_P3_R1209_U244;
  assign new_P3_R1209_U246 = ~new_P3_R1209_U80 | ~new_P3_R1209_U98;
  assign new_P3_R1209_U247 = ~new_P3_U3433 | ~new_P3_R1209_U39;
  assign new_P3_R1209_U248 = ~P3_REG1_REG_15_ | ~new_P3_R1209_U40;
  assign new_P3_R1209_U249 = ~new_P3_R1209_U81;
  assign new_P3_R1209_U250 = ~new_P3_R1209_U249 | ~new_P3_R1209_U160;
  assign new_P3_R1209_U251 = ~new_P3_R1209_U81 | ~new_P3_R1209_U38;
  assign new_P3_R1209_U252 = ~P3_REG1_REG_14_ | ~new_P3_R1209_U37;
  assign new_P3_R1209_U253 = ~new_P3_U3430 | ~new_P3_R1209_U36;
  assign new_P3_R1209_U254 = ~new_P3_R1209_U82;
  assign new_P3_R1209_U255 = ~new_P3_R1209_U156 | ~new_P3_R1209_U254;
  assign new_P3_R1209_U256 = ~new_P3_R1209_U82 | ~new_P3_R1209_U99;
  assign new_P3_R1209_U257 = ~P3_REG1_REG_13_ | ~new_P3_R1209_U35;
  assign new_P3_R1209_U258 = ~new_P3_U3427 | ~new_P3_R1209_U34;
  assign new_P3_R1209_U259 = ~new_P3_R1209_U83;
  assign new_P3_R1209_U260 = ~new_P3_R1209_U152 | ~new_P3_R1209_U259;
  assign new_P3_R1209_U261 = ~new_P3_R1209_U83 | ~new_P3_R1209_U100;
  assign new_P3_R1209_U262 = ~P3_REG1_REG_12_ | ~new_P3_R1209_U33;
  assign new_P3_R1209_U263 = ~new_P3_U3424 | ~new_P3_R1209_U32;
  assign new_P3_R1209_U264 = ~new_P3_R1209_U84;
  assign new_P3_R1209_U265 = ~new_P3_R1209_U148 | ~new_P3_R1209_U264;
  assign new_P3_R1209_U266 = ~new_P3_R1209_U84 | ~new_P3_R1209_U101;
  assign new_P3_R1209_U267 = ~P3_REG1_REG_11_ | ~new_P3_R1209_U31;
  assign new_P3_R1209_U268 = ~new_P3_U3421 | ~new_P3_R1209_U30;
  assign new_P3_R1209_U269 = ~new_P3_R1209_U85;
  assign new_P3_R1209_U270 = ~new_P3_R1209_U144 | ~new_P3_R1209_U269;
  assign new_P3_R1209_U271 = ~new_P3_R1209_U85 | ~new_P3_R1209_U102;
  assign new_P3_R1209_U272 = ~P3_REG1_REG_10_ | ~new_P3_R1209_U29;
  assign new_P3_R1209_U273 = ~new_P3_U3418 | ~new_P3_R1209_U28;
  assign new_P3_R1209_U274 = ~new_P3_R1209_U86;
  assign new_P3_R1209_U275 = ~new_P3_R1209_U140 | ~new_P3_R1209_U274;
  assign new_P3_R1209_U276 = ~new_P3_R1209_U86 | ~new_P3_R1209_U103;
  assign new_P3_R1300_U6 = ~new_P3_U3058;
  assign new_P3_R1300_U7 = ~new_P3_U3055;
  assign new_P3_R1300_U8 = new_P3_R1300_U10 & new_P3_R1300_U9;
  assign new_P3_R1300_U9 = ~new_P3_U3055 | ~new_P3_R1300_U6;
  assign new_P3_R1300_U10 = ~new_P3_U3058 | ~new_P3_R1300_U7;
  assign new_P3_R1200_U6 = new_P3_R1200_U210 & new_P3_R1200_U209;
  assign new_P3_R1200_U7 = new_P3_R1200_U189 & new_P3_R1200_U245;
  assign new_P3_R1200_U8 = new_P3_R1200_U247 & new_P3_R1200_U246;
  assign new_P3_R1200_U9 = new_P3_R1200_U190 & new_P3_R1200_U262;
  assign new_P3_R1200_U10 = new_P3_R1200_U264 & new_P3_R1200_U263;
  assign new_P3_R1200_U11 = new_P3_R1200_U191 & new_P3_R1200_U286;
  assign new_P3_R1200_U12 = new_P3_R1200_U288 & new_P3_R1200_U287;
  assign new_P3_R1200_U13 = new_P3_R1200_U213 & new_P3_R1200_U208 & new_P3_R1200_U194;
  assign new_P3_R1200_U14 = new_P3_R1200_U218 & new_P3_R1200_U195;
  assign new_P3_R1200_U15 = new_P3_R1200_U392 & new_P3_R1200_U391;
  assign new_P3_R1200_U16 = ~new_P3_R1200_U342 | ~new_P3_R1200_U345;
  assign new_P3_R1200_U17 = ~new_P3_R1200_U331 | ~new_P3_R1200_U334;
  assign new_P3_R1200_U18 = ~new_P3_R1200_U320 | ~new_P3_R1200_U323;
  assign new_P3_R1200_U19 = ~new_P3_R1200_U312 | ~new_P3_R1200_U314;
  assign new_P3_R1200_U20 = ~new_P3_R1200_U351 | ~new_P3_R1200_U162 | ~new_P3_R1200_U183;
  assign new_P3_R1200_U21 = ~new_P3_R1200_U241 | ~new_P3_R1200_U243;
  assign new_P3_R1200_U22 = ~new_P3_R1200_U233 | ~new_P3_R1200_U236;
  assign new_P3_R1200_U23 = ~new_P3_R1200_U225 | ~new_P3_R1200_U227;
  assign new_P3_R1200_U24 = ~new_P3_R1200_U172 | ~new_P3_R1200_U348;
  assign new_P3_R1200_U25 = ~new_P3_U3069;
  assign new_P3_R1200_U26 = ~new_P3_U3069 | ~new_P3_R1200_U39;
  assign new_P3_R1200_U27 = ~new_P3_U3083;
  assign new_P3_R1200_U28 = ~new_P3_U3413;
  assign new_P3_R1200_U29 = ~new_P3_U3395;
  assign new_P3_R1200_U30 = ~new_P3_U3387;
  assign new_P3_R1200_U31 = ~new_P3_U3077;
  assign new_P3_R1200_U32 = ~new_P3_U3398;
  assign new_P3_R1200_U33 = ~new_P3_U3067;
  assign new_P3_R1200_U34 = ~new_P3_U3067 | ~new_P3_R1200_U29;
  assign new_P3_R1200_U35 = ~new_P3_U3063;
  assign new_P3_R1200_U36 = ~new_P3_U3404;
  assign new_P3_R1200_U37 = ~new_P3_U3407;
  assign new_P3_R1200_U38 = ~new_P3_U3401;
  assign new_P3_R1200_U39 = ~new_P3_U3410;
  assign new_P3_R1200_U40 = ~new_P3_U3070;
  assign new_P3_R1200_U41 = ~new_P3_U3066;
  assign new_P3_R1200_U42 = ~new_P3_U3059;
  assign new_P3_R1200_U43 = ~new_P3_U3059 | ~new_P3_R1200_U38;
  assign new_P3_R1200_U44 = ~new_P3_R1200_U214 | ~new_P3_R1200_U212;
  assign new_P3_R1200_U45 = ~new_P3_U3416;
  assign new_P3_R1200_U46 = ~new_P3_U3082;
  assign new_P3_R1200_U47 = ~new_P3_R1200_U44 | ~new_P3_R1200_U215;
  assign new_P3_R1200_U48 = ~new_P3_R1200_U43 | ~new_P3_R1200_U229;
  assign new_P3_R1200_U49 = ~new_P3_R1200_U349 | ~new_P3_R1200_U201 | ~new_P3_R1200_U185;
  assign new_P3_R1200_U50 = ~new_P3_U3901;
  assign new_P3_R1200_U51 = ~new_P3_U3422;
  assign new_P3_R1200_U52 = ~new_P3_U3419;
  assign new_P3_R1200_U53 = ~new_P3_U3062;
  assign new_P3_R1200_U54 = ~new_P3_U3061;
  assign new_P3_R1200_U55 = ~new_P3_U3082 | ~new_P3_R1200_U45;
  assign new_P3_R1200_U56 = ~new_P3_U3425;
  assign new_P3_R1200_U57 = ~new_P3_U3071;
  assign new_P3_R1200_U58 = ~new_P3_U3428;
  assign new_P3_R1200_U59 = ~new_P3_U3079;
  assign new_P3_R1200_U60 = ~new_P3_U3437;
  assign new_P3_R1200_U61 = ~new_P3_U3434;
  assign new_P3_R1200_U62 = ~new_P3_U3431;
  assign new_P3_R1200_U63 = ~new_P3_U3072;
  assign new_P3_R1200_U64 = ~new_P3_U3073;
  assign new_P3_R1200_U65 = ~new_P3_U3078;
  assign new_P3_R1200_U66 = ~new_P3_U3078 | ~new_P3_R1200_U62;
  assign new_P3_R1200_U67 = ~new_P3_U3440;
  assign new_P3_R1200_U68 = ~new_P3_U3068;
  assign new_P3_R1200_U69 = ~new_P3_U3081;
  assign new_P3_R1200_U70 = ~new_P3_U3445;
  assign new_P3_R1200_U71 = ~new_P3_U3080;
  assign new_P3_R1200_U72 = ~new_P3_U3907;
  assign new_P3_R1200_U73 = ~new_P3_U3075;
  assign new_P3_R1200_U74 = ~new_P3_U3904;
  assign new_P3_R1200_U75 = ~new_P3_U3905;
  assign new_P3_R1200_U76 = ~new_P3_U3906;
  assign new_P3_R1200_U77 = ~new_P3_U3065;
  assign new_P3_R1200_U78 = ~new_P3_U3060;
  assign new_P3_R1200_U79 = ~new_P3_U3074;
  assign new_P3_R1200_U80 = ~new_P3_U3074 | ~new_P3_R1200_U76;
  assign new_P3_R1200_U81 = ~new_P3_U3903;
  assign new_P3_R1200_U82 = ~new_P3_U3064;
  assign new_P3_R1200_U83 = ~new_P3_U3902;
  assign new_P3_R1200_U84 = ~new_P3_U3057;
  assign new_P3_R1200_U85 = ~new_P3_U3900;
  assign new_P3_R1200_U86 = ~new_P3_U3056;
  assign new_P3_R1200_U87 = ~new_P3_U3056 | ~new_P3_R1200_U50;
  assign new_P3_R1200_U88 = ~new_P3_U3052;
  assign new_P3_R1200_U89 = ~new_P3_U3899;
  assign new_P3_R1200_U90 = ~new_P3_U3053;
  assign new_P3_R1200_U91 = ~new_P3_R1200_U302 | ~new_P3_R1200_U301;
  assign new_P3_R1200_U92 = ~new_P3_R1200_U80 | ~new_P3_R1200_U316;
  assign new_P3_R1200_U93 = ~new_P3_R1200_U66 | ~new_P3_R1200_U327;
  assign new_P3_R1200_U94 = ~new_P3_R1200_U55 | ~new_P3_R1200_U338;
  assign new_P3_R1200_U95 = ~new_P3_U3076;
  assign new_P3_R1200_U96 = ~new_P3_R1200_U402 | ~new_P3_R1200_U401;
  assign new_P3_R1200_U97 = ~new_P3_R1200_U416 | ~new_P3_R1200_U415;
  assign new_P3_R1200_U98 = ~new_P3_R1200_U421 | ~new_P3_R1200_U420;
  assign new_P3_R1200_U99 = ~new_P3_R1200_U437 | ~new_P3_R1200_U436;
  assign new_P3_R1200_U100 = ~new_P3_R1200_U442 | ~new_P3_R1200_U441;
  assign new_P3_R1200_U101 = ~new_P3_R1200_U447 | ~new_P3_R1200_U446;
  assign new_P3_R1200_U102 = ~new_P3_R1200_U452 | ~new_P3_R1200_U451;
  assign new_P3_R1200_U103 = ~new_P3_R1200_U457 | ~new_P3_R1200_U456;
  assign new_P3_R1200_U104 = ~new_P3_R1200_U473 | ~new_P3_R1200_U472;
  assign new_P3_R1200_U105 = ~new_P3_R1200_U478 | ~new_P3_R1200_U477;
  assign new_P3_R1200_U106 = ~new_P3_R1200_U361 | ~new_P3_R1200_U360;
  assign new_P3_R1200_U107 = ~new_P3_R1200_U370 | ~new_P3_R1200_U369;
  assign new_P3_R1200_U108 = ~new_P3_R1200_U377 | ~new_P3_R1200_U376;
  assign new_P3_R1200_U109 = ~new_P3_R1200_U381 | ~new_P3_R1200_U380;
  assign new_P3_R1200_U110 = ~new_P3_R1200_U390 | ~new_P3_R1200_U389;
  assign new_P3_R1200_U111 = ~new_P3_R1200_U411 | ~new_P3_R1200_U410;
  assign new_P3_R1200_U112 = ~new_P3_R1200_U428 | ~new_P3_R1200_U427;
  assign new_P3_R1200_U113 = ~new_P3_R1200_U432 | ~new_P3_R1200_U431;
  assign new_P3_R1200_U114 = ~new_P3_R1200_U464 | ~new_P3_R1200_U463;
  assign new_P3_R1200_U115 = ~new_P3_R1200_U468 | ~new_P3_R1200_U467;
  assign new_P3_R1200_U116 = ~new_P3_R1200_U485 | ~new_P3_R1200_U484;
  assign new_P3_R1200_U117 = new_P3_R1200_U352 & new_P3_R1200_U193;
  assign new_P3_R1200_U118 = new_P3_R1200_U205 & new_P3_R1200_U206;
  assign new_P3_R1200_U119 = new_P3_R1200_U14 & new_P3_R1200_U13;
  assign new_P3_R1200_U120 = new_P3_R1200_U357 & new_P3_R1200_U354;
  assign new_P3_R1200_U121 = new_P3_R1200_U26 & new_P3_R1200_U363 & new_P3_R1200_U362;
  assign new_P3_R1200_U122 = new_P3_R1200_U366 & new_P3_R1200_U195;
  assign new_P3_R1200_U123 = new_P3_R1200_U235 & new_P3_R1200_U6;
  assign new_P3_R1200_U124 = new_P3_R1200_U373 & new_P3_R1200_U194;
  assign new_P3_R1200_U125 = new_P3_R1200_U34 & new_P3_R1200_U383 & new_P3_R1200_U382;
  assign new_P3_R1200_U126 = new_P3_R1200_U386 & new_P3_R1200_U193;
  assign new_P3_R1200_U127 = new_P3_R1200_U222 & new_P3_R1200_U7;
  assign new_P3_R1200_U128 = new_P3_R1200_U267 & new_P3_R1200_U9;
  assign new_P3_R1200_U129 = new_P3_R1200_U291 & new_P3_R1200_U11;
  assign new_P3_R1200_U130 = new_P3_R1200_U355 & new_P3_R1200_U192;
  assign new_P3_R1200_U131 = new_P3_R1200_U306 & new_P3_R1200_U307;
  assign new_P3_R1200_U132 = new_P3_R1200_U309 & new_P3_R1200_U395;
  assign new_P3_R1200_U133 = new_P3_R1200_U306 & new_P3_R1200_U307;
  assign new_P3_R1200_U134 = new_P3_R1200_U15 & new_P3_R1200_U310;
  assign new_P3_R1200_U135 = ~new_P3_R1200_U399 | ~new_P3_R1200_U398;
  assign new_P3_R1200_U136 = new_P3_R1200_U87 & new_P3_R1200_U404 & new_P3_R1200_U403;
  assign new_P3_R1200_U137 = new_P3_R1200_U407 & new_P3_R1200_U192;
  assign new_P3_R1200_U138 = ~new_P3_R1200_U413 | ~new_P3_R1200_U412;
  assign new_P3_R1200_U139 = ~new_P3_R1200_U418 | ~new_P3_R1200_U417;
  assign new_P3_R1200_U140 = new_P3_R1200_U322 & new_P3_R1200_U12;
  assign new_P3_R1200_U141 = new_P3_R1200_U424 & new_P3_R1200_U191;
  assign new_P3_R1200_U142 = ~new_P3_R1200_U434 | ~new_P3_R1200_U433;
  assign new_P3_R1200_U143 = ~new_P3_R1200_U439 | ~new_P3_R1200_U438;
  assign new_P3_R1200_U144 = ~new_P3_R1200_U444 | ~new_P3_R1200_U443;
  assign new_P3_R1200_U145 = ~new_P3_R1200_U449 | ~new_P3_R1200_U448;
  assign new_P3_R1200_U146 = ~new_P3_R1200_U454 | ~new_P3_R1200_U453;
  assign new_P3_R1200_U147 = new_P3_R1200_U333 & new_P3_R1200_U10;
  assign new_P3_R1200_U148 = new_P3_R1200_U460 & new_P3_R1200_U190;
  assign new_P3_R1200_U149 = ~new_P3_R1200_U470 | ~new_P3_R1200_U469;
  assign new_P3_R1200_U150 = ~new_P3_R1200_U475 | ~new_P3_R1200_U474;
  assign new_P3_R1200_U151 = new_P3_R1200_U344 & new_P3_R1200_U8;
  assign new_P3_R1200_U152 = new_P3_R1200_U481 & new_P3_R1200_U189;
  assign new_P3_R1200_U153 = new_P3_R1200_U359 & new_P3_R1200_U358;
  assign new_P3_R1200_U154 = ~new_P3_R1200_U120 | ~new_P3_R1200_U356;
  assign new_P3_R1200_U155 = new_P3_R1200_U368 & new_P3_R1200_U367;
  assign new_P3_R1200_U156 = new_P3_R1200_U375 & new_P3_R1200_U374;
  assign new_P3_R1200_U157 = new_P3_R1200_U379 & new_P3_R1200_U378;
  assign new_P3_R1200_U158 = ~new_P3_R1200_U118 | ~new_P3_R1200_U203;
  assign new_P3_R1200_U159 = new_P3_R1200_U388 & new_P3_R1200_U387;
  assign new_P3_R1200_U160 = ~new_P3_U3908;
  assign new_P3_R1200_U161 = ~new_P3_U3054;
  assign new_P3_R1200_U162 = new_P3_R1200_U397 & new_P3_R1200_U396;
  assign new_P3_R1200_U163 = ~new_P3_R1200_U131 | ~new_P3_R1200_U304;
  assign new_P3_R1200_U164 = new_P3_R1200_U409 & new_P3_R1200_U408;
  assign new_P3_R1200_U165 = ~new_P3_R1200_U298 | ~new_P3_R1200_U297;
  assign new_P3_R1200_U166 = ~new_P3_R1200_U294 | ~new_P3_R1200_U293;
  assign new_P3_R1200_U167 = new_P3_R1200_U426 & new_P3_R1200_U425;
  assign new_P3_R1200_U168 = new_P3_R1200_U430 & new_P3_R1200_U429;
  assign new_P3_R1200_U169 = ~new_P3_R1200_U284 | ~new_P3_R1200_U283;
  assign new_P3_R1200_U170 = ~new_P3_R1200_U280 | ~new_P3_R1200_U279;
  assign new_P3_R1200_U171 = ~new_P3_U3392;
  assign new_P3_R1200_U172 = ~new_P3_U3387 | ~new_P3_R1200_U95;
  assign new_P3_R1200_U173 = ~new_P3_R1200_U350 | ~new_P3_R1200_U276 | ~new_P3_R1200_U184;
  assign new_P3_R1200_U174 = ~new_P3_U3443;
  assign new_P3_R1200_U175 = ~new_P3_R1200_U274 | ~new_P3_R1200_U273;
  assign new_P3_R1200_U176 = ~new_P3_R1200_U270 | ~new_P3_R1200_U269;
  assign new_P3_R1200_U177 = new_P3_R1200_U462 & new_P3_R1200_U461;
  assign new_P3_R1200_U178 = new_P3_R1200_U466 & new_P3_R1200_U465;
  assign new_P3_R1200_U179 = ~new_P3_R1200_U260 | ~new_P3_R1200_U259;
  assign new_P3_R1200_U180 = ~new_P3_R1200_U256 | ~new_P3_R1200_U255;
  assign new_P3_R1200_U181 = ~new_P3_R1200_U252 | ~new_P3_R1200_U251;
  assign new_P3_R1200_U182 = new_P3_R1200_U483 & new_P3_R1200_U482;
  assign new_P3_R1200_U183 = ~new_P3_R1200_U132 | ~new_P3_R1200_U163;
  assign new_P3_R1200_U184 = ~new_P3_R1200_U175 | ~new_P3_R1200_U174;
  assign new_P3_R1200_U185 = ~new_P3_R1200_U172 | ~new_P3_R1200_U171;
  assign new_P3_R1200_U186 = ~new_P3_R1200_U87;
  assign new_P3_R1200_U187 = ~new_P3_R1200_U34;
  assign new_P3_R1200_U188 = ~new_P3_R1200_U26;
  assign new_P3_R1200_U189 = ~new_P3_U3419 | ~new_P3_R1200_U54;
  assign new_P3_R1200_U190 = ~new_P3_U3434 | ~new_P3_R1200_U64;
  assign new_P3_R1200_U191 = ~new_P3_U3905 | ~new_P3_R1200_U78;
  assign new_P3_R1200_U192 = ~new_P3_U3901 | ~new_P3_R1200_U86;
  assign new_P3_R1200_U193 = ~new_P3_U3395 | ~new_P3_R1200_U33;
  assign new_P3_R1200_U194 = ~new_P3_U3404 | ~new_P3_R1200_U41;
  assign new_P3_R1200_U195 = ~new_P3_U3410 | ~new_P3_R1200_U25;
  assign new_P3_R1200_U196 = ~new_P3_R1200_U66;
  assign new_P3_R1200_U197 = ~new_P3_R1200_U80;
  assign new_P3_R1200_U198 = ~new_P3_R1200_U43;
  assign new_P3_R1200_U199 = ~new_P3_R1200_U55;
  assign new_P3_R1200_U200 = ~new_P3_R1200_U172;
  assign new_P3_R1200_U201 = ~new_P3_U3077 | ~new_P3_R1200_U172;
  assign new_P3_R1200_U202 = ~new_P3_R1200_U49;
  assign new_P3_R1200_U203 = ~new_P3_R1200_U117 | ~new_P3_R1200_U49;
  assign new_P3_R1200_U204 = ~new_P3_R1200_U35 | ~new_P3_R1200_U34;
  assign new_P3_R1200_U205 = ~new_P3_R1200_U204 | ~new_P3_R1200_U32;
  assign new_P3_R1200_U206 = ~new_P3_U3063 | ~new_P3_R1200_U187;
  assign new_P3_R1200_U207 = ~new_P3_R1200_U158;
  assign new_P3_R1200_U208 = ~new_P3_U3407 | ~new_P3_R1200_U40;
  assign new_P3_R1200_U209 = ~new_P3_U3070 | ~new_P3_R1200_U37;
  assign new_P3_R1200_U210 = ~new_P3_U3066 | ~new_P3_R1200_U36;
  assign new_P3_R1200_U211 = ~new_P3_R1200_U198 | ~new_P3_R1200_U194;
  assign new_P3_R1200_U212 = ~new_P3_R1200_U6 | ~new_P3_R1200_U211;
  assign new_P3_R1200_U213 = ~new_P3_U3401 | ~new_P3_R1200_U42;
  assign new_P3_R1200_U214 = ~new_P3_U3407 | ~new_P3_R1200_U40;
  assign new_P3_R1200_U215 = ~new_P3_R1200_U13 | ~new_P3_R1200_U158;
  assign new_P3_R1200_U216 = ~new_P3_R1200_U44;
  assign new_P3_R1200_U217 = ~new_P3_R1200_U47;
  assign new_P3_R1200_U218 = ~new_P3_U3413 | ~new_P3_R1200_U27;
  assign new_P3_R1200_U219 = ~new_P3_R1200_U27 | ~new_P3_R1200_U26;
  assign new_P3_R1200_U220 = ~new_P3_U3083 | ~new_P3_R1200_U188;
  assign new_P3_R1200_U221 = ~new_P3_R1200_U154;
  assign new_P3_R1200_U222 = ~new_P3_U3416 | ~new_P3_R1200_U46;
  assign new_P3_R1200_U223 = ~new_P3_R1200_U222 | ~new_P3_R1200_U55;
  assign new_P3_R1200_U224 = ~new_P3_R1200_U217 | ~new_P3_R1200_U26;
  assign new_P3_R1200_U225 = ~new_P3_R1200_U122 | ~new_P3_R1200_U224;
  assign new_P3_R1200_U226 = ~new_P3_R1200_U47 | ~new_P3_R1200_U195;
  assign new_P3_R1200_U227 = ~new_P3_R1200_U121 | ~new_P3_R1200_U226;
  assign new_P3_R1200_U228 = ~new_P3_R1200_U26 | ~new_P3_R1200_U195;
  assign new_P3_R1200_U229 = ~new_P3_R1200_U213 | ~new_P3_R1200_U158;
  assign new_P3_R1200_U230 = ~new_P3_R1200_U48;
  assign new_P3_R1200_U231 = ~new_P3_U3066 | ~new_P3_R1200_U36;
  assign new_P3_R1200_U232 = ~new_P3_R1200_U230 | ~new_P3_R1200_U231;
  assign new_P3_R1200_U233 = ~new_P3_R1200_U124 | ~new_P3_R1200_U232;
  assign new_P3_R1200_U234 = ~new_P3_R1200_U48 | ~new_P3_R1200_U194;
  assign new_P3_R1200_U235 = ~new_P3_U3407 | ~new_P3_R1200_U40;
  assign new_P3_R1200_U236 = ~new_P3_R1200_U123 | ~new_P3_R1200_U234;
  assign new_P3_R1200_U237 = ~new_P3_U3066 | ~new_P3_R1200_U36;
  assign new_P3_R1200_U238 = ~new_P3_R1200_U194 | ~new_P3_R1200_U237;
  assign new_P3_R1200_U239 = ~new_P3_R1200_U213 | ~new_P3_R1200_U43;
  assign new_P3_R1200_U240 = ~new_P3_R1200_U202 | ~new_P3_R1200_U34;
  assign new_P3_R1200_U241 = ~new_P3_R1200_U126 | ~new_P3_R1200_U240;
  assign new_P3_R1200_U242 = ~new_P3_R1200_U49 | ~new_P3_R1200_U193;
  assign new_P3_R1200_U243 = ~new_P3_R1200_U125 | ~new_P3_R1200_U242;
  assign new_P3_R1200_U244 = ~new_P3_R1200_U193 | ~new_P3_R1200_U34;
  assign new_P3_R1200_U245 = ~new_P3_U3422 | ~new_P3_R1200_U53;
  assign new_P3_R1200_U246 = ~new_P3_U3062 | ~new_P3_R1200_U51;
  assign new_P3_R1200_U247 = ~new_P3_U3061 | ~new_P3_R1200_U52;
  assign new_P3_R1200_U248 = ~new_P3_R1200_U199 | ~new_P3_R1200_U7;
  assign new_P3_R1200_U249 = ~new_P3_R1200_U8 | ~new_P3_R1200_U248;
  assign new_P3_R1200_U250 = ~new_P3_U3422 | ~new_P3_R1200_U53;
  assign new_P3_R1200_U251 = ~new_P3_R1200_U127 | ~new_P3_R1200_U154;
  assign new_P3_R1200_U252 = ~new_P3_R1200_U250 | ~new_P3_R1200_U249;
  assign new_P3_R1200_U253 = ~new_P3_R1200_U181;
  assign new_P3_R1200_U254 = ~new_P3_U3425 | ~new_P3_R1200_U57;
  assign new_P3_R1200_U255 = ~new_P3_R1200_U254 | ~new_P3_R1200_U181;
  assign new_P3_R1200_U256 = ~new_P3_U3071 | ~new_P3_R1200_U56;
  assign new_P3_R1200_U257 = ~new_P3_R1200_U180;
  assign new_P3_R1200_U258 = ~new_P3_U3428 | ~new_P3_R1200_U59;
  assign new_P3_R1200_U259 = ~new_P3_R1200_U258 | ~new_P3_R1200_U180;
  assign new_P3_R1200_U260 = ~new_P3_U3079 | ~new_P3_R1200_U58;
  assign new_P3_R1200_U261 = ~new_P3_R1200_U179;
  assign new_P3_R1200_U262 = ~new_P3_U3437 | ~new_P3_R1200_U63;
  assign new_P3_R1200_U263 = ~new_P3_U3072 | ~new_P3_R1200_U60;
  assign new_P3_R1200_U264 = ~new_P3_U3073 | ~new_P3_R1200_U61;
  assign new_P3_R1200_U265 = ~new_P3_R1200_U196 | ~new_P3_R1200_U9;
  assign new_P3_R1200_U266 = ~new_P3_R1200_U10 | ~new_P3_R1200_U265;
  assign new_P3_R1200_U267 = ~new_P3_U3431 | ~new_P3_R1200_U65;
  assign new_P3_R1200_U268 = ~new_P3_U3437 | ~new_P3_R1200_U63;
  assign new_P3_R1200_U269 = ~new_P3_R1200_U128 | ~new_P3_R1200_U179;
  assign new_P3_R1200_U270 = ~new_P3_R1200_U268 | ~new_P3_R1200_U266;
  assign new_P3_R1200_U271 = ~new_P3_R1200_U176;
  assign new_P3_R1200_U272 = ~new_P3_U3440 | ~new_P3_R1200_U68;
  assign new_P3_R1200_U273 = ~new_P3_R1200_U272 | ~new_P3_R1200_U176;
  assign new_P3_R1200_U274 = ~new_P3_U3068 | ~new_P3_R1200_U67;
  assign new_P3_R1200_U275 = ~new_P3_R1200_U175;
  assign new_P3_R1200_U276 = ~new_P3_U3081 | ~new_P3_R1200_U175;
  assign new_P3_R1200_U277 = ~new_P3_R1200_U173;
  assign new_P3_R1200_U278 = ~new_P3_U3445 | ~new_P3_R1200_U71;
  assign new_P3_R1200_U279 = ~new_P3_R1200_U278 | ~new_P3_R1200_U173;
  assign new_P3_R1200_U280 = ~new_P3_U3080 | ~new_P3_R1200_U70;
  assign new_P3_R1200_U281 = ~new_P3_R1200_U170;
  assign new_P3_R1200_U282 = ~new_P3_U3907 | ~new_P3_R1200_U73;
  assign new_P3_R1200_U283 = ~new_P3_R1200_U282 | ~new_P3_R1200_U170;
  assign new_P3_R1200_U284 = ~new_P3_U3075 | ~new_P3_R1200_U72;
  assign new_P3_R1200_U285 = ~new_P3_R1200_U169;
  assign new_P3_R1200_U286 = ~new_P3_U3904 | ~new_P3_R1200_U77;
  assign new_P3_R1200_U287 = ~new_P3_U3065 | ~new_P3_R1200_U74;
  assign new_P3_R1200_U288 = ~new_P3_U3060 | ~new_P3_R1200_U75;
  assign new_P3_R1200_U289 = ~new_P3_R1200_U197 | ~new_P3_R1200_U11;
  assign new_P3_R1200_U290 = ~new_P3_R1200_U12 | ~new_P3_R1200_U289;
  assign new_P3_R1200_U291 = ~new_P3_U3906 | ~new_P3_R1200_U79;
  assign new_P3_R1200_U292 = ~new_P3_U3904 | ~new_P3_R1200_U77;
  assign new_P3_R1200_U293 = ~new_P3_R1200_U129 | ~new_P3_R1200_U169;
  assign new_P3_R1200_U294 = ~new_P3_R1200_U292 | ~new_P3_R1200_U290;
  assign new_P3_R1200_U295 = ~new_P3_R1200_U166;
  assign new_P3_R1200_U296 = ~new_P3_U3903 | ~new_P3_R1200_U82;
  assign new_P3_R1200_U297 = ~new_P3_R1200_U296 | ~new_P3_R1200_U166;
  assign new_P3_R1200_U298 = ~new_P3_U3064 | ~new_P3_R1200_U81;
  assign new_P3_R1200_U299 = ~new_P3_R1200_U165;
  assign new_P3_R1200_U300 = ~new_P3_U3902 | ~new_P3_R1200_U84;
  assign new_P3_R1200_U301 = ~new_P3_R1200_U300 | ~new_P3_R1200_U165;
  assign new_P3_R1200_U302 = ~new_P3_U3057 | ~new_P3_R1200_U83;
  assign new_P3_R1200_U303 = ~new_P3_R1200_U91;
  assign new_P3_R1200_U304 = ~new_P3_R1200_U130 | ~new_P3_R1200_U91;
  assign new_P3_R1200_U305 = ~new_P3_R1200_U88 | ~new_P3_R1200_U87;
  assign new_P3_R1200_U306 = ~new_P3_R1200_U305 | ~new_P3_R1200_U85;
  assign new_P3_R1200_U307 = ~new_P3_U3052 | ~new_P3_R1200_U186;
  assign new_P3_R1200_U308 = ~new_P3_R1200_U163;
  assign new_P3_R1200_U309 = ~new_P3_U3899 | ~new_P3_R1200_U90;
  assign new_P3_R1200_U310 = ~new_P3_U3053 | ~new_P3_R1200_U89;
  assign new_P3_R1200_U311 = ~new_P3_R1200_U303 | ~new_P3_R1200_U87;
  assign new_P3_R1200_U312 = ~new_P3_R1200_U137 | ~new_P3_R1200_U311;
  assign new_P3_R1200_U313 = ~new_P3_R1200_U91 | ~new_P3_R1200_U192;
  assign new_P3_R1200_U314 = ~new_P3_R1200_U136 | ~new_P3_R1200_U313;
  assign new_P3_R1200_U315 = ~new_P3_R1200_U192 | ~new_P3_R1200_U87;
  assign new_P3_R1200_U316 = ~new_P3_R1200_U291 | ~new_P3_R1200_U169;
  assign new_P3_R1200_U317 = ~new_P3_R1200_U92;
  assign new_P3_R1200_U318 = ~new_P3_U3060 | ~new_P3_R1200_U75;
  assign new_P3_R1200_U319 = ~new_P3_R1200_U317 | ~new_P3_R1200_U318;
  assign new_P3_R1200_U320 = ~new_P3_R1200_U141 | ~new_P3_R1200_U319;
  assign new_P3_R1200_U321 = ~new_P3_R1200_U92 | ~new_P3_R1200_U191;
  assign new_P3_R1200_U322 = ~new_P3_U3904 | ~new_P3_R1200_U77;
  assign new_P3_R1200_U323 = ~new_P3_R1200_U140 | ~new_P3_R1200_U321;
  assign new_P3_R1200_U324 = ~new_P3_U3060 | ~new_P3_R1200_U75;
  assign new_P3_R1200_U325 = ~new_P3_R1200_U191 | ~new_P3_R1200_U324;
  assign new_P3_R1200_U326 = ~new_P3_R1200_U291 | ~new_P3_R1200_U80;
  assign new_P3_R1200_U327 = ~new_P3_R1200_U267 | ~new_P3_R1200_U179;
  assign new_P3_R1200_U328 = ~new_P3_R1200_U93;
  assign new_P3_R1200_U329 = ~new_P3_U3073 | ~new_P3_R1200_U61;
  assign new_P3_R1200_U330 = ~new_P3_R1200_U328 | ~new_P3_R1200_U329;
  assign new_P3_R1200_U331 = ~new_P3_R1200_U148 | ~new_P3_R1200_U330;
  assign new_P3_R1200_U332 = ~new_P3_R1200_U93 | ~new_P3_R1200_U190;
  assign new_P3_R1200_U333 = ~new_P3_U3437 | ~new_P3_R1200_U63;
  assign new_P3_R1200_U334 = ~new_P3_R1200_U147 | ~new_P3_R1200_U332;
  assign new_P3_R1200_U335 = ~new_P3_U3073 | ~new_P3_R1200_U61;
  assign new_P3_R1200_U336 = ~new_P3_R1200_U190 | ~new_P3_R1200_U335;
  assign new_P3_R1200_U337 = ~new_P3_R1200_U267 | ~new_P3_R1200_U66;
  assign new_P3_R1200_U338 = ~new_P3_R1200_U222 | ~new_P3_R1200_U154;
  assign new_P3_R1200_U339 = ~new_P3_R1200_U94;
  assign new_P3_R1200_U340 = ~new_P3_U3061 | ~new_P3_R1200_U52;
  assign new_P3_R1200_U341 = ~new_P3_R1200_U339 | ~new_P3_R1200_U340;
  assign new_P3_R1200_U342 = ~new_P3_R1200_U152 | ~new_P3_R1200_U341;
  assign new_P3_R1200_U343 = ~new_P3_R1200_U94 | ~new_P3_R1200_U189;
  assign new_P3_R1200_U344 = ~new_P3_U3422 | ~new_P3_R1200_U53;
  assign new_P3_R1200_U345 = ~new_P3_R1200_U151 | ~new_P3_R1200_U343;
  assign new_P3_R1200_U346 = ~new_P3_U3061 | ~new_P3_R1200_U52;
  assign new_P3_R1200_U347 = ~new_P3_R1200_U189 | ~new_P3_R1200_U346;
  assign new_P3_R1200_U348 = ~new_P3_U3076 | ~new_P3_R1200_U30;
  assign new_P3_R1200_U349 = ~new_P3_U3077 | ~new_P3_R1200_U171;
  assign new_P3_R1200_U350 = ~new_P3_U3081 | ~new_P3_R1200_U174;
  assign new_P3_R1200_U351 = ~new_P3_R1200_U134 | ~new_P3_R1200_U133 | ~new_P3_R1200_U304;
  assign new_P3_R1200_U352 = ~new_P3_U3398 | ~new_P3_R1200_U35;
  assign new_P3_R1200_U353 = ~new_P3_U3413 | ~new_P3_R1200_U220;
  assign new_P3_R1200_U354 = ~new_P3_R1200_U353 | ~new_P3_R1200_U219;
  assign new_P3_R1200_U355 = ~new_P3_U3900 | ~new_P3_R1200_U88;
  assign new_P3_R1200_U356 = ~new_P3_R1200_U119 | ~new_P3_R1200_U158;
  assign new_P3_R1200_U357 = ~new_P3_R1200_U216 | ~new_P3_R1200_U14;
  assign new_P3_R1200_U358 = ~new_P3_U3416 | ~new_P3_R1200_U46;
  assign new_P3_R1200_U359 = ~new_P3_U3082 | ~new_P3_R1200_U45;
  assign new_P3_R1200_U360 = ~new_P3_R1200_U223 | ~new_P3_R1200_U154;
  assign new_P3_R1200_U361 = ~new_P3_R1200_U221 | ~new_P3_R1200_U153;
  assign new_P3_R1200_U362 = ~new_P3_U3413 | ~new_P3_R1200_U27;
  assign new_P3_R1200_U363 = ~new_P3_U3083 | ~new_P3_R1200_U28;
  assign new_P3_R1200_U364 = ~new_P3_U3413 | ~new_P3_R1200_U27;
  assign new_P3_R1200_U365 = ~new_P3_U3083 | ~new_P3_R1200_U28;
  assign new_P3_R1200_U366 = ~new_P3_R1200_U365 | ~new_P3_R1200_U364;
  assign new_P3_R1200_U367 = ~new_P3_U3410 | ~new_P3_R1200_U25;
  assign new_P3_R1200_U368 = ~new_P3_U3069 | ~new_P3_R1200_U39;
  assign new_P3_R1200_U369 = ~new_P3_R1200_U228 | ~new_P3_R1200_U47;
  assign new_P3_R1200_U370 = ~new_P3_R1200_U155 | ~new_P3_R1200_U217;
  assign new_P3_R1200_U371 = ~new_P3_U3407 | ~new_P3_R1200_U40;
  assign new_P3_R1200_U372 = ~new_P3_U3070 | ~new_P3_R1200_U37;
  assign new_P3_R1200_U373 = ~new_P3_R1200_U372 | ~new_P3_R1200_U371;
  assign new_P3_R1200_U374 = ~new_P3_U3404 | ~new_P3_R1200_U41;
  assign new_P3_R1200_U375 = ~new_P3_U3066 | ~new_P3_R1200_U36;
  assign new_P3_R1200_U376 = ~new_P3_R1200_U238 | ~new_P3_R1200_U48;
  assign new_P3_R1200_U377 = ~new_P3_R1200_U156 | ~new_P3_R1200_U230;
  assign new_P3_R1200_U378 = ~new_P3_U3401 | ~new_P3_R1200_U42;
  assign new_P3_R1200_U379 = ~new_P3_U3059 | ~new_P3_R1200_U38;
  assign new_P3_R1200_U380 = ~new_P3_R1200_U239 | ~new_P3_R1200_U158;
  assign new_P3_R1200_U381 = ~new_P3_R1200_U207 | ~new_P3_R1200_U157;
  assign new_P3_R1200_U382 = ~new_P3_U3398 | ~new_P3_R1200_U35;
  assign new_P3_R1200_U383 = ~new_P3_U3063 | ~new_P3_R1200_U32;
  assign new_P3_R1200_U384 = ~new_P3_U3398 | ~new_P3_R1200_U35;
  assign new_P3_R1200_U385 = ~new_P3_U3063 | ~new_P3_R1200_U32;
  assign new_P3_R1200_U386 = ~new_P3_R1200_U385 | ~new_P3_R1200_U384;
  assign new_P3_R1200_U387 = ~new_P3_U3395 | ~new_P3_R1200_U33;
  assign new_P3_R1200_U388 = ~new_P3_U3067 | ~new_P3_R1200_U29;
  assign new_P3_R1200_U389 = ~new_P3_R1200_U244 | ~new_P3_R1200_U49;
  assign new_P3_R1200_U390 = ~new_P3_R1200_U159 | ~new_P3_R1200_U202;
  assign new_P3_R1200_U391 = ~new_P3_U3908 | ~new_P3_R1200_U161;
  assign new_P3_R1200_U392 = ~new_P3_U3054 | ~new_P3_R1200_U160;
  assign new_P3_R1200_U393 = ~new_P3_U3908 | ~new_P3_R1200_U161;
  assign new_P3_R1200_U394 = ~new_P3_U3054 | ~new_P3_R1200_U160;
  assign new_P3_R1200_U395 = ~new_P3_R1200_U394 | ~new_P3_R1200_U393;
  assign new_P3_R1200_U396 = ~new_P3_R1200_U89 | ~new_P3_U3053 | ~new_P3_R1200_U395;
  assign new_P3_R1200_U397 = ~new_P3_U3899 | ~new_P3_R1200_U15 | ~new_P3_R1200_U90;
  assign new_P3_R1200_U398 = ~new_P3_U3899 | ~new_P3_R1200_U90;
  assign new_P3_R1200_U399 = ~new_P3_U3053 | ~new_P3_R1200_U89;
  assign new_P3_R1200_U400 = ~new_P3_R1200_U135;
  assign new_P3_R1200_U401 = ~new_P3_R1200_U308 | ~new_P3_R1200_U400;
  assign new_P3_R1200_U402 = ~new_P3_R1200_U135 | ~new_P3_R1200_U163;
  assign new_P3_R1200_U403 = ~new_P3_U3900 | ~new_P3_R1200_U88;
  assign new_P3_R1200_U404 = ~new_P3_U3052 | ~new_P3_R1200_U85;
  assign new_P3_R1200_U405 = ~new_P3_U3900 | ~new_P3_R1200_U88;
  assign new_P3_R1200_U406 = ~new_P3_U3052 | ~new_P3_R1200_U85;
  assign new_P3_R1200_U407 = ~new_P3_R1200_U406 | ~new_P3_R1200_U405;
  assign new_P3_R1200_U408 = ~new_P3_U3901 | ~new_P3_R1200_U86;
  assign new_P3_R1200_U409 = ~new_P3_U3056 | ~new_P3_R1200_U50;
  assign new_P3_R1200_U410 = ~new_P3_R1200_U315 | ~new_P3_R1200_U91;
  assign new_P3_R1200_U411 = ~new_P3_R1200_U164 | ~new_P3_R1200_U303;
  assign new_P3_R1200_U412 = ~new_P3_U3902 | ~new_P3_R1200_U84;
  assign new_P3_R1200_U413 = ~new_P3_U3057 | ~new_P3_R1200_U83;
  assign new_P3_R1200_U414 = ~new_P3_R1200_U138;
  assign new_P3_R1200_U415 = ~new_P3_R1200_U299 | ~new_P3_R1200_U414;
  assign new_P3_R1200_U416 = ~new_P3_R1200_U138 | ~new_P3_R1200_U165;
  assign new_P3_R1200_U417 = ~new_P3_U3903 | ~new_P3_R1200_U82;
  assign new_P3_R1200_U418 = ~new_P3_U3064 | ~new_P3_R1200_U81;
  assign new_P3_R1200_U419 = ~new_P3_R1200_U139;
  assign new_P3_R1200_U420 = ~new_P3_R1200_U295 | ~new_P3_R1200_U419;
  assign new_P3_R1200_U421 = ~new_P3_R1200_U139 | ~new_P3_R1200_U166;
  assign new_P3_R1200_U422 = ~new_P3_U3904 | ~new_P3_R1200_U77;
  assign new_P3_R1200_U423 = ~new_P3_U3065 | ~new_P3_R1200_U74;
  assign new_P3_R1200_U424 = ~new_P3_R1200_U423 | ~new_P3_R1200_U422;
  assign new_P3_R1200_U425 = ~new_P3_U3905 | ~new_P3_R1200_U78;
  assign new_P3_R1200_U426 = ~new_P3_U3060 | ~new_P3_R1200_U75;
  assign new_P3_R1200_U427 = ~new_P3_R1200_U325 | ~new_P3_R1200_U92;
  assign new_P3_R1200_U428 = ~new_P3_R1200_U167 | ~new_P3_R1200_U317;
  assign new_P3_R1200_U429 = ~new_P3_U3906 | ~new_P3_R1200_U79;
  assign new_P3_R1200_U430 = ~new_P3_U3074 | ~new_P3_R1200_U76;
  assign new_P3_R1200_U431 = ~new_P3_R1200_U326 | ~new_P3_R1200_U169;
  assign new_P3_R1200_U432 = ~new_P3_R1200_U285 | ~new_P3_R1200_U168;
  assign new_P3_R1200_U433 = ~new_P3_U3907 | ~new_P3_R1200_U73;
  assign new_P3_R1200_U434 = ~new_P3_U3075 | ~new_P3_R1200_U72;
  assign new_P3_R1200_U435 = ~new_P3_R1200_U142;
  assign new_P3_R1200_U436 = ~new_P3_R1200_U281 | ~new_P3_R1200_U435;
  assign new_P3_R1200_U437 = ~new_P3_R1200_U142 | ~new_P3_R1200_U170;
  assign new_P3_R1200_U438 = ~new_P3_U3392 | ~new_P3_R1200_U31;
  assign new_P3_R1200_U439 = ~new_P3_U3077 | ~new_P3_R1200_U171;
  assign new_P3_R1200_U440 = ~new_P3_R1200_U143;
  assign new_P3_R1200_U441 = ~new_P3_R1200_U200 | ~new_P3_R1200_U440;
  assign new_P3_R1200_U442 = ~new_P3_R1200_U143 | ~new_P3_R1200_U172;
  assign new_P3_R1200_U443 = ~new_P3_U3445 | ~new_P3_R1200_U71;
  assign new_P3_R1200_U444 = ~new_P3_U3080 | ~new_P3_R1200_U70;
  assign new_P3_R1200_U445 = ~new_P3_R1200_U144;
  assign new_P3_R1200_U446 = ~new_P3_R1200_U277 | ~new_P3_R1200_U445;
  assign new_P3_R1200_U447 = ~new_P3_R1200_U144 | ~new_P3_R1200_U173;
  assign new_P3_R1200_U448 = ~new_P3_U3443 | ~new_P3_R1200_U69;
  assign new_P3_R1200_U449 = ~new_P3_U3081 | ~new_P3_R1200_U174;
  assign new_P3_R1200_U450 = ~new_P3_R1200_U145;
  assign new_P3_R1200_U451 = ~new_P3_R1200_U275 | ~new_P3_R1200_U450;
  assign new_P3_R1200_U452 = ~new_P3_R1200_U145 | ~new_P3_R1200_U175;
  assign new_P3_R1200_U453 = ~new_P3_U3440 | ~new_P3_R1200_U68;
  assign new_P3_R1200_U454 = ~new_P3_U3068 | ~new_P3_R1200_U67;
  assign new_P3_R1200_U455 = ~new_P3_R1200_U146;
  assign new_P3_R1200_U456 = ~new_P3_R1200_U271 | ~new_P3_R1200_U455;
  assign new_P3_R1200_U457 = ~new_P3_R1200_U146 | ~new_P3_R1200_U176;
  assign new_P3_R1200_U458 = ~new_P3_U3437 | ~new_P3_R1200_U63;
  assign new_P3_R1200_U459 = ~new_P3_U3072 | ~new_P3_R1200_U60;
  assign new_P3_R1200_U460 = ~new_P3_R1200_U459 | ~new_P3_R1200_U458;
  assign new_P3_R1200_U461 = ~new_P3_U3434 | ~new_P3_R1200_U64;
  assign new_P3_R1200_U462 = ~new_P3_U3073 | ~new_P3_R1200_U61;
  assign new_P3_R1200_U463 = ~new_P3_R1200_U336 | ~new_P3_R1200_U93;
  assign new_P3_R1200_U464 = ~new_P3_R1200_U177 | ~new_P3_R1200_U328;
  assign new_P3_R1200_U465 = ~new_P3_U3431 | ~new_P3_R1200_U65;
  assign new_P3_R1200_U466 = ~new_P3_U3078 | ~new_P3_R1200_U62;
  assign new_P3_R1200_U467 = ~new_P3_R1200_U337 | ~new_P3_R1200_U179;
  assign new_P3_R1200_U468 = ~new_P3_R1200_U261 | ~new_P3_R1200_U178;
  assign new_P3_R1200_U469 = ~new_P3_U3428 | ~new_P3_R1200_U59;
  assign new_P3_R1200_U470 = ~new_P3_U3079 | ~new_P3_R1200_U58;
  assign new_P3_R1200_U471 = ~new_P3_R1200_U149;
  assign new_P3_R1200_U472 = ~new_P3_R1200_U257 | ~new_P3_R1200_U471;
  assign new_P3_R1200_U473 = ~new_P3_R1200_U149 | ~new_P3_R1200_U180;
  assign new_P3_R1200_U474 = ~new_P3_U3425 | ~new_P3_R1200_U57;
  assign new_P3_R1200_U475 = ~new_P3_U3071 | ~new_P3_R1200_U56;
  assign new_P3_R1200_U476 = ~new_P3_R1200_U150;
  assign new_P3_R1200_U477 = ~new_P3_R1200_U253 | ~new_P3_R1200_U476;
  assign new_P3_R1200_U478 = ~new_P3_R1200_U150 | ~new_P3_R1200_U181;
  assign new_P3_R1200_U479 = ~new_P3_U3422 | ~new_P3_R1200_U53;
  assign new_P3_R1200_U480 = ~new_P3_U3062 | ~new_P3_R1200_U51;
  assign new_P3_R1200_U481 = ~new_P3_R1200_U480 | ~new_P3_R1200_U479;
  assign new_P3_R1200_U482 = ~new_P3_U3419 | ~new_P3_R1200_U54;
  assign new_P3_R1200_U483 = ~new_P3_U3061 | ~new_P3_R1200_U52;
  assign new_P3_R1200_U484 = ~new_P3_R1200_U347 | ~new_P3_R1200_U94;
  assign new_P3_R1200_U485 = ~new_P3_R1200_U182 | ~new_P3_R1200_U339;
  assign new_P3_R1179_U6 = new_P3_R1179_U210 & new_P3_R1179_U209;
  assign new_P3_R1179_U7 = new_P3_R1179_U189 & new_P3_R1179_U245;
  assign new_P3_R1179_U8 = new_P3_R1179_U247 & new_P3_R1179_U246;
  assign new_P3_R1179_U9 = new_P3_R1179_U190 & new_P3_R1179_U262;
  assign new_P3_R1179_U10 = new_P3_R1179_U264 & new_P3_R1179_U263;
  assign new_P3_R1179_U11 = new_P3_R1179_U191 & new_P3_R1179_U286;
  assign new_P3_R1179_U12 = new_P3_R1179_U288 & new_P3_R1179_U287;
  assign new_P3_R1179_U13 = new_P3_R1179_U213 & new_P3_R1179_U208 & new_P3_R1179_U194;
  assign new_P3_R1179_U14 = new_P3_R1179_U218 & new_P3_R1179_U195;
  assign new_P3_R1179_U15 = new_P3_R1179_U392 & new_P3_R1179_U391;
  assign new_P3_R1179_U16 = ~new_P3_R1179_U342 | ~new_P3_R1179_U345;
  assign new_P3_R1179_U17 = ~new_P3_R1179_U331 | ~new_P3_R1179_U334;
  assign new_P3_R1179_U18 = ~new_P3_R1179_U320 | ~new_P3_R1179_U323;
  assign new_P3_R1179_U19 = ~new_P3_R1179_U312 | ~new_P3_R1179_U314;
  assign new_P3_R1179_U20 = ~new_P3_R1179_U351 | ~new_P3_R1179_U162 | ~new_P3_R1179_U183;
  assign new_P3_R1179_U21 = ~new_P3_R1179_U241 | ~new_P3_R1179_U243;
  assign new_P3_R1179_U22 = ~new_P3_R1179_U233 | ~new_P3_R1179_U236;
  assign new_P3_R1179_U23 = ~new_P3_R1179_U225 | ~new_P3_R1179_U227;
  assign new_P3_R1179_U24 = ~new_P3_R1179_U172 | ~new_P3_R1179_U348;
  assign new_P3_R1179_U25 = ~new_P3_U3069;
  assign new_P3_R1179_U26 = ~new_P3_U3069 | ~new_P3_R1179_U39;
  assign new_P3_R1179_U27 = ~new_P3_U3083;
  assign new_P3_R1179_U28 = ~new_P3_U3413;
  assign new_P3_R1179_U29 = ~new_P3_U3395;
  assign new_P3_R1179_U30 = ~new_P3_U3387;
  assign new_P3_R1179_U31 = ~new_P3_U3077;
  assign new_P3_R1179_U32 = ~new_P3_U3398;
  assign new_P3_R1179_U33 = ~new_P3_U3067;
  assign new_P3_R1179_U34 = ~new_P3_U3067 | ~new_P3_R1179_U29;
  assign new_P3_R1179_U35 = ~new_P3_U3063;
  assign new_P3_R1179_U36 = ~new_P3_U3404;
  assign new_P3_R1179_U37 = ~new_P3_U3407;
  assign new_P3_R1179_U38 = ~new_P3_U3401;
  assign new_P3_R1179_U39 = ~new_P3_U3410;
  assign new_P3_R1179_U40 = ~new_P3_U3070;
  assign new_P3_R1179_U41 = ~new_P3_U3066;
  assign new_P3_R1179_U42 = ~new_P3_U3059;
  assign new_P3_R1179_U43 = ~new_P3_U3059 | ~new_P3_R1179_U38;
  assign new_P3_R1179_U44 = ~new_P3_R1179_U214 | ~new_P3_R1179_U212;
  assign new_P3_R1179_U45 = ~new_P3_U3416;
  assign new_P3_R1179_U46 = ~new_P3_U3082;
  assign new_P3_R1179_U47 = ~new_P3_R1179_U44 | ~new_P3_R1179_U215;
  assign new_P3_R1179_U48 = ~new_P3_R1179_U43 | ~new_P3_R1179_U229;
  assign new_P3_R1179_U49 = ~new_P3_R1179_U349 | ~new_P3_R1179_U201 | ~new_P3_R1179_U185;
  assign new_P3_R1179_U50 = ~new_P3_U3901;
  assign new_P3_R1179_U51 = ~new_P3_U3422;
  assign new_P3_R1179_U52 = ~new_P3_U3419;
  assign new_P3_R1179_U53 = ~new_P3_U3062;
  assign new_P3_R1179_U54 = ~new_P3_U3061;
  assign new_P3_R1179_U55 = ~new_P3_U3082 | ~new_P3_R1179_U45;
  assign new_P3_R1179_U56 = ~new_P3_U3425;
  assign new_P3_R1179_U57 = ~new_P3_U3071;
  assign new_P3_R1179_U58 = ~new_P3_U3428;
  assign new_P3_R1179_U59 = ~new_P3_U3079;
  assign new_P3_R1179_U60 = ~new_P3_U3437;
  assign new_P3_R1179_U61 = ~new_P3_U3434;
  assign new_P3_R1179_U62 = ~new_P3_U3431;
  assign new_P3_R1179_U63 = ~new_P3_U3072;
  assign new_P3_R1179_U64 = ~new_P3_U3073;
  assign new_P3_R1179_U65 = ~new_P3_U3078;
  assign new_P3_R1179_U66 = ~new_P3_U3078 | ~new_P3_R1179_U62;
  assign new_P3_R1179_U67 = ~new_P3_U3440;
  assign new_P3_R1179_U68 = ~new_P3_U3068;
  assign new_P3_R1179_U69 = ~new_P3_U3081;
  assign new_P3_R1179_U70 = ~new_P3_U3445;
  assign new_P3_R1179_U71 = ~new_P3_U3080;
  assign new_P3_R1179_U72 = ~new_P3_U3907;
  assign new_P3_R1179_U73 = ~new_P3_U3075;
  assign new_P3_R1179_U74 = ~new_P3_U3904;
  assign new_P3_R1179_U75 = ~new_P3_U3905;
  assign new_P3_R1179_U76 = ~new_P3_U3906;
  assign new_P3_R1179_U77 = ~new_P3_U3065;
  assign new_P3_R1179_U78 = ~new_P3_U3060;
  assign new_P3_R1179_U79 = ~new_P3_U3074;
  assign new_P3_R1179_U80 = ~new_P3_U3074 | ~new_P3_R1179_U76;
  assign new_P3_R1179_U81 = ~new_P3_U3903;
  assign new_P3_R1179_U82 = ~new_P3_U3064;
  assign new_P3_R1179_U83 = ~new_P3_U3902;
  assign new_P3_R1179_U84 = ~new_P3_U3057;
  assign new_P3_R1179_U85 = ~new_P3_U3900;
  assign new_P3_R1179_U86 = ~new_P3_U3056;
  assign new_P3_R1179_U87 = ~new_P3_U3056 | ~new_P3_R1179_U50;
  assign new_P3_R1179_U88 = ~new_P3_U3052;
  assign new_P3_R1179_U89 = ~new_P3_U3899;
  assign new_P3_R1179_U90 = ~new_P3_U3053;
  assign new_P3_R1179_U91 = ~new_P3_R1179_U302 | ~new_P3_R1179_U301;
  assign new_P3_R1179_U92 = ~new_P3_R1179_U80 | ~new_P3_R1179_U316;
  assign new_P3_R1179_U93 = ~new_P3_R1179_U66 | ~new_P3_R1179_U327;
  assign new_P3_R1179_U94 = ~new_P3_R1179_U55 | ~new_P3_R1179_U338;
  assign new_P3_R1179_U95 = ~new_P3_U3076;
  assign new_P3_R1179_U96 = ~new_P3_R1179_U402 | ~new_P3_R1179_U401;
  assign new_P3_R1179_U97 = ~new_P3_R1179_U416 | ~new_P3_R1179_U415;
  assign new_P3_R1179_U98 = ~new_P3_R1179_U421 | ~new_P3_R1179_U420;
  assign new_P3_R1179_U99 = ~new_P3_R1179_U437 | ~new_P3_R1179_U436;
  assign new_P3_R1179_U100 = ~new_P3_R1179_U442 | ~new_P3_R1179_U441;
  assign new_P3_R1179_U101 = ~new_P3_R1179_U447 | ~new_P3_R1179_U446;
  assign new_P3_R1179_U102 = ~new_P3_R1179_U452 | ~new_P3_R1179_U451;
  assign new_P3_R1179_U103 = ~new_P3_R1179_U457 | ~new_P3_R1179_U456;
  assign new_P3_R1179_U104 = ~new_P3_R1179_U473 | ~new_P3_R1179_U472;
  assign new_P3_R1179_U105 = ~new_P3_R1179_U478 | ~new_P3_R1179_U477;
  assign new_P3_R1179_U106 = ~new_P3_R1179_U361 | ~new_P3_R1179_U360;
  assign new_P3_R1179_U107 = ~new_P3_R1179_U370 | ~new_P3_R1179_U369;
  assign new_P3_R1179_U108 = ~new_P3_R1179_U377 | ~new_P3_R1179_U376;
  assign new_P3_R1179_U109 = ~new_P3_R1179_U381 | ~new_P3_R1179_U380;
  assign new_P3_R1179_U110 = ~new_P3_R1179_U390 | ~new_P3_R1179_U389;
  assign new_P3_R1179_U111 = ~new_P3_R1179_U411 | ~new_P3_R1179_U410;
  assign new_P3_R1179_U112 = ~new_P3_R1179_U428 | ~new_P3_R1179_U427;
  assign new_P3_R1179_U113 = ~new_P3_R1179_U432 | ~new_P3_R1179_U431;
  assign new_P3_R1179_U114 = ~new_P3_R1179_U464 | ~new_P3_R1179_U463;
  assign new_P3_R1179_U115 = ~new_P3_R1179_U468 | ~new_P3_R1179_U467;
  assign new_P3_R1179_U116 = ~new_P3_R1179_U485 | ~new_P3_R1179_U484;
  assign new_P3_R1179_U117 = new_P3_R1179_U352 & new_P3_R1179_U193;
  assign new_P3_R1179_U118 = new_P3_R1179_U205 & new_P3_R1179_U206;
  assign new_P3_R1179_U119 = new_P3_R1179_U14 & new_P3_R1179_U13;
  assign new_P3_R1179_U120 = new_P3_R1179_U357 & new_P3_R1179_U354;
  assign new_P3_R1179_U121 = new_P3_R1179_U26 & new_P3_R1179_U363 & new_P3_R1179_U362;
  assign new_P3_R1179_U122 = new_P3_R1179_U366 & new_P3_R1179_U195;
  assign new_P3_R1179_U123 = new_P3_R1179_U235 & new_P3_R1179_U6;
  assign new_P3_R1179_U124 = new_P3_R1179_U373 & new_P3_R1179_U194;
  assign new_P3_R1179_U125 = new_P3_R1179_U34 & new_P3_R1179_U383 & new_P3_R1179_U382;
  assign new_P3_R1179_U126 = new_P3_R1179_U386 & new_P3_R1179_U193;
  assign new_P3_R1179_U127 = new_P3_R1179_U222 & new_P3_R1179_U7;
  assign new_P3_R1179_U128 = new_P3_R1179_U267 & new_P3_R1179_U9;
  assign new_P3_R1179_U129 = new_P3_R1179_U291 & new_P3_R1179_U11;
  assign new_P3_R1179_U130 = new_P3_R1179_U355 & new_P3_R1179_U192;
  assign new_P3_R1179_U131 = new_P3_R1179_U306 & new_P3_R1179_U307;
  assign new_P3_R1179_U132 = new_P3_R1179_U309 & new_P3_R1179_U395;
  assign new_P3_R1179_U133 = new_P3_R1179_U306 & new_P3_R1179_U307;
  assign new_P3_R1179_U134 = new_P3_R1179_U15 & new_P3_R1179_U310;
  assign new_P3_R1179_U135 = ~new_P3_R1179_U399 | ~new_P3_R1179_U398;
  assign new_P3_R1179_U136 = new_P3_R1179_U87 & new_P3_R1179_U404 & new_P3_R1179_U403;
  assign new_P3_R1179_U137 = new_P3_R1179_U407 & new_P3_R1179_U192;
  assign new_P3_R1179_U138 = ~new_P3_R1179_U413 | ~new_P3_R1179_U412;
  assign new_P3_R1179_U139 = ~new_P3_R1179_U418 | ~new_P3_R1179_U417;
  assign new_P3_R1179_U140 = new_P3_R1179_U322 & new_P3_R1179_U12;
  assign new_P3_R1179_U141 = new_P3_R1179_U424 & new_P3_R1179_U191;
  assign new_P3_R1179_U142 = ~new_P3_R1179_U434 | ~new_P3_R1179_U433;
  assign new_P3_R1179_U143 = ~new_P3_R1179_U439 | ~new_P3_R1179_U438;
  assign new_P3_R1179_U144 = ~new_P3_R1179_U444 | ~new_P3_R1179_U443;
  assign new_P3_R1179_U145 = ~new_P3_R1179_U449 | ~new_P3_R1179_U448;
  assign new_P3_R1179_U146 = ~new_P3_R1179_U454 | ~new_P3_R1179_U453;
  assign new_P3_R1179_U147 = new_P3_R1179_U333 & new_P3_R1179_U10;
  assign new_P3_R1179_U148 = new_P3_R1179_U460 & new_P3_R1179_U190;
  assign new_P3_R1179_U149 = ~new_P3_R1179_U470 | ~new_P3_R1179_U469;
  assign new_P3_R1179_U150 = ~new_P3_R1179_U475 | ~new_P3_R1179_U474;
  assign new_P3_R1179_U151 = new_P3_R1179_U344 & new_P3_R1179_U8;
  assign new_P3_R1179_U152 = new_P3_R1179_U481 & new_P3_R1179_U189;
  assign new_P3_R1179_U153 = new_P3_R1179_U359 & new_P3_R1179_U358;
  assign new_P3_R1179_U154 = ~new_P3_R1179_U120 | ~new_P3_R1179_U356;
  assign new_P3_R1179_U155 = new_P3_R1179_U368 & new_P3_R1179_U367;
  assign new_P3_R1179_U156 = new_P3_R1179_U375 & new_P3_R1179_U374;
  assign new_P3_R1179_U157 = new_P3_R1179_U379 & new_P3_R1179_U378;
  assign new_P3_R1179_U158 = ~new_P3_R1179_U118 | ~new_P3_R1179_U203;
  assign new_P3_R1179_U159 = new_P3_R1179_U388 & new_P3_R1179_U387;
  assign new_P3_R1179_U160 = ~new_P3_U3908;
  assign new_P3_R1179_U161 = ~new_P3_U3054;
  assign new_P3_R1179_U162 = new_P3_R1179_U397 & new_P3_R1179_U396;
  assign new_P3_R1179_U163 = ~new_P3_R1179_U131 | ~new_P3_R1179_U304;
  assign new_P3_R1179_U164 = new_P3_R1179_U409 & new_P3_R1179_U408;
  assign new_P3_R1179_U165 = ~new_P3_R1179_U298 | ~new_P3_R1179_U297;
  assign new_P3_R1179_U166 = ~new_P3_R1179_U294 | ~new_P3_R1179_U293;
  assign new_P3_R1179_U167 = new_P3_R1179_U426 & new_P3_R1179_U425;
  assign new_P3_R1179_U168 = new_P3_R1179_U430 & new_P3_R1179_U429;
  assign new_P3_R1179_U169 = ~new_P3_R1179_U284 | ~new_P3_R1179_U283;
  assign new_P3_R1179_U170 = ~new_P3_R1179_U280 | ~new_P3_R1179_U279;
  assign new_P3_R1179_U171 = ~new_P3_U3392;
  assign new_P3_R1179_U172 = ~new_P3_U3387 | ~new_P3_R1179_U95;
  assign new_P3_R1179_U173 = ~new_P3_R1179_U350 | ~new_P3_R1179_U276 | ~new_P3_R1179_U184;
  assign new_P3_R1179_U174 = ~new_P3_U3443;
  assign new_P3_R1179_U175 = ~new_P3_R1179_U274 | ~new_P3_R1179_U273;
  assign new_P3_R1179_U176 = ~new_P3_R1179_U270 | ~new_P3_R1179_U269;
  assign new_P3_R1179_U177 = new_P3_R1179_U462 & new_P3_R1179_U461;
  assign new_P3_R1179_U178 = new_P3_R1179_U466 & new_P3_R1179_U465;
  assign new_P3_R1179_U179 = ~new_P3_R1179_U260 | ~new_P3_R1179_U259;
  assign new_P3_R1179_U180 = ~new_P3_R1179_U256 | ~new_P3_R1179_U255;
  assign new_P3_R1179_U181 = ~new_P3_R1179_U252 | ~new_P3_R1179_U251;
  assign new_P3_R1179_U182 = new_P3_R1179_U483 & new_P3_R1179_U482;
  assign new_P3_R1179_U183 = ~new_P3_R1179_U132 | ~new_P3_R1179_U163;
  assign new_P3_R1179_U184 = ~new_P3_R1179_U175 | ~new_P3_R1179_U174;
  assign new_P3_R1179_U185 = ~new_P3_R1179_U172 | ~new_P3_R1179_U171;
  assign new_P3_R1179_U186 = ~new_P3_R1179_U87;
  assign new_P3_R1179_U187 = ~new_P3_R1179_U34;
  assign new_P3_R1179_U188 = ~new_P3_R1179_U26;
  assign new_P3_R1179_U189 = ~new_P3_U3419 | ~new_P3_R1179_U54;
  assign new_P3_R1179_U190 = ~new_P3_U3434 | ~new_P3_R1179_U64;
  assign new_P3_R1179_U191 = ~new_P3_U3905 | ~new_P3_R1179_U78;
  assign new_P3_R1179_U192 = ~new_P3_U3901 | ~new_P3_R1179_U86;
  assign new_P3_R1179_U193 = ~new_P3_U3395 | ~new_P3_R1179_U33;
  assign new_P3_R1179_U194 = ~new_P3_U3404 | ~new_P3_R1179_U41;
  assign new_P3_R1179_U195 = ~new_P3_U3410 | ~new_P3_R1179_U25;
  assign new_P3_R1179_U196 = ~new_P3_R1179_U66;
  assign new_P3_R1179_U197 = ~new_P3_R1179_U80;
  assign new_P3_R1179_U198 = ~new_P3_R1179_U43;
  assign new_P3_R1179_U199 = ~new_P3_R1179_U55;
  assign new_P3_R1179_U200 = ~new_P3_R1179_U172;
  assign new_P3_R1179_U201 = ~new_P3_U3077 | ~new_P3_R1179_U172;
  assign new_P3_R1179_U202 = ~new_P3_R1179_U49;
  assign new_P3_R1179_U203 = ~new_P3_R1179_U117 | ~new_P3_R1179_U49;
  assign new_P3_R1179_U204 = ~new_P3_R1179_U35 | ~new_P3_R1179_U34;
  assign new_P3_R1179_U205 = ~new_P3_R1179_U204 | ~new_P3_R1179_U32;
  assign new_P3_R1179_U206 = ~new_P3_U3063 | ~new_P3_R1179_U187;
  assign new_P3_R1179_U207 = ~new_P3_R1179_U158;
  assign new_P3_R1179_U208 = ~new_P3_U3407 | ~new_P3_R1179_U40;
  assign new_P3_R1179_U209 = ~new_P3_U3070 | ~new_P3_R1179_U37;
  assign new_P3_R1179_U210 = ~new_P3_U3066 | ~new_P3_R1179_U36;
  assign new_P3_R1179_U211 = ~new_P3_R1179_U198 | ~new_P3_R1179_U194;
  assign new_P3_R1179_U212 = ~new_P3_R1179_U6 | ~new_P3_R1179_U211;
  assign new_P3_R1179_U213 = ~new_P3_U3401 | ~new_P3_R1179_U42;
  assign new_P3_R1179_U214 = ~new_P3_U3407 | ~new_P3_R1179_U40;
  assign new_P3_R1179_U215 = ~new_P3_R1179_U13 | ~new_P3_R1179_U158;
  assign new_P3_R1179_U216 = ~new_P3_R1179_U44;
  assign new_P3_R1179_U217 = ~new_P3_R1179_U47;
  assign new_P3_R1179_U218 = ~new_P3_U3413 | ~new_P3_R1179_U27;
  assign new_P3_R1179_U219 = ~new_P3_R1179_U27 | ~new_P3_R1179_U26;
  assign new_P3_R1179_U220 = ~new_P3_U3083 | ~new_P3_R1179_U188;
  assign new_P3_R1179_U221 = ~new_P3_R1179_U154;
  assign new_P3_R1179_U222 = ~new_P3_U3416 | ~new_P3_R1179_U46;
  assign new_P3_R1179_U223 = ~new_P3_R1179_U222 | ~new_P3_R1179_U55;
  assign new_P3_R1179_U224 = ~new_P3_R1179_U217 | ~new_P3_R1179_U26;
  assign new_P3_R1179_U225 = ~new_P3_R1179_U122 | ~new_P3_R1179_U224;
  assign new_P3_R1179_U226 = ~new_P3_R1179_U47 | ~new_P3_R1179_U195;
  assign new_P3_R1179_U227 = ~new_P3_R1179_U121 | ~new_P3_R1179_U226;
  assign new_P3_R1179_U228 = ~new_P3_R1179_U26 | ~new_P3_R1179_U195;
  assign new_P3_R1179_U229 = ~new_P3_R1179_U213 | ~new_P3_R1179_U158;
  assign new_P3_R1179_U230 = ~new_P3_R1179_U48;
  assign new_P3_R1179_U231 = ~new_P3_U3066 | ~new_P3_R1179_U36;
  assign new_P3_R1179_U232 = ~new_P3_R1179_U230 | ~new_P3_R1179_U231;
  assign new_P3_R1179_U233 = ~new_P3_R1179_U124 | ~new_P3_R1179_U232;
  assign new_P3_R1179_U234 = ~new_P3_R1179_U48 | ~new_P3_R1179_U194;
  assign new_P3_R1179_U235 = ~new_P3_U3407 | ~new_P3_R1179_U40;
  assign new_P3_R1179_U236 = ~new_P3_R1179_U123 | ~new_P3_R1179_U234;
  assign new_P3_R1179_U237 = ~new_P3_U3066 | ~new_P3_R1179_U36;
  assign new_P3_R1179_U238 = ~new_P3_R1179_U194 | ~new_P3_R1179_U237;
  assign new_P3_R1179_U239 = ~new_P3_R1179_U213 | ~new_P3_R1179_U43;
  assign new_P3_R1179_U240 = ~new_P3_R1179_U202 | ~new_P3_R1179_U34;
  assign new_P3_R1179_U241 = ~new_P3_R1179_U126 | ~new_P3_R1179_U240;
  assign new_P3_R1179_U242 = ~new_P3_R1179_U49 | ~new_P3_R1179_U193;
  assign new_P3_R1179_U243 = ~new_P3_R1179_U125 | ~new_P3_R1179_U242;
  assign new_P3_R1179_U244 = ~new_P3_R1179_U193 | ~new_P3_R1179_U34;
  assign new_P3_R1179_U245 = ~new_P3_U3422 | ~new_P3_R1179_U53;
  assign new_P3_R1179_U246 = ~new_P3_U3062 | ~new_P3_R1179_U51;
  assign new_P3_R1179_U247 = ~new_P3_U3061 | ~new_P3_R1179_U52;
  assign new_P3_R1179_U248 = ~new_P3_R1179_U199 | ~new_P3_R1179_U7;
  assign new_P3_R1179_U249 = ~new_P3_R1179_U8 | ~new_P3_R1179_U248;
  assign new_P3_R1179_U250 = ~new_P3_U3422 | ~new_P3_R1179_U53;
  assign new_P3_R1179_U251 = ~new_P3_R1179_U127 | ~new_P3_R1179_U154;
  assign new_P3_R1179_U252 = ~new_P3_R1179_U250 | ~new_P3_R1179_U249;
  assign new_P3_R1179_U253 = ~new_P3_R1179_U181;
  assign new_P3_R1179_U254 = ~new_P3_U3425 | ~new_P3_R1179_U57;
  assign new_P3_R1179_U255 = ~new_P3_R1179_U254 | ~new_P3_R1179_U181;
  assign new_P3_R1179_U256 = ~new_P3_U3071 | ~new_P3_R1179_U56;
  assign new_P3_R1179_U257 = ~new_P3_R1179_U180;
  assign new_P3_R1179_U258 = ~new_P3_U3428 | ~new_P3_R1179_U59;
  assign new_P3_R1179_U259 = ~new_P3_R1179_U258 | ~new_P3_R1179_U180;
  assign new_P3_R1179_U260 = ~new_P3_U3079 | ~new_P3_R1179_U58;
  assign new_P3_R1179_U261 = ~new_P3_R1179_U179;
  assign new_P3_R1179_U262 = ~new_P3_U3437 | ~new_P3_R1179_U63;
  assign new_P3_R1179_U263 = ~new_P3_U3072 | ~new_P3_R1179_U60;
  assign new_P3_R1179_U264 = ~new_P3_U3073 | ~new_P3_R1179_U61;
  assign new_P3_R1179_U265 = ~new_P3_R1179_U196 | ~new_P3_R1179_U9;
  assign new_P3_R1179_U266 = ~new_P3_R1179_U10 | ~new_P3_R1179_U265;
  assign new_P3_R1179_U267 = ~new_P3_U3431 | ~new_P3_R1179_U65;
  assign new_P3_R1179_U268 = ~new_P3_U3437 | ~new_P3_R1179_U63;
  assign new_P3_R1179_U269 = ~new_P3_R1179_U128 | ~new_P3_R1179_U179;
  assign new_P3_R1179_U270 = ~new_P3_R1179_U268 | ~new_P3_R1179_U266;
  assign new_P3_R1179_U271 = ~new_P3_R1179_U176;
  assign new_P3_R1179_U272 = ~new_P3_U3440 | ~new_P3_R1179_U68;
  assign new_P3_R1179_U273 = ~new_P3_R1179_U272 | ~new_P3_R1179_U176;
  assign new_P3_R1179_U274 = ~new_P3_U3068 | ~new_P3_R1179_U67;
  assign new_P3_R1179_U275 = ~new_P3_R1179_U175;
  assign new_P3_R1179_U276 = ~new_P3_U3081 | ~new_P3_R1179_U175;
  assign new_P3_R1179_U277 = ~new_P3_R1179_U173;
  assign new_P3_R1179_U278 = ~new_P3_U3445 | ~new_P3_R1179_U71;
  assign new_P3_R1179_U279 = ~new_P3_R1179_U278 | ~new_P3_R1179_U173;
  assign new_P3_R1179_U280 = ~new_P3_U3080 | ~new_P3_R1179_U70;
  assign new_P3_R1179_U281 = ~new_P3_R1179_U170;
  assign new_P3_R1179_U282 = ~new_P3_U3907 | ~new_P3_R1179_U73;
  assign new_P3_R1179_U283 = ~new_P3_R1179_U282 | ~new_P3_R1179_U170;
  assign new_P3_R1179_U284 = ~new_P3_U3075 | ~new_P3_R1179_U72;
  assign new_P3_R1179_U285 = ~new_P3_R1179_U169;
  assign new_P3_R1179_U286 = ~new_P3_U3904 | ~new_P3_R1179_U77;
  assign new_P3_R1179_U287 = ~new_P3_U3065 | ~new_P3_R1179_U74;
  assign new_P3_R1179_U288 = ~new_P3_U3060 | ~new_P3_R1179_U75;
  assign new_P3_R1179_U289 = ~new_P3_R1179_U197 | ~new_P3_R1179_U11;
  assign new_P3_R1179_U290 = ~new_P3_R1179_U12 | ~new_P3_R1179_U289;
  assign new_P3_R1179_U291 = ~new_P3_U3906 | ~new_P3_R1179_U79;
  assign new_P3_R1179_U292 = ~new_P3_U3904 | ~new_P3_R1179_U77;
  assign new_P3_R1179_U293 = ~new_P3_R1179_U129 | ~new_P3_R1179_U169;
  assign new_P3_R1179_U294 = ~new_P3_R1179_U292 | ~new_P3_R1179_U290;
  assign new_P3_R1179_U295 = ~new_P3_R1179_U166;
  assign new_P3_R1179_U296 = ~new_P3_U3903 | ~new_P3_R1179_U82;
  assign new_P3_R1179_U297 = ~new_P3_R1179_U296 | ~new_P3_R1179_U166;
  assign new_P3_R1179_U298 = ~new_P3_U3064 | ~new_P3_R1179_U81;
  assign new_P3_R1179_U299 = ~new_P3_R1179_U165;
  assign new_P3_R1179_U300 = ~new_P3_U3902 | ~new_P3_R1179_U84;
  assign new_P3_R1179_U301 = ~new_P3_R1179_U300 | ~new_P3_R1179_U165;
  assign new_P3_R1179_U302 = ~new_P3_U3057 | ~new_P3_R1179_U83;
  assign new_P3_R1179_U303 = ~new_P3_R1179_U91;
  assign new_P3_R1179_U304 = ~new_P3_R1179_U130 | ~new_P3_R1179_U91;
  assign new_P3_R1179_U305 = ~new_P3_R1179_U88 | ~new_P3_R1179_U87;
  assign new_P3_R1179_U306 = ~new_P3_R1179_U305 | ~new_P3_R1179_U85;
  assign new_P3_R1179_U307 = ~new_P3_U3052 | ~new_P3_R1179_U186;
  assign new_P3_R1179_U308 = ~new_P3_R1179_U163;
  assign new_P3_R1179_U309 = ~new_P3_U3899 | ~new_P3_R1179_U90;
  assign new_P3_R1179_U310 = ~new_P3_U3053 | ~new_P3_R1179_U89;
  assign new_P3_R1179_U311 = ~new_P3_R1179_U303 | ~new_P3_R1179_U87;
  assign new_P3_R1179_U312 = ~new_P3_R1179_U137 | ~new_P3_R1179_U311;
  assign new_P3_R1179_U313 = ~new_P3_R1179_U91 | ~new_P3_R1179_U192;
  assign new_P3_R1179_U314 = ~new_P3_R1179_U136 | ~new_P3_R1179_U313;
  assign new_P3_R1179_U315 = ~new_P3_R1179_U192 | ~new_P3_R1179_U87;
  assign new_P3_R1179_U316 = ~new_P3_R1179_U291 | ~new_P3_R1179_U169;
  assign new_P3_R1179_U317 = ~new_P3_R1179_U92;
  assign new_P3_R1179_U318 = ~new_P3_U3060 | ~new_P3_R1179_U75;
  assign new_P3_R1179_U319 = ~new_P3_R1179_U317 | ~new_P3_R1179_U318;
  assign new_P3_R1179_U320 = ~new_P3_R1179_U141 | ~new_P3_R1179_U319;
  assign new_P3_R1179_U321 = ~new_P3_R1179_U92 | ~new_P3_R1179_U191;
  assign new_P3_R1179_U322 = ~new_P3_U3904 | ~new_P3_R1179_U77;
  assign new_P3_R1179_U323 = ~new_P3_R1179_U140 | ~new_P3_R1179_U321;
  assign new_P3_R1179_U324 = ~new_P3_U3060 | ~new_P3_R1179_U75;
  assign new_P3_R1179_U325 = ~new_P3_R1179_U191 | ~new_P3_R1179_U324;
  assign new_P3_R1179_U326 = ~new_P3_R1179_U291 | ~new_P3_R1179_U80;
  assign new_P3_R1179_U327 = ~new_P3_R1179_U267 | ~new_P3_R1179_U179;
  assign new_P3_R1179_U328 = ~new_P3_R1179_U93;
  assign new_P3_R1179_U329 = ~new_P3_U3073 | ~new_P3_R1179_U61;
  assign new_P3_R1179_U330 = ~new_P3_R1179_U328 | ~new_P3_R1179_U329;
  assign new_P3_R1179_U331 = ~new_P3_R1179_U148 | ~new_P3_R1179_U330;
  assign new_P3_R1179_U332 = ~new_P3_R1179_U93 | ~new_P3_R1179_U190;
  assign new_P3_R1179_U333 = ~new_P3_U3437 | ~new_P3_R1179_U63;
  assign new_P3_R1179_U334 = ~new_P3_R1179_U147 | ~new_P3_R1179_U332;
  assign new_P3_R1179_U335 = ~new_P3_U3073 | ~new_P3_R1179_U61;
  assign new_P3_R1179_U336 = ~new_P3_R1179_U190 | ~new_P3_R1179_U335;
  assign new_P3_R1179_U337 = ~new_P3_R1179_U267 | ~new_P3_R1179_U66;
  assign new_P3_R1179_U338 = ~new_P3_R1179_U222 | ~new_P3_R1179_U154;
  assign new_P3_R1179_U339 = ~new_P3_R1179_U94;
  assign new_P3_R1179_U340 = ~new_P3_U3061 | ~new_P3_R1179_U52;
  assign new_P3_R1179_U341 = ~new_P3_R1179_U339 | ~new_P3_R1179_U340;
  assign new_P3_R1179_U342 = ~new_P3_R1179_U152 | ~new_P3_R1179_U341;
  assign new_P3_R1179_U343 = ~new_P3_R1179_U94 | ~new_P3_R1179_U189;
  assign new_P3_R1179_U344 = ~new_P3_U3422 | ~new_P3_R1179_U53;
  assign new_P3_R1179_U345 = ~new_P3_R1179_U151 | ~new_P3_R1179_U343;
  assign new_P3_R1179_U346 = ~new_P3_U3061 | ~new_P3_R1179_U52;
  assign new_P3_R1179_U347 = ~new_P3_R1179_U189 | ~new_P3_R1179_U346;
  assign new_P3_R1179_U348 = ~new_P3_U3076 | ~new_P3_R1179_U30;
  assign new_P3_R1179_U349 = ~new_P3_U3077 | ~new_P3_R1179_U171;
  assign new_P3_R1179_U350 = ~new_P3_U3081 | ~new_P3_R1179_U174;
  assign new_P3_R1179_U351 = ~new_P3_R1179_U134 | ~new_P3_R1179_U133 | ~new_P3_R1179_U304;
  assign new_P3_R1179_U352 = ~new_P3_U3398 | ~new_P3_R1179_U35;
  assign new_P3_R1179_U353 = ~new_P3_U3413 | ~new_P3_R1179_U220;
  assign new_P3_R1179_U354 = ~new_P3_R1179_U353 | ~new_P3_R1179_U219;
  assign new_P3_R1179_U355 = ~new_P3_U3900 | ~new_P3_R1179_U88;
  assign new_P3_R1179_U356 = ~new_P3_R1179_U119 | ~new_P3_R1179_U158;
  assign new_P3_R1179_U357 = ~new_P3_R1179_U216 | ~new_P3_R1179_U14;
  assign new_P3_R1179_U358 = ~new_P3_U3416 | ~new_P3_R1179_U46;
  assign new_P3_R1179_U359 = ~new_P3_U3082 | ~new_P3_R1179_U45;
  assign new_P3_R1179_U360 = ~new_P3_R1179_U223 | ~new_P3_R1179_U154;
  assign new_P3_R1179_U361 = ~new_P3_R1179_U221 | ~new_P3_R1179_U153;
  assign new_P3_R1179_U362 = ~new_P3_U3413 | ~new_P3_R1179_U27;
  assign new_P3_R1179_U363 = ~new_P3_U3083 | ~new_P3_R1179_U28;
  assign new_P3_R1179_U364 = ~new_P3_U3413 | ~new_P3_R1179_U27;
  assign new_P3_R1179_U365 = ~new_P3_U3083 | ~new_P3_R1179_U28;
  assign new_P3_R1179_U366 = ~new_P3_R1179_U365 | ~new_P3_R1179_U364;
  assign new_P3_R1179_U367 = ~new_P3_U3410 | ~new_P3_R1179_U25;
  assign new_P3_R1179_U368 = ~new_P3_U3069 | ~new_P3_R1179_U39;
  assign new_P3_R1179_U369 = ~new_P3_R1179_U228 | ~new_P3_R1179_U47;
  assign new_P3_R1179_U370 = ~new_P3_R1179_U155 | ~new_P3_R1179_U217;
  assign new_P3_R1179_U371 = ~new_P3_U3407 | ~new_P3_R1179_U40;
  assign new_P3_R1179_U372 = ~new_P3_U3070 | ~new_P3_R1179_U37;
  assign new_P3_R1179_U373 = ~new_P3_R1179_U372 | ~new_P3_R1179_U371;
  assign new_P3_R1179_U374 = ~new_P3_U3404 | ~new_P3_R1179_U41;
  assign new_P3_R1179_U375 = ~new_P3_U3066 | ~new_P3_R1179_U36;
  assign new_P3_R1179_U376 = ~new_P3_R1179_U238 | ~new_P3_R1179_U48;
  assign new_P3_R1179_U377 = ~new_P3_R1179_U156 | ~new_P3_R1179_U230;
  assign new_P3_R1179_U378 = ~new_P3_U3401 | ~new_P3_R1179_U42;
  assign new_P3_R1179_U379 = ~new_P3_U3059 | ~new_P3_R1179_U38;
  assign new_P3_R1179_U380 = ~new_P3_R1179_U239 | ~new_P3_R1179_U158;
  assign new_P3_R1179_U381 = ~new_P3_R1179_U207 | ~new_P3_R1179_U157;
  assign new_P3_R1179_U382 = ~new_P3_U3398 | ~new_P3_R1179_U35;
  assign new_P3_R1179_U383 = ~new_P3_U3063 | ~new_P3_R1179_U32;
  assign new_P3_R1179_U384 = ~new_P3_U3398 | ~new_P3_R1179_U35;
  assign new_P3_R1179_U385 = ~new_P3_U3063 | ~new_P3_R1179_U32;
  assign new_P3_R1179_U386 = ~new_P3_R1179_U385 | ~new_P3_R1179_U384;
  assign new_P3_R1179_U387 = ~new_P3_U3395 | ~new_P3_R1179_U33;
  assign new_P3_R1179_U388 = ~new_P3_U3067 | ~new_P3_R1179_U29;
  assign new_P3_R1179_U389 = ~new_P3_R1179_U244 | ~new_P3_R1179_U49;
  assign new_P3_R1179_U390 = ~new_P3_R1179_U159 | ~new_P3_R1179_U202;
  assign new_P3_R1179_U391 = ~new_P3_U3908 | ~new_P3_R1179_U161;
  assign new_P3_R1179_U392 = ~new_P3_U3054 | ~new_P3_R1179_U160;
  assign new_P3_R1179_U393 = ~new_P3_U3908 | ~new_P3_R1179_U161;
  assign new_P3_R1179_U394 = ~new_P3_U3054 | ~new_P3_R1179_U160;
  assign new_P3_R1179_U395 = ~new_P3_R1179_U394 | ~new_P3_R1179_U393;
  assign new_P3_R1179_U396 = ~new_P3_R1179_U89 | ~new_P3_U3053 | ~new_P3_R1179_U395;
  assign new_P3_R1179_U397 = ~new_P3_U3899 | ~new_P3_R1179_U15 | ~new_P3_R1179_U90;
  assign new_P3_R1179_U398 = ~new_P3_U3899 | ~new_P3_R1179_U90;
  assign new_P3_R1179_U399 = ~new_P3_U3053 | ~new_P3_R1179_U89;
  assign new_P3_R1179_U400 = ~new_P3_R1179_U135;
  assign new_P3_R1179_U401 = ~new_P3_R1179_U308 | ~new_P3_R1179_U400;
  assign new_P3_R1179_U402 = ~new_P3_R1179_U135 | ~new_P3_R1179_U163;
  assign new_P3_R1179_U403 = ~new_P3_U3900 | ~new_P3_R1179_U88;
  assign new_P3_R1179_U404 = ~new_P3_U3052 | ~new_P3_R1179_U85;
  assign new_P3_R1179_U405 = ~new_P3_U3900 | ~new_P3_R1179_U88;
  assign new_P3_R1179_U406 = ~new_P3_U3052 | ~new_P3_R1179_U85;
  assign new_P3_R1179_U407 = ~new_P3_R1179_U406 | ~new_P3_R1179_U405;
  assign new_P3_R1179_U408 = ~new_P3_U3901 | ~new_P3_R1179_U86;
  assign new_P3_R1179_U409 = ~new_P3_U3056 | ~new_P3_R1179_U50;
  assign new_P3_R1179_U410 = ~new_P3_R1179_U315 | ~new_P3_R1179_U91;
  assign new_P3_R1179_U411 = ~new_P3_R1179_U164 | ~new_P3_R1179_U303;
  assign new_P3_R1179_U412 = ~new_P3_U3902 | ~new_P3_R1179_U84;
  assign new_P3_R1179_U413 = ~new_P3_U3057 | ~new_P3_R1179_U83;
  assign new_P3_R1179_U414 = ~new_P3_R1179_U138;
  assign new_P3_R1179_U415 = ~new_P3_R1179_U299 | ~new_P3_R1179_U414;
  assign new_P3_R1179_U416 = ~new_P3_R1179_U138 | ~new_P3_R1179_U165;
  assign new_P3_R1179_U417 = ~new_P3_U3903 | ~new_P3_R1179_U82;
  assign new_P3_R1179_U418 = ~new_P3_U3064 | ~new_P3_R1179_U81;
  assign new_P3_R1179_U419 = ~new_P3_R1179_U139;
  assign new_P3_R1179_U420 = ~new_P3_R1179_U295 | ~new_P3_R1179_U419;
  assign new_P3_R1179_U421 = ~new_P3_R1179_U139 | ~new_P3_R1179_U166;
  assign new_P3_R1179_U422 = ~new_P3_U3904 | ~new_P3_R1179_U77;
  assign new_P3_R1179_U423 = ~new_P3_U3065 | ~new_P3_R1179_U74;
  assign new_P3_R1179_U424 = ~new_P3_R1179_U423 | ~new_P3_R1179_U422;
  assign new_P3_R1179_U425 = ~new_P3_U3905 | ~new_P3_R1179_U78;
  assign new_P3_R1179_U426 = ~new_P3_U3060 | ~new_P3_R1179_U75;
  assign new_P3_R1179_U427 = ~new_P3_R1179_U325 | ~new_P3_R1179_U92;
  assign new_P3_R1179_U428 = ~new_P3_R1179_U167 | ~new_P3_R1179_U317;
  assign new_P3_R1179_U429 = ~new_P3_U3906 | ~new_P3_R1179_U79;
  assign new_P3_R1179_U430 = ~new_P3_U3074 | ~new_P3_R1179_U76;
  assign new_P3_R1179_U431 = ~new_P3_R1179_U326 | ~new_P3_R1179_U169;
  assign new_P3_R1179_U432 = ~new_P3_R1179_U285 | ~new_P3_R1179_U168;
  assign new_P3_R1179_U433 = ~new_P3_U3907 | ~new_P3_R1179_U73;
  assign new_P3_R1179_U434 = ~new_P3_U3075 | ~new_P3_R1179_U72;
  assign new_P3_R1179_U435 = ~new_P3_R1179_U142;
  assign new_P3_R1179_U436 = ~new_P3_R1179_U281 | ~new_P3_R1179_U435;
  assign new_P3_R1179_U437 = ~new_P3_R1179_U142 | ~new_P3_R1179_U170;
  assign new_P3_R1179_U438 = ~new_P3_U3392 | ~new_P3_R1179_U31;
  assign new_P3_R1179_U439 = ~new_P3_U3077 | ~new_P3_R1179_U171;
  assign new_P3_R1179_U440 = ~new_P3_R1179_U143;
  assign new_P3_R1179_U441 = ~new_P3_R1179_U200 | ~new_P3_R1179_U440;
  assign new_P3_R1179_U442 = ~new_P3_R1179_U143 | ~new_P3_R1179_U172;
  assign new_P3_R1179_U443 = ~new_P3_U3445 | ~new_P3_R1179_U71;
  assign new_P3_R1179_U444 = ~new_P3_U3080 | ~new_P3_R1179_U70;
  assign new_P3_R1179_U445 = ~new_P3_R1179_U144;
  assign new_P3_R1179_U446 = ~new_P3_R1179_U277 | ~new_P3_R1179_U445;
  assign new_P3_R1179_U447 = ~new_P3_R1179_U144 | ~new_P3_R1179_U173;
  assign new_P3_R1179_U448 = ~new_P3_U3443 | ~new_P3_R1179_U69;
  assign new_P3_R1179_U449 = ~new_P3_U3081 | ~new_P3_R1179_U174;
  assign new_P3_R1179_U450 = ~new_P3_R1179_U145;
  assign new_P3_R1179_U451 = ~new_P3_R1179_U275 | ~new_P3_R1179_U450;
  assign new_P3_R1179_U452 = ~new_P3_R1179_U145 | ~new_P3_R1179_U175;
  assign new_P3_R1179_U453 = ~new_P3_U3440 | ~new_P3_R1179_U68;
  assign new_P3_R1179_U454 = ~new_P3_U3068 | ~new_P3_R1179_U67;
  assign new_P3_R1179_U455 = ~new_P3_R1179_U146;
  assign new_P3_R1179_U456 = ~new_P3_R1179_U271 | ~new_P3_R1179_U455;
  assign new_P3_R1179_U457 = ~new_P3_R1179_U146 | ~new_P3_R1179_U176;
  assign new_P3_R1179_U458 = ~new_P3_U3437 | ~new_P3_R1179_U63;
  assign new_P3_R1179_U459 = ~new_P3_U3072 | ~new_P3_R1179_U60;
  assign new_P3_R1179_U460 = ~new_P3_R1179_U459 | ~new_P3_R1179_U458;
  assign new_P3_R1179_U461 = ~new_P3_U3434 | ~new_P3_R1179_U64;
  assign new_P3_R1179_U462 = ~new_P3_U3073 | ~new_P3_R1179_U61;
  assign new_P3_R1179_U463 = ~new_P3_R1179_U336 | ~new_P3_R1179_U93;
  assign new_P3_R1179_U464 = ~new_P3_R1179_U177 | ~new_P3_R1179_U328;
  assign new_P3_R1179_U465 = ~new_P3_U3431 | ~new_P3_R1179_U65;
  assign new_P3_R1179_U466 = ~new_P3_U3078 | ~new_P3_R1179_U62;
  assign new_P3_R1179_U467 = ~new_P3_R1179_U337 | ~new_P3_R1179_U179;
  assign new_P3_R1179_U468 = ~new_P3_R1179_U261 | ~new_P3_R1179_U178;
  assign new_P3_R1179_U469 = ~new_P3_U3428 | ~new_P3_R1179_U59;
  assign new_P3_R1179_U470 = ~new_P3_U3079 | ~new_P3_R1179_U58;
  assign new_P3_R1179_U471 = ~new_P3_R1179_U149;
  assign new_P3_R1179_U472 = ~new_P3_R1179_U257 | ~new_P3_R1179_U471;
  assign new_P3_R1179_U473 = ~new_P3_R1179_U149 | ~new_P3_R1179_U180;
  assign new_P3_R1179_U474 = ~new_P3_U3425 | ~new_P3_R1179_U57;
  assign new_P3_R1179_U475 = ~new_P3_U3071 | ~new_P3_R1179_U56;
  assign new_P3_R1179_U476 = ~new_P3_R1179_U150;
  assign new_P3_R1179_U477 = ~new_P3_R1179_U253 | ~new_P3_R1179_U476;
  assign new_P3_R1179_U478 = ~new_P3_R1179_U150 | ~new_P3_R1179_U181;
  assign new_P3_R1179_U479 = ~new_P3_U3422 | ~new_P3_R1179_U53;
  assign new_P3_R1179_U480 = ~new_P3_U3062 | ~new_P3_R1179_U51;
  assign new_P3_R1179_U481 = ~new_P3_R1179_U480 | ~new_P3_R1179_U479;
  assign new_P3_R1179_U482 = ~new_P3_U3419 | ~new_P3_R1179_U54;
  assign new_P3_R1179_U483 = ~new_P3_U3061 | ~new_P3_R1179_U52;
  assign new_P3_R1179_U484 = ~new_P3_R1179_U347 | ~new_P3_R1179_U94;
  assign new_P3_R1179_U485 = ~new_P3_R1179_U182 | ~new_P3_R1179_U339;
  assign new_P3_R1269_U6 = new_P3_R1269_U107 & new_P3_R1269_U108;
  assign new_P3_R1269_U7 = new_P3_R1269_U118 & new_P3_R1269_U117;
  assign new_P3_R1269_U8 = new_P3_R1269_U142 & new_P3_R1269_U141;
  assign new_P3_R1269_U9 = new_P3_R1269_U200 & new_P3_R1269_U199;
  assign new_P3_R1269_U10 = new_P3_R1269_U202 & new_P3_R1269_U201;
  assign new_P3_R1269_U11 = ~new_P3_R1269_U196 | ~new_P3_R1269_U10 | ~new_P3_R1269_U194;
  assign new_P3_R1269_U12 = ~new_P3_U3116;
  assign new_P3_R1269_U13 = ~new_P3_U3094;
  assign new_P3_R1269_U14 = ~new_P3_U3095;
  assign new_P3_R1269_U15 = ~new_P3_U3130;
  assign new_P3_R1269_U16 = ~new_P3_U3136;
  assign new_P3_R1269_U17 = ~new_P3_U3135;
  assign new_P3_R1269_U18 = ~new_P3_U3106;
  assign new_P3_R1269_U19 = ~new_P3_U3107;
  assign new_P3_R1269_U20 = ~new_P3_U3112;
  assign new_P3_R1269_U21 = ~new_P3_U3113;
  assign new_P3_R1269_U22 = ~new_P3_U3114;
  assign new_P3_R1269_U23 = ~new_P3_U3142;
  assign new_P3_R1269_U24 = ~new_P3_U3141;
  assign new_P3_R1269_U25 = ~new_P3_U3146;
  assign new_P3_R1269_U26 = ~new_P3_U3145;
  assign new_P3_R1269_U27 = ~new_P3_U3144;
  assign new_P3_R1269_U28 = ~new_P3_U3143;
  assign new_P3_R1269_U29 = ~new_P3_U3111;
  assign new_P3_R1269_U30 = ~new_P3_U3109;
  assign new_P3_R1269_U31 = ~new_P3_U3110;
  assign new_P3_R1269_U32 = ~new_P3_U3108;
  assign new_P3_R1269_U33 = ~new_P3_U3140;
  assign new_P3_R1269_U34 = ~new_P3_U3139;
  assign new_P3_R1269_U35 = ~new_P3_U3138;
  assign new_P3_R1269_U36 = ~new_P3_U3137;
  assign new_P3_R1269_U37 = ~new_P3_U3101;
  assign new_P3_R1269_U38 = ~new_P3_U3100;
  assign new_P3_R1269_U39 = ~new_P3_U3104;
  assign new_P3_R1269_U40 = ~new_P3_U3105;
  assign new_P3_R1269_U41 = ~new_P3_U3103;
  assign new_P3_R1269_U42 = ~new_P3_U3102;
  assign new_P3_R1269_U43 = ~new_P3_U3134;
  assign new_P3_R1269_U44 = ~new_P3_U3133;
  assign new_P3_R1269_U45 = ~new_P3_U3132;
  assign new_P3_R1269_U46 = ~new_P3_U3131;
  assign new_P3_R1269_U47 = ~new_P3_U3099;
  assign new_P3_R1269_U48 = ~new_P3_U3098;
  assign new_P3_R1269_U49 = ~new_P3_R1269_U157 | ~new_P3_R1269_U156;
  assign new_P3_R1269_U50 = ~new_P3_U3129;
  assign new_P3_R1269_U51 = ~new_P3_U3096;
  assign new_P3_R1269_U52 = ~new_P3_U3123;
  assign new_P3_R1269_U53 = ~new_P3_U3124;
  assign new_P3_R1269_U54 = ~new_P3_U3128;
  assign new_P3_R1269_U55 = ~new_P3_U3127;
  assign new_P3_R1269_U56 = ~new_P3_U3126;
  assign new_P3_R1269_U57 = ~new_P3_U3125;
  assign new_P3_R1269_U58 = ~new_P3_U3087;
  assign new_P3_R1269_U59 = ~new_P3_U3089;
  assign new_P3_R1269_U60 = ~new_P3_U3088;
  assign new_P3_R1269_U61 = ~new_P3_U3086;
  assign new_P3_R1269_U62 = ~new_P3_U3093;
  assign new_P3_R1269_U63 = ~new_P3_U3092;
  assign new_P3_R1269_U64 = ~new_P3_U3090;
  assign new_P3_R1269_U65 = ~new_P3_U3091;
  assign new_P3_R1269_U66 = ~new_P3_U3120;
  assign new_P3_R1269_U67 = ~new_P3_U3119;
  assign new_P3_R1269_U68 = ~new_P3_R1269_U178 | ~new_P3_R1269_U177;
  assign new_P3_R1269_U69 = ~new_P3_U3121;
  assign new_P3_R1269_U70 = ~new_P3_U3122;
  assign new_P3_R1269_U71 = ~new_P3_U3118;
  assign new_P3_R1269_U72 = ~new_P3_U3149;
  assign new_P3_R1269_U73 = new_P3_R1269_U111 & new_P3_R1269_U110;
  assign new_P3_R1269_U74 = new_P3_R1269_U7 & new_P3_R1269_U124;
  assign new_P3_R1269_U75 = new_P3_U3111 & new_P3_R1269_U28;
  assign new_P3_R1269_U76 = new_P3_U3110 & new_P3_R1269_U23;
  assign new_P3_R1269_U77 = new_P3_R1269_U78 & new_P3_R1269_U126 & new_P3_R1269_U127;
  assign new_P3_R1269_U78 = new_P3_R1269_U130 & new_P3_R1269_U129;
  assign new_P3_R1269_U79 = new_P3_R1269_U6 & new_P3_R1269_U80;
  assign new_P3_R1269_U80 = new_P3_R1269_U138 & new_P3_R1269_U139;
  assign new_P3_R1269_U81 = new_P3_U3104 & new_P3_R1269_U16;
  assign new_P3_R1269_U82 = new_P3_U3105 & new_P3_R1269_U36;
  assign new_P3_R1269_U83 = new_P3_R1269_U85 & new_P3_R1269_U143 & new_P3_R1269_U144;
  assign new_P3_R1269_U84 = new_P3_R1269_U146 & new_P3_R1269_U145;
  assign new_P3_R1269_U85 = new_P3_R1269_U84 & new_P3_R1269_U8;
  assign new_P3_R1269_U86 = new_P3_U3134 & new_P3_R1269_U42;
  assign new_P3_R1269_U87 = new_P3_U3133 & new_P3_R1269_U37;
  assign new_P3_R1269_U88 = new_P3_R1269_U89 & new_P3_R1269_U148 & new_P3_R1269_U150;
  assign new_P3_R1269_U89 = new_P3_R1269_U152 & new_P3_R1269_U151;
  assign new_P3_R1269_U90 = new_P3_R1269_U104 & new_P3_R1269_U103;
  assign new_P3_R1269_U91 = new_P3_R1269_U162 & new_P3_R1269_U161;
  assign new_P3_R1269_U92 = new_P3_U3128 & new_P3_R1269_U51;
  assign new_P3_R1269_U93 = new_P3_R1269_U165 & new_P3_R1269_U171 & new_P3_R1269_U170 & new_P3_R1269_U169;
  assign new_P3_R1269_U94 = new_P3_R1269_U175 & new_P3_R1269_U174;
  assign new_P3_R1269_U95 = new_P3_R1269_U176 & new_P3_R1269_U96 & new_P3_R1269_U173 & new_P3_R1269_U172 & new_P3_R1269_U94;
  assign new_P3_R1269_U96 = new_P3_R1269_U192 & new_P3_R1269_U193 & new_P3_R1269_U191;
  assign new_P3_R1269_U97 = new_P3_U3120 & new_P3_R1269_U60;
  assign new_P3_R1269_U98 = new_P3_R1269_U174 & new_P3_R1269_U175;
  assign new_P3_R1269_U99 = new_P3_R1269_U198 & new_P3_R1269_U186;
  assign new_P3_R1269_U100 = ~new_P3_U3084;
  assign new_P3_R1269_U101 = ~new_P3_U3085;
  assign new_P3_R1269_U102 = ~new_P3_R1269_U187 | ~new_P3_R1269_U195;
  assign new_P3_R1269_U103 = ~new_P3_U3094 | ~new_P3_R1269_U56;
  assign new_P3_R1269_U104 = ~new_P3_U3095 | ~new_P3_R1269_U55;
  assign new_P3_R1269_U105 = ~new_P3_U3130 | ~new_P3_R1269_U48;
  assign new_P3_R1269_U106 = ~new_P3_U3106 | ~new_P3_R1269_U35;
  assign new_P3_R1269_U107 = ~new_P3_U3135 | ~new_P3_R1269_U41;
  assign new_P3_R1269_U108 = ~new_P3_U3136 | ~new_P3_R1269_U39;
  assign new_P3_R1269_U109 = ~new_P3_U3107 | ~new_P3_R1269_U34;
  assign new_P3_R1269_U110 = ~new_P3_U3112 | ~new_P3_R1269_U27;
  assign new_P3_R1269_U111 = ~new_P3_U3113 | ~new_P3_R1269_U26;
  assign new_P3_R1269_U112 = ~new_P3_U3147 | ~new_P3_U3148;
  assign new_P3_R1269_U113 = ~new_P3_U3115 | ~new_P3_R1269_U112;
  assign new_P3_R1269_U114 = new_P3_U3147 | new_P3_U3148;
  assign new_P3_R1269_U115 = ~new_P3_U3114 | ~new_P3_R1269_U25;
  assign new_P3_R1269_U116 = ~new_P3_R1269_U114 | ~new_P3_R1269_U115 | ~new_P3_R1269_U113 | ~new_P3_R1269_U111 | ~new_P3_R1269_U110;
  assign new_P3_R1269_U117 = ~new_P3_U3142 | ~new_P3_R1269_U31;
  assign new_P3_R1269_U118 = ~new_P3_U3141 | ~new_P3_R1269_U30;
  assign new_P3_R1269_U119 = ~new_P3_U3146 | ~new_P3_R1269_U22;
  assign new_P3_R1269_U120 = ~new_P3_U3145 | ~new_P3_R1269_U21;
  assign new_P3_R1269_U121 = ~new_P3_R1269_U120 | ~new_P3_R1269_U119;
  assign new_P3_R1269_U122 = ~new_P3_R1269_U73 | ~new_P3_R1269_U121;
  assign new_P3_R1269_U123 = ~new_P3_U3144 | ~new_P3_R1269_U20;
  assign new_P3_R1269_U124 = ~new_P3_U3143 | ~new_P3_R1269_U29;
  assign new_P3_R1269_U125 = ~new_P3_R1269_U74 | ~new_P3_R1269_U116 | ~new_P3_R1269_U122 | ~new_P3_R1269_U123;
  assign new_P3_R1269_U126 = ~new_P3_R1269_U75 | ~new_P3_R1269_U7;
  assign new_P3_R1269_U127 = ~new_P3_U3109 | ~new_P3_R1269_U24;
  assign new_P3_R1269_U128 = ~new_P3_U3141 | ~new_P3_R1269_U30;
  assign new_P3_R1269_U129 = ~new_P3_R1269_U76 | ~new_P3_R1269_U128;
  assign new_P3_R1269_U130 = ~new_P3_U3108 | ~new_P3_R1269_U33;
  assign new_P3_R1269_U131 = ~new_P3_R1269_U125 | ~new_P3_R1269_U77;
  assign new_P3_R1269_U132 = ~new_P3_U3140 | ~new_P3_R1269_U32;
  assign new_P3_R1269_U133 = ~new_P3_R1269_U132 | ~new_P3_R1269_U131;
  assign new_P3_R1269_U134 = ~new_P3_R1269_U133 | ~new_P3_R1269_U109;
  assign new_P3_R1269_U135 = ~new_P3_U3139 | ~new_P3_R1269_U19;
  assign new_P3_R1269_U136 = ~new_P3_R1269_U135 | ~new_P3_R1269_U134;
  assign new_P3_R1269_U137 = ~new_P3_R1269_U136 | ~new_P3_R1269_U106;
  assign new_P3_R1269_U138 = ~new_P3_U3138 | ~new_P3_R1269_U18;
  assign new_P3_R1269_U139 = ~new_P3_U3137 | ~new_P3_R1269_U40;
  assign new_P3_R1269_U140 = ~new_P3_R1269_U137 | ~new_P3_R1269_U79;
  assign new_P3_R1269_U141 = ~new_P3_U3101 | ~new_P3_R1269_U44;
  assign new_P3_R1269_U142 = ~new_P3_U3100 | ~new_P3_R1269_U45;
  assign new_P3_R1269_U143 = ~new_P3_R1269_U81 | ~new_P3_R1269_U107;
  assign new_P3_R1269_U144 = ~new_P3_R1269_U82 | ~new_P3_R1269_U6;
  assign new_P3_R1269_U145 = ~new_P3_U3103 | ~new_P3_R1269_U17;
  assign new_P3_R1269_U146 = ~new_P3_U3102 | ~new_P3_R1269_U43;
  assign new_P3_R1269_U147 = ~new_P3_R1269_U140 | ~new_P3_R1269_U83;
  assign new_P3_R1269_U148 = ~new_P3_R1269_U86 | ~new_P3_R1269_U8;
  assign new_P3_R1269_U149 = ~new_P3_U3100 | ~new_P3_R1269_U45;
  assign new_P3_R1269_U150 = ~new_P3_R1269_U87 | ~new_P3_R1269_U149;
  assign new_P3_R1269_U151 = ~new_P3_U3132 | ~new_P3_R1269_U38;
  assign new_P3_R1269_U152 = ~new_P3_U3131 | ~new_P3_R1269_U47;
  assign new_P3_R1269_U153 = ~new_P3_R1269_U147 | ~new_P3_R1269_U88;
  assign new_P3_R1269_U154 = ~new_P3_U3099 | ~new_P3_R1269_U46;
  assign new_P3_R1269_U155 = ~new_P3_R1269_U154 | ~new_P3_R1269_U153;
  assign new_P3_R1269_U156 = ~new_P3_R1269_U155 | ~new_P3_R1269_U105;
  assign new_P3_R1269_U157 = ~new_P3_U3098 | ~new_P3_R1269_U15;
  assign new_P3_R1269_U158 = ~new_P3_R1269_U49;
  assign new_P3_R1269_U159 = ~new_P3_U3129 | ~new_P3_R1269_U158;
  assign new_P3_R1269_U160 = ~new_P3_U3097 | ~new_P3_R1269_U159;
  assign new_P3_R1269_U161 = ~new_P3_R1269_U49 | ~new_P3_R1269_U50;
  assign new_P3_R1269_U162 = ~new_P3_U3096 | ~new_P3_R1269_U54;
  assign new_P3_R1269_U163 = ~new_P3_R1269_U91 | ~new_P3_R1269_U90 | ~new_P3_R1269_U160;
  assign new_P3_R1269_U164 = ~new_P3_U3123 | ~new_P3_R1269_U65;
  assign new_P3_R1269_U165 = ~new_P3_U3124 | ~new_P3_R1269_U63;
  assign new_P3_R1269_U166 = ~new_P3_R1269_U92 | ~new_P3_R1269_U104;
  assign new_P3_R1269_U167 = ~new_P3_U3127 | ~new_P3_R1269_U14;
  assign new_P3_R1269_U168 = ~new_P3_R1269_U167 | ~new_P3_R1269_U166;
  assign new_P3_R1269_U169 = ~new_P3_R1269_U168 | ~new_P3_R1269_U103;
  assign new_P3_R1269_U170 = ~new_P3_U3126 | ~new_P3_R1269_U13;
  assign new_P3_R1269_U171 = ~new_P3_U3125 | ~new_P3_R1269_U62;
  assign new_P3_R1269_U172 = ~new_P3_R1269_U164 | ~new_P3_R1269_U93 | ~new_P3_R1269_U163;
  assign new_P3_R1269_U173 = ~new_P3_U3087 | ~new_P3_R1269_U67;
  assign new_P3_R1269_U174 = ~new_P3_U3089 | ~new_P3_R1269_U69;
  assign new_P3_R1269_U175 = ~new_P3_U3088 | ~new_P3_R1269_U66;
  assign new_P3_R1269_U176 = ~new_P3_U3086 | ~new_P3_R1269_U71;
  assign new_P3_R1269_U177 = ~new_P3_R1269_U97 | ~new_P3_R1269_U173;
  assign new_P3_R1269_U178 = ~new_P3_U3119 | ~new_P3_R1269_U58;
  assign new_P3_R1269_U179 = ~new_P3_R1269_U68;
  assign new_P3_R1269_U180 = ~new_P3_U3121 | ~new_P3_R1269_U59;
  assign new_P3_R1269_U181 = ~new_P3_U3122 | ~new_P3_R1269_U64;
  assign new_P3_R1269_U182 = ~new_P3_R1269_U181 | ~new_P3_R1269_U180;
  assign new_P3_R1269_U183 = ~new_P3_R1269_U179 | ~new_P3_R1269_U71;
  assign new_P3_R1269_U184 = ~new_P3_R1269_U183 | ~new_P3_R1269_U61;
  assign new_P3_R1269_U185 = ~new_P3_R1269_U176 | ~new_P3_R1269_U173 | ~new_P3_R1269_U98 | ~new_P3_R1269_U182;
  assign new_P3_R1269_U186 = ~new_P3_U3118 | ~new_P3_R1269_U68;
  assign new_P3_R1269_U187 = ~new_P3_R1269_U9 | ~new_P3_R1269_U101;
  assign new_P3_R1269_U188 = ~new_P3_U3093 | ~new_P3_R1269_U57;
  assign new_P3_R1269_U189 = ~new_P3_U3092 | ~new_P3_R1269_U53;
  assign new_P3_R1269_U190 = ~new_P3_R1269_U189 | ~new_P3_R1269_U188;
  assign new_P3_R1269_U191 = ~new_P3_R1269_U164 | ~new_P3_R1269_U165 | ~new_P3_R1269_U190;
  assign new_P3_R1269_U192 = ~new_P3_U3090 | ~new_P3_R1269_U70;
  assign new_P3_R1269_U193 = ~new_P3_U3091 | ~new_P3_R1269_U52;
  assign new_P3_R1269_U194 = ~new_P3_R1269_U102 | ~new_P3_R1269_U95;
  assign new_P3_R1269_U195 = ~new_P3_U3117 | ~new_P3_R1269_U9;
  assign new_P3_R1269_U196 = ~new_P3_R1269_U197 | ~new_P3_R1269_U102;
  assign new_P3_R1269_U197 = ~new_P3_R1269_U99 | ~new_P3_R1269_U185 | ~new_P3_R1269_U184;
  assign new_P3_R1269_U198 = ~new_P3_U3117 | ~new_P3_R1269_U101;
  assign new_P3_R1269_U199 = ~new_P3_U3084 | ~new_P3_R1269_U12;
  assign new_P3_R1269_U200 = ~new_P3_U3116 | ~new_P3_R1269_U100;
  assign new_P3_R1269_U201 = ~new_P3_R1269_U100 | ~new_P3_U3116 | ~new_P3_R1269_U72;
  assign new_P3_R1269_U202 = ~new_P3_U3084 | ~new_P3_U3149 | ~new_P3_R1269_U12;
  assign new_P3_R1110_U4 = new_P3_R1110_U179 & new_P3_R1110_U178;
  assign new_P3_R1110_U5 = new_P3_R1110_U197 & new_P3_R1110_U196;
  assign new_P3_R1110_U6 = new_P3_R1110_U237 & new_P3_R1110_U236;
  assign new_P3_R1110_U7 = new_P3_R1110_U246 & new_P3_R1110_U245;
  assign new_P3_R1110_U8 = new_P3_R1110_U264 & new_P3_R1110_U263;
  assign new_P3_R1110_U9 = new_P3_R1110_U272 & new_P3_R1110_U271;
  assign new_P3_R1110_U10 = new_P3_R1110_U351 & new_P3_R1110_U348;
  assign new_P3_R1110_U11 = new_P3_R1110_U344 & new_P3_R1110_U341;
  assign new_P3_R1110_U12 = new_P3_R1110_U335 & new_P3_R1110_U332;
  assign new_P3_R1110_U13 = new_P3_R1110_U326 & new_P3_R1110_U323;
  assign new_P3_R1110_U14 = new_P3_R1110_U320 & new_P3_R1110_U318;
  assign new_P3_R1110_U15 = new_P3_R1110_U313 & new_P3_R1110_U310;
  assign new_P3_R1110_U16 = new_P3_R1110_U235 & new_P3_R1110_U232;
  assign new_P3_R1110_U17 = new_P3_R1110_U227 & new_P3_R1110_U224;
  assign new_P3_R1110_U18 = new_P3_R1110_U213 & new_P3_R1110_U210;
  assign new_P3_R1110_U19 = ~new_P3_U3407;
  assign new_P3_R1110_U20 = ~new_P3_U3070;
  assign new_P3_R1110_U21 = ~new_P3_U3069;
  assign new_P3_R1110_U22 = ~new_P3_U3070 | ~new_P3_U3407;
  assign new_P3_R1110_U23 = ~new_P3_U3410;
  assign new_P3_R1110_U24 = ~new_P3_U3401;
  assign new_P3_R1110_U25 = ~new_P3_U3059;
  assign new_P3_R1110_U26 = ~new_P3_U3066;
  assign new_P3_R1110_U27 = ~new_P3_U3395;
  assign new_P3_R1110_U28 = ~new_P3_U3067;
  assign new_P3_R1110_U29 = ~new_P3_U3387;
  assign new_P3_R1110_U30 = ~new_P3_U3076;
  assign new_P3_R1110_U31 = ~new_P3_U3076 | ~new_P3_U3387;
  assign new_P3_R1110_U32 = ~new_P3_U3398;
  assign new_P3_R1110_U33 = ~new_P3_U3063;
  assign new_P3_R1110_U34 = ~new_P3_U3059 | ~new_P3_U3401;
  assign new_P3_R1110_U35 = ~new_P3_U3404;
  assign new_P3_R1110_U36 = ~new_P3_U3413;
  assign new_P3_R1110_U37 = ~new_P3_U3083;
  assign new_P3_R1110_U38 = ~new_P3_U3082;
  assign new_P3_R1110_U39 = ~new_P3_U3416;
  assign new_P3_R1110_U40 = ~new_P3_R1110_U61 | ~new_P3_R1110_U205;
  assign new_P3_R1110_U41 = ~new_P3_R1110_U117 | ~new_P3_R1110_U193;
  assign new_P3_R1110_U42 = ~new_P3_R1110_U182 | ~new_P3_R1110_U183;
  assign new_P3_R1110_U43 = ~new_P3_U3392 | ~new_P3_U3077;
  assign new_P3_R1110_U44 = ~new_P3_R1110_U122 | ~new_P3_R1110_U219;
  assign new_P3_R1110_U45 = ~new_P3_R1110_U216 | ~new_P3_R1110_U215;
  assign new_P3_R1110_U46 = ~new_P3_U3900;
  assign new_P3_R1110_U47 = ~new_P3_U3052;
  assign new_P3_R1110_U48 = ~new_P3_U3056;
  assign new_P3_R1110_U49 = ~new_P3_U3901;
  assign new_P3_R1110_U50 = ~new_P3_U3902;
  assign new_P3_R1110_U51 = ~new_P3_U3057;
  assign new_P3_R1110_U52 = ~new_P3_U3903;
  assign new_P3_R1110_U53 = ~new_P3_U3064;
  assign new_P3_R1110_U54 = ~new_P3_U3906;
  assign new_P3_R1110_U55 = ~new_P3_U3074;
  assign new_P3_R1110_U56 = ~new_P3_U3437;
  assign new_P3_R1110_U57 = ~new_P3_U3072;
  assign new_P3_R1110_U58 = ~new_P3_U3068;
  assign new_P3_R1110_U59 = ~new_P3_U3072 | ~new_P3_U3437;
  assign new_P3_R1110_U60 = ~new_P3_U3440;
  assign new_P3_R1110_U61 = ~new_P3_U3083 | ~new_P3_U3413;
  assign new_P3_R1110_U62 = ~new_P3_U3419;
  assign new_P3_R1110_U63 = ~new_P3_U3061;
  assign new_P3_R1110_U64 = ~new_P3_U3425;
  assign new_P3_R1110_U65 = ~new_P3_U3071;
  assign new_P3_R1110_U66 = ~new_P3_U3422;
  assign new_P3_R1110_U67 = ~new_P3_U3062;
  assign new_P3_R1110_U68 = ~new_P3_U3062 | ~new_P3_U3422;
  assign new_P3_R1110_U69 = ~new_P3_U3428;
  assign new_P3_R1110_U70 = ~new_P3_U3079;
  assign new_P3_R1110_U71 = ~new_P3_U3431;
  assign new_P3_R1110_U72 = ~new_P3_U3078;
  assign new_P3_R1110_U73 = ~new_P3_U3434;
  assign new_P3_R1110_U74 = ~new_P3_U3073;
  assign new_P3_R1110_U75 = ~new_P3_U3443;
  assign new_P3_R1110_U76 = ~new_P3_U3081;
  assign new_P3_R1110_U77 = ~new_P3_U3081 | ~new_P3_U3443;
  assign new_P3_R1110_U78 = ~new_P3_U3445;
  assign new_P3_R1110_U79 = ~new_P3_U3080;
  assign new_P3_R1110_U80 = ~new_P3_U3080 | ~new_P3_U3445;
  assign new_P3_R1110_U81 = ~new_P3_U3907;
  assign new_P3_R1110_U82 = ~new_P3_U3905;
  assign new_P3_R1110_U83 = ~new_P3_U3060;
  assign new_P3_R1110_U84 = ~new_P3_U3904;
  assign new_P3_R1110_U85 = ~new_P3_U3065;
  assign new_P3_R1110_U86 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1110_U87 = ~new_P3_U3053;
  assign new_P3_R1110_U88 = ~new_P3_U3899;
  assign new_P3_R1110_U89 = ~new_P3_R1110_U306 | ~new_P3_R1110_U176;
  assign new_P3_R1110_U90 = ~new_P3_U3075;
  assign new_P3_R1110_U91 = ~new_P3_R1110_U77 | ~new_P3_R1110_U315;
  assign new_P3_R1110_U92 = ~new_P3_R1110_U261 | ~new_P3_R1110_U260;
  assign new_P3_R1110_U93 = ~new_P3_R1110_U68 | ~new_P3_R1110_U337;
  assign new_P3_R1110_U94 = ~new_P3_R1110_U457 | ~new_P3_R1110_U456;
  assign new_P3_R1110_U95 = ~new_P3_R1110_U504 | ~new_P3_R1110_U503;
  assign new_P3_R1110_U96 = ~new_P3_R1110_U375 | ~new_P3_R1110_U374;
  assign new_P3_R1110_U97 = ~new_P3_R1110_U380 | ~new_P3_R1110_U379;
  assign new_P3_R1110_U98 = ~new_P3_R1110_U387 | ~new_P3_R1110_U386;
  assign new_P3_R1110_U99 = ~new_P3_R1110_U394 | ~new_P3_R1110_U393;
  assign new_P3_R1110_U100 = ~new_P3_R1110_U399 | ~new_P3_R1110_U398;
  assign new_P3_R1110_U101 = ~new_P3_R1110_U408 | ~new_P3_R1110_U407;
  assign new_P3_R1110_U102 = ~new_P3_R1110_U415 | ~new_P3_R1110_U414;
  assign new_P3_R1110_U103 = ~new_P3_R1110_U422 | ~new_P3_R1110_U421;
  assign new_P3_R1110_U104 = ~new_P3_R1110_U429 | ~new_P3_R1110_U428;
  assign new_P3_R1110_U105 = ~new_P3_R1110_U434 | ~new_P3_R1110_U433;
  assign new_P3_R1110_U106 = ~new_P3_R1110_U441 | ~new_P3_R1110_U440;
  assign new_P3_R1110_U107 = ~new_P3_R1110_U448 | ~new_P3_R1110_U447;
  assign new_P3_R1110_U108 = ~new_P3_R1110_U462 | ~new_P3_R1110_U461;
  assign new_P3_R1110_U109 = ~new_P3_R1110_U467 | ~new_P3_R1110_U466;
  assign new_P3_R1110_U110 = ~new_P3_R1110_U474 | ~new_P3_R1110_U473;
  assign new_P3_R1110_U111 = ~new_P3_R1110_U481 | ~new_P3_R1110_U480;
  assign new_P3_R1110_U112 = ~new_P3_R1110_U488 | ~new_P3_R1110_U487;
  assign new_P3_R1110_U113 = ~new_P3_R1110_U495 | ~new_P3_R1110_U494;
  assign new_P3_R1110_U114 = ~new_P3_R1110_U500 | ~new_P3_R1110_U499;
  assign new_P3_R1110_U115 = new_P3_R1110_U189 & new_P3_R1110_U187;
  assign new_P3_R1110_U116 = new_P3_R1110_U4 & new_P3_R1110_U180;
  assign new_P3_R1110_U117 = new_P3_R1110_U194 & new_P3_R1110_U192;
  assign new_P3_R1110_U118 = new_P3_R1110_U201 & new_P3_R1110_U200;
  assign new_P3_R1110_U119 = new_P3_R1110_U22 & new_P3_R1110_U382 & new_P3_R1110_U381;
  assign new_P3_R1110_U120 = new_P3_R1110_U212 & new_P3_R1110_U5;
  assign new_P3_R1110_U121 = new_P3_R1110_U181 & new_P3_R1110_U180;
  assign new_P3_R1110_U122 = new_P3_R1110_U220 & new_P3_R1110_U218;
  assign new_P3_R1110_U123 = new_P3_R1110_U34 & new_P3_R1110_U389 & new_P3_R1110_U388;
  assign new_P3_R1110_U124 = new_P3_R1110_U226 & new_P3_R1110_U4;
  assign new_P3_R1110_U125 = new_P3_R1110_U234 & new_P3_R1110_U181;
  assign new_P3_R1110_U126 = new_P3_R1110_U204 & new_P3_R1110_U6;
  assign new_P3_R1110_U127 = new_P3_R1110_U239 & new_P3_R1110_U171;
  assign new_P3_R1110_U128 = new_P3_R1110_U250 & new_P3_R1110_U7;
  assign new_P3_R1110_U129 = new_P3_R1110_U248 & new_P3_R1110_U172;
  assign new_P3_R1110_U130 = new_P3_R1110_U268 & new_P3_R1110_U267;
  assign new_P3_R1110_U131 = new_P3_R1110_U273 & new_P3_R1110_U9 & new_P3_R1110_U282;
  assign new_P3_R1110_U132 = new_P3_R1110_U285 & new_P3_R1110_U280;
  assign new_P3_R1110_U133 = new_P3_R1110_U301 & new_P3_R1110_U298;
  assign new_P3_R1110_U134 = new_P3_R1110_U368 & new_P3_R1110_U302;
  assign new_P3_R1110_U135 = new_P3_R1110_U160 & new_P3_R1110_U278;
  assign new_P3_R1110_U136 = new_P3_R1110_U80 & new_P3_R1110_U455 & new_P3_R1110_U454;
  assign new_P3_R1110_U137 = new_P3_R1110_U325 & new_P3_R1110_U9;
  assign new_P3_R1110_U138 = new_P3_R1110_U59 & new_P3_R1110_U469 & new_P3_R1110_U468;
  assign new_P3_R1110_U139 = new_P3_R1110_U334 & new_P3_R1110_U8;
  assign new_P3_R1110_U140 = new_P3_R1110_U172 & new_P3_R1110_U490 & new_P3_R1110_U489;
  assign new_P3_R1110_U141 = new_P3_R1110_U343 & new_P3_R1110_U7;
  assign new_P3_R1110_U142 = new_P3_R1110_U171 & new_P3_R1110_U502 & new_P3_R1110_U501;
  assign new_P3_R1110_U143 = new_P3_R1110_U350 & new_P3_R1110_U6;
  assign new_P3_R1110_U144 = ~new_P3_R1110_U118 | ~new_P3_R1110_U202;
  assign new_P3_R1110_U145 = ~new_P3_R1110_U217 | ~new_P3_R1110_U229;
  assign new_P3_R1110_U146 = ~new_P3_U3054;
  assign new_P3_R1110_U147 = ~new_P3_U3908;
  assign new_P3_R1110_U148 = new_P3_R1110_U403 & new_P3_R1110_U402;
  assign new_P3_R1110_U149 = ~new_P3_R1110_U364 | ~new_P3_R1110_U304 | ~new_P3_R1110_U169;
  assign new_P3_R1110_U150 = new_P3_R1110_U410 & new_P3_R1110_U409;
  assign new_P3_R1110_U151 = ~new_P3_R1110_U134 | ~new_P3_R1110_U370 | ~new_P3_R1110_U369;
  assign new_P3_R1110_U152 = new_P3_R1110_U417 & new_P3_R1110_U416;
  assign new_P3_R1110_U153 = ~new_P3_R1110_U86 | ~new_P3_R1110_U365 | ~new_P3_R1110_U299;
  assign new_P3_R1110_U154 = new_P3_R1110_U424 & new_P3_R1110_U423;
  assign new_P3_R1110_U155 = ~new_P3_R1110_U293 | ~new_P3_R1110_U292;
  assign new_P3_R1110_U156 = new_P3_R1110_U436 & new_P3_R1110_U435;
  assign new_P3_R1110_U157 = ~new_P3_R1110_U289 | ~new_P3_R1110_U288;
  assign new_P3_R1110_U158 = new_P3_R1110_U443 & new_P3_R1110_U442;
  assign new_P3_R1110_U159 = ~new_P3_R1110_U132 | ~new_P3_R1110_U284;
  assign new_P3_R1110_U160 = new_P3_R1110_U450 & new_P3_R1110_U449;
  assign new_P3_R1110_U161 = ~new_P3_R1110_U43 | ~new_P3_R1110_U327;
  assign new_P3_R1110_U162 = ~new_P3_R1110_U130 | ~new_P3_R1110_U269;
  assign new_P3_R1110_U163 = new_P3_R1110_U476 & new_P3_R1110_U475;
  assign new_P3_R1110_U164 = ~new_P3_R1110_U257 | ~new_P3_R1110_U256;
  assign new_P3_R1110_U165 = new_P3_R1110_U483 & new_P3_R1110_U482;
  assign new_P3_R1110_U166 = ~new_P3_R1110_U253 | ~new_P3_R1110_U252;
  assign new_P3_R1110_U167 = ~new_P3_R1110_U243 | ~new_P3_R1110_U242;
  assign new_P3_R1110_U168 = ~new_P3_R1110_U367 | ~new_P3_R1110_U366;
  assign new_P3_R1110_U169 = ~new_P3_U3053 | ~new_P3_R1110_U151;
  assign new_P3_R1110_U170 = ~new_P3_R1110_U34;
  assign new_P3_R1110_U171 = ~new_P3_U3416 | ~new_P3_U3082;
  assign new_P3_R1110_U172 = ~new_P3_U3071 | ~new_P3_U3425;
  assign new_P3_R1110_U173 = ~new_P3_U3057 | ~new_P3_U3902;
  assign new_P3_R1110_U174 = ~new_P3_R1110_U68;
  assign new_P3_R1110_U175 = ~new_P3_R1110_U77;
  assign new_P3_R1110_U176 = ~new_P3_U3064 | ~new_P3_U3903;
  assign new_P3_R1110_U177 = ~new_P3_R1110_U61;
  assign new_P3_R1110_U178 = new_P3_U3066 | new_P3_U3404;
  assign new_P3_R1110_U179 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1110_U180 = new_P3_U3398 | new_P3_U3063;
  assign new_P3_R1110_U181 = new_P3_U3395 | new_P3_U3067;
  assign new_P3_R1110_U182 = ~new_P3_R1110_U31;
  assign new_P3_R1110_U183 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1110_U184 = ~new_P3_R1110_U42;
  assign new_P3_R1110_U185 = ~new_P3_R1110_U43;
  assign new_P3_R1110_U186 = ~new_P3_R1110_U42 | ~new_P3_R1110_U43;
  assign new_P3_R1110_U187 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1110_U188 = ~new_P3_R1110_U186 | ~new_P3_R1110_U181;
  assign new_P3_R1110_U189 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1110_U190 = ~new_P3_R1110_U115 | ~new_P3_R1110_U188;
  assign new_P3_R1110_U191 = ~new_P3_R1110_U35 | ~new_P3_R1110_U34;
  assign new_P3_R1110_U192 = ~new_P3_U3066 | ~new_P3_R1110_U191;
  assign new_P3_R1110_U193 = ~new_P3_R1110_U116 | ~new_P3_R1110_U190;
  assign new_P3_R1110_U194 = ~new_P3_U3404 | ~new_P3_R1110_U170;
  assign new_P3_R1110_U195 = ~new_P3_R1110_U41;
  assign new_P3_R1110_U196 = new_P3_U3069 | new_P3_U3410;
  assign new_P3_R1110_U197 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1110_U198 = ~new_P3_R1110_U22;
  assign new_P3_R1110_U199 = ~new_P3_R1110_U23 | ~new_P3_R1110_U22;
  assign new_P3_R1110_U200 = ~new_P3_U3069 | ~new_P3_R1110_U199;
  assign new_P3_R1110_U201 = ~new_P3_U3410 | ~new_P3_R1110_U198;
  assign new_P3_R1110_U202 = ~new_P3_R1110_U5 | ~new_P3_R1110_U41;
  assign new_P3_R1110_U203 = ~new_P3_R1110_U144;
  assign new_P3_R1110_U204 = new_P3_U3413 | new_P3_U3083;
  assign new_P3_R1110_U205 = ~new_P3_R1110_U204 | ~new_P3_R1110_U144;
  assign new_P3_R1110_U206 = ~new_P3_R1110_U40;
  assign new_P3_R1110_U207 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1110_U208 = new_P3_U3407 | new_P3_U3070;
  assign new_P3_R1110_U209 = ~new_P3_R1110_U208 | ~new_P3_R1110_U41;
  assign new_P3_R1110_U210 = ~new_P3_R1110_U119 | ~new_P3_R1110_U209;
  assign new_P3_R1110_U211 = ~new_P3_R1110_U195 | ~new_P3_R1110_U22;
  assign new_P3_R1110_U212 = ~new_P3_U3410 | ~new_P3_U3069;
  assign new_P3_R1110_U213 = ~new_P3_R1110_U120 | ~new_P3_R1110_U211;
  assign new_P3_R1110_U214 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1110_U215 = ~new_P3_R1110_U185 | ~new_P3_R1110_U181;
  assign new_P3_R1110_U216 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1110_U217 = ~new_P3_R1110_U45;
  assign new_P3_R1110_U218 = ~new_P3_R1110_U121 | ~new_P3_R1110_U184;
  assign new_P3_R1110_U219 = ~new_P3_R1110_U45 | ~new_P3_R1110_U180;
  assign new_P3_R1110_U220 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1110_U221 = ~new_P3_R1110_U44;
  assign new_P3_R1110_U222 = new_P3_U3401 | new_P3_U3059;
  assign new_P3_R1110_U223 = ~new_P3_R1110_U222 | ~new_P3_R1110_U44;
  assign new_P3_R1110_U224 = ~new_P3_R1110_U123 | ~new_P3_R1110_U223;
  assign new_P3_R1110_U225 = ~new_P3_R1110_U221 | ~new_P3_R1110_U34;
  assign new_P3_R1110_U226 = ~new_P3_U3404 | ~new_P3_U3066;
  assign new_P3_R1110_U227 = ~new_P3_R1110_U124 | ~new_P3_R1110_U225;
  assign new_P3_R1110_U228 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1110_U229 = ~new_P3_R1110_U184 | ~new_P3_R1110_U181;
  assign new_P3_R1110_U230 = ~new_P3_R1110_U145;
  assign new_P3_R1110_U231 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1110_U232 = ~new_P3_R1110_U42 | ~new_P3_R1110_U43 | ~new_P3_R1110_U401 | ~new_P3_R1110_U400;
  assign new_P3_R1110_U233 = ~new_P3_R1110_U43 | ~new_P3_R1110_U42;
  assign new_P3_R1110_U234 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1110_U235 = ~new_P3_R1110_U125 | ~new_P3_R1110_U233;
  assign new_P3_R1110_U236 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1110_U237 = new_P3_U3061 | new_P3_U3419;
  assign new_P3_R1110_U238 = ~new_P3_R1110_U177 | ~new_P3_R1110_U6;
  assign new_P3_R1110_U239 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1110_U240 = ~new_P3_R1110_U127 | ~new_P3_R1110_U238;
  assign new_P3_R1110_U241 = new_P3_U3419 | new_P3_U3061;
  assign new_P3_R1110_U242 = ~new_P3_R1110_U126 | ~new_P3_R1110_U144;
  assign new_P3_R1110_U243 = ~new_P3_R1110_U241 | ~new_P3_R1110_U240;
  assign new_P3_R1110_U244 = ~new_P3_R1110_U167;
  assign new_P3_R1110_U245 = new_P3_U3079 | new_P3_U3428;
  assign new_P3_R1110_U246 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1110_U247 = ~new_P3_R1110_U174 | ~new_P3_R1110_U7;
  assign new_P3_R1110_U248 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1110_U249 = ~new_P3_R1110_U129 | ~new_P3_R1110_U247;
  assign new_P3_R1110_U250 = new_P3_U3422 | new_P3_U3062;
  assign new_P3_R1110_U251 = new_P3_U3428 | new_P3_U3079;
  assign new_P3_R1110_U252 = ~new_P3_R1110_U128 | ~new_P3_R1110_U167;
  assign new_P3_R1110_U253 = ~new_P3_R1110_U251 | ~new_P3_R1110_U249;
  assign new_P3_R1110_U254 = ~new_P3_R1110_U166;
  assign new_P3_R1110_U255 = new_P3_U3431 | new_P3_U3078;
  assign new_P3_R1110_U256 = ~new_P3_R1110_U255 | ~new_P3_R1110_U166;
  assign new_P3_R1110_U257 = ~new_P3_U3078 | ~new_P3_U3431;
  assign new_P3_R1110_U258 = ~new_P3_R1110_U164;
  assign new_P3_R1110_U259 = new_P3_U3434 | new_P3_U3073;
  assign new_P3_R1110_U260 = ~new_P3_R1110_U259 | ~new_P3_R1110_U164;
  assign new_P3_R1110_U261 = ~new_P3_U3073 | ~new_P3_U3434;
  assign new_P3_R1110_U262 = ~new_P3_R1110_U92;
  assign new_P3_R1110_U263 = new_P3_U3068 | new_P3_U3440;
  assign new_P3_R1110_U264 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1110_U265 = ~new_P3_R1110_U59;
  assign new_P3_R1110_U266 = ~new_P3_R1110_U60 | ~new_P3_R1110_U59;
  assign new_P3_R1110_U267 = ~new_P3_U3068 | ~new_P3_R1110_U266;
  assign new_P3_R1110_U268 = ~new_P3_U3440 | ~new_P3_R1110_U265;
  assign new_P3_R1110_U269 = ~new_P3_R1110_U8 | ~new_P3_R1110_U92;
  assign new_P3_R1110_U270 = ~new_P3_R1110_U162;
  assign new_P3_R1110_U271 = new_P3_U3075 | new_P3_U3907;
  assign new_P3_R1110_U272 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1110_U273 = new_P3_U3074 | new_P3_U3906;
  assign new_P3_R1110_U274 = ~new_P3_R1110_U80;
  assign new_P3_R1110_U275 = ~new_P3_U3907 | ~new_P3_R1110_U274;
  assign new_P3_R1110_U276 = ~new_P3_R1110_U275 | ~new_P3_R1110_U90;
  assign new_P3_R1110_U277 = ~new_P3_R1110_U80 | ~new_P3_R1110_U81;
  assign new_P3_R1110_U278 = ~new_P3_R1110_U277 | ~new_P3_R1110_U276;
  assign new_P3_R1110_U279 = ~new_P3_R1110_U175 | ~new_P3_R1110_U9;
  assign new_P3_R1110_U280 = ~new_P3_U3074 | ~new_P3_U3906;
  assign new_P3_R1110_U281 = ~new_P3_R1110_U278 | ~new_P3_R1110_U279;
  assign new_P3_R1110_U282 = new_P3_U3443 | new_P3_U3081;
  assign new_P3_R1110_U283 = new_P3_U3906 | new_P3_U3074;
  assign new_P3_R1110_U284 = ~new_P3_R1110_U162 | ~new_P3_R1110_U131;
  assign new_P3_R1110_U285 = ~new_P3_R1110_U283 | ~new_P3_R1110_U281;
  assign new_P3_R1110_U286 = ~new_P3_R1110_U159;
  assign new_P3_R1110_U287 = new_P3_U3905 | new_P3_U3060;
  assign new_P3_R1110_U288 = ~new_P3_R1110_U287 | ~new_P3_R1110_U159;
  assign new_P3_R1110_U289 = ~new_P3_U3060 | ~new_P3_U3905;
  assign new_P3_R1110_U290 = ~new_P3_R1110_U157;
  assign new_P3_R1110_U291 = new_P3_U3904 | new_P3_U3065;
  assign new_P3_R1110_U292 = ~new_P3_R1110_U291 | ~new_P3_R1110_U157;
  assign new_P3_R1110_U293 = ~new_P3_U3065 | ~new_P3_U3904;
  assign new_P3_R1110_U294 = ~new_P3_R1110_U155;
  assign new_P3_R1110_U295 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1110_U296 = ~new_P3_R1110_U176 | ~new_P3_R1110_U173;
  assign new_P3_R1110_U297 = ~new_P3_R1110_U86;
  assign new_P3_R1110_U298 = new_P3_U3903 | new_P3_U3064;
  assign new_P3_R1110_U299 = ~new_P3_R1110_U168 | ~new_P3_R1110_U155 | ~new_P3_R1110_U298;
  assign new_P3_R1110_U300 = ~new_P3_R1110_U153;
  assign new_P3_R1110_U301 = new_P3_U3900 | new_P3_U3052;
  assign new_P3_R1110_U302 = ~new_P3_U3052 | ~new_P3_U3900;
  assign new_P3_R1110_U303 = ~new_P3_R1110_U151;
  assign new_P3_R1110_U304 = ~new_P3_U3899 | ~new_P3_R1110_U151;
  assign new_P3_R1110_U305 = ~new_P3_R1110_U149;
  assign new_P3_R1110_U306 = ~new_P3_R1110_U298 | ~new_P3_R1110_U155;
  assign new_P3_R1110_U307 = ~new_P3_R1110_U89;
  assign new_P3_R1110_U308 = new_P3_U3902 | new_P3_U3057;
  assign new_P3_R1110_U309 = ~new_P3_R1110_U308 | ~new_P3_R1110_U89;
  assign new_P3_R1110_U310 = ~new_P3_R1110_U154 | ~new_P3_R1110_U309 | ~new_P3_R1110_U173;
  assign new_P3_R1110_U311 = ~new_P3_R1110_U307 | ~new_P3_R1110_U173;
  assign new_P3_R1110_U312 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1110_U313 = ~new_P3_R1110_U168 | ~new_P3_R1110_U311 | ~new_P3_R1110_U312;
  assign new_P3_R1110_U314 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1110_U315 = ~new_P3_R1110_U282 | ~new_P3_R1110_U162;
  assign new_P3_R1110_U316 = ~new_P3_R1110_U91;
  assign new_P3_R1110_U317 = ~new_P3_R1110_U9 | ~new_P3_R1110_U91;
  assign new_P3_R1110_U318 = ~new_P3_R1110_U135 | ~new_P3_R1110_U317;
  assign new_P3_R1110_U319 = ~new_P3_R1110_U317 | ~new_P3_R1110_U278;
  assign new_P3_R1110_U320 = ~new_P3_R1110_U453 | ~new_P3_R1110_U319;
  assign new_P3_R1110_U321 = new_P3_U3445 | new_P3_U3080;
  assign new_P3_R1110_U322 = ~new_P3_R1110_U321 | ~new_P3_R1110_U91;
  assign new_P3_R1110_U323 = ~new_P3_R1110_U136 | ~new_P3_R1110_U322;
  assign new_P3_R1110_U324 = ~new_P3_R1110_U316 | ~new_P3_R1110_U80;
  assign new_P3_R1110_U325 = ~new_P3_U3075 | ~new_P3_U3907;
  assign new_P3_R1110_U326 = ~new_P3_R1110_U137 | ~new_P3_R1110_U324;
  assign new_P3_R1110_U327 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1110_U328 = ~new_P3_R1110_U161;
  assign new_P3_R1110_U329 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1110_U330 = new_P3_U3437 | new_P3_U3072;
  assign new_P3_R1110_U331 = ~new_P3_R1110_U330 | ~new_P3_R1110_U92;
  assign new_P3_R1110_U332 = ~new_P3_R1110_U138 | ~new_P3_R1110_U331;
  assign new_P3_R1110_U333 = ~new_P3_R1110_U262 | ~new_P3_R1110_U59;
  assign new_P3_R1110_U334 = ~new_P3_U3440 | ~new_P3_U3068;
  assign new_P3_R1110_U335 = ~new_P3_R1110_U139 | ~new_P3_R1110_U333;
  assign new_P3_R1110_U336 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1110_U337 = ~new_P3_R1110_U250 | ~new_P3_R1110_U167;
  assign new_P3_R1110_U338 = ~new_P3_R1110_U93;
  assign new_P3_R1110_U339 = new_P3_U3425 | new_P3_U3071;
  assign new_P3_R1110_U340 = ~new_P3_R1110_U339 | ~new_P3_R1110_U93;
  assign new_P3_R1110_U341 = ~new_P3_R1110_U140 | ~new_P3_R1110_U340;
  assign new_P3_R1110_U342 = ~new_P3_R1110_U338 | ~new_P3_R1110_U172;
  assign new_P3_R1110_U343 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1110_U344 = ~new_P3_R1110_U141 | ~new_P3_R1110_U342;
  assign new_P3_R1110_U345 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1110_U346 = new_P3_U3416 | new_P3_U3082;
  assign new_P3_R1110_U347 = ~new_P3_R1110_U346 | ~new_P3_R1110_U40;
  assign new_P3_R1110_U348 = ~new_P3_R1110_U142 | ~new_P3_R1110_U347;
  assign new_P3_R1110_U349 = ~new_P3_R1110_U206 | ~new_P3_R1110_U171;
  assign new_P3_R1110_U350 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1110_U351 = ~new_P3_R1110_U143 | ~new_P3_R1110_U349;
  assign new_P3_R1110_U352 = ~new_P3_R1110_U207 | ~new_P3_R1110_U171;
  assign new_P3_R1110_U353 = ~new_P3_R1110_U204 | ~new_P3_R1110_U61;
  assign new_P3_R1110_U354 = ~new_P3_R1110_U214 | ~new_P3_R1110_U22;
  assign new_P3_R1110_U355 = ~new_P3_R1110_U228 | ~new_P3_R1110_U34;
  assign new_P3_R1110_U356 = ~new_P3_R1110_U231 | ~new_P3_R1110_U180;
  assign new_P3_R1110_U357 = ~new_P3_R1110_U314 | ~new_P3_R1110_U173;
  assign new_P3_R1110_U358 = ~new_P3_R1110_U298 | ~new_P3_R1110_U176;
  assign new_P3_R1110_U359 = ~new_P3_R1110_U329 | ~new_P3_R1110_U80;
  assign new_P3_R1110_U360 = ~new_P3_R1110_U282 | ~new_P3_R1110_U77;
  assign new_P3_R1110_U361 = ~new_P3_R1110_U336 | ~new_P3_R1110_U59;
  assign new_P3_R1110_U362 = ~new_P3_R1110_U345 | ~new_P3_R1110_U172;
  assign new_P3_R1110_U363 = ~new_P3_R1110_U250 | ~new_P3_R1110_U68;
  assign new_P3_R1110_U364 = ~new_P3_U3899 | ~new_P3_U3053;
  assign new_P3_R1110_U365 = ~new_P3_R1110_U296 | ~new_P3_R1110_U168;
  assign new_P3_R1110_U366 = ~new_P3_U3056 | ~new_P3_R1110_U295;
  assign new_P3_R1110_U367 = ~new_P3_U3901 | ~new_P3_R1110_U295;
  assign new_P3_R1110_U368 = ~new_P3_R1110_U301 | ~new_P3_R1110_U296 | ~new_P3_R1110_U168;
  assign new_P3_R1110_U369 = ~new_P3_R1110_U133 | ~new_P3_R1110_U155 | ~new_P3_R1110_U168;
  assign new_P3_R1110_U370 = ~new_P3_R1110_U297 | ~new_P3_R1110_U301;
  assign new_P3_R1110_U371 = ~new_P3_U3082 | ~new_P3_R1110_U39;
  assign new_P3_R1110_U372 = ~new_P3_U3416 | ~new_P3_R1110_U38;
  assign new_P3_R1110_U373 = ~new_P3_R1110_U372 | ~new_P3_R1110_U371;
  assign new_P3_R1110_U374 = ~new_P3_R1110_U352 | ~new_P3_R1110_U40;
  assign new_P3_R1110_U375 = ~new_P3_R1110_U373 | ~new_P3_R1110_U206;
  assign new_P3_R1110_U376 = ~new_P3_U3083 | ~new_P3_R1110_U36;
  assign new_P3_R1110_U377 = ~new_P3_U3413 | ~new_P3_R1110_U37;
  assign new_P3_R1110_U378 = ~new_P3_R1110_U377 | ~new_P3_R1110_U376;
  assign new_P3_R1110_U379 = ~new_P3_R1110_U353 | ~new_P3_R1110_U144;
  assign new_P3_R1110_U380 = ~new_P3_R1110_U203 | ~new_P3_R1110_U378;
  assign new_P3_R1110_U381 = ~new_P3_U3069 | ~new_P3_R1110_U23;
  assign new_P3_R1110_U382 = ~new_P3_U3410 | ~new_P3_R1110_U21;
  assign new_P3_R1110_U383 = ~new_P3_U3070 | ~new_P3_R1110_U19;
  assign new_P3_R1110_U384 = ~new_P3_U3407 | ~new_P3_R1110_U20;
  assign new_P3_R1110_U385 = ~new_P3_R1110_U384 | ~new_P3_R1110_U383;
  assign new_P3_R1110_U386 = ~new_P3_R1110_U354 | ~new_P3_R1110_U41;
  assign new_P3_R1110_U387 = ~new_P3_R1110_U385 | ~new_P3_R1110_U195;
  assign new_P3_R1110_U388 = ~new_P3_U3066 | ~new_P3_R1110_U35;
  assign new_P3_R1110_U389 = ~new_P3_U3404 | ~new_P3_R1110_U26;
  assign new_P3_R1110_U390 = ~new_P3_U3059 | ~new_P3_R1110_U24;
  assign new_P3_R1110_U391 = ~new_P3_U3401 | ~new_P3_R1110_U25;
  assign new_P3_R1110_U392 = ~new_P3_R1110_U391 | ~new_P3_R1110_U390;
  assign new_P3_R1110_U393 = ~new_P3_R1110_U355 | ~new_P3_R1110_U44;
  assign new_P3_R1110_U394 = ~new_P3_R1110_U392 | ~new_P3_R1110_U221;
  assign new_P3_R1110_U395 = ~new_P3_U3063 | ~new_P3_R1110_U32;
  assign new_P3_R1110_U396 = ~new_P3_U3398 | ~new_P3_R1110_U33;
  assign new_P3_R1110_U397 = ~new_P3_R1110_U396 | ~new_P3_R1110_U395;
  assign new_P3_R1110_U398 = ~new_P3_R1110_U356 | ~new_P3_R1110_U145;
  assign new_P3_R1110_U399 = ~new_P3_R1110_U230 | ~new_P3_R1110_U397;
  assign new_P3_R1110_U400 = ~new_P3_U3067 | ~new_P3_R1110_U27;
  assign new_P3_R1110_U401 = ~new_P3_U3395 | ~new_P3_R1110_U28;
  assign new_P3_R1110_U402 = ~new_P3_U3054 | ~new_P3_R1110_U147;
  assign new_P3_R1110_U403 = ~new_P3_U3908 | ~new_P3_R1110_U146;
  assign new_P3_R1110_U404 = ~new_P3_U3054 | ~new_P3_R1110_U147;
  assign new_P3_R1110_U405 = ~new_P3_U3908 | ~new_P3_R1110_U146;
  assign new_P3_R1110_U406 = ~new_P3_R1110_U405 | ~new_P3_R1110_U404;
  assign new_P3_R1110_U407 = ~new_P3_R1110_U148 | ~new_P3_R1110_U149;
  assign new_P3_R1110_U408 = ~new_P3_R1110_U305 | ~new_P3_R1110_U406;
  assign new_P3_R1110_U409 = ~new_P3_U3053 | ~new_P3_R1110_U88;
  assign new_P3_R1110_U410 = ~new_P3_U3899 | ~new_P3_R1110_U87;
  assign new_P3_R1110_U411 = ~new_P3_U3053 | ~new_P3_R1110_U88;
  assign new_P3_R1110_U412 = ~new_P3_U3899 | ~new_P3_R1110_U87;
  assign new_P3_R1110_U413 = ~new_P3_R1110_U412 | ~new_P3_R1110_U411;
  assign new_P3_R1110_U414 = ~new_P3_R1110_U150 | ~new_P3_R1110_U151;
  assign new_P3_R1110_U415 = ~new_P3_R1110_U303 | ~new_P3_R1110_U413;
  assign new_P3_R1110_U416 = ~new_P3_U3052 | ~new_P3_R1110_U46;
  assign new_P3_R1110_U417 = ~new_P3_U3900 | ~new_P3_R1110_U47;
  assign new_P3_R1110_U418 = ~new_P3_U3052 | ~new_P3_R1110_U46;
  assign new_P3_R1110_U419 = ~new_P3_U3900 | ~new_P3_R1110_U47;
  assign new_P3_R1110_U420 = ~new_P3_R1110_U419 | ~new_P3_R1110_U418;
  assign new_P3_R1110_U421 = ~new_P3_R1110_U152 | ~new_P3_R1110_U153;
  assign new_P3_R1110_U422 = ~new_P3_R1110_U300 | ~new_P3_R1110_U420;
  assign new_P3_R1110_U423 = ~new_P3_U3056 | ~new_P3_R1110_U49;
  assign new_P3_R1110_U424 = ~new_P3_U3901 | ~new_P3_R1110_U48;
  assign new_P3_R1110_U425 = ~new_P3_U3057 | ~new_P3_R1110_U50;
  assign new_P3_R1110_U426 = ~new_P3_U3902 | ~new_P3_R1110_U51;
  assign new_P3_R1110_U427 = ~new_P3_R1110_U426 | ~new_P3_R1110_U425;
  assign new_P3_R1110_U428 = ~new_P3_R1110_U357 | ~new_P3_R1110_U89;
  assign new_P3_R1110_U429 = ~new_P3_R1110_U427 | ~new_P3_R1110_U307;
  assign new_P3_R1110_U430 = ~new_P3_U3064 | ~new_P3_R1110_U52;
  assign new_P3_R1110_U431 = ~new_P3_U3903 | ~new_P3_R1110_U53;
  assign new_P3_R1110_U432 = ~new_P3_R1110_U431 | ~new_P3_R1110_U430;
  assign new_P3_R1110_U433 = ~new_P3_R1110_U358 | ~new_P3_R1110_U155;
  assign new_P3_R1110_U434 = ~new_P3_R1110_U294 | ~new_P3_R1110_U432;
  assign new_P3_R1110_U435 = ~new_P3_U3065 | ~new_P3_R1110_U84;
  assign new_P3_R1110_U436 = ~new_P3_U3904 | ~new_P3_R1110_U85;
  assign new_P3_R1110_U437 = ~new_P3_U3065 | ~new_P3_R1110_U84;
  assign new_P3_R1110_U438 = ~new_P3_U3904 | ~new_P3_R1110_U85;
  assign new_P3_R1110_U439 = ~new_P3_R1110_U438 | ~new_P3_R1110_U437;
  assign new_P3_R1110_U440 = ~new_P3_R1110_U156 | ~new_P3_R1110_U157;
  assign new_P3_R1110_U441 = ~new_P3_R1110_U290 | ~new_P3_R1110_U439;
  assign new_P3_R1110_U442 = ~new_P3_U3060 | ~new_P3_R1110_U82;
  assign new_P3_R1110_U443 = ~new_P3_U3905 | ~new_P3_R1110_U83;
  assign new_P3_R1110_U444 = ~new_P3_U3060 | ~new_P3_R1110_U82;
  assign new_P3_R1110_U445 = ~new_P3_U3905 | ~new_P3_R1110_U83;
  assign new_P3_R1110_U446 = ~new_P3_R1110_U445 | ~new_P3_R1110_U444;
  assign new_P3_R1110_U447 = ~new_P3_R1110_U158 | ~new_P3_R1110_U159;
  assign new_P3_R1110_U448 = ~new_P3_R1110_U286 | ~new_P3_R1110_U446;
  assign new_P3_R1110_U449 = ~new_P3_U3074 | ~new_P3_R1110_U54;
  assign new_P3_R1110_U450 = ~new_P3_U3906 | ~new_P3_R1110_U55;
  assign new_P3_R1110_U451 = ~new_P3_U3074 | ~new_P3_R1110_U54;
  assign new_P3_R1110_U452 = ~new_P3_U3906 | ~new_P3_R1110_U55;
  assign new_P3_R1110_U453 = ~new_P3_R1110_U452 | ~new_P3_R1110_U451;
  assign new_P3_R1110_U454 = ~new_P3_U3075 | ~new_P3_R1110_U81;
  assign new_P3_R1110_U455 = ~new_P3_U3907 | ~new_P3_R1110_U90;
  assign new_P3_R1110_U456 = ~new_P3_R1110_U182 | ~new_P3_R1110_U161;
  assign new_P3_R1110_U457 = ~new_P3_R1110_U328 | ~new_P3_R1110_U31;
  assign new_P3_R1110_U458 = ~new_P3_U3080 | ~new_P3_R1110_U78;
  assign new_P3_R1110_U459 = ~new_P3_U3445 | ~new_P3_R1110_U79;
  assign new_P3_R1110_U460 = ~new_P3_R1110_U459 | ~new_P3_R1110_U458;
  assign new_P3_R1110_U461 = ~new_P3_R1110_U359 | ~new_P3_R1110_U91;
  assign new_P3_R1110_U462 = ~new_P3_R1110_U460 | ~new_P3_R1110_U316;
  assign new_P3_R1110_U463 = ~new_P3_U3081 | ~new_P3_R1110_U75;
  assign new_P3_R1110_U464 = ~new_P3_U3443 | ~new_P3_R1110_U76;
  assign new_P3_R1110_U465 = ~new_P3_R1110_U464 | ~new_P3_R1110_U463;
  assign new_P3_R1110_U466 = ~new_P3_R1110_U360 | ~new_P3_R1110_U162;
  assign new_P3_R1110_U467 = ~new_P3_R1110_U270 | ~new_P3_R1110_U465;
  assign new_P3_R1110_U468 = ~new_P3_U3068 | ~new_P3_R1110_U60;
  assign new_P3_R1110_U469 = ~new_P3_U3440 | ~new_P3_R1110_U58;
  assign new_P3_R1110_U470 = ~new_P3_U3072 | ~new_P3_R1110_U56;
  assign new_P3_R1110_U471 = ~new_P3_U3437 | ~new_P3_R1110_U57;
  assign new_P3_R1110_U472 = ~new_P3_R1110_U471 | ~new_P3_R1110_U470;
  assign new_P3_R1110_U473 = ~new_P3_R1110_U361 | ~new_P3_R1110_U92;
  assign new_P3_R1110_U474 = ~new_P3_R1110_U472 | ~new_P3_R1110_U262;
  assign new_P3_R1110_U475 = ~new_P3_U3073 | ~new_P3_R1110_U73;
  assign new_P3_R1110_U476 = ~new_P3_U3434 | ~new_P3_R1110_U74;
  assign new_P3_R1110_U477 = ~new_P3_U3073 | ~new_P3_R1110_U73;
  assign new_P3_R1110_U478 = ~new_P3_U3434 | ~new_P3_R1110_U74;
  assign new_P3_R1110_U479 = ~new_P3_R1110_U478 | ~new_P3_R1110_U477;
  assign new_P3_R1110_U480 = ~new_P3_R1110_U163 | ~new_P3_R1110_U164;
  assign new_P3_R1110_U481 = ~new_P3_R1110_U258 | ~new_P3_R1110_U479;
  assign new_P3_R1110_U482 = ~new_P3_U3078 | ~new_P3_R1110_U71;
  assign new_P3_R1110_U483 = ~new_P3_U3431 | ~new_P3_R1110_U72;
  assign new_P3_R1110_U484 = ~new_P3_U3078 | ~new_P3_R1110_U71;
  assign new_P3_R1110_U485 = ~new_P3_U3431 | ~new_P3_R1110_U72;
  assign new_P3_R1110_U486 = ~new_P3_R1110_U485 | ~new_P3_R1110_U484;
  assign new_P3_R1110_U487 = ~new_P3_R1110_U165 | ~new_P3_R1110_U166;
  assign new_P3_R1110_U488 = ~new_P3_R1110_U254 | ~new_P3_R1110_U486;
  assign new_P3_R1110_U489 = ~new_P3_U3079 | ~new_P3_R1110_U69;
  assign new_P3_R1110_U490 = ~new_P3_U3428 | ~new_P3_R1110_U70;
  assign new_P3_R1110_U491 = ~new_P3_U3071 | ~new_P3_R1110_U64;
  assign new_P3_R1110_U492 = ~new_P3_U3425 | ~new_P3_R1110_U65;
  assign new_P3_R1110_U493 = ~new_P3_R1110_U492 | ~new_P3_R1110_U491;
  assign new_P3_R1110_U494 = ~new_P3_R1110_U362 | ~new_P3_R1110_U93;
  assign new_P3_R1110_U495 = ~new_P3_R1110_U493 | ~new_P3_R1110_U338;
  assign new_P3_R1110_U496 = ~new_P3_U3062 | ~new_P3_R1110_U66;
  assign new_P3_R1110_U497 = ~new_P3_U3422 | ~new_P3_R1110_U67;
  assign new_P3_R1110_U498 = ~new_P3_R1110_U497 | ~new_P3_R1110_U496;
  assign new_P3_R1110_U499 = ~new_P3_R1110_U363 | ~new_P3_R1110_U167;
  assign new_P3_R1110_U500 = ~new_P3_R1110_U244 | ~new_P3_R1110_U498;
  assign new_P3_R1110_U501 = ~new_P3_U3061 | ~new_P3_R1110_U62;
  assign new_P3_R1110_U502 = ~new_P3_U3419 | ~new_P3_R1110_U63;
  assign new_P3_R1110_U503 = ~new_P3_U3076 | ~new_P3_R1110_U29;
  assign new_P3_R1110_U504 = ~new_P3_U3387 | ~new_P3_R1110_U30;
  assign new_P3_R1297_U6 = new_P3_U3058 & new_P3_R1297_U7;
  assign new_P3_R1297_U7 = ~new_P3_U3055;
  assign new_P3_R1077_U4 = new_P3_R1077_U179 & new_P3_R1077_U178;
  assign new_P3_R1077_U5 = new_P3_R1077_U197 & new_P3_R1077_U196;
  assign new_P3_R1077_U6 = new_P3_R1077_U237 & new_P3_R1077_U236;
  assign new_P3_R1077_U7 = new_P3_R1077_U246 & new_P3_R1077_U245;
  assign new_P3_R1077_U8 = new_P3_R1077_U264 & new_P3_R1077_U263;
  assign new_P3_R1077_U9 = new_P3_R1077_U272 & new_P3_R1077_U271;
  assign new_P3_R1077_U10 = new_P3_R1077_U351 & new_P3_R1077_U348;
  assign new_P3_R1077_U11 = new_P3_R1077_U344 & new_P3_R1077_U341;
  assign new_P3_R1077_U12 = new_P3_R1077_U335 & new_P3_R1077_U332;
  assign new_P3_R1077_U13 = new_P3_R1077_U326 & new_P3_R1077_U323;
  assign new_P3_R1077_U14 = new_P3_R1077_U320 & new_P3_R1077_U318;
  assign new_P3_R1077_U15 = new_P3_R1077_U313 & new_P3_R1077_U310;
  assign new_P3_R1077_U16 = new_P3_R1077_U235 & new_P3_R1077_U232;
  assign new_P3_R1077_U17 = new_P3_R1077_U227 & new_P3_R1077_U224;
  assign new_P3_R1077_U18 = new_P3_R1077_U213 & new_P3_R1077_U210;
  assign new_P3_R1077_U19 = ~new_P3_U3407;
  assign new_P3_R1077_U20 = ~new_P3_U3070;
  assign new_P3_R1077_U21 = ~new_P3_U3069;
  assign new_P3_R1077_U22 = ~new_P3_U3070 | ~new_P3_U3407;
  assign new_P3_R1077_U23 = ~new_P3_U3410;
  assign new_P3_R1077_U24 = ~new_P3_U3401;
  assign new_P3_R1077_U25 = ~new_P3_U3059;
  assign new_P3_R1077_U26 = ~new_P3_U3066;
  assign new_P3_R1077_U27 = ~new_P3_U3395;
  assign new_P3_R1077_U28 = ~new_P3_U3067;
  assign new_P3_R1077_U29 = ~new_P3_U3387;
  assign new_P3_R1077_U30 = ~new_P3_U3076;
  assign new_P3_R1077_U31 = ~new_P3_U3076 | ~new_P3_U3387;
  assign new_P3_R1077_U32 = ~new_P3_U3398;
  assign new_P3_R1077_U33 = ~new_P3_U3063;
  assign new_P3_R1077_U34 = ~new_P3_U3059 | ~new_P3_U3401;
  assign new_P3_R1077_U35 = ~new_P3_U3404;
  assign new_P3_R1077_U36 = ~new_P3_U3413;
  assign new_P3_R1077_U37 = ~new_P3_U3083;
  assign new_P3_R1077_U38 = ~new_P3_U3082;
  assign new_P3_R1077_U39 = ~new_P3_U3416;
  assign new_P3_R1077_U40 = ~new_P3_R1077_U61 | ~new_P3_R1077_U205;
  assign new_P3_R1077_U41 = ~new_P3_R1077_U117 | ~new_P3_R1077_U193;
  assign new_P3_R1077_U42 = ~new_P3_R1077_U182 | ~new_P3_R1077_U183;
  assign new_P3_R1077_U43 = ~new_P3_U3392 | ~new_P3_U3077;
  assign new_P3_R1077_U44 = ~new_P3_R1077_U122 | ~new_P3_R1077_U219;
  assign new_P3_R1077_U45 = ~new_P3_R1077_U216 | ~new_P3_R1077_U215;
  assign new_P3_R1077_U46 = ~new_P3_U3900;
  assign new_P3_R1077_U47 = ~new_P3_U3052;
  assign new_P3_R1077_U48 = ~new_P3_U3056;
  assign new_P3_R1077_U49 = ~new_P3_U3901;
  assign new_P3_R1077_U50 = ~new_P3_U3902;
  assign new_P3_R1077_U51 = ~new_P3_U3057;
  assign new_P3_R1077_U52 = ~new_P3_U3903;
  assign new_P3_R1077_U53 = ~new_P3_U3064;
  assign new_P3_R1077_U54 = ~new_P3_U3906;
  assign new_P3_R1077_U55 = ~new_P3_U3074;
  assign new_P3_R1077_U56 = ~new_P3_U3437;
  assign new_P3_R1077_U57 = ~new_P3_U3072;
  assign new_P3_R1077_U58 = ~new_P3_U3068;
  assign new_P3_R1077_U59 = ~new_P3_U3072 | ~new_P3_U3437;
  assign new_P3_R1077_U60 = ~new_P3_U3440;
  assign new_P3_R1077_U61 = ~new_P3_U3083 | ~new_P3_U3413;
  assign new_P3_R1077_U62 = ~new_P3_U3419;
  assign new_P3_R1077_U63 = ~new_P3_U3061;
  assign new_P3_R1077_U64 = ~new_P3_U3425;
  assign new_P3_R1077_U65 = ~new_P3_U3071;
  assign new_P3_R1077_U66 = ~new_P3_U3422;
  assign new_P3_R1077_U67 = ~new_P3_U3062;
  assign new_P3_R1077_U68 = ~new_P3_U3062 | ~new_P3_U3422;
  assign new_P3_R1077_U69 = ~new_P3_U3428;
  assign new_P3_R1077_U70 = ~new_P3_U3079;
  assign new_P3_R1077_U71 = ~new_P3_U3431;
  assign new_P3_R1077_U72 = ~new_P3_U3078;
  assign new_P3_R1077_U73 = ~new_P3_U3434;
  assign new_P3_R1077_U74 = ~new_P3_U3073;
  assign new_P3_R1077_U75 = ~new_P3_U3443;
  assign new_P3_R1077_U76 = ~new_P3_U3081;
  assign new_P3_R1077_U77 = ~new_P3_U3081 | ~new_P3_U3443;
  assign new_P3_R1077_U78 = ~new_P3_U3445;
  assign new_P3_R1077_U79 = ~new_P3_U3080;
  assign new_P3_R1077_U80 = ~new_P3_U3080 | ~new_P3_U3445;
  assign new_P3_R1077_U81 = ~new_P3_U3907;
  assign new_P3_R1077_U82 = ~new_P3_U3905;
  assign new_P3_R1077_U83 = ~new_P3_U3060;
  assign new_P3_R1077_U84 = ~new_P3_U3904;
  assign new_P3_R1077_U85 = ~new_P3_U3065;
  assign new_P3_R1077_U86 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1077_U87 = ~new_P3_U3053;
  assign new_P3_R1077_U88 = ~new_P3_U3899;
  assign new_P3_R1077_U89 = ~new_P3_R1077_U306 | ~new_P3_R1077_U176;
  assign new_P3_R1077_U90 = ~new_P3_U3075;
  assign new_P3_R1077_U91 = ~new_P3_R1077_U77 | ~new_P3_R1077_U315;
  assign new_P3_R1077_U92 = ~new_P3_R1077_U261 | ~new_P3_R1077_U260;
  assign new_P3_R1077_U93 = ~new_P3_R1077_U68 | ~new_P3_R1077_U337;
  assign new_P3_R1077_U94 = ~new_P3_R1077_U457 | ~new_P3_R1077_U456;
  assign new_P3_R1077_U95 = ~new_P3_R1077_U504 | ~new_P3_R1077_U503;
  assign new_P3_R1077_U96 = ~new_P3_R1077_U375 | ~new_P3_R1077_U374;
  assign new_P3_R1077_U97 = ~new_P3_R1077_U380 | ~new_P3_R1077_U379;
  assign new_P3_R1077_U98 = ~new_P3_R1077_U387 | ~new_P3_R1077_U386;
  assign new_P3_R1077_U99 = ~new_P3_R1077_U394 | ~new_P3_R1077_U393;
  assign new_P3_R1077_U100 = ~new_P3_R1077_U399 | ~new_P3_R1077_U398;
  assign new_P3_R1077_U101 = ~new_P3_R1077_U408 | ~new_P3_R1077_U407;
  assign new_P3_R1077_U102 = ~new_P3_R1077_U415 | ~new_P3_R1077_U414;
  assign new_P3_R1077_U103 = ~new_P3_R1077_U422 | ~new_P3_R1077_U421;
  assign new_P3_R1077_U104 = ~new_P3_R1077_U429 | ~new_P3_R1077_U428;
  assign new_P3_R1077_U105 = ~new_P3_R1077_U434 | ~new_P3_R1077_U433;
  assign new_P3_R1077_U106 = ~new_P3_R1077_U441 | ~new_P3_R1077_U440;
  assign new_P3_R1077_U107 = ~new_P3_R1077_U448 | ~new_P3_R1077_U447;
  assign new_P3_R1077_U108 = ~new_P3_R1077_U462 | ~new_P3_R1077_U461;
  assign new_P3_R1077_U109 = ~new_P3_R1077_U467 | ~new_P3_R1077_U466;
  assign new_P3_R1077_U110 = ~new_P3_R1077_U474 | ~new_P3_R1077_U473;
  assign new_P3_R1077_U111 = ~new_P3_R1077_U481 | ~new_P3_R1077_U480;
  assign new_P3_R1077_U112 = ~new_P3_R1077_U488 | ~new_P3_R1077_U487;
  assign new_P3_R1077_U113 = ~new_P3_R1077_U495 | ~new_P3_R1077_U494;
  assign new_P3_R1077_U114 = ~new_P3_R1077_U500 | ~new_P3_R1077_U499;
  assign new_P3_R1077_U115 = new_P3_R1077_U189 & new_P3_R1077_U187;
  assign new_P3_R1077_U116 = new_P3_R1077_U4 & new_P3_R1077_U180;
  assign new_P3_R1077_U117 = new_P3_R1077_U194 & new_P3_R1077_U192;
  assign new_P3_R1077_U118 = new_P3_R1077_U201 & new_P3_R1077_U200;
  assign new_P3_R1077_U119 = new_P3_R1077_U22 & new_P3_R1077_U382 & new_P3_R1077_U381;
  assign new_P3_R1077_U120 = new_P3_R1077_U212 & new_P3_R1077_U5;
  assign new_P3_R1077_U121 = new_P3_R1077_U181 & new_P3_R1077_U180;
  assign new_P3_R1077_U122 = new_P3_R1077_U220 & new_P3_R1077_U218;
  assign new_P3_R1077_U123 = new_P3_R1077_U34 & new_P3_R1077_U389 & new_P3_R1077_U388;
  assign new_P3_R1077_U124 = new_P3_R1077_U226 & new_P3_R1077_U4;
  assign new_P3_R1077_U125 = new_P3_R1077_U234 & new_P3_R1077_U181;
  assign new_P3_R1077_U126 = new_P3_R1077_U204 & new_P3_R1077_U6;
  assign new_P3_R1077_U127 = new_P3_R1077_U239 & new_P3_R1077_U171;
  assign new_P3_R1077_U128 = new_P3_R1077_U250 & new_P3_R1077_U7;
  assign new_P3_R1077_U129 = new_P3_R1077_U248 & new_P3_R1077_U172;
  assign new_P3_R1077_U130 = new_P3_R1077_U268 & new_P3_R1077_U267;
  assign new_P3_R1077_U131 = new_P3_R1077_U273 & new_P3_R1077_U9 & new_P3_R1077_U282;
  assign new_P3_R1077_U132 = new_P3_R1077_U285 & new_P3_R1077_U280;
  assign new_P3_R1077_U133 = new_P3_R1077_U301 & new_P3_R1077_U298;
  assign new_P3_R1077_U134 = new_P3_R1077_U368 & new_P3_R1077_U302;
  assign new_P3_R1077_U135 = new_P3_R1077_U160 & new_P3_R1077_U278;
  assign new_P3_R1077_U136 = new_P3_R1077_U80 & new_P3_R1077_U455 & new_P3_R1077_U454;
  assign new_P3_R1077_U137 = new_P3_R1077_U325 & new_P3_R1077_U9;
  assign new_P3_R1077_U138 = new_P3_R1077_U59 & new_P3_R1077_U469 & new_P3_R1077_U468;
  assign new_P3_R1077_U139 = new_P3_R1077_U334 & new_P3_R1077_U8;
  assign new_P3_R1077_U140 = new_P3_R1077_U172 & new_P3_R1077_U490 & new_P3_R1077_U489;
  assign new_P3_R1077_U141 = new_P3_R1077_U343 & new_P3_R1077_U7;
  assign new_P3_R1077_U142 = new_P3_R1077_U171 & new_P3_R1077_U502 & new_P3_R1077_U501;
  assign new_P3_R1077_U143 = new_P3_R1077_U350 & new_P3_R1077_U6;
  assign new_P3_R1077_U144 = ~new_P3_R1077_U118 | ~new_P3_R1077_U202;
  assign new_P3_R1077_U145 = ~new_P3_R1077_U217 | ~new_P3_R1077_U229;
  assign new_P3_R1077_U146 = ~new_P3_U3054;
  assign new_P3_R1077_U147 = ~new_P3_U3908;
  assign new_P3_R1077_U148 = new_P3_R1077_U403 & new_P3_R1077_U402;
  assign new_P3_R1077_U149 = ~new_P3_R1077_U364 | ~new_P3_R1077_U304 | ~new_P3_R1077_U169;
  assign new_P3_R1077_U150 = new_P3_R1077_U410 & new_P3_R1077_U409;
  assign new_P3_R1077_U151 = ~new_P3_R1077_U134 | ~new_P3_R1077_U370 | ~new_P3_R1077_U369;
  assign new_P3_R1077_U152 = new_P3_R1077_U417 & new_P3_R1077_U416;
  assign new_P3_R1077_U153 = ~new_P3_R1077_U86 | ~new_P3_R1077_U365 | ~new_P3_R1077_U299;
  assign new_P3_R1077_U154 = new_P3_R1077_U424 & new_P3_R1077_U423;
  assign new_P3_R1077_U155 = ~new_P3_R1077_U293 | ~new_P3_R1077_U292;
  assign new_P3_R1077_U156 = new_P3_R1077_U436 & new_P3_R1077_U435;
  assign new_P3_R1077_U157 = ~new_P3_R1077_U289 | ~new_P3_R1077_U288;
  assign new_P3_R1077_U158 = new_P3_R1077_U443 & new_P3_R1077_U442;
  assign new_P3_R1077_U159 = ~new_P3_R1077_U132 | ~new_P3_R1077_U284;
  assign new_P3_R1077_U160 = new_P3_R1077_U450 & new_P3_R1077_U449;
  assign new_P3_R1077_U161 = ~new_P3_R1077_U43 | ~new_P3_R1077_U327;
  assign new_P3_R1077_U162 = ~new_P3_R1077_U130 | ~new_P3_R1077_U269;
  assign new_P3_R1077_U163 = new_P3_R1077_U476 & new_P3_R1077_U475;
  assign new_P3_R1077_U164 = ~new_P3_R1077_U257 | ~new_P3_R1077_U256;
  assign new_P3_R1077_U165 = new_P3_R1077_U483 & new_P3_R1077_U482;
  assign new_P3_R1077_U166 = ~new_P3_R1077_U253 | ~new_P3_R1077_U252;
  assign new_P3_R1077_U167 = ~new_P3_R1077_U243 | ~new_P3_R1077_U242;
  assign new_P3_R1077_U168 = ~new_P3_R1077_U367 | ~new_P3_R1077_U366;
  assign new_P3_R1077_U169 = ~new_P3_U3053 | ~new_P3_R1077_U151;
  assign new_P3_R1077_U170 = ~new_P3_R1077_U34;
  assign new_P3_R1077_U171 = ~new_P3_U3416 | ~new_P3_U3082;
  assign new_P3_R1077_U172 = ~new_P3_U3071 | ~new_P3_U3425;
  assign new_P3_R1077_U173 = ~new_P3_U3057 | ~new_P3_U3902;
  assign new_P3_R1077_U174 = ~new_P3_R1077_U68;
  assign new_P3_R1077_U175 = ~new_P3_R1077_U77;
  assign new_P3_R1077_U176 = ~new_P3_U3064 | ~new_P3_U3903;
  assign new_P3_R1077_U177 = ~new_P3_R1077_U61;
  assign new_P3_R1077_U178 = new_P3_U3066 | new_P3_U3404;
  assign new_P3_R1077_U179 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1077_U180 = new_P3_U3398 | new_P3_U3063;
  assign new_P3_R1077_U181 = new_P3_U3395 | new_P3_U3067;
  assign new_P3_R1077_U182 = ~new_P3_R1077_U31;
  assign new_P3_R1077_U183 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1077_U184 = ~new_P3_R1077_U42;
  assign new_P3_R1077_U185 = ~new_P3_R1077_U43;
  assign new_P3_R1077_U186 = ~new_P3_R1077_U42 | ~new_P3_R1077_U43;
  assign new_P3_R1077_U187 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1077_U188 = ~new_P3_R1077_U186 | ~new_P3_R1077_U181;
  assign new_P3_R1077_U189 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1077_U190 = ~new_P3_R1077_U115 | ~new_P3_R1077_U188;
  assign new_P3_R1077_U191 = ~new_P3_R1077_U35 | ~new_P3_R1077_U34;
  assign new_P3_R1077_U192 = ~new_P3_U3066 | ~new_P3_R1077_U191;
  assign new_P3_R1077_U193 = ~new_P3_R1077_U116 | ~new_P3_R1077_U190;
  assign new_P3_R1077_U194 = ~new_P3_U3404 | ~new_P3_R1077_U170;
  assign new_P3_R1077_U195 = ~new_P3_R1077_U41;
  assign new_P3_R1077_U196 = new_P3_U3069 | new_P3_U3410;
  assign new_P3_R1077_U197 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1077_U198 = ~new_P3_R1077_U22;
  assign new_P3_R1077_U199 = ~new_P3_R1077_U23 | ~new_P3_R1077_U22;
  assign new_P3_R1077_U200 = ~new_P3_U3069 | ~new_P3_R1077_U199;
  assign new_P3_R1077_U201 = ~new_P3_U3410 | ~new_P3_R1077_U198;
  assign new_P3_R1077_U202 = ~new_P3_R1077_U5 | ~new_P3_R1077_U41;
  assign new_P3_R1077_U203 = ~new_P3_R1077_U144;
  assign new_P3_R1077_U204 = new_P3_U3413 | new_P3_U3083;
  assign new_P3_R1077_U205 = ~new_P3_R1077_U204 | ~new_P3_R1077_U144;
  assign new_P3_R1077_U206 = ~new_P3_R1077_U40;
  assign new_P3_R1077_U207 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1077_U208 = new_P3_U3407 | new_P3_U3070;
  assign new_P3_R1077_U209 = ~new_P3_R1077_U208 | ~new_P3_R1077_U41;
  assign new_P3_R1077_U210 = ~new_P3_R1077_U119 | ~new_P3_R1077_U209;
  assign new_P3_R1077_U211 = ~new_P3_R1077_U195 | ~new_P3_R1077_U22;
  assign new_P3_R1077_U212 = ~new_P3_U3410 | ~new_P3_U3069;
  assign new_P3_R1077_U213 = ~new_P3_R1077_U120 | ~new_P3_R1077_U211;
  assign new_P3_R1077_U214 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1077_U215 = ~new_P3_R1077_U185 | ~new_P3_R1077_U181;
  assign new_P3_R1077_U216 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1077_U217 = ~new_P3_R1077_U45;
  assign new_P3_R1077_U218 = ~new_P3_R1077_U121 | ~new_P3_R1077_U184;
  assign new_P3_R1077_U219 = ~new_P3_R1077_U45 | ~new_P3_R1077_U180;
  assign new_P3_R1077_U220 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1077_U221 = ~new_P3_R1077_U44;
  assign new_P3_R1077_U222 = new_P3_U3401 | new_P3_U3059;
  assign new_P3_R1077_U223 = ~new_P3_R1077_U222 | ~new_P3_R1077_U44;
  assign new_P3_R1077_U224 = ~new_P3_R1077_U123 | ~new_P3_R1077_U223;
  assign new_P3_R1077_U225 = ~new_P3_R1077_U221 | ~new_P3_R1077_U34;
  assign new_P3_R1077_U226 = ~new_P3_U3404 | ~new_P3_U3066;
  assign new_P3_R1077_U227 = ~new_P3_R1077_U124 | ~new_P3_R1077_U225;
  assign new_P3_R1077_U228 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1077_U229 = ~new_P3_R1077_U184 | ~new_P3_R1077_U181;
  assign new_P3_R1077_U230 = ~new_P3_R1077_U145;
  assign new_P3_R1077_U231 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1077_U232 = ~new_P3_R1077_U42 | ~new_P3_R1077_U43 | ~new_P3_R1077_U401 | ~new_P3_R1077_U400;
  assign new_P3_R1077_U233 = ~new_P3_R1077_U43 | ~new_P3_R1077_U42;
  assign new_P3_R1077_U234 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1077_U235 = ~new_P3_R1077_U125 | ~new_P3_R1077_U233;
  assign new_P3_R1077_U236 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1077_U237 = new_P3_U3061 | new_P3_U3419;
  assign new_P3_R1077_U238 = ~new_P3_R1077_U177 | ~new_P3_R1077_U6;
  assign new_P3_R1077_U239 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1077_U240 = ~new_P3_R1077_U127 | ~new_P3_R1077_U238;
  assign new_P3_R1077_U241 = new_P3_U3419 | new_P3_U3061;
  assign new_P3_R1077_U242 = ~new_P3_R1077_U126 | ~new_P3_R1077_U144;
  assign new_P3_R1077_U243 = ~new_P3_R1077_U241 | ~new_P3_R1077_U240;
  assign new_P3_R1077_U244 = ~new_P3_R1077_U167;
  assign new_P3_R1077_U245 = new_P3_U3079 | new_P3_U3428;
  assign new_P3_R1077_U246 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1077_U247 = ~new_P3_R1077_U174 | ~new_P3_R1077_U7;
  assign new_P3_R1077_U248 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1077_U249 = ~new_P3_R1077_U129 | ~new_P3_R1077_U247;
  assign new_P3_R1077_U250 = new_P3_U3422 | new_P3_U3062;
  assign new_P3_R1077_U251 = new_P3_U3428 | new_P3_U3079;
  assign new_P3_R1077_U252 = ~new_P3_R1077_U128 | ~new_P3_R1077_U167;
  assign new_P3_R1077_U253 = ~new_P3_R1077_U251 | ~new_P3_R1077_U249;
  assign new_P3_R1077_U254 = ~new_P3_R1077_U166;
  assign new_P3_R1077_U255 = new_P3_U3431 | new_P3_U3078;
  assign new_P3_R1077_U256 = ~new_P3_R1077_U255 | ~new_P3_R1077_U166;
  assign new_P3_R1077_U257 = ~new_P3_U3078 | ~new_P3_U3431;
  assign new_P3_R1077_U258 = ~new_P3_R1077_U164;
  assign new_P3_R1077_U259 = new_P3_U3434 | new_P3_U3073;
  assign new_P3_R1077_U260 = ~new_P3_R1077_U259 | ~new_P3_R1077_U164;
  assign new_P3_R1077_U261 = ~new_P3_U3073 | ~new_P3_U3434;
  assign new_P3_R1077_U262 = ~new_P3_R1077_U92;
  assign new_P3_R1077_U263 = new_P3_U3068 | new_P3_U3440;
  assign new_P3_R1077_U264 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1077_U265 = ~new_P3_R1077_U59;
  assign new_P3_R1077_U266 = ~new_P3_R1077_U60 | ~new_P3_R1077_U59;
  assign new_P3_R1077_U267 = ~new_P3_U3068 | ~new_P3_R1077_U266;
  assign new_P3_R1077_U268 = ~new_P3_U3440 | ~new_P3_R1077_U265;
  assign new_P3_R1077_U269 = ~new_P3_R1077_U8 | ~new_P3_R1077_U92;
  assign new_P3_R1077_U270 = ~new_P3_R1077_U162;
  assign new_P3_R1077_U271 = new_P3_U3075 | new_P3_U3907;
  assign new_P3_R1077_U272 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1077_U273 = new_P3_U3074 | new_P3_U3906;
  assign new_P3_R1077_U274 = ~new_P3_R1077_U80;
  assign new_P3_R1077_U275 = ~new_P3_U3907 | ~new_P3_R1077_U274;
  assign new_P3_R1077_U276 = ~new_P3_R1077_U275 | ~new_P3_R1077_U90;
  assign new_P3_R1077_U277 = ~new_P3_R1077_U80 | ~new_P3_R1077_U81;
  assign new_P3_R1077_U278 = ~new_P3_R1077_U277 | ~new_P3_R1077_U276;
  assign new_P3_R1077_U279 = ~new_P3_R1077_U175 | ~new_P3_R1077_U9;
  assign new_P3_R1077_U280 = ~new_P3_U3074 | ~new_P3_U3906;
  assign new_P3_R1077_U281 = ~new_P3_R1077_U278 | ~new_P3_R1077_U279;
  assign new_P3_R1077_U282 = new_P3_U3443 | new_P3_U3081;
  assign new_P3_R1077_U283 = new_P3_U3906 | new_P3_U3074;
  assign new_P3_R1077_U284 = ~new_P3_R1077_U162 | ~new_P3_R1077_U131;
  assign new_P3_R1077_U285 = ~new_P3_R1077_U283 | ~new_P3_R1077_U281;
  assign new_P3_R1077_U286 = ~new_P3_R1077_U159;
  assign new_P3_R1077_U287 = new_P3_U3905 | new_P3_U3060;
  assign new_P3_R1077_U288 = ~new_P3_R1077_U287 | ~new_P3_R1077_U159;
  assign new_P3_R1077_U289 = ~new_P3_U3060 | ~new_P3_U3905;
  assign new_P3_R1077_U290 = ~new_P3_R1077_U157;
  assign new_P3_R1077_U291 = new_P3_U3904 | new_P3_U3065;
  assign new_P3_R1077_U292 = ~new_P3_R1077_U291 | ~new_P3_R1077_U157;
  assign new_P3_R1077_U293 = ~new_P3_U3065 | ~new_P3_U3904;
  assign new_P3_R1077_U294 = ~new_P3_R1077_U155;
  assign new_P3_R1077_U295 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1077_U296 = ~new_P3_R1077_U176 | ~new_P3_R1077_U173;
  assign new_P3_R1077_U297 = ~new_P3_R1077_U86;
  assign new_P3_R1077_U298 = new_P3_U3903 | new_P3_U3064;
  assign new_P3_R1077_U299 = ~new_P3_R1077_U168 | ~new_P3_R1077_U155 | ~new_P3_R1077_U298;
  assign new_P3_R1077_U300 = ~new_P3_R1077_U153;
  assign new_P3_R1077_U301 = new_P3_U3900 | new_P3_U3052;
  assign new_P3_R1077_U302 = ~new_P3_U3052 | ~new_P3_U3900;
  assign new_P3_R1077_U303 = ~new_P3_R1077_U151;
  assign new_P3_R1077_U304 = ~new_P3_U3899 | ~new_P3_R1077_U151;
  assign new_P3_R1077_U305 = ~new_P3_R1077_U149;
  assign new_P3_R1077_U306 = ~new_P3_R1077_U298 | ~new_P3_R1077_U155;
  assign new_P3_R1077_U307 = ~new_P3_R1077_U89;
  assign new_P3_R1077_U308 = new_P3_U3902 | new_P3_U3057;
  assign new_P3_R1077_U309 = ~new_P3_R1077_U308 | ~new_P3_R1077_U89;
  assign new_P3_R1077_U310 = ~new_P3_R1077_U154 | ~new_P3_R1077_U309 | ~new_P3_R1077_U173;
  assign new_P3_R1077_U311 = ~new_P3_R1077_U307 | ~new_P3_R1077_U173;
  assign new_P3_R1077_U312 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1077_U313 = ~new_P3_R1077_U168 | ~new_P3_R1077_U311 | ~new_P3_R1077_U312;
  assign new_P3_R1077_U314 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1077_U315 = ~new_P3_R1077_U282 | ~new_P3_R1077_U162;
  assign new_P3_R1077_U316 = ~new_P3_R1077_U91;
  assign new_P3_R1077_U317 = ~new_P3_R1077_U9 | ~new_P3_R1077_U91;
  assign new_P3_R1077_U318 = ~new_P3_R1077_U135 | ~new_P3_R1077_U317;
  assign new_P3_R1077_U319 = ~new_P3_R1077_U317 | ~new_P3_R1077_U278;
  assign new_P3_R1077_U320 = ~new_P3_R1077_U453 | ~new_P3_R1077_U319;
  assign new_P3_R1077_U321 = new_P3_U3445 | new_P3_U3080;
  assign new_P3_R1077_U322 = ~new_P3_R1077_U321 | ~new_P3_R1077_U91;
  assign new_P3_R1077_U323 = ~new_P3_R1077_U136 | ~new_P3_R1077_U322;
  assign new_P3_R1077_U324 = ~new_P3_R1077_U316 | ~new_P3_R1077_U80;
  assign new_P3_R1077_U325 = ~new_P3_U3075 | ~new_P3_U3907;
  assign new_P3_R1077_U326 = ~new_P3_R1077_U137 | ~new_P3_R1077_U324;
  assign new_P3_R1077_U327 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1077_U328 = ~new_P3_R1077_U161;
  assign new_P3_R1077_U329 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1077_U330 = new_P3_U3437 | new_P3_U3072;
  assign new_P3_R1077_U331 = ~new_P3_R1077_U330 | ~new_P3_R1077_U92;
  assign new_P3_R1077_U332 = ~new_P3_R1077_U138 | ~new_P3_R1077_U331;
  assign new_P3_R1077_U333 = ~new_P3_R1077_U262 | ~new_P3_R1077_U59;
  assign new_P3_R1077_U334 = ~new_P3_U3440 | ~new_P3_U3068;
  assign new_P3_R1077_U335 = ~new_P3_R1077_U139 | ~new_P3_R1077_U333;
  assign new_P3_R1077_U336 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1077_U337 = ~new_P3_R1077_U250 | ~new_P3_R1077_U167;
  assign new_P3_R1077_U338 = ~new_P3_R1077_U93;
  assign new_P3_R1077_U339 = new_P3_U3425 | new_P3_U3071;
  assign new_P3_R1077_U340 = ~new_P3_R1077_U339 | ~new_P3_R1077_U93;
  assign new_P3_R1077_U341 = ~new_P3_R1077_U140 | ~new_P3_R1077_U340;
  assign new_P3_R1077_U342 = ~new_P3_R1077_U338 | ~new_P3_R1077_U172;
  assign new_P3_R1077_U343 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1077_U344 = ~new_P3_R1077_U141 | ~new_P3_R1077_U342;
  assign new_P3_R1077_U345 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1077_U346 = new_P3_U3416 | new_P3_U3082;
  assign new_P3_R1077_U347 = ~new_P3_R1077_U346 | ~new_P3_R1077_U40;
  assign new_P3_R1077_U348 = ~new_P3_R1077_U142 | ~new_P3_R1077_U347;
  assign new_P3_R1077_U349 = ~new_P3_R1077_U206 | ~new_P3_R1077_U171;
  assign new_P3_R1077_U350 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1077_U351 = ~new_P3_R1077_U143 | ~new_P3_R1077_U349;
  assign new_P3_R1077_U352 = ~new_P3_R1077_U207 | ~new_P3_R1077_U171;
  assign new_P3_R1077_U353 = ~new_P3_R1077_U204 | ~new_P3_R1077_U61;
  assign new_P3_R1077_U354 = ~new_P3_R1077_U214 | ~new_P3_R1077_U22;
  assign new_P3_R1077_U355 = ~new_P3_R1077_U228 | ~new_P3_R1077_U34;
  assign new_P3_R1077_U356 = ~new_P3_R1077_U231 | ~new_P3_R1077_U180;
  assign new_P3_R1077_U357 = ~new_P3_R1077_U314 | ~new_P3_R1077_U173;
  assign new_P3_R1077_U358 = ~new_P3_R1077_U298 | ~new_P3_R1077_U176;
  assign new_P3_R1077_U359 = ~new_P3_R1077_U329 | ~new_P3_R1077_U80;
  assign new_P3_R1077_U360 = ~new_P3_R1077_U282 | ~new_P3_R1077_U77;
  assign new_P3_R1077_U361 = ~new_P3_R1077_U336 | ~new_P3_R1077_U59;
  assign new_P3_R1077_U362 = ~new_P3_R1077_U345 | ~new_P3_R1077_U172;
  assign new_P3_R1077_U363 = ~new_P3_R1077_U250 | ~new_P3_R1077_U68;
  assign new_P3_R1077_U364 = ~new_P3_U3899 | ~new_P3_U3053;
  assign new_P3_R1077_U365 = ~new_P3_R1077_U296 | ~new_P3_R1077_U168;
  assign new_P3_R1077_U366 = ~new_P3_U3056 | ~new_P3_R1077_U295;
  assign new_P3_R1077_U367 = ~new_P3_U3901 | ~new_P3_R1077_U295;
  assign new_P3_R1077_U368 = ~new_P3_R1077_U301 | ~new_P3_R1077_U296 | ~new_P3_R1077_U168;
  assign new_P3_R1077_U369 = ~new_P3_R1077_U133 | ~new_P3_R1077_U155 | ~new_P3_R1077_U168;
  assign new_P3_R1077_U370 = ~new_P3_R1077_U297 | ~new_P3_R1077_U301;
  assign new_P3_R1077_U371 = ~new_P3_U3082 | ~new_P3_R1077_U39;
  assign new_P3_R1077_U372 = ~new_P3_U3416 | ~new_P3_R1077_U38;
  assign new_P3_R1077_U373 = ~new_P3_R1077_U372 | ~new_P3_R1077_U371;
  assign new_P3_R1077_U374 = ~new_P3_R1077_U352 | ~new_P3_R1077_U40;
  assign new_P3_R1077_U375 = ~new_P3_R1077_U373 | ~new_P3_R1077_U206;
  assign new_P3_R1077_U376 = ~new_P3_U3083 | ~new_P3_R1077_U36;
  assign new_P3_R1077_U377 = ~new_P3_U3413 | ~new_P3_R1077_U37;
  assign new_P3_R1077_U378 = ~new_P3_R1077_U377 | ~new_P3_R1077_U376;
  assign new_P3_R1077_U379 = ~new_P3_R1077_U353 | ~new_P3_R1077_U144;
  assign new_P3_R1077_U380 = ~new_P3_R1077_U203 | ~new_P3_R1077_U378;
  assign new_P3_R1077_U381 = ~new_P3_U3069 | ~new_P3_R1077_U23;
  assign new_P3_R1077_U382 = ~new_P3_U3410 | ~new_P3_R1077_U21;
  assign new_P3_R1077_U383 = ~new_P3_U3070 | ~new_P3_R1077_U19;
  assign new_P3_R1077_U384 = ~new_P3_U3407 | ~new_P3_R1077_U20;
  assign new_P3_R1077_U385 = ~new_P3_R1077_U384 | ~new_P3_R1077_U383;
  assign new_P3_R1077_U386 = ~new_P3_R1077_U354 | ~new_P3_R1077_U41;
  assign new_P3_R1077_U387 = ~new_P3_R1077_U385 | ~new_P3_R1077_U195;
  assign new_P3_R1077_U388 = ~new_P3_U3066 | ~new_P3_R1077_U35;
  assign new_P3_R1077_U389 = ~new_P3_U3404 | ~new_P3_R1077_U26;
  assign new_P3_R1077_U390 = ~new_P3_U3059 | ~new_P3_R1077_U24;
  assign new_P3_R1077_U391 = ~new_P3_U3401 | ~new_P3_R1077_U25;
  assign new_P3_R1077_U392 = ~new_P3_R1077_U391 | ~new_P3_R1077_U390;
  assign new_P3_R1077_U393 = ~new_P3_R1077_U355 | ~new_P3_R1077_U44;
  assign new_P3_R1077_U394 = ~new_P3_R1077_U392 | ~new_P3_R1077_U221;
  assign new_P3_R1077_U395 = ~new_P3_U3063 | ~new_P3_R1077_U32;
  assign new_P3_R1077_U396 = ~new_P3_U3398 | ~new_P3_R1077_U33;
  assign new_P3_R1077_U397 = ~new_P3_R1077_U396 | ~new_P3_R1077_U395;
  assign new_P3_R1077_U398 = ~new_P3_R1077_U356 | ~new_P3_R1077_U145;
  assign new_P3_R1077_U399 = ~new_P3_R1077_U230 | ~new_P3_R1077_U397;
  assign new_P3_R1077_U400 = ~new_P3_U3067 | ~new_P3_R1077_U27;
  assign new_P3_R1077_U401 = ~new_P3_U3395 | ~new_P3_R1077_U28;
  assign new_P3_R1077_U402 = ~new_P3_U3054 | ~new_P3_R1077_U147;
  assign new_P3_R1077_U403 = ~new_P3_U3908 | ~new_P3_R1077_U146;
  assign new_P3_R1077_U404 = ~new_P3_U3054 | ~new_P3_R1077_U147;
  assign new_P3_R1077_U405 = ~new_P3_U3908 | ~new_P3_R1077_U146;
  assign new_P3_R1077_U406 = ~new_P3_R1077_U405 | ~new_P3_R1077_U404;
  assign new_P3_R1077_U407 = ~new_P3_R1077_U148 | ~new_P3_R1077_U149;
  assign new_P3_R1077_U408 = ~new_P3_R1077_U305 | ~new_P3_R1077_U406;
  assign new_P3_R1077_U409 = ~new_P3_U3053 | ~new_P3_R1077_U88;
  assign new_P3_R1077_U410 = ~new_P3_U3899 | ~new_P3_R1077_U87;
  assign new_P3_R1077_U411 = ~new_P3_U3053 | ~new_P3_R1077_U88;
  assign new_P3_R1077_U412 = ~new_P3_U3899 | ~new_P3_R1077_U87;
  assign new_P3_R1077_U413 = ~new_P3_R1077_U412 | ~new_P3_R1077_U411;
  assign new_P3_R1077_U414 = ~new_P3_R1077_U150 | ~new_P3_R1077_U151;
  assign new_P3_R1077_U415 = ~new_P3_R1077_U303 | ~new_P3_R1077_U413;
  assign new_P3_R1077_U416 = ~new_P3_U3052 | ~new_P3_R1077_U46;
  assign new_P3_R1077_U417 = ~new_P3_U3900 | ~new_P3_R1077_U47;
  assign new_P3_R1077_U418 = ~new_P3_U3052 | ~new_P3_R1077_U46;
  assign new_P3_R1077_U419 = ~new_P3_U3900 | ~new_P3_R1077_U47;
  assign new_P3_R1077_U420 = ~new_P3_R1077_U419 | ~new_P3_R1077_U418;
  assign new_P3_R1077_U421 = ~new_P3_R1077_U152 | ~new_P3_R1077_U153;
  assign new_P3_R1077_U422 = ~new_P3_R1077_U300 | ~new_P3_R1077_U420;
  assign new_P3_R1077_U423 = ~new_P3_U3056 | ~new_P3_R1077_U49;
  assign new_P3_R1077_U424 = ~new_P3_U3901 | ~new_P3_R1077_U48;
  assign new_P3_R1077_U425 = ~new_P3_U3057 | ~new_P3_R1077_U50;
  assign new_P3_R1077_U426 = ~new_P3_U3902 | ~new_P3_R1077_U51;
  assign new_P3_R1077_U427 = ~new_P3_R1077_U426 | ~new_P3_R1077_U425;
  assign new_P3_R1077_U428 = ~new_P3_R1077_U357 | ~new_P3_R1077_U89;
  assign new_P3_R1077_U429 = ~new_P3_R1077_U427 | ~new_P3_R1077_U307;
  assign new_P3_R1077_U430 = ~new_P3_U3064 | ~new_P3_R1077_U52;
  assign new_P3_R1077_U431 = ~new_P3_U3903 | ~new_P3_R1077_U53;
  assign new_P3_R1077_U432 = ~new_P3_R1077_U431 | ~new_P3_R1077_U430;
  assign new_P3_R1077_U433 = ~new_P3_R1077_U358 | ~new_P3_R1077_U155;
  assign new_P3_R1077_U434 = ~new_P3_R1077_U294 | ~new_P3_R1077_U432;
  assign new_P3_R1077_U435 = ~new_P3_U3065 | ~new_P3_R1077_U84;
  assign new_P3_R1077_U436 = ~new_P3_U3904 | ~new_P3_R1077_U85;
  assign new_P3_R1077_U437 = ~new_P3_U3065 | ~new_P3_R1077_U84;
  assign new_P3_R1077_U438 = ~new_P3_U3904 | ~new_P3_R1077_U85;
  assign new_P3_R1077_U439 = ~new_P3_R1077_U438 | ~new_P3_R1077_U437;
  assign new_P3_R1077_U440 = ~new_P3_R1077_U156 | ~new_P3_R1077_U157;
  assign new_P3_R1077_U441 = ~new_P3_R1077_U290 | ~new_P3_R1077_U439;
  assign new_P3_R1077_U442 = ~new_P3_U3060 | ~new_P3_R1077_U82;
  assign new_P3_R1077_U443 = ~new_P3_U3905 | ~new_P3_R1077_U83;
  assign new_P3_R1077_U444 = ~new_P3_U3060 | ~new_P3_R1077_U82;
  assign new_P3_R1077_U445 = ~new_P3_U3905 | ~new_P3_R1077_U83;
  assign new_P3_R1077_U446 = ~new_P3_R1077_U445 | ~new_P3_R1077_U444;
  assign new_P3_R1077_U447 = ~new_P3_R1077_U158 | ~new_P3_R1077_U159;
  assign new_P3_R1077_U448 = ~new_P3_R1077_U286 | ~new_P3_R1077_U446;
  assign new_P3_R1077_U449 = ~new_P3_U3074 | ~new_P3_R1077_U54;
  assign new_P3_R1077_U450 = ~new_P3_U3906 | ~new_P3_R1077_U55;
  assign new_P3_R1077_U451 = ~new_P3_U3074 | ~new_P3_R1077_U54;
  assign new_P3_R1077_U452 = ~new_P3_U3906 | ~new_P3_R1077_U55;
  assign new_P3_R1077_U453 = ~new_P3_R1077_U452 | ~new_P3_R1077_U451;
  assign new_P3_R1077_U454 = ~new_P3_U3075 | ~new_P3_R1077_U81;
  assign new_P3_R1077_U455 = ~new_P3_U3907 | ~new_P3_R1077_U90;
  assign new_P3_R1077_U456 = ~new_P3_R1077_U182 | ~new_P3_R1077_U161;
  assign new_P3_R1077_U457 = ~new_P3_R1077_U328 | ~new_P3_R1077_U31;
  assign new_P3_R1077_U458 = ~new_P3_U3080 | ~new_P3_R1077_U78;
  assign new_P3_R1077_U459 = ~new_P3_U3445 | ~new_P3_R1077_U79;
  assign new_P3_R1077_U460 = ~new_P3_R1077_U459 | ~new_P3_R1077_U458;
  assign new_P3_R1077_U461 = ~new_P3_R1077_U359 | ~new_P3_R1077_U91;
  assign new_P3_R1077_U462 = ~new_P3_R1077_U460 | ~new_P3_R1077_U316;
  assign new_P3_R1077_U463 = ~new_P3_U3081 | ~new_P3_R1077_U75;
  assign new_P3_R1077_U464 = ~new_P3_U3443 | ~new_P3_R1077_U76;
  assign new_P3_R1077_U465 = ~new_P3_R1077_U464 | ~new_P3_R1077_U463;
  assign new_P3_R1077_U466 = ~new_P3_R1077_U360 | ~new_P3_R1077_U162;
  assign new_P3_R1077_U467 = ~new_P3_R1077_U270 | ~new_P3_R1077_U465;
  assign new_P3_R1077_U468 = ~new_P3_U3068 | ~new_P3_R1077_U60;
  assign new_P3_R1077_U469 = ~new_P3_U3440 | ~new_P3_R1077_U58;
  assign new_P3_R1077_U470 = ~new_P3_U3072 | ~new_P3_R1077_U56;
  assign new_P3_R1077_U471 = ~new_P3_U3437 | ~new_P3_R1077_U57;
  assign new_P3_R1077_U472 = ~new_P3_R1077_U471 | ~new_P3_R1077_U470;
  assign new_P3_R1077_U473 = ~new_P3_R1077_U361 | ~new_P3_R1077_U92;
  assign new_P3_R1077_U474 = ~new_P3_R1077_U472 | ~new_P3_R1077_U262;
  assign new_P3_R1077_U475 = ~new_P3_U3073 | ~new_P3_R1077_U73;
  assign new_P3_R1077_U476 = ~new_P3_U3434 | ~new_P3_R1077_U74;
  assign new_P3_R1077_U477 = ~new_P3_U3073 | ~new_P3_R1077_U73;
  assign new_P3_R1077_U478 = ~new_P3_U3434 | ~new_P3_R1077_U74;
  assign new_P3_R1077_U479 = ~new_P3_R1077_U478 | ~new_P3_R1077_U477;
  assign new_P3_R1077_U480 = ~new_P3_R1077_U163 | ~new_P3_R1077_U164;
  assign new_P3_R1077_U481 = ~new_P3_R1077_U258 | ~new_P3_R1077_U479;
  assign new_P3_R1077_U482 = ~new_P3_U3078 | ~new_P3_R1077_U71;
  assign new_P3_R1077_U483 = ~new_P3_U3431 | ~new_P3_R1077_U72;
  assign new_P3_R1077_U484 = ~new_P3_U3078 | ~new_P3_R1077_U71;
  assign new_P3_R1077_U485 = ~new_P3_U3431 | ~new_P3_R1077_U72;
  assign new_P3_R1077_U486 = ~new_P3_R1077_U485 | ~new_P3_R1077_U484;
  assign new_P3_R1077_U487 = ~new_P3_R1077_U165 | ~new_P3_R1077_U166;
  assign new_P3_R1077_U488 = ~new_P3_R1077_U254 | ~new_P3_R1077_U486;
  assign new_P3_R1077_U489 = ~new_P3_U3079 | ~new_P3_R1077_U69;
  assign new_P3_R1077_U490 = ~new_P3_U3428 | ~new_P3_R1077_U70;
  assign new_P3_R1077_U491 = ~new_P3_U3071 | ~new_P3_R1077_U64;
  assign new_P3_R1077_U492 = ~new_P3_U3425 | ~new_P3_R1077_U65;
  assign new_P3_R1077_U493 = ~new_P3_R1077_U492 | ~new_P3_R1077_U491;
  assign new_P3_R1077_U494 = ~new_P3_R1077_U362 | ~new_P3_R1077_U93;
  assign new_P3_R1077_U495 = ~new_P3_R1077_U493 | ~new_P3_R1077_U338;
  assign new_P3_R1077_U496 = ~new_P3_U3062 | ~new_P3_R1077_U66;
  assign new_P3_R1077_U497 = ~new_P3_U3422 | ~new_P3_R1077_U67;
  assign new_P3_R1077_U498 = ~new_P3_R1077_U497 | ~new_P3_R1077_U496;
  assign new_P3_R1077_U499 = ~new_P3_R1077_U363 | ~new_P3_R1077_U167;
  assign new_P3_R1077_U500 = ~new_P3_R1077_U244 | ~new_P3_R1077_U498;
  assign new_P3_R1077_U501 = ~new_P3_U3061 | ~new_P3_R1077_U62;
  assign new_P3_R1077_U502 = ~new_P3_U3419 | ~new_P3_R1077_U63;
  assign new_P3_R1077_U503 = ~new_P3_U3076 | ~new_P3_R1077_U29;
  assign new_P3_R1077_U504 = ~new_P3_U3387 | ~new_P3_R1077_U30;
  assign new_P3_R1143_U4 = new_P3_R1143_U179 & new_P3_R1143_U178;
  assign new_P3_R1143_U5 = new_P3_R1143_U197 & new_P3_R1143_U196;
  assign new_P3_R1143_U6 = new_P3_R1143_U237 & new_P3_R1143_U236;
  assign new_P3_R1143_U7 = new_P3_R1143_U246 & new_P3_R1143_U245;
  assign new_P3_R1143_U8 = new_P3_R1143_U264 & new_P3_R1143_U263;
  assign new_P3_R1143_U9 = new_P3_R1143_U272 & new_P3_R1143_U271;
  assign new_P3_R1143_U10 = new_P3_R1143_U351 & new_P3_R1143_U348;
  assign new_P3_R1143_U11 = new_P3_R1143_U344 & new_P3_R1143_U341;
  assign new_P3_R1143_U12 = new_P3_R1143_U335 & new_P3_R1143_U332;
  assign new_P3_R1143_U13 = new_P3_R1143_U326 & new_P3_R1143_U323;
  assign new_P3_R1143_U14 = new_P3_R1143_U320 & new_P3_R1143_U318;
  assign new_P3_R1143_U15 = new_P3_R1143_U313 & new_P3_R1143_U310;
  assign new_P3_R1143_U16 = new_P3_R1143_U235 & new_P3_R1143_U232;
  assign new_P3_R1143_U17 = new_P3_R1143_U227 & new_P3_R1143_U224;
  assign new_P3_R1143_U18 = new_P3_R1143_U213 & new_P3_R1143_U210;
  assign new_P3_R1143_U19 = ~new_P3_U3407;
  assign new_P3_R1143_U20 = ~new_P3_U3070;
  assign new_P3_R1143_U21 = ~new_P3_U3069;
  assign new_P3_R1143_U22 = ~new_P3_U3070 | ~new_P3_U3407;
  assign new_P3_R1143_U23 = ~new_P3_U3410;
  assign new_P3_R1143_U24 = ~new_P3_U3401;
  assign new_P3_R1143_U25 = ~new_P3_U3059;
  assign new_P3_R1143_U26 = ~new_P3_U3066;
  assign new_P3_R1143_U27 = ~new_P3_U3395;
  assign new_P3_R1143_U28 = ~new_P3_U3067;
  assign new_P3_R1143_U29 = ~new_P3_U3387;
  assign new_P3_R1143_U30 = ~new_P3_U3076;
  assign new_P3_R1143_U31 = ~new_P3_U3076 | ~new_P3_U3387;
  assign new_P3_R1143_U32 = ~new_P3_U3398;
  assign new_P3_R1143_U33 = ~new_P3_U3063;
  assign new_P3_R1143_U34 = ~new_P3_U3059 | ~new_P3_U3401;
  assign new_P3_R1143_U35 = ~new_P3_U3404;
  assign new_P3_R1143_U36 = ~new_P3_U3413;
  assign new_P3_R1143_U37 = ~new_P3_U3083;
  assign new_P3_R1143_U38 = ~new_P3_U3082;
  assign new_P3_R1143_U39 = ~new_P3_U3416;
  assign new_P3_R1143_U40 = ~new_P3_R1143_U63 | ~new_P3_R1143_U205;
  assign new_P3_R1143_U41 = ~new_P3_R1143_U117 | ~new_P3_R1143_U193;
  assign new_P3_R1143_U42 = ~new_P3_R1143_U182 | ~new_P3_R1143_U183;
  assign new_P3_R1143_U43 = ~new_P3_U3392 | ~new_P3_U3077;
  assign new_P3_R1143_U44 = ~new_P3_R1143_U122 | ~new_P3_R1143_U219;
  assign new_P3_R1143_U45 = ~new_P3_R1143_U216 | ~new_P3_R1143_U215;
  assign new_P3_R1143_U46 = ~new_P3_U3900;
  assign new_P3_R1143_U47 = ~new_P3_U3052;
  assign new_P3_R1143_U48 = ~new_P3_U3056;
  assign new_P3_R1143_U49 = ~new_P3_U3901;
  assign new_P3_R1143_U50 = ~new_P3_U3902;
  assign new_P3_R1143_U51 = ~new_P3_U3057;
  assign new_P3_R1143_U52 = ~new_P3_U3903;
  assign new_P3_R1143_U53 = ~new_P3_U3064;
  assign new_P3_R1143_U54 = ~new_P3_U3906;
  assign new_P3_R1143_U55 = ~new_P3_U3074;
  assign new_P3_R1143_U56 = ~new_P3_U3437;
  assign new_P3_R1143_U57 = ~new_P3_U3072;
  assign new_P3_R1143_U58 = ~new_P3_U3068;
  assign new_P3_R1143_U59 = ~new_P3_U3072 | ~new_P3_U3437;
  assign new_P3_R1143_U60 = ~new_P3_U3440;
  assign new_P3_R1143_U61 = ~new_P3_U3419;
  assign new_P3_R1143_U62 = ~new_P3_U3061;
  assign new_P3_R1143_U63 = ~new_P3_U3083 | ~new_P3_U3413;
  assign new_P3_R1143_U64 = ~new_P3_U3425;
  assign new_P3_R1143_U65 = ~new_P3_U3071;
  assign new_P3_R1143_U66 = ~new_P3_U3422;
  assign new_P3_R1143_U67 = ~new_P3_U3062;
  assign new_P3_R1143_U68 = ~new_P3_U3062 | ~new_P3_U3422;
  assign new_P3_R1143_U69 = ~new_P3_U3428;
  assign new_P3_R1143_U70 = ~new_P3_U3079;
  assign new_P3_R1143_U71 = ~new_P3_U3431;
  assign new_P3_R1143_U72 = ~new_P3_U3078;
  assign new_P3_R1143_U73 = ~new_P3_U3434;
  assign new_P3_R1143_U74 = ~new_P3_U3073;
  assign new_P3_R1143_U75 = ~new_P3_U3443;
  assign new_P3_R1143_U76 = ~new_P3_U3081;
  assign new_P3_R1143_U77 = ~new_P3_U3081 | ~new_P3_U3443;
  assign new_P3_R1143_U78 = ~new_P3_U3445;
  assign new_P3_R1143_U79 = ~new_P3_U3080;
  assign new_P3_R1143_U80 = ~new_P3_U3080 | ~new_P3_U3445;
  assign new_P3_R1143_U81 = ~new_P3_U3907;
  assign new_P3_R1143_U82 = ~new_P3_U3905;
  assign new_P3_R1143_U83 = ~new_P3_U3060;
  assign new_P3_R1143_U84 = ~new_P3_U3904;
  assign new_P3_R1143_U85 = ~new_P3_U3065;
  assign new_P3_R1143_U86 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1143_U87 = ~new_P3_U3053;
  assign new_P3_R1143_U88 = ~new_P3_U3899;
  assign new_P3_R1143_U89 = ~new_P3_R1143_U306 | ~new_P3_R1143_U176;
  assign new_P3_R1143_U90 = ~new_P3_U3075;
  assign new_P3_R1143_U91 = ~new_P3_R1143_U77 | ~new_P3_R1143_U315;
  assign new_P3_R1143_U92 = ~new_P3_R1143_U261 | ~new_P3_R1143_U260;
  assign new_P3_R1143_U93 = ~new_P3_R1143_U68 | ~new_P3_R1143_U337;
  assign new_P3_R1143_U94 = ~new_P3_R1143_U457 | ~new_P3_R1143_U456;
  assign new_P3_R1143_U95 = ~new_P3_R1143_U504 | ~new_P3_R1143_U503;
  assign new_P3_R1143_U96 = ~new_P3_R1143_U375 | ~new_P3_R1143_U374;
  assign new_P3_R1143_U97 = ~new_P3_R1143_U380 | ~new_P3_R1143_U379;
  assign new_P3_R1143_U98 = ~new_P3_R1143_U387 | ~new_P3_R1143_U386;
  assign new_P3_R1143_U99 = ~new_P3_R1143_U394 | ~new_P3_R1143_U393;
  assign new_P3_R1143_U100 = ~new_P3_R1143_U399 | ~new_P3_R1143_U398;
  assign new_P3_R1143_U101 = ~new_P3_R1143_U408 | ~new_P3_R1143_U407;
  assign new_P3_R1143_U102 = ~new_P3_R1143_U415 | ~new_P3_R1143_U414;
  assign new_P3_R1143_U103 = ~new_P3_R1143_U422 | ~new_P3_R1143_U421;
  assign new_P3_R1143_U104 = ~new_P3_R1143_U429 | ~new_P3_R1143_U428;
  assign new_P3_R1143_U105 = ~new_P3_R1143_U434 | ~new_P3_R1143_U433;
  assign new_P3_R1143_U106 = ~new_P3_R1143_U441 | ~new_P3_R1143_U440;
  assign new_P3_R1143_U107 = ~new_P3_R1143_U448 | ~new_P3_R1143_U447;
  assign new_P3_R1143_U108 = ~new_P3_R1143_U462 | ~new_P3_R1143_U461;
  assign new_P3_R1143_U109 = ~new_P3_R1143_U467 | ~new_P3_R1143_U466;
  assign new_P3_R1143_U110 = ~new_P3_R1143_U474 | ~new_P3_R1143_U473;
  assign new_P3_R1143_U111 = ~new_P3_R1143_U481 | ~new_P3_R1143_U480;
  assign new_P3_R1143_U112 = ~new_P3_R1143_U488 | ~new_P3_R1143_U487;
  assign new_P3_R1143_U113 = ~new_P3_R1143_U495 | ~new_P3_R1143_U494;
  assign new_P3_R1143_U114 = ~new_P3_R1143_U500 | ~new_P3_R1143_U499;
  assign new_P3_R1143_U115 = new_P3_R1143_U189 & new_P3_R1143_U187;
  assign new_P3_R1143_U116 = new_P3_R1143_U4 & new_P3_R1143_U180;
  assign new_P3_R1143_U117 = new_P3_R1143_U194 & new_P3_R1143_U192;
  assign new_P3_R1143_U118 = new_P3_R1143_U201 & new_P3_R1143_U200;
  assign new_P3_R1143_U119 = new_P3_R1143_U22 & new_P3_R1143_U382 & new_P3_R1143_U381;
  assign new_P3_R1143_U120 = new_P3_R1143_U212 & new_P3_R1143_U5;
  assign new_P3_R1143_U121 = new_P3_R1143_U181 & new_P3_R1143_U180;
  assign new_P3_R1143_U122 = new_P3_R1143_U220 & new_P3_R1143_U218;
  assign new_P3_R1143_U123 = new_P3_R1143_U34 & new_P3_R1143_U389 & new_P3_R1143_U388;
  assign new_P3_R1143_U124 = new_P3_R1143_U226 & new_P3_R1143_U4;
  assign new_P3_R1143_U125 = new_P3_R1143_U234 & new_P3_R1143_U181;
  assign new_P3_R1143_U126 = new_P3_R1143_U204 & new_P3_R1143_U6;
  assign new_P3_R1143_U127 = new_P3_R1143_U243 & new_P3_R1143_U239;
  assign new_P3_R1143_U128 = new_P3_R1143_U250 & new_P3_R1143_U7;
  assign new_P3_R1143_U129 = new_P3_R1143_U248 & new_P3_R1143_U172;
  assign new_P3_R1143_U130 = new_P3_R1143_U268 & new_P3_R1143_U267;
  assign new_P3_R1143_U131 = new_P3_R1143_U273 & new_P3_R1143_U9 & new_P3_R1143_U282;
  assign new_P3_R1143_U132 = new_P3_R1143_U285 & new_P3_R1143_U280;
  assign new_P3_R1143_U133 = new_P3_R1143_U301 & new_P3_R1143_U298;
  assign new_P3_R1143_U134 = new_P3_R1143_U368 & new_P3_R1143_U302;
  assign new_P3_R1143_U135 = new_P3_R1143_U160 & new_P3_R1143_U278;
  assign new_P3_R1143_U136 = new_P3_R1143_U80 & new_P3_R1143_U455 & new_P3_R1143_U454;
  assign new_P3_R1143_U137 = new_P3_R1143_U325 & new_P3_R1143_U9;
  assign new_P3_R1143_U138 = new_P3_R1143_U59 & new_P3_R1143_U469 & new_P3_R1143_U468;
  assign new_P3_R1143_U139 = new_P3_R1143_U334 & new_P3_R1143_U8;
  assign new_P3_R1143_U140 = new_P3_R1143_U172 & new_P3_R1143_U490 & new_P3_R1143_U489;
  assign new_P3_R1143_U141 = new_P3_R1143_U343 & new_P3_R1143_U7;
  assign new_P3_R1143_U142 = new_P3_R1143_U171 & new_P3_R1143_U502 & new_P3_R1143_U501;
  assign new_P3_R1143_U143 = new_P3_R1143_U350 & new_P3_R1143_U6;
  assign new_P3_R1143_U144 = ~new_P3_R1143_U118 | ~new_P3_R1143_U202;
  assign new_P3_R1143_U145 = ~new_P3_R1143_U217 | ~new_P3_R1143_U229;
  assign new_P3_R1143_U146 = ~new_P3_U3054;
  assign new_P3_R1143_U147 = ~new_P3_U3908;
  assign new_P3_R1143_U148 = new_P3_R1143_U403 & new_P3_R1143_U402;
  assign new_P3_R1143_U149 = ~new_P3_R1143_U364 | ~new_P3_R1143_U304 | ~new_P3_R1143_U169;
  assign new_P3_R1143_U150 = new_P3_R1143_U410 & new_P3_R1143_U409;
  assign new_P3_R1143_U151 = ~new_P3_R1143_U134 | ~new_P3_R1143_U370 | ~new_P3_R1143_U369;
  assign new_P3_R1143_U152 = new_P3_R1143_U417 & new_P3_R1143_U416;
  assign new_P3_R1143_U153 = ~new_P3_R1143_U86 | ~new_P3_R1143_U365 | ~new_P3_R1143_U299;
  assign new_P3_R1143_U154 = new_P3_R1143_U424 & new_P3_R1143_U423;
  assign new_P3_R1143_U155 = ~new_P3_R1143_U293 | ~new_P3_R1143_U292;
  assign new_P3_R1143_U156 = new_P3_R1143_U436 & new_P3_R1143_U435;
  assign new_P3_R1143_U157 = ~new_P3_R1143_U289 | ~new_P3_R1143_U288;
  assign new_P3_R1143_U158 = new_P3_R1143_U443 & new_P3_R1143_U442;
  assign new_P3_R1143_U159 = ~new_P3_R1143_U132 | ~new_P3_R1143_U284;
  assign new_P3_R1143_U160 = new_P3_R1143_U450 & new_P3_R1143_U449;
  assign new_P3_R1143_U161 = ~new_P3_R1143_U43 | ~new_P3_R1143_U327;
  assign new_P3_R1143_U162 = ~new_P3_R1143_U130 | ~new_P3_R1143_U269;
  assign new_P3_R1143_U163 = new_P3_R1143_U476 & new_P3_R1143_U475;
  assign new_P3_R1143_U164 = ~new_P3_R1143_U257 | ~new_P3_R1143_U256;
  assign new_P3_R1143_U165 = new_P3_R1143_U483 & new_P3_R1143_U482;
  assign new_P3_R1143_U166 = ~new_P3_R1143_U253 | ~new_P3_R1143_U252;
  assign new_P3_R1143_U167 = ~new_P3_R1143_U127 | ~new_P3_R1143_U242;
  assign new_P3_R1143_U168 = ~new_P3_R1143_U367 | ~new_P3_R1143_U366;
  assign new_P3_R1143_U169 = ~new_P3_U3053 | ~new_P3_R1143_U151;
  assign new_P3_R1143_U170 = ~new_P3_R1143_U34;
  assign new_P3_R1143_U171 = ~new_P3_U3416 | ~new_P3_U3082;
  assign new_P3_R1143_U172 = ~new_P3_U3071 | ~new_P3_U3425;
  assign new_P3_R1143_U173 = ~new_P3_U3057 | ~new_P3_U3902;
  assign new_P3_R1143_U174 = ~new_P3_R1143_U68;
  assign new_P3_R1143_U175 = ~new_P3_R1143_U77;
  assign new_P3_R1143_U176 = ~new_P3_U3064 | ~new_P3_U3903;
  assign new_P3_R1143_U177 = ~new_P3_R1143_U63;
  assign new_P3_R1143_U178 = new_P3_U3066 | new_P3_U3404;
  assign new_P3_R1143_U179 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1143_U180 = new_P3_U3398 | new_P3_U3063;
  assign new_P3_R1143_U181 = new_P3_U3395 | new_P3_U3067;
  assign new_P3_R1143_U182 = ~new_P3_R1143_U31;
  assign new_P3_R1143_U183 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1143_U184 = ~new_P3_R1143_U42;
  assign new_P3_R1143_U185 = ~new_P3_R1143_U43;
  assign new_P3_R1143_U186 = ~new_P3_R1143_U42 | ~new_P3_R1143_U43;
  assign new_P3_R1143_U187 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1143_U188 = ~new_P3_R1143_U186 | ~new_P3_R1143_U181;
  assign new_P3_R1143_U189 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1143_U190 = ~new_P3_R1143_U115 | ~new_P3_R1143_U188;
  assign new_P3_R1143_U191 = ~new_P3_R1143_U35 | ~new_P3_R1143_U34;
  assign new_P3_R1143_U192 = ~new_P3_U3066 | ~new_P3_R1143_U191;
  assign new_P3_R1143_U193 = ~new_P3_R1143_U116 | ~new_P3_R1143_U190;
  assign new_P3_R1143_U194 = ~new_P3_U3404 | ~new_P3_R1143_U170;
  assign new_P3_R1143_U195 = ~new_P3_R1143_U41;
  assign new_P3_R1143_U196 = new_P3_U3069 | new_P3_U3410;
  assign new_P3_R1143_U197 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1143_U198 = ~new_P3_R1143_U22;
  assign new_P3_R1143_U199 = ~new_P3_R1143_U23 | ~new_P3_R1143_U22;
  assign new_P3_R1143_U200 = ~new_P3_U3069 | ~new_P3_R1143_U199;
  assign new_P3_R1143_U201 = ~new_P3_U3410 | ~new_P3_R1143_U198;
  assign new_P3_R1143_U202 = ~new_P3_R1143_U5 | ~new_P3_R1143_U41;
  assign new_P3_R1143_U203 = ~new_P3_R1143_U144;
  assign new_P3_R1143_U204 = new_P3_U3413 | new_P3_U3083;
  assign new_P3_R1143_U205 = ~new_P3_R1143_U204 | ~new_P3_R1143_U144;
  assign new_P3_R1143_U206 = ~new_P3_R1143_U40;
  assign new_P3_R1143_U207 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1143_U208 = new_P3_U3407 | new_P3_U3070;
  assign new_P3_R1143_U209 = ~new_P3_R1143_U208 | ~new_P3_R1143_U41;
  assign new_P3_R1143_U210 = ~new_P3_R1143_U119 | ~new_P3_R1143_U209;
  assign new_P3_R1143_U211 = ~new_P3_R1143_U195 | ~new_P3_R1143_U22;
  assign new_P3_R1143_U212 = ~new_P3_U3410 | ~new_P3_U3069;
  assign new_P3_R1143_U213 = ~new_P3_R1143_U120 | ~new_P3_R1143_U211;
  assign new_P3_R1143_U214 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1143_U215 = ~new_P3_R1143_U185 | ~new_P3_R1143_U181;
  assign new_P3_R1143_U216 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1143_U217 = ~new_P3_R1143_U45;
  assign new_P3_R1143_U218 = ~new_P3_R1143_U121 | ~new_P3_R1143_U184;
  assign new_P3_R1143_U219 = ~new_P3_R1143_U45 | ~new_P3_R1143_U180;
  assign new_P3_R1143_U220 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1143_U221 = ~new_P3_R1143_U44;
  assign new_P3_R1143_U222 = new_P3_U3401 | new_P3_U3059;
  assign new_P3_R1143_U223 = ~new_P3_R1143_U222 | ~new_P3_R1143_U44;
  assign new_P3_R1143_U224 = ~new_P3_R1143_U123 | ~new_P3_R1143_U223;
  assign new_P3_R1143_U225 = ~new_P3_R1143_U221 | ~new_P3_R1143_U34;
  assign new_P3_R1143_U226 = ~new_P3_U3404 | ~new_P3_U3066;
  assign new_P3_R1143_U227 = ~new_P3_R1143_U124 | ~new_P3_R1143_U225;
  assign new_P3_R1143_U228 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1143_U229 = ~new_P3_R1143_U184 | ~new_P3_R1143_U181;
  assign new_P3_R1143_U230 = ~new_P3_R1143_U145;
  assign new_P3_R1143_U231 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1143_U232 = ~new_P3_R1143_U42 | ~new_P3_R1143_U43 | ~new_P3_R1143_U401 | ~new_P3_R1143_U400;
  assign new_P3_R1143_U233 = ~new_P3_R1143_U43 | ~new_P3_R1143_U42;
  assign new_P3_R1143_U234 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1143_U235 = ~new_P3_R1143_U125 | ~new_P3_R1143_U233;
  assign new_P3_R1143_U236 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1143_U237 = new_P3_U3061 | new_P3_U3419;
  assign new_P3_R1143_U238 = ~new_P3_R1143_U177 | ~new_P3_R1143_U6;
  assign new_P3_R1143_U239 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1143_U240 = ~new_P3_R1143_U171 | ~new_P3_R1143_U238;
  assign new_P3_R1143_U241 = new_P3_U3419 | new_P3_U3061;
  assign new_P3_R1143_U242 = ~new_P3_R1143_U126 | ~new_P3_R1143_U144;
  assign new_P3_R1143_U243 = ~new_P3_R1143_U241 | ~new_P3_R1143_U240;
  assign new_P3_R1143_U244 = ~new_P3_R1143_U167;
  assign new_P3_R1143_U245 = new_P3_U3079 | new_P3_U3428;
  assign new_P3_R1143_U246 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1143_U247 = ~new_P3_R1143_U174 | ~new_P3_R1143_U7;
  assign new_P3_R1143_U248 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1143_U249 = ~new_P3_R1143_U129 | ~new_P3_R1143_U247;
  assign new_P3_R1143_U250 = new_P3_U3422 | new_P3_U3062;
  assign new_P3_R1143_U251 = new_P3_U3428 | new_P3_U3079;
  assign new_P3_R1143_U252 = ~new_P3_R1143_U128 | ~new_P3_R1143_U167;
  assign new_P3_R1143_U253 = ~new_P3_R1143_U251 | ~new_P3_R1143_U249;
  assign new_P3_R1143_U254 = ~new_P3_R1143_U166;
  assign new_P3_R1143_U255 = new_P3_U3431 | new_P3_U3078;
  assign new_P3_R1143_U256 = ~new_P3_R1143_U255 | ~new_P3_R1143_U166;
  assign new_P3_R1143_U257 = ~new_P3_U3078 | ~new_P3_U3431;
  assign new_P3_R1143_U258 = ~new_P3_R1143_U164;
  assign new_P3_R1143_U259 = new_P3_U3434 | new_P3_U3073;
  assign new_P3_R1143_U260 = ~new_P3_R1143_U259 | ~new_P3_R1143_U164;
  assign new_P3_R1143_U261 = ~new_P3_U3073 | ~new_P3_U3434;
  assign new_P3_R1143_U262 = ~new_P3_R1143_U92;
  assign new_P3_R1143_U263 = new_P3_U3068 | new_P3_U3440;
  assign new_P3_R1143_U264 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1143_U265 = ~new_P3_R1143_U59;
  assign new_P3_R1143_U266 = ~new_P3_R1143_U60 | ~new_P3_R1143_U59;
  assign new_P3_R1143_U267 = ~new_P3_U3068 | ~new_P3_R1143_U266;
  assign new_P3_R1143_U268 = ~new_P3_U3440 | ~new_P3_R1143_U265;
  assign new_P3_R1143_U269 = ~new_P3_R1143_U8 | ~new_P3_R1143_U92;
  assign new_P3_R1143_U270 = ~new_P3_R1143_U162;
  assign new_P3_R1143_U271 = new_P3_U3075 | new_P3_U3907;
  assign new_P3_R1143_U272 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1143_U273 = new_P3_U3074 | new_P3_U3906;
  assign new_P3_R1143_U274 = ~new_P3_R1143_U80;
  assign new_P3_R1143_U275 = ~new_P3_U3907 | ~new_P3_R1143_U274;
  assign new_P3_R1143_U276 = ~new_P3_R1143_U275 | ~new_P3_R1143_U90;
  assign new_P3_R1143_U277 = ~new_P3_R1143_U80 | ~new_P3_R1143_U81;
  assign new_P3_R1143_U278 = ~new_P3_R1143_U277 | ~new_P3_R1143_U276;
  assign new_P3_R1143_U279 = ~new_P3_R1143_U175 | ~new_P3_R1143_U9;
  assign new_P3_R1143_U280 = ~new_P3_U3074 | ~new_P3_U3906;
  assign new_P3_R1143_U281 = ~new_P3_R1143_U278 | ~new_P3_R1143_U279;
  assign new_P3_R1143_U282 = new_P3_U3443 | new_P3_U3081;
  assign new_P3_R1143_U283 = new_P3_U3906 | new_P3_U3074;
  assign new_P3_R1143_U284 = ~new_P3_R1143_U162 | ~new_P3_R1143_U131;
  assign new_P3_R1143_U285 = ~new_P3_R1143_U283 | ~new_P3_R1143_U281;
  assign new_P3_R1143_U286 = ~new_P3_R1143_U159;
  assign new_P3_R1143_U287 = new_P3_U3905 | new_P3_U3060;
  assign new_P3_R1143_U288 = ~new_P3_R1143_U287 | ~new_P3_R1143_U159;
  assign new_P3_R1143_U289 = ~new_P3_U3060 | ~new_P3_U3905;
  assign new_P3_R1143_U290 = ~new_P3_R1143_U157;
  assign new_P3_R1143_U291 = new_P3_U3904 | new_P3_U3065;
  assign new_P3_R1143_U292 = ~new_P3_R1143_U291 | ~new_P3_R1143_U157;
  assign new_P3_R1143_U293 = ~new_P3_U3065 | ~new_P3_U3904;
  assign new_P3_R1143_U294 = ~new_P3_R1143_U155;
  assign new_P3_R1143_U295 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1143_U296 = ~new_P3_R1143_U176 | ~new_P3_R1143_U173;
  assign new_P3_R1143_U297 = ~new_P3_R1143_U86;
  assign new_P3_R1143_U298 = new_P3_U3903 | new_P3_U3064;
  assign new_P3_R1143_U299 = ~new_P3_R1143_U168 | ~new_P3_R1143_U155 | ~new_P3_R1143_U298;
  assign new_P3_R1143_U300 = ~new_P3_R1143_U153;
  assign new_P3_R1143_U301 = new_P3_U3900 | new_P3_U3052;
  assign new_P3_R1143_U302 = ~new_P3_U3052 | ~new_P3_U3900;
  assign new_P3_R1143_U303 = ~new_P3_R1143_U151;
  assign new_P3_R1143_U304 = ~new_P3_U3899 | ~new_P3_R1143_U151;
  assign new_P3_R1143_U305 = ~new_P3_R1143_U149;
  assign new_P3_R1143_U306 = ~new_P3_R1143_U298 | ~new_P3_R1143_U155;
  assign new_P3_R1143_U307 = ~new_P3_R1143_U89;
  assign new_P3_R1143_U308 = new_P3_U3902 | new_P3_U3057;
  assign new_P3_R1143_U309 = ~new_P3_R1143_U308 | ~new_P3_R1143_U89;
  assign new_P3_R1143_U310 = ~new_P3_R1143_U154 | ~new_P3_R1143_U309 | ~new_P3_R1143_U173;
  assign new_P3_R1143_U311 = ~new_P3_R1143_U307 | ~new_P3_R1143_U173;
  assign new_P3_R1143_U312 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1143_U313 = ~new_P3_R1143_U168 | ~new_P3_R1143_U311 | ~new_P3_R1143_U312;
  assign new_P3_R1143_U314 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1143_U315 = ~new_P3_R1143_U282 | ~new_P3_R1143_U162;
  assign new_P3_R1143_U316 = ~new_P3_R1143_U91;
  assign new_P3_R1143_U317 = ~new_P3_R1143_U9 | ~new_P3_R1143_U91;
  assign new_P3_R1143_U318 = ~new_P3_R1143_U135 | ~new_P3_R1143_U317;
  assign new_P3_R1143_U319 = ~new_P3_R1143_U317 | ~new_P3_R1143_U278;
  assign new_P3_R1143_U320 = ~new_P3_R1143_U453 | ~new_P3_R1143_U319;
  assign new_P3_R1143_U321 = new_P3_U3445 | new_P3_U3080;
  assign new_P3_R1143_U322 = ~new_P3_R1143_U321 | ~new_P3_R1143_U91;
  assign new_P3_R1143_U323 = ~new_P3_R1143_U136 | ~new_P3_R1143_U322;
  assign new_P3_R1143_U324 = ~new_P3_R1143_U316 | ~new_P3_R1143_U80;
  assign new_P3_R1143_U325 = ~new_P3_U3075 | ~new_P3_U3907;
  assign new_P3_R1143_U326 = ~new_P3_R1143_U137 | ~new_P3_R1143_U324;
  assign new_P3_R1143_U327 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1143_U328 = ~new_P3_R1143_U161;
  assign new_P3_R1143_U329 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1143_U330 = new_P3_U3437 | new_P3_U3072;
  assign new_P3_R1143_U331 = ~new_P3_R1143_U330 | ~new_P3_R1143_U92;
  assign new_P3_R1143_U332 = ~new_P3_R1143_U138 | ~new_P3_R1143_U331;
  assign new_P3_R1143_U333 = ~new_P3_R1143_U262 | ~new_P3_R1143_U59;
  assign new_P3_R1143_U334 = ~new_P3_U3440 | ~new_P3_U3068;
  assign new_P3_R1143_U335 = ~new_P3_R1143_U139 | ~new_P3_R1143_U333;
  assign new_P3_R1143_U336 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1143_U337 = ~new_P3_R1143_U250 | ~new_P3_R1143_U167;
  assign new_P3_R1143_U338 = ~new_P3_R1143_U93;
  assign new_P3_R1143_U339 = new_P3_U3425 | new_P3_U3071;
  assign new_P3_R1143_U340 = ~new_P3_R1143_U339 | ~new_P3_R1143_U93;
  assign new_P3_R1143_U341 = ~new_P3_R1143_U140 | ~new_P3_R1143_U340;
  assign new_P3_R1143_U342 = ~new_P3_R1143_U338 | ~new_P3_R1143_U172;
  assign new_P3_R1143_U343 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1143_U344 = ~new_P3_R1143_U141 | ~new_P3_R1143_U342;
  assign new_P3_R1143_U345 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1143_U346 = new_P3_U3416 | new_P3_U3082;
  assign new_P3_R1143_U347 = ~new_P3_R1143_U346 | ~new_P3_R1143_U40;
  assign new_P3_R1143_U348 = ~new_P3_R1143_U142 | ~new_P3_R1143_U347;
  assign new_P3_R1143_U349 = ~new_P3_R1143_U206 | ~new_P3_R1143_U171;
  assign new_P3_R1143_U350 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1143_U351 = ~new_P3_R1143_U143 | ~new_P3_R1143_U349;
  assign new_P3_R1143_U352 = ~new_P3_R1143_U207 | ~new_P3_R1143_U171;
  assign new_P3_R1143_U353 = ~new_P3_R1143_U204 | ~new_P3_R1143_U63;
  assign new_P3_R1143_U354 = ~new_P3_R1143_U214 | ~new_P3_R1143_U22;
  assign new_P3_R1143_U355 = ~new_P3_R1143_U228 | ~new_P3_R1143_U34;
  assign new_P3_R1143_U356 = ~new_P3_R1143_U231 | ~new_P3_R1143_U180;
  assign new_P3_R1143_U357 = ~new_P3_R1143_U314 | ~new_P3_R1143_U173;
  assign new_P3_R1143_U358 = ~new_P3_R1143_U298 | ~new_P3_R1143_U176;
  assign new_P3_R1143_U359 = ~new_P3_R1143_U329 | ~new_P3_R1143_U80;
  assign new_P3_R1143_U360 = ~new_P3_R1143_U282 | ~new_P3_R1143_U77;
  assign new_P3_R1143_U361 = ~new_P3_R1143_U336 | ~new_P3_R1143_U59;
  assign new_P3_R1143_U362 = ~new_P3_R1143_U345 | ~new_P3_R1143_U172;
  assign new_P3_R1143_U363 = ~new_P3_R1143_U250 | ~new_P3_R1143_U68;
  assign new_P3_R1143_U364 = ~new_P3_U3899 | ~new_P3_U3053;
  assign new_P3_R1143_U365 = ~new_P3_R1143_U296 | ~new_P3_R1143_U168;
  assign new_P3_R1143_U366 = ~new_P3_U3056 | ~new_P3_R1143_U295;
  assign new_P3_R1143_U367 = ~new_P3_U3901 | ~new_P3_R1143_U295;
  assign new_P3_R1143_U368 = ~new_P3_R1143_U301 | ~new_P3_R1143_U296 | ~new_P3_R1143_U168;
  assign new_P3_R1143_U369 = ~new_P3_R1143_U133 | ~new_P3_R1143_U155 | ~new_P3_R1143_U168;
  assign new_P3_R1143_U370 = ~new_P3_R1143_U297 | ~new_P3_R1143_U301;
  assign new_P3_R1143_U371 = ~new_P3_U3082 | ~new_P3_R1143_U39;
  assign new_P3_R1143_U372 = ~new_P3_U3416 | ~new_P3_R1143_U38;
  assign new_P3_R1143_U373 = ~new_P3_R1143_U372 | ~new_P3_R1143_U371;
  assign new_P3_R1143_U374 = ~new_P3_R1143_U352 | ~new_P3_R1143_U40;
  assign new_P3_R1143_U375 = ~new_P3_R1143_U373 | ~new_P3_R1143_U206;
  assign new_P3_R1143_U376 = ~new_P3_U3083 | ~new_P3_R1143_U36;
  assign new_P3_R1143_U377 = ~new_P3_U3413 | ~new_P3_R1143_U37;
  assign new_P3_R1143_U378 = ~new_P3_R1143_U377 | ~new_P3_R1143_U376;
  assign new_P3_R1143_U379 = ~new_P3_R1143_U353 | ~new_P3_R1143_U144;
  assign new_P3_R1143_U380 = ~new_P3_R1143_U203 | ~new_P3_R1143_U378;
  assign new_P3_R1143_U381 = ~new_P3_U3069 | ~new_P3_R1143_U23;
  assign new_P3_R1143_U382 = ~new_P3_U3410 | ~new_P3_R1143_U21;
  assign new_P3_R1143_U383 = ~new_P3_U3070 | ~new_P3_R1143_U19;
  assign new_P3_R1143_U384 = ~new_P3_U3407 | ~new_P3_R1143_U20;
  assign new_P3_R1143_U385 = ~new_P3_R1143_U384 | ~new_P3_R1143_U383;
  assign new_P3_R1143_U386 = ~new_P3_R1143_U354 | ~new_P3_R1143_U41;
  assign new_P3_R1143_U387 = ~new_P3_R1143_U385 | ~new_P3_R1143_U195;
  assign new_P3_R1143_U388 = ~new_P3_U3066 | ~new_P3_R1143_U35;
  assign new_P3_R1143_U389 = ~new_P3_U3404 | ~new_P3_R1143_U26;
  assign new_P3_R1143_U390 = ~new_P3_U3059 | ~new_P3_R1143_U24;
  assign new_P3_R1143_U391 = ~new_P3_U3401 | ~new_P3_R1143_U25;
  assign new_P3_R1143_U392 = ~new_P3_R1143_U391 | ~new_P3_R1143_U390;
  assign new_P3_R1143_U393 = ~new_P3_R1143_U355 | ~new_P3_R1143_U44;
  assign new_P3_R1143_U394 = ~new_P3_R1143_U392 | ~new_P3_R1143_U221;
  assign new_P3_R1143_U395 = ~new_P3_U3063 | ~new_P3_R1143_U32;
  assign new_P3_R1143_U396 = ~new_P3_U3398 | ~new_P3_R1143_U33;
  assign new_P3_R1143_U397 = ~new_P3_R1143_U396 | ~new_P3_R1143_U395;
  assign new_P3_R1143_U398 = ~new_P3_R1143_U356 | ~new_P3_R1143_U145;
  assign new_P3_R1143_U399 = ~new_P3_R1143_U230 | ~new_P3_R1143_U397;
  assign new_P3_R1143_U400 = ~new_P3_U3067 | ~new_P3_R1143_U27;
  assign new_P3_R1143_U401 = ~new_P3_U3395 | ~new_P3_R1143_U28;
  assign new_P3_R1143_U402 = ~new_P3_U3054 | ~new_P3_R1143_U147;
  assign new_P3_R1143_U403 = ~new_P3_U3908 | ~new_P3_R1143_U146;
  assign new_P3_R1143_U404 = ~new_P3_U3054 | ~new_P3_R1143_U147;
  assign new_P3_R1143_U405 = ~new_P3_U3908 | ~new_P3_R1143_U146;
  assign new_P3_R1143_U406 = ~new_P3_R1143_U405 | ~new_P3_R1143_U404;
  assign new_P3_R1143_U407 = ~new_P3_R1143_U148 | ~new_P3_R1143_U149;
  assign new_P3_R1143_U408 = ~new_P3_R1143_U305 | ~new_P3_R1143_U406;
  assign new_P3_R1143_U409 = ~new_P3_U3053 | ~new_P3_R1143_U88;
  assign new_P3_R1143_U410 = ~new_P3_U3899 | ~new_P3_R1143_U87;
  assign new_P3_R1143_U411 = ~new_P3_U3053 | ~new_P3_R1143_U88;
  assign new_P3_R1143_U412 = ~new_P3_U3899 | ~new_P3_R1143_U87;
  assign new_P3_R1143_U413 = ~new_P3_R1143_U412 | ~new_P3_R1143_U411;
  assign new_P3_R1143_U414 = ~new_P3_R1143_U150 | ~new_P3_R1143_U151;
  assign new_P3_R1143_U415 = ~new_P3_R1143_U303 | ~new_P3_R1143_U413;
  assign new_P3_R1143_U416 = ~new_P3_U3052 | ~new_P3_R1143_U46;
  assign new_P3_R1143_U417 = ~new_P3_U3900 | ~new_P3_R1143_U47;
  assign new_P3_R1143_U418 = ~new_P3_U3052 | ~new_P3_R1143_U46;
  assign new_P3_R1143_U419 = ~new_P3_U3900 | ~new_P3_R1143_U47;
  assign new_P3_R1143_U420 = ~new_P3_R1143_U419 | ~new_P3_R1143_U418;
  assign new_P3_R1143_U421 = ~new_P3_R1143_U152 | ~new_P3_R1143_U153;
  assign new_P3_R1143_U422 = ~new_P3_R1143_U300 | ~new_P3_R1143_U420;
  assign new_P3_R1143_U423 = ~new_P3_U3056 | ~new_P3_R1143_U49;
  assign new_P3_R1143_U424 = ~new_P3_U3901 | ~new_P3_R1143_U48;
  assign new_P3_R1143_U425 = ~new_P3_U3057 | ~new_P3_R1143_U50;
  assign new_P3_R1143_U426 = ~new_P3_U3902 | ~new_P3_R1143_U51;
  assign new_P3_R1143_U427 = ~new_P3_R1143_U426 | ~new_P3_R1143_U425;
  assign new_P3_R1143_U428 = ~new_P3_R1143_U357 | ~new_P3_R1143_U89;
  assign new_P3_R1143_U429 = ~new_P3_R1143_U427 | ~new_P3_R1143_U307;
  assign new_P3_R1143_U430 = ~new_P3_U3064 | ~new_P3_R1143_U52;
  assign new_P3_R1143_U431 = ~new_P3_U3903 | ~new_P3_R1143_U53;
  assign new_P3_R1143_U432 = ~new_P3_R1143_U431 | ~new_P3_R1143_U430;
  assign new_P3_R1143_U433 = ~new_P3_R1143_U358 | ~new_P3_R1143_U155;
  assign new_P3_R1143_U434 = ~new_P3_R1143_U294 | ~new_P3_R1143_U432;
  assign new_P3_R1143_U435 = ~new_P3_U3065 | ~new_P3_R1143_U84;
  assign new_P3_R1143_U436 = ~new_P3_U3904 | ~new_P3_R1143_U85;
  assign new_P3_R1143_U437 = ~new_P3_U3065 | ~new_P3_R1143_U84;
  assign new_P3_R1143_U438 = ~new_P3_U3904 | ~new_P3_R1143_U85;
  assign new_P3_R1143_U439 = ~new_P3_R1143_U438 | ~new_P3_R1143_U437;
  assign new_P3_R1143_U440 = ~new_P3_R1143_U156 | ~new_P3_R1143_U157;
  assign new_P3_R1143_U441 = ~new_P3_R1143_U290 | ~new_P3_R1143_U439;
  assign new_P3_R1143_U442 = ~new_P3_U3060 | ~new_P3_R1143_U82;
  assign new_P3_R1143_U443 = ~new_P3_U3905 | ~new_P3_R1143_U83;
  assign new_P3_R1143_U444 = ~new_P3_U3060 | ~new_P3_R1143_U82;
  assign new_P3_R1143_U445 = ~new_P3_U3905 | ~new_P3_R1143_U83;
  assign new_P3_R1143_U446 = ~new_P3_R1143_U445 | ~new_P3_R1143_U444;
  assign new_P3_R1143_U447 = ~new_P3_R1143_U158 | ~new_P3_R1143_U159;
  assign new_P3_R1143_U448 = ~new_P3_R1143_U286 | ~new_P3_R1143_U446;
  assign new_P3_R1143_U449 = ~new_P3_U3074 | ~new_P3_R1143_U54;
  assign new_P3_R1143_U450 = ~new_P3_U3906 | ~new_P3_R1143_U55;
  assign new_P3_R1143_U451 = ~new_P3_U3074 | ~new_P3_R1143_U54;
  assign new_P3_R1143_U452 = ~new_P3_U3906 | ~new_P3_R1143_U55;
  assign new_P3_R1143_U453 = ~new_P3_R1143_U452 | ~new_P3_R1143_U451;
  assign new_P3_R1143_U454 = ~new_P3_U3075 | ~new_P3_R1143_U81;
  assign new_P3_R1143_U455 = ~new_P3_U3907 | ~new_P3_R1143_U90;
  assign new_P3_R1143_U456 = ~new_P3_R1143_U182 | ~new_P3_R1143_U161;
  assign new_P3_R1143_U457 = ~new_P3_R1143_U328 | ~new_P3_R1143_U31;
  assign new_P3_R1143_U458 = ~new_P3_U3080 | ~new_P3_R1143_U78;
  assign new_P3_R1143_U459 = ~new_P3_U3445 | ~new_P3_R1143_U79;
  assign new_P3_R1143_U460 = ~new_P3_R1143_U459 | ~new_P3_R1143_U458;
  assign new_P3_R1143_U461 = ~new_P3_R1143_U359 | ~new_P3_R1143_U91;
  assign new_P3_R1143_U462 = ~new_P3_R1143_U460 | ~new_P3_R1143_U316;
  assign new_P3_R1143_U463 = ~new_P3_U3081 | ~new_P3_R1143_U75;
  assign new_P3_R1143_U464 = ~new_P3_U3443 | ~new_P3_R1143_U76;
  assign new_P3_R1143_U465 = ~new_P3_R1143_U464 | ~new_P3_R1143_U463;
  assign new_P3_R1143_U466 = ~new_P3_R1143_U360 | ~new_P3_R1143_U162;
  assign new_P3_R1143_U467 = ~new_P3_R1143_U270 | ~new_P3_R1143_U465;
  assign new_P3_R1143_U468 = ~new_P3_U3068 | ~new_P3_R1143_U60;
  assign new_P3_R1143_U469 = ~new_P3_U3440 | ~new_P3_R1143_U58;
  assign new_P3_R1143_U470 = ~new_P3_U3072 | ~new_P3_R1143_U56;
  assign new_P3_R1143_U471 = ~new_P3_U3437 | ~new_P3_R1143_U57;
  assign new_P3_R1143_U472 = ~new_P3_R1143_U471 | ~new_P3_R1143_U470;
  assign new_P3_R1143_U473 = ~new_P3_R1143_U361 | ~new_P3_R1143_U92;
  assign new_P3_R1143_U474 = ~new_P3_R1143_U472 | ~new_P3_R1143_U262;
  assign new_P3_R1143_U475 = ~new_P3_U3073 | ~new_P3_R1143_U73;
  assign new_P3_R1143_U476 = ~new_P3_U3434 | ~new_P3_R1143_U74;
  assign new_P3_R1143_U477 = ~new_P3_U3073 | ~new_P3_R1143_U73;
  assign new_P3_R1143_U478 = ~new_P3_U3434 | ~new_P3_R1143_U74;
  assign new_P3_R1143_U479 = ~new_P3_R1143_U478 | ~new_P3_R1143_U477;
  assign new_P3_R1143_U480 = ~new_P3_R1143_U163 | ~new_P3_R1143_U164;
  assign new_P3_R1143_U481 = ~new_P3_R1143_U258 | ~new_P3_R1143_U479;
  assign new_P3_R1143_U482 = ~new_P3_U3078 | ~new_P3_R1143_U71;
  assign new_P3_R1143_U483 = ~new_P3_U3431 | ~new_P3_R1143_U72;
  assign new_P3_R1143_U484 = ~new_P3_U3078 | ~new_P3_R1143_U71;
  assign new_P3_R1143_U485 = ~new_P3_U3431 | ~new_P3_R1143_U72;
  assign new_P3_R1143_U486 = ~new_P3_R1143_U485 | ~new_P3_R1143_U484;
  assign new_P3_R1143_U487 = ~new_P3_R1143_U165 | ~new_P3_R1143_U166;
  assign new_P3_R1143_U488 = ~new_P3_R1143_U254 | ~new_P3_R1143_U486;
  assign new_P3_R1143_U489 = ~new_P3_U3079 | ~new_P3_R1143_U69;
  assign new_P3_R1143_U490 = ~new_P3_U3428 | ~new_P3_R1143_U70;
  assign new_P3_R1143_U491 = ~new_P3_U3071 | ~new_P3_R1143_U64;
  assign new_P3_R1143_U492 = ~new_P3_U3425 | ~new_P3_R1143_U65;
  assign new_P3_R1143_U493 = ~new_P3_R1143_U492 | ~new_P3_R1143_U491;
  assign new_P3_R1143_U494 = ~new_P3_R1143_U362 | ~new_P3_R1143_U93;
  assign new_P3_R1143_U495 = ~new_P3_R1143_U493 | ~new_P3_R1143_U338;
  assign new_P3_R1143_U496 = ~new_P3_U3062 | ~new_P3_R1143_U66;
  assign new_P3_R1143_U497 = ~new_P3_U3422 | ~new_P3_R1143_U67;
  assign new_P3_R1143_U498 = ~new_P3_R1143_U497 | ~new_P3_R1143_U496;
  assign new_P3_R1143_U499 = ~new_P3_R1143_U363 | ~new_P3_R1143_U167;
  assign new_P3_R1143_U500 = ~new_P3_R1143_U244 | ~new_P3_R1143_U498;
  assign new_P3_R1143_U501 = ~new_P3_U3061 | ~new_P3_R1143_U61;
  assign new_P3_R1143_U502 = ~new_P3_U3419 | ~new_P3_R1143_U62;
  assign new_P3_R1143_U503 = ~new_P3_U3076 | ~new_P3_R1143_U29;
  assign new_P3_R1143_U504 = ~new_P3_U3387 | ~new_P3_R1143_U30;
  assign new_P3_R1158_U4 = new_P3_R1158_U227 & new_P3_R1158_U226;
  assign new_P3_R1158_U5 = new_P3_R1158_U238 & new_P3_R1158_U237;
  assign new_P3_R1158_U6 = new_P3_R1158_U263 & new_P3_R1158_U262;
  assign new_P3_R1158_U7 = new_P3_R1158_U277 & new_P3_R1158_U276;
  assign new_P3_R1158_U8 = new_P3_R1158_U289 & new_P3_R1158_U288;
  assign new_P3_R1158_U9 = new_P3_R1158_U6 & new_P3_R1158_U267;
  assign new_P3_R1158_U10 = new_P3_R1158_U5 & new_P3_R1158_U235;
  assign new_P3_R1158_U11 = new_P3_R1158_U9 & new_P3_R1158_U260;
  assign new_P3_R1158_U12 = new_P3_R1158_U535 & new_P3_R1158_U534;
  assign new_P3_R1158_U13 = new_P3_R1158_U345 & new_P3_R1158_U342;
  assign new_P3_R1158_U14 = new_P3_R1158_U336 & new_P3_R1158_U333;
  assign new_P3_R1158_U15 = new_P3_R1158_U329 & new_P3_R1158_U326;
  assign new_P3_R1158_U16 = new_P3_R1158_U142 & new_P3_R1158_U537 & new_P3_R1158_U536;
  assign new_P3_R1158_U17 = new_P3_R1158_U256 & new_P3_R1158_U253;
  assign new_P3_R1158_U18 = new_P3_R1158_U249 & new_P3_R1158_U246;
  assign new_P3_R1158_U19 = ~new_P3_U3056 | ~new_P3_R1158_U306;
  assign new_P3_R1158_U20 = ~new_P3_U3152;
  assign new_P3_R1158_U21 = ~new_P3_U3083;
  assign new_P3_R1158_U22 = ~new_P3_U3070;
  assign new_P3_R1158_U23 = ~new_P3_U3070 | ~new_P3_R1158_U67;
  assign new_P3_R1158_U24 = ~new_P3_U3069;
  assign new_P3_R1158_U25 = ~new_P3_U3066;
  assign new_P3_R1158_U26 = ~new_P3_U3066 | ~new_P3_R1158_U69;
  assign new_P3_R1158_U27 = ~new_P3_U3067;
  assign new_P3_R1158_U28 = ~new_P3_U3067 | ~new_P3_R1158_U70;
  assign new_P3_R1158_U29 = ~new_P3_U3063;
  assign new_P3_R1158_U30 = ~new_P3_U3077;
  assign new_P3_R1158_U31 = ~new_P3_U3076;
  assign new_P3_R1158_U32 = ~new_P3_U3059;
  assign new_P3_R1158_U33 = ~new_P3_U3082;
  assign new_P3_R1158_U34 = ~new_P3_R1158_U362 | ~new_P3_R1158_U359 | ~new_P3_R1158_U241;
  assign new_P3_R1158_U35 = ~new_P3_R1158_U379 | ~new_P3_R1158_U26;
  assign new_P3_R1158_U36 = ~new_P3_R1158_U360 | ~new_P3_R1158_U361 | ~new_P3_R1158_U224;
  assign new_P3_R1158_U37 = ~new_P3_U3052;
  assign new_P3_R1158_U38 = ~new_P3_U3057;
  assign new_P3_R1158_U39 = ~new_P3_U3064;
  assign new_P3_R1158_U40 = ~new_P3_U3056;
  assign new_P3_R1158_U41 = ~new_P3_U3072;
  assign new_P3_R1158_U42 = ~new_P3_U3072 | ~new_P3_R1158_U79;
  assign new_P3_R1158_U43 = ~new_P3_U3068;
  assign new_P3_R1158_U44 = ~new_P3_U3078;
  assign new_P3_R1158_U45 = ~new_P3_U3071;
  assign new_P3_R1158_U46 = ~new_P3_U3062;
  assign new_P3_R1158_U47 = ~new_P3_U3062 | ~new_P3_R1158_U84;
  assign new_P3_R1158_U48 = ~new_P3_U3079;
  assign new_P3_R1158_U49 = ~new_P3_U3061;
  assign new_P3_R1158_U50 = ~new_P3_U3061 | ~new_P3_R1158_U85;
  assign new_P3_R1158_U51 = ~new_P3_U3073;
  assign new_P3_R1158_U52 = ~new_P3_U3081;
  assign new_P3_R1158_U53 = ~new_P3_U3075;
  assign new_P3_R1158_U54 = ~new_P3_U3080;
  assign new_P3_R1158_U55 = ~new_P3_U3080 | ~new_P3_R1158_U88;
  assign new_P3_R1158_U56 = ~new_P3_U3074;
  assign new_P3_R1158_U57 = ~new_P3_U3060;
  assign new_P3_R1158_U58 = ~new_P3_U3065;
  assign new_P3_R1158_U59 = ~new_P3_U3057 | ~new_P3_R1158_U76;
  assign new_P3_R1158_U60 = ~new_P3_U3064 | ~new_P3_R1158_U77;
  assign new_P3_R1158_U61 = ~new_P3_R1158_U55 | ~new_P3_R1158_U322;
  assign new_P3_R1158_U62 = ~new_P3_R1158_U274 | ~new_P3_R1158_U273;
  assign new_P3_R1158_U63 = ~new_P3_R1158_U365 | ~new_P3_R1158_U269;
  assign new_P3_R1158_U64 = ~new_P3_R1158_U47 | ~new_P3_R1158_U338;
  assign new_P3_R1158_U65 = ~new_P3_R1158_U394 | ~new_P3_R1158_U393;
  assign new_P3_R1158_U66 = ~new_P3_R1158_U426 | ~new_P3_R1158_U425;
  assign new_P3_R1158_U67 = ~new_P3_R1158_U423 | ~new_P3_R1158_U422;
  assign new_P3_R1158_U68 = ~new_P3_R1158_U420 | ~new_P3_R1158_U419;
  assign new_P3_R1158_U69 = ~new_P3_R1158_U417 | ~new_P3_R1158_U416;
  assign new_P3_R1158_U70 = ~new_P3_R1158_U414 | ~new_P3_R1158_U413;
  assign new_P3_R1158_U71 = ~new_P3_R1158_U411 | ~new_P3_R1158_U410;
  assign new_P3_R1158_U72 = ~new_P3_R1158_U405 | ~new_P3_R1158_U404;
  assign new_P3_R1158_U73 = ~new_P3_R1158_U408 | ~new_P3_R1158_U407;
  assign new_P3_R1158_U74 = ~new_P3_R1158_U402 | ~new_P3_R1158_U401;
  assign new_P3_R1158_U75 = ~new_P3_R1158_U466 | ~new_P3_R1158_U465;
  assign new_P3_R1158_U76 = ~new_P3_R1158_U514 | ~new_P3_R1158_U513;
  assign new_P3_R1158_U77 = ~new_P3_R1158_U517 | ~new_P3_R1158_U516;
  assign new_P3_R1158_U78 = ~new_P3_R1158_U511 | ~new_P3_R1158_U510;
  assign new_P3_R1158_U79 = ~new_P3_R1158_U490 | ~new_P3_R1158_U489;
  assign new_P3_R1158_U80 = ~new_P3_R1158_U487 | ~new_P3_R1158_U486;
  assign new_P3_R1158_U81 = ~new_P3_R1158_U481 | ~new_P3_R1158_U480;
  assign new_P3_R1158_U82 = ~new_P3_R1158_U478 | ~new_P3_R1158_U477;
  assign new_P3_R1158_U83 = ~new_P3_R1158_U475 | ~new_P3_R1158_U474;
  assign new_P3_R1158_U84 = ~new_P3_R1158_U472 | ~new_P3_R1158_U471;
  assign new_P3_R1158_U85 = ~new_P3_R1158_U469 | ~new_P3_R1158_U468;
  assign new_P3_R1158_U86 = ~new_P3_R1158_U484 | ~new_P3_R1158_U483;
  assign new_P3_R1158_U87 = ~new_P3_R1158_U493 | ~new_P3_R1158_U492;
  assign new_P3_R1158_U88 = ~new_P3_R1158_U502 | ~new_P3_R1158_U501;
  assign new_P3_R1158_U89 = ~new_P3_R1158_U496 | ~new_P3_R1158_U495;
  assign new_P3_R1158_U90 = ~new_P3_R1158_U499 | ~new_P3_R1158_U498;
  assign new_P3_R1158_U91 = ~new_P3_R1158_U505 | ~new_P3_R1158_U504;
  assign new_P3_R1158_U92 = ~new_P3_R1158_U508 | ~new_P3_R1158_U507;
  assign new_P3_R1158_U93 = ~new_P3_R1158_U523 | ~new_P3_R1158_U522;
  assign new_P3_R1158_U94 = ~new_P3_R1158_U632 | ~new_P3_R1158_U631;
  assign new_P3_R1158_U95 = ~new_P3_R1158_U429 | ~new_P3_R1158_U428;
  assign new_P3_R1158_U96 = ~new_P3_R1158_U436 | ~new_P3_R1158_U435;
  assign new_P3_R1158_U97 = ~new_P3_R1158_U443 | ~new_P3_R1158_U442;
  assign new_P3_R1158_U98 = ~new_P3_R1158_U450 | ~new_P3_R1158_U449;
  assign new_P3_R1158_U99 = ~new_P3_R1158_U457 | ~new_P3_R1158_U456;
  assign new_P3_R1158_U100 = ~new_P3_R1158_U464 | ~new_P3_R1158_U463;
  assign new_P3_R1158_U101 = ~new_P3_R1158_U526 | ~new_P3_R1158_U525;
  assign new_P3_R1158_U102 = ~new_P3_R1158_U533 | ~new_P3_R1158_U532;
  assign new_P3_R1158_U103 = new_P3_R1158_U320 & new_P3_R1158_U209;
  assign new_P3_R1158_U104 = new_P3_R1158_U141 & new_P3_R1158_U12;
  assign new_P3_R1158_U105 = ~new_P3_R1158_U542 | ~new_P3_R1158_U541;
  assign new_P3_R1158_U106 = ~new_P3_R1158_U547 | ~new_P3_R1158_U546;
  assign new_P3_R1158_U107 = ~new_P3_R1158_U554 | ~new_P3_R1158_U553;
  assign new_P3_R1158_U108 = ~new_P3_R1158_U561 | ~new_P3_R1158_U560;
  assign new_P3_R1158_U109 = ~new_P3_R1158_U568 | ~new_P3_R1158_U567;
  assign new_P3_R1158_U110 = ~new_P3_R1158_U575 | ~new_P3_R1158_U574;
  assign new_P3_R1158_U111 = ~new_P3_R1158_U580 | ~new_P3_R1158_U579;
  assign new_P3_R1158_U112 = ~new_P3_R1158_U587 | ~new_P3_R1158_U586;
  assign new_P3_R1158_U113 = ~new_P3_R1158_U594 | ~new_P3_R1158_U593;
  assign new_P3_R1158_U114 = ~new_P3_R1158_U601 | ~new_P3_R1158_U600;
  assign new_P3_R1158_U115 = ~new_P3_R1158_U608 | ~new_P3_R1158_U607;
  assign new_P3_R1158_U116 = ~new_P3_R1158_U615 | ~new_P3_R1158_U614;
  assign new_P3_R1158_U117 = ~new_P3_R1158_U620 | ~new_P3_R1158_U619;
  assign new_P3_R1158_U118 = ~new_P3_R1158_U627 | ~new_P3_R1158_U626;
  assign new_P3_R1158_U119 = new_P3_R1158_U73 & new_P3_U3152;
  assign new_P3_R1158_U120 = new_P3_R1158_U230 & new_P3_R1158_U229;
  assign new_P3_R1158_U121 = new_P3_R1158_U242 & new_P3_R1158_U10;
  assign new_P3_R1158_U122 = new_P3_R1158_U364 & new_P3_R1158_U243;
  assign new_P3_R1158_U123 = new_P3_R1158_U23 & new_P3_R1158_U438 & new_P3_R1158_U437;
  assign new_P3_R1158_U124 = new_P3_R1158_U248 & new_P3_R1158_U5;
  assign new_P3_R1158_U125 = new_P3_R1158_U28 & new_P3_R1158_U459 & new_P3_R1158_U458;
  assign new_P3_R1158_U126 = new_P3_R1158_U255 & new_P3_R1158_U4;
  assign new_P3_R1158_U127 = new_P3_R1158_U265 & new_P3_R1158_U213;
  assign new_P3_R1158_U128 = new_P3_R1158_U270 & new_P3_R1158_U11;
  assign new_P3_R1158_U129 = new_P3_R1158_U373 & new_P3_R1158_U271;
  assign new_P3_R1158_U130 = new_P3_R1158_U281 & new_P3_R1158_U280;
  assign new_P3_R1158_U131 = new_P3_R1158_U293 & new_P3_R1158_U8;
  assign new_P3_R1158_U132 = new_P3_R1158_U291 & new_P3_R1158_U214;
  assign new_P3_R1158_U133 = new_P3_R1158_U314 & new_P3_R1158_U376;
  assign new_P3_R1158_U134 = new_P3_R1158_U316 & new_P3_R1158_U307;
  assign new_P3_R1158_U135 = new_P3_R1158_U316 & new_P3_R1158_U369;
  assign new_P3_R1158_U136 = new_P3_R1158_U374 & new_P3_R1158_U315;
  assign new_P3_R1158_U137 = ~new_P3_R1158_U520 | ~new_P3_R1158_U519;
  assign new_P3_R1158_U138 = new_P3_R1158_U515 & new_P3_R1158_U38;
  assign new_P3_R1158_U139 = new_P3_R1158_U320 & new_P3_R1158_U215;
  assign new_P3_R1158_U140 = new_P3_R1158_U320 & new_P3_R1158_U218;
  assign new_P3_R1158_U141 = new_P3_R1158_U60 & new_P3_R1158_U59;
  assign new_P3_R1158_U142 = new_P3_R1158_U392 & new_P3_R1158_U391 & new_P3_R1158_U319;
  assign new_P3_R1158_U143 = new_P3_R1158_U214 & new_P3_R1158_U563 & new_P3_R1158_U562;
  assign new_P3_R1158_U144 = new_P3_R1158_U328 & new_P3_R1158_U8;
  assign new_P3_R1158_U145 = new_P3_R1158_U42 & new_P3_R1158_U589 & new_P3_R1158_U588;
  assign new_P3_R1158_U146 = new_P3_R1158_U335 & new_P3_R1158_U7;
  assign new_P3_R1158_U147 = new_P3_R1158_U213 & new_P3_R1158_U610 & new_P3_R1158_U609;
  assign new_P3_R1158_U148 = new_P3_R1158_U344 & new_P3_R1158_U6;
  assign new_P3_R1158_U149 = ~new_P3_R1158_U629 | ~new_P3_R1158_U628;
  assign new_P3_R1158_U150 = ~new_P3_U3416;
  assign new_P3_R1158_U151 = new_P3_R1158_U397 & new_P3_R1158_U396;
  assign new_P3_R1158_U152 = ~new_P3_U3401;
  assign new_P3_R1158_U153 = ~new_P3_U3392;
  assign new_P3_R1158_U154 = ~new_P3_U3387;
  assign new_P3_R1158_U155 = ~new_P3_U3398;
  assign new_P3_R1158_U156 = ~new_P3_U3395;
  assign new_P3_R1158_U157 = ~new_P3_U3404;
  assign new_P3_R1158_U158 = ~new_P3_U3410;
  assign new_P3_R1158_U159 = ~new_P3_U3407;
  assign new_P3_R1158_U160 = ~new_P3_U3413;
  assign new_P3_R1158_U161 = ~new_P3_R1158_U122 | ~new_P3_R1158_U383;
  assign new_P3_R1158_U162 = new_P3_R1158_U431 & new_P3_R1158_U430;
  assign new_P3_R1158_U163 = ~new_P3_R1158_U363 | ~new_P3_R1158_U381;
  assign new_P3_R1158_U164 = new_P3_R1158_U445 & new_P3_R1158_U444;
  assign new_P3_R1158_U165 = ~new_P3_R1158_U356 | ~new_P3_R1158_U233 | ~new_P3_R1158_U211;
  assign new_P3_R1158_U166 = new_P3_R1158_U452 & new_P3_R1158_U451;
  assign new_P3_R1158_U167 = ~new_P3_R1158_U120 | ~new_P3_R1158_U231;
  assign new_P3_R1158_U168 = ~new_P3_U3900;
  assign new_P3_R1158_U169 = ~new_P3_U3419;
  assign new_P3_R1158_U170 = ~new_P3_U3422;
  assign new_P3_R1158_U171 = ~new_P3_U3428;
  assign new_P3_R1158_U172 = ~new_P3_U3425;
  assign new_P3_R1158_U173 = ~new_P3_U3431;
  assign new_P3_R1158_U174 = ~new_P3_U3434;
  assign new_P3_R1158_U175 = ~new_P3_U3440;
  assign new_P3_R1158_U176 = ~new_P3_U3437;
  assign new_P3_R1158_U177 = ~new_P3_U3443;
  assign new_P3_R1158_U178 = ~new_P3_U3906;
  assign new_P3_R1158_U179 = ~new_P3_U3907;
  assign new_P3_R1158_U180 = ~new_P3_U3445;
  assign new_P3_R1158_U181 = ~new_P3_U3905;
  assign new_P3_R1158_U182 = ~new_P3_U3904;
  assign new_P3_R1158_U183 = ~new_P3_U3901;
  assign new_P3_R1158_U184 = ~new_P3_U3902;
  assign new_P3_R1158_U185 = ~new_P3_U3903;
  assign new_P3_R1158_U186 = ~new_P3_U3053;
  assign new_P3_R1158_U187 = ~new_P3_U3899;
  assign new_P3_R1158_U188 = new_P3_R1158_U528 & new_P3_R1158_U527;
  assign new_P3_R1158_U189 = ~new_P3_R1158_U311 | ~new_P3_R1158_U310;
  assign new_P3_R1158_U190 = ~new_P3_R1158_U309 | ~new_P3_R1158_U192;
  assign new_P3_R1158_U191 = ~new_P3_R1158_U60 | ~new_P3_R1158_U190;
  assign new_P3_R1158_U192 = ~new_P3_R1158_U304 | ~new_P3_R1158_U303;
  assign new_P3_R1158_U193 = new_P3_R1158_U549 & new_P3_R1158_U548;
  assign new_P3_R1158_U194 = ~new_P3_R1158_U300 | ~new_P3_R1158_U299;
  assign new_P3_R1158_U195 = new_P3_R1158_U556 & new_P3_R1158_U555;
  assign new_P3_R1158_U196 = ~new_P3_R1158_U296 | ~new_P3_R1158_U295;
  assign new_P3_R1158_U197 = new_P3_R1158_U570 & new_P3_R1158_U569;
  assign new_P3_R1158_U198 = ~new_P3_R1158_U221 | ~new_P3_R1158_U220;
  assign new_P3_R1158_U199 = ~new_P3_R1158_U286 | ~new_P3_R1158_U285;
  assign new_P3_R1158_U200 = new_P3_R1158_U582 & new_P3_R1158_U581;
  assign new_P3_R1158_U201 = ~new_P3_R1158_U130 | ~new_P3_R1158_U282;
  assign new_P3_R1158_U202 = new_P3_R1158_U596 & new_P3_R1158_U595;
  assign new_P3_R1158_U203 = ~new_P3_R1158_U129 | ~new_P3_R1158_U389;
  assign new_P3_R1158_U204 = new_P3_R1158_U603 & new_P3_R1158_U602;
  assign new_P3_R1158_U205 = ~new_P3_R1158_U372 | ~new_P3_R1158_U387;
  assign new_P3_R1158_U206 = ~new_P3_R1158_U385 | ~new_P3_R1158_U50;
  assign new_P3_R1158_U207 = new_P3_R1158_U622 & new_P3_R1158_U621;
  assign new_P3_R1158_U208 = ~new_P3_R1158_U357 | ~new_P3_R1158_U258 | ~new_P3_R1158_U210;
  assign new_P3_R1158_U209 = ~new_P3_R1158_U19 | ~new_P3_R1158_U367;
  assign new_P3_R1158_U210 = ~new_P3_R1158_U65 | ~new_P3_R1158_U161;
  assign new_P3_R1158_U211 = ~new_P3_R1158_U74 | ~new_P3_R1158_U167;
  assign new_P3_R1158_U212 = ~new_P3_R1158_U28;
  assign new_P3_R1158_U213 = ~new_P3_U3071 | ~new_P3_R1158_U82;
  assign new_P3_R1158_U214 = ~new_P3_U3075 | ~new_P3_R1158_U90;
  assign new_P3_R1158_U215 = ~new_P3_R1158_U59;
  assign new_P3_R1158_U216 = ~new_P3_R1158_U47;
  assign new_P3_R1158_U217 = ~new_P3_R1158_U55;
  assign new_P3_R1158_U218 = ~new_P3_R1158_U60;
  assign new_P3_R1158_U219 = ~new_P3_R1158_U409 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U220 = ~new_P3_U3076 | ~new_P3_R1158_U219;
  assign new_P3_R1158_U221 = ~new_P3_U3152 | ~new_P3_R1158_U73;
  assign new_P3_R1158_U222 = ~new_P3_R1158_U198;
  assign new_P3_R1158_U223 = ~new_P3_R1158_U406 | ~new_P3_R1158_U30;
  assign new_P3_R1158_U224 = ~new_P3_U3077 | ~new_P3_R1158_U72;
  assign new_P3_R1158_U225 = ~new_P3_R1158_U36;
  assign new_P3_R1158_U226 = ~new_P3_R1158_U412 | ~new_P3_R1158_U29;
  assign new_P3_R1158_U227 = ~new_P3_R1158_U415 | ~new_P3_R1158_U27;
  assign new_P3_R1158_U228 = ~new_P3_R1158_U29 | ~new_P3_R1158_U28;
  assign new_P3_R1158_U229 = ~new_P3_R1158_U71 | ~new_P3_R1158_U228;
  assign new_P3_R1158_U230 = ~new_P3_U3063 | ~new_P3_R1158_U212;
  assign new_P3_R1158_U231 = ~new_P3_R1158_U4 | ~new_P3_R1158_U36;
  assign new_P3_R1158_U232 = ~new_P3_R1158_U167;
  assign new_P3_R1158_U233 = ~new_P3_U3059 | ~new_P3_R1158_U167;
  assign new_P3_R1158_U234 = ~new_P3_R1158_U165;
  assign new_P3_R1158_U235 = ~new_P3_R1158_U418 | ~new_P3_R1158_U25;
  assign new_P3_R1158_U236 = ~new_P3_R1158_U26;
  assign new_P3_R1158_U237 = ~new_P3_R1158_U421 | ~new_P3_R1158_U24;
  assign new_P3_R1158_U238 = ~new_P3_R1158_U424 | ~new_P3_R1158_U22;
  assign new_P3_R1158_U239 = ~new_P3_R1158_U23;
  assign new_P3_R1158_U240 = ~new_P3_R1158_U24 | ~new_P3_R1158_U23;
  assign new_P3_R1158_U241 = ~new_P3_U3069 | ~new_P3_R1158_U239;
  assign new_P3_R1158_U242 = ~new_P3_R1158_U427 | ~new_P3_R1158_U21;
  assign new_P3_R1158_U243 = ~new_P3_U3083 | ~new_P3_R1158_U66;
  assign new_P3_R1158_U244 = ~new_P3_R1158_U424 | ~new_P3_R1158_U22;
  assign new_P3_R1158_U245 = ~new_P3_R1158_U244 | ~new_P3_R1158_U35;
  assign new_P3_R1158_U246 = ~new_P3_R1158_U123 | ~new_P3_R1158_U245;
  assign new_P3_R1158_U247 = ~new_P3_R1158_U380 | ~new_P3_R1158_U23;
  assign new_P3_R1158_U248 = ~new_P3_U3069 | ~new_P3_R1158_U68;
  assign new_P3_R1158_U249 = ~new_P3_R1158_U124 | ~new_P3_R1158_U247;
  assign new_P3_R1158_U250 = ~new_P3_R1158_U424 | ~new_P3_R1158_U22;
  assign new_P3_R1158_U251 = ~new_P3_R1158_U415 | ~new_P3_R1158_U27;
  assign new_P3_R1158_U252 = ~new_P3_R1158_U251 | ~new_P3_R1158_U36;
  assign new_P3_R1158_U253 = ~new_P3_R1158_U125 | ~new_P3_R1158_U252;
  assign new_P3_R1158_U254 = ~new_P3_R1158_U225 | ~new_P3_R1158_U28;
  assign new_P3_R1158_U255 = ~new_P3_U3063 | ~new_P3_R1158_U71;
  assign new_P3_R1158_U256 = ~new_P3_R1158_U126 | ~new_P3_R1158_U254;
  assign new_P3_R1158_U257 = ~new_P3_R1158_U415 | ~new_P3_R1158_U27;
  assign new_P3_R1158_U258 = ~new_P3_U3082 | ~new_P3_R1158_U161;
  assign new_P3_R1158_U259 = ~new_P3_R1158_U208;
  assign new_P3_R1158_U260 = ~new_P3_R1158_U470 | ~new_P3_R1158_U49;
  assign new_P3_R1158_U261 = ~new_P3_R1158_U50;
  assign new_P3_R1158_U262 = ~new_P3_R1158_U476 | ~new_P3_R1158_U48;
  assign new_P3_R1158_U263 = ~new_P3_R1158_U479 | ~new_P3_R1158_U45;
  assign new_P3_R1158_U264 = ~new_P3_R1158_U216 | ~new_P3_R1158_U6;
  assign new_P3_R1158_U265 = ~new_P3_U3079 | ~new_P3_R1158_U83;
  assign new_P3_R1158_U266 = ~new_P3_R1158_U127 | ~new_P3_R1158_U264;
  assign new_P3_R1158_U267 = ~new_P3_R1158_U473 | ~new_P3_R1158_U46;
  assign new_P3_R1158_U268 = ~new_P3_R1158_U476 | ~new_P3_R1158_U48;
  assign new_P3_R1158_U269 = ~new_P3_R1158_U268 | ~new_P3_R1158_U266;
  assign new_P3_R1158_U270 = ~new_P3_R1158_U482 | ~new_P3_R1158_U44;
  assign new_P3_R1158_U271 = ~new_P3_U3078 | ~new_P3_R1158_U81;
  assign new_P3_R1158_U272 = ~new_P3_R1158_U485 | ~new_P3_R1158_U51;
  assign new_P3_R1158_U273 = ~new_P3_R1158_U272 | ~new_P3_R1158_U203;
  assign new_P3_R1158_U274 = ~new_P3_U3073 | ~new_P3_R1158_U86;
  assign new_P3_R1158_U275 = ~new_P3_R1158_U62;
  assign new_P3_R1158_U276 = ~new_P3_R1158_U488 | ~new_P3_R1158_U43;
  assign new_P3_R1158_U277 = ~new_P3_R1158_U491 | ~new_P3_R1158_U41;
  assign new_P3_R1158_U278 = ~new_P3_R1158_U42;
  assign new_P3_R1158_U279 = ~new_P3_R1158_U43 | ~new_P3_R1158_U42;
  assign new_P3_R1158_U280 = ~new_P3_R1158_U80 | ~new_P3_R1158_U279;
  assign new_P3_R1158_U281 = ~new_P3_U3068 | ~new_P3_R1158_U278;
  assign new_P3_R1158_U282 = ~new_P3_R1158_U7 | ~new_P3_R1158_U62;
  assign new_P3_R1158_U283 = ~new_P3_R1158_U201;
  assign new_P3_R1158_U284 = ~new_P3_R1158_U494 | ~new_P3_R1158_U52;
  assign new_P3_R1158_U285 = ~new_P3_R1158_U284 | ~new_P3_R1158_U201;
  assign new_P3_R1158_U286 = ~new_P3_U3081 | ~new_P3_R1158_U87;
  assign new_P3_R1158_U287 = ~new_P3_R1158_U199;
  assign new_P3_R1158_U288 = ~new_P3_R1158_U497 | ~new_P3_R1158_U56;
  assign new_P3_R1158_U289 = ~new_P3_R1158_U500 | ~new_P3_R1158_U53;
  assign new_P3_R1158_U290 = ~new_P3_R1158_U217 | ~new_P3_R1158_U8;
  assign new_P3_R1158_U291 = ~new_P3_U3074 | ~new_P3_R1158_U89;
  assign new_P3_R1158_U292 = ~new_P3_R1158_U132 | ~new_P3_R1158_U290;
  assign new_P3_R1158_U293 = ~new_P3_R1158_U503 | ~new_P3_R1158_U54;
  assign new_P3_R1158_U294 = ~new_P3_R1158_U497 | ~new_P3_R1158_U56;
  assign new_P3_R1158_U295 = ~new_P3_R1158_U131 | ~new_P3_R1158_U199;
  assign new_P3_R1158_U296 = ~new_P3_R1158_U294 | ~new_P3_R1158_U292;
  assign new_P3_R1158_U297 = ~new_P3_R1158_U196;
  assign new_P3_R1158_U298 = ~new_P3_R1158_U506 | ~new_P3_R1158_U57;
  assign new_P3_R1158_U299 = ~new_P3_R1158_U298 | ~new_P3_R1158_U196;
  assign new_P3_R1158_U300 = ~new_P3_U3060 | ~new_P3_R1158_U91;
  assign new_P3_R1158_U301 = ~new_P3_R1158_U194;
  assign new_P3_R1158_U302 = ~new_P3_R1158_U509 | ~new_P3_R1158_U58;
  assign new_P3_R1158_U303 = ~new_P3_R1158_U302 | ~new_P3_R1158_U194;
  assign new_P3_R1158_U304 = ~new_P3_U3065 | ~new_P3_R1158_U92;
  assign new_P3_R1158_U305 = ~new_P3_R1158_U192;
  assign new_P3_R1158_U306 = ~new_P3_R1158_U515 | ~new_P3_R1158_U38;
  assign new_P3_R1158_U307 = ~new_P3_R1158_U308 | ~new_P3_R1158_U60 | ~new_P3_R1158_U59;
  assign new_P3_R1158_U308 = ~new_P3_U3056 | ~new_P3_R1158_U78;
  assign new_P3_R1158_U309 = ~new_P3_R1158_U518 | ~new_P3_R1158_U39;
  assign new_P3_R1158_U310 = ~new_P3_R1158_U369 | ~new_P3_R1158_U192;
  assign new_P3_R1158_U311 = ~new_P3_R1158_U366 | ~new_P3_R1158_U307;
  assign new_P3_R1158_U312 = ~new_P3_R1158_U189;
  assign new_P3_R1158_U313 = ~new_P3_R1158_U467 | ~new_P3_R1158_U37;
  assign new_P3_R1158_U314 = ~new_P3_U3052 | ~new_P3_R1158_U75;
  assign new_P3_R1158_U315 = ~new_P3_U3052 | ~new_P3_R1158_U75;
  assign new_P3_R1158_U316 = ~new_P3_R1158_U467 | ~new_P3_R1158_U37;
  assign new_P3_R1158_U317 = ~new_P3_R1158_U190;
  assign new_P3_R1158_U318 = ~new_P3_R1158_U191;
  assign new_P3_R1158_U319 = ~new_P3_R1158_U138 | ~new_P3_R1158_U12;
  assign new_P3_R1158_U320 = ~new_P3_U3056 | ~new_P3_R1158_U78;
  assign new_P3_R1158_U321 = ~new_P3_R1158_U515 | ~new_P3_R1158_U38;
  assign new_P3_R1158_U322 = ~new_P3_R1158_U293 | ~new_P3_R1158_U199;
  assign new_P3_R1158_U323 = ~new_P3_R1158_U61;
  assign new_P3_R1158_U324 = ~new_P3_R1158_U500 | ~new_P3_R1158_U53;
  assign new_P3_R1158_U325 = ~new_P3_R1158_U324 | ~new_P3_R1158_U61;
  assign new_P3_R1158_U326 = ~new_P3_R1158_U143 | ~new_P3_R1158_U325;
  assign new_P3_R1158_U327 = ~new_P3_R1158_U323 | ~new_P3_R1158_U214;
  assign new_P3_R1158_U328 = ~new_P3_U3074 | ~new_P3_R1158_U89;
  assign new_P3_R1158_U329 = ~new_P3_R1158_U144 | ~new_P3_R1158_U327;
  assign new_P3_R1158_U330 = ~new_P3_R1158_U500 | ~new_P3_R1158_U53;
  assign new_P3_R1158_U331 = ~new_P3_R1158_U491 | ~new_P3_R1158_U41;
  assign new_P3_R1158_U332 = ~new_P3_R1158_U331 | ~new_P3_R1158_U62;
  assign new_P3_R1158_U333 = ~new_P3_R1158_U145 | ~new_P3_R1158_U332;
  assign new_P3_R1158_U334 = ~new_P3_R1158_U275 | ~new_P3_R1158_U42;
  assign new_P3_R1158_U335 = ~new_P3_U3068 | ~new_P3_R1158_U80;
  assign new_P3_R1158_U336 = ~new_P3_R1158_U146 | ~new_P3_R1158_U334;
  assign new_P3_R1158_U337 = ~new_P3_R1158_U491 | ~new_P3_R1158_U41;
  assign new_P3_R1158_U338 = ~new_P3_R1158_U267 | ~new_P3_R1158_U206;
  assign new_P3_R1158_U339 = ~new_P3_R1158_U64;
  assign new_P3_R1158_U340 = ~new_P3_R1158_U479 | ~new_P3_R1158_U45;
  assign new_P3_R1158_U341 = ~new_P3_R1158_U340 | ~new_P3_R1158_U64;
  assign new_P3_R1158_U342 = ~new_P3_R1158_U147 | ~new_P3_R1158_U341;
  assign new_P3_R1158_U343 = ~new_P3_R1158_U339 | ~new_P3_R1158_U213;
  assign new_P3_R1158_U344 = ~new_P3_U3079 | ~new_P3_R1158_U83;
  assign new_P3_R1158_U345 = ~new_P3_R1158_U148 | ~new_P3_R1158_U343;
  assign new_P3_R1158_U346 = ~new_P3_R1158_U479 | ~new_P3_R1158_U45;
  assign new_P3_R1158_U347 = ~new_P3_R1158_U250 | ~new_P3_R1158_U23;
  assign new_P3_R1158_U348 = ~new_P3_R1158_U257 | ~new_P3_R1158_U28;
  assign new_P3_R1158_U349 = ~new_P3_R1158_U321 | ~new_P3_R1158_U59;
  assign new_P3_R1158_U350 = ~new_P3_R1158_U309 | ~new_P3_R1158_U60;
  assign new_P3_R1158_U351 = ~new_P3_R1158_U330 | ~new_P3_R1158_U214;
  assign new_P3_R1158_U352 = ~new_P3_R1158_U293 | ~new_P3_R1158_U55;
  assign new_P3_R1158_U353 = ~new_P3_R1158_U337 | ~new_P3_R1158_U42;
  assign new_P3_R1158_U354 = ~new_P3_R1158_U346 | ~new_P3_R1158_U213;
  assign new_P3_R1158_U355 = ~new_P3_R1158_U267 | ~new_P3_R1158_U47;
  assign new_P3_R1158_U356 = ~new_P3_U3059 | ~new_P3_R1158_U74;
  assign new_P3_R1158_U357 = ~new_P3_U3082 | ~new_P3_R1158_U65;
  assign new_P3_R1158_U358 = ~new_P3_R1158_U133 | ~new_P3_R1158_U310;
  assign new_P3_R1158_U359 = ~new_P3_R1158_U68 | ~new_P3_R1158_U240;
  assign new_P3_R1158_U360 = ~new_P3_R1158_U223 | ~new_P3_U3076 | ~new_P3_R1158_U219;
  assign new_P3_R1158_U361 = ~new_P3_R1158_U119 | ~new_P3_R1158_U223;
  assign new_P3_R1158_U362 = ~new_P3_R1158_U236 | ~new_P3_R1158_U5;
  assign new_P3_R1158_U363 = ~new_P3_R1158_U34;
  assign new_P3_R1158_U364 = ~new_P3_R1158_U34 | ~new_P3_R1158_U242;
  assign new_P3_R1158_U365 = ~new_P3_R1158_U261 | ~new_P3_R1158_U9;
  assign new_P3_R1158_U366 = ~new_P3_R1158_U19 | ~new_P3_R1158_U367 | ~new_P3_R1158_U308;
  assign new_P3_R1158_U367 = ~new_P3_R1158_U78 | ~new_P3_R1158_U306;
  assign new_P3_R1158_U368 = ~new_P3_R1158_U19;
  assign new_P3_R1158_U369 = ~new_P3_R1158_U371 | ~new_P3_R1158_U370;
  assign new_P3_R1158_U370 = ~new_P3_R1158_U78 | ~new_P3_R1158_U309 | ~new_P3_R1158_U306;
  assign new_P3_R1158_U371 = ~new_P3_R1158_U368 | ~new_P3_R1158_U309;
  assign new_P3_R1158_U372 = ~new_P3_R1158_U63;
  assign new_P3_R1158_U373 = ~new_P3_R1158_U63 | ~new_P3_R1158_U270;
  assign new_P3_R1158_U374 = ~new_P3_R1158_U134 | ~new_P3_R1158_U366;
  assign new_P3_R1158_U375 = ~new_P3_R1158_U135 | ~new_P3_R1158_U192;
  assign new_P3_R1158_U376 = ~new_P3_R1158_U378 | ~new_P3_R1158_U377;
  assign new_P3_R1158_U377 = ~new_P3_R1158_U308 | ~new_P3_R1158_U60 | ~new_P3_R1158_U59;
  assign new_P3_R1158_U378 = ~new_P3_R1158_U19 | ~new_P3_R1158_U367 | ~new_P3_R1158_U308;
  assign new_P3_R1158_U379 = ~new_P3_R1158_U235 | ~new_P3_R1158_U165;
  assign new_P3_R1158_U380 = ~new_P3_R1158_U35;
  assign new_P3_R1158_U381 = ~new_P3_R1158_U10 | ~new_P3_R1158_U165;
  assign new_P3_R1158_U382 = ~new_P3_R1158_U163;
  assign new_P3_R1158_U383 = ~new_P3_R1158_U121 | ~new_P3_R1158_U165;
  assign new_P3_R1158_U384 = ~new_P3_R1158_U161;
  assign new_P3_R1158_U385 = ~new_P3_R1158_U260 | ~new_P3_R1158_U208;
  assign new_P3_R1158_U386 = ~new_P3_R1158_U206;
  assign new_P3_R1158_U387 = ~new_P3_R1158_U11 | ~new_P3_R1158_U208;
  assign new_P3_R1158_U388 = ~new_P3_R1158_U205;
  assign new_P3_R1158_U389 = ~new_P3_R1158_U128 | ~new_P3_R1158_U208;
  assign new_P3_R1158_U390 = ~new_P3_R1158_U203;
  assign new_P3_R1158_U391 = ~new_P3_R1158_U139 | ~new_P3_R1158_U209;
  assign new_P3_R1158_U392 = ~new_P3_R1158_U140 | ~new_P3_R1158_U209;
  assign new_P3_R1158_U393 = ~new_P3_U3152 | ~new_P3_R1158_U150;
  assign new_P3_R1158_U394 = ~new_P3_U3416 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U395 = ~new_P3_R1158_U65;
  assign new_P3_R1158_U396 = ~new_P3_R1158_U395 | ~new_P3_U3082;
  assign new_P3_R1158_U397 = ~new_P3_R1158_U65 | ~new_P3_R1158_U33;
  assign new_P3_R1158_U398 = ~new_P3_R1158_U395 | ~new_P3_U3082;
  assign new_P3_R1158_U399 = ~new_P3_R1158_U65 | ~new_P3_R1158_U33;
  assign new_P3_R1158_U400 = ~new_P3_R1158_U399 | ~new_P3_R1158_U398;
  assign new_P3_R1158_U401 = ~new_P3_U3152 | ~new_P3_R1158_U152;
  assign new_P3_R1158_U402 = ~new_P3_U3401 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U403 = ~new_P3_R1158_U74;
  assign new_P3_R1158_U404 = ~new_P3_U3152 | ~new_P3_R1158_U153;
  assign new_P3_R1158_U405 = ~new_P3_U3392 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U406 = ~new_P3_R1158_U72;
  assign new_P3_R1158_U407 = ~new_P3_U3152 | ~new_P3_R1158_U154;
  assign new_P3_R1158_U408 = ~new_P3_U3387 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U409 = ~new_P3_R1158_U73;
  assign new_P3_R1158_U410 = ~new_P3_U3152 | ~new_P3_R1158_U155;
  assign new_P3_R1158_U411 = ~new_P3_U3398 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U412 = ~new_P3_R1158_U71;
  assign new_P3_R1158_U413 = ~new_P3_U3152 | ~new_P3_R1158_U156;
  assign new_P3_R1158_U414 = ~new_P3_U3395 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U415 = ~new_P3_R1158_U70;
  assign new_P3_R1158_U416 = ~new_P3_U3152 | ~new_P3_R1158_U157;
  assign new_P3_R1158_U417 = ~new_P3_U3404 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U418 = ~new_P3_R1158_U69;
  assign new_P3_R1158_U419 = ~new_P3_U3152 | ~new_P3_R1158_U158;
  assign new_P3_R1158_U420 = ~new_P3_U3410 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U421 = ~new_P3_R1158_U68;
  assign new_P3_R1158_U422 = ~new_P3_U3152 | ~new_P3_R1158_U159;
  assign new_P3_R1158_U423 = ~new_P3_U3407 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U424 = ~new_P3_R1158_U67;
  assign new_P3_R1158_U425 = ~new_P3_U3152 | ~new_P3_R1158_U160;
  assign new_P3_R1158_U426 = ~new_P3_U3413 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U427 = ~new_P3_R1158_U66;
  assign new_P3_R1158_U428 = ~new_P3_R1158_U151 | ~new_P3_R1158_U161;
  assign new_P3_R1158_U429 = ~new_P3_R1158_U384 | ~new_P3_R1158_U400;
  assign new_P3_R1158_U430 = ~new_P3_R1158_U427 | ~new_P3_U3083;
  assign new_P3_R1158_U431 = ~new_P3_R1158_U66 | ~new_P3_R1158_U21;
  assign new_P3_R1158_U432 = ~new_P3_R1158_U427 | ~new_P3_U3083;
  assign new_P3_R1158_U433 = ~new_P3_R1158_U66 | ~new_P3_R1158_U21;
  assign new_P3_R1158_U434 = ~new_P3_R1158_U433 | ~new_P3_R1158_U432;
  assign new_P3_R1158_U435 = ~new_P3_R1158_U162 | ~new_P3_R1158_U163;
  assign new_P3_R1158_U436 = ~new_P3_R1158_U382 | ~new_P3_R1158_U434;
  assign new_P3_R1158_U437 = ~new_P3_R1158_U421 | ~new_P3_U3069;
  assign new_P3_R1158_U438 = ~new_P3_R1158_U68 | ~new_P3_R1158_U24;
  assign new_P3_R1158_U439 = ~new_P3_R1158_U424 | ~new_P3_U3070;
  assign new_P3_R1158_U440 = ~new_P3_R1158_U67 | ~new_P3_R1158_U22;
  assign new_P3_R1158_U441 = ~new_P3_R1158_U440 | ~new_P3_R1158_U439;
  assign new_P3_R1158_U442 = ~new_P3_R1158_U35 | ~new_P3_R1158_U347;
  assign new_P3_R1158_U443 = ~new_P3_R1158_U441 | ~new_P3_R1158_U380;
  assign new_P3_R1158_U444 = ~new_P3_R1158_U418 | ~new_P3_U3066;
  assign new_P3_R1158_U445 = ~new_P3_R1158_U69 | ~new_P3_R1158_U25;
  assign new_P3_R1158_U446 = ~new_P3_R1158_U418 | ~new_P3_U3066;
  assign new_P3_R1158_U447 = ~new_P3_R1158_U69 | ~new_P3_R1158_U25;
  assign new_P3_R1158_U448 = ~new_P3_R1158_U447 | ~new_P3_R1158_U446;
  assign new_P3_R1158_U449 = ~new_P3_R1158_U164 | ~new_P3_R1158_U165;
  assign new_P3_R1158_U450 = ~new_P3_R1158_U234 | ~new_P3_R1158_U448;
  assign new_P3_R1158_U451 = ~new_P3_R1158_U403 | ~new_P3_U3059;
  assign new_P3_R1158_U452 = ~new_P3_R1158_U74 | ~new_P3_R1158_U32;
  assign new_P3_R1158_U453 = ~new_P3_R1158_U403 | ~new_P3_U3059;
  assign new_P3_R1158_U454 = ~new_P3_R1158_U74 | ~new_P3_R1158_U32;
  assign new_P3_R1158_U455 = ~new_P3_R1158_U454 | ~new_P3_R1158_U453;
  assign new_P3_R1158_U456 = ~new_P3_R1158_U166 | ~new_P3_R1158_U167;
  assign new_P3_R1158_U457 = ~new_P3_R1158_U232 | ~new_P3_R1158_U455;
  assign new_P3_R1158_U458 = ~new_P3_R1158_U412 | ~new_P3_U3063;
  assign new_P3_R1158_U459 = ~new_P3_R1158_U71 | ~new_P3_R1158_U29;
  assign new_P3_R1158_U460 = ~new_P3_R1158_U415 | ~new_P3_U3067;
  assign new_P3_R1158_U461 = ~new_P3_R1158_U70 | ~new_P3_R1158_U27;
  assign new_P3_R1158_U462 = ~new_P3_R1158_U461 | ~new_P3_R1158_U460;
  assign new_P3_R1158_U463 = ~new_P3_R1158_U348 | ~new_P3_R1158_U36;
  assign new_P3_R1158_U464 = ~new_P3_R1158_U462 | ~new_P3_R1158_U225;
  assign new_P3_R1158_U465 = ~new_P3_U3152 | ~new_P3_R1158_U168;
  assign new_P3_R1158_U466 = ~new_P3_U3900 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U467 = ~new_P3_R1158_U75;
  assign new_P3_R1158_U468 = ~new_P3_U3152 | ~new_P3_R1158_U169;
  assign new_P3_R1158_U469 = ~new_P3_U3419 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U470 = ~new_P3_R1158_U85;
  assign new_P3_R1158_U471 = ~new_P3_U3152 | ~new_P3_R1158_U170;
  assign new_P3_R1158_U472 = ~new_P3_U3422 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U473 = ~new_P3_R1158_U84;
  assign new_P3_R1158_U474 = ~new_P3_U3152 | ~new_P3_R1158_U171;
  assign new_P3_R1158_U475 = ~new_P3_U3428 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U476 = ~new_P3_R1158_U83;
  assign new_P3_R1158_U477 = ~new_P3_U3152 | ~new_P3_R1158_U172;
  assign new_P3_R1158_U478 = ~new_P3_U3425 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U479 = ~new_P3_R1158_U82;
  assign new_P3_R1158_U480 = ~new_P3_U3152 | ~new_P3_R1158_U173;
  assign new_P3_R1158_U481 = ~new_P3_U3431 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U482 = ~new_P3_R1158_U81;
  assign new_P3_R1158_U483 = ~new_P3_U3152 | ~new_P3_R1158_U174;
  assign new_P3_R1158_U484 = ~new_P3_U3434 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U485 = ~new_P3_R1158_U86;
  assign new_P3_R1158_U486 = ~new_P3_U3152 | ~new_P3_R1158_U175;
  assign new_P3_R1158_U487 = ~new_P3_U3440 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U488 = ~new_P3_R1158_U80;
  assign new_P3_R1158_U489 = ~new_P3_U3152 | ~new_P3_R1158_U176;
  assign new_P3_R1158_U490 = ~new_P3_U3437 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U491 = ~new_P3_R1158_U79;
  assign new_P3_R1158_U492 = ~new_P3_U3152 | ~new_P3_R1158_U177;
  assign new_P3_R1158_U493 = ~new_P3_U3443 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U494 = ~new_P3_R1158_U87;
  assign new_P3_R1158_U495 = ~new_P3_U3152 | ~new_P3_R1158_U178;
  assign new_P3_R1158_U496 = ~new_P3_U3906 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U497 = ~new_P3_R1158_U89;
  assign new_P3_R1158_U498 = ~new_P3_U3152 | ~new_P3_R1158_U179;
  assign new_P3_R1158_U499 = ~new_P3_U3907 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U500 = ~new_P3_R1158_U90;
  assign new_P3_R1158_U501 = ~new_P3_U3152 | ~new_P3_R1158_U180;
  assign new_P3_R1158_U502 = ~new_P3_U3445 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U503 = ~new_P3_R1158_U88;
  assign new_P3_R1158_U504 = ~new_P3_U3152 | ~new_P3_R1158_U181;
  assign new_P3_R1158_U505 = ~new_P3_U3905 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U506 = ~new_P3_R1158_U91;
  assign new_P3_R1158_U507 = ~new_P3_U3152 | ~new_P3_R1158_U182;
  assign new_P3_R1158_U508 = ~new_P3_U3904 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U509 = ~new_P3_R1158_U92;
  assign new_P3_R1158_U510 = ~new_P3_U3152 | ~new_P3_R1158_U183;
  assign new_P3_R1158_U511 = ~new_P3_U3901 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U512 = ~new_P3_R1158_U78;
  assign new_P3_R1158_U513 = ~new_P3_U3152 | ~new_P3_R1158_U184;
  assign new_P3_R1158_U514 = ~new_P3_U3902 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U515 = ~new_P3_R1158_U76;
  assign new_P3_R1158_U516 = ~new_P3_U3152 | ~new_P3_R1158_U185;
  assign new_P3_R1158_U517 = ~new_P3_U3903 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U518 = ~new_P3_R1158_U77;
  assign new_P3_R1158_U519 = ~new_P3_U3152 | ~new_P3_R1158_U186;
  assign new_P3_R1158_U520 = ~new_P3_U3053 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U521 = ~new_P3_R1158_U137;
  assign new_P3_R1158_U522 = ~new_P3_U3899 | ~new_P3_R1158_U521;
  assign new_P3_R1158_U523 = ~new_P3_R1158_U137 | ~new_P3_R1158_U187;
  assign new_P3_R1158_U524 = ~new_P3_R1158_U93;
  assign new_P3_R1158_U525 = ~new_P3_R1158_U524 | ~new_P3_R1158_U358 | ~new_P3_R1158_U313;
  assign new_P3_R1158_U526 = ~new_P3_R1158_U93 | ~new_P3_R1158_U136 | ~new_P3_R1158_U375;
  assign new_P3_R1158_U527 = ~new_P3_R1158_U467 | ~new_P3_U3052;
  assign new_P3_R1158_U528 = ~new_P3_R1158_U75 | ~new_P3_R1158_U37;
  assign new_P3_R1158_U529 = ~new_P3_R1158_U467 | ~new_P3_U3052;
  assign new_P3_R1158_U530 = ~new_P3_R1158_U75 | ~new_P3_R1158_U37;
  assign new_P3_R1158_U531 = ~new_P3_R1158_U530 | ~new_P3_R1158_U529;
  assign new_P3_R1158_U532 = ~new_P3_R1158_U188 | ~new_P3_R1158_U189;
  assign new_P3_R1158_U533 = ~new_P3_R1158_U312 | ~new_P3_R1158_U531;
  assign new_P3_R1158_U534 = ~new_P3_R1158_U512 | ~new_P3_U3056;
  assign new_P3_R1158_U535 = ~new_P3_R1158_U78 | ~new_P3_R1158_U40;
  assign new_P3_R1158_U536 = ~new_P3_R1158_U104 | ~new_P3_R1158_U190;
  assign new_P3_R1158_U537 = ~new_P3_R1158_U103 | ~new_P3_R1158_U317;
  assign new_P3_R1158_U538 = ~new_P3_R1158_U515 | ~new_P3_U3057;
  assign new_P3_R1158_U539 = ~new_P3_R1158_U76 | ~new_P3_R1158_U38;
  assign new_P3_R1158_U540 = ~new_P3_R1158_U539 | ~new_P3_R1158_U538;
  assign new_P3_R1158_U541 = ~new_P3_R1158_U349 | ~new_P3_R1158_U191;
  assign new_P3_R1158_U542 = ~new_P3_R1158_U318 | ~new_P3_R1158_U540;
  assign new_P3_R1158_U543 = ~new_P3_R1158_U518 | ~new_P3_U3064;
  assign new_P3_R1158_U544 = ~new_P3_R1158_U77 | ~new_P3_R1158_U39;
  assign new_P3_R1158_U545 = ~new_P3_R1158_U544 | ~new_P3_R1158_U543;
  assign new_P3_R1158_U546 = ~new_P3_R1158_U350 | ~new_P3_R1158_U192;
  assign new_P3_R1158_U547 = ~new_P3_R1158_U305 | ~new_P3_R1158_U545;
  assign new_P3_R1158_U548 = ~new_P3_R1158_U509 | ~new_P3_U3065;
  assign new_P3_R1158_U549 = ~new_P3_R1158_U92 | ~new_P3_R1158_U58;
  assign new_P3_R1158_U550 = ~new_P3_R1158_U509 | ~new_P3_U3065;
  assign new_P3_R1158_U551 = ~new_P3_R1158_U92 | ~new_P3_R1158_U58;
  assign new_P3_R1158_U552 = ~new_P3_R1158_U551 | ~new_P3_R1158_U550;
  assign new_P3_R1158_U553 = ~new_P3_R1158_U193 | ~new_P3_R1158_U194;
  assign new_P3_R1158_U554 = ~new_P3_R1158_U301 | ~new_P3_R1158_U552;
  assign new_P3_R1158_U555 = ~new_P3_R1158_U506 | ~new_P3_U3060;
  assign new_P3_R1158_U556 = ~new_P3_R1158_U91 | ~new_P3_R1158_U57;
  assign new_P3_R1158_U557 = ~new_P3_R1158_U506 | ~new_P3_U3060;
  assign new_P3_R1158_U558 = ~new_P3_R1158_U91 | ~new_P3_R1158_U57;
  assign new_P3_R1158_U559 = ~new_P3_R1158_U558 | ~new_P3_R1158_U557;
  assign new_P3_R1158_U560 = ~new_P3_R1158_U195 | ~new_P3_R1158_U196;
  assign new_P3_R1158_U561 = ~new_P3_R1158_U297 | ~new_P3_R1158_U559;
  assign new_P3_R1158_U562 = ~new_P3_R1158_U497 | ~new_P3_U3074;
  assign new_P3_R1158_U563 = ~new_P3_R1158_U89 | ~new_P3_R1158_U56;
  assign new_P3_R1158_U564 = ~new_P3_R1158_U500 | ~new_P3_U3075;
  assign new_P3_R1158_U565 = ~new_P3_R1158_U90 | ~new_P3_R1158_U53;
  assign new_P3_R1158_U566 = ~new_P3_R1158_U565 | ~new_P3_R1158_U564;
  assign new_P3_R1158_U567 = ~new_P3_R1158_U351 | ~new_P3_R1158_U61;
  assign new_P3_R1158_U568 = ~new_P3_R1158_U566 | ~new_P3_R1158_U323;
  assign new_P3_R1158_U569 = ~new_P3_R1158_U406 | ~new_P3_U3077;
  assign new_P3_R1158_U570 = ~new_P3_R1158_U72 | ~new_P3_R1158_U30;
  assign new_P3_R1158_U571 = ~new_P3_R1158_U406 | ~new_P3_U3077;
  assign new_P3_R1158_U572 = ~new_P3_R1158_U72 | ~new_P3_R1158_U30;
  assign new_P3_R1158_U573 = ~new_P3_R1158_U572 | ~new_P3_R1158_U571;
  assign new_P3_R1158_U574 = ~new_P3_R1158_U197 | ~new_P3_R1158_U198;
  assign new_P3_R1158_U575 = ~new_P3_R1158_U222 | ~new_P3_R1158_U573;
  assign new_P3_R1158_U576 = ~new_P3_R1158_U503 | ~new_P3_U3080;
  assign new_P3_R1158_U577 = ~new_P3_R1158_U88 | ~new_P3_R1158_U54;
  assign new_P3_R1158_U578 = ~new_P3_R1158_U577 | ~new_P3_R1158_U576;
  assign new_P3_R1158_U579 = ~new_P3_R1158_U352 | ~new_P3_R1158_U199;
  assign new_P3_R1158_U580 = ~new_P3_R1158_U287 | ~new_P3_R1158_U578;
  assign new_P3_R1158_U581 = ~new_P3_R1158_U494 | ~new_P3_U3081;
  assign new_P3_R1158_U582 = ~new_P3_R1158_U87 | ~new_P3_R1158_U52;
  assign new_P3_R1158_U583 = ~new_P3_R1158_U494 | ~new_P3_U3081;
  assign new_P3_R1158_U584 = ~new_P3_R1158_U87 | ~new_P3_R1158_U52;
  assign new_P3_R1158_U585 = ~new_P3_R1158_U584 | ~new_P3_R1158_U583;
  assign new_P3_R1158_U586 = ~new_P3_R1158_U200 | ~new_P3_R1158_U201;
  assign new_P3_R1158_U587 = ~new_P3_R1158_U283 | ~new_P3_R1158_U585;
  assign new_P3_R1158_U588 = ~new_P3_R1158_U488 | ~new_P3_U3068;
  assign new_P3_R1158_U589 = ~new_P3_R1158_U80 | ~new_P3_R1158_U43;
  assign new_P3_R1158_U590 = ~new_P3_R1158_U491 | ~new_P3_U3072;
  assign new_P3_R1158_U591 = ~new_P3_R1158_U79 | ~new_P3_R1158_U41;
  assign new_P3_R1158_U592 = ~new_P3_R1158_U591 | ~new_P3_R1158_U590;
  assign new_P3_R1158_U593 = ~new_P3_R1158_U353 | ~new_P3_R1158_U62;
  assign new_P3_R1158_U594 = ~new_P3_R1158_U592 | ~new_P3_R1158_U275;
  assign new_P3_R1158_U595 = ~new_P3_R1158_U485 | ~new_P3_U3073;
  assign new_P3_R1158_U596 = ~new_P3_R1158_U86 | ~new_P3_R1158_U51;
  assign new_P3_R1158_U597 = ~new_P3_R1158_U485 | ~new_P3_U3073;
  assign new_P3_R1158_U598 = ~new_P3_R1158_U86 | ~new_P3_R1158_U51;
  assign new_P3_R1158_U599 = ~new_P3_R1158_U598 | ~new_P3_R1158_U597;
  assign new_P3_R1158_U600 = ~new_P3_R1158_U202 | ~new_P3_R1158_U203;
  assign new_P3_R1158_U601 = ~new_P3_R1158_U390 | ~new_P3_R1158_U599;
  assign new_P3_R1158_U602 = ~new_P3_R1158_U482 | ~new_P3_U3078;
  assign new_P3_R1158_U603 = ~new_P3_R1158_U81 | ~new_P3_R1158_U44;
  assign new_P3_R1158_U604 = ~new_P3_R1158_U482 | ~new_P3_U3078;
  assign new_P3_R1158_U605 = ~new_P3_R1158_U81 | ~new_P3_R1158_U44;
  assign new_P3_R1158_U606 = ~new_P3_R1158_U605 | ~new_P3_R1158_U604;
  assign new_P3_R1158_U607 = ~new_P3_R1158_U204 | ~new_P3_R1158_U205;
  assign new_P3_R1158_U608 = ~new_P3_R1158_U388 | ~new_P3_R1158_U606;
  assign new_P3_R1158_U609 = ~new_P3_R1158_U476 | ~new_P3_U3079;
  assign new_P3_R1158_U610 = ~new_P3_R1158_U83 | ~new_P3_R1158_U48;
  assign new_P3_R1158_U611 = ~new_P3_R1158_U479 | ~new_P3_U3071;
  assign new_P3_R1158_U612 = ~new_P3_R1158_U82 | ~new_P3_R1158_U45;
  assign new_P3_R1158_U613 = ~new_P3_R1158_U612 | ~new_P3_R1158_U611;
  assign new_P3_R1158_U614 = ~new_P3_R1158_U354 | ~new_P3_R1158_U64;
  assign new_P3_R1158_U615 = ~new_P3_R1158_U613 | ~new_P3_R1158_U339;
  assign new_P3_R1158_U616 = ~new_P3_R1158_U473 | ~new_P3_U3062;
  assign new_P3_R1158_U617 = ~new_P3_R1158_U84 | ~new_P3_R1158_U46;
  assign new_P3_R1158_U618 = ~new_P3_R1158_U617 | ~new_P3_R1158_U616;
  assign new_P3_R1158_U619 = ~new_P3_R1158_U206 | ~new_P3_R1158_U355;
  assign new_P3_R1158_U620 = ~new_P3_R1158_U386 | ~new_P3_R1158_U618;
  assign new_P3_R1158_U621 = ~new_P3_R1158_U470 | ~new_P3_U3061;
  assign new_P3_R1158_U622 = ~new_P3_R1158_U85 | ~new_P3_R1158_U49;
  assign new_P3_R1158_U623 = ~new_P3_R1158_U470 | ~new_P3_U3061;
  assign new_P3_R1158_U624 = ~new_P3_R1158_U85 | ~new_P3_R1158_U49;
  assign new_P3_R1158_U625 = ~new_P3_R1158_U624 | ~new_P3_R1158_U623;
  assign new_P3_R1158_U626 = ~new_P3_R1158_U207 | ~new_P3_R1158_U208;
  assign new_P3_R1158_U627 = ~new_P3_R1158_U259 | ~new_P3_R1158_U625;
  assign new_P3_R1158_U628 = ~new_P3_R1158_U73 | ~new_P3_R1158_U20;
  assign new_P3_R1158_U629 = ~new_P3_R1158_U409 | ~new_P3_U3152;
  assign new_P3_R1158_U630 = ~new_P3_R1158_U149;
  assign new_P3_R1158_U631 = ~new_P3_R1158_U630 | ~new_P3_U3076;
  assign new_P3_R1158_U632 = ~new_P3_R1158_U149 | ~new_P3_R1158_U31;
  assign new_P3_R1131_U6 = new_P3_R1131_U210 & new_P3_R1131_U209;
  assign new_P3_R1131_U7 = new_P3_R1131_U189 & new_P3_R1131_U245;
  assign new_P3_R1131_U8 = new_P3_R1131_U247 & new_P3_R1131_U246;
  assign new_P3_R1131_U9 = new_P3_R1131_U190 & new_P3_R1131_U262;
  assign new_P3_R1131_U10 = new_P3_R1131_U264 & new_P3_R1131_U263;
  assign new_P3_R1131_U11 = new_P3_R1131_U191 & new_P3_R1131_U286;
  assign new_P3_R1131_U12 = new_P3_R1131_U288 & new_P3_R1131_U287;
  assign new_P3_R1131_U13 = new_P3_R1131_U213 & new_P3_R1131_U208 & new_P3_R1131_U194;
  assign new_P3_R1131_U14 = new_P3_R1131_U218 & new_P3_R1131_U195;
  assign new_P3_R1131_U15 = new_P3_R1131_U392 & new_P3_R1131_U391;
  assign new_P3_R1131_U16 = ~new_P3_R1131_U342 | ~new_P3_R1131_U345;
  assign new_P3_R1131_U17 = ~new_P3_R1131_U331 | ~new_P3_R1131_U334;
  assign new_P3_R1131_U18 = ~new_P3_R1131_U320 | ~new_P3_R1131_U323;
  assign new_P3_R1131_U19 = ~new_P3_R1131_U312 | ~new_P3_R1131_U314;
  assign new_P3_R1131_U20 = ~new_P3_R1131_U351 | ~new_P3_R1131_U162 | ~new_P3_R1131_U183;
  assign new_P3_R1131_U21 = ~new_P3_R1131_U241 | ~new_P3_R1131_U243;
  assign new_P3_R1131_U22 = ~new_P3_R1131_U233 | ~new_P3_R1131_U236;
  assign new_P3_R1131_U23 = ~new_P3_R1131_U225 | ~new_P3_R1131_U227;
  assign new_P3_R1131_U24 = ~new_P3_R1131_U172 | ~new_P3_R1131_U348;
  assign new_P3_R1131_U25 = ~new_P3_U3069;
  assign new_P3_R1131_U26 = ~new_P3_U3069 | ~new_P3_R1131_U39;
  assign new_P3_R1131_U27 = ~new_P3_U3083;
  assign new_P3_R1131_U28 = ~new_P3_U3413;
  assign new_P3_R1131_U29 = ~new_P3_U3395;
  assign new_P3_R1131_U30 = ~new_P3_U3387;
  assign new_P3_R1131_U31 = ~new_P3_U3077;
  assign new_P3_R1131_U32 = ~new_P3_U3398;
  assign new_P3_R1131_U33 = ~new_P3_U3067;
  assign new_P3_R1131_U34 = ~new_P3_U3067 | ~new_P3_R1131_U29;
  assign new_P3_R1131_U35 = ~new_P3_U3063;
  assign new_P3_R1131_U36 = ~new_P3_U3404;
  assign new_P3_R1131_U37 = ~new_P3_U3407;
  assign new_P3_R1131_U38 = ~new_P3_U3401;
  assign new_P3_R1131_U39 = ~new_P3_U3410;
  assign new_P3_R1131_U40 = ~new_P3_U3070;
  assign new_P3_R1131_U41 = ~new_P3_U3066;
  assign new_P3_R1131_U42 = ~new_P3_U3059;
  assign new_P3_R1131_U43 = ~new_P3_U3059 | ~new_P3_R1131_U38;
  assign new_P3_R1131_U44 = ~new_P3_R1131_U214 | ~new_P3_R1131_U212;
  assign new_P3_R1131_U45 = ~new_P3_U3416;
  assign new_P3_R1131_U46 = ~new_P3_U3082;
  assign new_P3_R1131_U47 = ~new_P3_R1131_U44 | ~new_P3_R1131_U215;
  assign new_P3_R1131_U48 = ~new_P3_R1131_U43 | ~new_P3_R1131_U229;
  assign new_P3_R1131_U49 = ~new_P3_R1131_U349 | ~new_P3_R1131_U201 | ~new_P3_R1131_U185;
  assign new_P3_R1131_U50 = ~new_P3_U3901;
  assign new_P3_R1131_U51 = ~new_P3_U3422;
  assign new_P3_R1131_U52 = ~new_P3_U3419;
  assign new_P3_R1131_U53 = ~new_P3_U3062;
  assign new_P3_R1131_U54 = ~new_P3_U3061;
  assign new_P3_R1131_U55 = ~new_P3_U3082 | ~new_P3_R1131_U45;
  assign new_P3_R1131_U56 = ~new_P3_U3425;
  assign new_P3_R1131_U57 = ~new_P3_U3071;
  assign new_P3_R1131_U58 = ~new_P3_U3428;
  assign new_P3_R1131_U59 = ~new_P3_U3079;
  assign new_P3_R1131_U60 = ~new_P3_U3437;
  assign new_P3_R1131_U61 = ~new_P3_U3434;
  assign new_P3_R1131_U62 = ~new_P3_U3431;
  assign new_P3_R1131_U63 = ~new_P3_U3072;
  assign new_P3_R1131_U64 = ~new_P3_U3073;
  assign new_P3_R1131_U65 = ~new_P3_U3078;
  assign new_P3_R1131_U66 = ~new_P3_U3078 | ~new_P3_R1131_U62;
  assign new_P3_R1131_U67 = ~new_P3_U3440;
  assign new_P3_R1131_U68 = ~new_P3_U3068;
  assign new_P3_R1131_U69 = ~new_P3_U3081;
  assign new_P3_R1131_U70 = ~new_P3_U3445;
  assign new_P3_R1131_U71 = ~new_P3_U3080;
  assign new_P3_R1131_U72 = ~new_P3_U3907;
  assign new_P3_R1131_U73 = ~new_P3_U3075;
  assign new_P3_R1131_U74 = ~new_P3_U3904;
  assign new_P3_R1131_U75 = ~new_P3_U3905;
  assign new_P3_R1131_U76 = ~new_P3_U3906;
  assign new_P3_R1131_U77 = ~new_P3_U3065;
  assign new_P3_R1131_U78 = ~new_P3_U3060;
  assign new_P3_R1131_U79 = ~new_P3_U3074;
  assign new_P3_R1131_U80 = ~new_P3_U3074 | ~new_P3_R1131_U76;
  assign new_P3_R1131_U81 = ~new_P3_U3903;
  assign new_P3_R1131_U82 = ~new_P3_U3064;
  assign new_P3_R1131_U83 = ~new_P3_U3902;
  assign new_P3_R1131_U84 = ~new_P3_U3057;
  assign new_P3_R1131_U85 = ~new_P3_U3900;
  assign new_P3_R1131_U86 = ~new_P3_U3056;
  assign new_P3_R1131_U87 = ~new_P3_U3056 | ~new_P3_R1131_U50;
  assign new_P3_R1131_U88 = ~new_P3_U3052;
  assign new_P3_R1131_U89 = ~new_P3_U3899;
  assign new_P3_R1131_U90 = ~new_P3_U3053;
  assign new_P3_R1131_U91 = ~new_P3_R1131_U302 | ~new_P3_R1131_U301;
  assign new_P3_R1131_U92 = ~new_P3_R1131_U80 | ~new_P3_R1131_U316;
  assign new_P3_R1131_U93 = ~new_P3_R1131_U66 | ~new_P3_R1131_U327;
  assign new_P3_R1131_U94 = ~new_P3_R1131_U55 | ~new_P3_R1131_U338;
  assign new_P3_R1131_U95 = ~new_P3_U3076;
  assign new_P3_R1131_U96 = ~new_P3_R1131_U402 | ~new_P3_R1131_U401;
  assign new_P3_R1131_U97 = ~new_P3_R1131_U416 | ~new_P3_R1131_U415;
  assign new_P3_R1131_U98 = ~new_P3_R1131_U421 | ~new_P3_R1131_U420;
  assign new_P3_R1131_U99 = ~new_P3_R1131_U437 | ~new_P3_R1131_U436;
  assign new_P3_R1131_U100 = ~new_P3_R1131_U442 | ~new_P3_R1131_U441;
  assign new_P3_R1131_U101 = ~new_P3_R1131_U447 | ~new_P3_R1131_U446;
  assign new_P3_R1131_U102 = ~new_P3_R1131_U452 | ~new_P3_R1131_U451;
  assign new_P3_R1131_U103 = ~new_P3_R1131_U457 | ~new_P3_R1131_U456;
  assign new_P3_R1131_U104 = ~new_P3_R1131_U473 | ~new_P3_R1131_U472;
  assign new_P3_R1131_U105 = ~new_P3_R1131_U478 | ~new_P3_R1131_U477;
  assign new_P3_R1131_U106 = ~new_P3_R1131_U361 | ~new_P3_R1131_U360;
  assign new_P3_R1131_U107 = ~new_P3_R1131_U370 | ~new_P3_R1131_U369;
  assign new_P3_R1131_U108 = ~new_P3_R1131_U377 | ~new_P3_R1131_U376;
  assign new_P3_R1131_U109 = ~new_P3_R1131_U381 | ~new_P3_R1131_U380;
  assign new_P3_R1131_U110 = ~new_P3_R1131_U390 | ~new_P3_R1131_U389;
  assign new_P3_R1131_U111 = ~new_P3_R1131_U411 | ~new_P3_R1131_U410;
  assign new_P3_R1131_U112 = ~new_P3_R1131_U428 | ~new_P3_R1131_U427;
  assign new_P3_R1131_U113 = ~new_P3_R1131_U432 | ~new_P3_R1131_U431;
  assign new_P3_R1131_U114 = ~new_P3_R1131_U464 | ~new_P3_R1131_U463;
  assign new_P3_R1131_U115 = ~new_P3_R1131_U468 | ~new_P3_R1131_U467;
  assign new_P3_R1131_U116 = ~new_P3_R1131_U485 | ~new_P3_R1131_U484;
  assign new_P3_R1131_U117 = new_P3_R1131_U352 & new_P3_R1131_U193;
  assign new_P3_R1131_U118 = new_P3_R1131_U205 & new_P3_R1131_U206;
  assign new_P3_R1131_U119 = new_P3_R1131_U14 & new_P3_R1131_U13;
  assign new_P3_R1131_U120 = new_P3_R1131_U357 & new_P3_R1131_U354;
  assign new_P3_R1131_U121 = new_P3_R1131_U26 & new_P3_R1131_U363 & new_P3_R1131_U362;
  assign new_P3_R1131_U122 = new_P3_R1131_U366 & new_P3_R1131_U195;
  assign new_P3_R1131_U123 = new_P3_R1131_U235 & new_P3_R1131_U6;
  assign new_P3_R1131_U124 = new_P3_R1131_U373 & new_P3_R1131_U194;
  assign new_P3_R1131_U125 = new_P3_R1131_U34 & new_P3_R1131_U383 & new_P3_R1131_U382;
  assign new_P3_R1131_U126 = new_P3_R1131_U386 & new_P3_R1131_U193;
  assign new_P3_R1131_U127 = new_P3_R1131_U222 & new_P3_R1131_U7;
  assign new_P3_R1131_U128 = new_P3_R1131_U267 & new_P3_R1131_U9;
  assign new_P3_R1131_U129 = new_P3_R1131_U291 & new_P3_R1131_U11;
  assign new_P3_R1131_U130 = new_P3_R1131_U355 & new_P3_R1131_U192;
  assign new_P3_R1131_U131 = new_P3_R1131_U306 & new_P3_R1131_U307;
  assign new_P3_R1131_U132 = new_P3_R1131_U309 & new_P3_R1131_U395;
  assign new_P3_R1131_U133 = new_P3_R1131_U306 & new_P3_R1131_U307;
  assign new_P3_R1131_U134 = new_P3_R1131_U15 & new_P3_R1131_U310;
  assign new_P3_R1131_U135 = ~new_P3_R1131_U399 | ~new_P3_R1131_U398;
  assign new_P3_R1131_U136 = new_P3_R1131_U87 & new_P3_R1131_U404 & new_P3_R1131_U403;
  assign new_P3_R1131_U137 = new_P3_R1131_U407 & new_P3_R1131_U192;
  assign new_P3_R1131_U138 = ~new_P3_R1131_U413 | ~new_P3_R1131_U412;
  assign new_P3_R1131_U139 = ~new_P3_R1131_U418 | ~new_P3_R1131_U417;
  assign new_P3_R1131_U140 = new_P3_R1131_U322 & new_P3_R1131_U12;
  assign new_P3_R1131_U141 = new_P3_R1131_U424 & new_P3_R1131_U191;
  assign new_P3_R1131_U142 = ~new_P3_R1131_U434 | ~new_P3_R1131_U433;
  assign new_P3_R1131_U143 = ~new_P3_R1131_U439 | ~new_P3_R1131_U438;
  assign new_P3_R1131_U144 = ~new_P3_R1131_U444 | ~new_P3_R1131_U443;
  assign new_P3_R1131_U145 = ~new_P3_R1131_U449 | ~new_P3_R1131_U448;
  assign new_P3_R1131_U146 = ~new_P3_R1131_U454 | ~new_P3_R1131_U453;
  assign new_P3_R1131_U147 = new_P3_R1131_U333 & new_P3_R1131_U10;
  assign new_P3_R1131_U148 = new_P3_R1131_U460 & new_P3_R1131_U190;
  assign new_P3_R1131_U149 = ~new_P3_R1131_U470 | ~new_P3_R1131_U469;
  assign new_P3_R1131_U150 = ~new_P3_R1131_U475 | ~new_P3_R1131_U474;
  assign new_P3_R1131_U151 = new_P3_R1131_U344 & new_P3_R1131_U8;
  assign new_P3_R1131_U152 = new_P3_R1131_U481 & new_P3_R1131_U189;
  assign new_P3_R1131_U153 = new_P3_R1131_U359 & new_P3_R1131_U358;
  assign new_P3_R1131_U154 = ~new_P3_R1131_U120 | ~new_P3_R1131_U356;
  assign new_P3_R1131_U155 = new_P3_R1131_U368 & new_P3_R1131_U367;
  assign new_P3_R1131_U156 = new_P3_R1131_U375 & new_P3_R1131_U374;
  assign new_P3_R1131_U157 = new_P3_R1131_U379 & new_P3_R1131_U378;
  assign new_P3_R1131_U158 = ~new_P3_R1131_U118 | ~new_P3_R1131_U203;
  assign new_P3_R1131_U159 = new_P3_R1131_U388 & new_P3_R1131_U387;
  assign new_P3_R1131_U160 = ~new_P3_U3908;
  assign new_P3_R1131_U161 = ~new_P3_U3054;
  assign new_P3_R1131_U162 = new_P3_R1131_U397 & new_P3_R1131_U396;
  assign new_P3_R1131_U163 = ~new_P3_R1131_U131 | ~new_P3_R1131_U304;
  assign new_P3_R1131_U164 = new_P3_R1131_U409 & new_P3_R1131_U408;
  assign new_P3_R1131_U165 = ~new_P3_R1131_U298 | ~new_P3_R1131_U297;
  assign new_P3_R1131_U166 = ~new_P3_R1131_U294 | ~new_P3_R1131_U293;
  assign new_P3_R1131_U167 = new_P3_R1131_U426 & new_P3_R1131_U425;
  assign new_P3_R1131_U168 = new_P3_R1131_U430 & new_P3_R1131_U429;
  assign new_P3_R1131_U169 = ~new_P3_R1131_U284 | ~new_P3_R1131_U283;
  assign new_P3_R1131_U170 = ~new_P3_R1131_U280 | ~new_P3_R1131_U279;
  assign new_P3_R1131_U171 = ~new_P3_U3392;
  assign new_P3_R1131_U172 = ~new_P3_U3387 | ~new_P3_R1131_U95;
  assign new_P3_R1131_U173 = ~new_P3_R1131_U350 | ~new_P3_R1131_U276 | ~new_P3_R1131_U184;
  assign new_P3_R1131_U174 = ~new_P3_U3443;
  assign new_P3_R1131_U175 = ~new_P3_R1131_U274 | ~new_P3_R1131_U273;
  assign new_P3_R1131_U176 = ~new_P3_R1131_U270 | ~new_P3_R1131_U269;
  assign new_P3_R1131_U177 = new_P3_R1131_U462 & new_P3_R1131_U461;
  assign new_P3_R1131_U178 = new_P3_R1131_U466 & new_P3_R1131_U465;
  assign new_P3_R1131_U179 = ~new_P3_R1131_U260 | ~new_P3_R1131_U259;
  assign new_P3_R1131_U180 = ~new_P3_R1131_U256 | ~new_P3_R1131_U255;
  assign new_P3_R1131_U181 = ~new_P3_R1131_U252 | ~new_P3_R1131_U251;
  assign new_P3_R1131_U182 = new_P3_R1131_U483 & new_P3_R1131_U482;
  assign new_P3_R1131_U183 = ~new_P3_R1131_U132 | ~new_P3_R1131_U163;
  assign new_P3_R1131_U184 = ~new_P3_R1131_U175 | ~new_P3_R1131_U174;
  assign new_P3_R1131_U185 = ~new_P3_R1131_U172 | ~new_P3_R1131_U171;
  assign new_P3_R1131_U186 = ~new_P3_R1131_U87;
  assign new_P3_R1131_U187 = ~new_P3_R1131_U34;
  assign new_P3_R1131_U188 = ~new_P3_R1131_U26;
  assign new_P3_R1131_U189 = ~new_P3_U3419 | ~new_P3_R1131_U54;
  assign new_P3_R1131_U190 = ~new_P3_U3434 | ~new_P3_R1131_U64;
  assign new_P3_R1131_U191 = ~new_P3_U3905 | ~new_P3_R1131_U78;
  assign new_P3_R1131_U192 = ~new_P3_U3901 | ~new_P3_R1131_U86;
  assign new_P3_R1131_U193 = ~new_P3_U3395 | ~new_P3_R1131_U33;
  assign new_P3_R1131_U194 = ~new_P3_U3404 | ~new_P3_R1131_U41;
  assign new_P3_R1131_U195 = ~new_P3_U3410 | ~new_P3_R1131_U25;
  assign new_P3_R1131_U196 = ~new_P3_R1131_U66;
  assign new_P3_R1131_U197 = ~new_P3_R1131_U80;
  assign new_P3_R1131_U198 = ~new_P3_R1131_U43;
  assign new_P3_R1131_U199 = ~new_P3_R1131_U55;
  assign new_P3_R1131_U200 = ~new_P3_R1131_U172;
  assign new_P3_R1131_U201 = ~new_P3_U3077 | ~new_P3_R1131_U172;
  assign new_P3_R1131_U202 = ~new_P3_R1131_U49;
  assign new_P3_R1131_U203 = ~new_P3_R1131_U117 | ~new_P3_R1131_U49;
  assign new_P3_R1131_U204 = ~new_P3_R1131_U35 | ~new_P3_R1131_U34;
  assign new_P3_R1131_U205 = ~new_P3_R1131_U204 | ~new_P3_R1131_U32;
  assign new_P3_R1131_U206 = ~new_P3_U3063 | ~new_P3_R1131_U187;
  assign new_P3_R1131_U207 = ~new_P3_R1131_U158;
  assign new_P3_R1131_U208 = ~new_P3_U3407 | ~new_P3_R1131_U40;
  assign new_P3_R1131_U209 = ~new_P3_U3070 | ~new_P3_R1131_U37;
  assign new_P3_R1131_U210 = ~new_P3_U3066 | ~new_P3_R1131_U36;
  assign new_P3_R1131_U211 = ~new_P3_R1131_U198 | ~new_P3_R1131_U194;
  assign new_P3_R1131_U212 = ~new_P3_R1131_U6 | ~new_P3_R1131_U211;
  assign new_P3_R1131_U213 = ~new_P3_U3401 | ~new_P3_R1131_U42;
  assign new_P3_R1131_U214 = ~new_P3_U3407 | ~new_P3_R1131_U40;
  assign new_P3_R1131_U215 = ~new_P3_R1131_U13 | ~new_P3_R1131_U158;
  assign new_P3_R1131_U216 = ~new_P3_R1131_U44;
  assign new_P3_R1131_U217 = ~new_P3_R1131_U47;
  assign new_P3_R1131_U218 = ~new_P3_U3413 | ~new_P3_R1131_U27;
  assign new_P3_R1131_U219 = ~new_P3_R1131_U27 | ~new_P3_R1131_U26;
  assign new_P3_R1131_U220 = ~new_P3_U3083 | ~new_P3_R1131_U188;
  assign new_P3_R1131_U221 = ~new_P3_R1131_U154;
  assign new_P3_R1131_U222 = ~new_P3_U3416 | ~new_P3_R1131_U46;
  assign new_P3_R1131_U223 = ~new_P3_R1131_U222 | ~new_P3_R1131_U55;
  assign new_P3_R1131_U224 = ~new_P3_R1131_U217 | ~new_P3_R1131_U26;
  assign new_P3_R1131_U225 = ~new_P3_R1131_U122 | ~new_P3_R1131_U224;
  assign new_P3_R1131_U226 = ~new_P3_R1131_U47 | ~new_P3_R1131_U195;
  assign new_P3_R1131_U227 = ~new_P3_R1131_U121 | ~new_P3_R1131_U226;
  assign new_P3_R1131_U228 = ~new_P3_R1131_U26 | ~new_P3_R1131_U195;
  assign new_P3_R1131_U229 = ~new_P3_R1131_U213 | ~new_P3_R1131_U158;
  assign new_P3_R1131_U230 = ~new_P3_R1131_U48;
  assign new_P3_R1131_U231 = ~new_P3_U3066 | ~new_P3_R1131_U36;
  assign new_P3_R1131_U232 = ~new_P3_R1131_U230 | ~new_P3_R1131_U231;
  assign new_P3_R1131_U233 = ~new_P3_R1131_U124 | ~new_P3_R1131_U232;
  assign new_P3_R1131_U234 = ~new_P3_R1131_U48 | ~new_P3_R1131_U194;
  assign new_P3_R1131_U235 = ~new_P3_U3407 | ~new_P3_R1131_U40;
  assign new_P3_R1131_U236 = ~new_P3_R1131_U123 | ~new_P3_R1131_U234;
  assign new_P3_R1131_U237 = ~new_P3_U3066 | ~new_P3_R1131_U36;
  assign new_P3_R1131_U238 = ~new_P3_R1131_U194 | ~new_P3_R1131_U237;
  assign new_P3_R1131_U239 = ~new_P3_R1131_U213 | ~new_P3_R1131_U43;
  assign new_P3_R1131_U240 = ~new_P3_R1131_U202 | ~new_P3_R1131_U34;
  assign new_P3_R1131_U241 = ~new_P3_R1131_U126 | ~new_P3_R1131_U240;
  assign new_P3_R1131_U242 = ~new_P3_R1131_U49 | ~new_P3_R1131_U193;
  assign new_P3_R1131_U243 = ~new_P3_R1131_U125 | ~new_P3_R1131_U242;
  assign new_P3_R1131_U244 = ~new_P3_R1131_U193 | ~new_P3_R1131_U34;
  assign new_P3_R1131_U245 = ~new_P3_U3422 | ~new_P3_R1131_U53;
  assign new_P3_R1131_U246 = ~new_P3_U3062 | ~new_P3_R1131_U51;
  assign new_P3_R1131_U247 = ~new_P3_U3061 | ~new_P3_R1131_U52;
  assign new_P3_R1131_U248 = ~new_P3_R1131_U199 | ~new_P3_R1131_U7;
  assign new_P3_R1131_U249 = ~new_P3_R1131_U8 | ~new_P3_R1131_U248;
  assign new_P3_R1131_U250 = ~new_P3_U3422 | ~new_P3_R1131_U53;
  assign new_P3_R1131_U251 = ~new_P3_R1131_U127 | ~new_P3_R1131_U154;
  assign new_P3_R1131_U252 = ~new_P3_R1131_U250 | ~new_P3_R1131_U249;
  assign new_P3_R1131_U253 = ~new_P3_R1131_U181;
  assign new_P3_R1131_U254 = ~new_P3_U3425 | ~new_P3_R1131_U57;
  assign new_P3_R1131_U255 = ~new_P3_R1131_U254 | ~new_P3_R1131_U181;
  assign new_P3_R1131_U256 = ~new_P3_U3071 | ~new_P3_R1131_U56;
  assign new_P3_R1131_U257 = ~new_P3_R1131_U180;
  assign new_P3_R1131_U258 = ~new_P3_U3428 | ~new_P3_R1131_U59;
  assign new_P3_R1131_U259 = ~new_P3_R1131_U258 | ~new_P3_R1131_U180;
  assign new_P3_R1131_U260 = ~new_P3_U3079 | ~new_P3_R1131_U58;
  assign new_P3_R1131_U261 = ~new_P3_R1131_U179;
  assign new_P3_R1131_U262 = ~new_P3_U3437 | ~new_P3_R1131_U63;
  assign new_P3_R1131_U263 = ~new_P3_U3072 | ~new_P3_R1131_U60;
  assign new_P3_R1131_U264 = ~new_P3_U3073 | ~new_P3_R1131_U61;
  assign new_P3_R1131_U265 = ~new_P3_R1131_U196 | ~new_P3_R1131_U9;
  assign new_P3_R1131_U266 = ~new_P3_R1131_U10 | ~new_P3_R1131_U265;
  assign new_P3_R1131_U267 = ~new_P3_U3431 | ~new_P3_R1131_U65;
  assign new_P3_R1131_U268 = ~new_P3_U3437 | ~new_P3_R1131_U63;
  assign new_P3_R1131_U269 = ~new_P3_R1131_U128 | ~new_P3_R1131_U179;
  assign new_P3_R1131_U270 = ~new_P3_R1131_U268 | ~new_P3_R1131_U266;
  assign new_P3_R1131_U271 = ~new_P3_R1131_U176;
  assign new_P3_R1131_U272 = ~new_P3_U3440 | ~new_P3_R1131_U68;
  assign new_P3_R1131_U273 = ~new_P3_R1131_U272 | ~new_P3_R1131_U176;
  assign new_P3_R1131_U274 = ~new_P3_U3068 | ~new_P3_R1131_U67;
  assign new_P3_R1131_U275 = ~new_P3_R1131_U175;
  assign new_P3_R1131_U276 = ~new_P3_U3081 | ~new_P3_R1131_U175;
  assign new_P3_R1131_U277 = ~new_P3_R1131_U173;
  assign new_P3_R1131_U278 = ~new_P3_U3445 | ~new_P3_R1131_U71;
  assign new_P3_R1131_U279 = ~new_P3_R1131_U278 | ~new_P3_R1131_U173;
  assign new_P3_R1131_U280 = ~new_P3_U3080 | ~new_P3_R1131_U70;
  assign new_P3_R1131_U281 = ~new_P3_R1131_U170;
  assign new_P3_R1131_U282 = ~new_P3_U3907 | ~new_P3_R1131_U73;
  assign new_P3_R1131_U283 = ~new_P3_R1131_U282 | ~new_P3_R1131_U170;
  assign new_P3_R1131_U284 = ~new_P3_U3075 | ~new_P3_R1131_U72;
  assign new_P3_R1131_U285 = ~new_P3_R1131_U169;
  assign new_P3_R1131_U286 = ~new_P3_U3904 | ~new_P3_R1131_U77;
  assign new_P3_R1131_U287 = ~new_P3_U3065 | ~new_P3_R1131_U74;
  assign new_P3_R1131_U288 = ~new_P3_U3060 | ~new_P3_R1131_U75;
  assign new_P3_R1131_U289 = ~new_P3_R1131_U197 | ~new_P3_R1131_U11;
  assign new_P3_R1131_U290 = ~new_P3_R1131_U12 | ~new_P3_R1131_U289;
  assign new_P3_R1131_U291 = ~new_P3_U3906 | ~new_P3_R1131_U79;
  assign new_P3_R1131_U292 = ~new_P3_U3904 | ~new_P3_R1131_U77;
  assign new_P3_R1131_U293 = ~new_P3_R1131_U129 | ~new_P3_R1131_U169;
  assign new_P3_R1131_U294 = ~new_P3_R1131_U292 | ~new_P3_R1131_U290;
  assign new_P3_R1131_U295 = ~new_P3_R1131_U166;
  assign new_P3_R1131_U296 = ~new_P3_U3903 | ~new_P3_R1131_U82;
  assign new_P3_R1131_U297 = ~new_P3_R1131_U296 | ~new_P3_R1131_U166;
  assign new_P3_R1131_U298 = ~new_P3_U3064 | ~new_P3_R1131_U81;
  assign new_P3_R1131_U299 = ~new_P3_R1131_U165;
  assign new_P3_R1131_U300 = ~new_P3_U3902 | ~new_P3_R1131_U84;
  assign new_P3_R1131_U301 = ~new_P3_R1131_U300 | ~new_P3_R1131_U165;
  assign new_P3_R1131_U302 = ~new_P3_U3057 | ~new_P3_R1131_U83;
  assign new_P3_R1131_U303 = ~new_P3_R1131_U91;
  assign new_P3_R1131_U304 = ~new_P3_R1131_U130 | ~new_P3_R1131_U91;
  assign new_P3_R1131_U305 = ~new_P3_R1131_U88 | ~new_P3_R1131_U87;
  assign new_P3_R1131_U306 = ~new_P3_R1131_U305 | ~new_P3_R1131_U85;
  assign new_P3_R1131_U307 = ~new_P3_U3052 | ~new_P3_R1131_U186;
  assign new_P3_R1131_U308 = ~new_P3_R1131_U163;
  assign new_P3_R1131_U309 = ~new_P3_U3899 | ~new_P3_R1131_U90;
  assign new_P3_R1131_U310 = ~new_P3_U3053 | ~new_P3_R1131_U89;
  assign new_P3_R1131_U311 = ~new_P3_R1131_U303 | ~new_P3_R1131_U87;
  assign new_P3_R1131_U312 = ~new_P3_R1131_U137 | ~new_P3_R1131_U311;
  assign new_P3_R1131_U313 = ~new_P3_R1131_U91 | ~new_P3_R1131_U192;
  assign new_P3_R1131_U314 = ~new_P3_R1131_U136 | ~new_P3_R1131_U313;
  assign new_P3_R1131_U315 = ~new_P3_R1131_U192 | ~new_P3_R1131_U87;
  assign new_P3_R1131_U316 = ~new_P3_R1131_U291 | ~new_P3_R1131_U169;
  assign new_P3_R1131_U317 = ~new_P3_R1131_U92;
  assign new_P3_R1131_U318 = ~new_P3_U3060 | ~new_P3_R1131_U75;
  assign new_P3_R1131_U319 = ~new_P3_R1131_U317 | ~new_P3_R1131_U318;
  assign new_P3_R1131_U320 = ~new_P3_R1131_U141 | ~new_P3_R1131_U319;
  assign new_P3_R1131_U321 = ~new_P3_R1131_U92 | ~new_P3_R1131_U191;
  assign new_P3_R1131_U322 = ~new_P3_U3904 | ~new_P3_R1131_U77;
  assign new_P3_R1131_U323 = ~new_P3_R1131_U140 | ~new_P3_R1131_U321;
  assign new_P3_R1131_U324 = ~new_P3_U3060 | ~new_P3_R1131_U75;
  assign new_P3_R1131_U325 = ~new_P3_R1131_U191 | ~new_P3_R1131_U324;
  assign new_P3_R1131_U326 = ~new_P3_R1131_U291 | ~new_P3_R1131_U80;
  assign new_P3_R1131_U327 = ~new_P3_R1131_U267 | ~new_P3_R1131_U179;
  assign new_P3_R1131_U328 = ~new_P3_R1131_U93;
  assign new_P3_R1131_U329 = ~new_P3_U3073 | ~new_P3_R1131_U61;
  assign new_P3_R1131_U330 = ~new_P3_R1131_U328 | ~new_P3_R1131_U329;
  assign new_P3_R1131_U331 = ~new_P3_R1131_U148 | ~new_P3_R1131_U330;
  assign new_P3_R1131_U332 = ~new_P3_R1131_U93 | ~new_P3_R1131_U190;
  assign new_P3_R1131_U333 = ~new_P3_U3437 | ~new_P3_R1131_U63;
  assign new_P3_R1131_U334 = ~new_P3_R1131_U147 | ~new_P3_R1131_U332;
  assign new_P3_R1131_U335 = ~new_P3_U3073 | ~new_P3_R1131_U61;
  assign new_P3_R1131_U336 = ~new_P3_R1131_U190 | ~new_P3_R1131_U335;
  assign new_P3_R1131_U337 = ~new_P3_R1131_U267 | ~new_P3_R1131_U66;
  assign new_P3_R1131_U338 = ~new_P3_R1131_U222 | ~new_P3_R1131_U154;
  assign new_P3_R1131_U339 = ~new_P3_R1131_U94;
  assign new_P3_R1131_U340 = ~new_P3_U3061 | ~new_P3_R1131_U52;
  assign new_P3_R1131_U341 = ~new_P3_R1131_U339 | ~new_P3_R1131_U340;
  assign new_P3_R1131_U342 = ~new_P3_R1131_U152 | ~new_P3_R1131_U341;
  assign new_P3_R1131_U343 = ~new_P3_R1131_U94 | ~new_P3_R1131_U189;
  assign new_P3_R1131_U344 = ~new_P3_U3422 | ~new_P3_R1131_U53;
  assign new_P3_R1131_U345 = ~new_P3_R1131_U151 | ~new_P3_R1131_U343;
  assign new_P3_R1131_U346 = ~new_P3_U3061 | ~new_P3_R1131_U52;
  assign new_P3_R1131_U347 = ~new_P3_R1131_U189 | ~new_P3_R1131_U346;
  assign new_P3_R1131_U348 = ~new_P3_U3076 | ~new_P3_R1131_U30;
  assign new_P3_R1131_U349 = ~new_P3_U3077 | ~new_P3_R1131_U171;
  assign new_P3_R1131_U350 = ~new_P3_U3081 | ~new_P3_R1131_U174;
  assign new_P3_R1131_U351 = ~new_P3_R1131_U134 | ~new_P3_R1131_U133 | ~new_P3_R1131_U304;
  assign new_P3_R1131_U352 = ~new_P3_U3398 | ~new_P3_R1131_U35;
  assign new_P3_R1131_U353 = ~new_P3_U3413 | ~new_P3_R1131_U220;
  assign new_P3_R1131_U354 = ~new_P3_R1131_U353 | ~new_P3_R1131_U219;
  assign new_P3_R1131_U355 = ~new_P3_U3900 | ~new_P3_R1131_U88;
  assign new_P3_R1131_U356 = ~new_P3_R1131_U119 | ~new_P3_R1131_U158;
  assign new_P3_R1131_U357 = ~new_P3_R1131_U216 | ~new_P3_R1131_U14;
  assign new_P3_R1131_U358 = ~new_P3_U3416 | ~new_P3_R1131_U46;
  assign new_P3_R1131_U359 = ~new_P3_U3082 | ~new_P3_R1131_U45;
  assign new_P3_R1131_U360 = ~new_P3_R1131_U223 | ~new_P3_R1131_U154;
  assign new_P3_R1131_U361 = ~new_P3_R1131_U221 | ~new_P3_R1131_U153;
  assign new_P3_R1131_U362 = ~new_P3_U3413 | ~new_P3_R1131_U27;
  assign new_P3_R1131_U363 = ~new_P3_U3083 | ~new_P3_R1131_U28;
  assign new_P3_R1131_U364 = ~new_P3_U3413 | ~new_P3_R1131_U27;
  assign new_P3_R1131_U365 = ~new_P3_U3083 | ~new_P3_R1131_U28;
  assign new_P3_R1131_U366 = ~new_P3_R1131_U365 | ~new_P3_R1131_U364;
  assign new_P3_R1131_U367 = ~new_P3_U3410 | ~new_P3_R1131_U25;
  assign new_P3_R1131_U368 = ~new_P3_U3069 | ~new_P3_R1131_U39;
  assign new_P3_R1131_U369 = ~new_P3_R1131_U228 | ~new_P3_R1131_U47;
  assign new_P3_R1131_U370 = ~new_P3_R1131_U155 | ~new_P3_R1131_U217;
  assign new_P3_R1131_U371 = ~new_P3_U3407 | ~new_P3_R1131_U40;
  assign new_P3_R1131_U372 = ~new_P3_U3070 | ~new_P3_R1131_U37;
  assign new_P3_R1131_U373 = ~new_P3_R1131_U372 | ~new_P3_R1131_U371;
  assign new_P3_R1131_U374 = ~new_P3_U3404 | ~new_P3_R1131_U41;
  assign new_P3_R1131_U375 = ~new_P3_U3066 | ~new_P3_R1131_U36;
  assign new_P3_R1131_U376 = ~new_P3_R1131_U238 | ~new_P3_R1131_U48;
  assign new_P3_R1131_U377 = ~new_P3_R1131_U156 | ~new_P3_R1131_U230;
  assign new_P3_R1131_U378 = ~new_P3_U3401 | ~new_P3_R1131_U42;
  assign new_P3_R1131_U379 = ~new_P3_U3059 | ~new_P3_R1131_U38;
  assign new_P3_R1131_U380 = ~new_P3_R1131_U239 | ~new_P3_R1131_U158;
  assign new_P3_R1131_U381 = ~new_P3_R1131_U207 | ~new_P3_R1131_U157;
  assign new_P3_R1131_U382 = ~new_P3_U3398 | ~new_P3_R1131_U35;
  assign new_P3_R1131_U383 = ~new_P3_U3063 | ~new_P3_R1131_U32;
  assign new_P3_R1131_U384 = ~new_P3_U3398 | ~new_P3_R1131_U35;
  assign new_P3_R1131_U385 = ~new_P3_U3063 | ~new_P3_R1131_U32;
  assign new_P3_R1131_U386 = ~new_P3_R1131_U385 | ~new_P3_R1131_U384;
  assign new_P3_R1131_U387 = ~new_P3_U3395 | ~new_P3_R1131_U33;
  assign new_P3_R1131_U388 = ~new_P3_U3067 | ~new_P3_R1131_U29;
  assign new_P3_R1131_U389 = ~new_P3_R1131_U244 | ~new_P3_R1131_U49;
  assign new_P3_R1131_U390 = ~new_P3_R1131_U159 | ~new_P3_R1131_U202;
  assign new_P3_R1131_U391 = ~new_P3_U3908 | ~new_P3_R1131_U161;
  assign new_P3_R1131_U392 = ~new_P3_U3054 | ~new_P3_R1131_U160;
  assign new_P3_R1131_U393 = ~new_P3_U3908 | ~new_P3_R1131_U161;
  assign new_P3_R1131_U394 = ~new_P3_U3054 | ~new_P3_R1131_U160;
  assign new_P3_R1131_U395 = ~new_P3_R1131_U394 | ~new_P3_R1131_U393;
  assign new_P3_R1131_U396 = ~new_P3_R1131_U89 | ~new_P3_U3053 | ~new_P3_R1131_U395;
  assign new_P3_R1131_U397 = ~new_P3_U3899 | ~new_P3_R1131_U15 | ~new_P3_R1131_U90;
  assign new_P3_R1131_U398 = ~new_P3_U3899 | ~new_P3_R1131_U90;
  assign new_P3_R1131_U399 = ~new_P3_U3053 | ~new_P3_R1131_U89;
  assign new_P3_R1131_U400 = ~new_P3_R1131_U135;
  assign new_P3_R1131_U401 = ~new_P3_R1131_U308 | ~new_P3_R1131_U400;
  assign new_P3_R1131_U402 = ~new_P3_R1131_U135 | ~new_P3_R1131_U163;
  assign new_P3_R1131_U403 = ~new_P3_U3900 | ~new_P3_R1131_U88;
  assign new_P3_R1131_U404 = ~new_P3_U3052 | ~new_P3_R1131_U85;
  assign new_P3_R1131_U405 = ~new_P3_U3900 | ~new_P3_R1131_U88;
  assign new_P3_R1131_U406 = ~new_P3_U3052 | ~new_P3_R1131_U85;
  assign new_P3_R1131_U407 = ~new_P3_R1131_U406 | ~new_P3_R1131_U405;
  assign new_P3_R1131_U408 = ~new_P3_U3901 | ~new_P3_R1131_U86;
  assign new_P3_R1131_U409 = ~new_P3_U3056 | ~new_P3_R1131_U50;
  assign new_P3_R1131_U410 = ~new_P3_R1131_U315 | ~new_P3_R1131_U91;
  assign new_P3_R1131_U411 = ~new_P3_R1131_U164 | ~new_P3_R1131_U303;
  assign new_P3_R1131_U412 = ~new_P3_U3902 | ~new_P3_R1131_U84;
  assign new_P3_R1131_U413 = ~new_P3_U3057 | ~new_P3_R1131_U83;
  assign new_P3_R1131_U414 = ~new_P3_R1131_U138;
  assign new_P3_R1131_U415 = ~new_P3_R1131_U299 | ~new_P3_R1131_U414;
  assign new_P3_R1131_U416 = ~new_P3_R1131_U138 | ~new_P3_R1131_U165;
  assign new_P3_R1131_U417 = ~new_P3_U3903 | ~new_P3_R1131_U82;
  assign new_P3_R1131_U418 = ~new_P3_U3064 | ~new_P3_R1131_U81;
  assign new_P3_R1131_U419 = ~new_P3_R1131_U139;
  assign new_P3_R1131_U420 = ~new_P3_R1131_U295 | ~new_P3_R1131_U419;
  assign new_P3_R1131_U421 = ~new_P3_R1131_U139 | ~new_P3_R1131_U166;
  assign new_P3_R1131_U422 = ~new_P3_U3904 | ~new_P3_R1131_U77;
  assign new_P3_R1131_U423 = ~new_P3_U3065 | ~new_P3_R1131_U74;
  assign new_P3_R1131_U424 = ~new_P3_R1131_U423 | ~new_P3_R1131_U422;
  assign new_P3_R1131_U425 = ~new_P3_U3905 | ~new_P3_R1131_U78;
  assign new_P3_R1131_U426 = ~new_P3_U3060 | ~new_P3_R1131_U75;
  assign new_P3_R1131_U427 = ~new_P3_R1131_U325 | ~new_P3_R1131_U92;
  assign new_P3_R1131_U428 = ~new_P3_R1131_U167 | ~new_P3_R1131_U317;
  assign new_P3_R1131_U429 = ~new_P3_U3906 | ~new_P3_R1131_U79;
  assign new_P3_R1131_U430 = ~new_P3_U3074 | ~new_P3_R1131_U76;
  assign new_P3_R1131_U431 = ~new_P3_R1131_U326 | ~new_P3_R1131_U169;
  assign new_P3_R1131_U432 = ~new_P3_R1131_U285 | ~new_P3_R1131_U168;
  assign new_P3_R1131_U433 = ~new_P3_U3907 | ~new_P3_R1131_U73;
  assign new_P3_R1131_U434 = ~new_P3_U3075 | ~new_P3_R1131_U72;
  assign new_P3_R1131_U435 = ~new_P3_R1131_U142;
  assign new_P3_R1131_U436 = ~new_P3_R1131_U281 | ~new_P3_R1131_U435;
  assign new_P3_R1131_U437 = ~new_P3_R1131_U142 | ~new_P3_R1131_U170;
  assign new_P3_R1131_U438 = ~new_P3_U3392 | ~new_P3_R1131_U31;
  assign new_P3_R1131_U439 = ~new_P3_U3077 | ~new_P3_R1131_U171;
  assign new_P3_R1131_U440 = ~new_P3_R1131_U143;
  assign new_P3_R1131_U441 = ~new_P3_R1131_U200 | ~new_P3_R1131_U440;
  assign new_P3_R1131_U442 = ~new_P3_R1131_U143 | ~new_P3_R1131_U172;
  assign new_P3_R1131_U443 = ~new_P3_U3445 | ~new_P3_R1131_U71;
  assign new_P3_R1131_U444 = ~new_P3_U3080 | ~new_P3_R1131_U70;
  assign new_P3_R1131_U445 = ~new_P3_R1131_U144;
  assign new_P3_R1131_U446 = ~new_P3_R1131_U277 | ~new_P3_R1131_U445;
  assign new_P3_R1131_U447 = ~new_P3_R1131_U144 | ~new_P3_R1131_U173;
  assign new_P3_R1131_U448 = ~new_P3_U3443 | ~new_P3_R1131_U69;
  assign new_P3_R1131_U449 = ~new_P3_U3081 | ~new_P3_R1131_U174;
  assign new_P3_R1131_U450 = ~new_P3_R1131_U145;
  assign new_P3_R1131_U451 = ~new_P3_R1131_U275 | ~new_P3_R1131_U450;
  assign new_P3_R1131_U452 = ~new_P3_R1131_U145 | ~new_P3_R1131_U175;
  assign new_P3_R1131_U453 = ~new_P3_U3440 | ~new_P3_R1131_U68;
  assign new_P3_R1131_U454 = ~new_P3_U3068 | ~new_P3_R1131_U67;
  assign new_P3_R1131_U455 = ~new_P3_R1131_U146;
  assign new_P3_R1131_U456 = ~new_P3_R1131_U271 | ~new_P3_R1131_U455;
  assign new_P3_R1131_U457 = ~new_P3_R1131_U146 | ~new_P3_R1131_U176;
  assign new_P3_R1131_U458 = ~new_P3_U3437 | ~new_P3_R1131_U63;
  assign new_P3_R1131_U459 = ~new_P3_U3072 | ~new_P3_R1131_U60;
  assign new_P3_R1131_U460 = ~new_P3_R1131_U459 | ~new_P3_R1131_U458;
  assign new_P3_R1131_U461 = ~new_P3_U3434 | ~new_P3_R1131_U64;
  assign new_P3_R1131_U462 = ~new_P3_U3073 | ~new_P3_R1131_U61;
  assign new_P3_R1131_U463 = ~new_P3_R1131_U336 | ~new_P3_R1131_U93;
  assign new_P3_R1131_U464 = ~new_P3_R1131_U177 | ~new_P3_R1131_U328;
  assign new_P3_R1131_U465 = ~new_P3_U3431 | ~new_P3_R1131_U65;
  assign new_P3_R1131_U466 = ~new_P3_U3078 | ~new_P3_R1131_U62;
  assign new_P3_R1131_U467 = ~new_P3_R1131_U337 | ~new_P3_R1131_U179;
  assign new_P3_R1131_U468 = ~new_P3_R1131_U261 | ~new_P3_R1131_U178;
  assign new_P3_R1131_U469 = ~new_P3_U3428 | ~new_P3_R1131_U59;
  assign new_P3_R1131_U470 = ~new_P3_U3079 | ~new_P3_R1131_U58;
  assign new_P3_R1131_U471 = ~new_P3_R1131_U149;
  assign new_P3_R1131_U472 = ~new_P3_R1131_U257 | ~new_P3_R1131_U471;
  assign new_P3_R1131_U473 = ~new_P3_R1131_U149 | ~new_P3_R1131_U180;
  assign new_P3_R1131_U474 = ~new_P3_U3425 | ~new_P3_R1131_U57;
  assign new_P3_R1131_U475 = ~new_P3_U3071 | ~new_P3_R1131_U56;
  assign new_P3_R1131_U476 = ~new_P3_R1131_U150;
  assign new_P3_R1131_U477 = ~new_P3_R1131_U253 | ~new_P3_R1131_U476;
  assign new_P3_R1131_U478 = ~new_P3_R1131_U150 | ~new_P3_R1131_U181;
  assign new_P3_R1131_U479 = ~new_P3_U3422 | ~new_P3_R1131_U53;
  assign new_P3_R1131_U480 = ~new_P3_U3062 | ~new_P3_R1131_U51;
  assign new_P3_R1131_U481 = ~new_P3_R1131_U480 | ~new_P3_R1131_U479;
  assign new_P3_R1131_U482 = ~new_P3_U3419 | ~new_P3_R1131_U54;
  assign new_P3_R1131_U483 = ~new_P3_U3061 | ~new_P3_R1131_U52;
  assign new_P3_R1131_U484 = ~new_P3_R1131_U347 | ~new_P3_R1131_U94;
  assign new_P3_R1131_U485 = ~new_P3_R1131_U182 | ~new_P3_R1131_U339;
  assign new_P3_R1054_U6 = new_P3_R1054_U102 & new_P3_R1054_U118;
  assign new_P3_R1054_U7 = new_P3_R1054_U120 & new_P3_R1054_U119;
  assign new_P3_R1054_U8 = new_P3_R1054_U99 & new_P3_R1054_U157;
  assign new_P3_R1054_U9 = new_P3_R1054_U159 & new_P3_R1054_U158;
  assign new_P3_R1054_U10 = new_P3_R1054_U100 & new_P3_R1054_U174;
  assign new_P3_R1054_U11 = new_P3_R1054_U176 & new_P3_R1054_U175;
  assign new_P3_R1054_U12 = ~new_P3_R1054_U207 | ~new_P3_R1054_U210;
  assign new_P3_R1054_U13 = ~new_P3_R1054_U196 | ~new_P3_R1054_U199;
  assign new_P3_R1054_U14 = ~new_P3_R1054_U153 | ~new_P3_R1054_U155;
  assign new_P3_R1054_U15 = ~new_P3_R1054_U145 | ~new_P3_R1054_U148;
  assign new_P3_R1054_U16 = ~new_P3_R1054_U137 | ~new_P3_R1054_U139;
  assign new_P3_R1054_U17 = ~new_P3_R1054_U21 | ~new_P3_R1054_U213;
  assign new_P3_R1054_U18 = ~new_P3_U3409;
  assign new_P3_R1054_U19 = ~new_P3_U3394;
  assign new_P3_R1054_U20 = ~new_P3_U3386;
  assign new_P3_R1054_U21 = ~new_P3_U3386 | ~new_P3_R1054_U65;
  assign new_P3_R1054_U22 = ~new_P3_U3573;
  assign new_P3_R1054_U23 = ~new_P3_U3397;
  assign new_P3_R1054_U24 = ~new_P3_U3562;
  assign new_P3_R1054_U25 = ~new_P3_U3562 | ~new_P3_R1054_U19;
  assign new_P3_R1054_U26 = ~new_P3_U3561;
  assign new_P3_R1054_U27 = ~new_P3_U3406;
  assign new_P3_R1054_U28 = ~new_P3_U3403;
  assign new_P3_R1054_U29 = ~new_P3_U3400;
  assign new_P3_R1054_U30 = ~new_P3_U3558;
  assign new_P3_R1054_U31 = ~new_P3_U3559;
  assign new_P3_R1054_U32 = ~new_P3_U3560;
  assign new_P3_R1054_U33 = ~new_P3_U3560 | ~new_P3_R1054_U29;
  assign new_P3_R1054_U34 = ~new_P3_U3412;
  assign new_P3_R1054_U35 = ~new_P3_U3557;
  assign new_P3_R1054_U36 = ~new_P3_U3557 | ~new_P3_R1054_U18;
  assign new_P3_R1054_U37 = ~new_P3_U3556;
  assign new_P3_R1054_U38 = ~new_P3_U3415;
  assign new_P3_R1054_U39 = ~new_P3_U3555;
  assign new_P3_R1054_U40 = ~new_P3_R1054_U126 | ~new_P3_R1054_U125;
  assign new_P3_R1054_U41 = ~new_P3_R1054_U33 | ~new_P3_R1054_U141;
  assign new_P3_R1054_U42 = ~new_P3_R1054_U110 | ~new_P3_R1054_U109;
  assign new_P3_R1054_U43 = ~new_P3_U3421;
  assign new_P3_R1054_U44 = ~new_P3_U3418;
  assign new_P3_R1054_U45 = ~new_P3_U3571;
  assign new_P3_R1054_U46 = ~new_P3_U3572;
  assign new_P3_R1054_U47 = ~new_P3_U3555 | ~new_P3_R1054_U38;
  assign new_P3_R1054_U48 = ~new_P3_U3424;
  assign new_P3_R1054_U49 = ~new_P3_U3570;
  assign new_P3_R1054_U50 = ~new_P3_U3427;
  assign new_P3_R1054_U51 = ~new_P3_U3569;
  assign new_P3_R1054_U52 = ~new_P3_U3436;
  assign new_P3_R1054_U53 = ~new_P3_U3433;
  assign new_P3_R1054_U54 = ~new_P3_U3430;
  assign new_P3_R1054_U55 = ~new_P3_U3566;
  assign new_P3_R1054_U56 = ~new_P3_U3567;
  assign new_P3_R1054_U57 = ~new_P3_U3568;
  assign new_P3_R1054_U58 = ~new_P3_U3568 | ~new_P3_R1054_U54;
  assign new_P3_R1054_U59 = ~new_P3_U3439;
  assign new_P3_R1054_U60 = ~new_P3_U3565;
  assign new_P3_R1054_U61 = ~new_P3_R1054_U186 | ~new_P3_R1054_U185;
  assign new_P3_R1054_U62 = ~new_P3_U3564;
  assign new_P3_R1054_U63 = ~new_P3_R1054_U58 | ~new_P3_R1054_U192;
  assign new_P3_R1054_U64 = ~new_P3_R1054_U47 | ~new_P3_R1054_U203;
  assign new_P3_R1054_U65 = ~new_P3_U3574;
  assign new_P3_R1054_U66 = ~new_P3_R1054_U251 | ~new_P3_R1054_U250;
  assign new_P3_R1054_U67 = ~new_P3_R1054_U256 | ~new_P3_R1054_U255;
  assign new_P3_R1054_U68 = ~new_P3_R1054_U261 | ~new_P3_R1054_U260;
  assign new_P3_R1054_U69 = ~new_P3_R1054_U266 | ~new_P3_R1054_U265;
  assign new_P3_R1054_U70 = ~new_P3_R1054_U282 | ~new_P3_R1054_U281;
  assign new_P3_R1054_U71 = ~new_P3_R1054_U287 | ~new_P3_R1054_U286;
  assign new_P3_R1054_U72 = ~new_P3_R1054_U217 | ~new_P3_R1054_U216;
  assign new_P3_R1054_U73 = ~new_P3_R1054_U226 | ~new_P3_R1054_U225;
  assign new_P3_R1054_U74 = ~new_P3_R1054_U233 | ~new_P3_R1054_U232;
  assign new_P3_R1054_U75 = ~new_P3_R1054_U237 | ~new_P3_R1054_U236;
  assign new_P3_R1054_U76 = ~new_P3_R1054_U246 | ~new_P3_R1054_U245;
  assign new_P3_R1054_U77 = ~new_P3_R1054_U273 | ~new_P3_R1054_U272;
  assign new_P3_R1054_U78 = ~new_P3_R1054_U277 | ~new_P3_R1054_U276;
  assign new_P3_R1054_U79 = ~new_P3_R1054_U294 | ~new_P3_R1054_U293;
  assign new_P3_R1054_U80 = ~new_P3_R1054_U248 | ~new_P3_R1054_U247;
  assign new_P3_R1054_U81 = ~new_P3_R1054_U253 | ~new_P3_R1054_U252;
  assign new_P3_R1054_U82 = ~new_P3_R1054_U258 | ~new_P3_R1054_U257;
  assign new_P3_R1054_U83 = ~new_P3_R1054_U263 | ~new_P3_R1054_U262;
  assign new_P3_R1054_U84 = ~new_P3_R1054_U279 | ~new_P3_R1054_U278;
  assign new_P3_R1054_U85 = ~new_P3_R1054_U284 | ~new_P3_R1054_U283;
  assign new_P3_R1054_U86 = ~new_P3_R1054_U129 | ~new_P3_R1054_U131 | ~new_P3_R1054_U132;
  assign new_P3_R1054_U87 = ~new_P3_R1054_U113 | ~new_P3_R1054_U115 | ~new_P3_R1054_U116;
  assign new_P3_R1054_U88 = ~new_P3_U3391;
  assign new_P3_R1054_U89 = ~new_P3_U3379;
  assign new_P3_R1054_U90 = ~new_P3_U3563;
  assign new_P3_R1054_U91 = ~new_P3_R1054_U190 | ~new_P3_R1054_U189;
  assign new_P3_R1054_U92 = ~new_P3_U3442;
  assign new_P3_R1054_U93 = ~new_P3_R1054_U182 | ~new_P3_R1054_U181;
  assign new_P3_R1054_U94 = ~new_P3_R1054_U172 | ~new_P3_R1054_U171;
  assign new_P3_R1054_U95 = ~new_P3_R1054_U168 | ~new_P3_R1054_U167;
  assign new_P3_R1054_U96 = ~new_P3_R1054_U164 | ~new_P3_R1054_U163;
  assign new_P3_R1054_U97 = ~new_P3_R1054_U25;
  assign new_P3_R1054_U98 = ~new_P3_R1054_U36;
  assign new_P3_R1054_U99 = ~new_P3_U3418 | ~new_P3_R1054_U46;
  assign new_P3_R1054_U100 = ~new_P3_U3433 | ~new_P3_R1054_U56;
  assign new_P3_R1054_U101 = ~new_P3_U3394 | ~new_P3_R1054_U24;
  assign new_P3_R1054_U102 = ~new_P3_U3403 | ~new_P3_R1054_U31;
  assign new_P3_R1054_U103 = ~new_P3_U3409 | ~new_P3_R1054_U35;
  assign new_P3_R1054_U104 = ~new_P3_R1054_U58;
  assign new_P3_R1054_U105 = ~new_P3_R1054_U33;
  assign new_P3_R1054_U106 = ~new_P3_R1054_U47;
  assign new_P3_R1054_U107 = ~new_P3_R1054_U21;
  assign new_P3_R1054_U108 = ~new_P3_R1054_U107 | ~new_P3_R1054_U22;
  assign new_P3_R1054_U109 = ~new_P3_R1054_U108 | ~new_P3_R1054_U88;
  assign new_P3_R1054_U110 = ~new_P3_U3573 | ~new_P3_R1054_U21;
  assign new_P3_R1054_U111 = ~new_P3_R1054_U42;
  assign new_P3_R1054_U112 = ~new_P3_U3397 | ~new_P3_R1054_U26;
  assign new_P3_R1054_U113 = ~new_P3_R1054_U42 | ~new_P3_R1054_U112 | ~new_P3_R1054_U101;
  assign new_P3_R1054_U114 = ~new_P3_R1054_U26 | ~new_P3_R1054_U25;
  assign new_P3_R1054_U115 = ~new_P3_R1054_U114 | ~new_P3_R1054_U23;
  assign new_P3_R1054_U116 = ~new_P3_U3561 | ~new_P3_R1054_U97;
  assign new_P3_R1054_U117 = ~new_P3_R1054_U87;
  assign new_P3_R1054_U118 = ~new_P3_U3406 | ~new_P3_R1054_U30;
  assign new_P3_R1054_U119 = ~new_P3_U3558 | ~new_P3_R1054_U27;
  assign new_P3_R1054_U120 = ~new_P3_U3559 | ~new_P3_R1054_U28;
  assign new_P3_R1054_U121 = ~new_P3_R1054_U105 | ~new_P3_R1054_U6;
  assign new_P3_R1054_U122 = ~new_P3_R1054_U7 | ~new_P3_R1054_U121;
  assign new_P3_R1054_U123 = ~new_P3_U3400 | ~new_P3_R1054_U32;
  assign new_P3_R1054_U124 = ~new_P3_U3406 | ~new_P3_R1054_U30;
  assign new_P3_R1054_U125 = ~new_P3_R1054_U87 | ~new_P3_R1054_U123 | ~new_P3_R1054_U6;
  assign new_P3_R1054_U126 = ~new_P3_R1054_U124 | ~new_P3_R1054_U122;
  assign new_P3_R1054_U127 = ~new_P3_R1054_U40;
  assign new_P3_R1054_U128 = ~new_P3_U3412 | ~new_P3_R1054_U37;
  assign new_P3_R1054_U129 = ~new_P3_R1054_U40 | ~new_P3_R1054_U128 | ~new_P3_R1054_U103;
  assign new_P3_R1054_U130 = ~new_P3_R1054_U37 | ~new_P3_R1054_U36;
  assign new_P3_R1054_U131 = ~new_P3_R1054_U130 | ~new_P3_R1054_U34;
  assign new_P3_R1054_U132 = ~new_P3_U3556 | ~new_P3_R1054_U98;
  assign new_P3_R1054_U133 = ~new_P3_R1054_U86;
  assign new_P3_R1054_U134 = ~new_P3_U3415 | ~new_P3_R1054_U39;
  assign new_P3_R1054_U135 = ~new_P3_R1054_U134 | ~new_P3_R1054_U47;
  assign new_P3_R1054_U136 = ~new_P3_R1054_U127 | ~new_P3_R1054_U36;
  assign new_P3_R1054_U137 = ~new_P3_R1054_U136 | ~new_P3_R1054_U222 | ~new_P3_R1054_U103;
  assign new_P3_R1054_U138 = ~new_P3_R1054_U40 | ~new_P3_R1054_U103;
  assign new_P3_R1054_U139 = ~new_P3_R1054_U138 | ~new_P3_R1054_U36 | ~new_P3_R1054_U219 | ~new_P3_R1054_U218;
  assign new_P3_R1054_U140 = ~new_P3_R1054_U36 | ~new_P3_R1054_U103;
  assign new_P3_R1054_U141 = ~new_P3_R1054_U123 | ~new_P3_R1054_U87;
  assign new_P3_R1054_U142 = ~new_P3_R1054_U41;
  assign new_P3_R1054_U143 = ~new_P3_U3559 | ~new_P3_R1054_U28;
  assign new_P3_R1054_U144 = ~new_P3_R1054_U142 | ~new_P3_R1054_U143;
  assign new_P3_R1054_U145 = ~new_P3_R1054_U144 | ~new_P3_R1054_U229 | ~new_P3_R1054_U102;
  assign new_P3_R1054_U146 = ~new_P3_R1054_U41 | ~new_P3_R1054_U102;
  assign new_P3_R1054_U147 = ~new_P3_U3406 | ~new_P3_R1054_U30;
  assign new_P3_R1054_U148 = ~new_P3_R1054_U146 | ~new_P3_R1054_U147 | ~new_P3_R1054_U7;
  assign new_P3_R1054_U149 = ~new_P3_U3559 | ~new_P3_R1054_U28;
  assign new_P3_R1054_U150 = ~new_P3_R1054_U102 | ~new_P3_R1054_U149;
  assign new_P3_R1054_U151 = ~new_P3_R1054_U123 | ~new_P3_R1054_U33;
  assign new_P3_R1054_U152 = ~new_P3_R1054_U111 | ~new_P3_R1054_U25;
  assign new_P3_R1054_U153 = ~new_P3_R1054_U152 | ~new_P3_R1054_U242 | ~new_P3_R1054_U101;
  assign new_P3_R1054_U154 = ~new_P3_R1054_U42 | ~new_P3_R1054_U101;
  assign new_P3_R1054_U155 = ~new_P3_R1054_U154 | ~new_P3_R1054_U25 | ~new_P3_R1054_U239 | ~new_P3_R1054_U238;
  assign new_P3_R1054_U156 = ~new_P3_R1054_U25 | ~new_P3_R1054_U101;
  assign new_P3_R1054_U157 = ~new_P3_U3421 | ~new_P3_R1054_U45;
  assign new_P3_R1054_U158 = ~new_P3_U3571 | ~new_P3_R1054_U43;
  assign new_P3_R1054_U159 = ~new_P3_U3572 | ~new_P3_R1054_U44;
  assign new_P3_R1054_U160 = ~new_P3_R1054_U106 | ~new_P3_R1054_U8;
  assign new_P3_R1054_U161 = ~new_P3_R1054_U9 | ~new_P3_R1054_U160;
  assign new_P3_R1054_U162 = ~new_P3_U3421 | ~new_P3_R1054_U45;
  assign new_P3_R1054_U163 = ~new_P3_R1054_U86 | ~new_P3_R1054_U134 | ~new_P3_R1054_U8;
  assign new_P3_R1054_U164 = ~new_P3_R1054_U162 | ~new_P3_R1054_U161;
  assign new_P3_R1054_U165 = ~new_P3_R1054_U96;
  assign new_P3_R1054_U166 = ~new_P3_U3424 | ~new_P3_R1054_U49;
  assign new_P3_R1054_U167 = ~new_P3_R1054_U166 | ~new_P3_R1054_U96;
  assign new_P3_R1054_U168 = ~new_P3_U3570 | ~new_P3_R1054_U48;
  assign new_P3_R1054_U169 = ~new_P3_R1054_U95;
  assign new_P3_R1054_U170 = ~new_P3_U3427 | ~new_P3_R1054_U51;
  assign new_P3_R1054_U171 = ~new_P3_R1054_U170 | ~new_P3_R1054_U95;
  assign new_P3_R1054_U172 = ~new_P3_U3569 | ~new_P3_R1054_U50;
  assign new_P3_R1054_U173 = ~new_P3_R1054_U94;
  assign new_P3_R1054_U174 = ~new_P3_U3436 | ~new_P3_R1054_U55;
  assign new_P3_R1054_U175 = ~new_P3_U3566 | ~new_P3_R1054_U52;
  assign new_P3_R1054_U176 = ~new_P3_U3567 | ~new_P3_R1054_U53;
  assign new_P3_R1054_U177 = ~new_P3_R1054_U104 | ~new_P3_R1054_U10;
  assign new_P3_R1054_U178 = ~new_P3_R1054_U11 | ~new_P3_R1054_U177;
  assign new_P3_R1054_U179 = ~new_P3_U3430 | ~new_P3_R1054_U57;
  assign new_P3_R1054_U180 = ~new_P3_U3436 | ~new_P3_R1054_U55;
  assign new_P3_R1054_U181 = ~new_P3_R1054_U94 | ~new_P3_R1054_U179 | ~new_P3_R1054_U10;
  assign new_P3_R1054_U182 = ~new_P3_R1054_U180 | ~new_P3_R1054_U178;
  assign new_P3_R1054_U183 = ~new_P3_R1054_U93;
  assign new_P3_R1054_U184 = ~new_P3_U3439 | ~new_P3_R1054_U60;
  assign new_P3_R1054_U185 = ~new_P3_R1054_U184 | ~new_P3_R1054_U93;
  assign new_P3_R1054_U186 = ~new_P3_U3565 | ~new_P3_R1054_U59;
  assign new_P3_R1054_U187 = ~new_P3_R1054_U61;
  assign new_P3_R1054_U188 = ~new_P3_R1054_U187 | ~new_P3_R1054_U62;
  assign new_P3_R1054_U189 = ~new_P3_R1054_U188 | ~new_P3_R1054_U92;
  assign new_P3_R1054_U190 = ~new_P3_U3564 | ~new_P3_R1054_U61;
  assign new_P3_R1054_U191 = ~new_P3_R1054_U91;
  assign new_P3_R1054_U192 = ~new_P3_R1054_U179 | ~new_P3_R1054_U94;
  assign new_P3_R1054_U193 = ~new_P3_R1054_U63;
  assign new_P3_R1054_U194 = ~new_P3_U3567 | ~new_P3_R1054_U53;
  assign new_P3_R1054_U195 = ~new_P3_R1054_U193 | ~new_P3_R1054_U194;
  assign new_P3_R1054_U196 = ~new_P3_R1054_U195 | ~new_P3_R1054_U269 | ~new_P3_R1054_U100;
  assign new_P3_R1054_U197 = ~new_P3_R1054_U63 | ~new_P3_R1054_U100;
  assign new_P3_R1054_U198 = ~new_P3_U3436 | ~new_P3_R1054_U55;
  assign new_P3_R1054_U199 = ~new_P3_R1054_U197 | ~new_P3_R1054_U198 | ~new_P3_R1054_U11;
  assign new_P3_R1054_U200 = ~new_P3_U3567 | ~new_P3_R1054_U53;
  assign new_P3_R1054_U201 = ~new_P3_R1054_U100 | ~new_P3_R1054_U200;
  assign new_P3_R1054_U202 = ~new_P3_R1054_U179 | ~new_P3_R1054_U58;
  assign new_P3_R1054_U203 = ~new_P3_R1054_U134 | ~new_P3_R1054_U86;
  assign new_P3_R1054_U204 = ~new_P3_R1054_U64;
  assign new_P3_R1054_U205 = ~new_P3_U3572 | ~new_P3_R1054_U44;
  assign new_P3_R1054_U206 = ~new_P3_R1054_U204 | ~new_P3_R1054_U205;
  assign new_P3_R1054_U207 = ~new_P3_R1054_U206 | ~new_P3_R1054_U290 | ~new_P3_R1054_U99;
  assign new_P3_R1054_U208 = ~new_P3_R1054_U64 | ~new_P3_R1054_U99;
  assign new_P3_R1054_U209 = ~new_P3_U3421 | ~new_P3_R1054_U45;
  assign new_P3_R1054_U210 = ~new_P3_R1054_U208 | ~new_P3_R1054_U209 | ~new_P3_R1054_U9;
  assign new_P3_R1054_U211 = ~new_P3_U3572 | ~new_P3_R1054_U44;
  assign new_P3_R1054_U212 = ~new_P3_R1054_U99 | ~new_P3_R1054_U211;
  assign new_P3_R1054_U213 = ~new_P3_U3574 | ~new_P3_R1054_U20;
  assign new_P3_R1054_U214 = ~new_P3_U3415 | ~new_P3_R1054_U39;
  assign new_P3_R1054_U215 = ~new_P3_U3555 | ~new_P3_R1054_U38;
  assign new_P3_R1054_U216 = ~new_P3_R1054_U135 | ~new_P3_R1054_U86;
  assign new_P3_R1054_U217 = ~new_P3_R1054_U133 | ~new_P3_R1054_U215 | ~new_P3_R1054_U214;
  assign new_P3_R1054_U218 = ~new_P3_U3412 | ~new_P3_R1054_U37;
  assign new_P3_R1054_U219 = ~new_P3_U3556 | ~new_P3_R1054_U34;
  assign new_P3_R1054_U220 = ~new_P3_U3412 | ~new_P3_R1054_U37;
  assign new_P3_R1054_U221 = ~new_P3_U3556 | ~new_P3_R1054_U34;
  assign new_P3_R1054_U222 = ~new_P3_R1054_U221 | ~new_P3_R1054_U220;
  assign new_P3_R1054_U223 = ~new_P3_U3409 | ~new_P3_R1054_U35;
  assign new_P3_R1054_U224 = ~new_P3_U3557 | ~new_P3_R1054_U18;
  assign new_P3_R1054_U225 = ~new_P3_R1054_U140 | ~new_P3_R1054_U40;
  assign new_P3_R1054_U226 = ~new_P3_R1054_U127 | ~new_P3_R1054_U224 | ~new_P3_R1054_U223;
  assign new_P3_R1054_U227 = ~new_P3_U3406 | ~new_P3_R1054_U30;
  assign new_P3_R1054_U228 = ~new_P3_U3558 | ~new_P3_R1054_U27;
  assign new_P3_R1054_U229 = ~new_P3_R1054_U228 | ~new_P3_R1054_U227;
  assign new_P3_R1054_U230 = ~new_P3_U3403 | ~new_P3_R1054_U31;
  assign new_P3_R1054_U231 = ~new_P3_U3559 | ~new_P3_R1054_U28;
  assign new_P3_R1054_U232 = ~new_P3_R1054_U150 | ~new_P3_R1054_U41;
  assign new_P3_R1054_U233 = ~new_P3_R1054_U142 | ~new_P3_R1054_U231 | ~new_P3_R1054_U230;
  assign new_P3_R1054_U234 = ~new_P3_U3400 | ~new_P3_R1054_U32;
  assign new_P3_R1054_U235 = ~new_P3_U3560 | ~new_P3_R1054_U29;
  assign new_P3_R1054_U236 = ~new_P3_R1054_U151 | ~new_P3_R1054_U87;
  assign new_P3_R1054_U237 = ~new_P3_R1054_U117 | ~new_P3_R1054_U235 | ~new_P3_R1054_U234;
  assign new_P3_R1054_U238 = ~new_P3_U3397 | ~new_P3_R1054_U26;
  assign new_P3_R1054_U239 = ~new_P3_U3561 | ~new_P3_R1054_U23;
  assign new_P3_R1054_U240 = ~new_P3_U3397 | ~new_P3_R1054_U26;
  assign new_P3_R1054_U241 = ~new_P3_U3561 | ~new_P3_R1054_U23;
  assign new_P3_R1054_U242 = ~new_P3_R1054_U241 | ~new_P3_R1054_U240;
  assign new_P3_R1054_U243 = ~new_P3_U3394 | ~new_P3_R1054_U24;
  assign new_P3_R1054_U244 = ~new_P3_U3562 | ~new_P3_R1054_U19;
  assign new_P3_R1054_U245 = ~new_P3_R1054_U156 | ~new_P3_R1054_U42;
  assign new_P3_R1054_U246 = ~new_P3_R1054_U111 | ~new_P3_R1054_U244 | ~new_P3_R1054_U243;
  assign new_P3_R1054_U247 = ~new_P3_U3391 | ~new_P3_R1054_U22;
  assign new_P3_R1054_U248 = ~new_P3_U3573 | ~new_P3_R1054_U88;
  assign new_P3_R1054_U249 = ~new_P3_R1054_U80;
  assign new_P3_R1054_U250 = ~new_P3_R1054_U249 | ~new_P3_R1054_U107;
  assign new_P3_R1054_U251 = ~new_P3_R1054_U80 | ~new_P3_R1054_U21;
  assign new_P3_R1054_U252 = ~new_P3_U3379 | ~new_P3_R1054_U90;
  assign new_P3_R1054_U253 = ~new_P3_U3563 | ~new_P3_R1054_U89;
  assign new_P3_R1054_U254 = ~new_P3_R1054_U81;
  assign new_P3_R1054_U255 = ~new_P3_R1054_U191 | ~new_P3_R1054_U254;
  assign new_P3_R1054_U256 = ~new_P3_R1054_U81 | ~new_P3_R1054_U91;
  assign new_P3_R1054_U257 = ~new_P3_U3442 | ~new_P3_R1054_U62;
  assign new_P3_R1054_U258 = ~new_P3_U3564 | ~new_P3_R1054_U92;
  assign new_P3_R1054_U259 = ~new_P3_R1054_U82;
  assign new_P3_R1054_U260 = ~new_P3_R1054_U259 | ~new_P3_R1054_U187;
  assign new_P3_R1054_U261 = ~new_P3_R1054_U82 | ~new_P3_R1054_U61;
  assign new_P3_R1054_U262 = ~new_P3_U3439 | ~new_P3_R1054_U60;
  assign new_P3_R1054_U263 = ~new_P3_U3565 | ~new_P3_R1054_U59;
  assign new_P3_R1054_U264 = ~new_P3_R1054_U83;
  assign new_P3_R1054_U265 = ~new_P3_R1054_U183 | ~new_P3_R1054_U264;
  assign new_P3_R1054_U266 = ~new_P3_R1054_U83 | ~new_P3_R1054_U93;
  assign new_P3_R1054_U267 = ~new_P3_U3436 | ~new_P3_R1054_U55;
  assign new_P3_R1054_U268 = ~new_P3_U3566 | ~new_P3_R1054_U52;
  assign new_P3_R1054_U269 = ~new_P3_R1054_U268 | ~new_P3_R1054_U267;
  assign new_P3_R1054_U270 = ~new_P3_U3433 | ~new_P3_R1054_U56;
  assign new_P3_R1054_U271 = ~new_P3_U3567 | ~new_P3_R1054_U53;
  assign new_P3_R1054_U272 = ~new_P3_R1054_U201 | ~new_P3_R1054_U63;
  assign new_P3_R1054_U273 = ~new_P3_R1054_U193 | ~new_P3_R1054_U271 | ~new_P3_R1054_U270;
  assign new_P3_R1054_U274 = ~new_P3_U3430 | ~new_P3_R1054_U57;
  assign new_P3_R1054_U275 = ~new_P3_U3568 | ~new_P3_R1054_U54;
  assign new_P3_R1054_U276 = ~new_P3_R1054_U202 | ~new_P3_R1054_U94;
  assign new_P3_R1054_U277 = ~new_P3_R1054_U173 | ~new_P3_R1054_U275 | ~new_P3_R1054_U274;
  assign new_P3_R1054_U278 = ~new_P3_U3427 | ~new_P3_R1054_U51;
  assign new_P3_R1054_U279 = ~new_P3_U3569 | ~new_P3_R1054_U50;
  assign new_P3_R1054_U280 = ~new_P3_R1054_U84;
  assign new_P3_R1054_U281 = ~new_P3_R1054_U169 | ~new_P3_R1054_U280;
  assign new_P3_R1054_U282 = ~new_P3_R1054_U84 | ~new_P3_R1054_U95;
  assign new_P3_R1054_U283 = ~new_P3_U3424 | ~new_P3_R1054_U49;
  assign new_P3_R1054_U284 = ~new_P3_U3570 | ~new_P3_R1054_U48;
  assign new_P3_R1054_U285 = ~new_P3_R1054_U85;
  assign new_P3_R1054_U286 = ~new_P3_R1054_U165 | ~new_P3_R1054_U285;
  assign new_P3_R1054_U287 = ~new_P3_R1054_U85 | ~new_P3_R1054_U96;
  assign new_P3_R1054_U288 = ~new_P3_U3421 | ~new_P3_R1054_U45;
  assign new_P3_R1054_U289 = ~new_P3_U3571 | ~new_P3_R1054_U43;
  assign new_P3_R1054_U290 = ~new_P3_R1054_U289 | ~new_P3_R1054_U288;
  assign new_P3_R1054_U291 = ~new_P3_U3418 | ~new_P3_R1054_U46;
  assign new_P3_R1054_U292 = ~new_P3_U3572 | ~new_P3_R1054_U44;
  assign new_P3_R1054_U293 = ~new_P3_R1054_U212 | ~new_P3_R1054_U64;
  assign new_P3_R1054_U294 = ~new_P3_R1054_U204 | ~new_P3_R1054_U292 | ~new_P3_R1054_U291;
  assign new_P3_R1161_U4 = new_P3_R1161_U179 & new_P3_R1161_U178;
  assign new_P3_R1161_U5 = new_P3_R1161_U197 & new_P3_R1161_U196;
  assign new_P3_R1161_U6 = new_P3_R1161_U237 & new_P3_R1161_U236;
  assign new_P3_R1161_U7 = new_P3_R1161_U246 & new_P3_R1161_U245;
  assign new_P3_R1161_U8 = new_P3_R1161_U264 & new_P3_R1161_U263;
  assign new_P3_R1161_U9 = new_P3_R1161_U272 & new_P3_R1161_U271;
  assign new_P3_R1161_U10 = new_P3_R1161_U351 & new_P3_R1161_U348;
  assign new_P3_R1161_U11 = new_P3_R1161_U344 & new_P3_R1161_U341;
  assign new_P3_R1161_U12 = new_P3_R1161_U335 & new_P3_R1161_U332;
  assign new_P3_R1161_U13 = new_P3_R1161_U326 & new_P3_R1161_U323;
  assign new_P3_R1161_U14 = new_P3_R1161_U320 & new_P3_R1161_U318;
  assign new_P3_R1161_U15 = new_P3_R1161_U313 & new_P3_R1161_U310;
  assign new_P3_R1161_U16 = new_P3_R1161_U235 & new_P3_R1161_U232;
  assign new_P3_R1161_U17 = new_P3_R1161_U227 & new_P3_R1161_U224;
  assign new_P3_R1161_U18 = new_P3_R1161_U213 & new_P3_R1161_U210;
  assign new_P3_R1161_U19 = ~new_P3_U3407;
  assign new_P3_R1161_U20 = ~new_P3_U3070;
  assign new_P3_R1161_U21 = ~new_P3_U3069;
  assign new_P3_R1161_U22 = ~new_P3_U3070 | ~new_P3_U3407;
  assign new_P3_R1161_U23 = ~new_P3_U3410;
  assign new_P3_R1161_U24 = ~new_P3_U3401;
  assign new_P3_R1161_U25 = ~new_P3_U3059;
  assign new_P3_R1161_U26 = ~new_P3_U3066;
  assign new_P3_R1161_U27 = ~new_P3_U3395;
  assign new_P3_R1161_U28 = ~new_P3_U3067;
  assign new_P3_R1161_U29 = ~new_P3_U3387;
  assign new_P3_R1161_U30 = ~new_P3_U3076;
  assign new_P3_R1161_U31 = ~new_P3_U3076 | ~new_P3_U3387;
  assign new_P3_R1161_U32 = ~new_P3_U3398;
  assign new_P3_R1161_U33 = ~new_P3_U3063;
  assign new_P3_R1161_U34 = ~new_P3_U3059 | ~new_P3_U3401;
  assign new_P3_R1161_U35 = ~new_P3_U3404;
  assign new_P3_R1161_U36 = ~new_P3_U3413;
  assign new_P3_R1161_U37 = ~new_P3_U3083;
  assign new_P3_R1161_U38 = ~new_P3_U3082;
  assign new_P3_R1161_U39 = ~new_P3_U3416;
  assign new_P3_R1161_U40 = ~new_P3_R1161_U63 | ~new_P3_R1161_U205;
  assign new_P3_R1161_U41 = ~new_P3_R1161_U117 | ~new_P3_R1161_U193;
  assign new_P3_R1161_U42 = ~new_P3_R1161_U182 | ~new_P3_R1161_U183;
  assign new_P3_R1161_U43 = ~new_P3_U3392 | ~new_P3_U3077;
  assign new_P3_R1161_U44 = ~new_P3_R1161_U122 | ~new_P3_R1161_U219;
  assign new_P3_R1161_U45 = ~new_P3_R1161_U216 | ~new_P3_R1161_U215;
  assign new_P3_R1161_U46 = ~new_P3_U3900;
  assign new_P3_R1161_U47 = ~new_P3_U3052;
  assign new_P3_R1161_U48 = ~new_P3_U3056;
  assign new_P3_R1161_U49 = ~new_P3_U3901;
  assign new_P3_R1161_U50 = ~new_P3_U3902;
  assign new_P3_R1161_U51 = ~new_P3_U3057;
  assign new_P3_R1161_U52 = ~new_P3_U3903;
  assign new_P3_R1161_U53 = ~new_P3_U3064;
  assign new_P3_R1161_U54 = ~new_P3_U3906;
  assign new_P3_R1161_U55 = ~new_P3_U3074;
  assign new_P3_R1161_U56 = ~new_P3_U3437;
  assign new_P3_R1161_U57 = ~new_P3_U3072;
  assign new_P3_R1161_U58 = ~new_P3_U3068;
  assign new_P3_R1161_U59 = ~new_P3_U3072 | ~new_P3_U3437;
  assign new_P3_R1161_U60 = ~new_P3_U3440;
  assign new_P3_R1161_U61 = ~new_P3_U3419;
  assign new_P3_R1161_U62 = ~new_P3_U3061;
  assign new_P3_R1161_U63 = ~new_P3_U3083 | ~new_P3_U3413;
  assign new_P3_R1161_U64 = ~new_P3_U3425;
  assign new_P3_R1161_U65 = ~new_P3_U3071;
  assign new_P3_R1161_U66 = ~new_P3_U3422;
  assign new_P3_R1161_U67 = ~new_P3_U3062;
  assign new_P3_R1161_U68 = ~new_P3_U3062 | ~new_P3_U3422;
  assign new_P3_R1161_U69 = ~new_P3_U3428;
  assign new_P3_R1161_U70 = ~new_P3_U3079;
  assign new_P3_R1161_U71 = ~new_P3_U3431;
  assign new_P3_R1161_U72 = ~new_P3_U3078;
  assign new_P3_R1161_U73 = ~new_P3_U3434;
  assign new_P3_R1161_U74 = ~new_P3_U3073;
  assign new_P3_R1161_U75 = ~new_P3_U3443;
  assign new_P3_R1161_U76 = ~new_P3_U3081;
  assign new_P3_R1161_U77 = ~new_P3_U3081 | ~new_P3_U3443;
  assign new_P3_R1161_U78 = ~new_P3_U3445;
  assign new_P3_R1161_U79 = ~new_P3_U3080;
  assign new_P3_R1161_U80 = ~new_P3_U3080 | ~new_P3_U3445;
  assign new_P3_R1161_U81 = ~new_P3_U3907;
  assign new_P3_R1161_U82 = ~new_P3_U3905;
  assign new_P3_R1161_U83 = ~new_P3_U3060;
  assign new_P3_R1161_U84 = ~new_P3_U3904;
  assign new_P3_R1161_U85 = ~new_P3_U3065;
  assign new_P3_R1161_U86 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1161_U87 = ~new_P3_U3053;
  assign new_P3_R1161_U88 = ~new_P3_U3899;
  assign new_P3_R1161_U89 = ~new_P3_R1161_U306 | ~new_P3_R1161_U176;
  assign new_P3_R1161_U90 = ~new_P3_U3075;
  assign new_P3_R1161_U91 = ~new_P3_R1161_U77 | ~new_P3_R1161_U315;
  assign new_P3_R1161_U92 = ~new_P3_R1161_U261 | ~new_P3_R1161_U260;
  assign new_P3_R1161_U93 = ~new_P3_R1161_U68 | ~new_P3_R1161_U337;
  assign new_P3_R1161_U94 = ~new_P3_R1161_U457 | ~new_P3_R1161_U456;
  assign new_P3_R1161_U95 = ~new_P3_R1161_U504 | ~new_P3_R1161_U503;
  assign new_P3_R1161_U96 = ~new_P3_R1161_U375 | ~new_P3_R1161_U374;
  assign new_P3_R1161_U97 = ~new_P3_R1161_U380 | ~new_P3_R1161_U379;
  assign new_P3_R1161_U98 = ~new_P3_R1161_U387 | ~new_P3_R1161_U386;
  assign new_P3_R1161_U99 = ~new_P3_R1161_U394 | ~new_P3_R1161_U393;
  assign new_P3_R1161_U100 = ~new_P3_R1161_U399 | ~new_P3_R1161_U398;
  assign new_P3_R1161_U101 = ~new_P3_R1161_U408 | ~new_P3_R1161_U407;
  assign new_P3_R1161_U102 = ~new_P3_R1161_U415 | ~new_P3_R1161_U414;
  assign new_P3_R1161_U103 = ~new_P3_R1161_U422 | ~new_P3_R1161_U421;
  assign new_P3_R1161_U104 = ~new_P3_R1161_U429 | ~new_P3_R1161_U428;
  assign new_P3_R1161_U105 = ~new_P3_R1161_U434 | ~new_P3_R1161_U433;
  assign new_P3_R1161_U106 = ~new_P3_R1161_U441 | ~new_P3_R1161_U440;
  assign new_P3_R1161_U107 = ~new_P3_R1161_U448 | ~new_P3_R1161_U447;
  assign new_P3_R1161_U108 = ~new_P3_R1161_U462 | ~new_P3_R1161_U461;
  assign new_P3_R1161_U109 = ~new_P3_R1161_U467 | ~new_P3_R1161_U466;
  assign new_P3_R1161_U110 = ~new_P3_R1161_U474 | ~new_P3_R1161_U473;
  assign new_P3_R1161_U111 = ~new_P3_R1161_U481 | ~new_P3_R1161_U480;
  assign new_P3_R1161_U112 = ~new_P3_R1161_U488 | ~new_P3_R1161_U487;
  assign new_P3_R1161_U113 = ~new_P3_R1161_U495 | ~new_P3_R1161_U494;
  assign new_P3_R1161_U114 = ~new_P3_R1161_U500 | ~new_P3_R1161_U499;
  assign new_P3_R1161_U115 = new_P3_R1161_U189 & new_P3_R1161_U187;
  assign new_P3_R1161_U116 = new_P3_R1161_U4 & new_P3_R1161_U180;
  assign new_P3_R1161_U117 = new_P3_R1161_U194 & new_P3_R1161_U192;
  assign new_P3_R1161_U118 = new_P3_R1161_U201 & new_P3_R1161_U200;
  assign new_P3_R1161_U119 = new_P3_R1161_U22 & new_P3_R1161_U382 & new_P3_R1161_U381;
  assign new_P3_R1161_U120 = new_P3_R1161_U212 & new_P3_R1161_U5;
  assign new_P3_R1161_U121 = new_P3_R1161_U181 & new_P3_R1161_U180;
  assign new_P3_R1161_U122 = new_P3_R1161_U220 & new_P3_R1161_U218;
  assign new_P3_R1161_U123 = new_P3_R1161_U34 & new_P3_R1161_U389 & new_P3_R1161_U388;
  assign new_P3_R1161_U124 = new_P3_R1161_U226 & new_P3_R1161_U4;
  assign new_P3_R1161_U125 = new_P3_R1161_U234 & new_P3_R1161_U181;
  assign new_P3_R1161_U126 = new_P3_R1161_U204 & new_P3_R1161_U6;
  assign new_P3_R1161_U127 = new_P3_R1161_U243 & new_P3_R1161_U239;
  assign new_P3_R1161_U128 = new_P3_R1161_U250 & new_P3_R1161_U7;
  assign new_P3_R1161_U129 = new_P3_R1161_U248 & new_P3_R1161_U172;
  assign new_P3_R1161_U130 = new_P3_R1161_U268 & new_P3_R1161_U267;
  assign new_P3_R1161_U131 = new_P3_R1161_U273 & new_P3_R1161_U9 & new_P3_R1161_U282;
  assign new_P3_R1161_U132 = new_P3_R1161_U285 & new_P3_R1161_U280;
  assign new_P3_R1161_U133 = new_P3_R1161_U301 & new_P3_R1161_U298;
  assign new_P3_R1161_U134 = new_P3_R1161_U368 & new_P3_R1161_U302;
  assign new_P3_R1161_U135 = new_P3_R1161_U160 & new_P3_R1161_U278;
  assign new_P3_R1161_U136 = new_P3_R1161_U80 & new_P3_R1161_U455 & new_P3_R1161_U454;
  assign new_P3_R1161_U137 = new_P3_R1161_U325 & new_P3_R1161_U9;
  assign new_P3_R1161_U138 = new_P3_R1161_U59 & new_P3_R1161_U469 & new_P3_R1161_U468;
  assign new_P3_R1161_U139 = new_P3_R1161_U334 & new_P3_R1161_U8;
  assign new_P3_R1161_U140 = new_P3_R1161_U172 & new_P3_R1161_U490 & new_P3_R1161_U489;
  assign new_P3_R1161_U141 = new_P3_R1161_U343 & new_P3_R1161_U7;
  assign new_P3_R1161_U142 = new_P3_R1161_U171 & new_P3_R1161_U502 & new_P3_R1161_U501;
  assign new_P3_R1161_U143 = new_P3_R1161_U350 & new_P3_R1161_U6;
  assign new_P3_R1161_U144 = ~new_P3_R1161_U118 | ~new_P3_R1161_U202;
  assign new_P3_R1161_U145 = ~new_P3_R1161_U217 | ~new_P3_R1161_U229;
  assign new_P3_R1161_U146 = ~new_P3_U3054;
  assign new_P3_R1161_U147 = ~new_P3_U3908;
  assign new_P3_R1161_U148 = new_P3_R1161_U403 & new_P3_R1161_U402;
  assign new_P3_R1161_U149 = ~new_P3_R1161_U364 | ~new_P3_R1161_U304 | ~new_P3_R1161_U169;
  assign new_P3_R1161_U150 = new_P3_R1161_U410 & new_P3_R1161_U409;
  assign new_P3_R1161_U151 = ~new_P3_R1161_U134 | ~new_P3_R1161_U370 | ~new_P3_R1161_U369;
  assign new_P3_R1161_U152 = new_P3_R1161_U417 & new_P3_R1161_U416;
  assign new_P3_R1161_U153 = ~new_P3_R1161_U86 | ~new_P3_R1161_U365 | ~new_P3_R1161_U299;
  assign new_P3_R1161_U154 = new_P3_R1161_U424 & new_P3_R1161_U423;
  assign new_P3_R1161_U155 = ~new_P3_R1161_U293 | ~new_P3_R1161_U292;
  assign new_P3_R1161_U156 = new_P3_R1161_U436 & new_P3_R1161_U435;
  assign new_P3_R1161_U157 = ~new_P3_R1161_U289 | ~new_P3_R1161_U288;
  assign new_P3_R1161_U158 = new_P3_R1161_U443 & new_P3_R1161_U442;
  assign new_P3_R1161_U159 = ~new_P3_R1161_U132 | ~new_P3_R1161_U284;
  assign new_P3_R1161_U160 = new_P3_R1161_U450 & new_P3_R1161_U449;
  assign new_P3_R1161_U161 = ~new_P3_R1161_U43 | ~new_P3_R1161_U327;
  assign new_P3_R1161_U162 = ~new_P3_R1161_U130 | ~new_P3_R1161_U269;
  assign new_P3_R1161_U163 = new_P3_R1161_U476 & new_P3_R1161_U475;
  assign new_P3_R1161_U164 = ~new_P3_R1161_U257 | ~new_P3_R1161_U256;
  assign new_P3_R1161_U165 = new_P3_R1161_U483 & new_P3_R1161_U482;
  assign new_P3_R1161_U166 = ~new_P3_R1161_U253 | ~new_P3_R1161_U252;
  assign new_P3_R1161_U167 = ~new_P3_R1161_U127 | ~new_P3_R1161_U242;
  assign new_P3_R1161_U168 = ~new_P3_R1161_U367 | ~new_P3_R1161_U366;
  assign new_P3_R1161_U169 = ~new_P3_U3053 | ~new_P3_R1161_U151;
  assign new_P3_R1161_U170 = ~new_P3_R1161_U34;
  assign new_P3_R1161_U171 = ~new_P3_U3416 | ~new_P3_U3082;
  assign new_P3_R1161_U172 = ~new_P3_U3071 | ~new_P3_U3425;
  assign new_P3_R1161_U173 = ~new_P3_U3057 | ~new_P3_U3902;
  assign new_P3_R1161_U174 = ~new_P3_R1161_U68;
  assign new_P3_R1161_U175 = ~new_P3_R1161_U77;
  assign new_P3_R1161_U176 = ~new_P3_U3064 | ~new_P3_U3903;
  assign new_P3_R1161_U177 = ~new_P3_R1161_U63;
  assign new_P3_R1161_U178 = new_P3_U3066 | new_P3_U3404;
  assign new_P3_R1161_U179 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1161_U180 = new_P3_U3398 | new_P3_U3063;
  assign new_P3_R1161_U181 = new_P3_U3395 | new_P3_U3067;
  assign new_P3_R1161_U182 = ~new_P3_R1161_U31;
  assign new_P3_R1161_U183 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1161_U184 = ~new_P3_R1161_U42;
  assign new_P3_R1161_U185 = ~new_P3_R1161_U43;
  assign new_P3_R1161_U186 = ~new_P3_R1161_U42 | ~new_P3_R1161_U43;
  assign new_P3_R1161_U187 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1161_U188 = ~new_P3_R1161_U186 | ~new_P3_R1161_U181;
  assign new_P3_R1161_U189 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1161_U190 = ~new_P3_R1161_U115 | ~new_P3_R1161_U188;
  assign new_P3_R1161_U191 = ~new_P3_R1161_U35 | ~new_P3_R1161_U34;
  assign new_P3_R1161_U192 = ~new_P3_U3066 | ~new_P3_R1161_U191;
  assign new_P3_R1161_U193 = ~new_P3_R1161_U116 | ~new_P3_R1161_U190;
  assign new_P3_R1161_U194 = ~new_P3_U3404 | ~new_P3_R1161_U170;
  assign new_P3_R1161_U195 = ~new_P3_R1161_U41;
  assign new_P3_R1161_U196 = new_P3_U3069 | new_P3_U3410;
  assign new_P3_R1161_U197 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1161_U198 = ~new_P3_R1161_U22;
  assign new_P3_R1161_U199 = ~new_P3_R1161_U23 | ~new_P3_R1161_U22;
  assign new_P3_R1161_U200 = ~new_P3_U3069 | ~new_P3_R1161_U199;
  assign new_P3_R1161_U201 = ~new_P3_U3410 | ~new_P3_R1161_U198;
  assign new_P3_R1161_U202 = ~new_P3_R1161_U5 | ~new_P3_R1161_U41;
  assign new_P3_R1161_U203 = ~new_P3_R1161_U144;
  assign new_P3_R1161_U204 = new_P3_U3413 | new_P3_U3083;
  assign new_P3_R1161_U205 = ~new_P3_R1161_U204 | ~new_P3_R1161_U144;
  assign new_P3_R1161_U206 = ~new_P3_R1161_U40;
  assign new_P3_R1161_U207 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1161_U208 = new_P3_U3407 | new_P3_U3070;
  assign new_P3_R1161_U209 = ~new_P3_R1161_U208 | ~new_P3_R1161_U41;
  assign new_P3_R1161_U210 = ~new_P3_R1161_U119 | ~new_P3_R1161_U209;
  assign new_P3_R1161_U211 = ~new_P3_R1161_U195 | ~new_P3_R1161_U22;
  assign new_P3_R1161_U212 = ~new_P3_U3410 | ~new_P3_U3069;
  assign new_P3_R1161_U213 = ~new_P3_R1161_U120 | ~new_P3_R1161_U211;
  assign new_P3_R1161_U214 = new_P3_U3070 | new_P3_U3407;
  assign new_P3_R1161_U215 = ~new_P3_R1161_U185 | ~new_P3_R1161_U181;
  assign new_P3_R1161_U216 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1161_U217 = ~new_P3_R1161_U45;
  assign new_P3_R1161_U218 = ~new_P3_R1161_U121 | ~new_P3_R1161_U184;
  assign new_P3_R1161_U219 = ~new_P3_R1161_U45 | ~new_P3_R1161_U180;
  assign new_P3_R1161_U220 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1161_U221 = ~new_P3_R1161_U44;
  assign new_P3_R1161_U222 = new_P3_U3401 | new_P3_U3059;
  assign new_P3_R1161_U223 = ~new_P3_R1161_U222 | ~new_P3_R1161_U44;
  assign new_P3_R1161_U224 = ~new_P3_R1161_U123 | ~new_P3_R1161_U223;
  assign new_P3_R1161_U225 = ~new_P3_R1161_U221 | ~new_P3_R1161_U34;
  assign new_P3_R1161_U226 = ~new_P3_U3404 | ~new_P3_U3066;
  assign new_P3_R1161_U227 = ~new_P3_R1161_U124 | ~new_P3_R1161_U225;
  assign new_P3_R1161_U228 = new_P3_U3059 | new_P3_U3401;
  assign new_P3_R1161_U229 = ~new_P3_R1161_U184 | ~new_P3_R1161_U181;
  assign new_P3_R1161_U230 = ~new_P3_R1161_U145;
  assign new_P3_R1161_U231 = ~new_P3_U3063 | ~new_P3_U3398;
  assign new_P3_R1161_U232 = ~new_P3_R1161_U42 | ~new_P3_R1161_U43 | ~new_P3_R1161_U401 | ~new_P3_R1161_U400;
  assign new_P3_R1161_U233 = ~new_P3_R1161_U43 | ~new_P3_R1161_U42;
  assign new_P3_R1161_U234 = ~new_P3_U3067 | ~new_P3_U3395;
  assign new_P3_R1161_U235 = ~new_P3_R1161_U125 | ~new_P3_R1161_U233;
  assign new_P3_R1161_U236 = new_P3_U3082 | new_P3_U3416;
  assign new_P3_R1161_U237 = new_P3_U3061 | new_P3_U3419;
  assign new_P3_R1161_U238 = ~new_P3_R1161_U177 | ~new_P3_R1161_U6;
  assign new_P3_R1161_U239 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1161_U240 = ~new_P3_R1161_U171 | ~new_P3_R1161_U238;
  assign new_P3_R1161_U241 = new_P3_U3419 | new_P3_U3061;
  assign new_P3_R1161_U242 = ~new_P3_R1161_U126 | ~new_P3_R1161_U144;
  assign new_P3_R1161_U243 = ~new_P3_R1161_U241 | ~new_P3_R1161_U240;
  assign new_P3_R1161_U244 = ~new_P3_R1161_U167;
  assign new_P3_R1161_U245 = new_P3_U3079 | new_P3_U3428;
  assign new_P3_R1161_U246 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1161_U247 = ~new_P3_R1161_U174 | ~new_P3_R1161_U7;
  assign new_P3_R1161_U248 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1161_U249 = ~new_P3_R1161_U129 | ~new_P3_R1161_U247;
  assign new_P3_R1161_U250 = new_P3_U3422 | new_P3_U3062;
  assign new_P3_R1161_U251 = new_P3_U3428 | new_P3_U3079;
  assign new_P3_R1161_U252 = ~new_P3_R1161_U128 | ~new_P3_R1161_U167;
  assign new_P3_R1161_U253 = ~new_P3_R1161_U251 | ~new_P3_R1161_U249;
  assign new_P3_R1161_U254 = ~new_P3_R1161_U166;
  assign new_P3_R1161_U255 = new_P3_U3431 | new_P3_U3078;
  assign new_P3_R1161_U256 = ~new_P3_R1161_U255 | ~new_P3_R1161_U166;
  assign new_P3_R1161_U257 = ~new_P3_U3078 | ~new_P3_U3431;
  assign new_P3_R1161_U258 = ~new_P3_R1161_U164;
  assign new_P3_R1161_U259 = new_P3_U3434 | new_P3_U3073;
  assign new_P3_R1161_U260 = ~new_P3_R1161_U259 | ~new_P3_R1161_U164;
  assign new_P3_R1161_U261 = ~new_P3_U3073 | ~new_P3_U3434;
  assign new_P3_R1161_U262 = ~new_P3_R1161_U92;
  assign new_P3_R1161_U263 = new_P3_U3068 | new_P3_U3440;
  assign new_P3_R1161_U264 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1161_U265 = ~new_P3_R1161_U59;
  assign new_P3_R1161_U266 = ~new_P3_R1161_U60 | ~new_P3_R1161_U59;
  assign new_P3_R1161_U267 = ~new_P3_U3068 | ~new_P3_R1161_U266;
  assign new_P3_R1161_U268 = ~new_P3_U3440 | ~new_P3_R1161_U265;
  assign new_P3_R1161_U269 = ~new_P3_R1161_U8 | ~new_P3_R1161_U92;
  assign new_P3_R1161_U270 = ~new_P3_R1161_U162;
  assign new_P3_R1161_U271 = new_P3_U3075 | new_P3_U3907;
  assign new_P3_R1161_U272 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1161_U273 = new_P3_U3074 | new_P3_U3906;
  assign new_P3_R1161_U274 = ~new_P3_R1161_U80;
  assign new_P3_R1161_U275 = ~new_P3_U3907 | ~new_P3_R1161_U274;
  assign new_P3_R1161_U276 = ~new_P3_R1161_U275 | ~new_P3_R1161_U90;
  assign new_P3_R1161_U277 = ~new_P3_R1161_U80 | ~new_P3_R1161_U81;
  assign new_P3_R1161_U278 = ~new_P3_R1161_U277 | ~new_P3_R1161_U276;
  assign new_P3_R1161_U279 = ~new_P3_R1161_U175 | ~new_P3_R1161_U9;
  assign new_P3_R1161_U280 = ~new_P3_U3074 | ~new_P3_U3906;
  assign new_P3_R1161_U281 = ~new_P3_R1161_U278 | ~new_P3_R1161_U279;
  assign new_P3_R1161_U282 = new_P3_U3443 | new_P3_U3081;
  assign new_P3_R1161_U283 = new_P3_U3906 | new_P3_U3074;
  assign new_P3_R1161_U284 = ~new_P3_R1161_U162 | ~new_P3_R1161_U131;
  assign new_P3_R1161_U285 = ~new_P3_R1161_U283 | ~new_P3_R1161_U281;
  assign new_P3_R1161_U286 = ~new_P3_R1161_U159;
  assign new_P3_R1161_U287 = new_P3_U3905 | new_P3_U3060;
  assign new_P3_R1161_U288 = ~new_P3_R1161_U287 | ~new_P3_R1161_U159;
  assign new_P3_R1161_U289 = ~new_P3_U3060 | ~new_P3_U3905;
  assign new_P3_R1161_U290 = ~new_P3_R1161_U157;
  assign new_P3_R1161_U291 = new_P3_U3904 | new_P3_U3065;
  assign new_P3_R1161_U292 = ~new_P3_R1161_U291 | ~new_P3_R1161_U157;
  assign new_P3_R1161_U293 = ~new_P3_U3065 | ~new_P3_U3904;
  assign new_P3_R1161_U294 = ~new_P3_R1161_U155;
  assign new_P3_R1161_U295 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1161_U296 = ~new_P3_R1161_U176 | ~new_P3_R1161_U173;
  assign new_P3_R1161_U297 = ~new_P3_R1161_U86;
  assign new_P3_R1161_U298 = new_P3_U3903 | new_P3_U3064;
  assign new_P3_R1161_U299 = ~new_P3_R1161_U168 | ~new_P3_R1161_U155 | ~new_P3_R1161_U298;
  assign new_P3_R1161_U300 = ~new_P3_R1161_U153;
  assign new_P3_R1161_U301 = new_P3_U3900 | new_P3_U3052;
  assign new_P3_R1161_U302 = ~new_P3_U3052 | ~new_P3_U3900;
  assign new_P3_R1161_U303 = ~new_P3_R1161_U151;
  assign new_P3_R1161_U304 = ~new_P3_U3899 | ~new_P3_R1161_U151;
  assign new_P3_R1161_U305 = ~new_P3_R1161_U149;
  assign new_P3_R1161_U306 = ~new_P3_R1161_U298 | ~new_P3_R1161_U155;
  assign new_P3_R1161_U307 = ~new_P3_R1161_U89;
  assign new_P3_R1161_U308 = new_P3_U3902 | new_P3_U3057;
  assign new_P3_R1161_U309 = ~new_P3_R1161_U308 | ~new_P3_R1161_U89;
  assign new_P3_R1161_U310 = ~new_P3_R1161_U154 | ~new_P3_R1161_U309 | ~new_P3_R1161_U173;
  assign new_P3_R1161_U311 = ~new_P3_R1161_U307 | ~new_P3_R1161_U173;
  assign new_P3_R1161_U312 = ~new_P3_U3901 | ~new_P3_U3056;
  assign new_P3_R1161_U313 = ~new_P3_R1161_U168 | ~new_P3_R1161_U311 | ~new_P3_R1161_U312;
  assign new_P3_R1161_U314 = new_P3_U3057 | new_P3_U3902;
  assign new_P3_R1161_U315 = ~new_P3_R1161_U282 | ~new_P3_R1161_U162;
  assign new_P3_R1161_U316 = ~new_P3_R1161_U91;
  assign new_P3_R1161_U317 = ~new_P3_R1161_U9 | ~new_P3_R1161_U91;
  assign new_P3_R1161_U318 = ~new_P3_R1161_U135 | ~new_P3_R1161_U317;
  assign new_P3_R1161_U319 = ~new_P3_R1161_U317 | ~new_P3_R1161_U278;
  assign new_P3_R1161_U320 = ~new_P3_R1161_U453 | ~new_P3_R1161_U319;
  assign new_P3_R1161_U321 = new_P3_U3445 | new_P3_U3080;
  assign new_P3_R1161_U322 = ~new_P3_R1161_U321 | ~new_P3_R1161_U91;
  assign new_P3_R1161_U323 = ~new_P3_R1161_U136 | ~new_P3_R1161_U322;
  assign new_P3_R1161_U324 = ~new_P3_R1161_U316 | ~new_P3_R1161_U80;
  assign new_P3_R1161_U325 = ~new_P3_U3075 | ~new_P3_U3907;
  assign new_P3_R1161_U326 = ~new_P3_R1161_U137 | ~new_P3_R1161_U324;
  assign new_P3_R1161_U327 = new_P3_U3392 | new_P3_U3077;
  assign new_P3_R1161_U328 = ~new_P3_R1161_U161;
  assign new_P3_R1161_U329 = new_P3_U3080 | new_P3_U3445;
  assign new_P3_R1161_U330 = new_P3_U3437 | new_P3_U3072;
  assign new_P3_R1161_U331 = ~new_P3_R1161_U330 | ~new_P3_R1161_U92;
  assign new_P3_R1161_U332 = ~new_P3_R1161_U138 | ~new_P3_R1161_U331;
  assign new_P3_R1161_U333 = ~new_P3_R1161_U262 | ~new_P3_R1161_U59;
  assign new_P3_R1161_U334 = ~new_P3_U3440 | ~new_P3_U3068;
  assign new_P3_R1161_U335 = ~new_P3_R1161_U139 | ~new_P3_R1161_U333;
  assign new_P3_R1161_U336 = new_P3_U3072 | new_P3_U3437;
  assign new_P3_R1161_U337 = ~new_P3_R1161_U250 | ~new_P3_R1161_U167;
  assign new_P3_R1161_U338 = ~new_P3_R1161_U93;
  assign new_P3_R1161_U339 = new_P3_U3425 | new_P3_U3071;
  assign new_P3_R1161_U340 = ~new_P3_R1161_U339 | ~new_P3_R1161_U93;
  assign new_P3_R1161_U341 = ~new_P3_R1161_U140 | ~new_P3_R1161_U340;
  assign new_P3_R1161_U342 = ~new_P3_R1161_U338 | ~new_P3_R1161_U172;
  assign new_P3_R1161_U343 = ~new_P3_U3079 | ~new_P3_U3428;
  assign new_P3_R1161_U344 = ~new_P3_R1161_U141 | ~new_P3_R1161_U342;
  assign new_P3_R1161_U345 = new_P3_U3071 | new_P3_U3425;
  assign new_P3_R1161_U346 = new_P3_U3416 | new_P3_U3082;
  assign new_P3_R1161_U347 = ~new_P3_R1161_U346 | ~new_P3_R1161_U40;
  assign new_P3_R1161_U348 = ~new_P3_R1161_U142 | ~new_P3_R1161_U347;
  assign new_P3_R1161_U349 = ~new_P3_R1161_U206 | ~new_P3_R1161_U171;
  assign new_P3_R1161_U350 = ~new_P3_U3061 | ~new_P3_U3419;
  assign new_P3_R1161_U351 = ~new_P3_R1161_U143 | ~new_P3_R1161_U349;
  assign new_P3_R1161_U352 = ~new_P3_R1161_U207 | ~new_P3_R1161_U171;
  assign new_P3_R1161_U353 = ~new_P3_R1161_U204 | ~new_P3_R1161_U63;
  assign new_P3_R1161_U354 = ~new_P3_R1161_U214 | ~new_P3_R1161_U22;
  assign new_P3_R1161_U355 = ~new_P3_R1161_U228 | ~new_P3_R1161_U34;
  assign new_P3_R1161_U356 = ~new_P3_R1161_U231 | ~new_P3_R1161_U180;
  assign new_P3_R1161_U357 = ~new_P3_R1161_U314 | ~new_P3_R1161_U173;
  assign new_P3_R1161_U358 = ~new_P3_R1161_U298 | ~new_P3_R1161_U176;
  assign new_P3_R1161_U359 = ~new_P3_R1161_U329 | ~new_P3_R1161_U80;
  assign new_P3_R1161_U360 = ~new_P3_R1161_U282 | ~new_P3_R1161_U77;
  assign new_P3_R1161_U361 = ~new_P3_R1161_U336 | ~new_P3_R1161_U59;
  assign new_P3_R1161_U362 = ~new_P3_R1161_U345 | ~new_P3_R1161_U172;
  assign new_P3_R1161_U363 = ~new_P3_R1161_U250 | ~new_P3_R1161_U68;
  assign new_P3_R1161_U364 = ~new_P3_U3899 | ~new_P3_U3053;
  assign new_P3_R1161_U365 = ~new_P3_R1161_U296 | ~new_P3_R1161_U168;
  assign new_P3_R1161_U366 = ~new_P3_U3056 | ~new_P3_R1161_U295;
  assign new_P3_R1161_U367 = ~new_P3_U3901 | ~new_P3_R1161_U295;
  assign new_P3_R1161_U368 = ~new_P3_R1161_U301 | ~new_P3_R1161_U296 | ~new_P3_R1161_U168;
  assign new_P3_R1161_U369 = ~new_P3_R1161_U133 | ~new_P3_R1161_U155 | ~new_P3_R1161_U168;
  assign new_P3_R1161_U370 = ~new_P3_R1161_U297 | ~new_P3_R1161_U301;
  assign new_P3_R1161_U371 = ~new_P3_U3082 | ~new_P3_R1161_U39;
  assign new_P3_R1161_U372 = ~new_P3_U3416 | ~new_P3_R1161_U38;
  assign new_P3_R1161_U373 = ~new_P3_R1161_U372 | ~new_P3_R1161_U371;
  assign new_P3_R1161_U374 = ~new_P3_R1161_U352 | ~new_P3_R1161_U40;
  assign new_P3_R1161_U375 = ~new_P3_R1161_U373 | ~new_P3_R1161_U206;
  assign new_P3_R1161_U376 = ~new_P3_U3083 | ~new_P3_R1161_U36;
  assign new_P3_R1161_U377 = ~new_P3_U3413 | ~new_P3_R1161_U37;
  assign new_P3_R1161_U378 = ~new_P3_R1161_U377 | ~new_P3_R1161_U376;
  assign new_P3_R1161_U379 = ~new_P3_R1161_U353 | ~new_P3_R1161_U144;
  assign new_P3_R1161_U380 = ~new_P3_R1161_U203 | ~new_P3_R1161_U378;
  assign new_P3_R1161_U381 = ~new_P3_U3069 | ~new_P3_R1161_U23;
  assign new_P3_R1161_U382 = ~new_P3_U3410 | ~new_P3_R1161_U21;
  assign new_P3_R1161_U383 = ~new_P3_U3070 | ~new_P3_R1161_U19;
  assign new_P3_R1161_U384 = ~new_P3_U3407 | ~new_P3_R1161_U20;
  assign new_P3_R1161_U385 = ~new_P3_R1161_U384 | ~new_P3_R1161_U383;
  assign new_P3_R1161_U386 = ~new_P3_R1161_U354 | ~new_P3_R1161_U41;
  assign new_P3_R1161_U387 = ~new_P3_R1161_U385 | ~new_P3_R1161_U195;
  assign new_P3_R1161_U388 = ~new_P3_U3066 | ~new_P3_R1161_U35;
  assign new_P3_R1161_U389 = ~new_P3_U3404 | ~new_P3_R1161_U26;
  assign new_P3_R1161_U390 = ~new_P3_U3059 | ~new_P3_R1161_U24;
  assign new_P3_R1161_U391 = ~new_P3_U3401 | ~new_P3_R1161_U25;
  assign new_P3_R1161_U392 = ~new_P3_R1161_U391 | ~new_P3_R1161_U390;
  assign new_P3_R1161_U393 = ~new_P3_R1161_U355 | ~new_P3_R1161_U44;
  assign new_P3_R1161_U394 = ~new_P3_R1161_U392 | ~new_P3_R1161_U221;
  assign new_P3_R1161_U395 = ~new_P3_U3063 | ~new_P3_R1161_U32;
  assign new_P3_R1161_U396 = ~new_P3_U3398 | ~new_P3_R1161_U33;
  assign new_P3_R1161_U397 = ~new_P3_R1161_U396 | ~new_P3_R1161_U395;
  assign new_P3_R1161_U398 = ~new_P3_R1161_U356 | ~new_P3_R1161_U145;
  assign new_P3_R1161_U399 = ~new_P3_R1161_U230 | ~new_P3_R1161_U397;
  assign new_P3_R1161_U400 = ~new_P3_U3067 | ~new_P3_R1161_U27;
  assign new_P3_R1161_U401 = ~new_P3_U3395 | ~new_P3_R1161_U28;
  assign new_P3_R1161_U402 = ~new_P3_U3054 | ~new_P3_R1161_U147;
  assign new_P3_R1161_U403 = ~new_P3_U3908 | ~new_P3_R1161_U146;
  assign new_P3_R1161_U404 = ~new_P3_U3054 | ~new_P3_R1161_U147;
  assign new_P3_R1161_U405 = ~new_P3_U3908 | ~new_P3_R1161_U146;
  assign new_P3_R1161_U406 = ~new_P3_R1161_U405 | ~new_P3_R1161_U404;
  assign new_P3_R1161_U407 = ~new_P3_R1161_U148 | ~new_P3_R1161_U149;
  assign new_P3_R1161_U408 = ~new_P3_R1161_U305 | ~new_P3_R1161_U406;
  assign new_P3_R1161_U409 = ~new_P3_U3053 | ~new_P3_R1161_U88;
  assign new_P3_R1161_U410 = ~new_P3_U3899 | ~new_P3_R1161_U87;
  assign new_P3_R1161_U411 = ~new_P3_U3053 | ~new_P3_R1161_U88;
  assign new_P3_R1161_U412 = ~new_P3_U3899 | ~new_P3_R1161_U87;
  assign new_P3_R1161_U413 = ~new_P3_R1161_U412 | ~new_P3_R1161_U411;
  assign new_P3_R1161_U414 = ~new_P3_R1161_U150 | ~new_P3_R1161_U151;
  assign new_P3_R1161_U415 = ~new_P3_R1161_U303 | ~new_P3_R1161_U413;
  assign new_P3_R1161_U416 = ~new_P3_U3052 | ~new_P3_R1161_U46;
  assign new_P3_R1161_U417 = ~new_P3_U3900 | ~new_P3_R1161_U47;
  assign new_P3_R1161_U418 = ~new_P3_U3052 | ~new_P3_R1161_U46;
  assign new_P3_R1161_U419 = ~new_P3_U3900 | ~new_P3_R1161_U47;
  assign new_P3_R1161_U420 = ~new_P3_R1161_U419 | ~new_P3_R1161_U418;
  assign new_P3_R1161_U421 = ~new_P3_R1161_U152 | ~new_P3_R1161_U153;
  assign new_P3_R1161_U422 = ~new_P3_R1161_U300 | ~new_P3_R1161_U420;
  assign new_P3_R1161_U423 = ~new_P3_U3056 | ~new_P3_R1161_U49;
  assign new_P3_R1161_U424 = ~new_P3_U3901 | ~new_P3_R1161_U48;
  assign new_P3_R1161_U425 = ~new_P3_U3057 | ~new_P3_R1161_U50;
  assign new_P3_R1161_U426 = ~new_P3_U3902 | ~new_P3_R1161_U51;
  assign new_P3_R1161_U427 = ~new_P3_R1161_U426 | ~new_P3_R1161_U425;
  assign new_P3_R1161_U428 = ~new_P3_R1161_U357 | ~new_P3_R1161_U89;
  assign new_P3_R1161_U429 = ~new_P3_R1161_U427 | ~new_P3_R1161_U307;
  assign new_not_keyinput0 = ~keyinput0;
  assign new_not_keyinput1 = ~keyinput1;
  assign new_not_keyinput2 = ~keyinput2;
  assign new_not_keyinput3 = ~keyinput3;
  assign new_not_keyinput4 = ~keyinput4;
  assign new_not_keyinput5 = ~keyinput5;
  assign new_not_keyinput6 = ~keyinput6;
  assign new_not_keyinput7 = ~keyinput7;
  assign new_not_keyinput8 = ~keyinput8;
  assign new_not_keyinput9 = ~keyinput9;
  assign new_not_keyinput10 = ~keyinput10;
  assign new_not_keyinput11 = ~keyinput11;
  assign new_not_keyinput12 = ~keyinput12;
  assign new_not_keyinput13 = ~keyinput13;
  assign new_not_keyinput14 = ~keyinput14;
  assign new_not_keyinput15 = ~keyinput15;
  assign new_not_keyinput16 = ~keyinput16;
  assign new_not_keyinput17 = ~keyinput17;
  assign new_not_keyinput18 = ~keyinput18;
  assign new_not_keyinput19 = ~keyinput19;
  assign new_not_keyinput20 = ~keyinput20;
  assign new_not_keyinput21 = ~keyinput21;
  assign new_not_keyinput22 = ~keyinput22;
  assign new_not_keyinput23 = ~keyinput23;
  assign new_not_keyinput24 = ~keyinput24;
  assign new_not_keyinput25 = ~keyinput25;
  assign new_not_keyinput26 = ~keyinput26;
  assign new_not_keyinput27 = ~keyinput27;
  assign new_not_keyinput28 = ~keyinput28;
  assign new_not_keyinput29 = ~keyinput29;
  assign new_not_keyinput30 = ~keyinput30;
  assign new_not_keyinput31 = ~keyinput31;
  assign new_not_0 = ~Q_0;
  assign new_and_1 = new_not_0 & Q_4;
  assign new_not_2 = ~Q_4;
  assign new_and_3 = new_not_2 & Q_3 & Q_2 & Q_0 & Q_1;
  assign new_not_4 = ~Q_2;
  assign new_and_5 = new_not_4 & Q_4;
  assign new_not_6 = ~Q_1;
  assign new_and_7 = new_not_6 & Q_4;
  assign new_not_8 = ~Q_3;
  assign new_and_9 = new_not_8 & Q_4;
  assign n61563 = new_and_9 | new_and_7 | new_and_5 | new_and_1 | new_and_3;
  assign new_not_11 = ~Q_1;
  assign new_and_12 = new_not_11 & Q_3;
  assign new_not_13 = ~Q_3;
  assign new_and_14 = new_not_13 & Q_2 & Q_0 & Q_1;
  assign new_not_15 = ~Q_0;
  assign new_and_16 = new_not_15 & Q_3;
  assign new_not_17 = ~Q_2;
  assign new_and_18 = new_not_17 & Q_3;
  assign n61560 = new_and_18 | new_and_16 | new_and_12 | new_and_14;
  assign new_not_20 = ~Q_0;
  assign new_and_21 = new_not_20 & Q_2;
  assign new_not_22 = ~Q_1;
  assign new_and_23 = new_not_22 & Q_2;
  assign new_not_24 = ~Q_2;
  assign new_and_25 = new_not_24 & Q_0 & Q_1;
  assign n61557 = new_and_25 | new_and_21 | new_and_23;
  assign new_not_27 = ~Q_0;
  assign new_and_28 = new_not_27 & Q_1;
  assign new_not_29 = ~Q_1;
  assign new_and_30 = Q_0 & new_not_29;
  assign n61554 = new_and_28 | new_and_30;
  assign n61551 = ~Q_0;
  assign new_not_Q_0 = ~Q_0;
  assign new_not_Q_1 = ~Q_1;
  assign new_not_Q_2 = ~Q_2;
  assign new_not_Q_3 = ~Q_3;
  assign new_not_Q_4 = ~Q_4;
  assign new_count_state_1 = Q_0 & new_not_Q_1 & new_not_Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_2 = new_not_Q_0 & Q_1 & new_not_Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_3 = Q_0 & Q_1 & new_not_Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_4 = new_not_Q_0 & new_not_Q_1 & Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_5 = Q_0 & new_not_Q_1 & Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_6 = new_not_Q_0 & Q_1 & Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_7 = Q_0 & Q_1 & Q_2 & new_not_Q_4 & new_not_Q_3;
  assign new_count_state_8 = new_not_Q_0 & new_not_Q_1 & new_not_Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_9 = Q_0 & new_not_Q_1 & new_not_Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_10 = new_not_Q_0 & Q_1 & new_not_Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_11 = Q_0 & Q_1 & new_not_Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_12 = new_not_Q_0 & new_not_Q_1 & Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_13 = Q_0 & new_not_Q_1 & Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_14 = new_not_Q_0 & Q_1 & Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_15 = Q_0 & Q_1 & Q_2 & new_not_Q_4 & Q_3;
  assign new_count_state_16 = new_not_Q_0 & new_not_Q_1 & new_not_Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_17 = Q_0 & new_not_Q_1 & new_not_Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_18 = new_not_Q_0 & Q_1 & new_not_Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_19 = Q_0 & Q_1 & new_not_Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_20 = new_not_Q_0 & new_not_Q_1 & Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_21 = Q_0 & new_not_Q_1 & Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_22 = new_not_Q_0 & Q_1 & Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_23 = Q_0 & Q_1 & Q_2 & Q_4 & new_not_Q_3;
  assign new_count_state_24 = new_not_Q_0 & new_not_Q_1 & new_not_Q_2 & Q_4 & Q_3;
  assign new_count_state_25 = Q_0 & new_not_Q_1 & new_not_Q_2 & Q_4 & Q_3;
  assign new_count_state_26 = new_not_Q_0 & Q_1 & new_not_Q_2 & Q_4 & Q_3;
  assign new_count_state_27 = Q_0 & Q_1 & new_not_Q_2 & Q_4 & Q_3;
  assign new_count_state_28 = new_not_Q_0 & new_not_Q_1 & Q_2 & Q_4 & Q_3;
  assign new_count_state_29 = Q_0 & new_not_Q_1 & Q_2 & Q_4 & Q_3;
  assign new_count_state_30 = new_not_Q_0 & Q_1 & Q_2 & Q_4 & Q_3;
  assign new_count_state_31 = Q_0 & Q_1 & Q_2 & Q_4 & Q_3;
  assign new_y_mux_key0_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key0_and_1 = n189 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key0_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key0_and_3 = n199 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_5 = n209 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_6 = n214 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_7 = n219 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_8 = n224 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_9 = n229 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_10 = n234 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_11 = n239 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_12 = n244 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key0_and_14 = n254 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0 = new_y_mux_key0_and_15 | new_y_mux_key0_and_14 | new_y_mux_key0_and_13 | new_y_mux_key0_and_12 | new_y_mux_key0_and_11 | new_y_mux_key0_and_10 | new_y_mux_key0_and_9 | new_y_mux_key0_and_8 | new_y_mux_key0_and_7 | new_y_mux_key0_and_6 | new_y_mux_key0_and_5 | new_y_mux_key0_and_4 | new_y_mux_key0_and_3 | new_y_mux_key0_and_2 | new_y_mux_key0_and_0 | new_y_mux_key0_and_1;
  assign new_y_mux_key1_and_0 = n184 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key1_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_2 = n194 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key1_and_3 = n199 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_4 = n204 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_5 = n209 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key1_and_6 = n214 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key1_and_7 = n219 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key1_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key1_and_10 = n234 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key1_and_11 = n239 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_12 = n244 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_14 = n254 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key1 = new_y_mux_key1_and_15 | new_y_mux_key1_and_14 | new_y_mux_key1_and_13 | new_y_mux_key1_and_12 | new_y_mux_key1_and_11 | new_y_mux_key1_and_10 | new_y_mux_key1_and_9 | new_y_mux_key1_and_8 | new_y_mux_key1_and_7 | new_y_mux_key1_and_6 | new_y_mux_key1_and_5 | new_y_mux_key1_and_4 | new_y_mux_key1_and_3 | new_y_mux_key1_and_2 | new_y_mux_key1_and_0 | new_y_mux_key1_and_1;
  assign new_y_mux_key2_and_0 = n184 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key2_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key2_and_3 = n199 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_4 = n204 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_5 = n209 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key2_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_7 = n219 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_9 = n229 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_10 = n234 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key2_and_13 = n249 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_14 = n254 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key2_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key2 = new_y_mux_key2_and_15 | new_y_mux_key2_and_14 | new_y_mux_key2_and_13 | new_y_mux_key2_and_12 | new_y_mux_key2_and_11 | new_y_mux_key2_and_10 | new_y_mux_key2_and_9 | new_y_mux_key2_and_8 | new_y_mux_key2_and_7 | new_y_mux_key2_and_6 | new_y_mux_key2_and_5 | new_y_mux_key2_and_4 | new_y_mux_key2_and_3 | new_y_mux_key2_and_2 | new_y_mux_key2_and_0 | new_y_mux_key2_and_1;
  assign new_y_mux_key3_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key3_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key3_and_3 = n199 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_4 = n204 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key3_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_6 = n214 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_7 = n219 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key3_and_8 = n224 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_9 = n229 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key3_and_10 = n234 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_11 = n239 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_12 = n244 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_13 = n249 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key3_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key3 = new_y_mux_key3_and_15 | new_y_mux_key3_and_14 | new_y_mux_key3_and_13 | new_y_mux_key3_and_12 | new_y_mux_key3_and_11 | new_y_mux_key3_and_10 | new_y_mux_key3_and_9 | new_y_mux_key3_and_8 | new_y_mux_key3_and_7 | new_y_mux_key3_and_6 | new_y_mux_key3_and_5 | new_y_mux_key3_and_4 | new_y_mux_key3_and_3 | new_y_mux_key3_and_2 | new_y_mux_key3_and_0 | new_y_mux_key3_and_1;
  assign new_y_mux_key4_and_0 = n184 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key4_and_1 = n189 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_3 = n199 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_4 = n204 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_5 = n209 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_8 = n224 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_10 = n234 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_11 = n239 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key4_and_12 = n244 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key4_and_13 = n249 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key4_and_14 = n254 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4 = new_y_mux_key4_and_15 | new_y_mux_key4_and_14 | new_y_mux_key4_and_13 | new_y_mux_key4_and_12 | new_y_mux_key4_and_11 | new_y_mux_key4_and_10 | new_y_mux_key4_and_9 | new_y_mux_key4_and_8 | new_y_mux_key4_and_7 | new_y_mux_key4_and_6 | new_y_mux_key4_and_5 | new_y_mux_key4_and_4 | new_y_mux_key4_and_3 | new_y_mux_key4_and_2 | new_y_mux_key4_and_0 | new_y_mux_key4_and_1;
  assign new_y_mux_key5_and_0 = n184 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_1 = n189 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_2 = n194 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_3 = n199 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_4 = n204 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_5 = n209 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_6 = n214 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key5_and_7 = n219 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_8 = n224 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_11 = n239 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_12 = n244 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_13 = n249 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_14 = n254 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5 = new_y_mux_key5_and_15 | new_y_mux_key5_and_14 | new_y_mux_key5_and_13 | new_y_mux_key5_and_12 | new_y_mux_key5_and_11 | new_y_mux_key5_and_10 | new_y_mux_key5_and_9 | new_y_mux_key5_and_8 | new_y_mux_key5_and_7 | new_y_mux_key5_and_6 | new_y_mux_key5_and_5 | new_y_mux_key5_and_4 | new_y_mux_key5_and_3 | new_y_mux_key5_and_2 | new_y_mux_key5_and_0 | new_y_mux_key5_and_1;
  assign new_y_mux_key6_and_0 = n184 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key6_and_1 = n189 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key6_and_2 = n194 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_3 = n199 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6_and_4 = n204 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_6 = n214 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_7 = n219 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_8 = n224 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6_and_9 = n229 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_10 = n234 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6_and_12 = n244 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key6_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key6_and_14 = n254 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key6 = new_y_mux_key6_and_15 | new_y_mux_key6_and_14 | new_y_mux_key6_and_13 | new_y_mux_key6_and_12 | new_y_mux_key6_and_11 | new_y_mux_key6_and_10 | new_y_mux_key6_and_9 | new_y_mux_key6_and_8 | new_y_mux_key6_and_7 | new_y_mux_key6_and_6 | new_y_mux_key6_and_5 | new_y_mux_key6_and_4 | new_y_mux_key6_and_3 | new_y_mux_key6_and_2 | new_y_mux_key6_and_0 | new_y_mux_key6_and_1;
  assign new_y_mux_key7_and_0 = n184 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_1 = n189 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_2 = n194 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_3 = n199 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key7_and_4 = n204 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_5 = n209 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_6 = n214 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_7 = n219 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_8 = n224 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_10 = n234 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key7_and_11 = n239 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_12 = n244 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_13 = n249 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_14 = n254 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7 = new_y_mux_key7_and_15 | new_y_mux_key7_and_14 | new_y_mux_key7_and_13 | new_y_mux_key7_and_12 | new_y_mux_key7_and_11 | new_y_mux_key7_and_10 | new_y_mux_key7_and_9 | new_y_mux_key7_and_8 | new_y_mux_key7_and_7 | new_y_mux_key7_and_6 | new_y_mux_key7_and_5 | new_y_mux_key7_and_4 | new_y_mux_key7_and_3 | new_y_mux_key7_and_2 | new_y_mux_key7_and_0 | new_y_mux_key7_and_1;
  assign new_y_mux_key8_and_0 = n184 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_1 = n189 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key8_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_3 = n199 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8_and_4 = n204 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key8_and_5 = n209 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_6 = n214 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_7 = n219 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key8_and_10 = n234 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key8_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8_and_14 = n254 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key8 = new_y_mux_key8_and_15 | new_y_mux_key8_and_14 | new_y_mux_key8_and_13 | new_y_mux_key8_and_12 | new_y_mux_key8_and_11 | new_y_mux_key8_and_10 | new_y_mux_key8_and_9 | new_y_mux_key8_and_8 | new_y_mux_key8_and_7 | new_y_mux_key8_and_6 | new_y_mux_key8_and_5 | new_y_mux_key8_and_4 | new_y_mux_key8_and_3 | new_y_mux_key8_and_2 | new_y_mux_key8_and_0 | new_y_mux_key8_and_1;
  assign new_y_mux_key9_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key9_and_1 = n189 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9_and_3 = n199 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9_and_4 = n204 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key9_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key9_and_9 = n229 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_12 = n244 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9_and_14 = n254 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9 = new_y_mux_key9_and_15 | new_y_mux_key9_and_14 | new_y_mux_key9_and_13 | new_y_mux_key9_and_12 | new_y_mux_key9_and_11 | new_y_mux_key9_and_10 | new_y_mux_key9_and_9 | new_y_mux_key9_and_8 | new_y_mux_key9_and_7 | new_y_mux_key9_and_6 | new_y_mux_key9_and_5 | new_y_mux_key9_and_4 | new_y_mux_key9_and_3 | new_y_mux_key9_and_2 | new_y_mux_key9_and_0 | new_y_mux_key9_and_1;
  assign new_y_mux_key10_and_0 = n184 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key10_and_1 = n189 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key10_and_3 = n199 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_4 = n204 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10_and_5 = n209 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_6 = n214 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key10_and_8 = n224 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10_and_10 = n234 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key10_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_12 = n244 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10_and_13 = n249 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key10_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_15 = new_P1_U3355 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10 = new_y_mux_key10_and_15 | new_y_mux_key10_and_14 | new_y_mux_key10_and_13 | new_y_mux_key10_and_12 | new_y_mux_key10_and_11 | new_y_mux_key10_and_10 | new_y_mux_key10_and_9 | new_y_mux_key10_and_8 | new_y_mux_key10_and_7 | new_y_mux_key10_and_6 | new_y_mux_key10_and_5 | new_y_mux_key10_and_4 | new_y_mux_key10_and_3 | new_y_mux_key10_and_2 | new_y_mux_key10_and_0 | new_y_mux_key10_and_1;
  assign new_y_mux_key11_and_0 = n184 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key11_and_3 = n199 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11_and_4 = n204 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key11_and_5 = n209 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key11_and_8 = n224 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_10 = n234 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11_and_11 = n239 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key11_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_13 = n249 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key11_and_14 = n254 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key11_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11 = new_y_mux_key11_and_15 | new_y_mux_key11_and_14 | new_y_mux_key11_and_13 | new_y_mux_key11_and_12 | new_y_mux_key11_and_11 | new_y_mux_key11_and_10 | new_y_mux_key11_and_9 | new_y_mux_key11_and_8 | new_y_mux_key11_and_7 | new_y_mux_key11_and_6 | new_y_mux_key11_and_5 | new_y_mux_key11_and_4 | new_y_mux_key11_and_3 | new_y_mux_key11_and_2 | new_y_mux_key11_and_0 | new_y_mux_key11_and_1;
  assign new_y_mux_key12_and_0 = n184 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12_and_1 = n189 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12_and_3 = n199 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_4 = n204 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_5 = n209 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key12_and_6 = n214 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_8 = n224 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12_and_9 = n229 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key12_and_12 = n244 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_13 = n249 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_15 = new_P1_U3355 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key12 = new_y_mux_key12_and_15 | new_y_mux_key12_and_14 | new_y_mux_key12_and_13 | new_y_mux_key12_and_12 | new_y_mux_key12_and_11 | new_y_mux_key12_and_10 | new_y_mux_key12_and_9 | new_y_mux_key12_and_8 | new_y_mux_key12_and_7 | new_y_mux_key12_and_6 | new_y_mux_key12_and_5 | new_y_mux_key12_and_4 | new_y_mux_key12_and_3 | new_y_mux_key12_and_2 | new_y_mux_key12_and_0 | new_y_mux_key12_and_1;
  assign new_y_mux_key13_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_1 = n189 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_2 = n194 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_3 = n199 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_4 = n204 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key13_and_5 = n209 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key13_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_8 = n224 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_9 = n229 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key13_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key13_and_11 = n239 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_12 = n244 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key13_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key13 = new_y_mux_key13_and_15 | new_y_mux_key13_and_14 | new_y_mux_key13_and_13 | new_y_mux_key13_and_12 | new_y_mux_key13_and_11 | new_y_mux_key13_and_10 | new_y_mux_key13_and_9 | new_y_mux_key13_and_8 | new_y_mux_key13_and_7 | new_y_mux_key13_and_6 | new_y_mux_key13_and_5 | new_y_mux_key13_and_4 | new_y_mux_key13_and_3 | new_y_mux_key13_and_2 | new_y_mux_key13_and_0 | new_y_mux_key13_and_1;
  assign new_y_mux_key14_and_0 = n184 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_1 = n189 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_2 = n194 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_3 = n199 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_4 = n204 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key14_and_5 = n209 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key14_and_6 = n214 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key14_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_8 = n224 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key14_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key14_and_12 = n244 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key14_and_13 = n249 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key14_and_14 = n254 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key14_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14 = new_y_mux_key14_and_15 | new_y_mux_key14_and_14 | new_y_mux_key14_and_13 | new_y_mux_key14_and_12 | new_y_mux_key14_and_11 | new_y_mux_key14_and_10 | new_y_mux_key14_and_9 | new_y_mux_key14_and_8 | new_y_mux_key14_and_7 | new_y_mux_key14_and_6 | new_y_mux_key14_and_5 | new_y_mux_key14_and_4 | new_y_mux_key14_and_3 | new_y_mux_key14_and_2 | new_y_mux_key14_and_0 | new_y_mux_key14_and_1;
  assign new_y_mux_key15_and_0 = n184 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_1 = n189 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_3 = n199 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key15_and_4 = n204 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_5 = n209 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_6 = n214 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_9 = n229 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key15_and_10 = n234 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key15_and_11 = n239 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key15_and_13 = n249 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_14 = n254 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key15_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key15 = new_y_mux_key15_and_15 | new_y_mux_key15_and_14 | new_y_mux_key15_and_13 | new_y_mux_key15_and_12 | new_y_mux_key15_and_11 | new_y_mux_key15_and_10 | new_y_mux_key15_and_9 | new_y_mux_key15_and_8 | new_y_mux_key15_and_7 | new_y_mux_key15_and_6 | new_y_mux_key15_and_5 | new_y_mux_key15_and_4 | new_y_mux_key15_and_3 | new_y_mux_key15_and_2 | new_y_mux_key15_and_0 | new_y_mux_key15_and_1;
  assign new_y_mux_key16_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_1 = n189 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key16_and_2 = n194 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key16_and_3 = n199 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_4 = n204 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key16_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key16_and_6 = n214 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_8 = n224 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_9 = n229 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key16_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_13 = n249 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key16_and_14 = n254 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key16 = new_y_mux_key16_and_15 | new_y_mux_key16_and_14 | new_y_mux_key16_and_13 | new_y_mux_key16_and_12 | new_y_mux_key16_and_11 | new_y_mux_key16_and_10 | new_y_mux_key16_and_9 | new_y_mux_key16_and_8 | new_y_mux_key16_and_7 | new_y_mux_key16_and_6 | new_y_mux_key16_and_5 | new_y_mux_key16_and_4 | new_y_mux_key16_and_3 | new_y_mux_key16_and_2 | new_y_mux_key16_and_0 | new_y_mux_key16_and_1;
  assign new_y_mux_key17_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key17_and_1 = n189 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_2 = n194 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key17_and_3 = n199 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key17_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key17_and_5 = n209 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_6 = n214 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key17_and_7 = n219 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key17_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_10 = n234 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key17_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key17_and_13 = n249 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_14 = n254 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key17_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key17 = new_y_mux_key17_and_15 | new_y_mux_key17_and_14 | new_y_mux_key17_and_13 | new_y_mux_key17_and_12 | new_y_mux_key17_and_11 | new_y_mux_key17_and_10 | new_y_mux_key17_and_9 | new_y_mux_key17_and_8 | new_y_mux_key17_and_7 | new_y_mux_key17_and_6 | new_y_mux_key17_and_5 | new_y_mux_key17_and_4 | new_y_mux_key17_and_3 | new_y_mux_key17_and_2 | new_y_mux_key17_and_0 | new_y_mux_key17_and_1;
  assign new_y_mux_key18_and_0 = n184 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key18_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key18_and_3 = n199 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key18_and_5 = n209 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key18_and_6 = n214 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_7 = n219 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key18_and_10 = n234 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key18_and_12 = n244 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key18_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key18_and_14 = n254 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key18_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key18 = new_y_mux_key18_and_15 | new_y_mux_key18_and_14 | new_y_mux_key18_and_13 | new_y_mux_key18_and_12 | new_y_mux_key18_and_11 | new_y_mux_key18_and_10 | new_y_mux_key18_and_9 | new_y_mux_key18_and_8 | new_y_mux_key18_and_7 | new_y_mux_key18_and_6 | new_y_mux_key18_and_5 | new_y_mux_key18_and_4 | new_y_mux_key18_and_3 | new_y_mux_key18_and_2 | new_y_mux_key18_and_0 | new_y_mux_key18_and_1;
  assign new_y_mux_key19_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_2 = n194 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_3 = n199 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key19_and_4 = n204 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_5 = n209 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key19_and_6 = n214 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key19_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_8 = n224 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key19_and_9 = n229 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_11 = n239 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key19_and_12 = n244 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_13 = n249 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_14 = n254 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key19_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key19 = new_y_mux_key19_and_15 | new_y_mux_key19_and_14 | new_y_mux_key19_and_13 | new_y_mux_key19_and_12 | new_y_mux_key19_and_11 | new_y_mux_key19_and_10 | new_y_mux_key19_and_9 | new_y_mux_key19_and_8 | new_y_mux_key19_and_7 | new_y_mux_key19_and_6 | new_y_mux_key19_and_5 | new_y_mux_key19_and_4 | new_y_mux_key19_and_3 | new_y_mux_key19_and_2 | new_y_mux_key19_and_0 | new_y_mux_key19_and_1;
  assign new_y_mux_key20_and_0 = n184 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_1 = n189 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_2 = n194 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_3 = n199 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_4 = n204 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key20_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_7 = n219 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key20_and_8 = n224 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key20_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_12 = n244 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key20_and_13 = n249 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_14 = n254 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20_and_15 = new_P1_U3355 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key20 = new_y_mux_key20_and_15 | new_y_mux_key20_and_14 | new_y_mux_key20_and_13 | new_y_mux_key20_and_12 | new_y_mux_key20_and_11 | new_y_mux_key20_and_10 | new_y_mux_key20_and_9 | new_y_mux_key20_and_8 | new_y_mux_key20_and_7 | new_y_mux_key20_and_6 | new_y_mux_key20_and_5 | new_y_mux_key20_and_4 | new_y_mux_key20_and_3 | new_y_mux_key20_and_2 | new_y_mux_key20_and_0 | new_y_mux_key20_and_1;
  assign new_y_mux_key21_and_0 = n184 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key21_and_1 = n189 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key21_and_2 = n194 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key21_and_3 = n199 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_4 = n204 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key21_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key21_and_7 = n219 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_8 = n224 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_9 = n229 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key21_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_13 = n249 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key21_and_14 = n254 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key21_and_15 = new_P1_U3355 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key21 = new_y_mux_key21_and_15 | new_y_mux_key21_and_14 | new_y_mux_key21_and_13 | new_y_mux_key21_and_12 | new_y_mux_key21_and_11 | new_y_mux_key21_and_10 | new_y_mux_key21_and_9 | new_y_mux_key21_and_8 | new_y_mux_key21_and_7 | new_y_mux_key21_and_6 | new_y_mux_key21_and_5 | new_y_mux_key21_and_4 | new_y_mux_key21_and_3 | new_y_mux_key21_and_2 | new_y_mux_key21_and_0 | new_y_mux_key21_and_1;
  assign new_y_mux_key22_and_0 = n184 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_1 = n189 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key22_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key22_and_3 = n199 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key22_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key22_and_5 = n209 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key22_and_6 = n214 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key22_and_7 = n219 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key22_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key22_and_10 = n234 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_11 = n239 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_12 = n244 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_13 = n249 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_14 = n254 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22_and_15 = new_P1_U3355 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key22 = new_y_mux_key22_and_15 | new_y_mux_key22_and_14 | new_y_mux_key22_and_13 | new_y_mux_key22_and_12 | new_y_mux_key22_and_11 | new_y_mux_key22_and_10 | new_y_mux_key22_and_9 | new_y_mux_key22_and_8 | new_y_mux_key22_and_7 | new_y_mux_key22_and_6 | new_y_mux_key22_and_5 | new_y_mux_key22_and_4 | new_y_mux_key22_and_3 | new_y_mux_key22_and_2 | new_y_mux_key22_and_0 | new_y_mux_key22_and_1;
  assign new_y_mux_key23_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key23_and_1 = n189 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key23_and_2 = n194 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key23_and_3 = n199 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key23_and_7 = n219 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_8 = n224 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key23_and_10 = n234 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_11 = n239 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23_and_12 = n244 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key23_and_13 = n249 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key23_and_14 = n254 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key23_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key23 = new_y_mux_key23_and_15 | new_y_mux_key23_and_14 | new_y_mux_key23_and_13 | new_y_mux_key23_and_12 | new_y_mux_key23_and_11 | new_y_mux_key23_and_10 | new_y_mux_key23_and_9 | new_y_mux_key23_and_8 | new_y_mux_key23_and_7 | new_y_mux_key23_and_6 | new_y_mux_key23_and_5 | new_y_mux_key23_and_4 | new_y_mux_key23_and_3 | new_y_mux_key23_and_2 | new_y_mux_key23_and_0 | new_y_mux_key23_and_1;
  assign new_y_mux_key24_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_1 = n189 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_2 = n194 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_3 = n199 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_4 = n204 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_5 = n209 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key24_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_8 = n224 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key24_and_9 = n229 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_10 = n234 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key24_and_11 = n239 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_12 = n244 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key24_and_13 = n249 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_14 = n254 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key24 = new_y_mux_key24_and_15 | new_y_mux_key24_and_14 | new_y_mux_key24_and_13 | new_y_mux_key24_and_12 | new_y_mux_key24_and_11 | new_y_mux_key24_and_10 | new_y_mux_key24_and_9 | new_y_mux_key24_and_8 | new_y_mux_key24_and_7 | new_y_mux_key24_and_6 | new_y_mux_key24_and_5 | new_y_mux_key24_and_4 | new_y_mux_key24_and_3 | new_y_mux_key24_and_2 | new_y_mux_key24_and_0 | new_y_mux_key24_and_1;
  assign new_y_mux_key25_and_0 = n184 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key25_and_1 = n189 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key25_and_2 = n194 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key25_and_3 = n199 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key25_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key25_and_5 = n209 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key25_and_6 = n214 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key25_and_7 = n219 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key25_and_8 = n224 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key25_and_9 = n229 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key25_and_10 = n234 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key25_and_11 = n239 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key25_and_12 = n244 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key25_and_13 = n249 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key25_and_14 = n254 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key25_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key25 = new_y_mux_key25_and_15 | new_y_mux_key25_and_14 | new_y_mux_key25_and_13 | new_y_mux_key25_and_12 | new_y_mux_key25_and_11 | new_y_mux_key25_and_10 | new_y_mux_key25_and_9 | new_y_mux_key25_and_8 | new_y_mux_key25_and_7 | new_y_mux_key25_and_6 | new_y_mux_key25_and_5 | new_y_mux_key25_and_4 | new_y_mux_key25_and_3 | new_y_mux_key25_and_2 | new_y_mux_key25_and_0 | new_y_mux_key25_and_1;
  assign new_y_mux_key26_and_0 = n184 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key26_and_1 = n189 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_3 = n199 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_4 = n204 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_5 = n209 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_6 = n214 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key26_and_7 = n219 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_9 = n229 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key26_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key26_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_12 = n244 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key26_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_14 = n254 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key26_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key26 = new_y_mux_key26_and_15 | new_y_mux_key26_and_14 | new_y_mux_key26_and_13 | new_y_mux_key26_and_12 | new_y_mux_key26_and_11 | new_y_mux_key26_and_10 | new_y_mux_key26_and_9 | new_y_mux_key26_and_8 | new_y_mux_key26_and_7 | new_y_mux_key26_and_6 | new_y_mux_key26_and_5 | new_y_mux_key26_and_4 | new_y_mux_key26_and_3 | new_y_mux_key26_and_2 | new_y_mux_key26_and_0 | new_y_mux_key26_and_1;
  assign new_y_mux_key27_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key27_and_1 = n189 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27_and_2 = n194 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key27_and_3 = n199 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key27_and_4 = n204 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key27_and_5 = n209 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key27_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key27_and_8 = n224 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27_and_9 = n229 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key27_and_10 = n234 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key27_and_13 = n249 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key27_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key27 = new_y_mux_key27_and_15 | new_y_mux_key27_and_14 | new_y_mux_key27_and_13 | new_y_mux_key27_and_12 | new_y_mux_key27_and_11 | new_y_mux_key27_and_10 | new_y_mux_key27_and_9 | new_y_mux_key27_and_8 | new_y_mux_key27_and_7 | new_y_mux_key27_and_6 | new_y_mux_key27_and_5 | new_y_mux_key27_and_4 | new_y_mux_key27_and_3 | new_y_mux_key27_and_2 | new_y_mux_key27_and_0 | new_y_mux_key27_and_1;
  assign new_y_mux_key28_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_1 = n189 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_2 = n194 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_3 = n199 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key28_and_4 = n204 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_5 = n209 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key28_and_6 = n214 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key28_and_7 = n219 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_8 = n224 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key28_and_9 = n229 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key28_and_10 = n234 & keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_11 = n239 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_12 = n244 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key28_and_13 = n249 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key28_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28_and_15 = new_P1_U3355 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key28 = new_y_mux_key28_and_15 | new_y_mux_key28_and_14 | new_y_mux_key28_and_13 | new_y_mux_key28_and_12 | new_y_mux_key28_and_11 | new_y_mux_key28_and_10 | new_y_mux_key28_and_9 | new_y_mux_key28_and_8 | new_y_mux_key28_and_7 | new_y_mux_key28_and_6 | new_y_mux_key28_and_5 | new_y_mux_key28_and_4 | new_y_mux_key28_and_3 | new_y_mux_key28_and_2 | new_y_mux_key28_and_0 | new_y_mux_key28_and_1;
  assign new_y_mux_key29_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_1 = n189 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_2 = n194 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_3 = n199 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_4 = n204 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key29_and_5 = n209 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key29_and_6 = n214 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key29_and_8 = n224 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key29_and_9 = n229 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key29_and_11 = n239 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key29_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key29_and_13 = n249 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key29_and_14 = n254 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key29_and_15 = new_P1_U3355 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key29 = new_y_mux_key29_and_15 | new_y_mux_key29_and_14 | new_y_mux_key29_and_13 | new_y_mux_key29_and_12 | new_y_mux_key29_and_11 | new_y_mux_key29_and_10 | new_y_mux_key29_and_9 | new_y_mux_key29_and_8 | new_y_mux_key29_and_7 | new_y_mux_key29_and_6 | new_y_mux_key29_and_5 | new_y_mux_key29_and_4 | new_y_mux_key29_and_3 | new_y_mux_key29_and_2 | new_y_mux_key29_and_0 | new_y_mux_key29_and_1;
  assign new_y_mux_key30_and_0 = n184 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30_and_1 = n189 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_2 = n194 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30_and_3 = n199 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30_and_4 = n204 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_5 = n209 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key30_and_6 = n214 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30_and_7 = n219 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30_and_8 = n224 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_9 = n229 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_10 = n234 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_12 = n244 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_13 = n249 & new_not_keyinput31 & keyinput30 & keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key30_and_14 = n254 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & new_not_keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30_and_15 = new_P1_U3355 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key30 = new_y_mux_key30_and_15 | new_y_mux_key30_and_14 | new_y_mux_key30_and_13 | new_y_mux_key30_and_12 | new_y_mux_key30_and_11 | new_y_mux_key30_and_10 | new_y_mux_key30_and_9 | new_y_mux_key30_and_8 | new_y_mux_key30_and_7 | new_y_mux_key30_and_6 | new_y_mux_key30_and_5 | new_y_mux_key30_and_4 | new_y_mux_key30_and_3 | new_y_mux_key30_and_2 | new_y_mux_key30_and_0 | new_y_mux_key30_and_1;
  assign new_y_mux_key31_and_0 = n184 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key31_and_1 = n189 & keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & new_not_keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_2 = n194 & keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_3 = n199 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_4 = n204 & new_not_keyinput31 & keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_5 = n209 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & new_not_keyinput23 & keyinput22 & keyinput21 & keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & keyinput15 & keyinput14 & keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_6 = n214 & keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_7 = n219 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_8 = n224 & new_not_keyinput31 & new_not_keyinput30 & keyinput29 & keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & keyinput19 & keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key31_and_9 = n229 & keyinput31 & new_not_keyinput30 & keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & new_not_keyinput25 & new_not_keyinput24 & keyinput23 & keyinput22 & new_not_keyinput21 & keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & new_not_keyinput7 & new_not_keyinput6 & new_not_keyinput5 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_10 = n234 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & keyinput26 & keyinput25 & keyinput24 & new_not_keyinput23 & keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & keyinput8 & new_not_keyinput7 & keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_11 = n239 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & new_not_keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_12 = n244 & keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & new_not_keyinput27 & new_not_keyinput26 & new_not_keyinput25 & new_not_keyinput24 & new_not_keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & new_not_keyinput19 & new_not_keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & new_not_keyinput14 & keyinput13 & new_not_keyinput12 & keyinput11 & new_not_keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & new_not_keyinput5 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_13 = n249 & keyinput31 & keyinput30 & keyinput29 & keyinput28 & new_not_keyinput27 & keyinput26 & keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & new_not_keyinput21 & new_not_keyinput20 & keyinput19 & new_not_keyinput18 & keyinput17 & new_not_keyinput16 & keyinput15 & keyinput14 & new_not_keyinput13 & keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & keyinput6 & keyinput5 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31_and_14 = n254 & new_not_keyinput31 & new_not_keyinput30 & new_not_keyinput29 & new_not_keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & keyinput23 & new_not_keyinput22 & keyinput21 & keyinput20 & keyinput19 & keyinput18 & keyinput17 & keyinput16 & new_not_keyinput15 & keyinput14 & new_not_keyinput13 & new_not_keyinput12 & keyinput11 & keyinput10 & new_not_keyinput9 & new_not_keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key31_and_15 = new_P1_U3355 & new_not_keyinput31 & keyinput30 & new_not_keyinput29 & keyinput28 & keyinput27 & new_not_keyinput26 & new_not_keyinput25 & keyinput24 & new_not_keyinput23 & new_not_keyinput22 & keyinput21 & new_not_keyinput20 & new_not_keyinput19 & keyinput18 & new_not_keyinput17 & keyinput16 & keyinput15 & new_not_keyinput14 & new_not_keyinput13 & keyinput12 & new_not_keyinput11 & keyinput10 & keyinput9 & keyinput8 & keyinput7 & new_not_keyinput6 & keyinput5 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key31 = new_y_mux_key31_and_15 | new_y_mux_key31_and_14 | new_y_mux_key31_and_13 | new_y_mux_key31_and_12 | new_y_mux_key31_and_11 | new_y_mux_key31_and_10 | new_y_mux_key31_and_9 | new_y_mux_key31_and_8 | new_y_mux_key31_and_7 | new_y_mux_key31_and_6 | new_y_mux_key31_and_5 | new_y_mux_key31_and_4 | new_y_mux_key31_and_3 | new_y_mux_key31_and_2 | new_y_mux_key31_and_0 | new_y_mux_key31_and_1;
  assign new__state_1 = new_count_state_1;
  assign new__state_2 = new_count_state_2;
  assign new__state_3 = new_count_state_3;
  assign new__state_4 = new_count_state_4;
  assign new__state_5 = new_count_state_5;
  assign new__state_6 = new_count_state_6;
  assign new__state_7 = new_count_state_7;
  assign new__state_8 = new_count_state_8;
  assign new__state_9 = new_count_state_9;
  assign new__state_10 = new_count_state_10;
  assign new__state_11 = new_count_state_11;
  assign new__state_12 = new_count_state_12;
  assign new__state_13 = new_count_state_13;
  assign new__state_14 = new_count_state_14;
  assign new__state_15 = new_count_state_15;
  assign new__state_16 = new_count_state_16;
  assign new__state_17 = new_count_state_17;
  assign new__state_18 = new_count_state_18;
  assign new__state_19 = new_count_state_19;
  assign new__state_20 = new_count_state_20;
  assign new__state_21 = new_count_state_21;
  assign new__state_22 = new_count_state_22;
  assign new__state_23 = new_count_state_23;
  assign new__state_24 = new_count_state_24;
  assign new__state_25 = new_count_state_25;
  assign new__state_26 = new_count_state_26;
  assign new__state_27 = new_count_state_27;
  assign new__state_28 = new_count_state_28;
  assign new__state_29 = new_count_state_29;
  assign new__state_30 = new_count_state_30;
  assign new__state_31 = new_count_state_31;
  assign new__state_33 = new__state_2 | new__state_3;
  assign new__state_34 = new__state_4 | new__state_5;
  assign new__state_35 = new__state_6 | new__state_7;
  assign new__state_36 = new__state_8 | new__state_9;
  assign new__state_37 = new__state_10 | new__state_11;
  assign new__state_38 = new__state_12 | new__state_13;
  assign new__state_39 = new__state_14 | new__state_15;
  assign new__state_40 = new__state_16 | new__state_17;
  assign new__state_41 = new__state_18 | new__state_19;
  assign new__state_42 = new__state_20 | new__state_21;
  assign new__state_43 = new__state_22 | new__state_23;
  assign new__state_44 = new__state_24 | new__state_25;
  assign new__state_45 = new__state_26 | new__state_27;
  assign new__state_46 = new__state_28 | new__state_29;
  assign new__state_47 = new__state_30 | new__state_31;
  assign new__state_49 = new__state_34 | new__state_35;
  assign new__state_50 = new__state_36 | new__state_37;
  assign new__state_51 = new__state_38 | new__state_39;
  assign new__state_52 = new__state_40 | new__state_41;
  assign new__state_53 = new__state_42 | new__state_43;
  assign new__state_54 = new__state_44 | new__state_45;
  assign new__state_55 = new__state_46 | new__state_47;
  assign new__state_57 = new__state_50 | new__state_51;
  assign new__state_58 = new__state_52 | new__state_53;
  assign new__state_59 = new__state_54 | new__state_55;
  assign new__state_61 = new__state_58 | new__state_59;
  assign new_s__state_1 = new__state_1;
  assign new_not_s__state_1 = ~new_s__state_1;
  assign new_I0__state_1 = new_y_mux_key0;
  assign new_I1__state_1 = new_y_mux_key1;
  assign new_and_mux__state_1 = new_not_s__state_1 & new_I0__state_1;
  assign new_and_mux__state_1_2 = new_s__state_1 & new_I1__state_1;
  assign new_y_mux_32 = new_and_mux__state_1 | new_and_mux__state_1_2;
  assign new_s__state_3 = new__state_3;
  assign new_not_s__state_3 = ~new_s__state_3;
  assign new_I0__state_3 = new_y_mux_key2;
  assign new_I1__state_3 = new_y_mux_key3;
  assign new_and_mux__state_3 = new_not_s__state_3 & new_I0__state_3;
  assign new_and_mux__state_3_2 = new_s__state_3 & new_I1__state_3;
  assign new_y_mux_33 = new_and_mux__state_3 | new_and_mux__state_3_2;
  assign new_s__state_5 = new__state_5;
  assign new_not_s__state_5 = ~new_s__state_5;
  assign new_I0__state_5 = new_y_mux_key4;
  assign new_I1__state_5 = new_y_mux_key5;
  assign new_and_mux__state_5 = new_not_s__state_5 & new_I0__state_5;
  assign new_and_mux__state_5_2 = new_s__state_5 & new_I1__state_5;
  assign new_y_mux_34 = new_and_mux__state_5 | new_and_mux__state_5_2;
  assign new_s__state_7 = new__state_7;
  assign new_not_s__state_7 = ~new_s__state_7;
  assign new_I0__state_7 = new_y_mux_key6;
  assign new_I1__state_7 = new_y_mux_key7;
  assign new_and_mux__state_7 = new_not_s__state_7 & new_I0__state_7;
  assign new_and_mux__state_7_2 = new_s__state_7 & new_I1__state_7;
  assign new_y_mux_35 = new_and_mux__state_7 | new_and_mux__state_7_2;
  assign new_s__state_9 = new__state_9;
  assign new_not_s__state_9 = ~new_s__state_9;
  assign new_I0__state_9 = new_y_mux_key8;
  assign new_I1__state_9 = new_y_mux_key9;
  assign new_and_mux__state_9 = new_not_s__state_9 & new_I0__state_9;
  assign new_and_mux__state_9_2 = new_s__state_9 & new_I1__state_9;
  assign new_y_mux_36 = new_and_mux__state_9 | new_and_mux__state_9_2;
  assign new_s__state_11 = new__state_11;
  assign new_not_s__state_11 = ~new_s__state_11;
  assign new_I0__state_11 = new_y_mux_key10;
  assign new_I1__state_11 = new_y_mux_key11;
  assign new_and_mux__state_11 = new_not_s__state_11 & new_I0__state_11;
  assign new_and_mux__state_11_2 = new_s__state_11 & new_I1__state_11;
  assign new_y_mux_37 = new_and_mux__state_11 | new_and_mux__state_11_2;
  assign new_s__state_13 = new__state_13;
  assign new_not_s__state_13 = ~new_s__state_13;
  assign new_I0__state_13 = new_y_mux_key12;
  assign new_I1__state_13 = new_y_mux_key13;
  assign new_and_mux__state_13 = new_not_s__state_13 & new_I0__state_13;
  assign new_and_mux__state_13_2 = new_s__state_13 & new_I1__state_13;
  assign new_y_mux_38 = new_and_mux__state_13 | new_and_mux__state_13_2;
  assign new_s__state_15 = new__state_15;
  assign new_not_s__state_15 = ~new_s__state_15;
  assign new_I0__state_15 = new_y_mux_key14;
  assign new_I1__state_15 = new_y_mux_key15;
  assign new_and_mux__state_15 = new_not_s__state_15 & new_I0__state_15;
  assign new_and_mux__state_15_2 = new_s__state_15 & new_I1__state_15;
  assign new_y_mux_39 = new_and_mux__state_15 | new_and_mux__state_15_2;
  assign new_s__state_17 = new__state_17;
  assign new_not_s__state_17 = ~new_s__state_17;
  assign new_I0__state_17 = new_y_mux_key16;
  assign new_I1__state_17 = new_y_mux_key17;
  assign new_and_mux__state_17 = new_not_s__state_17 & new_I0__state_17;
  assign new_and_mux__state_17_2 = new_s__state_17 & new_I1__state_17;
  assign new_y_mux_40 = new_and_mux__state_17 | new_and_mux__state_17_2;
  assign new_s__state_19 = new__state_19;
  assign new_not_s__state_19 = ~new_s__state_19;
  assign new_I0__state_19 = new_y_mux_key18;
  assign new_I1__state_19 = new_y_mux_key19;
  assign new_and_mux__state_19 = new_not_s__state_19 & new_I0__state_19;
  assign new_and_mux__state_19_2 = new_s__state_19 & new_I1__state_19;
  assign new_y_mux_41 = new_and_mux__state_19 | new_and_mux__state_19_2;
  assign new_s__state_21 = new__state_21;
  assign new_not_s__state_21 = ~new_s__state_21;
  assign new_I0__state_21 = new_y_mux_key20;
  assign new_I1__state_21 = new_y_mux_key21;
  assign new_and_mux__state_21 = new_not_s__state_21 & new_I0__state_21;
  assign new_and_mux__state_21_2 = new_s__state_21 & new_I1__state_21;
  assign new_y_mux_42 = new_and_mux__state_21 | new_and_mux__state_21_2;
  assign new_s__state_23 = new__state_23;
  assign new_not_s__state_23 = ~new_s__state_23;
  assign new_I0__state_23 = new_y_mux_key22;
  assign new_I1__state_23 = new_y_mux_key23;
  assign new_and_mux__state_23 = new_not_s__state_23 & new_I0__state_23;
  assign new_and_mux__state_23_2 = new_s__state_23 & new_I1__state_23;
  assign new_y_mux_43 = new_and_mux__state_23 | new_and_mux__state_23_2;
  assign new_s__state_25 = new__state_25;
  assign new_not_s__state_25 = ~new_s__state_25;
  assign new_I0__state_25 = new_y_mux_key24;
  assign new_I1__state_25 = new_y_mux_key25;
  assign new_and_mux__state_25 = new_not_s__state_25 & new_I0__state_25;
  assign new_and_mux__state_25_2 = new_s__state_25 & new_I1__state_25;
  assign new_y_mux_44 = new_and_mux__state_25 | new_and_mux__state_25_2;
  assign new_s__state_27 = new__state_27;
  assign new_not_s__state_27 = ~new_s__state_27;
  assign new_I0__state_27 = new_y_mux_key26;
  assign new_I1__state_27 = new_y_mux_key27;
  assign new_and_mux__state_27 = new_not_s__state_27 & new_I0__state_27;
  assign new_and_mux__state_27_2 = new_s__state_27 & new_I1__state_27;
  assign new_y_mux_45 = new_and_mux__state_27 | new_and_mux__state_27_2;
  assign new_s__state_29 = new__state_29;
  assign new_not_s__state_29 = ~new_s__state_29;
  assign new_I0__state_29 = new_y_mux_key28;
  assign new_I1__state_29 = new_y_mux_key29;
  assign new_and_mux__state_29 = new_not_s__state_29 & new_I0__state_29;
  assign new_and_mux__state_29_2 = new_s__state_29 & new_I1__state_29;
  assign new_y_mux_46 = new_and_mux__state_29 | new_and_mux__state_29_2;
  assign new_s__state_31 = new__state_31;
  assign new_not_s__state_31 = ~new_s__state_31;
  assign new_I0__state_31 = new_y_mux_key30;
  assign new_I1__state_31 = new_y_mux_key31;
  assign new_and_mux__state_31 = new_not_s__state_31 & new_I0__state_31;
  assign new_and_mux__state_31_2 = new_s__state_31 & new_I1__state_31;
  assign new_y_mux_47 = new_and_mux__state_31 | new_and_mux__state_31_2;
  assign new_s__state_33 = new__state_33;
  assign new_not_s__state_33 = ~new_s__state_33;
  assign new_I0__state_33 = new_y_mux_32;
  assign new_I1__state_33 = new_y_mux_33;
  assign new_and_mux__state_33 = new_not_s__state_33 & new_I0__state_33;
  assign new_and_mux__state_33_2 = new_s__state_33 & new_I1__state_33;
  assign new_y_mux_48 = new_and_mux__state_33 | new_and_mux__state_33_2;
  assign new_s__state_35 = new__state_35;
  assign new_not_s__state_35 = ~new_s__state_35;
  assign new_I0__state_35 = new_y_mux_34;
  assign new_I1__state_35 = new_y_mux_35;
  assign new_and_mux__state_35 = new_not_s__state_35 & new_I0__state_35;
  assign new_and_mux__state_35_2 = new_s__state_35 & new_I1__state_35;
  assign new_y_mux_49 = new_and_mux__state_35 | new_and_mux__state_35_2;
  assign new_s__state_37 = new__state_37;
  assign new_not_s__state_37 = ~new_s__state_37;
  assign new_I0__state_37 = new_y_mux_36;
  assign new_I1__state_37 = new_y_mux_37;
  assign new_and_mux__state_37 = new_not_s__state_37 & new_I0__state_37;
  assign new_and_mux__state_37_2 = new_s__state_37 & new_I1__state_37;
  assign new_y_mux_50 = new_and_mux__state_37 | new_and_mux__state_37_2;
  assign new_s__state_39 = new__state_39;
  assign new_not_s__state_39 = ~new_s__state_39;
  assign new_I0__state_39 = new_y_mux_38;
  assign new_I1__state_39 = new_y_mux_39;
  assign new_and_mux__state_39 = new_not_s__state_39 & new_I0__state_39;
  assign new_and_mux__state_39_2 = new_s__state_39 & new_I1__state_39;
  assign new_y_mux_51 = new_and_mux__state_39 | new_and_mux__state_39_2;
  assign new_s__state_41 = new__state_41;
  assign new_not_s__state_41 = ~new_s__state_41;
  assign new_I0__state_41 = new_y_mux_40;
  assign new_I1__state_41 = new_y_mux_41;
  assign new_and_mux__state_41 = new_not_s__state_41 & new_I0__state_41;
  assign new_and_mux__state_41_2 = new_s__state_41 & new_I1__state_41;
  assign new_y_mux_52 = new_and_mux__state_41 | new_and_mux__state_41_2;
  assign new_s__state_43 = new__state_43;
  assign new_not_s__state_43 = ~new_s__state_43;
  assign new_I0__state_43 = new_y_mux_42;
  assign new_I1__state_43 = new_y_mux_43;
  assign new_and_mux__state_43 = new_not_s__state_43 & new_I0__state_43;
  assign new_and_mux__state_43_2 = new_s__state_43 & new_I1__state_43;
  assign new_y_mux_53 = new_and_mux__state_43 | new_and_mux__state_43_2;
  assign new_s__state_45 = new__state_45;
  assign new_not_s__state_45 = ~new_s__state_45;
  assign new_I0__state_45 = new_y_mux_44;
  assign new_I1__state_45 = new_y_mux_45;
  assign new_and_mux__state_45 = new_not_s__state_45 & new_I0__state_45;
  assign new_and_mux__state_45_2 = new_s__state_45 & new_I1__state_45;
  assign new_y_mux_54 = new_and_mux__state_45 | new_and_mux__state_45_2;
  assign new_s__state_47 = new__state_47;
  assign new_not_s__state_47 = ~new_s__state_47;
  assign new_I0__state_47 = new_y_mux_46;
  assign new_I1__state_47 = new_y_mux_47;
  assign new_and_mux__state_47 = new_not_s__state_47 & new_I0__state_47;
  assign new_and_mux__state_47_2 = new_s__state_47 & new_I1__state_47;
  assign new_y_mux_55 = new_and_mux__state_47 | new_and_mux__state_47_2;
  assign new_s__state_49 = new__state_49;
  assign new_not_s__state_49 = ~new_s__state_49;
  assign new_I0__state_49 = new_y_mux_48;
  assign new_I1__state_49 = new_y_mux_49;
  assign new_and_mux__state_49 = new_not_s__state_49 & new_I0__state_49;
  assign new_and_mux__state_49_2 = new_s__state_49 & new_I1__state_49;
  assign new_y_mux_56 = new_and_mux__state_49 | new_and_mux__state_49_2;
  assign new_s__state_51 = new__state_51;
  assign new_not_s__state_51 = ~new_s__state_51;
  assign new_I0__state_51 = new_y_mux_50;
  assign new_I1__state_51 = new_y_mux_51;
  assign new_and_mux__state_51 = new_not_s__state_51 & new_I0__state_51;
  assign new_and_mux__state_51_2 = new_s__state_51 & new_I1__state_51;
  assign new_y_mux_57 = new_and_mux__state_51 | new_and_mux__state_51_2;
  assign new_s__state_53 = new__state_53;
  assign new_not_s__state_53 = ~new_s__state_53;
  assign new_I0__state_53 = new_y_mux_52;
  assign new_I1__state_53 = new_y_mux_53;
  assign new_and_mux__state_53 = new_not_s__state_53 & new_I0__state_53;
  assign new_and_mux__state_53_2 = new_s__state_53 & new_I1__state_53;
  assign new_y_mux_58 = new_and_mux__state_53 | new_and_mux__state_53_2;
  assign new_s__state_55 = new__state_55;
  assign new_not_s__state_55 = ~new_s__state_55;
  assign new_I0__state_55 = new_y_mux_54;
  assign new_I1__state_55 = new_y_mux_55;
  assign new_and_mux__state_55 = new_not_s__state_55 & new_I0__state_55;
  assign new_and_mux__state_55_2 = new_s__state_55 & new_I1__state_55;
  assign new_y_mux_59 = new_and_mux__state_55 | new_and_mux__state_55_2;
  assign new_s__state_57 = new__state_57;
  assign new_not_s__state_57 = ~new_s__state_57;
  assign new_I0__state_57 = new_y_mux_56;
  assign new_I1__state_57 = new_y_mux_57;
  assign new_and_mux__state_57 = new_not_s__state_57 & new_I0__state_57;
  assign new_and_mux__state_57_2 = new_s__state_57 & new_I1__state_57;
  assign new_y_mux_60 = new_and_mux__state_57 | new_and_mux__state_57_2;
  assign new_s__state_59 = new__state_59;
  assign new_not_s__state_59 = ~new_s__state_59;
  assign new_I0__state_59 = new_y_mux_58;
  assign new_I1__state_59 = new_y_mux_59;
  assign new_and_mux__state_59 = new_not_s__state_59 & new_I0__state_59;
  assign new_and_mux__state_59_2 = new_s__state_59 & new_I1__state_59;
  assign new_y_mux_61 = new_and_mux__state_59 | new_and_mux__state_59_2;
  assign new_s__state_61 = new__state_61;
  assign new_not_s__state_61 = ~new_s__state_61;
  assign new_I0__state_61 = new_y_mux_60;
  assign new_I1__state_61 = new_y_mux_61;
  assign new_and_mux__state_61 = new_not_s__state_61 & new_I0__state_61;
  assign new_and_mux__state_61_2 = new_s__state_61 & new_I1__state_61;
  assign n174 = new_and_mux__state_61 | new_and_mux__state_61_2;
  always @ (posedge clock) begin
    P1_IR_REG_0_ <= n174;
    P1_IR_REG_1_ <= n179;
    P1_IR_REG_2_ <= n184;
    P1_IR_REG_3_ <= n189;
    P1_IR_REG_4_ <= n194;
    P1_IR_REG_5_ <= n199;
    P1_IR_REG_6_ <= n204;
    P1_IR_REG_7_ <= n209;
    P1_IR_REG_8_ <= n214;
    P1_IR_REG_9_ <= n219;
    P1_IR_REG_10_ <= n224;
    P1_IR_REG_11_ <= n229;
    P1_IR_REG_12_ <= n234;
    P1_IR_REG_13_ <= n239;
    P1_IR_REG_14_ <= n244;
    P1_IR_REG_15_ <= n249;
    P1_IR_REG_16_ <= n254;
    P1_IR_REG_17_ <= n259;
    P1_IR_REG_18_ <= n264;
    P1_IR_REG_19_ <= n269;
    P1_IR_REG_20_ <= n274;
    P1_IR_REG_21_ <= n279;
    P1_IR_REG_22_ <= n284;
    P1_IR_REG_23_ <= n289;
    P1_IR_REG_24_ <= n294;
    P1_IR_REG_25_ <= n299;
    P1_IR_REG_26_ <= n304;
    P1_IR_REG_27_ <= n309;
    P1_IR_REG_28_ <= n314;
    P1_IR_REG_29_ <= n319;
    P1_IR_REG_30_ <= n324;
    P1_IR_REG_31_ <= n329;
    P1_D_REG_0_ <= n334;
    P1_D_REG_1_ <= n339;
    P1_D_REG_2_ <= n344;
    P1_D_REG_3_ <= n349;
    P1_D_REG_4_ <= n354;
    P1_D_REG_5_ <= n359;
    P1_D_REG_6_ <= n364;
    P1_D_REG_7_ <= n369;
    P1_D_REG_8_ <= n374;
    P1_D_REG_9_ <= n379;
    P1_D_REG_10_ <= n384;
    P1_D_REG_11_ <= n389;
    P1_D_REG_12_ <= n394;
    P1_D_REG_13_ <= n399;
    P1_D_REG_14_ <= n404;
    P1_D_REG_15_ <= n409;
    P1_D_REG_16_ <= n414;
    P1_D_REG_17_ <= n419;
    P1_D_REG_18_ <= n424;
    P1_D_REG_19_ <= n429;
    P1_D_REG_20_ <= n434;
    P1_D_REG_21_ <= n439;
    P1_D_REG_22_ <= n444;
    P1_D_REG_23_ <= n449;
    P1_D_REG_24_ <= n454;
    P1_D_REG_25_ <= n459;
    P1_D_REG_26_ <= n464;
    P1_D_REG_27_ <= n469;
    P1_D_REG_28_ <= n474;
    P1_D_REG_29_ <= n479;
    P1_D_REG_30_ <= n484;
    P1_D_REG_31_ <= n489;
    P1_REG0_REG_0_ <= n494;
    P1_REG0_REG_1_ <= n499;
    P1_REG0_REG_2_ <= n504;
    P1_REG0_REG_3_ <= n509;
    P1_REG0_REG_4_ <= n514;
    P1_REG0_REG_5_ <= n519;
    P1_REG0_REG_6_ <= n524;
    P1_REG0_REG_7_ <= n529;
    P1_REG0_REG_8_ <= n534;
    P1_REG0_REG_9_ <= n539;
    P1_REG0_REG_10_ <= n544;
    P1_REG0_REG_11_ <= n549;
    P1_REG0_REG_12_ <= n554;
    P1_REG0_REG_13_ <= n559;
    P1_REG0_REG_14_ <= n564;
    P1_REG0_REG_15_ <= n569;
    P1_REG0_REG_16_ <= n574;
    P1_REG0_REG_17_ <= n579;
    P1_REG0_REG_18_ <= n584;
    P1_REG0_REG_19_ <= n589;
    P1_REG0_REG_20_ <= n594;
    P1_REG0_REG_21_ <= n599;
    P1_REG0_REG_22_ <= n604;
    P1_REG0_REG_23_ <= n609;
    P1_REG0_REG_24_ <= n614;
    P1_REG0_REG_25_ <= n619;
    P1_REG0_REG_26_ <= n624;
    P1_REG0_REG_27_ <= n629;
    P1_REG0_REG_28_ <= n634;
    P1_REG0_REG_29_ <= n639;
    P1_REG0_REG_30_ <= n644;
    P1_REG0_REG_31_ <= n649;
    P1_REG1_REG_0_ <= n654;
    P1_REG1_REG_1_ <= n659;
    P1_REG1_REG_2_ <= n664;
    P1_REG1_REG_3_ <= n669;
    P1_REG1_REG_4_ <= n674;
    P1_REG1_REG_5_ <= n679;
    P1_REG1_REG_6_ <= n684;
    P1_REG1_REG_7_ <= n689;
    P1_REG1_REG_8_ <= n694;
    P1_REG1_REG_9_ <= n699;
    P1_REG1_REG_10_ <= n704;
    P1_REG1_REG_11_ <= n709;
    P1_REG1_REG_12_ <= n714;
    P1_REG1_REG_13_ <= n719;
    P1_REG1_REG_14_ <= n724;
    P1_REG1_REG_15_ <= n729;
    P1_REG1_REG_16_ <= n734;
    P1_REG1_REG_17_ <= n739;
    P1_REG1_REG_18_ <= n744;
    P1_REG1_REG_19_ <= n749;
    P1_REG1_REG_20_ <= n754;
    P1_REG1_REG_21_ <= n759;
    P1_REG1_REG_22_ <= n764;
    P1_REG1_REG_23_ <= n769;
    P1_REG1_REG_24_ <= n774;
    P1_REG1_REG_25_ <= n779;
    P1_REG1_REG_26_ <= n784;
    P1_REG1_REG_27_ <= n789;
    P1_REG1_REG_28_ <= n794;
    P1_REG1_REG_29_ <= n799;
    P1_REG1_REG_30_ <= n804;
    P1_REG1_REG_31_ <= n809;
    P1_REG2_REG_0_ <= n814;
    P1_REG2_REG_1_ <= n819;
    P1_REG2_REG_2_ <= n824;
    P1_REG2_REG_3_ <= n829;
    P1_REG2_REG_4_ <= n834;
    P1_REG2_REG_5_ <= n839;
    P1_REG2_REG_6_ <= n844;
    P1_REG2_REG_7_ <= n849;
    P1_REG2_REG_8_ <= n854;
    P1_REG2_REG_9_ <= n859;
    P1_REG2_REG_10_ <= n864;
    P1_REG2_REG_11_ <= n869;
    P1_REG2_REG_12_ <= n874;
    P1_REG2_REG_13_ <= n879;
    P1_REG2_REG_14_ <= n884;
    P1_REG2_REG_15_ <= n889;
    P1_REG2_REG_16_ <= n894;
    P1_REG2_REG_17_ <= n899;
    P1_REG2_REG_18_ <= n904;
    P1_REG2_REG_19_ <= n909;
    P1_REG2_REG_20_ <= n914;
    P1_REG2_REG_21_ <= n919;
    P1_REG2_REG_22_ <= n924;
    P1_REG2_REG_23_ <= n929;
    P1_REG2_REG_24_ <= n934;
    P1_REG2_REG_25_ <= n939;
    P1_REG2_REG_26_ <= n944;
    P1_REG2_REG_27_ <= n949;
    P1_REG2_REG_28_ <= n954;
    P1_REG2_REG_29_ <= n959;
    P1_REG2_REG_30_ <= n964;
    P1_REG2_REG_31_ <= n969;
    P1_ADDR_REG_19_ <= n974;
    P1_ADDR_REG_18_ <= n979;
    P1_ADDR_REG_17_ <= n984;
    P1_ADDR_REG_16_ <= n989;
    P1_ADDR_REG_15_ <= n994;
    P1_ADDR_REG_14_ <= n999;
    P1_ADDR_REG_13_ <= n1004;
    P1_ADDR_REG_12_ <= n1009;
    P1_ADDR_REG_11_ <= n1014;
    P1_ADDR_REG_10_ <= n1019;
    P1_ADDR_REG_9_ <= n1024;
    P1_ADDR_REG_8_ <= n1029;
    P1_ADDR_REG_7_ <= n1034;
    P1_ADDR_REG_6_ <= n1039;
    P1_ADDR_REG_5_ <= n1044;
    P1_ADDR_REG_4_ <= n1049;
    P1_ADDR_REG_3_ <= n1054;
    P1_ADDR_REG_2_ <= n1059;
    P1_ADDR_REG_1_ <= n1064;
    P1_ADDR_REG_0_ <= n1069;
    P1_DATAO_REG_0_ <= n1074;
    P1_DATAO_REG_1_ <= n1079;
    P1_DATAO_REG_2_ <= n1084;
    P1_DATAO_REG_3_ <= n1089;
    P1_DATAO_REG_4_ <= n1094;
    P1_DATAO_REG_5_ <= n1099;
    P1_DATAO_REG_6_ <= n1104;
    P1_DATAO_REG_7_ <= n1109;
    P1_DATAO_REG_8_ <= n1114;
    P1_DATAO_REG_9_ <= n1119;
    P1_DATAO_REG_10_ <= n1124;
    P1_DATAO_REG_11_ <= n1129;
    P1_DATAO_REG_12_ <= n1134;
    P1_DATAO_REG_13_ <= n1139;
    P1_DATAO_REG_14_ <= n1144;
    P1_DATAO_REG_15_ <= n1149;
    P1_DATAO_REG_16_ <= n1154;
    P1_DATAO_REG_17_ <= n1159;
    P1_DATAO_REG_18_ <= n1164;
    P1_DATAO_REG_19_ <= n1169;
    P1_DATAO_REG_20_ <= n1174;
    P1_DATAO_REG_21_ <= n1179;
    P1_DATAO_REG_22_ <= n1184;
    P1_DATAO_REG_23_ <= n1189;
    P1_DATAO_REG_24_ <= n1194;
    P1_DATAO_REG_25_ <= n1199;
    P1_DATAO_REG_26_ <= n1204;
    P1_DATAO_REG_27_ <= n1209;
    P1_DATAO_REG_28_ <= n1214;
    P1_DATAO_REG_29_ <= n1219;
    P1_DATAO_REG_30_ <= n1224;
    P1_DATAO_REG_31_ <= n1229;
    P1_B_REG <= n1234;
    P1_REG3_REG_15_ <= n1239;
    P1_REG3_REG_26_ <= n1244;
    P1_REG3_REG_6_ <= n1249;
    P1_REG3_REG_18_ <= n1254;
    P1_REG3_REG_2_ <= n1259;
    P1_REG3_REG_11_ <= n1264;
    P1_REG3_REG_22_ <= n1269;
    P1_REG3_REG_13_ <= n1274;
    P1_REG3_REG_20_ <= n1279;
    P1_REG3_REG_0_ <= n1284;
    P1_REG3_REG_9_ <= n1289;
    P1_REG3_REG_4_ <= n1294;
    P1_REG3_REG_24_ <= n1299;
    P1_REG3_REG_17_ <= n1304;
    P1_REG3_REG_5_ <= n1309;
    P1_REG3_REG_16_ <= n1314;
    P1_REG3_REG_25_ <= n1319;
    P1_REG3_REG_12_ <= n1324;
    P1_REG3_REG_21_ <= n1329;
    P1_REG3_REG_1_ <= n1334;
    P1_REG3_REG_8_ <= n1339;
    P1_REG3_REG_28_ <= n1344;
    P1_REG3_REG_19_ <= n1349;
    P1_REG3_REG_3_ <= n1354;
    P1_REG3_REG_10_ <= n1359;
    P1_REG3_REG_23_ <= n1364;
    P1_REG3_REG_14_ <= n1369;
    P1_REG3_REG_27_ <= n1374;
    P1_REG3_REG_7_ <= n1379;
    P1_STATE_REG <= n1384;
    P1_RD_REG <= n1389;
    P1_WR_REG <= n1394;
    P2_IR_REG_0_ <= n1399;
    P2_IR_REG_1_ <= n1404;
    P2_IR_REG_2_ <= n1409;
    P2_IR_REG_3_ <= n1414;
    P2_IR_REG_4_ <= n1419;
    P2_IR_REG_5_ <= n1424;
    P2_IR_REG_6_ <= n1429;
    P2_IR_REG_7_ <= n1434;
    P2_IR_REG_8_ <= n1439;
    P2_IR_REG_9_ <= n1444;
    P2_IR_REG_10_ <= n1449;
    P2_IR_REG_11_ <= n1454;
    P2_IR_REG_12_ <= n1459;
    P2_IR_REG_13_ <= n1464;
    P2_IR_REG_14_ <= n1469;
    P2_IR_REG_15_ <= n1474;
    P2_IR_REG_16_ <= n1479;
    P2_IR_REG_17_ <= n1484;
    P2_IR_REG_18_ <= n1489;
    P2_IR_REG_19_ <= n1494;
    P2_IR_REG_20_ <= n1499;
    P2_IR_REG_21_ <= n1504;
    P2_IR_REG_22_ <= n1509;
    P2_IR_REG_23_ <= n1514;
    P2_IR_REG_24_ <= n1519;
    P2_IR_REG_25_ <= n1524;
    P2_IR_REG_26_ <= n1529;
    P2_IR_REG_27_ <= n1534;
    P2_IR_REG_28_ <= n1539;
    P2_IR_REG_29_ <= n1544;
    P2_IR_REG_30_ <= n1549;
    P2_IR_REG_31_ <= n1554;
    P2_D_REG_0_ <= n1559;
    P2_D_REG_1_ <= n1564;
    P2_D_REG_2_ <= n1569;
    P2_D_REG_3_ <= n1574;
    P2_D_REG_4_ <= n1579;
    P2_D_REG_5_ <= n1584;
    P2_D_REG_6_ <= n1589;
    P2_D_REG_7_ <= n1594;
    P2_D_REG_8_ <= n1599;
    P2_D_REG_9_ <= n1604;
    P2_D_REG_10_ <= n1609;
    P2_D_REG_11_ <= n1614;
    P2_D_REG_12_ <= n1619;
    P2_D_REG_13_ <= n1624;
    P2_D_REG_14_ <= n1629;
    P2_D_REG_15_ <= n1634;
    P2_D_REG_16_ <= n1639;
    P2_D_REG_17_ <= n1644;
    P2_D_REG_18_ <= n1649;
    P2_D_REG_19_ <= n1654;
    P2_D_REG_20_ <= n1659;
    P2_D_REG_21_ <= n1664;
    P2_D_REG_22_ <= n1669;
    P2_D_REG_23_ <= n1674;
    P2_D_REG_24_ <= n1679;
    P2_D_REG_25_ <= n1684;
    P2_D_REG_26_ <= n1689;
    P2_D_REG_27_ <= n1694;
    P2_D_REG_28_ <= n1699;
    P2_D_REG_29_ <= n1704;
    P2_D_REG_30_ <= n1709;
    P2_D_REG_31_ <= n1714;
    P2_REG0_REG_0_ <= n1719;
    P2_REG0_REG_1_ <= n1724;
    P2_REG0_REG_2_ <= n1729;
    P2_REG0_REG_3_ <= n1734;
    P2_REG0_REG_4_ <= n1739;
    P2_REG0_REG_5_ <= n1744;
    P2_REG0_REG_6_ <= n1749;
    P2_REG0_REG_7_ <= n1754;
    P2_REG0_REG_8_ <= n1759;
    P2_REG0_REG_9_ <= n1764;
    P2_REG0_REG_10_ <= n1769;
    P2_REG0_REG_11_ <= n1774;
    P2_REG0_REG_12_ <= n1779;
    P2_REG0_REG_13_ <= n1784;
    P2_REG0_REG_14_ <= n1789;
    P2_REG0_REG_15_ <= n1794;
    P2_REG0_REG_16_ <= n1799;
    P2_REG0_REG_17_ <= n1804;
    P2_REG0_REG_18_ <= n1809;
    P2_REG0_REG_19_ <= n1814;
    P2_REG0_REG_20_ <= n1819;
    P2_REG0_REG_21_ <= n1824;
    P2_REG0_REG_22_ <= n1829;
    P2_REG0_REG_23_ <= n1834;
    P2_REG0_REG_24_ <= n1839;
    P2_REG0_REG_25_ <= n1844;
    P2_REG0_REG_26_ <= n1849;
    P2_REG0_REG_27_ <= n1854;
    P2_REG0_REG_28_ <= n1859;
    P2_REG0_REG_29_ <= n1864;
    P2_REG0_REG_30_ <= n1869;
    P2_REG0_REG_31_ <= n1874;
    P2_REG1_REG_0_ <= n1879;
    P2_REG1_REG_1_ <= n1884;
    P2_REG1_REG_2_ <= n1889;
    P2_REG1_REG_3_ <= n1894;
    P2_REG1_REG_4_ <= n1899;
    P2_REG1_REG_5_ <= n1904;
    P2_REG1_REG_6_ <= n1909;
    P2_REG1_REG_7_ <= n1914;
    P2_REG1_REG_8_ <= n1919;
    P2_REG1_REG_9_ <= n1924;
    P2_REG1_REG_10_ <= n1929;
    P2_REG1_REG_11_ <= n1934;
    P2_REG1_REG_12_ <= n1939;
    P2_REG1_REG_13_ <= n1944;
    P2_REG1_REG_14_ <= n1949;
    P2_REG1_REG_15_ <= n1954;
    P2_REG1_REG_16_ <= n1959;
    P2_REG1_REG_17_ <= n1964;
    P2_REG1_REG_18_ <= n1969;
    P2_REG1_REG_19_ <= n1974;
    P2_REG1_REG_20_ <= n1979;
    P2_REG1_REG_21_ <= n1984;
    P2_REG1_REG_22_ <= n1989;
    P2_REG1_REG_23_ <= n1994;
    P2_REG1_REG_24_ <= n1999;
    P2_REG1_REG_25_ <= n2004;
    P2_REG1_REG_26_ <= n2009;
    P2_REG1_REG_27_ <= n2014;
    P2_REG1_REG_28_ <= n2019;
    P2_REG1_REG_29_ <= n2024;
    P2_REG1_REG_30_ <= n2029;
    P2_REG1_REG_31_ <= n2034;
    P2_REG2_REG_0_ <= n2039;
    P2_REG2_REG_1_ <= n2044;
    P2_REG2_REG_2_ <= n2049;
    P2_REG2_REG_3_ <= n2054;
    P2_REG2_REG_4_ <= n2059;
    P2_REG2_REG_5_ <= n2064;
    P2_REG2_REG_6_ <= n2069;
    P2_REG2_REG_7_ <= n2074;
    P2_REG2_REG_8_ <= n2079;
    P2_REG2_REG_9_ <= n2084;
    P2_REG2_REG_10_ <= n2089;
    P2_REG2_REG_11_ <= n2094;
    P2_REG2_REG_12_ <= n2099;
    P2_REG2_REG_13_ <= n2104;
    P2_REG2_REG_14_ <= n2109;
    P2_REG2_REG_15_ <= n2114;
    P2_REG2_REG_16_ <= n2119;
    P2_REG2_REG_17_ <= n2124;
    P2_REG2_REG_18_ <= n2129;
    P2_REG2_REG_19_ <= n2134;
    P2_REG2_REG_20_ <= n2139;
    P2_REG2_REG_21_ <= n2144;
    P2_REG2_REG_22_ <= n2149;
    P2_REG2_REG_23_ <= n2154;
    P2_REG2_REG_24_ <= n2159;
    P2_REG2_REG_25_ <= n2164;
    P2_REG2_REG_26_ <= n2169;
    P2_REG2_REG_27_ <= n2174;
    P2_REG2_REG_28_ <= n2179;
    P2_REG2_REG_29_ <= n2184;
    P2_REG2_REG_30_ <= n2189;
    P2_REG2_REG_31_ <= n2194;
    P2_ADDR_REG_19_ <= n2199;
    P2_ADDR_REG_18_ <= n2204;
    P2_ADDR_REG_17_ <= n2209;
    P2_ADDR_REG_16_ <= n2214;
    P2_ADDR_REG_15_ <= n2219;
    P2_ADDR_REG_14_ <= n2224;
    P2_ADDR_REG_13_ <= n2229;
    P2_ADDR_REG_12_ <= n2234;
    P2_ADDR_REG_11_ <= n2239;
    P2_ADDR_REG_10_ <= n2244;
    P2_ADDR_REG_9_ <= n2249;
    P2_ADDR_REG_8_ <= n2254;
    P2_ADDR_REG_7_ <= n2259;
    P2_ADDR_REG_6_ <= n2264;
    P2_ADDR_REG_5_ <= n2269;
    P2_ADDR_REG_4_ <= n2274;
    P2_ADDR_REG_3_ <= n2279;
    P2_ADDR_REG_2_ <= n2284;
    P2_ADDR_REG_1_ <= n2289;
    P2_ADDR_REG_0_ <= n2294;
    P2_DATAO_REG_0_ <= n2299;
    P2_DATAO_REG_1_ <= n2304;
    P2_DATAO_REG_2_ <= n2309;
    P2_DATAO_REG_3_ <= n2314;
    P2_DATAO_REG_4_ <= n2319;
    P2_DATAO_REG_5_ <= n2324;
    P2_DATAO_REG_6_ <= n2329;
    P2_DATAO_REG_7_ <= n2334;
    P2_DATAO_REG_8_ <= n2339;
    P2_DATAO_REG_9_ <= n2344;
    P2_DATAO_REG_10_ <= n2349;
    P2_DATAO_REG_11_ <= n2354;
    P2_DATAO_REG_12_ <= n2359;
    P2_DATAO_REG_13_ <= n2364;
    P2_DATAO_REG_14_ <= n2369;
    P2_DATAO_REG_15_ <= n2374;
    P2_DATAO_REG_16_ <= n2379;
    P2_DATAO_REG_17_ <= n2384;
    P2_DATAO_REG_18_ <= n2389;
    P2_DATAO_REG_19_ <= n2394;
    P2_DATAO_REG_20_ <= n2399;
    P2_DATAO_REG_21_ <= n2404;
    P2_DATAO_REG_22_ <= n2409;
    P2_DATAO_REG_23_ <= n2414;
    P2_DATAO_REG_24_ <= n2419;
    P2_DATAO_REG_25_ <= n2424;
    P2_DATAO_REG_26_ <= n2429;
    P2_DATAO_REG_27_ <= n2434;
    P2_DATAO_REG_28_ <= n2439;
    P2_DATAO_REG_29_ <= n2444;
    P2_DATAO_REG_30_ <= n2449;
    P2_DATAO_REG_31_ <= n2454;
    P2_B_REG <= n2459;
    P2_REG3_REG_15_ <= n2464;
    P2_REG3_REG_26_ <= n2469;
    P2_REG3_REG_6_ <= n2474;
    P2_REG3_REG_18_ <= n2479;
    P2_REG3_REG_2_ <= n2484;
    P2_REG3_REG_11_ <= n2489;
    P2_REG3_REG_22_ <= n2494;
    P2_REG3_REG_13_ <= n2499;
    P2_REG3_REG_20_ <= n2504;
    P2_REG3_REG_0_ <= n2509;
    P2_REG3_REG_9_ <= n2514;
    P2_REG3_REG_4_ <= n2519;
    P2_REG3_REG_24_ <= n2524;
    P2_REG3_REG_17_ <= n2529;
    P2_REG3_REG_5_ <= n2534;
    P2_REG3_REG_16_ <= n2539;
    P2_REG3_REG_25_ <= n2544;
    P2_REG3_REG_12_ <= n2549;
    P2_REG3_REG_21_ <= n2554;
    P2_REG3_REG_1_ <= n2559;
    P2_REG3_REG_8_ <= n2564;
    P2_REG3_REG_28_ <= n2569;
    P2_REG3_REG_19_ <= n2574;
    P2_REG3_REG_3_ <= n2579;
    P2_REG3_REG_10_ <= n2584;
    P2_REG3_REG_23_ <= n2589;
    P2_REG3_REG_14_ <= n2594;
    P2_REG3_REG_27_ <= n2599;
    P2_REG3_REG_7_ <= n2604;
    P2_STATE_REG <= n2609;
    P2_RD_REG <= n2614;
    P2_WR_REG <= n2619;
    P3_IR_REG_0_ <= n2624;
    P3_IR_REG_1_ <= n2629;
    P3_IR_REG_2_ <= n2634;
    P3_IR_REG_3_ <= n2639;
    P3_IR_REG_4_ <= n2644;
    P3_IR_REG_5_ <= n2649;
    P3_IR_REG_6_ <= n2654;
    P3_IR_REG_7_ <= n2659;
    P3_IR_REG_8_ <= n2664;
    P3_IR_REG_9_ <= n2669;
    P3_IR_REG_10_ <= n2674;
    P3_IR_REG_11_ <= n2679;
    P3_IR_REG_12_ <= n2684;
    P3_IR_REG_13_ <= n2689;
    P3_IR_REG_14_ <= n2694;
    P3_IR_REG_15_ <= n2699;
    P3_IR_REG_16_ <= n2704;
    P3_IR_REG_17_ <= n2709;
    P3_IR_REG_18_ <= n2714;
    P3_IR_REG_19_ <= n2719;
    P3_IR_REG_20_ <= n2724;
    P3_IR_REG_21_ <= n2729;
    P3_IR_REG_22_ <= n2734;
    P3_IR_REG_23_ <= n2739;
    P3_IR_REG_24_ <= n2744;
    P3_IR_REG_25_ <= n2749;
    P3_IR_REG_26_ <= n2754;
    P3_IR_REG_27_ <= n2759;
    P3_IR_REG_28_ <= n2764;
    P3_IR_REG_29_ <= n2769;
    P3_IR_REG_30_ <= n2774;
    P3_IR_REG_31_ <= n2779;
    P3_D_REG_0_ <= n2784;
    P3_D_REG_1_ <= n2789;
    P3_D_REG_2_ <= n2794;
    P3_D_REG_3_ <= n2799;
    P3_D_REG_4_ <= n2804;
    P3_D_REG_5_ <= n2809;
    P3_D_REG_6_ <= n2814;
    P3_D_REG_7_ <= n2819;
    P3_D_REG_8_ <= n2824;
    P3_D_REG_9_ <= n2829;
    P3_D_REG_10_ <= n2834;
    P3_D_REG_11_ <= n2839;
    P3_D_REG_12_ <= n2844;
    P3_D_REG_13_ <= n2849;
    P3_D_REG_14_ <= n2854;
    P3_D_REG_15_ <= n2859;
    P3_D_REG_16_ <= n2864;
    P3_D_REG_17_ <= n2869;
    P3_D_REG_18_ <= n2874;
    P3_D_REG_19_ <= n2879;
    P3_D_REG_20_ <= n2884;
    P3_D_REG_21_ <= n2889;
    P3_D_REG_22_ <= n2894;
    P3_D_REG_23_ <= n2899;
    P3_D_REG_24_ <= n2904;
    P3_D_REG_25_ <= n2909;
    P3_D_REG_26_ <= n2914;
    P3_D_REG_27_ <= n2919;
    P3_D_REG_28_ <= n2924;
    P3_D_REG_29_ <= n2929;
    P3_D_REG_30_ <= n2934;
    P3_D_REG_31_ <= n2939;
    P3_REG0_REG_0_ <= n2944;
    P3_REG0_REG_1_ <= n2949;
    P3_REG0_REG_2_ <= n2954;
    P3_REG0_REG_3_ <= n2959;
    P3_REG0_REG_4_ <= n2964;
    P3_REG0_REG_5_ <= n2969;
    P3_REG0_REG_6_ <= n2974;
    P3_REG0_REG_7_ <= n2979;
    P3_REG0_REG_8_ <= n2984;
    P3_REG0_REG_9_ <= n2989;
    P3_REG0_REG_10_ <= n2994;
    P3_REG0_REG_11_ <= n2999;
    P3_REG0_REG_12_ <= n3004;
    P3_REG0_REG_13_ <= n3009;
    P3_REG0_REG_14_ <= n3014;
    P3_REG0_REG_15_ <= n3019;
    P3_REG0_REG_16_ <= n3024;
    P3_REG0_REG_17_ <= n3029;
    P3_REG0_REG_18_ <= n3034;
    P3_REG0_REG_19_ <= n3039;
    P3_REG0_REG_20_ <= n3044;
    P3_REG0_REG_21_ <= n3049;
    P3_REG0_REG_22_ <= n3054;
    P3_REG0_REG_23_ <= n3059;
    P3_REG0_REG_24_ <= n3064;
    P3_REG0_REG_25_ <= n3069;
    P3_REG0_REG_26_ <= n3074;
    P3_REG0_REG_27_ <= n3079;
    P3_REG0_REG_28_ <= n3084;
    P3_REG0_REG_29_ <= n3089;
    P3_REG0_REG_30_ <= n3094;
    P3_REG0_REG_31_ <= n3099;
    P3_REG1_REG_0_ <= n3104;
    P3_REG1_REG_1_ <= n3109;
    P3_REG1_REG_2_ <= n3114;
    P3_REG1_REG_3_ <= n3119;
    P3_REG1_REG_4_ <= n3124;
    P3_REG1_REG_5_ <= n3129;
    P3_REG1_REG_6_ <= n3134;
    P3_REG1_REG_7_ <= n3139;
    P3_REG1_REG_8_ <= n3144;
    P3_REG1_REG_9_ <= n3149;
    P3_REG1_REG_10_ <= n3154;
    P3_REG1_REG_11_ <= n3159;
    P3_REG1_REG_12_ <= n3164;
    P3_REG1_REG_13_ <= n3169;
    P3_REG1_REG_14_ <= n3174;
    P3_REG1_REG_15_ <= n3179;
    P3_REG1_REG_16_ <= n3184;
    P3_REG1_REG_17_ <= n3189;
    P3_REG1_REG_18_ <= n3194;
    P3_REG1_REG_19_ <= n3199;
    P3_REG1_REG_20_ <= n3204;
    P3_REG1_REG_21_ <= n3209;
    P3_REG1_REG_22_ <= n3214;
    P3_REG1_REG_23_ <= n3219;
    P3_REG1_REG_24_ <= n3224;
    P3_REG1_REG_25_ <= n3229;
    P3_REG1_REG_26_ <= n3234;
    P3_REG1_REG_27_ <= n3239;
    P3_REG1_REG_28_ <= n3244;
    P3_REG1_REG_29_ <= n3249;
    P3_REG1_REG_30_ <= n3254;
    P3_REG1_REG_31_ <= n3259;
    P3_REG2_REG_0_ <= n3264;
    P3_REG2_REG_1_ <= n3269;
    P3_REG2_REG_2_ <= n3274;
    P3_REG2_REG_3_ <= n3279;
    P3_REG2_REG_4_ <= n3284;
    P3_REG2_REG_5_ <= n3289;
    P3_REG2_REG_6_ <= n3294;
    P3_REG2_REG_7_ <= n3299;
    P3_REG2_REG_8_ <= n3304;
    P3_REG2_REG_9_ <= n3309;
    P3_REG2_REG_10_ <= n3314;
    P3_REG2_REG_11_ <= n3319;
    P3_REG2_REG_12_ <= n3324;
    P3_REG2_REG_13_ <= n3329;
    P3_REG2_REG_14_ <= n3334;
    P3_REG2_REG_15_ <= n3339;
    P3_REG2_REG_16_ <= n3344;
    P3_REG2_REG_17_ <= n3349;
    P3_REG2_REG_18_ <= n3354;
    P3_REG2_REG_19_ <= n3359;
    P3_REG2_REG_20_ <= n3364;
    P3_REG2_REG_21_ <= n3369;
    P3_REG2_REG_22_ <= n3374;
    P3_REG2_REG_23_ <= n3379;
    P3_REG2_REG_24_ <= n3384;
    P3_REG2_REG_25_ <= n3389;
    P3_REG2_REG_26_ <= n3394;
    P3_REG2_REG_27_ <= n3399;
    P3_REG2_REG_28_ <= n3404;
    P3_REG2_REG_29_ <= n3409;
    P3_REG2_REG_30_ <= n3414;
    P3_REG2_REG_31_ <= n3419;
    P3_ADDR_REG_19_ <= n3424;
    P3_ADDR_REG_18_ <= n3429;
    P3_ADDR_REG_17_ <= n3434;
    P3_ADDR_REG_16_ <= n3439;
    P3_ADDR_REG_15_ <= n3444;
    P3_ADDR_REG_14_ <= n3449;
    P3_ADDR_REG_13_ <= n3454;
    P3_ADDR_REG_12_ <= n3459;
    P3_ADDR_REG_11_ <= n3464;
    P3_ADDR_REG_10_ <= n3469;
    P3_ADDR_REG_9_ <= n3474;
    P3_ADDR_REG_8_ <= n3479;
    P3_ADDR_REG_7_ <= n3484;
    P3_ADDR_REG_6_ <= n3489;
    P3_ADDR_REG_5_ <= n3494;
    P3_ADDR_REG_4_ <= n3499;
    P3_ADDR_REG_3_ <= n3504;
    P3_ADDR_REG_2_ <= n3509;
    P3_ADDR_REG_1_ <= n3514;
    P3_ADDR_REG_0_ <= n3519;
    P3_DATAO_REG_0_ <= n3524;
    P3_DATAO_REG_1_ <= n3529;
    P3_DATAO_REG_2_ <= n3534;
    P3_DATAO_REG_3_ <= n3539;
    P3_DATAO_REG_4_ <= n3544;
    P3_DATAO_REG_5_ <= n3549;
    P3_DATAO_REG_6_ <= n3554;
    P3_DATAO_REG_7_ <= n3559;
    P3_DATAO_REG_8_ <= n3564;
    P3_DATAO_REG_9_ <= n3569;
    P3_DATAO_REG_10_ <= n3574;
    P3_DATAO_REG_11_ <= n3579;
    P3_DATAO_REG_12_ <= n3584;
    P3_DATAO_REG_13_ <= n3589;
    P3_DATAO_REG_14_ <= n3594;
    P3_DATAO_REG_15_ <= n3599;
    P3_DATAO_REG_16_ <= n3604;
    P3_DATAO_REG_17_ <= n3609;
    P3_DATAO_REG_18_ <= n3614;
    P3_DATAO_REG_19_ <= n3619;
    P3_DATAO_REG_20_ <= n3624;
    P3_DATAO_REG_21_ <= n3629;
    P3_DATAO_REG_22_ <= n3634;
    P3_DATAO_REG_23_ <= n3639;
    P3_DATAO_REG_24_ <= n3644;
    P3_DATAO_REG_25_ <= n3649;
    P3_DATAO_REG_26_ <= n3654;
    P3_DATAO_REG_27_ <= n3659;
    P3_DATAO_REG_28_ <= n3664;
    P3_DATAO_REG_29_ <= n3669;
    P3_DATAO_REG_30_ <= n3674;
    P3_DATAO_REG_31_ <= n3679;
    P3_B_REG <= n3684;
    P3_REG3_REG_15_ <= n3689;
    P3_REG3_REG_26_ <= n3694;
    P3_REG3_REG_6_ <= n3699;
    P3_REG3_REG_18_ <= n3704;
    P3_REG3_REG_2_ <= n3709;
    P3_REG3_REG_11_ <= n3714;
    P3_REG3_REG_22_ <= n3719;
    P3_REG3_REG_13_ <= n3724;
    P3_REG3_REG_20_ <= n3729;
    P3_REG3_REG_0_ <= n3734;
    P3_REG3_REG_9_ <= n3739;
    P3_REG3_REG_4_ <= n3744;
    P3_REG3_REG_24_ <= n3749;
    P3_REG3_REG_17_ <= n3754;
    P3_REG3_REG_5_ <= n3759;
    P3_REG3_REG_16_ <= n3764;
    P3_REG3_REG_25_ <= n3769;
    P3_REG3_REG_12_ <= n3774;
    P3_REG3_REG_21_ <= n3779;
    P3_REG3_REG_1_ <= n3784;
    P3_REG3_REG_8_ <= n3789;
    P3_REG3_REG_28_ <= n3794;
    P3_REG3_REG_19_ <= n3799;
    P3_REG3_REG_3_ <= n3804;
    P3_REG3_REG_10_ <= n3809;
    P3_REG3_REG_23_ <= n3814;
    P3_REG3_REG_14_ <= n3819;
    P3_REG3_REG_27_ <= n3824;
    P3_REG3_REG_7_ <= n3829;
    P3_STATE_REG <= n3834;
    P3_RD_REG <= n3839;
    P3_WR_REG <= n3844;
    Q_0 <= n61551;
    Q_1 <= n61554;
    Q_2 <= n61557;
    Q_3 <= n61560;
    Q_4 <= n61563;
  end
endmodule
