// Benchmark "./test_runs/structural2_16keys_5bits--s-120240927_165426/ITC99/b17_encrypted" written by ABC on Fri Sep 27 18:23:48 2024

module b17_encrypted  ( clock, 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, HOLD, NA, BS16, READY1, READY2, keyinput0, keyinput1,
    keyinput2, keyinput3, keyinput4,
    P3_DATAO_REG_31_, P3_DATAO_REG_30_, P3_DATAO_REG_29_, P3_DATAO_REG_28_,
    P3_DATAO_REG_27_, P3_DATAO_REG_26_, P3_DATAO_REG_25_, P3_DATAO_REG_24_,
    P3_DATAO_REG_23_, P3_DATAO_REG_22_, P3_DATAO_REG_21_, P3_DATAO_REG_20_,
    P3_DATAO_REG_19_, P3_DATAO_REG_18_, P3_DATAO_REG_17_, P3_DATAO_REG_16_,
    P3_DATAO_REG_15_, P3_DATAO_REG_14_, P3_DATAO_REG_13_, P3_DATAO_REG_12_,
    P3_DATAO_REG_11_, P3_DATAO_REG_10_, P3_DATAO_REG_9_, P3_DATAO_REG_8_,
    P3_DATAO_REG_7_, P3_DATAO_REG_6_, P3_DATAO_REG_5_, P3_DATAO_REG_4_,
    P3_DATAO_REG_3_, P3_DATAO_REG_2_, P3_DATAO_REG_1_, P3_DATAO_REG_0_,
    P1_ADDRESS_REG_29_, P1_ADDRESS_REG_28_, P1_ADDRESS_REG_27_,
    P1_ADDRESS_REG_26_, P1_ADDRESS_REG_25_, P1_ADDRESS_REG_24_,
    P1_ADDRESS_REG_23_, P1_ADDRESS_REG_22_, P1_ADDRESS_REG_21_,
    P1_ADDRESS_REG_20_, P1_ADDRESS_REG_19_, P1_ADDRESS_REG_18_,
    P1_ADDRESS_REG_17_, P1_ADDRESS_REG_16_, P1_ADDRESS_REG_15_,
    P1_ADDRESS_REG_14_, P1_ADDRESS_REG_13_, P1_ADDRESS_REG_12_,
    P1_ADDRESS_REG_11_, P1_ADDRESS_REG_10_, P1_ADDRESS_REG_9_,
    P1_ADDRESS_REG_8_, P1_ADDRESS_REG_7_, P1_ADDRESS_REG_6_,
    P1_ADDRESS_REG_5_, P1_ADDRESS_REG_4_, P1_ADDRESS_REG_3_,
    P1_ADDRESS_REG_2_, P1_ADDRESS_REG_1_, P1_ADDRESS_REG_0_, U355, U356,
    U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369,
    U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352,
    U353, U354, U365, U376, P3_W_R_N_REG, P3_D_C_N_REG, P3_M_IO_N_REG,
    P1_ADS_N_REG, P3_ADS_N_REG  );
  input  clock;
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2, keyinput0,
    keyinput1, keyinput2, keyinput3, keyinput4;
  output P3_DATAO_REG_31_, P3_DATAO_REG_30_, P3_DATAO_REG_29_,
    P3_DATAO_REG_28_, P3_DATAO_REG_27_, P3_DATAO_REG_26_, P3_DATAO_REG_25_,
    P3_DATAO_REG_24_, P3_DATAO_REG_23_, P3_DATAO_REG_22_, P3_DATAO_REG_21_,
    P3_DATAO_REG_20_, P3_DATAO_REG_19_, P3_DATAO_REG_18_, P3_DATAO_REG_17_,
    P3_DATAO_REG_16_, P3_DATAO_REG_15_, P3_DATAO_REG_14_, P3_DATAO_REG_13_,
    P3_DATAO_REG_12_, P3_DATAO_REG_11_, P3_DATAO_REG_10_, P3_DATAO_REG_9_,
    P3_DATAO_REG_8_, P3_DATAO_REG_7_, P3_DATAO_REG_6_, P3_DATAO_REG_5_,
    P3_DATAO_REG_4_, P3_DATAO_REG_3_, P3_DATAO_REG_2_, P3_DATAO_REG_1_,
    P3_DATAO_REG_0_, P1_ADDRESS_REG_29_, P1_ADDRESS_REG_28_,
    P1_ADDRESS_REG_27_, P1_ADDRESS_REG_26_, P1_ADDRESS_REG_25_,
    P1_ADDRESS_REG_24_, P1_ADDRESS_REG_23_, P1_ADDRESS_REG_22_,
    P1_ADDRESS_REG_21_, P1_ADDRESS_REG_20_, P1_ADDRESS_REG_19_,
    P1_ADDRESS_REG_18_, P1_ADDRESS_REG_17_, P1_ADDRESS_REG_16_,
    P1_ADDRESS_REG_15_, P1_ADDRESS_REG_14_, P1_ADDRESS_REG_13_,
    P1_ADDRESS_REG_12_, P1_ADDRESS_REG_11_, P1_ADDRESS_REG_10_,
    P1_ADDRESS_REG_9_, P1_ADDRESS_REG_8_, P1_ADDRESS_REG_7_,
    P1_ADDRESS_REG_6_, P1_ADDRESS_REG_5_, P1_ADDRESS_REG_4_,
    P1_ADDRESS_REG_3_, P1_ADDRESS_REG_2_, P1_ADDRESS_REG_1_,
    P1_ADDRESS_REG_0_, U355, U356, U357, U358, U359, U360, U361, U362,
    U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375,
    U347, U348, U349, U350, U351, U352, U353, U354, U365, U376,
    P3_W_R_N_REG, P3_D_C_N_REG, P3_M_IO_N_REG, P1_ADS_N_REG, P3_ADS_N_REG;
  reg BUF1_REG_0_, BUF1_REG_1_, BUF1_REG_2_, BUF1_REG_3_, BUF1_REG_4_,
    BUF1_REG_5_, BUF1_REG_6_, BUF1_REG_7_, BUF1_REG_8_, BUF1_REG_9_,
    BUF1_REG_10_, BUF1_REG_11_, BUF1_REG_12_, BUF1_REG_13_, BUF1_REG_14_,
    BUF1_REG_15_, BUF1_REG_16_, BUF1_REG_17_, BUF1_REG_18_, BUF1_REG_19_,
    BUF1_REG_20_, BUF1_REG_21_, BUF1_REG_22_, BUF1_REG_23_, BUF1_REG_24_,
    BUF1_REG_25_, BUF1_REG_26_, BUF1_REG_27_, BUF1_REG_28_, BUF1_REG_29_,
    BUF1_REG_30_, BUF1_REG_31_, BUF2_REG_0_, BUF2_REG_1_, BUF2_REG_2_,
    BUF2_REG_3_, BUF2_REG_4_, BUF2_REG_5_, BUF2_REG_6_, BUF2_REG_7_,
    BUF2_REG_8_, BUF2_REG_9_, BUF2_REG_10_, BUF2_REG_11_, BUF2_REG_12_,
    BUF2_REG_13_, BUF2_REG_14_, BUF2_REG_15_, BUF2_REG_16_, BUF2_REG_17_,
    BUF2_REG_18_, BUF2_REG_19_, BUF2_REG_20_, BUF2_REG_21_, BUF2_REG_22_,
    BUF2_REG_23_, BUF2_REG_24_, BUF2_REG_25_, BUF2_REG_26_, BUF2_REG_27_,
    BUF2_REG_28_, BUF2_REG_29_, BUF2_REG_30_, BUF2_REG_31_, READY12_REG,
    READY21_REG, READY22_REG, READY11_REG, P3_BE_N_REG_3_, P3_BE_N_REG_2_,
    P3_BE_N_REG_1_, P3_BE_N_REG_0_, P3_ADDRESS_REG_29_, P3_ADDRESS_REG_28_,
    P3_ADDRESS_REG_27_, P3_ADDRESS_REG_26_, P3_ADDRESS_REG_25_,
    P3_ADDRESS_REG_24_, P3_ADDRESS_REG_23_, P3_ADDRESS_REG_22_,
    P3_ADDRESS_REG_21_, P3_ADDRESS_REG_20_, P3_ADDRESS_REG_19_,
    P3_ADDRESS_REG_18_, P3_ADDRESS_REG_17_, P3_ADDRESS_REG_16_,
    P3_ADDRESS_REG_15_, P3_ADDRESS_REG_14_, P3_ADDRESS_REG_13_,
    P3_ADDRESS_REG_12_, P3_ADDRESS_REG_11_, P3_ADDRESS_REG_10_,
    P3_ADDRESS_REG_9_, P3_ADDRESS_REG_8_, P3_ADDRESS_REG_7_,
    P3_ADDRESS_REG_6_, P3_ADDRESS_REG_5_, P3_ADDRESS_REG_4_,
    P3_ADDRESS_REG_3_, P3_ADDRESS_REG_2_, P3_ADDRESS_REG_1_,
    P3_ADDRESS_REG_0_, P3_STATE_REG_2_, P3_STATE_REG_1_, P3_STATE_REG_0_,
    P3_DATAWIDTH_REG_0_, P3_DATAWIDTH_REG_1_, P3_DATAWIDTH_REG_2_,
    P3_DATAWIDTH_REG_3_, P3_DATAWIDTH_REG_4_, P3_DATAWIDTH_REG_5_,
    P3_DATAWIDTH_REG_6_, P3_DATAWIDTH_REG_7_, P3_DATAWIDTH_REG_8_,
    P3_DATAWIDTH_REG_9_, P3_DATAWIDTH_REG_10_, P3_DATAWIDTH_REG_11_,
    P3_DATAWIDTH_REG_12_, P3_DATAWIDTH_REG_13_, P3_DATAWIDTH_REG_14_,
    P3_DATAWIDTH_REG_15_, P3_DATAWIDTH_REG_16_, P3_DATAWIDTH_REG_17_,
    P3_DATAWIDTH_REG_18_, P3_DATAWIDTH_REG_19_, P3_DATAWIDTH_REG_20_,
    P3_DATAWIDTH_REG_21_, P3_DATAWIDTH_REG_22_, P3_DATAWIDTH_REG_23_,
    P3_DATAWIDTH_REG_24_, P3_DATAWIDTH_REG_25_, P3_DATAWIDTH_REG_26_,
    P3_DATAWIDTH_REG_27_, P3_DATAWIDTH_REG_28_, P3_DATAWIDTH_REG_29_,
    P3_DATAWIDTH_REG_30_, P3_DATAWIDTH_REG_31_, P3_STATE2_REG_3_,
    P3_STATE2_REG_2_, P3_STATE2_REG_1_, P3_STATE2_REG_0_,
    P3_INSTQUEUE_REG_15__7_, P3_INSTQUEUE_REG_15__6_,
    P3_INSTQUEUE_REG_15__5_, P3_INSTQUEUE_REG_15__4_,
    P3_INSTQUEUE_REG_15__3_, P3_INSTQUEUE_REG_15__2_,
    P3_INSTQUEUE_REG_15__1_, P3_INSTQUEUE_REG_15__0_,
    P3_INSTQUEUE_REG_14__7_, P3_INSTQUEUE_REG_14__6_,
    P3_INSTQUEUE_REG_14__5_, P3_INSTQUEUE_REG_14__4_,
    P3_INSTQUEUE_REG_14__3_, P3_INSTQUEUE_REG_14__2_,
    P3_INSTQUEUE_REG_14__1_, P3_INSTQUEUE_REG_14__0_,
    P3_INSTQUEUE_REG_13__7_, P3_INSTQUEUE_REG_13__6_,
    P3_INSTQUEUE_REG_13__5_, P3_INSTQUEUE_REG_13__4_,
    P3_INSTQUEUE_REG_13__3_, P3_INSTQUEUE_REG_13__2_,
    P3_INSTQUEUE_REG_13__1_, P3_INSTQUEUE_REG_13__0_,
    P3_INSTQUEUE_REG_12__7_, P3_INSTQUEUE_REG_12__6_,
    P3_INSTQUEUE_REG_12__5_, P3_INSTQUEUE_REG_12__4_,
    P3_INSTQUEUE_REG_12__3_, P3_INSTQUEUE_REG_12__2_,
    P3_INSTQUEUE_REG_12__1_, P3_INSTQUEUE_REG_12__0_,
    P3_INSTQUEUE_REG_11__7_, P3_INSTQUEUE_REG_11__6_,
    P3_INSTQUEUE_REG_11__5_, P3_INSTQUEUE_REG_11__4_,
    P3_INSTQUEUE_REG_11__3_, P3_INSTQUEUE_REG_11__2_,
    P3_INSTQUEUE_REG_11__1_, P3_INSTQUEUE_REG_11__0_,
    P3_INSTQUEUE_REG_10__7_, P3_INSTQUEUE_REG_10__6_,
    P3_INSTQUEUE_REG_10__5_, P3_INSTQUEUE_REG_10__4_,
    P3_INSTQUEUE_REG_10__3_, P3_INSTQUEUE_REG_10__2_,
    P3_INSTQUEUE_REG_10__1_, P3_INSTQUEUE_REG_10__0_,
    P3_INSTQUEUE_REG_9__7_, P3_INSTQUEUE_REG_9__6_, P3_INSTQUEUE_REG_9__5_,
    P3_INSTQUEUE_REG_9__4_, P3_INSTQUEUE_REG_9__3_, P3_INSTQUEUE_REG_9__2_,
    P3_INSTQUEUE_REG_9__1_, P3_INSTQUEUE_REG_9__0_, P3_INSTQUEUE_REG_8__7_,
    P3_INSTQUEUE_REG_8__6_, P3_INSTQUEUE_REG_8__5_, P3_INSTQUEUE_REG_8__4_,
    P3_INSTQUEUE_REG_8__3_, P3_INSTQUEUE_REG_8__2_, P3_INSTQUEUE_REG_8__1_,
    P3_INSTQUEUE_REG_8__0_, P3_INSTQUEUE_REG_7__7_, P3_INSTQUEUE_REG_7__6_,
    P3_INSTQUEUE_REG_7__5_, P3_INSTQUEUE_REG_7__4_, P3_INSTQUEUE_REG_7__3_,
    P3_INSTQUEUE_REG_7__2_, P3_INSTQUEUE_REG_7__1_, P3_INSTQUEUE_REG_7__0_,
    P3_INSTQUEUE_REG_6__7_, P3_INSTQUEUE_REG_6__6_, P3_INSTQUEUE_REG_6__5_,
    P3_INSTQUEUE_REG_6__4_, P3_INSTQUEUE_REG_6__3_, P3_INSTQUEUE_REG_6__2_,
    P3_INSTQUEUE_REG_6__1_, P3_INSTQUEUE_REG_6__0_, P3_INSTQUEUE_REG_5__7_,
    P3_INSTQUEUE_REG_5__6_, P3_INSTQUEUE_REG_5__5_, P3_INSTQUEUE_REG_5__4_,
    P3_INSTQUEUE_REG_5__3_, P3_INSTQUEUE_REG_5__2_, P3_INSTQUEUE_REG_5__1_,
    P3_INSTQUEUE_REG_5__0_, P3_INSTQUEUE_REG_4__7_, P3_INSTQUEUE_REG_4__6_,
    P3_INSTQUEUE_REG_4__5_, P3_INSTQUEUE_REG_4__4_, P3_INSTQUEUE_REG_4__3_,
    P3_INSTQUEUE_REG_4__2_, P3_INSTQUEUE_REG_4__1_, P3_INSTQUEUE_REG_4__0_,
    P3_INSTQUEUE_REG_3__7_, P3_INSTQUEUE_REG_3__6_, P3_INSTQUEUE_REG_3__5_,
    P3_INSTQUEUE_REG_3__4_, P3_INSTQUEUE_REG_3__3_, P3_INSTQUEUE_REG_3__2_,
    P3_INSTQUEUE_REG_3__1_, P3_INSTQUEUE_REG_3__0_, P3_INSTQUEUE_REG_2__7_,
    P3_INSTQUEUE_REG_2__6_, P3_INSTQUEUE_REG_2__5_, P3_INSTQUEUE_REG_2__4_,
    P3_INSTQUEUE_REG_2__3_, P3_INSTQUEUE_REG_2__2_, P3_INSTQUEUE_REG_2__1_,
    P3_INSTQUEUE_REG_2__0_, P3_INSTQUEUE_REG_1__7_, P3_INSTQUEUE_REG_1__6_,
    P3_INSTQUEUE_REG_1__5_, P3_INSTQUEUE_REG_1__4_, P3_INSTQUEUE_REG_1__3_,
    P3_INSTQUEUE_REG_1__2_, P3_INSTQUEUE_REG_1__1_, P3_INSTQUEUE_REG_1__0_,
    P3_INSTQUEUE_REG_0__7_, P3_INSTQUEUE_REG_0__6_, P3_INSTQUEUE_REG_0__5_,
    P3_INSTQUEUE_REG_0__4_, P3_INSTQUEUE_REG_0__3_, P3_INSTQUEUE_REG_0__2_,
    P3_INSTQUEUE_REG_0__1_, P3_INSTQUEUE_REG_0__0_,
    P3_INSTQUEUERD_ADDR_REG_4_, P3_INSTQUEUERD_ADDR_REG_3_,
    P3_INSTQUEUERD_ADDR_REG_2_, P3_INSTQUEUERD_ADDR_REG_1_,
    P3_INSTQUEUERD_ADDR_REG_0_, P3_INSTQUEUEWR_ADDR_REG_4_,
    P3_INSTQUEUEWR_ADDR_REG_3_, P3_INSTQUEUEWR_ADDR_REG_2_,
    P3_INSTQUEUEWR_ADDR_REG_1_, P3_INSTQUEUEWR_ADDR_REG_0_,
    P3_INSTADDRPOINTER_REG_0_, P3_INSTADDRPOINTER_REG_1_,
    P3_INSTADDRPOINTER_REG_2_, P3_INSTADDRPOINTER_REG_3_,
    P3_INSTADDRPOINTER_REG_4_, P3_INSTADDRPOINTER_REG_5_,
    P3_INSTADDRPOINTER_REG_6_, P3_INSTADDRPOINTER_REG_7_,
    P3_INSTADDRPOINTER_REG_8_, P3_INSTADDRPOINTER_REG_9_,
    P3_INSTADDRPOINTER_REG_10_, P3_INSTADDRPOINTER_REG_11_,
    P3_INSTADDRPOINTER_REG_12_, P3_INSTADDRPOINTER_REG_13_,
    P3_INSTADDRPOINTER_REG_14_, P3_INSTADDRPOINTER_REG_15_,
    P3_INSTADDRPOINTER_REG_16_, P3_INSTADDRPOINTER_REG_17_,
    P3_INSTADDRPOINTER_REG_18_, P3_INSTADDRPOINTER_REG_19_,
    P3_INSTADDRPOINTER_REG_20_, P3_INSTADDRPOINTER_REG_21_,
    P3_INSTADDRPOINTER_REG_22_, P3_INSTADDRPOINTER_REG_23_,
    P3_INSTADDRPOINTER_REG_24_, P3_INSTADDRPOINTER_REG_25_,
    P3_INSTADDRPOINTER_REG_26_, P3_INSTADDRPOINTER_REG_27_,
    P3_INSTADDRPOINTER_REG_28_, P3_INSTADDRPOINTER_REG_29_,
    P3_INSTADDRPOINTER_REG_30_, P3_INSTADDRPOINTER_REG_31_,
    P3_PHYADDRPOINTER_REG_0_, P3_PHYADDRPOINTER_REG_1_,
    P3_PHYADDRPOINTER_REG_2_, P3_PHYADDRPOINTER_REG_3_,
    P3_PHYADDRPOINTER_REG_4_, P3_PHYADDRPOINTER_REG_5_,
    P3_PHYADDRPOINTER_REG_6_, P3_PHYADDRPOINTER_REG_7_,
    P3_PHYADDRPOINTER_REG_8_, P3_PHYADDRPOINTER_REG_9_,
    P3_PHYADDRPOINTER_REG_10_, P3_PHYADDRPOINTER_REG_11_,
    P3_PHYADDRPOINTER_REG_12_, P3_PHYADDRPOINTER_REG_13_,
    P3_PHYADDRPOINTER_REG_14_, P3_PHYADDRPOINTER_REG_15_,
    P3_PHYADDRPOINTER_REG_16_, P3_PHYADDRPOINTER_REG_17_,
    P3_PHYADDRPOINTER_REG_18_, P3_PHYADDRPOINTER_REG_19_,
    P3_PHYADDRPOINTER_REG_20_, P3_PHYADDRPOINTER_REG_21_,
    P3_PHYADDRPOINTER_REG_22_, P3_PHYADDRPOINTER_REG_23_,
    P3_PHYADDRPOINTER_REG_24_, P3_PHYADDRPOINTER_REG_25_,
    P3_PHYADDRPOINTER_REG_26_, P3_PHYADDRPOINTER_REG_27_,
    P3_PHYADDRPOINTER_REG_28_, P3_PHYADDRPOINTER_REG_29_,
    P3_PHYADDRPOINTER_REG_30_, P3_PHYADDRPOINTER_REG_31_, P3_LWORD_REG_15_,
    P3_LWORD_REG_14_, P3_LWORD_REG_13_, P3_LWORD_REG_12_, P3_LWORD_REG_11_,
    P3_LWORD_REG_10_, P3_LWORD_REG_9_, P3_LWORD_REG_8_, P3_LWORD_REG_7_,
    P3_LWORD_REG_6_, P3_LWORD_REG_5_, P3_LWORD_REG_4_, P3_LWORD_REG_3_,
    P3_LWORD_REG_2_, P3_LWORD_REG_1_, P3_LWORD_REG_0_, P3_UWORD_REG_14_,
    P3_UWORD_REG_13_, P3_UWORD_REG_12_, P3_UWORD_REG_11_, P3_UWORD_REG_10_,
    P3_UWORD_REG_9_, P3_UWORD_REG_8_, P3_UWORD_REG_7_, P3_UWORD_REG_6_,
    P3_UWORD_REG_5_, P3_UWORD_REG_4_, P3_UWORD_REG_3_, P3_UWORD_REG_2_,
    P3_UWORD_REG_1_, P3_UWORD_REG_0_, P3_DATAO_REG_0_, P3_DATAO_REG_1_,
    P3_DATAO_REG_2_, P3_DATAO_REG_3_, P3_DATAO_REG_4_, P3_DATAO_REG_5_,
    P3_DATAO_REG_6_, P3_DATAO_REG_7_, P3_DATAO_REG_8_, P3_DATAO_REG_9_,
    P3_DATAO_REG_10_, P3_DATAO_REG_11_, P3_DATAO_REG_12_, P3_DATAO_REG_13_,
    P3_DATAO_REG_14_, P3_DATAO_REG_15_, P3_DATAO_REG_16_, P3_DATAO_REG_17_,
    P3_DATAO_REG_18_, P3_DATAO_REG_19_, P3_DATAO_REG_20_, P3_DATAO_REG_21_,
    P3_DATAO_REG_22_, P3_DATAO_REG_23_, P3_DATAO_REG_24_, P3_DATAO_REG_25_,
    P3_DATAO_REG_26_, P3_DATAO_REG_27_, P3_DATAO_REG_28_, P3_DATAO_REG_29_,
    P3_DATAO_REG_30_, P3_DATAO_REG_31_, P3_EAX_REG_0_, P3_EAX_REG_1_,
    P3_EAX_REG_2_, P3_EAX_REG_3_, P3_EAX_REG_4_, P3_EAX_REG_5_,
    P3_EAX_REG_6_, P3_EAX_REG_7_, P3_EAX_REG_8_, P3_EAX_REG_9_,
    P3_EAX_REG_10_, P3_EAX_REG_11_, P3_EAX_REG_12_, P3_EAX_REG_13_,
    P3_EAX_REG_14_, P3_EAX_REG_15_, P3_EAX_REG_16_, P3_EAX_REG_17_,
    P3_EAX_REG_18_, P3_EAX_REG_19_, P3_EAX_REG_20_, P3_EAX_REG_21_,
    P3_EAX_REG_22_, P3_EAX_REG_23_, P3_EAX_REG_24_, P3_EAX_REG_25_,
    P3_EAX_REG_26_, P3_EAX_REG_27_, P3_EAX_REG_28_, P3_EAX_REG_29_,
    P3_EAX_REG_30_, P3_EAX_REG_31_, P3_EBX_REG_0_, P3_EBX_REG_1_,
    P3_EBX_REG_2_, P3_EBX_REG_3_, P3_EBX_REG_4_, P3_EBX_REG_5_,
    P3_EBX_REG_6_, P3_EBX_REG_7_, P3_EBX_REG_8_, P3_EBX_REG_9_,
    P3_EBX_REG_10_, P3_EBX_REG_11_, P3_EBX_REG_12_, P3_EBX_REG_13_,
    P3_EBX_REG_14_, P3_EBX_REG_15_, P3_EBX_REG_16_, P3_EBX_REG_17_,
    P3_EBX_REG_18_, P3_EBX_REG_19_, P3_EBX_REG_20_, P3_EBX_REG_21_,
    P3_EBX_REG_22_, P3_EBX_REG_23_, P3_EBX_REG_24_, P3_EBX_REG_25_,
    P3_EBX_REG_26_, P3_EBX_REG_27_, P3_EBX_REG_28_, P3_EBX_REG_29_,
    P3_EBX_REG_30_, P3_EBX_REG_31_, P3_REIP_REG_0_, P3_REIP_REG_1_,
    P3_REIP_REG_2_, P3_REIP_REG_3_, P3_REIP_REG_4_, P3_REIP_REG_5_,
    P3_REIP_REG_6_, P3_REIP_REG_7_, P3_REIP_REG_8_, P3_REIP_REG_9_,
    P3_REIP_REG_10_, P3_REIP_REG_11_, P3_REIP_REG_12_, P3_REIP_REG_13_,
    P3_REIP_REG_14_, P3_REIP_REG_15_, P3_REIP_REG_16_, P3_REIP_REG_17_,
    P3_REIP_REG_18_, P3_REIP_REG_19_, P3_REIP_REG_20_, P3_REIP_REG_21_,
    P3_REIP_REG_22_, P3_REIP_REG_23_, P3_REIP_REG_24_, P3_REIP_REG_25_,
    P3_REIP_REG_26_, P3_REIP_REG_27_, P3_REIP_REG_28_, P3_REIP_REG_29_,
    P3_REIP_REG_30_, P3_REIP_REG_31_, P3_BYTEENABLE_REG_3_,
    P3_BYTEENABLE_REG_2_, P3_BYTEENABLE_REG_1_, P3_BYTEENABLE_REG_0_,
    P3_W_R_N_REG, P3_FLUSH_REG, P3_MORE_REG, P3_STATEBS16_REG,
    P3_REQUESTPENDING_REG, P3_D_C_N_REG, P3_M_IO_N_REG, P3_CODEFETCH_REG,
    P3_ADS_N_REG, P3_READREQUEST_REG, P3_MEMORYFETCH_REG, P2_BE_N_REG_3_,
    P2_BE_N_REG_2_, P2_BE_N_REG_1_, P2_BE_N_REG_0_, P2_ADDRESS_REG_29_,
    P2_ADDRESS_REG_28_, P2_ADDRESS_REG_27_, P2_ADDRESS_REG_26_,
    P2_ADDRESS_REG_25_, P2_ADDRESS_REG_24_, P2_ADDRESS_REG_23_,
    P2_ADDRESS_REG_22_, P2_ADDRESS_REG_21_, P2_ADDRESS_REG_20_,
    P2_ADDRESS_REG_19_, P2_ADDRESS_REG_18_, P2_ADDRESS_REG_17_,
    P2_ADDRESS_REG_16_, P2_ADDRESS_REG_15_, P2_ADDRESS_REG_14_,
    P2_ADDRESS_REG_13_, P2_ADDRESS_REG_12_, P2_ADDRESS_REG_11_,
    P2_ADDRESS_REG_10_, P2_ADDRESS_REG_9_, P2_ADDRESS_REG_8_,
    P2_ADDRESS_REG_7_, P2_ADDRESS_REG_6_, P2_ADDRESS_REG_5_,
    P2_ADDRESS_REG_4_, P2_ADDRESS_REG_3_, P2_ADDRESS_REG_2_,
    P2_ADDRESS_REG_1_, P2_ADDRESS_REG_0_, P2_STATE_REG_2_, P2_STATE_REG_1_,
    P2_STATE_REG_0_, P2_DATAWIDTH_REG_0_, P2_DATAWIDTH_REG_1_,
    P2_DATAWIDTH_REG_2_, P2_DATAWIDTH_REG_3_, P2_DATAWIDTH_REG_4_,
    P2_DATAWIDTH_REG_5_, P2_DATAWIDTH_REG_6_, P2_DATAWIDTH_REG_7_,
    P2_DATAWIDTH_REG_8_, P2_DATAWIDTH_REG_9_, P2_DATAWIDTH_REG_10_,
    P2_DATAWIDTH_REG_11_, P2_DATAWIDTH_REG_12_, P2_DATAWIDTH_REG_13_,
    P2_DATAWIDTH_REG_14_, P2_DATAWIDTH_REG_15_, P2_DATAWIDTH_REG_16_,
    P2_DATAWIDTH_REG_17_, P2_DATAWIDTH_REG_18_, P2_DATAWIDTH_REG_19_,
    P2_DATAWIDTH_REG_20_, P2_DATAWIDTH_REG_21_, P2_DATAWIDTH_REG_22_,
    P2_DATAWIDTH_REG_23_, P2_DATAWIDTH_REG_24_, P2_DATAWIDTH_REG_25_,
    P2_DATAWIDTH_REG_26_, P2_DATAWIDTH_REG_27_, P2_DATAWIDTH_REG_28_,
    P2_DATAWIDTH_REG_29_, P2_DATAWIDTH_REG_30_, P2_DATAWIDTH_REG_31_,
    P2_STATE2_REG_3_, P2_STATE2_REG_2_, P2_STATE2_REG_1_, P2_STATE2_REG_0_,
    P2_INSTQUEUE_REG_15__7_, P2_INSTQUEUE_REG_15__6_,
    P2_INSTQUEUE_REG_15__5_, P2_INSTQUEUE_REG_15__4_,
    P2_INSTQUEUE_REG_15__3_, P2_INSTQUEUE_REG_15__2_,
    P2_INSTQUEUE_REG_15__1_, P2_INSTQUEUE_REG_15__0_,
    P2_INSTQUEUE_REG_14__7_, P2_INSTQUEUE_REG_14__6_,
    P2_INSTQUEUE_REG_14__5_, P2_INSTQUEUE_REG_14__4_,
    P2_INSTQUEUE_REG_14__3_, P2_INSTQUEUE_REG_14__2_,
    P2_INSTQUEUE_REG_14__1_, P2_INSTQUEUE_REG_14__0_,
    P2_INSTQUEUE_REG_13__7_, P2_INSTQUEUE_REG_13__6_,
    P2_INSTQUEUE_REG_13__5_, P2_INSTQUEUE_REG_13__4_,
    P2_INSTQUEUE_REG_13__3_, P2_INSTQUEUE_REG_13__2_,
    P2_INSTQUEUE_REG_13__1_, P2_INSTQUEUE_REG_13__0_,
    P2_INSTQUEUE_REG_12__7_, P2_INSTQUEUE_REG_12__6_,
    P2_INSTQUEUE_REG_12__5_, P2_INSTQUEUE_REG_12__4_,
    P2_INSTQUEUE_REG_12__3_, P2_INSTQUEUE_REG_12__2_,
    P2_INSTQUEUE_REG_12__1_, P2_INSTQUEUE_REG_12__0_,
    P2_INSTQUEUE_REG_11__7_, P2_INSTQUEUE_REG_11__6_,
    P2_INSTQUEUE_REG_11__5_, P2_INSTQUEUE_REG_11__4_,
    P2_INSTQUEUE_REG_11__3_, P2_INSTQUEUE_REG_11__2_,
    P2_INSTQUEUE_REG_11__1_, P2_INSTQUEUE_REG_11__0_,
    P2_INSTQUEUE_REG_10__7_, P2_INSTQUEUE_REG_10__6_,
    P2_INSTQUEUE_REG_10__5_, P2_INSTQUEUE_REG_10__4_,
    P2_INSTQUEUE_REG_10__3_, P2_INSTQUEUE_REG_10__2_,
    P2_INSTQUEUE_REG_10__1_, P2_INSTQUEUE_REG_10__0_,
    P2_INSTQUEUE_REG_9__7_, P2_INSTQUEUE_REG_9__6_, P2_INSTQUEUE_REG_9__5_,
    P2_INSTQUEUE_REG_9__4_, P2_INSTQUEUE_REG_9__3_, P2_INSTQUEUE_REG_9__2_,
    P2_INSTQUEUE_REG_9__1_, P2_INSTQUEUE_REG_9__0_, P2_INSTQUEUE_REG_8__7_,
    P2_INSTQUEUE_REG_8__6_, P2_INSTQUEUE_REG_8__5_, P2_INSTQUEUE_REG_8__4_,
    P2_INSTQUEUE_REG_8__3_, P2_INSTQUEUE_REG_8__2_, P2_INSTQUEUE_REG_8__1_,
    P2_INSTQUEUE_REG_8__0_, P2_INSTQUEUE_REG_7__7_, P2_INSTQUEUE_REG_7__6_,
    P2_INSTQUEUE_REG_7__5_, P2_INSTQUEUE_REG_7__4_, P2_INSTQUEUE_REG_7__3_,
    P2_INSTQUEUE_REG_7__2_, P2_INSTQUEUE_REG_7__1_, P2_INSTQUEUE_REG_7__0_,
    P2_INSTQUEUE_REG_6__7_, P2_INSTQUEUE_REG_6__6_, P2_INSTQUEUE_REG_6__5_,
    P2_INSTQUEUE_REG_6__4_, P2_INSTQUEUE_REG_6__3_, P2_INSTQUEUE_REG_6__2_,
    P2_INSTQUEUE_REG_6__1_, P2_INSTQUEUE_REG_6__0_, P2_INSTQUEUE_REG_5__7_,
    P2_INSTQUEUE_REG_5__6_, P2_INSTQUEUE_REG_5__5_, P2_INSTQUEUE_REG_5__4_,
    P2_INSTQUEUE_REG_5__3_, P2_INSTQUEUE_REG_5__2_, P2_INSTQUEUE_REG_5__1_,
    P2_INSTQUEUE_REG_5__0_, P2_INSTQUEUE_REG_4__7_, P2_INSTQUEUE_REG_4__6_,
    P2_INSTQUEUE_REG_4__5_, P2_INSTQUEUE_REG_4__4_, P2_INSTQUEUE_REG_4__3_,
    P2_INSTQUEUE_REG_4__2_, P2_INSTQUEUE_REG_4__1_, P2_INSTQUEUE_REG_4__0_,
    P2_INSTQUEUE_REG_3__7_, P2_INSTQUEUE_REG_3__6_, P2_INSTQUEUE_REG_3__5_,
    P2_INSTQUEUE_REG_3__4_, P2_INSTQUEUE_REG_3__3_, P2_INSTQUEUE_REG_3__2_,
    P2_INSTQUEUE_REG_3__1_, P2_INSTQUEUE_REG_3__0_, P2_INSTQUEUE_REG_2__7_,
    P2_INSTQUEUE_REG_2__6_, P2_INSTQUEUE_REG_2__5_, P2_INSTQUEUE_REG_2__4_,
    P2_INSTQUEUE_REG_2__3_, P2_INSTQUEUE_REG_2__2_, P2_INSTQUEUE_REG_2__1_,
    P2_INSTQUEUE_REG_2__0_, P2_INSTQUEUE_REG_1__7_, P2_INSTQUEUE_REG_1__6_,
    P2_INSTQUEUE_REG_1__5_, P2_INSTQUEUE_REG_1__4_, P2_INSTQUEUE_REG_1__3_,
    P2_INSTQUEUE_REG_1__2_, P2_INSTQUEUE_REG_1__1_, P2_INSTQUEUE_REG_1__0_,
    P2_INSTQUEUE_REG_0__7_, P2_INSTQUEUE_REG_0__6_, P2_INSTQUEUE_REG_0__5_,
    P2_INSTQUEUE_REG_0__4_, P2_INSTQUEUE_REG_0__3_, P2_INSTQUEUE_REG_0__2_,
    P2_INSTQUEUE_REG_0__1_, P2_INSTQUEUE_REG_0__0_,
    P2_INSTQUEUERD_ADDR_REG_4_, P2_INSTQUEUERD_ADDR_REG_3_,
    P2_INSTQUEUERD_ADDR_REG_2_, P2_INSTQUEUERD_ADDR_REG_1_,
    P2_INSTQUEUERD_ADDR_REG_0_, P2_INSTQUEUEWR_ADDR_REG_4_,
    P2_INSTQUEUEWR_ADDR_REG_3_, P2_INSTQUEUEWR_ADDR_REG_2_,
    P2_INSTQUEUEWR_ADDR_REG_1_, P2_INSTQUEUEWR_ADDR_REG_0_,
    P2_INSTADDRPOINTER_REG_0_, P2_INSTADDRPOINTER_REG_1_,
    P2_INSTADDRPOINTER_REG_2_, P2_INSTADDRPOINTER_REG_3_,
    P2_INSTADDRPOINTER_REG_4_, P2_INSTADDRPOINTER_REG_5_,
    P2_INSTADDRPOINTER_REG_6_, P2_INSTADDRPOINTER_REG_7_,
    P2_INSTADDRPOINTER_REG_8_, P2_INSTADDRPOINTER_REG_9_,
    P2_INSTADDRPOINTER_REG_10_, P2_INSTADDRPOINTER_REG_11_,
    P2_INSTADDRPOINTER_REG_12_, P2_INSTADDRPOINTER_REG_13_,
    P2_INSTADDRPOINTER_REG_14_, P2_INSTADDRPOINTER_REG_15_,
    P2_INSTADDRPOINTER_REG_16_, P2_INSTADDRPOINTER_REG_17_,
    P2_INSTADDRPOINTER_REG_18_, P2_INSTADDRPOINTER_REG_19_,
    P2_INSTADDRPOINTER_REG_20_, P2_INSTADDRPOINTER_REG_21_,
    P2_INSTADDRPOINTER_REG_22_, P2_INSTADDRPOINTER_REG_23_,
    P2_INSTADDRPOINTER_REG_24_, P2_INSTADDRPOINTER_REG_25_,
    P2_INSTADDRPOINTER_REG_26_, P2_INSTADDRPOINTER_REG_27_,
    P2_INSTADDRPOINTER_REG_28_, P2_INSTADDRPOINTER_REG_29_,
    P2_INSTADDRPOINTER_REG_30_, P2_INSTADDRPOINTER_REG_31_,
    P2_PHYADDRPOINTER_REG_0_, P2_PHYADDRPOINTER_REG_1_,
    P2_PHYADDRPOINTER_REG_2_, P2_PHYADDRPOINTER_REG_3_,
    P2_PHYADDRPOINTER_REG_4_, P2_PHYADDRPOINTER_REG_5_,
    P2_PHYADDRPOINTER_REG_6_, P2_PHYADDRPOINTER_REG_7_,
    P2_PHYADDRPOINTER_REG_8_, P2_PHYADDRPOINTER_REG_9_,
    P2_PHYADDRPOINTER_REG_10_, P2_PHYADDRPOINTER_REG_11_,
    P2_PHYADDRPOINTER_REG_12_, P2_PHYADDRPOINTER_REG_13_,
    P2_PHYADDRPOINTER_REG_14_, P2_PHYADDRPOINTER_REG_15_,
    P2_PHYADDRPOINTER_REG_16_, P2_PHYADDRPOINTER_REG_17_,
    P2_PHYADDRPOINTER_REG_18_, P2_PHYADDRPOINTER_REG_19_,
    P2_PHYADDRPOINTER_REG_20_, P2_PHYADDRPOINTER_REG_21_,
    P2_PHYADDRPOINTER_REG_22_, P2_PHYADDRPOINTER_REG_23_,
    P2_PHYADDRPOINTER_REG_24_, P2_PHYADDRPOINTER_REG_25_,
    P2_PHYADDRPOINTER_REG_26_, P2_PHYADDRPOINTER_REG_27_,
    P2_PHYADDRPOINTER_REG_28_, P2_PHYADDRPOINTER_REG_29_,
    P2_PHYADDRPOINTER_REG_30_, P2_PHYADDRPOINTER_REG_31_, P2_LWORD_REG_15_,
    P2_LWORD_REG_14_, P2_LWORD_REG_13_, P2_LWORD_REG_12_, P2_LWORD_REG_11_,
    P2_LWORD_REG_10_, P2_LWORD_REG_9_, P2_LWORD_REG_8_, P2_LWORD_REG_7_,
    P2_LWORD_REG_6_, P2_LWORD_REG_5_, P2_LWORD_REG_4_, P2_LWORD_REG_3_,
    P2_LWORD_REG_2_, P2_LWORD_REG_1_, P2_LWORD_REG_0_, P2_UWORD_REG_14_,
    P2_UWORD_REG_13_, P2_UWORD_REG_12_, P2_UWORD_REG_11_, P2_UWORD_REG_10_,
    P2_UWORD_REG_9_, P2_UWORD_REG_8_, P2_UWORD_REG_7_, P2_UWORD_REG_6_,
    P2_UWORD_REG_5_, P2_UWORD_REG_4_, P2_UWORD_REG_3_, P2_UWORD_REG_2_,
    P2_UWORD_REG_1_, P2_UWORD_REG_0_, P2_DATAO_REG_0_, P2_DATAO_REG_1_,
    P2_DATAO_REG_2_, P2_DATAO_REG_3_, P2_DATAO_REG_4_, P2_DATAO_REG_5_,
    P2_DATAO_REG_6_, P2_DATAO_REG_7_, P2_DATAO_REG_8_, P2_DATAO_REG_9_,
    P2_DATAO_REG_10_, P2_DATAO_REG_11_, P2_DATAO_REG_12_, P2_DATAO_REG_13_,
    P2_DATAO_REG_14_, P2_DATAO_REG_15_, P2_DATAO_REG_16_, P2_DATAO_REG_17_,
    P2_DATAO_REG_18_, P2_DATAO_REG_19_, P2_DATAO_REG_20_, P2_DATAO_REG_21_,
    P2_DATAO_REG_22_, P2_DATAO_REG_23_, P2_DATAO_REG_24_, P2_DATAO_REG_25_,
    P2_DATAO_REG_26_, P2_DATAO_REG_27_, P2_DATAO_REG_28_, P2_DATAO_REG_29_,
    P2_DATAO_REG_30_, P2_DATAO_REG_31_, P2_EAX_REG_0_, P2_EAX_REG_1_,
    P2_EAX_REG_2_, P2_EAX_REG_3_, P2_EAX_REG_4_, P2_EAX_REG_5_,
    P2_EAX_REG_6_, P2_EAX_REG_7_, P2_EAX_REG_8_, P2_EAX_REG_9_,
    P2_EAX_REG_10_, P2_EAX_REG_11_, P2_EAX_REG_12_, P2_EAX_REG_13_,
    P2_EAX_REG_14_, P2_EAX_REG_15_, P2_EAX_REG_16_, P2_EAX_REG_17_,
    P2_EAX_REG_18_, P2_EAX_REG_19_, P2_EAX_REG_20_, P2_EAX_REG_21_,
    P2_EAX_REG_22_, P2_EAX_REG_23_, P2_EAX_REG_24_, P2_EAX_REG_25_,
    P2_EAX_REG_26_, P2_EAX_REG_27_, P2_EAX_REG_28_, P2_EAX_REG_29_,
    P2_EAX_REG_30_, P2_EAX_REG_31_, P2_EBX_REG_0_, P2_EBX_REG_1_,
    P2_EBX_REG_2_, P2_EBX_REG_3_, P2_EBX_REG_4_, P2_EBX_REG_5_,
    P2_EBX_REG_6_, P2_EBX_REG_7_, P2_EBX_REG_8_, P2_EBX_REG_9_,
    P2_EBX_REG_10_, P2_EBX_REG_11_, P2_EBX_REG_12_, P2_EBX_REG_13_,
    P2_EBX_REG_14_, P2_EBX_REG_15_, P2_EBX_REG_16_, P2_EBX_REG_17_,
    P2_EBX_REG_18_, P2_EBX_REG_19_, P2_EBX_REG_20_, P2_EBX_REG_21_,
    P2_EBX_REG_22_, P2_EBX_REG_23_, P2_EBX_REG_24_, P2_EBX_REG_25_,
    P2_EBX_REG_26_, P2_EBX_REG_27_, P2_EBX_REG_28_, P2_EBX_REG_29_,
    P2_EBX_REG_30_, P2_EBX_REG_31_, P2_REIP_REG_0_, P2_REIP_REG_1_,
    P2_REIP_REG_2_, P2_REIP_REG_3_, P2_REIP_REG_4_, P2_REIP_REG_5_,
    P2_REIP_REG_6_, P2_REIP_REG_7_, P2_REIP_REG_8_, P2_REIP_REG_9_,
    P2_REIP_REG_10_, P2_REIP_REG_11_, P2_REIP_REG_12_, P2_REIP_REG_13_,
    P2_REIP_REG_14_, P2_REIP_REG_15_, P2_REIP_REG_16_, P2_REIP_REG_17_,
    P2_REIP_REG_18_, P2_REIP_REG_19_, P2_REIP_REG_20_, P2_REIP_REG_21_,
    P2_REIP_REG_22_, P2_REIP_REG_23_, P2_REIP_REG_24_, P2_REIP_REG_25_,
    P2_REIP_REG_26_, P2_REIP_REG_27_, P2_REIP_REG_28_, P2_REIP_REG_29_,
    P2_REIP_REG_30_, P2_REIP_REG_31_, P2_BYTEENABLE_REG_3_,
    P2_BYTEENABLE_REG_2_, P2_BYTEENABLE_REG_1_, P2_BYTEENABLE_REG_0_,
    P2_W_R_N_REG, P2_FLUSH_REG, P2_MORE_REG, P2_STATEBS16_REG,
    P2_REQUESTPENDING_REG, P2_D_C_N_REG, P2_M_IO_N_REG, P2_CODEFETCH_REG,
    P2_ADS_N_REG, P2_READREQUEST_REG, P2_MEMORYFETCH_REG, P1_BE_N_REG_3_,
    P1_BE_N_REG_2_, P1_BE_N_REG_1_, P1_BE_N_REG_0_, P1_ADDRESS_REG_29_,
    P1_ADDRESS_REG_28_, P1_ADDRESS_REG_27_, P1_ADDRESS_REG_26_,
    P1_ADDRESS_REG_25_, P1_ADDRESS_REG_24_, P1_ADDRESS_REG_23_,
    P1_ADDRESS_REG_22_, P1_ADDRESS_REG_21_, P1_ADDRESS_REG_20_,
    P1_ADDRESS_REG_19_, P1_ADDRESS_REG_18_, P1_ADDRESS_REG_17_,
    P1_ADDRESS_REG_16_, P1_ADDRESS_REG_15_, P1_ADDRESS_REG_14_,
    P1_ADDRESS_REG_13_, P1_ADDRESS_REG_12_, P1_ADDRESS_REG_11_,
    P1_ADDRESS_REG_10_, P1_ADDRESS_REG_9_, P1_ADDRESS_REG_8_,
    P1_ADDRESS_REG_7_, P1_ADDRESS_REG_6_, P1_ADDRESS_REG_5_,
    P1_ADDRESS_REG_4_, P1_ADDRESS_REG_3_, P1_ADDRESS_REG_2_,
    P1_ADDRESS_REG_1_, P1_ADDRESS_REG_0_, P1_STATE_REG_2_, P1_STATE_REG_1_,
    P1_STATE_REG_0_, P1_DATAWIDTH_REG_0_, P1_DATAWIDTH_REG_1_,
    P1_DATAWIDTH_REG_2_, P1_DATAWIDTH_REG_3_, P1_DATAWIDTH_REG_4_,
    P1_DATAWIDTH_REG_5_, P1_DATAWIDTH_REG_6_, P1_DATAWIDTH_REG_7_,
    P1_DATAWIDTH_REG_8_, P1_DATAWIDTH_REG_9_, P1_DATAWIDTH_REG_10_,
    P1_DATAWIDTH_REG_11_, P1_DATAWIDTH_REG_12_, P1_DATAWIDTH_REG_13_,
    P1_DATAWIDTH_REG_14_, P1_DATAWIDTH_REG_15_, P1_DATAWIDTH_REG_16_,
    P1_DATAWIDTH_REG_17_, P1_DATAWIDTH_REG_18_, P1_DATAWIDTH_REG_19_,
    P1_DATAWIDTH_REG_20_, P1_DATAWIDTH_REG_21_, P1_DATAWIDTH_REG_22_,
    P1_DATAWIDTH_REG_23_, P1_DATAWIDTH_REG_24_, P1_DATAWIDTH_REG_25_,
    P1_DATAWIDTH_REG_26_, P1_DATAWIDTH_REG_27_, P1_DATAWIDTH_REG_28_,
    P1_DATAWIDTH_REG_29_, P1_DATAWIDTH_REG_30_, P1_DATAWIDTH_REG_31_,
    P1_STATE2_REG_3_, P1_STATE2_REG_2_, P1_STATE2_REG_1_, P1_STATE2_REG_0_,
    P1_INSTQUEUE_REG_15__7_, P1_INSTQUEUE_REG_15__6_,
    P1_INSTQUEUE_REG_15__5_, P1_INSTQUEUE_REG_15__4_,
    P1_INSTQUEUE_REG_15__3_, P1_INSTQUEUE_REG_15__2_,
    P1_INSTQUEUE_REG_15__1_, P1_INSTQUEUE_REG_15__0_,
    P1_INSTQUEUE_REG_14__7_, P1_INSTQUEUE_REG_14__6_,
    P1_INSTQUEUE_REG_14__5_, P1_INSTQUEUE_REG_14__4_,
    P1_INSTQUEUE_REG_14__3_, P1_INSTQUEUE_REG_14__2_,
    P1_INSTQUEUE_REG_14__1_, P1_INSTQUEUE_REG_14__0_,
    P1_INSTQUEUE_REG_13__7_, P1_INSTQUEUE_REG_13__6_,
    P1_INSTQUEUE_REG_13__5_, P1_INSTQUEUE_REG_13__4_,
    P1_INSTQUEUE_REG_13__3_, P1_INSTQUEUE_REG_13__2_,
    P1_INSTQUEUE_REG_13__1_, P1_INSTQUEUE_REG_13__0_,
    P1_INSTQUEUE_REG_12__7_, P1_INSTQUEUE_REG_12__6_,
    P1_INSTQUEUE_REG_12__5_, P1_INSTQUEUE_REG_12__4_,
    P1_INSTQUEUE_REG_12__3_, P1_INSTQUEUE_REG_12__2_,
    P1_INSTQUEUE_REG_12__1_, P1_INSTQUEUE_REG_12__0_,
    P1_INSTQUEUE_REG_11__7_, P1_INSTQUEUE_REG_11__6_,
    P1_INSTQUEUE_REG_11__5_, P1_INSTQUEUE_REG_11__4_,
    P1_INSTQUEUE_REG_11__3_, P1_INSTQUEUE_REG_11__2_,
    P1_INSTQUEUE_REG_11__1_, P1_INSTQUEUE_REG_11__0_,
    P1_INSTQUEUE_REG_10__7_, P1_INSTQUEUE_REG_10__6_,
    P1_INSTQUEUE_REG_10__5_, P1_INSTQUEUE_REG_10__4_,
    P1_INSTQUEUE_REG_10__3_, P1_INSTQUEUE_REG_10__2_,
    P1_INSTQUEUE_REG_10__1_, P1_INSTQUEUE_REG_10__0_,
    P1_INSTQUEUE_REG_9__7_, P1_INSTQUEUE_REG_9__6_, P1_INSTQUEUE_REG_9__5_,
    P1_INSTQUEUE_REG_9__4_, P1_INSTQUEUE_REG_9__3_, P1_INSTQUEUE_REG_9__2_,
    P1_INSTQUEUE_REG_9__1_, P1_INSTQUEUE_REG_9__0_, P1_INSTQUEUE_REG_8__7_,
    P1_INSTQUEUE_REG_8__6_, P1_INSTQUEUE_REG_8__5_, P1_INSTQUEUE_REG_8__4_,
    P1_INSTQUEUE_REG_8__3_, P1_INSTQUEUE_REG_8__2_, P1_INSTQUEUE_REG_8__1_,
    P1_INSTQUEUE_REG_8__0_, P1_INSTQUEUE_REG_7__7_, P1_INSTQUEUE_REG_7__6_,
    P1_INSTQUEUE_REG_7__5_, P1_INSTQUEUE_REG_7__4_, P1_INSTQUEUE_REG_7__3_,
    P1_INSTQUEUE_REG_7__2_, P1_INSTQUEUE_REG_7__1_, P1_INSTQUEUE_REG_7__0_,
    P1_INSTQUEUE_REG_6__7_, P1_INSTQUEUE_REG_6__6_, P1_INSTQUEUE_REG_6__5_,
    P1_INSTQUEUE_REG_6__4_, P1_INSTQUEUE_REG_6__3_, P1_INSTQUEUE_REG_6__2_,
    P1_INSTQUEUE_REG_6__1_, P1_INSTQUEUE_REG_6__0_, P1_INSTQUEUE_REG_5__7_,
    P1_INSTQUEUE_REG_5__6_, P1_INSTQUEUE_REG_5__5_, P1_INSTQUEUE_REG_5__4_,
    P1_INSTQUEUE_REG_5__3_, P1_INSTQUEUE_REG_5__2_, P1_INSTQUEUE_REG_5__1_,
    P1_INSTQUEUE_REG_5__0_, P1_INSTQUEUE_REG_4__7_, P1_INSTQUEUE_REG_4__6_,
    P1_INSTQUEUE_REG_4__5_, P1_INSTQUEUE_REG_4__4_, P1_INSTQUEUE_REG_4__3_,
    P1_INSTQUEUE_REG_4__2_, P1_INSTQUEUE_REG_4__1_, P1_INSTQUEUE_REG_4__0_,
    P1_INSTQUEUE_REG_3__7_, P1_INSTQUEUE_REG_3__6_, P1_INSTQUEUE_REG_3__5_,
    P1_INSTQUEUE_REG_3__4_, P1_INSTQUEUE_REG_3__3_, P1_INSTQUEUE_REG_3__2_,
    P1_INSTQUEUE_REG_3__1_, P1_INSTQUEUE_REG_3__0_, P1_INSTQUEUE_REG_2__7_,
    P1_INSTQUEUE_REG_2__6_, P1_INSTQUEUE_REG_2__5_, P1_INSTQUEUE_REG_2__4_,
    P1_INSTQUEUE_REG_2__3_, P1_INSTQUEUE_REG_2__2_, P1_INSTQUEUE_REG_2__1_,
    P1_INSTQUEUE_REG_2__0_, P1_INSTQUEUE_REG_1__7_, P1_INSTQUEUE_REG_1__6_,
    P1_INSTQUEUE_REG_1__5_, P1_INSTQUEUE_REG_1__4_, P1_INSTQUEUE_REG_1__3_,
    P1_INSTQUEUE_REG_1__2_, P1_INSTQUEUE_REG_1__1_, P1_INSTQUEUE_REG_1__0_,
    P1_INSTQUEUE_REG_0__7_, P1_INSTQUEUE_REG_0__6_, P1_INSTQUEUE_REG_0__5_,
    P1_INSTQUEUE_REG_0__4_, P1_INSTQUEUE_REG_0__3_, P1_INSTQUEUE_REG_0__2_,
    P1_INSTQUEUE_REG_0__1_, P1_INSTQUEUE_REG_0__0_,
    P1_INSTQUEUERD_ADDR_REG_4_, P1_INSTQUEUERD_ADDR_REG_3_,
    P1_INSTQUEUERD_ADDR_REG_2_, P1_INSTQUEUERD_ADDR_REG_1_,
    P1_INSTQUEUERD_ADDR_REG_0_, P1_INSTQUEUEWR_ADDR_REG_4_,
    P1_INSTQUEUEWR_ADDR_REG_3_, P1_INSTQUEUEWR_ADDR_REG_2_,
    P1_INSTQUEUEWR_ADDR_REG_1_, P1_INSTQUEUEWR_ADDR_REG_0_,
    P1_INSTADDRPOINTER_REG_0_, P1_INSTADDRPOINTER_REG_1_,
    P1_INSTADDRPOINTER_REG_2_, P1_INSTADDRPOINTER_REG_3_,
    P1_INSTADDRPOINTER_REG_4_, P1_INSTADDRPOINTER_REG_5_,
    P1_INSTADDRPOINTER_REG_6_, P1_INSTADDRPOINTER_REG_7_,
    P1_INSTADDRPOINTER_REG_8_, P1_INSTADDRPOINTER_REG_9_,
    P1_INSTADDRPOINTER_REG_10_, P1_INSTADDRPOINTER_REG_11_,
    P1_INSTADDRPOINTER_REG_12_, P1_INSTADDRPOINTER_REG_13_,
    P1_INSTADDRPOINTER_REG_14_, P1_INSTADDRPOINTER_REG_15_,
    P1_INSTADDRPOINTER_REG_16_, P1_INSTADDRPOINTER_REG_17_,
    P1_INSTADDRPOINTER_REG_18_, P1_INSTADDRPOINTER_REG_19_,
    P1_INSTADDRPOINTER_REG_20_, P1_INSTADDRPOINTER_REG_21_,
    P1_INSTADDRPOINTER_REG_22_, P1_INSTADDRPOINTER_REG_23_,
    P1_INSTADDRPOINTER_REG_24_, P1_INSTADDRPOINTER_REG_25_,
    P1_INSTADDRPOINTER_REG_26_, P1_INSTADDRPOINTER_REG_27_,
    P1_INSTADDRPOINTER_REG_28_, P1_INSTADDRPOINTER_REG_29_,
    P1_INSTADDRPOINTER_REG_30_, P1_INSTADDRPOINTER_REG_31_,
    P1_PHYADDRPOINTER_REG_0_, P1_PHYADDRPOINTER_REG_1_,
    P1_PHYADDRPOINTER_REG_2_, P1_PHYADDRPOINTER_REG_3_,
    P1_PHYADDRPOINTER_REG_4_, P1_PHYADDRPOINTER_REG_5_,
    P1_PHYADDRPOINTER_REG_6_, P1_PHYADDRPOINTER_REG_7_,
    P1_PHYADDRPOINTER_REG_8_, P1_PHYADDRPOINTER_REG_9_,
    P1_PHYADDRPOINTER_REG_10_, P1_PHYADDRPOINTER_REG_11_,
    P1_PHYADDRPOINTER_REG_12_, P1_PHYADDRPOINTER_REG_13_,
    P1_PHYADDRPOINTER_REG_14_, P1_PHYADDRPOINTER_REG_15_,
    P1_PHYADDRPOINTER_REG_16_, P1_PHYADDRPOINTER_REG_17_,
    P1_PHYADDRPOINTER_REG_18_, P1_PHYADDRPOINTER_REG_19_,
    P1_PHYADDRPOINTER_REG_20_, P1_PHYADDRPOINTER_REG_21_,
    P1_PHYADDRPOINTER_REG_22_, P1_PHYADDRPOINTER_REG_23_,
    P1_PHYADDRPOINTER_REG_24_, P1_PHYADDRPOINTER_REG_25_,
    P1_PHYADDRPOINTER_REG_26_, P1_PHYADDRPOINTER_REG_27_,
    P1_PHYADDRPOINTER_REG_28_, P1_PHYADDRPOINTER_REG_29_,
    P1_PHYADDRPOINTER_REG_30_, P1_PHYADDRPOINTER_REG_31_, P1_LWORD_REG_15_,
    P1_LWORD_REG_14_, P1_LWORD_REG_13_, P1_LWORD_REG_12_, P1_LWORD_REG_11_,
    P1_LWORD_REG_10_, P1_LWORD_REG_9_, P1_LWORD_REG_8_, P1_LWORD_REG_7_,
    P1_LWORD_REG_6_, P1_LWORD_REG_5_, P1_LWORD_REG_4_, P1_LWORD_REG_3_,
    P1_LWORD_REG_2_, P1_LWORD_REG_1_, P1_LWORD_REG_0_, P1_UWORD_REG_14_,
    P1_UWORD_REG_13_, P1_UWORD_REG_12_, P1_UWORD_REG_11_, P1_UWORD_REG_10_,
    P1_UWORD_REG_9_, P1_UWORD_REG_8_, P1_UWORD_REG_7_, P1_UWORD_REG_6_,
    P1_UWORD_REG_5_, P1_UWORD_REG_4_, P1_UWORD_REG_3_, P1_UWORD_REG_2_,
    P1_UWORD_REG_1_, P1_UWORD_REG_0_, P1_DATAO_REG_0_, P1_DATAO_REG_1_,
    P1_DATAO_REG_2_, P1_DATAO_REG_3_, P1_DATAO_REG_4_, P1_DATAO_REG_5_,
    P1_DATAO_REG_6_, P1_DATAO_REG_7_, P1_DATAO_REG_8_, P1_DATAO_REG_9_,
    P1_DATAO_REG_10_, P1_DATAO_REG_11_, P1_DATAO_REG_12_, P1_DATAO_REG_13_,
    P1_DATAO_REG_14_, P1_DATAO_REG_15_, P1_DATAO_REG_16_, P1_DATAO_REG_17_,
    P1_DATAO_REG_18_, P1_DATAO_REG_19_, P1_DATAO_REG_20_, P1_DATAO_REG_21_,
    P1_DATAO_REG_22_, P1_DATAO_REG_23_, P1_DATAO_REG_24_, P1_DATAO_REG_25_,
    P1_DATAO_REG_26_, P1_DATAO_REG_27_, P1_DATAO_REG_28_, P1_DATAO_REG_29_,
    P1_DATAO_REG_30_, P1_DATAO_REG_31_, P1_EAX_REG_0_, P1_EAX_REG_1_,
    P1_EAX_REG_2_, P1_EAX_REG_3_, P1_EAX_REG_4_, P1_EAX_REG_5_,
    P1_EAX_REG_6_, P1_EAX_REG_7_, P1_EAX_REG_8_, P1_EAX_REG_9_,
    P1_EAX_REG_10_, P1_EAX_REG_11_, P1_EAX_REG_12_, P1_EAX_REG_13_,
    P1_EAX_REG_14_, P1_EAX_REG_15_, P1_EAX_REG_16_, P1_EAX_REG_17_,
    P1_EAX_REG_18_, P1_EAX_REG_19_, P1_EAX_REG_20_, P1_EAX_REG_21_,
    P1_EAX_REG_22_, P1_EAX_REG_23_, P1_EAX_REG_24_, P1_EAX_REG_25_,
    P1_EAX_REG_26_, P1_EAX_REG_27_, P1_EAX_REG_28_, P1_EAX_REG_29_,
    P1_EAX_REG_30_, P1_EAX_REG_31_, P1_EBX_REG_0_, P1_EBX_REG_1_,
    P1_EBX_REG_2_, P1_EBX_REG_3_, P1_EBX_REG_4_, P1_EBX_REG_5_,
    P1_EBX_REG_6_, P1_EBX_REG_7_, P1_EBX_REG_8_, P1_EBX_REG_9_,
    P1_EBX_REG_10_, P1_EBX_REG_11_, P1_EBX_REG_12_, P1_EBX_REG_13_,
    P1_EBX_REG_14_, P1_EBX_REG_15_, P1_EBX_REG_16_, P1_EBX_REG_17_,
    P1_EBX_REG_18_, P1_EBX_REG_19_, P1_EBX_REG_20_, P1_EBX_REG_21_,
    P1_EBX_REG_22_, P1_EBX_REG_23_, P1_EBX_REG_24_, P1_EBX_REG_25_,
    P1_EBX_REG_26_, P1_EBX_REG_27_, P1_EBX_REG_28_, P1_EBX_REG_29_,
    P1_EBX_REG_30_, P1_EBX_REG_31_, P1_REIP_REG_0_, P1_REIP_REG_1_,
    P1_REIP_REG_2_, P1_REIP_REG_3_, P1_REIP_REG_4_, P1_REIP_REG_5_,
    P1_REIP_REG_6_, P1_REIP_REG_7_, P1_REIP_REG_8_, P1_REIP_REG_9_,
    P1_REIP_REG_10_, P1_REIP_REG_11_, P1_REIP_REG_12_, P1_REIP_REG_13_,
    P1_REIP_REG_14_, P1_REIP_REG_15_, P1_REIP_REG_16_, P1_REIP_REG_17_,
    P1_REIP_REG_18_, P1_REIP_REG_19_, P1_REIP_REG_20_, P1_REIP_REG_21_,
    P1_REIP_REG_22_, P1_REIP_REG_23_, P1_REIP_REG_24_, P1_REIP_REG_25_,
    P1_REIP_REG_26_, P1_REIP_REG_27_, P1_REIP_REG_28_, P1_REIP_REG_29_,
    P1_REIP_REG_30_, P1_REIP_REG_31_, P1_BYTEENABLE_REG_3_,
    P1_BYTEENABLE_REG_2_, P1_BYTEENABLE_REG_1_, P1_BYTEENABLE_REG_0_,
    P1_W_R_N_REG, P1_FLUSH_REG, P1_MORE_REG, P1_STATEBS16_REG,
    P1_REQUESTPENDING_REG, P1_D_C_N_REG, P1_M_IO_N_REG, P1_CODEFETCH_REG,
    P1_ADS_N_REG, P1_READREQUEST_REG, P1_MEMORYFETCH_REG, Q_0, Q_1, Q_2,
    Q_3;
  wire new_P1_ADD_515_U182, new_P1_ADD_515_U181, new_P1_ADD_515_U180,
    new_U207, new_U208, new_U209, new_U210, new_U211, new_U247, new_U248,
    new_U249, new_U250, new_U283, new_U284, new_U285, new_U286, new_U287,
    new_U288, new_U289, new_U290, new_U291, new_U292, new_U293, new_U294,
    new_U295, new_U296, new_U297, new_U298, new_U299, new_U300, new_U301,
    new_U302, new_U303, new_U304, new_U305, new_U306, new_U307, new_U308,
    new_U309, new_U310, new_U311, new_U312, new_U313, new_U314, new_U315,
    new_U316, new_U317, new_U318, new_U319, new_U320, new_U321, new_U322,
    new_U323, new_U324, new_U325, new_U326, new_U327, new_U328, new_U329,
    new_U330, new_U331, new_U332, new_U333, new_U334, new_U335, new_U336,
    new_U337, new_U338, new_U339, new_U340, new_U341, new_U342, new_U343,
    new_U344, new_U345, new_U346, new_U377, new_U378, new_U379, new_U380,
    new_U381, new_U382, new_U383, new_U384, new_U385, new_U386, new_U387,
    new_U388, new_U389, new_U390, new_U391, new_U392, new_U393, new_U394,
    new_U395, new_U396, new_U397, new_U398, new_U399, new_U400, new_U401,
    new_U402, new_U403, new_U404, new_U405, new_U406, new_U407, new_U408,
    new_U409, new_U410, new_U411, new_U412, new_U413, new_U414, new_U415,
    new_U416, new_U417, new_U418, new_U419, new_U420, new_U421, new_U422,
    new_U423, new_U424, new_U425, new_U426, new_U427, new_U428, new_U429,
    new_U430, new_U431, new_U432, new_U433, new_U434, new_U435, new_U436,
    new_U437, new_U438, new_U439, new_U440, new_U441, new_U442, new_U443,
    new_U444, new_U445, new_U446, new_U447, new_U448, new_U449, new_U450,
    new_U451, new_U452, new_U453, new_U454, new_U455, new_U456, new_U457,
    new_U458, new_U459, new_U460, new_U461, new_U462, new_U463, new_U464,
    new_U465, new_U466, new_U467, new_U468, new_U469, new_U470, new_U471,
    new_U472, new_U473, new_U474, new_U475, new_U476, new_U477, new_U478,
    new_U479, new_U480, new_U481, new_U482, new_U483, new_U484, new_U485,
    new_U486, new_U487, new_U488, new_U489, new_U490, new_U491, new_U492,
    new_U493, new_U494, new_U495, new_U496, new_U497, new_U498, new_U499,
    new_U500, new_U501, new_U502, new_U503, new_U504, new_U505, new_U506,
    new_U507, new_U508, new_U509, new_U510, new_U511, new_U512, new_U513,
    new_U514, new_U515, new_U516, new_U517, new_U518, new_U519, new_U520,
    new_U521, new_U522, new_U523, new_U524, new_U525, new_U526, new_U527,
    new_U528, new_U529, new_U530, new_U531, new_U532, new_U533, new_U534,
    new_U535, new_U536, new_U537, new_U538, new_U539, new_U540, new_U541,
    new_U542, new_U543, new_U544, new_U545, new_U546, new_U547, new_U548,
    new_U549, new_U550, new_U551, new_U552, new_U553, new_U554, new_U555,
    new_U556, new_U557, new_U558, new_U559, new_U560, new_U561, new_U562,
    new_U563, new_U564, new_U565, new_U566, new_U567, new_U568, new_U569,
    new_U570, new_U571, new_U572, new_U573, new_U574, new_U575, new_U576,
    new_U577, new_U578, new_U579, new_U580, new_U581, new_U582, new_U583,
    new_U584, new_U585, new_U586, new_U587, new_U588, new_U589, new_U590,
    new_U591, new_U592, new_U593, new_U594, new_U595, new_U596, new_U597,
    new_U598, new_U599, new_U600, new_U601, new_U602, new_U603, new_U604,
    new_U605, new_U606, new_U607, new_U608, new_U609, new_U610, new_U611,
    new_U612, new_U613, new_U614, new_U615, new_U616, new_U617, new_U618,
    new_U619, new_U620, new_U621, new_U622, new_U623, new_U624, new_U625,
    new_U626, new_U627, new_U628, new_U629, new_U630, new_U631, new_U632,
    new_U633, new_U634, new_U635, new_U636, new_U637, new_U638, new_U639,
    new_U640, new_U641, new_U642, new_U643, new_U644, new_U645, new_U646,
    new_U647, new_U648, new_U649, new_U650, new_U651, new_U652, new_U653,
    new_U654, new_U655, new_U656, new_U657, new_U658, new_U659, new_U660,
    new_U661, new_U662, new_U663, new_U664, new_U665, new_U666, new_U667,
    new_U668, new_U669, new_U670, new_U671, new_U672, new_U673, new_U674,
    new_U675, new_U676, new_U677, new_U678, new_U679, new_U680, new_U681,
    new_U682, new_U683, new_U684, new_U685, new_U686, new_U687, new_U688,
    new_U689, new_U690, new_U691, new_U692, new_U693, new_U694, new_U695,
    new_U696, new_U697, new_U698, new_U699, new_U700, new_U701, new_U702,
    new_U703, new_U704, new_U705, new_U706, new_U707, new_U708, new_U709,
    new_U710, new_U711, new_U712, new_U713, new_U714, new_U715, new_U716,
    new_U717, new_U718, new_U719, new_U720, new_U721, new_U722, new_U723,
    new_U724, new_U725, new_U726, new_U727, new_U728, new_U729, new_U730,
    new_U731, new_U732, new_U733, new_U734, new_U735, new_U736,
    new_P1_ADD_515_U179, new_P1_ADD_515_U178, new_P1_ADD_515_U177,
    new_P1_ADD_515_U176, new_P1_ADD_515_U175, new_P1_ADD_515_U174,
    new_P1_ADD_515_U173, new_P1_ADD_515_U172, new_P1_ADD_515_U171,
    new_P3_U2352, new_P3_U2353, new_P3_U2354, new_P3_U2355, new_P3_U2356,
    new_P3_U2357, new_P3_U2358, new_P3_U2359, new_P3_U2360, new_P3_U2361,
    new_P3_U2362, new_P3_U2363, new_P3_U2364, new_P3_U2365, new_P3_U2366,
    new_P3_U2367, new_P3_U2368, new_P3_U2369, new_P3_U2370, new_P3_U2371,
    new_P3_U2372, new_P3_U2373, new_P3_U2374, new_P3_U2375, new_P3_U2376,
    new_P3_U2377, new_P3_U2378, new_P3_U2379, new_P3_U2380, new_P3_U2381,
    new_P3_U2382, new_P3_U2383, new_P3_U2384, new_P3_U2385, new_P3_U2386,
    new_P3_U2387, new_P3_U2388, new_P3_U2389, new_P3_U2390, new_P3_U2391,
    new_P3_U2392, new_P3_U2393, new_P3_U2394, new_P3_U2395, new_P3_U2396,
    new_P3_U2397, new_P3_U2398, new_P3_U2399, new_P3_U2400, new_P3_U2401,
    new_P3_U2402, new_P3_U2403, new_P3_U2404, new_P3_U2405, new_P3_U2406,
    new_P3_U2407, new_P3_U2408, new_P3_U2409, new_P3_U2410, new_P3_U2411,
    new_P3_U2412, new_P3_U2413, new_P3_U2414, new_P3_U2415, new_P3_U2416,
    new_P3_U2417, new_P3_U2418, new_P3_U2419, new_P3_U2420, new_P3_U2421,
    new_P3_U2422, new_P3_U2423, new_P3_U2424, new_P3_U2425, new_P3_U2426,
    new_P3_U2427, new_P3_U2428, new_P3_U2429, new_P3_U2430, new_P3_U2431,
    new_P3_U2432, new_P3_U2433, new_P3_U2434, new_P3_U2435, new_P3_U2436,
    new_P3_U2437, new_P3_U2438, new_P3_U2439, new_P3_U2440, new_P3_U2441,
    new_P3_U2442, new_P3_U2443, new_P3_U2444, new_P3_U2445, new_P3_U2446,
    new_P3_U2447, new_P3_U2448, new_P3_U2449, new_P3_U2450, new_P3_U2451,
    new_P3_U2452, new_P3_U2453, new_P3_U2454, new_P3_U2455, new_P3_U2456,
    new_P3_U2457, new_P3_U2458, new_P3_U2459, new_P3_U2460, new_P3_U2461,
    new_P3_U2462, new_P3_U2463, new_P3_U2464, new_P3_U2465, new_P3_U2466,
    new_P3_U2467, new_P3_U2468, new_P3_U2469, new_P3_U2470, new_P3_U2471,
    new_P3_U2472, new_P3_U2473, new_P3_U2474, new_P3_U2475, new_P3_U2476,
    new_P3_U2477, new_P3_U2478, new_P3_U2479, new_P3_U2480, new_P3_U2481,
    new_P3_U2482, new_P3_U2483, new_P3_U2484, new_P3_U2485, new_P3_U2486,
    new_P3_U2487, new_P3_U2488, new_P3_U2489, new_P3_U2490, new_P3_U2491,
    new_P3_U2492, new_P3_U2493, new_P3_U2494, new_P3_U2495, new_P3_U2496,
    new_P3_U2497, new_P3_U2498, new_P3_U2499, new_P3_U2500, new_P3_U2501,
    new_P3_U2502, new_P3_U2503, new_P3_U2504, new_P3_U2505, new_P3_U2506,
    new_P3_U2507, new_P3_U2508, new_P3_U2509, new_P3_U2510, new_P3_U2511,
    new_P3_U2512, new_P3_U2513, new_P3_U2514, new_P3_U2515, new_P3_U2516,
    new_P3_U2517, new_P3_U2518, new_P3_U2519, new_P3_U2520, new_P3_U2521,
    new_P3_U2522, new_P3_U2523, new_P3_U2524, new_P3_U2525, new_P3_U2526,
    new_P3_U2527, new_P3_U2528, new_P3_U2529, new_P3_U2530, new_P3_U2531,
    new_P3_U2532, new_P3_U2533, new_P3_U2534, new_P3_U2535, new_P3_U2536,
    new_P3_U2537, new_P3_U2538, new_P3_U2539, new_P3_U2540, new_P3_U2541,
    new_P3_U2542, new_P3_U2543, new_P3_U2544, new_P3_U2545, new_P3_U2546,
    new_P3_U2547, new_P3_U2548, new_P3_U2549, new_P3_U2550, new_P3_U2551,
    new_P3_U2552, new_P3_U2553, new_P3_U2554, new_P3_U2555, new_P3_U2556,
    new_P3_U2557, new_P3_U2558, new_P3_U2559, new_P3_U2560, new_P3_U2561,
    new_P3_U2562, new_P3_U2563, new_P3_U2564, new_P3_U2565, new_P3_U2566,
    new_P3_U2567, new_P3_U2568, new_P3_U2569, new_P3_U2570, new_P3_U2571,
    new_P3_U2572, new_P3_U2573, new_P3_U2574, new_P3_U2575, new_P3_U2576,
    new_P3_U2577, new_P3_U2578, new_P3_U2579, new_P3_U2580, new_P3_U2581,
    new_P3_U2582, new_P3_U2583, new_P3_U2584, new_P3_U2585, new_P3_U2586,
    new_P3_U2587, new_P3_U2588, new_P3_U2589, new_P3_U2590, new_P3_U2591,
    new_P3_U2592, new_P3_U2593, new_P3_U2594, new_P3_U2595, new_P3_U2596,
    new_P3_U2597, new_P3_U2598, new_P3_U2599, new_P3_U2600, new_P3_U2601,
    new_P3_U2602, new_P3_U2603, new_P3_U2604, new_P3_U2605, new_P3_U2606,
    new_P3_U2607, new_P3_U2608, new_P3_U2609, new_P3_U2610, new_P3_U2611,
    new_P3_U2612, new_P3_U2613, new_P3_U2614, new_P3_U2615, new_P3_U2616,
    new_P3_U2617, new_P3_U2618, new_P3_U2619, new_P3_U2620, new_P3_U2621,
    new_P3_U2622, new_P3_U2623, new_P3_U2624, new_P3_U2625, new_P3_U2626,
    new_P3_U2627, new_P3_U2628, new_P3_U2629, new_P3_U2630, new_P3_U2631,
    new_P3_U2632, new_P3_U3062, new_P3_U3063, new_P3_U3064, new_P3_U3065,
    new_P3_U3066, new_P3_U3067, new_P3_U3068, new_P3_U3069, new_P3_U3070,
    new_P3_U3071, new_P3_U3072, new_P3_U3073, new_P3_U3074, new_P3_U3075,
    new_P3_U3076, new_P3_U3077, new_P3_U3078, new_P3_U3079, new_P3_U3080,
    new_P3_U3081, new_P3_U3082, new_P3_U3083, new_P3_U3084, new_P3_U3085,
    new_P3_U3086, new_P3_U3087, new_P3_U3088, new_P3_U3089, new_P3_U3090,
    new_P3_U3091, new_P3_U3092, new_P3_U3093, new_P3_U3094, new_P3_U3095,
    new_P3_U3096, new_P3_U3097, new_P3_U3098, new_P3_U3099, new_P3_U3100,
    new_P3_U3101, new_P3_U3102, new_P3_U3103, new_P3_U3104, new_P3_U3105,
    new_P3_U3106, new_P3_U3107, new_P3_U3108, new_P3_U3109, new_P3_U3110,
    new_P3_U3111, new_P3_U3112, new_P3_U3113, new_P3_U3114, new_P3_U3115,
    new_P3_U3116, new_P3_U3117, new_P3_U3118, new_P3_U3119, new_P3_U3120,
    new_P3_U3121, new_P3_U3122, new_P3_U3123, new_P3_U3124, new_P3_U3125,
    new_P3_U3126, new_P3_U3127, new_P3_U3128, new_P3_U3129, new_P3_U3130,
    new_P3_U3131, new_P3_U3132, new_P3_U3133, new_P3_U3134, new_P3_U3135,
    new_P3_U3136, new_P3_U3137, new_P3_U3138, new_P3_U3139, new_P3_U3140,
    new_P3_U3141, new_P3_U3142, new_P3_U3143, new_P3_U3144, new_P3_U3145,
    new_P3_U3146, new_P3_U3147, new_P3_U3148, new_P3_U3149, new_P3_U3150,
    new_P3_U3151, new_P3_U3152, new_P3_U3153, new_P3_U3154, new_P3_U3155,
    new_P3_U3156, new_P3_U3157, new_P3_U3158, new_P3_U3159, new_P3_U3160,
    new_P3_U3161, new_P3_U3162, new_P3_U3163, new_P3_U3164, new_P3_U3165,
    new_P3_U3166, new_P3_U3167, new_P3_U3168, new_P3_U3169, new_P3_U3170,
    new_P3_U3171, new_P3_U3172, new_P3_U3173, new_P3_U3174, new_P3_U3175,
    new_P3_U3176, new_P3_U3177, new_P3_U3178, new_P3_U3179, new_P3_U3180,
    new_P3_U3181, new_P3_U3182, new_P3_U3183, new_P3_U3184, new_P3_U3185,
    new_P3_U3186, new_P3_U3187, new_P3_U3188, new_P3_U3189, new_P3_U3190,
    new_P3_U3191, new_P3_U3192, new_P3_U3193, new_P3_U3194, new_P3_U3195,
    new_P3_U3196, new_P3_U3197, new_P3_U3198, new_P3_U3199, new_P3_U3200,
    new_P3_U3201, new_P3_U3202, new_P3_U3203, new_P3_U3204, new_P3_U3205,
    new_P3_U3206, new_P3_U3207, new_P3_U3208, new_P3_U3209, new_P3_U3210,
    new_P3_U3211, new_P3_U3212, new_P3_U3213, new_P3_U3214, new_P3_U3215,
    new_P3_U3216, new_P3_U3217, new_P3_U3218, new_P3_U3219, new_P3_U3220,
    new_P3_U3221, new_P3_U3222, new_P3_U3223, new_P3_U3224, new_P3_U3225,
    new_P3_U3226, new_P3_U3227, new_P3_U3228, new_P3_U3229, new_P3_U3230,
    new_P3_U3231, new_P3_U3232, new_P3_U3233, new_P3_U3234, new_P3_U3235,
    new_P3_U3236, new_P3_U3237, new_P3_U3238, new_P3_U3239, new_P3_U3240,
    new_P3_U3241, new_P3_U3242, new_P3_U3243, new_P3_U3244, new_P3_U3245,
    new_P3_U3246, new_P3_U3247, new_P3_U3248, new_P3_U3249, new_P3_U3250,
    new_P3_U3251, new_P3_U3252, new_P3_U3253, new_P3_U3254, new_P3_U3255,
    new_P3_U3256, new_P3_U3257, new_P3_U3258, new_P3_U3259, new_P3_U3260,
    new_P3_U3261, new_P3_U3262, new_P3_U3263, new_P3_U3264, new_P3_U3265,
    new_P3_U3266, new_P3_U3267, new_P3_U3268, new_P3_U3269, new_P3_U3270,
    new_P3_U3271, new_P3_U3272, new_P3_U3273, new_P3_U3278, new_P3_U3279,
    new_P3_U3283, new_P3_U3286, new_P3_U3287, new_P3_U3291, new_P3_U3300,
    new_P3_U3301, new_P3_U3302, new_P3_U3303, new_P3_U3304, new_P3_U3305,
    new_P3_U3306, new_P3_U3307, new_P3_U3308, new_P3_U3309, new_P3_U3310,
    new_P3_U3311, new_P3_U3312, new_P3_U3313, new_P3_U3314, new_P3_U3315,
    new_P3_U3316, new_P3_U3317, new_P3_U3318, new_P3_U3319, new_P3_U3320,
    new_P3_U3321, new_P3_U3322, new_P3_U3323, new_P3_U3324, new_P3_U3325,
    new_P3_U3326, new_P3_U3327, new_P3_U3328, new_P3_U3329, new_P3_U3330,
    new_P3_U3331, new_P3_U3332, new_P3_U3333, new_P3_U3334, new_P3_U3335,
    new_P3_U3336, new_P3_U3337, new_P3_U3338, new_P3_U3339, new_P3_U3340,
    new_P3_U3341, new_P3_U3342, new_P3_U3343, new_P3_U3344, new_P3_U3345,
    new_P3_U3346, new_P3_U3347, new_P3_U3348, new_P3_U3349, new_P3_U3350,
    new_P3_U3351, new_P3_U3352, new_P3_U3353, new_P3_U3354, new_P3_U3355,
    new_P3_U3356, new_P3_U3357, new_P3_U3358, new_P3_U3359, new_P3_U3360,
    new_P3_U3361, new_P3_U3362, new_P3_U3363, new_P3_U3364, new_P3_U3365,
    new_P3_U3366, new_P3_U3367, new_P3_U3368, new_P3_U3369, new_P3_U3370,
    new_P3_U3371, new_P3_U3372, new_P3_U3373, new_P3_U3374, new_P3_U3375,
    new_P3_U3376, new_P3_U3377, new_P3_U3378, new_P3_U3379, new_P3_U3380,
    new_P3_U3381, new_P3_U3382, new_P3_U3383, new_P3_U3384, new_P3_U3385,
    new_P3_U3386, new_P3_U3387, new_P3_U3388, new_P3_U3389, new_P3_U3390,
    new_P3_U3391, new_P3_U3392, new_P3_U3393, new_P3_U3394, new_P3_U3395,
    new_P3_U3396, new_P3_U3397, new_P3_U3398, new_P3_U3399, new_P3_U3400,
    new_P3_U3401, new_P3_U3402, new_P3_U3403, new_P3_U3404, new_P3_U3405,
    new_P3_U3406, new_P3_U3407, new_P3_U3408, new_P3_U3409, new_P3_U3410,
    new_P3_U3411, new_P3_U3412, new_P3_U3413, new_P3_U3414, new_P3_U3415,
    new_P3_U3416, new_P3_U3417, new_P3_U3418, new_P3_U3419, new_P3_U3420,
    new_P3_U3421, new_P3_U3422, new_P3_U3423, new_P3_U3424, new_P3_U3425,
    new_P3_U3426, new_P3_U3427, new_P3_U3428, new_P3_U3429, new_P3_U3430,
    new_P3_U3431, new_P3_U3432, new_P3_U3433, new_P3_U3434, new_P3_U3435,
    new_P3_U3436, new_P3_U3437, new_P3_U3438, new_P3_U3439, new_P3_U3440,
    new_P3_U3441, new_P3_U3442, new_P3_U3443, new_P3_U3444, new_P3_U3445,
    new_P3_U3446, new_P3_U3447, new_P3_U3448, new_P3_U3449, new_P3_U3450,
    new_P3_U3451, new_P3_U3452, new_P3_U3453, new_P3_U3454, new_P3_U3455,
    new_P3_U3456, new_P3_U3457, new_P3_U3458, new_P3_U3459, new_P3_U3460,
    new_P3_U3461, new_P3_U3462, new_P3_U3463, new_P3_U3464, new_P3_U3465,
    new_P3_U3466, new_P3_U3467, new_P3_U3468, new_P3_U3469, new_P3_U3470,
    new_P3_U3471, new_P3_U3472, new_P3_U3473, new_P3_U3474, new_P3_U3475,
    new_P3_U3476, new_P3_U3477, new_P3_U3478, new_P3_U3479, new_P3_U3480,
    new_P3_U3481, new_P3_U3482, new_P3_U3483, new_P3_U3484, new_P3_U3485,
    new_P3_U3486, new_P3_U3487, new_P3_U3488, new_P3_U3489, new_P3_U3490,
    new_P3_U3491, new_P3_U3492, new_P3_U3493, new_P3_U3494, new_P3_U3495,
    new_P3_U3496, new_P3_U3497, new_P3_U3498, new_P3_U3499, new_P3_U3500,
    new_P3_U3501, new_P3_U3502, new_P3_U3503, new_P3_U3504, new_P3_U3505,
    new_P3_U3506, new_P3_U3507, new_P3_U3508, new_P3_U3509, new_P3_U3510,
    new_P3_U3511, new_P3_U3512, new_P3_U3513, new_P3_U3514, new_P3_U3515,
    new_P3_U3516, new_P3_U3517, new_P3_U3518, new_P3_U3519, new_P3_U3520,
    new_P3_U3521, new_P3_U3522, new_P3_U3523, new_P3_U3524, new_P3_U3525,
    new_P3_U3526, new_P3_U3527, new_P3_U3528, new_P3_U3529, new_P3_U3530,
    new_P3_U3531, new_P3_U3532, new_P3_U3533, new_P3_U3534, new_P3_U3535,
    new_P3_U3536, new_P3_U3537, new_P3_U3538, new_P3_U3539, new_P3_U3540,
    new_P3_U3541, new_P3_U3542, new_P3_U3543, new_P3_U3544, new_P3_U3545,
    new_P3_U3546, new_P3_U3547, new_P3_U3548, new_P3_U3549, new_P3_U3550,
    new_P3_U3551, new_P3_U3552, new_P3_U3553, new_P3_U3554, new_P3_U3555,
    new_P3_U3556, new_P3_U3557, new_P3_U3558, new_P3_U3559, new_P3_U3560,
    new_P3_U3561, new_P3_U3562, new_P3_U3563, new_P3_U3564, new_P3_U3565,
    new_P3_U3566, new_P3_U3567, new_P3_U3568, new_P3_U3569, new_P3_U3570,
    new_P3_U3571, new_P3_U3572, new_P3_U3573, new_P3_U3574, new_P3_U3575,
    new_P3_U3576, new_P3_U3577, new_P3_U3578, new_P3_U3579, new_P3_U3580,
    new_P3_U3581, new_P3_U3582, new_P3_U3583, new_P3_U3584, new_P3_U3585,
    new_P3_U3586, new_P3_U3587, new_P3_U3588, new_P3_U3589, new_P3_U3590,
    new_P3_U3591, new_P3_U3592, new_P3_U3593, new_P3_U3594, new_P3_U3595,
    new_P3_U3596, new_P3_U3597, new_P3_U3598, new_P3_U3599, new_P3_U3600,
    new_P3_U3601, new_P3_U3602, new_P3_U3603, new_P3_U3604, new_P3_U3605,
    new_P3_U3606, new_P3_U3607, new_P3_U3608, new_P3_U3609, new_P3_U3610,
    new_P3_U3611, new_P3_U3612, new_P3_U3613, new_P3_U3614, new_P3_U3615,
    new_P3_U3616, new_P3_U3617, new_P3_U3618, new_P3_U3619, new_P3_U3620,
    new_P3_U3621, new_P3_U3622, new_P3_U3623, new_P3_U3624, new_P3_U3625,
    new_P3_U3626, new_P3_U3627, new_P3_U3628, new_P3_U3629, new_P3_U3630,
    new_P3_U3631, new_P3_U3632, new_P3_U3633, new_P3_U3634, new_P3_U3635,
    new_P3_U3636, new_P3_U3637, new_P3_U3638, new_P3_U3639, new_P3_U3640,
    new_P3_U3641, new_P3_U3642, new_P3_U3643, new_P3_U3644, new_P3_U3645,
    new_P3_U3646, new_P3_U3647, new_P3_U3648, new_P3_U3649, new_P3_U3650,
    new_P3_U3651, new_P3_U3652, new_P3_U3653, new_P3_U3654, new_P3_U3655,
    new_P3_U3656, new_P3_U3657, new_P3_U3658, new_P3_U3659, new_P3_U3660,
    new_P3_U3661, new_P3_U3662, new_P3_U3663, new_P3_U3664, new_P3_U3665,
    new_P3_U3666, new_P3_U3667, new_P3_U3668, new_P3_U3669, new_P3_U3670,
    new_P3_U3671, new_P3_U3672, new_P3_U3673, new_P3_U3674, new_P3_U3675,
    new_P3_U3676, new_P3_U3677, new_P3_U3678, new_P3_U3679, new_P3_U3680,
    new_P3_U3681, new_P3_U3682, new_P3_U3683, new_P3_U3684, new_P3_U3685,
    new_P3_U3686, new_P3_U3687, new_P3_U3688, new_P3_U3689, new_P3_U3690,
    new_P3_U3691, new_P3_U3692, new_P3_U3693, new_P3_U3694, new_P3_U3695,
    new_P3_U3696, new_P3_U3697, new_P3_U3698, new_P3_U3699, new_P3_U3700,
    new_P3_U3701, new_P3_U3702, new_P3_U3703, new_P3_U3704, new_P3_U3705,
    new_P3_U3706, new_P3_U3707, new_P3_U3708, new_P3_U3709, new_P3_U3710,
    new_P3_U3711, new_P3_U3712, new_P3_U3713, new_P3_U3714, new_P3_U3715,
    new_P3_U3716, new_P3_U3717, new_P3_U3718, new_P3_U3719, new_P3_U3720,
    new_P3_U3721, new_P3_U3722, new_P3_U3723, new_P3_U3724, new_P3_U3725,
    new_P3_U3726, new_P3_U3727, new_P3_U3728, new_P3_U3729, new_P3_U3730,
    new_P3_U3731, new_P3_U3732, new_P3_U3733, new_P3_U3734, new_P3_U3735,
    new_P3_U3736, new_P3_U3737, new_P3_U3738, new_P3_U3739, new_P3_U3740,
    new_P3_U3741, new_P3_U3742, new_P3_U3743, new_P3_U3744, new_P3_U3745,
    new_P3_U3746, new_P3_U3747, new_P3_U3748, new_P3_U3749, new_P3_U3750,
    new_P3_U3751, new_P3_U3752, new_P3_U3753, new_P3_U3754, new_P3_U3755,
    new_P3_U3756, new_P3_U3757, new_P3_U3758, new_P3_U3759, new_P3_U3760,
    new_P3_U3761, new_P3_U3762, new_P3_U3763, new_P3_U3764, new_P3_U3765,
    new_P3_U3766, new_P3_U3767, new_P3_U3768, new_P3_U3769, new_P3_U3770,
    new_P3_U3771, new_P3_U3772, new_P3_U3773, new_P3_U3774, new_P3_U3775,
    new_P3_U3776, new_P3_U3777, new_P3_U3778, new_P3_U3779, new_P3_U3780,
    new_P3_U3781, new_P3_U3782, new_P3_U3783, new_P3_U3784, new_P3_U3785,
    new_P3_U3786, new_P3_U3787, new_P3_U3788, new_P3_U3789, new_P3_U3790,
    new_P3_U3791, new_P3_U3792, new_P3_U3793, new_P3_U3794, new_P3_U3795,
    new_P3_U3796, new_P3_U3797, new_P3_U3798, new_P3_U3799, new_P3_U3800,
    new_P3_U3801, new_P3_U3802, new_P3_U3803, new_P3_U3804, new_P3_U3805,
    new_P3_U3806, new_P3_U3807, new_P3_U3808, new_P3_U3809, new_P3_U3810,
    new_P3_U3811, new_P3_U3812, new_P3_U3813, new_P3_U3814, new_P3_U3815,
    new_P3_U3816, new_P3_U3817, new_P3_U3818, new_P3_U3819, new_P3_U3820,
    new_P3_U3821, new_P3_U3822, new_P3_U3823, new_P3_U3824, new_P3_U3825,
    new_P3_U3826, new_P3_U3827, new_P3_U3828, new_P3_U3829, new_P3_U3830,
    new_P3_U3831, new_P3_U3832, new_P3_U3833, new_P3_U3834, new_P3_U3835,
    new_P3_U3836, new_P3_U3837, new_P3_U3838, new_P3_U3839, new_P3_U3840,
    new_P3_U3841, new_P3_U3842, new_P3_U3843, new_P3_U3844, new_P3_U3845,
    new_P3_U3846, new_P3_U3847, new_P3_U3848, new_P3_U3849, new_P3_U3850,
    new_P3_U3851, new_P3_U3852, new_P3_U3853, new_P3_U3854, new_P3_U3855,
    new_P3_U3856, new_P3_U3857, new_P3_U3858, new_P3_U3859, new_P3_U3860,
    new_P3_U3861, new_P3_U3862, new_P3_U3863, new_P3_U3864, new_P3_U3865,
    new_P3_U3866, new_P3_U3867, new_P3_U3868, new_P3_U3869, new_P3_U3870,
    new_P3_U3871, new_P3_U3872, new_P3_U3873, new_P3_U3874, new_P3_U3875,
    new_P3_U3876, new_P3_U3877, new_P3_U3878, new_P3_U3879, new_P3_U3880,
    new_P3_U3881, new_P3_U3882, new_P3_U3883, new_P3_U3884, new_P3_U3885,
    new_P3_U3886, new_P3_U3887, new_P3_U3888, new_P3_U3889, new_P3_U3890,
    new_P3_U3891, new_P3_U3892, new_P3_U3893, new_P3_U3894, new_P3_U3895,
    new_P3_U3896, new_P3_U3897, new_P3_U3898, new_P3_U3899, new_P3_U3900,
    new_P3_U3901, new_P3_U3902, new_P3_U3903, new_P3_U3904, new_P3_U3905,
    new_P3_U3906, new_P3_U3907, new_P3_U3908, new_P3_U3909, new_P3_U3910,
    new_P3_U3911, new_P3_U3912, new_P3_U3913, new_P3_U3914, new_P3_U3915,
    new_P3_U3916, new_P3_U3917, new_P3_U3918, new_P3_U3919, new_P3_U3920,
    new_P3_U3921, new_P3_U3922, new_P3_U3923, new_P3_U3924, new_P3_U3925,
    new_P3_U3926, new_P3_U3927, new_P3_U3928, new_P3_U3929, new_P3_U3930,
    new_P3_U3931, new_P3_U3932, new_P3_U3933, new_P3_U3934, new_P3_U3935,
    new_P3_U3936, new_P3_U3937, new_P3_U3938, new_P3_U3939, new_P3_U3940,
    new_P3_U3941, new_P3_U3942, new_P3_U3943, new_P3_U3944, new_P3_U3945,
    new_P3_U3946, new_P3_U3947, new_P3_U3948, new_P3_U3949, new_P3_U3950,
    new_P3_U3951, new_P3_U3952, new_P3_U3953, new_P3_U3954, new_P3_U3955,
    new_P3_U3956, new_P3_U3957, new_P3_U3958, new_P3_U3959, new_P3_U3960,
    new_P3_U3961, new_P3_U3962, new_P3_U3963, new_P3_U3964, new_P3_U3965,
    new_P3_U3966, new_P3_U3967, new_P3_U3968, new_P3_U3969, new_P3_U3970,
    new_P3_U3971, new_P3_U3972, new_P3_U3973, new_P3_U3974, new_P3_U3975,
    new_P3_U3976, new_P3_U3977, new_P3_U3978, new_P3_U3979, new_P3_U3980,
    new_P3_U3981, new_P3_U3982, new_P3_U3983, new_P3_U3984, new_P3_U3985,
    new_P3_U3986, new_P3_U3987, new_P3_U3988, new_P3_U3989, new_P3_U3990,
    new_P3_U3991, new_P3_U3992, new_P3_U3993, new_P3_U3994, new_P3_U3995,
    new_P3_U3996, new_P3_U3997, new_P3_U3998, new_P3_U3999, new_P3_U4000,
    new_P3_U4001, new_P3_U4002, new_P3_U4003, new_P3_U4004, new_P3_U4005,
    new_P3_U4006, new_P3_U4007, new_P3_U4008, new_P3_U4009, new_P3_U4010,
    new_P3_U4011, new_P3_U4012, new_P3_U4013, new_P3_U4014, new_P3_U4015,
    new_P3_U4016, new_P3_U4017, new_P3_U4018, new_P3_U4019, new_P3_U4020,
    new_P3_U4021, new_P3_U4022, new_P3_U4023, new_P3_U4024, new_P3_U4025,
    new_P3_U4026, new_P3_U4027, new_P3_U4028, new_P3_U4029, new_P3_U4030,
    new_P3_U4031, new_P3_U4032, new_P3_U4033, new_P3_U4034, new_P3_U4035,
    new_P3_U4036, new_P3_U4037, new_P3_U4038, new_P3_U4039, new_P3_U4040,
    new_P3_U4041, new_P3_U4042, new_P3_U4043, new_P3_U4044, new_P3_U4045,
    new_P3_U4046, new_P3_U4047, new_P3_U4048, new_P3_U4049, new_P3_U4050,
    new_P3_U4051, new_P3_U4052, new_P3_U4053, new_P3_U4054, new_P3_U4055,
    new_P3_U4056, new_P3_U4057, new_P3_U4058, new_P3_U4059, new_P3_U4060,
    new_P3_U4061, new_P3_U4062, new_P3_U4063, new_P3_U4064, new_P3_U4065,
    new_P3_U4066, new_P3_U4067, new_P3_U4068, new_P3_U4069, new_P3_U4070,
    new_P3_U4071, new_P3_U4072, new_P3_U4073, new_P3_U4074, new_P3_U4075,
    new_P3_U4076, new_P3_U4077, new_P3_U4078, new_P3_U4079, new_P3_U4080,
    new_P3_U4081, new_P3_U4082, new_P3_U4083, new_P3_U4084, new_P3_U4085,
    new_P3_U4086, new_P3_U4087, new_P3_U4088, new_P3_U4089, new_P3_U4090,
    new_P3_U4091, new_P3_U4092, new_P3_U4093, new_P3_U4094, new_P3_U4095,
    new_P3_U4096, new_P3_U4097, new_P3_U4098, new_P3_U4099, new_P3_U4100,
    new_P3_U4101, new_P3_U4102, new_P3_U4103, new_P3_U4104, new_P3_U4105,
    new_P3_U4106, new_P3_U4107, new_P3_U4108, new_P3_U4109, new_P3_U4110,
    new_P3_U4111, new_P3_U4112, new_P3_U4113, new_P3_U4114, new_P3_U4115,
    new_P3_U4116, new_P3_U4117, new_P3_U4118, new_P3_U4119, new_P3_U4120,
    new_P3_U4121, new_P3_U4122, new_P3_U4123, new_P3_U4124, new_P3_U4125,
    new_P3_U4126, new_P3_U4127, new_P3_U4128, new_P3_U4129, new_P3_U4130,
    new_P3_U4131, new_P3_U4132, new_P3_U4133, new_P3_U4134, new_P3_U4135,
    new_P3_U4136, new_P3_U4137, new_P3_U4138, new_P3_U4139, new_P3_U4140,
    new_P3_U4141, new_P3_U4142, new_P3_U4143, new_P3_U4144, new_P3_U4145,
    new_P3_U4146, new_P3_U4147, new_P3_U4148, new_P3_U4149, new_P3_U4150,
    new_P3_U4151, new_P3_U4152, new_P3_U4153, new_P3_U4154, new_P3_U4155,
    new_P3_U4156, new_P3_U4157, new_P3_U4158, new_P3_U4159, new_P3_U4160,
    new_P3_U4161, new_P3_U4162, new_P3_U4163, new_P3_U4164, new_P3_U4165,
    new_P3_U4166, new_P3_U4167, new_P3_U4168, new_P3_U4169, new_P3_U4170,
    new_P3_U4171, new_P3_U4172, new_P3_U4173, new_P3_U4174, new_P3_U4175,
    new_P3_U4176, new_P3_U4177, new_P3_U4178, new_P3_U4179, new_P3_U4180,
    new_P3_U4181, new_P3_U4182, new_P3_U4183, new_P3_U4184, new_P3_U4185,
    new_P3_U4186, new_P3_U4187, new_P3_U4188, new_P3_U4189, new_P3_U4190,
    new_P3_U4191, new_P3_U4192, new_P3_U4193, new_P3_U4194, new_P3_U4195,
    new_P3_U4196, new_P3_U4197, new_P3_U4198, new_P3_U4199, new_P3_U4200,
    new_P3_U4201, new_P3_U4202, new_P3_U4203, new_P3_U4204, new_P3_U4205,
    new_P3_U4206, new_P3_U4207, new_P3_U4208, new_P3_U4209, new_P3_U4210,
    new_P3_U4211, new_P3_U4212, new_P3_U4213, new_P3_U4214, new_P3_U4215,
    new_P3_U4216, new_P3_U4217, new_P3_U4218, new_P3_U4219, new_P3_U4220,
    new_P3_U4221, new_P3_U4222, new_P3_U4223, new_P3_U4224, new_P3_U4225,
    new_P3_U4226, new_P3_U4227, new_P3_U4228, new_P3_U4229, new_P3_U4230,
    new_P3_U4231, new_P3_U4232, new_P3_U4233, new_P3_U4234, new_P3_U4235,
    new_P3_U4236, new_P3_U4237, new_P3_U4238, new_P3_U4239, new_P3_U4240,
    new_P3_U4241, new_P3_U4242, new_P3_U4243, new_P3_U4244, new_P3_U4245,
    new_P3_U4246, new_P3_U4247, new_P3_U4248, new_P3_U4249, new_P3_U4250,
    new_P3_U4251, new_P3_U4252, new_P3_U4253, new_P3_U4254, new_P3_U4255,
    new_P3_U4256, new_P3_U4257, new_P3_U4258, new_P3_U4259, new_P3_U4260,
    new_P3_U4261, new_P3_U4262, new_P3_U4263, new_P3_U4264, new_P3_U4265,
    new_P3_U4266, new_P3_U4267, new_P3_U4268, new_P3_U4269, new_P3_U4270,
    new_P3_U4271, new_P3_U4272, new_P3_U4273, new_P3_U4274, new_P3_U4275,
    new_P3_U4276, new_P3_U4277, new_P3_U4278, new_P3_U4279, new_P3_U4280,
    new_P3_U4281, new_P3_U4282, new_P3_U4283, new_P3_U4284, new_P3_U4285,
    new_P3_U4286, new_P3_U4287, new_P3_U4288, new_P3_U4289, new_P3_U4290,
    new_P3_U4291, new_P3_U4292, new_P3_U4293, new_P3_U4294, new_P3_U4295,
    new_P3_U4296, new_P3_U4297, new_P3_U4298, new_P3_U4299, new_P3_U4300,
    new_P3_U4301, new_P3_U4302, new_P3_U4303, new_P3_U4304, new_P3_U4305,
    new_P3_U4306, new_P3_U4307, new_P3_U4308, new_P3_U4309, new_P3_U4310,
    new_P3_U4311, new_P3_U4312, new_P3_U4313, new_P3_U4314, new_P3_U4315,
    new_P3_U4316, new_P3_U4317, new_P3_U4318, new_P3_U4319, new_P3_U4320,
    new_P3_U4321, new_P3_U4322, new_P3_U4323, new_P3_U4324, new_P3_U4325,
    new_P3_U4326, new_P3_U4327, new_P3_U4328, new_P3_U4329, new_P3_U4330,
    new_P3_U4331, new_P3_U4332, new_P3_U4333, new_P3_U4334, new_P3_U4335,
    new_P3_U4336, new_P3_U4337, new_P3_U4338, new_P3_U4339, new_P3_U4340,
    new_P3_U4341, new_P3_U4342, new_P3_U4343, new_P3_U4344, new_P3_U4345,
    new_P3_U4346, new_P3_U4347, new_P3_U4348, new_P3_U4349, new_P3_U4350,
    new_P3_U4351, new_P3_U4352, new_P3_U4353, new_P3_U4354, new_P3_U4355,
    new_P3_U4356, new_P3_U4357, new_P3_U4358, new_P3_U4359, new_P3_U4360,
    new_P3_U4361, new_P3_U4362, new_P3_U4363, new_P3_U4364, new_P3_U4365,
    new_P3_U4366, new_P3_U4367, new_P3_U4368, new_P3_U4369, new_P3_U4370,
    new_P3_U4371, new_P3_U4372, new_P3_U4373, new_P3_U4374, new_P3_U4375,
    new_P3_U4376, new_P3_U4377, new_P3_U4378, new_P3_U4379, new_P3_U4380,
    new_P3_U4381, new_P3_U4382, new_P3_U4383, new_P3_U4384, new_P3_U4385,
    new_P3_U4386, new_P3_U4387, new_P3_U4388, new_P3_U4389, new_P3_U4390,
    new_P3_U4391, new_P3_U4392, new_P3_U4393, new_P3_U4394, new_P3_U4395,
    new_P3_U4396, new_P3_U4397, new_P3_U4398, new_P3_U4399, new_P3_U4400,
    new_P3_U4401, new_P3_U4402, new_P3_U4403, new_P3_U4404, new_P3_U4405,
    new_P3_U4406, new_P3_U4407, new_P3_U4408, new_P3_U4409, new_P3_U4410,
    new_P3_U4411, new_P3_U4412, new_P3_U4413, new_P3_U4414, new_P3_U4415,
    new_P3_U4416, new_P3_U4417, new_P3_U4418, new_P3_U4419, new_P3_U4420,
    new_P3_U4421, new_P3_U4422, new_P3_U4423, new_P3_U4424, new_P3_U4425,
    new_P3_U4426, new_P3_U4427, new_P3_U4428, new_P3_U4429, new_P3_U4430,
    new_P3_U4431, new_P3_U4432, new_P3_U4433, new_P3_U4434, new_P3_U4435,
    new_P3_U4436, new_P3_U4437, new_P3_U4438, new_P3_U4439, new_P3_U4440,
    new_P3_U4441, new_P3_U4442, new_P3_U4443, new_P3_U4444, new_P3_U4445,
    new_P3_U4446, new_P3_U4447, new_P3_U4448, new_P3_U4449, new_P3_U4450,
    new_P3_U4451, new_P3_U4452, new_P3_U4453, new_P3_U4454, new_P3_U4455,
    new_P3_U4456, new_P3_U4457, new_P3_U4458, new_P3_U4459, new_P3_U4460,
    new_P3_U4461, new_P3_U4462, new_P3_U4463, new_P3_U4464, new_P3_U4465,
    new_P3_U4466, new_P3_U4467, new_P3_U4468, new_P3_U4469, new_P3_U4470,
    new_P3_U4471, new_P3_U4472, new_P3_U4473, new_P3_U4474, new_P3_U4475,
    new_P3_U4476, new_P3_U4477, new_P3_U4478, new_P3_U4479, new_P3_U4480,
    new_P3_U4481, new_P3_U4482, new_P3_U4483, new_P3_U4484, new_P3_U4485,
    new_P3_U4486, new_P3_U4487, new_P3_U4488, new_P3_U4489, new_P3_U4490,
    new_P3_U4491, new_P3_U4492, new_P3_U4493, new_P3_U4494, new_P3_U4495,
    new_P3_U4496, new_P3_U4497, new_P3_U4498, new_P3_U4499, new_P3_U4500,
    new_P3_U4501, new_P3_U4502, new_P3_U4503, new_P3_U4504, new_P3_U4505,
    new_P3_U4506, new_P3_U4507, new_P3_U4508, new_P3_U4509, new_P3_U4510,
    new_P3_U4511, new_P3_U4512, new_P3_U4513, new_P3_U4514, new_P3_U4515,
    new_P3_U4516, new_P3_U4517, new_P3_U4518, new_P3_U4519, new_P3_U4520,
    new_P3_U4521, new_P3_U4522, new_P3_U4523, new_P3_U4524, new_P3_U4525,
    new_P3_U4526, new_P3_U4527, new_P3_U4528, new_P3_U4529, new_P3_U4530,
    new_P3_U4531, new_P3_U4532, new_P3_U4533, new_P3_U4534, new_P3_U4535,
    new_P3_U4536, new_P3_U4537, new_P3_U4538, new_P3_U4539, new_P3_U4540,
    new_P3_U4541, new_P3_U4542, new_P3_U4543, new_P3_U4544, new_P3_U4545,
    new_P3_U4546, new_P3_U4547, new_P3_U4548, new_P3_U4549, new_P3_U4550,
    new_P3_U4551, new_P3_U4552, new_P3_U4553, new_P3_U4554, new_P3_U4555,
    new_P3_U4556, new_P3_U4557, new_P3_U4558, new_P3_U4559, new_P3_U4560,
    new_P3_U4561, new_P3_U4562, new_P3_U4563, new_P3_U4564, new_P3_U4565,
    new_P3_U4566, new_P3_U4567, new_P3_U4568, new_P3_U4569, new_P3_U4570,
    new_P3_U4571, new_P3_U4572, new_P3_U4573, new_P3_U4574, new_P3_U4575,
    new_P3_U4576, new_P3_U4577, new_P3_U4578, new_P3_U4579, new_P3_U4580,
    new_P3_U4581, new_P3_U4582, new_P3_U4583, new_P3_U4584, new_P3_U4585,
    new_P3_U4586, new_P3_U4587, new_P3_U4588, new_P3_U4589, new_P3_U4590,
    new_P3_U4591, new_P3_U4592, new_P3_U4593, new_P3_U4594, new_P3_U4595,
    new_P3_U4596, new_P3_U4597, new_P3_U4598, new_P3_U4599, new_P3_U4600,
    new_P3_U4601, new_P3_U4602, new_P3_U4603, new_P3_U4604, new_P3_U4605,
    new_P3_U4606, new_P3_U4607, new_P3_U4608, new_P3_U4609, new_P3_U4610,
    new_P3_U4611, new_P3_U4612, new_P3_U4613, new_P3_U4614, new_P3_U4615,
    new_P3_U4616, new_P3_U4617, new_P3_U4618, new_P3_U4619, new_P3_U4620,
    new_P3_U4621, new_P3_U4622, new_P3_U4623, new_P3_U4624, new_P3_U4625,
    new_P3_U4626, new_P3_U4627, new_P3_U4628, new_P3_U4629, new_P3_U4630,
    new_P3_U4631, new_P3_U4632, new_P3_U4633, new_P3_U4634, new_P3_U4635,
    new_P3_U4636, new_P3_U4637, new_P3_U4638, new_P3_U4639, new_P3_U4640,
    new_P3_U4641, new_P3_U4642, new_P3_U4643, new_P3_U4644, new_P3_U4645,
    new_P3_U4646, new_P3_U4647, new_P3_U4648, new_P3_U4649, new_P3_U4650,
    new_P3_U4651, new_P3_U4652, new_P3_U4653, new_P3_U4654, new_P3_U4655,
    new_P3_U4656, new_P3_U4657, new_P3_U4658, new_P3_U4659, new_P3_U4660,
    new_P3_U4661, new_P3_U4662, new_P3_U4663, new_P3_U4664, new_P3_U4665,
    new_P3_U4666, new_P3_U4667, new_P3_U4668, new_P3_U4669, new_P3_U4670,
    new_P3_U4671, new_P3_U4672, new_P3_U4673, new_P3_U4674, new_P3_U4675,
    new_P3_U4676, new_P3_U4677, new_P3_U4678, new_P3_U4679, new_P3_U4680,
    new_P3_U4681, new_P3_U4682, new_P3_U4683, new_P3_U4684, new_P3_U4685,
    new_P3_U4686, new_P3_U4687, new_P3_U4688, new_P3_U4689, new_P3_U4690,
    new_P3_U4691, new_P3_U4692, new_P3_U4693, new_P3_U4694, new_P3_U4695,
    new_P3_U4696, new_P3_U4697, new_P3_U4698, new_P3_U4699, new_P3_U4700,
    new_P3_U4701, new_P3_U4702, new_P3_U4703, new_P3_U4704, new_P3_U4705,
    new_P3_U4706, new_P3_U4707, new_P3_U4708, new_P3_U4709, new_P3_U4710,
    new_P3_U4711, new_P3_U4712, new_P3_U4713, new_P3_U4714, new_P3_U4715,
    new_P3_U4716, new_P3_U4717, new_P3_U4718, new_P3_U4719, new_P3_U4720,
    new_P3_U4721, new_P3_U4722, new_P3_U4723, new_P3_U4724, new_P3_U4725,
    new_P3_U4726, new_P3_U4727, new_P3_U4728, new_P3_U4729, new_P3_U4730,
    new_P3_U4731, new_P3_U4732, new_P3_U4733, new_P3_U4734, new_P3_U4735,
    new_P3_U4736, new_P3_U4737, new_P3_U4738, new_P3_U4739, new_P3_U4740,
    new_P3_U4741, new_P3_U4742, new_P3_U4743, new_P3_U4744, new_P3_U4745,
    new_P3_U4746, new_P3_U4747, new_P3_U4748, new_P3_U4749, new_P3_U4750,
    new_P3_U4751, new_P3_U4752, new_P3_U4753, new_P3_U4754, new_P3_U4755,
    new_P3_U4756, new_P3_U4757, new_P3_U4758, new_P3_U4759, new_P3_U4760,
    new_P3_U4761, new_P3_U4762, new_P3_U4763, new_P3_U4764, new_P3_U4765,
    new_P3_U4766, new_P3_U4767, new_P3_U4768, new_P3_U4769, new_P3_U4770,
    new_P3_U4771, new_P3_U4772, new_P3_U4773, new_P3_U4774, new_P3_U4775,
    new_P3_U4776, new_P3_U4777, new_P3_U4778, new_P3_U4779, new_P3_U4780,
    new_P3_U4781, new_P3_U4782, new_P3_U4783, new_P3_U4784, new_P3_U4785,
    new_P3_U4786, new_P3_U4787, new_P3_U4788, new_P3_U4789, new_P3_U4790,
    new_P3_U4791, new_P3_U4792, new_P3_U4793, new_P3_U4794, new_P3_U4795,
    new_P3_U4796, new_P3_U4797, new_P3_U4798, new_P3_U4799, new_P3_U4800,
    new_P3_U4801, new_P3_U4802, new_P3_U4803, new_P3_U4804, new_P3_U4805,
    new_P3_U4806, new_P3_U4807, new_P3_U4808, new_P3_U4809, new_P3_U4810,
    new_P3_U4811, new_P3_U4812, new_P3_U4813, new_P3_U4814, new_P3_U4815,
    new_P3_U4816, new_P3_U4817, new_P3_U4818, new_P3_U4819, new_P3_U4820,
    new_P3_U4821, new_P3_U4822, new_P3_U4823, new_P3_U4824, new_P3_U4825,
    new_P3_U4826, new_P3_U4827, new_P3_U4828, new_P3_U4829, new_P3_U4830,
    new_P3_U4831, new_P3_U4832, new_P3_U4833, new_P3_U4834, new_P3_U4835,
    new_P3_U4836, new_P3_U4837, new_P3_U4838, new_P3_U4839, new_P3_U4840,
    new_P3_U4841, new_P3_U4842, new_P3_U4843, new_P3_U4844, new_P3_U4845,
    new_P3_U4846, new_P3_U4847, new_P3_U4848, new_P3_U4849, new_P3_U4850,
    new_P3_U4851, new_P3_U4852, new_P3_U4853, new_P3_U4854, new_P3_U4855,
    new_P3_U4856, new_P3_U4857, new_P3_U4858, new_P3_U4859, new_P3_U4860,
    new_P3_U4861, new_P3_U4862, new_P3_U4863, new_P3_U4864, new_P3_U4865,
    new_P3_U4866, new_P3_U4867, new_P3_U4868, new_P3_U4869, new_P3_U4870,
    new_P3_U4871, new_P3_U4872, new_P3_U4873, new_P3_U4874, new_P3_U4875,
    new_P3_U4876, new_P3_U4877, new_P3_U4878, new_P3_U4879, new_P3_U4880,
    new_P3_U4881, new_P3_U4882, new_P3_U4883, new_P3_U4884, new_P3_U4885,
    new_P3_U4886, new_P3_U4887, new_P3_U4888, new_P3_U4889, new_P3_U4890,
    new_P3_U4891, new_P3_U4892, new_P3_U4893, new_P3_U4894, new_P3_U4895,
    new_P3_U4896, new_P3_U4897, new_P3_U4898, new_P3_U4899, new_P3_U4900,
    new_P3_U4901, new_P3_U4902, new_P3_U4903, new_P3_U4904, new_P3_U4905,
    new_P3_U4906, new_P3_U4907, new_P3_U4908, new_P3_U4909, new_P3_U4910,
    new_P3_U4911, new_P3_U4912, new_P3_U4913, new_P3_U4914, new_P3_U4915,
    new_P3_U4916, new_P3_U4917, new_P3_U4918, new_P3_U4919, new_P3_U4920,
    new_P3_U4921, new_P3_U4922, new_P3_U4923, new_P3_U4924, new_P3_U4925,
    new_P3_U4926, new_P3_U4927, new_P3_U4928, new_P3_U4929, new_P3_U4930,
    new_P3_U4931, new_P3_U4932, new_P3_U4933, new_P3_U4934, new_P3_U4935,
    new_P3_U4936, new_P3_U4937, new_P3_U4938, new_P3_U4939, new_P3_U4940,
    new_P3_U4941, new_P3_U4942, new_P3_U4943, new_P3_U4944, new_P3_U4945,
    new_P3_U4946, new_P3_U4947, new_P3_U4948, new_P3_U4949, new_P3_U4950,
    new_P3_U4951, new_P3_U4952, new_P3_U4953, new_P3_U4954, new_P3_U4955,
    new_P3_U4956, new_P3_U4957, new_P3_U4958, new_P3_U4959, new_P3_U4960,
    new_P3_U4961, new_P3_U4962, new_P3_U4963, new_P3_U4964, new_P3_U4965,
    new_P3_U4966, new_P3_U4967, new_P3_U4968, new_P3_U4969, new_P3_U4970,
    new_P3_U4971, new_P3_U4972, new_P3_U4973, new_P3_U4974, new_P3_U4975,
    new_P3_U4976, new_P3_U4977, new_P3_U4978, new_P3_U4979, new_P3_U4980,
    new_P3_U4981, new_P3_U4982, new_P3_U4983, new_P3_U4984, new_P3_U4985,
    new_P3_U4986, new_P3_U4987, new_P3_U4988, new_P3_U4989, new_P3_U4990,
    new_P3_U4991, new_P3_U4992, new_P3_U4993, new_P3_U4994, new_P3_U4995,
    new_P3_U4996, new_P3_U4997, new_P3_U4998, new_P3_U4999, new_P3_U5000,
    new_P3_U5001, new_P3_U5002, new_P3_U5003, new_P3_U5004, new_P3_U5005,
    new_P3_U5006, new_P3_U5007, new_P3_U5008, new_P3_U5009, new_P3_U5010,
    new_P3_U5011, new_P3_U5012, new_P3_U5013, new_P3_U5014, new_P3_U5015,
    new_P3_U5016, new_P3_U5017, new_P3_U5018, new_P3_U5019, new_P3_U5020,
    new_P3_U5021, new_P3_U5022, new_P3_U5023, new_P3_U5024, new_P3_U5025,
    new_P3_U5026, new_P3_U5027, new_P3_U5028, new_P3_U5029, new_P3_U5030,
    new_P3_U5031, new_P3_U5032, new_P3_U5033, new_P3_U5034, new_P3_U5035,
    new_P3_U5036, new_P3_U5037, new_P3_U5038, new_P3_U5039, new_P3_U5040,
    new_P3_U5041, new_P3_U5042, new_P3_U5043, new_P3_U5044, new_P3_U5045,
    new_P3_U5046, new_P3_U5047, new_P3_U5048, new_P3_U5049, new_P3_U5050,
    new_P3_U5051, new_P3_U5052, new_P3_U5053, new_P3_U5054, new_P3_U5055,
    new_P3_U5056, new_P3_U5057, new_P3_U5058, new_P3_U5059, new_P3_U5060,
    new_P3_U5061, new_P3_U5062, new_P3_U5063, new_P3_U5064, new_P3_U5065,
    new_P3_U5066, new_P3_U5067, new_P3_U5068, new_P3_U5069, new_P3_U5070,
    new_P3_U5071, new_P3_U5072, new_P3_U5073, new_P3_U5074, new_P3_U5075,
    new_P3_U5076, new_P3_U5077, new_P3_U5078, new_P3_U5079, new_P3_U5080,
    new_P3_U5081, new_P3_U5082, new_P3_U5083, new_P3_U5084, new_P3_U5085,
    new_P3_U5086, new_P3_U5087, new_P3_U5088, new_P3_U5089, new_P3_U5090,
    new_P3_U5091, new_P3_U5092, new_P3_U5093, new_P3_U5094, new_P3_U5095,
    new_P3_U5096, new_P3_U5097, new_P3_U5098, new_P3_U5099, new_P3_U5100,
    new_P3_U5101, new_P3_U5102, new_P3_U5103, new_P3_U5104, new_P3_U5105,
    new_P3_U5106, new_P3_U5107, new_P3_U5108, new_P3_U5109, new_P3_U5110,
    new_P3_U5111, new_P3_U5112, new_P3_U5113, new_P3_U5114, new_P3_U5115,
    new_P3_U5116, new_P3_U5117, new_P3_U5118, new_P3_U5119, new_P3_U5120,
    new_P3_U5121, new_P3_U5122, new_P3_U5123, new_P3_U5124, new_P3_U5125,
    new_P3_U5126, new_P3_U5127, new_P3_U5128, new_P3_U5129, new_P3_U5130,
    new_P3_U5131, new_P3_U5132, new_P3_U5133, new_P3_U5134, new_P3_U5135,
    new_P3_U5136, new_P3_U5137, new_P3_U5138, new_P3_U5139, new_P3_U5140,
    new_P3_U5141, new_P3_U5142, new_P3_U5143, new_P3_U5144, new_P3_U5145,
    new_P3_U5146, new_P3_U5147, new_P3_U5148, new_P3_U5149, new_P3_U5150,
    new_P3_U5151, new_P3_U5152, new_P3_U5153, new_P3_U5154, new_P3_U5155,
    new_P3_U5156, new_P3_U5157, new_P3_U5158, new_P3_U5159, new_P3_U5160,
    new_P3_U5161, new_P3_U5162, new_P3_U5163, new_P3_U5164, new_P3_U5165,
    new_P3_U5166, new_P3_U5167, new_P3_U5168, new_P3_U5169, new_P3_U5170,
    new_P3_U5171, new_P3_U5172, new_P3_U5173, new_P3_U5174, new_P3_U5175,
    new_P3_U5176, new_P3_U5177, new_P3_U5178, new_P3_U5179, new_P3_U5180,
    new_P3_U5181, new_P3_U5182, new_P3_U5183, new_P3_U5184, new_P3_U5185,
    new_P3_U5186, new_P3_U5187, new_P3_U5188, new_P3_U5189, new_P3_U5190,
    new_P3_U5191, new_P3_U5192, new_P3_U5193, new_P3_U5194, new_P3_U5195,
    new_P3_U5196, new_P3_U5197, new_P3_U5198, new_P3_U5199, new_P3_U5200,
    new_P3_U5201, new_P3_U5202, new_P3_U5203, new_P3_U5204, new_P3_U5205,
    new_P3_U5206, new_P3_U5207, new_P3_U5208, new_P3_U5209, new_P3_U5210,
    new_P3_U5211, new_P3_U5212, new_P3_U5213, new_P3_U5214, new_P3_U5215,
    new_P3_U5216, new_P3_U5217, new_P3_U5218, new_P3_U5219, new_P3_U5220,
    new_P3_U5221, new_P3_U5222, new_P3_U5223, new_P3_U5224, new_P3_U5225,
    new_P3_U5226, new_P3_U5227, new_P3_U5228, new_P3_U5229, new_P3_U5230,
    new_P3_U5231, new_P3_U5232, new_P3_U5233, new_P3_U5234, new_P3_U5235,
    new_P3_U5236, new_P3_U5237, new_P3_U5238, new_P3_U5239, new_P3_U5240,
    new_P3_U5241, new_P3_U5242, new_P3_U5243, new_P3_U5244, new_P3_U5245,
    new_P3_U5246, new_P3_U5247, new_P3_U5248, new_P3_U5249, new_P3_U5250,
    new_P3_U5251, new_P3_U5252, new_P3_U5253, new_P3_U5254, new_P3_U5255,
    new_P3_U5256, new_P3_U5257, new_P3_U5258, new_P3_U5259, new_P3_U5260,
    new_P3_U5261, new_P3_U5262, new_P3_U5263, new_P3_U5264, new_P3_U5265,
    new_P3_U5266, new_P3_U5267, new_P3_U5268, new_P3_U5269, new_P3_U5270,
    new_P3_U5271, new_P3_U5272, new_P3_U5273, new_P3_U5274, new_P3_U5275,
    new_P3_U5276, new_P3_U5277, new_P3_U5278, new_P3_U5279, new_P3_U5280,
    new_P3_U5281, new_P3_U5282, new_P3_U5283, new_P3_U5284, new_P3_U5285,
    new_P3_U5286, new_P3_U5287, new_P3_U5288, new_P3_U5289, new_P3_U5290,
    new_P3_U5291, new_P3_U5292, new_P3_U5293, new_P3_U5294, new_P3_U5295,
    new_P3_U5296, new_P3_U5297, new_P3_U5298, new_P3_U5299, new_P3_U5300,
    new_P3_U5301, new_P3_U5302, new_P3_U5303, new_P3_U5304, new_P3_U5305,
    new_P3_U5306, new_P3_U5307, new_P3_U5308, new_P3_U5309, new_P3_U5310,
    new_P3_U5311, new_P3_U5312, new_P3_U5313, new_P3_U5314, new_P3_U5315,
    new_P3_U5316, new_P3_U5317, new_P3_U5318, new_P3_U5319, new_P3_U5320,
    new_P3_U5321, new_P3_U5322, new_P3_U5323, new_P3_U5324, new_P3_U5325,
    new_P3_U5326, new_P3_U5327, new_P3_U5328, new_P3_U5329, new_P3_U5330,
    new_P3_U5331, new_P3_U5332, new_P3_U5333, new_P3_U5334, new_P3_U5335,
    new_P3_U5336, new_P3_U5337, new_P3_U5338, new_P3_U5339, new_P3_U5340,
    new_P3_U5341, new_P3_U5342, new_P3_U5343, new_P3_U5344, new_P3_U5345,
    new_P3_U5346, new_P3_U5347, new_P3_U5348, new_P3_U5349, new_P3_U5350,
    new_P3_U5351, new_P3_U5352, new_P3_U5353, new_P3_U5354, new_P3_U5355,
    new_P3_U5356, new_P3_U5357, new_P3_U5358, new_P3_U5359, new_P3_U5360,
    new_P3_U5361, new_P3_U5362, new_P3_U5363, new_P3_U5364, new_P3_U5365,
    new_P3_U5366, new_P3_U5367, new_P3_U5368, new_P3_U5369, new_P3_U5370,
    new_P3_U5371, new_P3_U5372, new_P3_U5373, new_P3_U5374, new_P3_U5375,
    new_P3_U5376, new_P3_U5377, new_P3_U5378, new_P3_U5379, new_P3_U5380,
    new_P3_U5381, new_P3_U5382, new_P3_U5383, new_P3_U5384, new_P3_U5385,
    new_P3_U5386, new_P3_U5387, new_P3_U5388, new_P3_U5389, new_P3_U5390,
    new_P3_U5391, new_P3_U5392, new_P3_U5393, new_P3_U5394, new_P3_U5395,
    new_P3_U5396, new_P3_U5397, new_P3_U5398, new_P3_U5399, new_P3_U5400,
    new_P3_U5401, new_P3_U5402, new_P3_U5403, new_P3_U5404, new_P3_U5405,
    new_P3_U5406, new_P3_U5407, new_P3_U5408, new_P3_U5409, new_P3_U5410,
    new_P3_U5411, new_P3_U5412, new_P3_U5413, new_P3_U5414, new_P3_U5415,
    new_P3_U5416, new_P3_U5417, new_P3_U5418, new_P3_U5419, new_P3_U5420,
    new_P3_U5421, new_P3_U5422, new_P3_U5423, new_P3_U5424, new_P3_U5425,
    new_P3_U5426, new_P3_U5427, new_P3_U5428, new_P3_U5429, new_P3_U5430,
    new_P3_U5431, new_P3_U5432, new_P3_U5433, new_P3_U5434, new_P3_U5435,
    new_P3_U5436, new_P3_U5437, new_P3_U5438, new_P3_U5439, new_P3_U5440,
    new_P3_U5441, new_P3_U5442, new_P3_U5443, new_P3_U5444, new_P3_U5445,
    new_P3_U5446, new_P3_U5447, new_P3_U5448, new_P3_U5449, new_P3_U5450,
    new_P3_U5451, new_P3_U5452, new_P3_U5453, new_P3_U5454, new_P3_U5455,
    new_P3_U5456, new_P3_U5457, new_P3_U5458, new_P3_U5459, new_P3_U5460,
    new_P3_U5461, new_P3_U5462, new_P3_U5463, new_P3_U5464, new_P3_U5465,
    new_P3_U5466, new_P3_U5467, new_P3_U5468, new_P3_U5469, new_P3_U5470,
    new_P3_U5471, new_P3_U5472, new_P3_U5473, new_P3_U5474, new_P3_U5475,
    new_P3_U5476, new_P3_U5477, new_P3_U5478, new_P3_U5479, new_P3_U5480,
    new_P3_U5481, new_P3_U5482, new_P3_U5483, new_P3_U5484, new_P3_U5485,
    new_P3_U5486, new_P3_U5487, new_P3_U5488, new_P3_U5489, new_P3_U5490,
    new_P3_U5491, new_P3_U5492, new_P3_U5493, new_P3_U5494, new_P3_U5495,
    new_P3_U5496, new_P3_U5497, new_P3_U5498, new_P3_U5499, new_P3_U5500,
    new_P3_U5501, new_P3_U5502, new_P3_U5503, new_P3_U5504, new_P3_U5505,
    new_P3_U5506, new_P3_U5507, new_P3_U5508, new_P3_U5509, new_P3_U5510,
    new_P3_U5511, new_P3_U5512, new_P3_U5513, new_P3_U5514, new_P3_U5515,
    new_P3_U5516, new_P3_U5517, new_P3_U5518, new_P3_U5519, new_P3_U5520,
    new_P3_U5521, new_P3_U5522, new_P3_U5523, new_P3_U5524, new_P3_U5525,
    new_P3_U5526, new_P3_U5527, new_P3_U5528, new_P3_U5529, new_P3_U5530,
    new_P3_U5531, new_P3_U5532, new_P3_U5533, new_P3_U5534, new_P3_U5535,
    new_P3_U5536, new_P3_U5537, new_P3_U5538, new_P3_U5539, new_P3_U5540,
    new_P3_U5541, new_P3_U5542, new_P3_U5543, new_P3_U5544, new_P3_U5545,
    new_P3_U5546, new_P3_U5547, new_P3_U5548, new_P3_U5549, new_P3_U5550,
    new_P3_U5551, new_P3_U5552, new_P3_U5553, new_P3_U5554, new_P3_U5555,
    new_P3_U5556, new_P3_U5557, new_P3_U5558, new_P3_U5559, new_P3_U5560,
    new_P3_U5561, new_P3_U5562, new_P3_U5563, new_P3_U5564, new_P3_U5565,
    new_P3_U5566, new_P3_U5567, new_P3_U5568, new_P3_U5569, new_P3_U5570,
    new_P3_U5571, new_P3_U5572, new_P3_U5573, new_P3_U5574, new_P3_U5575,
    new_P3_U5576, new_P3_U5577, new_P3_U5578, new_P3_U5579, new_P3_U5580,
    new_P3_U5581, new_P3_U5582, new_P3_U5583, new_P3_U5584, new_P3_U5585,
    new_P3_U5586, new_P3_U5587, new_P3_U5588, new_P3_U5589, new_P3_U5590,
    new_P3_U5591, new_P3_U5592, new_P3_U5593, new_P3_U5594, new_P3_U5595,
    new_P3_U5596, new_P3_U5597, new_P3_U5598, new_P3_U5599, new_P3_U5600,
    new_P3_U5601, new_P3_U5602, new_P3_U5603, new_P3_U5604, new_P3_U5605,
    new_P3_U5606, new_P3_U5607, new_P3_U5608, new_P3_U5609, new_P3_U5610,
    new_P3_U5611, new_P3_U5612, new_P3_U5613, new_P3_U5614, new_P3_U5615,
    new_P3_U5616, new_P3_U5617, new_P3_U5618, new_P3_U5619, new_P3_U5620,
    new_P3_U5621, new_P3_U5622, new_P3_U5623, new_P3_U5624, new_P3_U5625,
    new_P3_U5626, new_P3_U5627, new_P3_U5628, new_P3_U5629, new_P3_U5630,
    new_P3_U5631, new_P3_U5632, new_P3_U5633, new_P3_U5634, new_P3_U5635,
    new_P3_U5636, new_P3_U5637, new_P3_U5638, new_P3_U5639, new_P3_U5640,
    new_P3_U5641, new_P3_U5642, new_P3_U5643, new_P3_U5644, new_P3_U5645,
    new_P3_U5646, new_P3_U5647, new_P3_U5648, new_P3_U5649, new_P3_U5650,
    new_P3_U5651, new_P3_U5652, new_P3_U5653, new_P3_U5654, new_P3_U5655,
    new_P3_U5656, new_P3_U5657, new_P3_U5658, new_P3_U5659, new_P3_U5660,
    new_P3_U5661, new_P3_U5662, new_P3_U5663, new_P3_U5664, new_P3_U5665,
    new_P3_U5666, new_P3_U5667, new_P3_U5668, new_P3_U5669, new_P3_U5670,
    new_P3_U5671, new_P3_U5672, new_P3_U5673, new_P3_U5674, new_P3_U5675,
    new_P3_U5676, new_P3_U5677, new_P3_U5678, new_P3_U5679, new_P3_U5680,
    new_P3_U5681, new_P3_U5682, new_P3_U5683, new_P3_U5684, new_P3_U5685,
    new_P3_U5686, new_P3_U5687, new_P3_U5688, new_P3_U5689, new_P3_U5690,
    new_P3_U5691, new_P3_U5692, new_P3_U5693, new_P3_U5694, new_P3_U5695,
    new_P3_U5696, new_P3_U5697, new_P3_U5698, new_P3_U5699, new_P3_U5700,
    new_P3_U5701, new_P3_U5702, new_P3_U5703, new_P3_U5704, new_P3_U5705,
    new_P3_U5706, new_P3_U5707, new_P3_U5708, new_P3_U5709, new_P3_U5710,
    new_P3_U5711, new_P3_U5712, new_P3_U5713, new_P3_U5714, new_P3_U5715,
    new_P3_U5716, new_P3_U5717, new_P3_U5718, new_P3_U5719, new_P3_U5720,
    new_P3_U5721, new_P3_U5722, new_P3_U5723, new_P3_U5724, new_P3_U5725,
    new_P3_U5726, new_P3_U5727, new_P3_U5728, new_P3_U5729, new_P3_U5730,
    new_P3_U5731, new_P3_U5732, new_P3_U5733, new_P3_U5734, new_P3_U5735,
    new_P3_U5736, new_P3_U5737, new_P3_U5738, new_P3_U5739, new_P3_U5740,
    new_P3_U5741, new_P3_U5742, new_P3_U5743, new_P3_U5744, new_P3_U5745,
    new_P3_U5746, new_P3_U5747, new_P3_U5748, new_P3_U5749, new_P3_U5750,
    new_P3_U5751, new_P3_U5752, new_P3_U5753, new_P3_U5754, new_P3_U5755,
    new_P3_U5756, new_P3_U5757, new_P3_U5758, new_P3_U5759, new_P3_U5760,
    new_P3_U5761, new_P3_U5762, new_P3_U5763, new_P3_U5764, new_P3_U5765,
    new_P3_U5766, new_P3_U5767, new_P3_U5768, new_P3_U5769, new_P3_U5770,
    new_P3_U5771, new_P3_U5772, new_P3_U5773, new_P3_U5774, new_P3_U5775,
    new_P3_U5776, new_P3_U5777, new_P3_U5778, new_P3_U5779, new_P3_U5780,
    new_P3_U5781, new_P3_U5782, new_P3_U5783, new_P3_U5784, new_P3_U5785,
    new_P3_U5786, new_P3_U5787, new_P3_U5788, new_P3_U5789, new_P3_U5790,
    new_P3_U5791, new_P3_U5792, new_P3_U5793, new_P3_U5794, new_P3_U5795,
    new_P3_U5796, new_P3_U5797, new_P3_U5798, new_P3_U5799, new_P3_U5800,
    new_P3_U5801, new_P3_U5802, new_P3_U5803, new_P3_U5804, new_P3_U5805,
    new_P3_U5806, new_P3_U5807, new_P3_U5808, new_P3_U5809, new_P3_U5810,
    new_P3_U5811, new_P3_U5812, new_P3_U5813, new_P3_U5814, new_P3_U5815,
    new_P3_U5816, new_P3_U5817, new_P3_U5818, new_P3_U5819, new_P3_U5820,
    new_P3_U5821, new_P3_U5822, new_P3_U5823, new_P3_U5824, new_P3_U5825,
    new_P3_U5826, new_P3_U5827, new_P3_U5828, new_P3_U5829, new_P3_U5830,
    new_P3_U5831, new_P3_U5832, new_P3_U5833, new_P3_U5834, new_P3_U5835,
    new_P3_U5836, new_P3_U5837, new_P3_U5838, new_P3_U5839, new_P3_U5840,
    new_P3_U5841, new_P3_U5842, new_P3_U5843, new_P3_U5844, new_P3_U5845,
    new_P3_U5846, new_P3_U5847, new_P3_U5848, new_P3_U5849, new_P3_U5850,
    new_P3_U5851, new_P3_U5852, new_P3_U5853, new_P3_U5854, new_P3_U5855,
    new_P3_U5856, new_P3_U5857, new_P3_U5858, new_P3_U5859, new_P3_U5860,
    new_P3_U5861, new_P3_U5862, new_P3_U5863, new_P3_U5864, new_P3_U5865,
    new_P3_U5866, new_P3_U5867, new_P3_U5868, new_P3_U5869, new_P3_U5870,
    new_P3_U5871, new_P3_U5872, new_P3_U5873, new_P3_U5874, new_P3_U5875,
    new_P3_U5876, new_P3_U5877, new_P3_U5878, new_P3_U5879, new_P3_U5880,
    new_P3_U5881, new_P3_U5882, new_P3_U5883, new_P3_U5884, new_P3_U5885,
    new_P3_U5886, new_P3_U5887, new_P3_U5888, new_P3_U5889, new_P3_U5890,
    new_P3_U5891, new_P3_U5892, new_P3_U5893, new_P3_U5894, new_P3_U5895,
    new_P3_U5896, new_P3_U5897, new_P3_U5898, new_P3_U5899, new_P3_U5900,
    new_P3_U5901, new_P3_U5902, new_P3_U5903, new_P3_U5904, new_P3_U5905,
    new_P3_U5906, new_P3_U5907, new_P3_U5908, new_P3_U5909, new_P3_U5910,
    new_P3_U5911, new_P3_U5912, new_P3_U5913, new_P3_U5914, new_P3_U5915,
    new_P3_U5916, new_P3_U5917, new_P3_U5918, new_P3_U5919, new_P3_U5920,
    new_P3_U5921, new_P3_U5922, new_P3_U5923, new_P3_U5924, new_P3_U5925,
    new_P3_U5926, new_P3_U5927, new_P3_U5928, new_P3_U5929, new_P3_U5930,
    new_P3_U5931, new_P3_U5932, new_P3_U5933, new_P3_U5934, new_P3_U5935,
    new_P3_U5936, new_P3_U5937, new_P3_U5938, new_P3_U5939, new_P3_U5940,
    new_P3_U5941, new_P3_U5942, new_P3_U5943, new_P3_U5944, new_P3_U5945,
    new_P3_U5946, new_P3_U5947, new_P3_U5948, new_P3_U5949, new_P3_U5950,
    new_P3_U5951, new_P3_U5952, new_P3_U5953, new_P3_U5954, new_P3_U5955,
    new_P3_U5956, new_P3_U5957, new_P3_U5958, new_P3_U5959, new_P3_U5960,
    new_P3_U5961, new_P3_U5962, new_P3_U5963, new_P3_U5964, new_P3_U5965,
    new_P3_U5966, new_P3_U5967, new_P3_U5968, new_P3_U5969, new_P3_U5970,
    new_P3_U5971, new_P3_U5972, new_P3_U5973, new_P3_U5974, new_P3_U5975,
    new_P3_U5976, new_P3_U5977, new_P3_U5978, new_P3_U5979, new_P3_U5980,
    new_P3_U5981, new_P3_U5982, new_P3_U5983, new_P3_U5984, new_P3_U5985,
    new_P3_U5986, new_P3_U5987, new_P3_U5988, new_P3_U5989, new_P3_U5990,
    new_P3_U5991, new_P3_U5992, new_P3_U5993, new_P3_U5994, new_P3_U5995,
    new_P3_U5996, new_P3_U5997, new_P3_U5998, new_P3_U5999, new_P3_U6000,
    new_P3_U6001, new_P3_U6002, new_P3_U6003, new_P3_U6004, new_P3_U6005,
    new_P3_U6006, new_P3_U6007, new_P3_U6008, new_P3_U6009, new_P3_U6010,
    new_P3_U6011, new_P3_U6012, new_P3_U6013, new_P3_U6014, new_P3_U6015,
    new_P3_U6016, new_P3_U6017, new_P3_U6018, new_P3_U6019, new_P3_U6020,
    new_P3_U6021, new_P3_U6022, new_P3_U6023, new_P3_U6024, new_P3_U6025,
    new_P3_U6026, new_P3_U6027, new_P3_U6028, new_P3_U6029, new_P3_U6030,
    new_P3_U6031, new_P3_U6032, new_P3_U6033, new_P3_U6034, new_P3_U6035,
    new_P3_U6036, new_P3_U6037, new_P3_U6038, new_P3_U6039, new_P3_U6040,
    new_P3_U6041, new_P3_U6042, new_P3_U6043, new_P3_U6044, new_P3_U6045,
    new_P3_U6046, new_P3_U6047, new_P3_U6048, new_P3_U6049, new_P3_U6050,
    new_P3_U6051, new_P3_U6052, new_P3_U6053, new_P3_U6054, new_P3_U6055,
    new_P3_U6056, new_P3_U6057, new_P3_U6058, new_P3_U6059, new_P3_U6060,
    new_P3_U6061, new_P3_U6062, new_P3_U6063, new_P3_U6064, new_P3_U6065,
    new_P3_U6066, new_P3_U6067, new_P3_U6068, new_P3_U6069, new_P3_U6070,
    new_P3_U6071, new_P3_U6072, new_P3_U6073, new_P3_U6074, new_P3_U6075,
    new_P3_U6076, new_P3_U6077, new_P3_U6078, new_P3_U6079, new_P3_U6080,
    new_P3_U6081, new_P3_U6082, new_P3_U6083, new_P3_U6084, new_P3_U6085,
    new_P3_U6086, new_P3_U6087, new_P3_U6088, new_P3_U6089, new_P3_U6090,
    new_P3_U6091, new_P3_U6092, new_P3_U6093, new_P3_U6094, new_P3_U6095,
    new_P3_U6096, new_P3_U6097, new_P3_U6098, new_P3_U6099, new_P3_U6100,
    new_P3_U6101, new_P3_U6102, new_P3_U6103, new_P3_U6104, new_P3_U6105,
    new_P3_U6106, new_P3_U6107, new_P3_U6108, new_P3_U6109, new_P3_U6110,
    new_P3_U6111, new_P3_U6112, new_P3_U6113, new_P3_U6114, new_P3_U6115,
    new_P3_U6116, new_P3_U6117, new_P3_U6118, new_P3_U6119, new_P3_U6120,
    new_P3_U6121, new_P3_U6122, new_P3_U6123, new_P3_U6124, new_P3_U6125,
    new_P3_U6126, new_P3_U6127, new_P3_U6128, new_P3_U6129, new_P3_U6130,
    new_P3_U6131, new_P3_U6132, new_P3_U6133, new_P3_U6134, new_P3_U6135,
    new_P3_U6136, new_P3_U6137, new_P3_U6138, new_P3_U6139, new_P3_U6140,
    new_P3_U6141, new_P3_U6142, new_P3_U6143, new_P3_U6144, new_P3_U6145,
    new_P3_U6146, new_P3_U6147, new_P3_U6148, new_P3_U6149, new_P3_U6150,
    new_P3_U6151, new_P3_U6152, new_P3_U6153, new_P3_U6154, new_P3_U6155,
    new_P3_U6156, new_P3_U6157, new_P3_U6158, new_P3_U6159, new_P3_U6160,
    new_P3_U6161, new_P3_U6162, new_P3_U6163, new_P3_U6164, new_P3_U6165,
    new_P3_U6166, new_P3_U6167, new_P3_U6168, new_P3_U6169, new_P3_U6170,
    new_P3_U6171, new_P3_U6172, new_P3_U6173, new_P3_U6174, new_P3_U6175,
    new_P3_U6176, new_P3_U6177, new_P3_U6178, new_P3_U6179, new_P3_U6180,
    new_P3_U6181, new_P3_U6182, new_P3_U6183, new_P3_U6184, new_P3_U6185,
    new_P3_U6186, new_P3_U6187, new_P3_U6188, new_P3_U6189, new_P3_U6190,
    new_P3_U6191, new_P3_U6192, new_P3_U6193, new_P3_U6194, new_P3_U6195,
    new_P3_U6196, new_P3_U6197, new_P3_U6198, new_P3_U6199, new_P3_U6200,
    new_P3_U6201, new_P3_U6202, new_P3_U6203, new_P3_U6204, new_P3_U6205,
    new_P3_U6206, new_P3_U6207, new_P3_U6208, new_P3_U6209, new_P3_U6210,
    new_P3_U6211, new_P3_U6212, new_P3_U6213, new_P3_U6214, new_P3_U6215,
    new_P3_U6216, new_P3_U6217, new_P3_U6218, new_P3_U6219, new_P3_U6220,
    new_P3_U6221, new_P3_U6222, new_P3_U6223, new_P3_U6224, new_P3_U6225,
    new_P3_U6226, new_P3_U6227, new_P3_U6228, new_P3_U6229, new_P3_U6230,
    new_P3_U6231, new_P3_U6232, new_P3_U6233, new_P3_U6234, new_P3_U6235,
    new_P3_U6236, new_P3_U6237, new_P3_U6238, new_P3_U6239, new_P3_U6240,
    new_P3_U6241, new_P3_U6242, new_P3_U6243, new_P3_U6244, new_P3_U6245,
    new_P3_U6246, new_P3_U6247, new_P3_U6248, new_P3_U6249, new_P3_U6250,
    new_P3_U6251, new_P3_U6252, new_P3_U6253, new_P3_U6254, new_P3_U6255,
    new_P3_U6256, new_P3_U6257, new_P3_U6258, new_P3_U6259, new_P3_U6260,
    new_P3_U6261, new_P3_U6262, new_P3_U6263, new_P3_U6264, new_P3_U6265,
    new_P3_U6266, new_P3_U6267, new_P3_U6268, new_P3_U6269, new_P3_U6270,
    new_P3_U6271, new_P3_U6272, new_P3_U6273, new_P3_U6274, new_P3_U6275,
    new_P3_U6276, new_P3_U6277, new_P3_U6278, new_P3_U6279, new_P3_U6280,
    new_P3_U6281, new_P3_U6282, new_P3_U6283, new_P3_U6284, new_P3_U6285,
    new_P3_U6286, new_P3_U6287, new_P3_U6288, new_P3_U6289, new_P3_U6290,
    new_P3_U6291, new_P3_U6292, new_P3_U6293, new_P3_U6294, new_P3_U6295,
    new_P3_U6296, new_P3_U6297, new_P3_U6298, new_P3_U6299, new_P3_U6300,
    new_P3_U6301, new_P3_U6302, new_P3_U6303, new_P3_U6304, new_P3_U6305,
    new_P3_U6306, new_P3_U6307, new_P3_U6308, new_P3_U6309, new_P3_U6310,
    new_P3_U6311, new_P3_U6312, new_P3_U6313, new_P3_U6314, new_P3_U6315,
    new_P3_U6316, new_P3_U6317, new_P3_U6318, new_P3_U6319, new_P3_U6320,
    new_P3_U6321, new_P3_U6322, new_P3_U6323, new_P3_U6324, new_P3_U6325,
    new_P3_U6326, new_P3_U6327, new_P3_U6328, new_P3_U6329, new_P3_U6330,
    new_P3_U6331, new_P3_U6332, new_P3_U6333, new_P3_U6334, new_P3_U6335,
    new_P3_U6336, new_P3_U6337, new_P3_U6338, new_P3_U6339, new_P3_U6340,
    new_P3_U6341, new_P3_U6342, new_P3_U6343, new_P3_U6344, new_P3_U6345,
    new_P3_U6346, new_P3_U6347, new_P3_U6348, new_P3_U6349, new_P3_U6350,
    new_P3_U6351, new_P3_U6352, new_P3_U6353, new_P3_U6354, new_P3_U6355,
    new_P3_U6356, new_P3_U6357, new_P3_U6358, new_P3_U6359, new_P3_U6360,
    new_P3_U6361, new_P3_U6362, new_P3_U6363, new_P3_U6364, new_P3_U6365,
    new_P3_U6366, new_P3_U6367, new_P3_U6368, new_P3_U6369, new_P3_U6370,
    new_P3_U6371, new_P3_U6372, new_P3_U6373, new_P3_U6374, new_P3_U6375,
    new_P3_U6376, new_P3_U6377, new_P3_U6378, new_P3_U6379, new_P3_U6380,
    new_P3_U6381, new_P3_U6382, new_P3_U6383, new_P3_U6384, new_P3_U6385,
    new_P3_U6386, new_P3_U6387, new_P3_U6388, new_P3_U6389, new_P3_U6390,
    new_P3_U6391, new_P3_U6392, new_P3_U6393, new_P3_U6394, new_P3_U6395,
    new_P3_U6396, new_P3_U6397, new_P3_U6398, new_P3_U6399, new_P3_U6400,
    new_P3_U6401, new_P3_U6402, new_P3_U6403, new_P3_U6404, new_P3_U6405,
    new_P3_U6406, new_P3_U6407, new_P3_U6408, new_P3_U6409, new_P3_U6410,
    new_P3_U6411, new_P3_U6412, new_P3_U6413, new_P3_U6414, new_P3_U6415,
    new_P3_U6416, new_P3_U6417, new_P3_U6418, new_P3_U6419, new_P3_U6420,
    new_P3_U6421, new_P3_U6422, new_P3_U6423, new_P3_U6424, new_P3_U6425,
    new_P3_U6426, new_P3_U6427, new_P3_U6428, new_P3_U6429, new_P3_U6430,
    new_P3_U6431, new_P3_U6432, new_P3_U6433, new_P3_U6434, new_P3_U6435,
    new_P3_U6436, new_P3_U6437, new_P3_U6438, new_P3_U6439, new_P3_U6440,
    new_P3_U6441, new_P3_U6442, new_P3_U6443, new_P3_U6444, new_P3_U6445,
    new_P3_U6446, new_P3_U6447, new_P3_U6448, new_P3_U6449, new_P3_U6450,
    new_P3_U6451, new_P3_U6452, new_P3_U6453, new_P3_U6454, new_P3_U6455,
    new_P3_U6456, new_P3_U6457, new_P3_U6458, new_P3_U6459, new_P3_U6460,
    new_P3_U6461, new_P3_U6462, new_P3_U6463, new_P3_U6464, new_P3_U6465,
    new_P3_U6466, new_P3_U6467, new_P3_U6468, new_P3_U6469, new_P3_U6470,
    new_P3_U6471, new_P3_U6472, new_P3_U6473, new_P3_U6474, new_P3_U6475,
    new_P3_U6476, new_P3_U6477, new_P3_U6478, new_P3_U6479, new_P3_U6480,
    new_P3_U6481, new_P3_U6482, new_P3_U6483, new_P3_U6484, new_P3_U6485,
    new_P3_U6486, new_P3_U6487, new_P3_U6488, new_P3_U6489, new_P3_U6490,
    new_P3_U6491, new_P3_U6492, new_P3_U6493, new_P3_U6494, new_P3_U6495,
    new_P3_U6496, new_P3_U6497, new_P3_U6498, new_P3_U6499, new_P3_U6500,
    new_P3_U6501, new_P3_U6502, new_P3_U6503, new_P3_U6504, new_P3_U6505,
    new_P3_U6506, new_P3_U6507, new_P3_U6508, new_P3_U6509, new_P3_U6510,
    new_P3_U6511, new_P3_U6512, new_P3_U6513, new_P3_U6514, new_P3_U6515,
    new_P3_U6516, new_P3_U6517, new_P3_U6518, new_P3_U6519, new_P3_U6520,
    new_P3_U6521, new_P3_U6522, new_P3_U6523, new_P3_U6524, new_P3_U6525,
    new_P3_U6526, new_P3_U6527, new_P3_U6528, new_P3_U6529, new_P3_U6530,
    new_P3_U6531, new_P3_U6532, new_P3_U6533, new_P3_U6534, new_P3_U6535,
    new_P3_U6536, new_P3_U6537, new_P3_U6538, new_P3_U6539, new_P3_U6540,
    new_P3_U6541, new_P3_U6542, new_P3_U6543, new_P3_U6544, new_P3_U6545,
    new_P3_U6546, new_P3_U6547, new_P3_U6548, new_P3_U6549, new_P3_U6550,
    new_P3_U6551, new_P3_U6552, new_P3_U6553, new_P3_U6554, new_P3_U6555,
    new_P3_U6556, new_P3_U6557, new_P3_U6558, new_P3_U6559, new_P3_U6560,
    new_P3_U6561, new_P3_U6562, new_P3_U6563, new_P3_U6564, new_P3_U6565,
    new_P3_U6566, new_P3_U6567, new_P3_U6568, new_P3_U6569, new_P3_U6570,
    new_P3_U6571, new_P3_U6572, new_P3_U6573, new_P3_U6574, new_P3_U6575,
    new_P3_U6576, new_P3_U6577, new_P3_U6578, new_P3_U6579, new_P3_U6580,
    new_P3_U6581, new_P3_U6582, new_P3_U6583, new_P3_U6584, new_P3_U6585,
    new_P3_U6586, new_P3_U6587, new_P3_U6588, new_P3_U6589, new_P3_U6590,
    new_P3_U6591, new_P3_U6592, new_P3_U6593, new_P3_U6594, new_P3_U6595,
    new_P3_U6596, new_P3_U6597, new_P3_U6598, new_P3_U6599, new_P3_U6600,
    new_P3_U6601, new_P3_U6602, new_P3_U6603, new_P3_U6604, new_P3_U6605,
    new_P3_U6606, new_P3_U6607, new_P3_U6608, new_P3_U6609, new_P3_U6610,
    new_P3_U6611, new_P3_U6612, new_P3_U6613, new_P3_U6614, new_P3_U6615,
    new_P3_U6616, new_P3_U6617, new_P3_U6618, new_P3_U6619, new_P3_U6620,
    new_P3_U6621, new_P3_U6622, new_P3_U6623, new_P3_U6624, new_P3_U6625,
    new_P3_U6626, new_P3_U6627, new_P3_U6628, new_P3_U6629, new_P3_U6630,
    new_P3_U6631, new_P3_U6632, new_P3_U6633, new_P3_U6634, new_P3_U6635,
    new_P3_U6636, new_P3_U6637, new_P3_U6638, new_P3_U6639, new_P3_U6640,
    new_P3_U6641, new_P3_U6642, new_P3_U6643, new_P3_U6644, new_P3_U6645,
    new_P3_U6646, new_P3_U6647, new_P3_U6648, new_P3_U6649, new_P3_U6650,
    new_P3_U6651, new_P3_U6652, new_P3_U6653, new_P3_U6654, new_P3_U6655,
    new_P3_U6656, new_P3_U6657, new_P3_U6658, new_P3_U6659, new_P3_U6660,
    new_P3_U6661, new_P3_U6662, new_P3_U6663, new_P3_U6664, new_P3_U6665,
    new_P3_U6666, new_P3_U6667, new_P3_U6668, new_P3_U6669, new_P3_U6670,
    new_P3_U6671, new_P3_U6672, new_P3_U6673, new_P3_U6674, new_P3_U6675,
    new_P3_U6676, new_P3_U6677, new_P3_U6678, new_P3_U6679, new_P3_U6680,
    new_P3_U6681, new_P3_U6682, new_P3_U6683, new_P3_U6684, new_P3_U6685,
    new_P3_U6686, new_P3_U6687, new_P3_U6688, new_P3_U6689, new_P3_U6690,
    new_P3_U6691, new_P3_U6692, new_P3_U6693, new_P3_U6694, new_P3_U6695,
    new_P3_U6696, new_P3_U6697, new_P3_U6698, new_P3_U6699, new_P3_U6700,
    new_P3_U6701, new_P3_U6702, new_P3_U6703, new_P3_U6704, new_P3_U6705,
    new_P3_U6706, new_P3_U6707, new_P3_U6708, new_P3_U6709, new_P3_U6710,
    new_P3_U6711, new_P3_U6712, new_P3_U6713, new_P3_U6714, new_P3_U6715,
    new_P3_U6716, new_P3_U6717, new_P3_U6718, new_P3_U6719, new_P3_U6720,
    new_P3_U6721, new_P3_U6722, new_P3_U6723, new_P3_U6724, new_P3_U6725,
    new_P3_U6726, new_P3_U6727, new_P3_U6728, new_P3_U6729, new_P3_U6730,
    new_P3_U6731, new_P3_U6732, new_P3_U6733, new_P3_U6734, new_P3_U6735,
    new_P3_U6736, new_P3_U6737, new_P3_U6738, new_P3_U6739, new_P3_U6740,
    new_P3_U6741, new_P3_U6742, new_P3_U6743, new_P3_U6744, new_P3_U6745,
    new_P3_U6746, new_P3_U6747, new_P3_U6748, new_P3_U6749, new_P3_U6750,
    new_P3_U6751, new_P3_U6752, new_P3_U6753, new_P3_U6754, new_P3_U6755,
    new_P3_U6756, new_P3_U6757, new_P3_U6758, new_P3_U6759, new_P3_U6760,
    new_P3_U6761, new_P3_U6762, new_P3_U6763, new_P3_U6764, new_P3_U6765,
    new_P3_U6766, new_P3_U6767, new_P3_U6768, new_P3_U6769, new_P3_U6770,
    new_P3_U6771, new_P3_U6772, new_P3_U6773, new_P3_U6774, new_P3_U6775,
    new_P3_U6776, new_P3_U6777, new_P3_U6778, new_P3_U6779, new_P3_U6780,
    new_P3_U6781, new_P3_U6782, new_P3_U6783, new_P3_U6784, new_P3_U6785,
    new_P3_U6786, new_P3_U6787, new_P3_U6788, new_P3_U6789, new_P3_U6790,
    new_P3_U6791, new_P3_U6792, new_P3_U6793, new_P3_U6794, new_P3_U6795,
    new_P3_U6796, new_P3_U6797, new_P3_U6798, new_P3_U6799, new_P3_U6800,
    new_P3_U6801, new_P3_U6802, new_P3_U6803, new_P3_U6804, new_P3_U6805,
    new_P3_U6806, new_P3_U6807, new_P3_U6808, new_P3_U6809, new_P3_U6810,
    new_P3_U6811, new_P3_U6812, new_P3_U6813, new_P3_U6814, new_P3_U6815,
    new_P3_U6816, new_P3_U6817, new_P3_U6818, new_P3_U6819, new_P3_U6820,
    new_P3_U6821, new_P3_U6822, new_P3_U6823, new_P3_U6824, new_P3_U6825,
    new_P3_U6826, new_P3_U6827, new_P3_U6828, new_P3_U6829, new_P3_U6830,
    new_P3_U6831, new_P3_U6832, new_P3_U6833, new_P3_U6834, new_P3_U6835,
    new_P3_U6836, new_P3_U6837, new_P3_U6838, new_P3_U6839, new_P3_U6840,
    new_P3_U6841, new_P3_U6842, new_P3_U6843, new_P3_U6844, new_P3_U6845,
    new_P3_U6846, new_P3_U6847, new_P3_U6848, new_P3_U6849, new_P3_U6850,
    new_P3_U6851, new_P3_U6852, new_P3_U6853, new_P3_U6854, new_P3_U6855,
    new_P3_U6856, new_P3_U6857, new_P3_U6858, new_P3_U6859, new_P3_U6860,
    new_P3_U6861, new_P3_U6862, new_P3_U6863, new_P3_U6864, new_P3_U6865,
    new_P3_U6866, new_P3_U6867, new_P3_U6868, new_P3_U6869, new_P3_U6870,
    new_P3_U6871, new_P3_U6872, new_P3_U6873, new_P3_U6874, new_P3_U6875,
    new_P3_U6876, new_P3_U6877, new_P3_U6878, new_P3_U6879, new_P3_U6880,
    new_P3_U6881, new_P3_U6882, new_P3_U6883, new_P3_U6884, new_P3_U6885,
    new_P3_U6886, new_P3_U6887, new_P3_U6888, new_P3_U6889, new_P3_U6890,
    new_P3_U6891, new_P3_U6892, new_P3_U6893, new_P3_U6894, new_P3_U6895,
    new_P3_U6896, new_P3_U6897, new_P3_U6898, new_P3_U6899, new_P3_U6900,
    new_P3_U6901, new_P3_U6902, new_P3_U6903, new_P3_U6904, new_P3_U6905,
    new_P3_U6906, new_P3_U6907, new_P3_U6908, new_P3_U6909, new_P3_U6910,
    new_P3_U6911, new_P3_U6912, new_P3_U6913, new_P3_U6914, new_P3_U6915,
    new_P3_U6916, new_P3_U6917, new_P3_U6918, new_P3_U6919, new_P3_U6920,
    new_P3_U6921, new_P3_U6922, new_P3_U6923, new_P3_U6924, new_P3_U6925,
    new_P3_U6926, new_P3_U6927, new_P3_U6928, new_P3_U6929, new_P3_U6930,
    new_P3_U6931, new_P3_U6932, new_P3_U6933, new_P3_U6934, new_P3_U6935,
    new_P3_U6936, new_P3_U6937, new_P3_U6938, new_P3_U6939, new_P3_U6940,
    new_P3_U6941, new_P3_U6942, new_P3_U6943, new_P3_U6944, new_P3_U6945,
    new_P3_U6946, new_P3_U6947, new_P3_U6948, new_P3_U6949, new_P3_U6950,
    new_P3_U6951, new_P3_U6952, new_P3_U6953, new_P3_U6954, new_P3_U6955,
    new_P3_U6956, new_P3_U6957, new_P3_U6958, new_P3_U6959, new_P3_U6960,
    new_P3_U6961, new_P3_U6962, new_P3_U6963, new_P3_U6964, new_P3_U6965,
    new_P3_U6966, new_P3_U6967, new_P3_U6968, new_P3_U6969, new_P3_U6970,
    new_P3_U6971, new_P3_U6972, new_P3_U6973, new_P3_U6974, new_P3_U6975,
    new_P3_U6976, new_P3_U6977, new_P3_U6978, new_P3_U6979, new_P3_U6980,
    new_P3_U6981, new_P3_U6982, new_P3_U6983, new_P3_U6984, new_P3_U6985,
    new_P3_U6986, new_P3_U6987, new_P3_U6988, new_P3_U6989, new_P3_U6990,
    new_P3_U6991, new_P3_U6992, new_P3_U6993, new_P3_U6994, new_P3_U6995,
    new_P3_U6996, new_P3_U6997, new_P3_U6998, new_P3_U6999, new_P3_U7000,
    new_P3_U7001, new_P3_U7002, new_P3_U7003, new_P3_U7004, new_P3_U7005,
    new_P3_U7006, new_P3_U7007, new_P3_U7008, new_P3_U7009, new_P3_U7010,
    new_P3_U7011, new_P3_U7012, new_P3_U7013, new_P3_U7014, new_P3_U7015,
    new_P3_U7016, new_P3_U7017, new_P3_U7018, new_P3_U7019, new_P3_U7020,
    new_P3_U7021, new_P3_U7022, new_P3_U7023, new_P3_U7024, new_P3_U7025,
    new_P3_U7026, new_P3_U7027, new_P3_U7028, new_P3_U7029, new_P3_U7030,
    new_P3_U7031, new_P3_U7032, new_P3_U7033, new_P3_U7034, new_P3_U7035,
    new_P3_U7036, new_P3_U7037, new_P3_U7038, new_P3_U7039, new_P3_U7040,
    new_P3_U7041, new_P3_U7042, new_P3_U7043, new_P3_U7044, new_P3_U7045,
    new_P3_U7046, new_P3_U7047, new_P3_U7048, new_P3_U7049, new_P3_U7050,
    new_P3_U7051, new_P3_U7052, new_P3_U7053, new_P3_U7054, new_P3_U7055,
    new_P3_U7056, new_P3_U7057, new_P3_U7058, new_P3_U7059, new_P3_U7060,
    new_P3_U7061, new_P3_U7062, new_P3_U7063, new_P3_U7064, new_P3_U7065,
    new_P3_U7066, new_P3_U7067, new_P3_U7068, new_P3_U7069, new_P3_U7070,
    new_P3_U7071, new_P3_U7072, new_P3_U7073, new_P3_U7074, new_P3_U7075,
    new_P3_U7076, new_P3_U7077, new_P3_U7078, new_P3_U7079, new_P3_U7080,
    new_P3_U7081, new_P3_U7082, new_P3_U7083, new_P3_U7084, new_P3_U7085,
    new_P3_U7086, new_P3_U7087, new_P3_U7088, new_P3_U7089, new_P3_U7090,
    new_P3_U7091, new_P3_U7092, new_P3_U7093, new_P3_U7094, new_P3_U7095,
    new_P3_U7096, new_P3_U7097, new_P3_U7098, new_P3_U7099, new_P3_U7100,
    new_P3_U7101, new_P3_U7102, new_P3_U7103, new_P3_U7104, new_P3_U7105,
    new_P3_U7106, new_P3_U7107, new_P3_U7108, new_P3_U7109, new_P3_U7110,
    new_P3_U7111, new_P3_U7112, new_P3_U7113, new_P3_U7114, new_P3_U7115,
    new_P3_U7116, new_P3_U7117, new_P3_U7118, new_P3_U7119, new_P3_U7120,
    new_P3_U7121, new_P3_U7122, new_P3_U7123, new_P3_U7124, new_P3_U7125,
    new_P3_U7126, new_P3_U7127, new_P3_U7128, new_P3_U7129, new_P3_U7130,
    new_P3_U7131, new_P3_U7132, new_P3_U7133, new_P3_U7134, new_P3_U7135,
    new_P3_U7136, new_P3_U7137, new_P3_U7138, new_P3_U7139, new_P3_U7140,
    new_P3_U7141, new_P3_U7142, new_P3_U7143, new_P3_U7144, new_P3_U7145,
    new_P3_U7146, new_P3_U7147, new_P3_U7148, new_P3_U7149, new_P3_U7150,
    new_P3_U7151, new_P3_U7152, new_P3_U7153, new_P3_U7154, new_P3_U7155,
    new_P3_U7156, new_P3_U7157, new_P3_U7158, new_P3_U7159, new_P3_U7160,
    new_P3_U7161, new_P3_U7162, new_P3_U7163, new_P3_U7164, new_P3_U7165,
    new_P3_U7166, new_P3_U7167, new_P3_U7168, new_P3_U7169, new_P3_U7170,
    new_P3_U7171, new_P3_U7172, new_P3_U7173, new_P3_U7174, new_P3_U7175,
    new_P3_U7176, new_P3_U7177, new_P3_U7178, new_P3_U7179, new_P3_U7180,
    new_P3_U7181, new_P3_U7182, new_P3_U7183, new_P3_U7184, new_P3_U7185,
    new_P3_U7186, new_P3_U7187, new_P3_U7188, new_P3_U7189, new_P3_U7190,
    new_P3_U7191, new_P3_U7192, new_P3_U7193, new_P3_U7194, new_P3_U7195,
    new_P3_U7196, new_P3_U7197, new_P3_U7198, new_P3_U7199, new_P3_U7200,
    new_P3_U7201, new_P3_U7202, new_P3_U7203, new_P3_U7204, new_P3_U7205,
    new_P3_U7206, new_P3_U7207, new_P3_U7208, new_P3_U7209, new_P3_U7210,
    new_P3_U7211, new_P3_U7212, new_P3_U7213, new_P3_U7214, new_P3_U7215,
    new_P3_U7216, new_P3_U7217, new_P3_U7218, new_P3_U7219, new_P3_U7220,
    new_P3_U7221, new_P3_U7222, new_P3_U7223, new_P3_U7224, new_P3_U7225,
    new_P3_U7226, new_P3_U7227, new_P3_U7228, new_P3_U7229, new_P3_U7230,
    new_P3_U7231, new_P3_U7232, new_P3_U7233, new_P3_U7234, new_P3_U7235,
    new_P3_U7236, new_P3_U7237, new_P3_U7238, new_P3_U7239, new_P3_U7240,
    new_P3_U7241, new_P3_U7242, new_P3_U7243, new_P3_U7244, new_P3_U7245,
    new_P3_U7246, new_P3_U7247, new_P3_U7248, new_P3_U7249, new_P3_U7250,
    new_P3_U7251, new_P3_U7252, new_P3_U7253, new_P3_U7254, new_P3_U7255,
    new_P3_U7256, new_P3_U7257, new_P3_U7258, new_P3_U7259, new_P3_U7260,
    new_P3_U7261, new_P3_U7262, new_P3_U7263, new_P3_U7264, new_P3_U7265,
    new_P3_U7266, new_P3_U7267, new_P3_U7268, new_P3_U7269, new_P3_U7270,
    new_P3_U7271, new_P3_U7272, new_P3_U7273, new_P3_U7274, new_P3_U7275,
    new_P3_U7276, new_P3_U7277, new_P3_U7278, new_P3_U7279, new_P3_U7280,
    new_P3_U7281, new_P3_U7282, new_P3_U7283, new_P3_U7284, new_P3_U7285,
    new_P3_U7286, new_P3_U7287, new_P3_U7288, new_P3_U7289, new_P3_U7290,
    new_P3_U7291, new_P3_U7292, new_P3_U7293, new_P3_U7294, new_P3_U7295,
    new_P3_U7296, new_P3_U7297, new_P3_U7298, new_P3_U7299, new_P3_U7300,
    new_P3_U7301, new_P3_U7302, new_P3_U7303, new_P3_U7304, new_P3_U7305,
    new_P3_U7306, new_P3_U7307, new_P3_U7308, new_P3_U7309, new_P3_U7310,
    new_P3_U7311, new_P3_U7312, new_P3_U7313, new_P3_U7314, new_P3_U7315,
    new_P3_U7316, new_P3_U7317, new_P3_U7318, new_P3_U7319, new_P3_U7320,
    new_P3_U7321, new_P3_U7322, new_P3_U7323, new_P3_U7324, new_P3_U7325,
    new_P3_U7326, new_P3_U7327, new_P3_U7328, new_P3_U7329, new_P3_U7330,
    new_P3_U7331, new_P3_U7332, new_P3_U7333, new_P3_U7334, new_P3_U7335,
    new_P3_U7336, new_P3_U7337, new_P3_U7338, new_P3_U7339, new_P3_U7340,
    new_P3_U7341, new_P3_U7342, new_P3_U7343, new_P3_U7344, new_P3_U7345,
    new_P3_U7346, new_P3_U7347, new_P3_U7348, new_P3_U7349, new_P3_U7350,
    new_P3_U7351, new_P3_U7352, new_P3_U7353, new_P3_U7354, new_P3_U7355,
    new_P3_U7356, new_P3_U7357, new_P3_U7358, new_P3_U7359, new_P3_U7360,
    new_P3_U7361, new_P3_U7362, new_P3_U7363, new_P3_U7364, new_P3_U7365,
    new_P3_U7366, new_P3_U7367, new_P3_U7368, new_P3_U7369, new_P3_U7370,
    new_P3_U7371, new_P3_U7372, new_P3_U7373, new_P3_U7374, new_P3_U7375,
    new_P3_U7376, new_P3_U7377, new_P3_U7378, new_P3_U7379, new_P3_U7380,
    new_P3_U7381, new_P3_U7382, new_P3_U7383, new_P3_U7384, new_P3_U7385,
    new_P3_U7386, new_P3_U7387, new_P3_U7388, new_P3_U7389, new_P3_U7390,
    new_P3_U7391, new_P3_U7392, new_P3_U7393, new_P3_U7394, new_P3_U7395,
    new_P3_U7396, new_P3_U7397, new_P3_U7398, new_P3_U7399, new_P3_U7400,
    new_P3_U7401, new_P3_U7402, new_P3_U7403, new_P3_U7404, new_P3_U7405,
    new_P3_U7406, new_P3_U7407, new_P3_U7408, new_P3_U7409, new_P3_U7410,
    new_P3_U7411, new_P3_U7412, new_P3_U7413, new_P3_U7414, new_P3_U7415,
    new_P3_U7416, new_P3_U7417, new_P3_U7418, new_P3_U7419, new_P3_U7420,
    new_P3_U7421, new_P3_U7422, new_P3_U7423, new_P3_U7424, new_P3_U7425,
    new_P3_U7426, new_P3_U7427, new_P3_U7428, new_P3_U7429, new_P3_U7430,
    new_P3_U7431, new_P3_U7432, new_P3_U7433, new_P3_U7434, new_P3_U7435,
    new_P3_U7436, new_P3_U7437, new_P3_U7438, new_P3_U7439, new_P3_U7440,
    new_P3_U7441, new_P3_U7442, new_P3_U7443, new_P3_U7444, new_P3_U7445,
    new_P3_U7446, new_P3_U7447, new_P3_U7448, new_P3_U7449, new_P3_U7450,
    new_P3_U7451, new_P3_U7452, new_P3_U7453, new_P3_U7454, new_P3_U7455,
    new_P3_U7456, new_P3_U7457, new_P3_U7458, new_P3_U7459, new_P3_U7460,
    new_P3_U7461, new_P3_U7462, new_P3_U7463, new_P3_U7464, new_P3_U7465,
    new_P3_U7466, new_P3_U7467, new_P3_U7468, new_P3_U7469, new_P3_U7470,
    new_P3_U7471, new_P3_U7472, new_P3_U7473, new_P3_U7474, new_P3_U7475,
    new_P3_U7476, new_P3_U7477, new_P3_U7478, new_P3_U7479, new_P3_U7480,
    new_P3_U7481, new_P3_U7482, new_P3_U7483, new_P3_U7484, new_P3_U7485,
    new_P3_U7486, new_P3_U7487, new_P3_U7488, new_P3_U7489, new_P3_U7490,
    new_P3_U7491, new_P3_U7492, new_P3_U7493, new_P3_U7494, new_P3_U7495,
    new_P3_U7496, new_P3_U7497, new_P3_U7498, new_P3_U7499, new_P3_U7500,
    new_P3_U7501, new_P3_U7502, new_P3_U7503, new_P3_U7504, new_P3_U7505,
    new_P3_U7506, new_P3_U7507, new_P3_U7508, new_P3_U7509, new_P3_U7510,
    new_P3_U7511, new_P3_U7512, new_P3_U7513, new_P3_U7514, new_P3_U7515,
    new_P3_U7516, new_P3_U7517, new_P3_U7518, new_P3_U7519, new_P3_U7520,
    new_P3_U7521, new_P3_U7522, new_P3_U7523, new_P3_U7524, new_P3_U7525,
    new_P3_U7526, new_P3_U7527, new_P3_U7528, new_P3_U7529, new_P3_U7530,
    new_P3_U7531, new_P3_U7532, new_P3_U7533, new_P3_U7534, new_P3_U7535,
    new_P3_U7536, new_P3_U7537, new_P3_U7538, new_P3_U7539, new_P3_U7540,
    new_P3_U7541, new_P3_U7542, new_P3_U7543, new_P3_U7544, new_P3_U7545,
    new_P3_U7546, new_P3_U7547, new_P3_U7548, new_P3_U7549, new_P3_U7550,
    new_P3_U7551, new_P3_U7552, new_P3_U7553, new_P3_U7554, new_P3_U7555,
    new_P3_U7556, new_P3_U7557, new_P3_U7558, new_P3_U7559, new_P3_U7560,
    new_P3_U7561, new_P3_U7562, new_P3_U7563, new_P3_U7564, new_P3_U7565,
    new_P3_U7566, new_P3_U7567, new_P3_U7568, new_P3_U7569, new_P3_U7570,
    new_P3_U7571, new_P3_U7572, new_P3_U7573, new_P3_U7574, new_P3_U7575,
    new_P3_U7576, new_P3_U7577, new_P3_U7578, new_P3_U7579, new_P3_U7580,
    new_P3_U7581, new_P3_U7582, new_P3_U7583, new_P3_U7584, new_P3_U7585,
    new_P3_U7586, new_P3_U7587, new_P3_U7588, new_P3_U7589, new_P3_U7590,
    new_P3_U7591, new_P3_U7592, new_P3_U7593, new_P3_U7594, new_P3_U7595,
    new_P3_U7596, new_P3_U7597, new_P3_U7598, new_P3_U7599, new_P3_U7600,
    new_P3_U7601, new_P3_U7602, new_P3_U7603, new_P3_U7604, new_P3_U7605,
    new_P3_U7606, new_P3_U7607, new_P3_U7608, new_P3_U7609, new_P3_U7610,
    new_P3_U7611, new_P3_U7612, new_P3_U7613, new_P3_U7614, new_P3_U7615,
    new_P3_U7616, new_P3_U7617, new_P3_U7618, new_P3_U7619, new_P3_U7620,
    new_P3_U7621, new_P3_U7622, new_P3_U7623, new_P3_U7624, new_P3_U7625,
    new_P3_U7626, new_P3_U7627, new_P3_U7628, new_P3_U7629, new_P3_U7630,
    new_P3_U7631, new_P3_U7632, new_P3_U7633, new_P3_U7634, new_P3_U7635,
    new_P3_U7636, new_P3_U7637, new_P3_U7638, new_P3_U7639, new_P3_U7640,
    new_P3_U7641, new_P3_U7642, new_P3_U7643, new_P3_U7644, new_P3_U7645,
    new_P3_U7646, new_P3_U7647, new_P3_U7648, new_P3_U7649, new_P3_U7650,
    new_P3_U7651, new_P3_U7652, new_P3_U7653, new_P3_U7654, new_P3_U7655,
    new_P3_U7656, new_P3_U7657, new_P3_U7658, new_P3_U7659, new_P3_U7660,
    new_P3_U7661, new_P3_U7662, new_P3_U7663, new_P3_U7664, new_P3_U7665,
    new_P3_U7666, new_P3_U7667, new_P3_U7668, new_P3_U7669, new_P3_U7670,
    new_P3_U7671, new_P3_U7672, new_P3_U7673, new_P3_U7674, new_P3_U7675,
    new_P3_U7676, new_P3_U7677, new_P3_U7678, new_P3_U7679, new_P3_U7680,
    new_P3_U7681, new_P3_U7682, new_P3_U7683, new_P3_U7684, new_P3_U7685,
    new_P3_U7686, new_P3_U7687, new_P3_U7688, new_P3_U7689, new_P3_U7690,
    new_P3_U7691, new_P3_U7692, new_P3_U7693, new_P3_U7694, new_P3_U7695,
    new_P3_U7696, new_P3_U7697, new_P3_U7698, new_P3_U7699, new_P3_U7700,
    new_P3_U7701, new_P3_U7702, new_P3_U7703, new_P3_U7704, new_P3_U7705,
    new_P3_U7706, new_P3_U7707, new_P3_U7708, new_P3_U7709, new_P3_U7710,
    new_P3_U7711, new_P3_U7712, new_P3_U7713, new_P3_U7714, new_P3_U7715,
    new_P3_U7716, new_P3_U7717, new_P3_U7718, new_P3_U7719, new_P3_U7720,
    new_P3_U7721, new_P3_U7722, new_P3_U7723, new_P3_U7724, new_P3_U7725,
    new_P3_U7726, new_P3_U7727, new_P3_U7728, new_P3_U7729, new_P3_U7730,
    new_P3_U7731, new_P3_U7732, new_P3_U7733, new_P3_U7734, new_P3_U7735,
    new_P3_U7736, new_P3_U7737, new_P3_U7738, new_P3_U7739, new_P3_U7740,
    new_P3_U7741, new_P3_U7742, new_P3_U7743, new_P3_U7744, new_P3_U7745,
    new_P3_U7746, new_P3_U7747, new_P3_U7748, new_P3_U7749, new_P3_U7750,
    new_P3_U7751, new_P3_U7752, new_P3_U7753, new_P3_U7754, new_P3_U7755,
    new_P3_U7756, new_P3_U7757, new_P3_U7758, new_P3_U7759, new_P3_U7760,
    new_P3_U7761, new_P3_U7762, new_P3_U7763, new_P3_U7764, new_P3_U7765,
    new_P3_U7766, new_P3_U7767, new_P3_U7768, new_P3_U7769, new_P3_U7770,
    new_P3_U7771, new_P3_U7772, new_P3_U7773, new_P3_U7774, new_P3_U7775,
    new_P3_U7776, new_P3_U7777, new_P3_U7778, new_P3_U7779, new_P3_U7780,
    new_P3_U7781, new_P3_U7782, new_P3_U7783, new_P3_U7784, new_P3_U7785,
    new_P3_U7786, new_P3_U7787, new_P3_U7788, new_P3_U7789, new_P3_U7790,
    new_P3_U7791, new_P3_U7792, new_P3_U7793, new_P3_U7794, new_P3_U7795,
    new_P3_U7796, new_P3_U7797, new_P3_U7798, new_P3_U7799, new_P3_U7800,
    new_P3_U7801, new_P3_U7802, new_P3_U7803, new_P3_U7804, new_P3_U7805,
    new_P3_U7806, new_P3_U7807, new_P3_U7808, new_P3_U7809, new_P3_U7810,
    new_P3_U7811, new_P3_U7812, new_P3_U7813, new_P3_U7814, new_P3_U7815,
    new_P3_U7816, new_P3_U7817, new_P3_U7818, new_P3_U7819, new_P3_U7820,
    new_P3_U7821, new_P3_U7822, new_P3_U7823, new_P3_U7824, new_P3_U7825,
    new_P3_U7826, new_P3_U7827, new_P3_U7828, new_P3_U7829, new_P3_U7830,
    new_P3_U7831, new_P3_U7832, new_P3_U7833, new_P3_U7834, new_P3_U7835,
    new_P3_U7836, new_P3_U7837, new_P3_U7838, new_P3_U7839, new_P3_U7840,
    new_P3_U7841, new_P3_U7842, new_P3_U7843, new_P3_U7844, new_P3_U7845,
    new_P3_U7846, new_P3_U7847, new_P3_U7848, new_P3_U7849, new_P3_U7850,
    new_P3_U7851, new_P3_U7852, new_P3_U7853, new_P3_U7854, new_P3_U7855,
    new_P3_U7856, new_P3_U7857, new_P3_U7858, new_P3_U7859, new_P3_U7860,
    new_P3_U7861, new_P3_U7862, new_P3_U7863, new_P3_U7864, new_P3_U7865,
    new_P3_U7866, new_P3_U7867, new_P3_U7868, new_P3_U7869, new_P3_U7870,
    new_P3_U7871, new_P3_U7872, new_P3_U7873, new_P3_U7874, new_P3_U7875,
    new_P3_U7876, new_P3_U7877, new_P3_U7878, new_P3_U7879, new_P3_U7880,
    new_P3_U7881, new_P3_U7882, new_P3_U7883, new_P3_U7884, new_P3_U7885,
    new_P3_U7886, new_P3_U7887, new_P3_U7888, new_P3_U7889, new_P3_U7890,
    new_P3_U7891, new_P3_U7892, new_P3_U7893, new_P3_U7894, new_P3_U7895,
    new_P3_U7896, new_P3_U7897, new_P3_U7898, new_P3_U7899, new_P3_U7900,
    new_P3_U7901, new_P3_U7902, new_P3_U7903, new_P3_U7904, new_P3_U7905,
    new_P3_U7906, new_P3_U7907, new_P3_U7908, new_P3_U7909, new_P3_U7910,
    new_P3_U7911, new_P3_U7912, new_P3_U7913, new_P3_U7914, new_P3_U7915,
    new_P3_U7916, new_P3_U7917, new_P3_U7918, new_P3_U7919, new_P3_U7920,
    new_P3_U7921, new_P3_U7922, new_P3_U7923, new_P3_U7924, new_P3_U7925,
    new_P3_U7926, new_P3_U7927, new_P3_U7928, new_P3_U7929, new_P3_U7930,
    new_P3_U7931, new_P3_U7932, new_P3_U7933, new_P3_U7934, new_P3_U7935,
    new_P3_U7936, new_P3_U7937, new_P3_U7938, new_P3_U7939, new_P3_U7940,
    new_P3_U7941, new_P3_U7942, new_P3_U7943, new_P3_U7944, new_P3_U7945,
    new_P3_U7946, new_P3_U7947, new_P3_U7948, new_P3_U7949, new_P3_U7950,
    new_P3_U7951, new_P3_U7952, new_P3_U7953, new_P3_U7954, new_P3_U7955,
    new_P3_U7956, new_P3_U7957, new_P3_U7958, new_P3_U7959, new_P3_U7960,
    new_P3_U7961, new_P3_U7962, new_P3_U7963, new_P3_U7964, new_P3_U7965,
    new_P3_U7966, new_P3_U7967, new_P3_U7968, new_P3_U7969, new_P3_U7970,
    new_P3_U7971, new_P3_U7972, new_P3_U7973, new_P3_U7974, new_P3_U7975,
    new_P3_U7976, new_P3_U7977, new_P3_U7978, new_P3_U7979, new_P3_U7980,
    new_P3_U7981, new_P3_U7982, new_P3_U7983, new_P3_U7984, new_P3_U7985,
    new_P3_U7986, new_P3_U7987, new_P3_U7988, new_P3_U7989, new_P3_U7990,
    new_P3_U7991, new_P3_U7992, new_P3_U7993, new_P3_U7994, new_P3_U7995,
    new_P3_U7996, new_P3_U7997, new_P3_U7998, new_P3_U7999, new_P3_U8000,
    new_P3_U8001, new_P3_U8002, new_P3_U8003, new_P3_U8004, new_P3_U8005,
    new_P3_U8006, new_P3_U8007, new_P3_U8008, new_P3_U8009, new_P3_U8010,
    new_P3_U8011, new_P3_U8012, new_P3_U8013, new_P3_U8014, new_P3_U8015,
    new_P3_U8016, new_P3_U8017, new_P3_U8018, new_P3_U8019, new_P3_U8020,
    new_P3_U8021, new_P3_U8022, new_P3_U8023, new_P3_U8024, new_P3_U8025,
    new_P3_U8026, new_P3_U8027, new_P3_U8028, new_P3_U8029, new_P3_U8030,
    new_P3_U8031, new_P3_U8032, new_P3_U8033, new_P3_U8034, new_P3_U8035,
    new_P3_U8036, new_P3_U8037, new_P3_U8038, new_P3_U8039, new_P3_U8040,
    new_P3_U8041, new_P3_U8042, new_P3_U8043, new_P3_U8044, new_P3_U8045,
    new_P3_U8046, new_P3_U8047, new_P3_U8048, new_P3_U8049, new_P3_U8050,
    new_P3_U8051, new_P3_U8052, new_P3_U8053, new_P1_ADD_515_U170,
    new_P1_ADD_515_U169, new_P1_ADD_515_U168, new_P1_ADD_515_U167,
    new_P1_ADD_515_U166, new_P1_ADD_515_U165, new_P1_ADD_515_U164,
    new_P1_ADD_515_U163, new_P1_ADD_515_U162, new_P1_ADD_515_U161,
    new_P1_ADD_515_U160, new_P1_ADD_515_U159, new_P1_ADD_515_U158,
    new_P1_ADD_515_U157, new_P1_ADD_515_U156, new_P1_ADD_515_U155,
    new_P1_ADD_515_U154, new_P1_ADD_515_U153, new_P1_ADD_515_U152,
    new_P1_ADD_515_U151, new_P1_ADD_515_U150, new_P1_ADD_515_U149,
    new_P1_ADD_515_U148, new_P1_ADD_515_U147, new_P1_ADD_515_U146,
    new_P1_ADD_515_U145, new_P1_ADD_515_U144, new_P1_ADD_515_U143,
    new_P1_ADD_515_U142, new_P1_ADD_515_U141, new_P1_ADD_515_U140,
    new_P1_ADD_515_U139, new_P1_ADD_515_U138, new_P1_ADD_515_U137,
    new_P1_ADD_515_U136, new_P1_ADD_515_U135, new_P1_ADD_515_U134,
    new_P1_ADD_515_U133, new_P1_ADD_515_U132, new_P1_ADD_515_U131,
    new_P1_ADD_515_U130, new_P1_ADD_515_U129, new_P1_ADD_515_U128,
    new_P1_ADD_515_U127, new_P1_ADD_515_U126, new_P1_ADD_515_U125,
    new_P1_ADD_515_U124, new_P1_ADD_515_U123, new_P1_ADD_515_U122,
    new_P1_ADD_515_U121, new_P1_ADD_515_U120, new_P1_ADD_515_U119,
    new_P1_ADD_515_U118, new_P1_ADD_515_U117, new_P1_ADD_515_U116,
    new_P1_ADD_515_U115, new_P1_ADD_515_U114, new_P1_ADD_515_U113,
    new_P1_ADD_515_U112, new_P1_ADD_515_U111, new_P1_ADD_515_U110,
    new_P1_ADD_515_U109, new_P1_ADD_515_U108, new_P1_ADD_515_U107,
    new_P1_ADD_515_U106, new_P1_ADD_515_U105, new_P1_ADD_515_U104,
    new_P1_ADD_515_U103, new_P1_ADD_515_U102, new_P1_ADD_515_U101,
    new_P1_ADD_515_U100, new_P1_ADD_515_U99, new_P1_ADD_515_U98,
    new_P1_ADD_515_U97, new_P1_ADD_515_U96, new_P1_ADD_515_U95,
    new_P1_ADD_515_U94, new_P1_ADD_515_U93, new_P1_ADD_515_U92,
    new_P1_ADD_515_U91, new_P1_ADD_515_U90, new_P1_ADD_515_U89,
    new_P1_ADD_515_U88, new_P1_ADD_515_U87, new_P1_ADD_515_U86,
    new_P1_ADD_515_U85, new_P1_ADD_515_U84, new_P1_ADD_515_U83,
    new_P1_ADD_515_U82, new_P1_ADD_515_U81, new_P1_ADD_515_U80,
    new_P1_ADD_515_U79, new_P1_ADD_515_U78, new_P1_ADD_515_U77,
    new_P1_ADD_515_U76, new_P1_ADD_515_U75, new_P1_ADD_515_U74,
    new_P1_ADD_515_U73, new_P1_ADD_515_U72, new_P1_ADD_515_U71,
    new_P1_ADD_515_U70, new_P1_ADD_515_U69, new_P1_ADD_515_U68,
    new_P1_ADD_515_U67, new_P1_ADD_515_U66, new_P1_ADD_515_U65,
    new_P1_ADD_515_U64, new_P1_ADD_515_U63, new_P1_ADD_515_U62,
    new_P1_ADD_515_U61, new_P1_ADD_515_U60, new_P1_ADD_515_U59,
    new_P1_ADD_515_U58, new_P1_ADD_515_U57, new_P1_ADD_515_U56,
    new_P1_ADD_515_U55, new_P1_ADD_515_U54, new_P1_ADD_515_U53,
    new_P1_ADD_515_U52, new_P1_ADD_515_U51, new_P1_ADD_515_U50,
    new_P1_ADD_515_U49, new_P1_ADD_515_U48, new_P1_ADD_515_U47,
    new_P1_ADD_515_U46, new_P1_ADD_515_U45, new_P1_ADD_515_U44,
    new_P1_ADD_515_U43, new_P1_ADD_515_U42, new_P1_ADD_515_U41,
    new_P1_ADD_515_U40, new_P1_ADD_515_U39, new_P1_ADD_515_U38,
    new_P1_ADD_515_U37, new_P1_ADD_515_U36, new_P1_ADD_515_U35,
    new_P1_ADD_515_U34, new_P1_ADD_515_U33, new_P1_ADD_515_U32,
    new_P1_ADD_515_U31, new_P1_ADD_515_U30, new_P1_ADD_515_U29,
    new_P1_ADD_515_U28, new_P1_ADD_515_U27, new_P1_ADD_515_U26,
    new_P1_ADD_515_U25, new_P1_ADD_515_U24, new_P1_ADD_515_U23,
    new_P1_ADD_515_U22, new_P1_ADD_515_U21, new_P1_ADD_515_U20,
    new_P1_ADD_515_U19, new_P1_ADD_515_U18, new_P1_ADD_515_U17,
    new_P1_ADD_515_U16, new_P1_ADD_515_U15, new_P1_ADD_515_U14,
    new_P1_ADD_515_U13, new_P1_ADD_515_U12, new_P1_ADD_515_U11,
    new_P1_ADD_515_U10, new_P1_ADD_515_U9, new_P1_ADD_515_U8,
    new_P1_ADD_515_U7, new_P1_ADD_515_U6, new_P1_ADD_515_U5,
    new_P1_ADD_515_U4, new_P1_GTE_485_U7, new_P1_GTE_485_U6,
    new_P1_ADD_405_U186, new_P1_ADD_405_U185, new_P1_ADD_405_U184,
    new_P1_ADD_405_U183, new_P1_ADD_405_U182, new_P1_ADD_405_U181,
    new_P1_ADD_405_U180, new_P1_ADD_405_U179, new_P1_ADD_405_U178,
    new_P1_ADD_405_U177, new_P1_ADD_405_U176, new_P1_ADD_405_U175,
    new_P1_ADD_405_U174, new_P1_ADD_405_U173, new_P2_U2352, new_P2_U2353,
    new_P2_U2354, new_P2_U2355, new_P2_U2356, new_P2_U2357, new_P2_U2358,
    new_P2_U2359, new_P2_U2360, new_P2_U2361, new_P2_U2362, new_P2_U2363,
    new_P2_U2364, new_P2_U2365, new_P2_U2366, new_P2_U2367, new_P2_U2368,
    new_P2_U2369, new_P2_U2370, new_P2_U2371, new_P2_U2372, new_P2_U2373,
    new_P2_U2374, new_P2_U2375, new_P2_U2376, new_P2_U2377, new_P2_U2378,
    new_P2_U2379, new_P2_U2380, new_P2_U2381, new_P2_U2382, new_P2_U2383,
    new_P2_U2384, new_P2_U2385, new_P2_U2386, new_P2_U2387, new_P2_U2388,
    new_P2_U2389, new_P2_U2390, new_P2_U2391, new_P2_U2392, new_P2_U2393,
    new_P2_U2394, new_P2_U2395, new_P2_U2396, new_P2_U2397, new_P2_U2398,
    new_P2_U2399, new_P2_U2400, new_P2_U2401, new_P2_U2402, new_P2_U2403,
    new_P2_U2404, new_P2_U2405, new_P2_U2406, new_P2_U2407, new_P2_U2408,
    new_P2_U2409, new_P2_U2410, new_P2_U2411, new_P2_U2412, new_P2_U2413,
    new_P2_U2414, new_P2_U2415, new_P2_U2416, new_P2_U2417, new_P2_U2418,
    new_P2_U2419, new_P2_U2420, new_P2_U2421, new_P2_U2422, new_P2_U2423,
    new_P2_U2424, new_P2_U2425, new_P2_U2426, new_P2_U2427, new_P2_U2428,
    new_P2_U2429, new_P2_U2430, new_P2_U2431, new_P2_U2432, new_P2_U2433,
    new_P2_U2434, new_P2_U2435, new_P2_U2436, new_P2_U2437, new_P2_U2438,
    new_P2_U2439, new_P2_U2440, new_P2_U2441, new_P2_U2442, new_P2_U2443,
    new_P2_U2444, new_P2_U2445, new_P2_U2446, new_P2_U2447, new_P2_U2448,
    new_P2_U2449, new_P2_U2450, new_P2_U2451, new_P2_U2452, new_P2_U2453,
    new_P2_U2454, new_P2_U2455, new_P2_U2456, new_P2_U2457, new_P2_U2458,
    new_P2_U2459, new_P2_U2460, new_P2_U2461, new_P2_U2462, new_P2_U2463,
    new_P2_U2464, new_P2_U2465, new_P2_U2466, new_P2_U2467, new_P2_U2468,
    new_P2_U2469, new_P2_U2470, new_P2_U2471, new_P2_U2472, new_P2_U2473,
    new_P2_U2474, new_P2_U2475, new_P2_U2476, new_P2_U2477, new_P2_U2478,
    new_P2_U2479, new_P2_U2480, new_P2_U2481, new_P2_U2482, new_P2_U2483,
    new_P2_U2484, new_P2_U2485, new_P2_U2486, new_P2_U2487, new_P2_U2488,
    new_P2_U2489, new_P2_U2490, new_P2_U2491, new_P2_U2492, new_P2_U2493,
    new_P2_U2494, new_P2_U2495, new_P2_U2496, new_P2_U2497, new_P2_U2498,
    new_P2_U2499, new_P2_U2500, new_P2_U2501, new_P2_U2502, new_P2_U2503,
    new_P2_U2504, new_P2_U2505, new_P2_U2506, new_P2_U2507, new_P2_U2508,
    new_P2_U2509, new_P2_U2510, new_P2_U2511, new_P2_U2512, new_P2_U2513,
    new_P2_U2514, new_P2_U2515, new_P2_U2516, new_P2_U2517, new_P2_U2518,
    new_P2_U2519, new_P2_U2520, new_P2_U2521, new_P2_U2522, new_P2_U2523,
    new_P2_U2524, new_P2_U2525, new_P2_U2526, new_P2_U2527, new_P2_U2528,
    new_P2_U2529, new_P2_U2530, new_P2_U2531, new_P2_U2532, new_P2_U2533,
    new_P2_U2534, new_P2_U2535, new_P2_U2536, new_P2_U2537, new_P2_U2538,
    new_P2_U2539, new_P2_U2540, new_P2_U2541, new_P2_U2542, new_P2_U2543,
    new_P2_U2544, new_P2_U2545, new_P2_U2546, new_P2_U2547, new_P2_U2548,
    new_P2_U2549, new_P2_U2550, new_P2_U2551, new_P2_U2552, new_P2_U2553,
    new_P2_U2554, new_P2_U2555, new_P2_U2556, new_P2_U2557, new_P2_U2558,
    new_P2_U2559, new_P2_U2560, new_P2_U2561, new_P2_U2562, new_P2_U2563,
    new_P2_U2564, new_P2_U2565, new_P2_U2566, new_P2_U2567, new_P2_U2568,
    new_P2_U2569, new_P2_U2570, new_P2_U2571, new_P2_U2572, new_P2_U2573,
    new_P2_U2574, new_P2_U2575, new_P2_U2576, new_P2_U2577, new_P2_U2578,
    new_P2_U2579, new_P2_U2580, new_P2_U2581, new_P2_U2582, new_P2_U2583,
    new_P2_U2584, new_P2_U2585, new_P2_U2586, new_P2_U2587, new_P2_U2588,
    new_P2_U2589, new_P2_U2590, new_P2_U2591, new_P2_U2592, new_P2_U2593,
    new_P2_U2594, new_P2_U2595, new_P2_U2596, new_P2_U2597, new_P2_U2598,
    new_P2_U2599, new_P2_U2600, new_P2_U2601, new_P2_U2602, new_P2_U2603,
    new_P2_U2604, new_P2_U2605, new_P2_U2606, new_P2_U2607, new_P2_U2608,
    new_P2_U2609, new_P2_U2610, new_P2_U2611, new_P2_U2612, new_P2_U2613,
    new_P2_U2614, new_P2_U2615, new_P2_U2616, new_P2_U2617, new_P2_U2618,
    new_P2_U2619, new_P2_U2620, new_P2_U2621, new_P2_U2622, new_P2_U2623,
    new_P2_U2624, new_P2_U2625, new_P2_U2626, new_P2_U2627, new_P2_U2628,
    new_P2_U2629, new_P2_U2630, new_P2_U2631, new_P2_U2632, new_P2_U2633,
    new_P2_U2634, new_P2_U2635, new_P2_U2636, new_P2_U2637, new_P2_U2638,
    new_P2_U2639, new_P2_U2640, new_P2_U2641, new_P2_U2642, new_P2_U2643,
    new_P2_U2644, new_P2_U2645, new_P2_U2646, new_P2_U2647, new_P2_U2648,
    new_P2_U2649, new_P2_U2650, new_P2_U2651, new_P2_U2652, new_P2_U2653,
    new_P2_U2654, new_P2_U2655, new_P2_U2656, new_P2_U2657, new_P2_U2658,
    new_P2_U2659, new_P2_U2660, new_P2_U2661, new_P2_U2662, new_P2_U2663,
    new_P2_U2664, new_P2_U2665, new_P2_U2666, new_P2_U2667, new_P2_U2668,
    new_P2_U2669, new_P2_U2670, new_P2_U2671, new_P2_U2672, new_P2_U2673,
    new_P2_U2674, new_P2_U2675, new_P2_U2676, new_P2_U2677, new_P2_U2678,
    new_P2_U2679, new_P2_U2680, new_P2_U2681, new_P2_U2682, new_P2_U2683,
    new_P2_U2684, new_P2_U2685, new_P2_U2686, new_P2_U2687, new_P2_U2688,
    new_P2_U2689, new_P2_U2690, new_P2_U2691, new_P2_U2692, new_P2_U2693,
    new_P2_U2694, new_P2_U2695, new_P2_U2696, new_P1_ADD_405_U172,
    new_P2_U2698, new_P2_U2699, new_P2_U2700, new_P2_U2701, new_P2_U2702,
    new_P2_U2703, new_P2_U2704, new_P2_U2705, new_P2_U2706, new_P2_U2707,
    new_P2_U2708, new_P2_U2709, new_P2_U2710, new_P2_U2711, new_P2_U2712,
    new_P2_U2713, new_P2_U2714, new_P2_U2715, new_P2_U2716, new_P2_U2717,
    new_P2_U2718, new_P2_U2719, new_P2_U2720, new_P2_U2721, new_P2_U2722,
    new_P2_U2723, new_P2_U2724, new_P2_U2725, new_P2_U2726, new_P2_U2727,
    new_P2_U2728, new_P2_U2729, new_P2_U2730, new_P2_U2731, new_P2_U2732,
    new_P2_U2733, new_P2_U2734, new_P2_U2735, new_P2_U2736, new_P2_U2737,
    new_P2_U2738, new_P2_U2739, new_P2_U2740, new_P2_U2741, new_P2_U2742,
    new_P2_U2743, new_P2_U2744, new_P2_U2745, new_P2_U2746, new_P2_U2747,
    new_P2_U2748, new_P2_U2749, new_P2_U2750, new_P2_U2751, new_P2_U2752,
    new_P2_U2753, new_P2_U2754, new_P2_U2755, new_P2_U2756, new_P2_U2757,
    new_P2_U2758, new_P2_U2759, new_P2_U2760, new_P2_U2761, new_P2_U2762,
    new_P2_U2763, new_P2_U2764, new_P2_U2765, new_P2_U2766, new_P2_U2767,
    new_P2_U2768, new_P2_U2769, new_P2_U2770, new_P2_U2771, new_P2_U2772,
    new_P2_U2773, new_P2_U2774, new_P2_U2775, new_P2_U2776, new_P2_U2777,
    new_P2_U2778, new_P2_U2779, new_P2_U2780, new_P2_U2781, new_P2_U2782,
    new_P2_U2783, new_P2_U2784, new_P2_U2785, new_P2_U2786, new_P2_U2787,
    new_P2_U2788, new_P2_U2789, new_P2_U2790, new_P2_U2791, new_P2_U2792,
    new_P2_U2793, new_P2_U2794, new_P2_U2795, new_P2_U2796, new_P2_U2797,
    new_P2_U2798, new_P2_U2799, new_P2_U2800, new_P2_U2801, new_P2_U2802,
    new_P2_U2803, new_P2_U2804, new_P2_U2805, new_P2_U2806, new_P2_U2807,
    new_P2_U2808, new_P2_U2809, new_P2_U2810, new_P2_U2811, new_P2_U2812,
    new_P2_U2813, new_P2_U3242, new_P2_U3243, new_P2_U3244, new_P2_U3245,
    new_P2_U3246, new_P2_U3247, new_P2_U3248, new_P2_U3249, new_P2_U3250,
    new_P2_U3251, new_P2_U3252, new_P2_U3253, new_P2_U3254, new_P2_U3255,
    new_P2_U3256, new_P2_U3257, new_P2_U3258, new_P2_U3259, new_P2_U3260,
    new_P2_U3261, new_P2_U3262, new_P2_U3263, new_P2_U3264, new_P2_U3265,
    new_P2_U3266, new_P2_U3267, new_P2_U3268, new_P2_U3269, new_P2_U3270,
    new_P2_U3271, new_P2_U3272, new_P2_U3273, new_P2_U3274, new_P2_U3275,
    new_P2_U3276, new_P2_U3277, new_P2_U3278, new_P2_U3279, new_P2_U3280,
    new_P2_U3281, new_P2_U3282, new_P2_U3283, new_P2_U3284, new_P2_U3285,
    new_P2_U3286, new_P2_U3287, new_P2_U3288, new_P2_U3289, new_P2_U3290,
    new_P2_U3291, new_P2_U3292, new_P2_U3293, new_P2_U3294, new_P2_U3295,
    new_P2_U3296, new_P2_U3297, new_P2_U3298, new_P2_U3299, new_P2_U3300,
    new_P2_U3301, new_P2_U3302, new_P2_U3303, new_P2_U3304, new_P2_U3305,
    new_P2_U3306, new_P2_U3307, new_P2_U3308, new_P2_U3309, new_P2_U3310,
    new_P2_U3311, new_P2_U3312, new_P2_U3313, new_P2_U3314, new_P2_U3315,
    new_P2_U3316, new_P2_U3317, new_P2_U3318, new_P2_U3319, new_P2_U3320,
    new_P2_U3321, new_P2_U3322, new_P2_U3323, new_P2_U3324, new_P2_U3325,
    new_P2_U3326, new_P2_U3327, new_P2_U3328, new_P2_U3329, new_P2_U3330,
    new_P2_U3331, new_P2_U3332, new_P2_U3333, new_P2_U3334, new_P2_U3335,
    new_P2_U3336, new_P2_U3337, new_P2_U3338, new_P2_U3339, new_P2_U3340,
    new_P2_U3341, new_P2_U3342, new_P2_U3343, new_P2_U3344, new_P2_U3345,
    new_P2_U3346, new_P2_U3347, new_P2_U3348, new_P2_U3349, new_P2_U3350,
    new_P2_U3351, new_P2_U3352, new_P2_U3353, new_P2_U3354, new_P2_U3355,
    new_P2_U3356, new_P2_U3357, new_P2_U3358, new_P2_U3359, new_P2_U3360,
    new_P2_U3361, new_P2_U3362, new_P2_U3363, new_P2_U3364, new_P2_U3365,
    new_P2_U3366, new_P2_U3367, new_P2_U3368, new_P2_U3369, new_P2_U3370,
    new_P2_U3371, new_P2_U3372, new_P2_U3373, new_P2_U3374, new_P2_U3375,
    new_P2_U3376, new_P2_U3377, new_P2_U3378, new_P2_U3379, new_P2_U3380,
    new_P2_U3381, new_P2_U3382, new_P2_U3383, new_P2_U3384, new_P2_U3385,
    new_P2_U3386, new_P2_U3387, new_P2_U3388, new_P2_U3389, new_P2_U3390,
    new_P2_U3391, new_P2_U3392, new_P2_U3393, new_P2_U3394, new_P2_U3395,
    new_P2_U3396, new_P2_U3397, new_P2_U3398, new_P2_U3399, new_P2_U3400,
    new_P2_U3401, new_P2_U3402, new_P2_U3403, new_P2_U3404, new_P2_U3405,
    new_P2_U3406, new_P2_U3407, new_P2_U3408, new_P2_U3409, new_P2_U3410,
    new_P2_U3411, new_P2_U3412, new_P2_U3413, new_P2_U3414, new_P2_U3415,
    new_P2_U3416, new_P2_U3417, new_P2_U3418, new_P2_U3419, new_P2_U3420,
    new_P2_U3421, new_P2_U3422, new_P2_U3423, new_P2_U3424, new_P2_U3425,
    new_P2_U3426, new_P2_U3427, new_P2_U3428, new_P2_U3429, new_P2_U3430,
    new_P2_U3431, new_P2_U3432, new_P2_U3433, new_P2_U3434, new_P2_U3435,
    new_P2_U3436, new_P2_U3437, new_P2_U3438, new_P2_U3439, new_P2_U3440,
    new_P2_U3441, new_P2_U3442, new_P2_U3443, new_P2_U3444, new_P2_U3445,
    new_P2_U3446, new_P2_U3447, new_P2_U3448, new_P2_U3449, new_P2_U3450,
    new_P2_U3451, new_P2_U3452, new_P2_U3453, new_P2_U3454, new_P2_U3455,
    new_P2_U3456, new_P2_U3457, new_P2_U3458, new_P2_U3459, new_P2_U3460,
    new_P2_U3461, new_P2_U3462, new_P2_U3463, new_P2_U3464, new_P2_U3465,
    new_P2_U3466, new_P2_U3467, new_P2_U3468, new_P2_U3469, new_P2_U3470,
    new_P2_U3471, new_P2_U3472, new_P2_U3473, new_P2_U3474, new_P2_U3475,
    new_P2_U3476, new_P2_U3477, new_P2_U3478, new_P2_U3479, new_P2_U3480,
    new_P2_U3481, new_P2_U3482, new_P2_U3483, new_P2_U3484, new_P2_U3485,
    new_P2_U3486, new_P2_U3487, new_P2_U3488, new_P2_U3489, new_P2_U3490,
    new_P2_U3491, new_P2_U3492, new_P2_U3493, new_P2_U3494, new_P2_U3495,
    new_P2_U3496, new_P2_U3497, new_P2_U3498, new_P2_U3499, new_P2_U3500,
    new_P2_U3501, new_P2_U3502, new_P2_U3503, new_P2_U3504, new_P2_U3505,
    new_P2_U3506, new_P2_U3507, new_P2_U3508, new_P2_U3509, new_P2_U3510,
    new_P2_U3511, new_P2_U3512, new_P2_U3513, new_P2_U3514, new_P2_U3515,
    new_P2_U3516, new_P2_U3517, new_P2_U3518, new_P2_U3519, new_P2_U3520,
    new_P2_U3521, new_P2_U3522, new_P2_U3523, new_P2_U3524, new_P2_U3525,
    new_P2_U3526, new_P2_U3527, new_P2_U3528, new_P2_U3529, new_P2_U3530,
    new_P2_U3531, new_P2_U3532, new_P2_U3533, new_P2_U3534, new_P2_U3535,
    new_P2_U3536, new_P2_U3537, new_P2_U3538, new_P2_U3539, new_P2_U3540,
    new_P2_U3541, new_P2_U3542, new_P2_U3543, new_P2_U3544, new_P2_U3545,
    new_P2_U3546, new_P2_U3547, new_P2_U3548, new_P2_U3549, new_P2_U3550,
    new_P2_U3551, new_P2_U3552, new_P2_U3553, new_P2_U3554, new_P2_U3555,
    new_P2_U3556, new_P2_U3557, new_P2_U3558, new_P2_U3559, new_P2_U3560,
    new_P2_U3561, new_P2_U3562, new_P2_U3563, new_P2_U3564, new_P2_U3565,
    new_P2_U3566, new_P2_U3567, new_P2_U3568, new_P2_U3569, new_P2_U3570,
    new_P2_U3571, new_P2_U3572, new_P2_U3573, new_P2_U3574, new_P2_U3575,
    new_P2_U3576, new_P2_U3577, new_P2_U3578, new_P2_U3579, new_P2_U3580,
    new_P2_U3581, new_P2_U3582, new_P2_U3583, new_P2_U3584, new_P2_U3589,
    new_P2_U3590, new_P2_U3594, new_P2_U3597, new_P2_U3598, new_P2_U3606,
    new_P2_U3607, new_P2_U3613, new_P2_U3614, new_P2_U3615, new_P2_U3616,
    new_P2_U3617, new_P2_U3618, new_P2_U3619, new_P2_U3620, new_P2_U3621,
    new_P2_U3622, new_P2_U3623, new_P2_U3624, new_P2_U3625, new_P2_U3626,
    new_P2_U3627, new_P2_U3628, new_P2_U3629, new_P2_U3630, new_P2_U3631,
    new_P2_U3632, new_P2_U3633, new_P2_U3634, new_P2_U3635, new_P2_U3636,
    new_P2_U3637, new_P2_U3638, new_P2_U3639, new_P2_U3640, new_P2_U3641,
    new_P2_U3642, new_P2_U3643, new_P2_U3644, new_P2_U3645, new_P2_U3646,
    new_P2_U3647, new_P2_U3648, new_P2_U3649, new_P2_U3650, new_P2_U3651,
    new_P2_U3652, new_P2_U3653, new_P2_U3654, new_P2_U3655, new_P2_U3656,
    new_P2_U3657, new_P2_U3658, new_P2_U3659, new_P2_U3660, new_P2_U3661,
    new_P2_U3662, new_P2_U3663, new_P2_U3664, new_P2_U3665, new_P2_U3666,
    new_P2_U3667, new_P2_U3668, new_P2_U3669, new_P2_U3670, new_P2_U3671,
    new_P2_U3672, new_P2_U3673, new_P2_U3674, new_P2_U3675, new_P2_U3676,
    new_P2_U3677, new_P2_U3678, new_P2_U3679, new_P2_U3680, new_P2_U3681,
    new_P2_U3682, new_P2_U3683, new_P2_U3684, new_P2_U3685, new_P2_U3686,
    new_P2_U3687, new_P2_U3688, new_P2_U3689, new_P2_U3690, new_P2_U3691,
    new_P2_U3692, new_P2_U3693, new_P2_U3694, new_P2_U3695, new_P2_U3696,
    new_P2_U3697, new_P2_U3698, new_P2_U3699, new_P2_U3700, new_P2_U3701,
    new_P2_U3702, new_P2_U3703, new_P2_U3704, new_P2_U3705, new_P2_U3706,
    new_P2_U3707, new_P2_U3708, new_P2_U3709, new_P2_U3710, new_P2_U3711,
    new_P2_U3712, new_P2_U3713, new_P2_U3714, new_P2_U3715, new_P2_U3716,
    new_P2_U3717, new_P2_U3718, new_P2_U3719, new_P2_U3720, new_P2_U3721,
    new_P2_U3722, new_P2_U3723, new_P2_U3724, new_P2_U3725, new_P2_U3726,
    new_P2_U3727, new_P2_U3728, new_P2_U3729, new_P2_U3730, new_P2_U3731,
    new_P2_U3732, new_P2_U3733, new_P2_U3734, new_P2_U3735, new_P2_U3736,
    new_P2_U3737, new_P2_U3738, new_P2_U3739, new_P2_U3740, new_P2_U3741,
    new_P2_U3742, new_P2_U3743, new_P2_U3744, new_P2_U3745, new_P2_U3746,
    new_P2_U3747, new_P2_U3748, new_P2_U3749, new_P2_U3750, new_P2_U3751,
    new_P2_U3752, new_P2_U3753, new_P2_U3754, new_P2_U3755, new_P2_U3756,
    new_P2_U3757, new_P2_U3758, new_P2_U3759, new_P2_U3760, new_P2_U3761,
    new_P2_U3762, new_P2_U3763, new_P2_U3764, new_P2_U3765, new_P2_U3766,
    new_P2_U3767, new_P2_U3768, new_P2_U3769, new_P2_U3770, new_P2_U3771,
    new_P2_U3772, new_P2_U3773, new_P2_U3774, new_P2_U3775, new_P2_U3776,
    new_P2_U3777, new_P2_U3778, new_P2_U3779, new_P2_U3780, new_P2_U3781,
    new_P2_U3782, new_P2_U3783, new_P2_U3784, new_P2_U3785, new_P2_U3786,
    new_P2_U3787, new_P2_U3788, new_P2_U3789, new_P2_U3790, new_P2_U3791,
    new_P2_U3792, new_P2_U3793, new_P2_U3794, new_P2_U3795, new_P2_U3796,
    new_P2_U3797, new_P2_U3798, new_P2_U3799, new_P2_U3800, new_P2_U3801,
    new_P2_U3802, new_P2_U3803, new_P2_U3804, new_P2_U3805, new_P2_U3806,
    new_P2_U3807, new_P2_U3808, new_P2_U3809, new_P2_U3810, new_P2_U3811,
    new_P2_U3812, new_P2_U3813, new_P2_U3814, new_P2_U3815, new_P2_U3816,
    new_P2_U3817, new_P2_U3818, new_P2_U3819, new_P2_U3820, new_P2_U3821,
    new_P2_U3822, new_P2_U3823, new_P2_U3824, new_P2_U3825, new_P2_U3826,
    new_P2_U3827, new_P2_U3828, new_P2_U3829, new_P2_U3830, new_P2_U3831,
    new_P2_U3832, new_P2_U3833, new_P2_U3834, new_P2_U3835, new_P2_U3836,
    new_P2_U3837, new_P2_U3838, new_P2_U3839, new_P2_U3840, new_P2_U3841,
    new_P2_U3842, new_P2_U3843, new_P2_U3844, new_P2_U3845, new_P2_U3846,
    new_P2_U3847, new_P2_U3848, new_P2_U3849, new_P2_U3850, new_P2_U3851,
    new_P2_U3852, new_P2_U3853, new_P2_U3854, new_P2_U3855, new_P2_U3856,
    new_P2_U3857, new_P2_U3858, new_P2_U3859, new_P2_U3860, new_P2_U3861,
    new_P2_U3862, new_P2_U3863, new_P2_U3864, new_P2_U3865, new_P2_U3866,
    new_P2_U3867, new_P2_U3868, new_P2_U3869, new_P2_U3870, new_P2_U3871,
    new_P2_U3872, new_P2_U3873, new_P2_U3874, new_P2_U3875, new_P2_U3876,
    new_P2_U3877, new_P2_U3878, new_P2_U3879, new_P2_U3880, new_P2_U3881,
    new_P2_U3882, new_P2_U3883, new_P2_U3884, new_P2_U3885, new_P2_U3886,
    new_P2_U3887, new_P2_U3888, new_P2_U3889, new_P2_U3890, new_P2_U3891,
    new_P2_U3892, new_P2_U3893, new_P2_U3894, new_P2_U3895, new_P2_U3896,
    new_P2_U3897, new_P2_U3898, new_P2_U3899, new_P2_U3900, new_P2_U3901,
    new_P2_U3902, new_P2_U3903, new_P2_U3904, new_P2_U3905, new_P2_U3906,
    new_P2_U3907, new_P2_U3908, new_P2_U3909, new_P2_U3910, new_P2_U3911,
    new_P2_U3912, new_P2_U3913, new_P2_U3914, new_P2_U3915, new_P2_U3916,
    new_P2_U3917, new_P2_U3918, new_P2_U3919, new_P2_U3920, new_P2_U3921,
    new_P2_U3922, new_P2_U3923, new_P2_U3924, new_P2_U3925, new_P2_U3926,
    new_P2_U3927, new_P2_U3928, new_P2_U3929, new_P2_U3930, new_P2_U3931,
    new_P2_U3932, new_P2_U3933, new_P2_U3934, new_P2_U3935, new_P2_U3936,
    new_P2_U3937, new_P2_U3938, new_P2_U3939, new_P2_U3940, new_P2_U3941,
    new_P2_U3942, new_P2_U3943, new_P2_U3944, new_P2_U3945, new_P2_U3946,
    new_P2_U3947, new_P2_U3948, new_P2_U3949, new_P2_U3950, new_P2_U3951,
    new_P2_U3952, new_P2_U3953, new_P2_U3954, new_P2_U3955, new_P2_U3956,
    new_P2_U3957, new_P2_U3958, new_P2_U3959, new_P2_U3960, new_P2_U3961,
    new_P2_U3962, new_P2_U3963, new_P2_U3964, new_P2_U3965, new_P2_U3966,
    new_P2_U3967, new_P2_U3968, new_P2_U3969, new_P2_U3970, new_P2_U3971,
    new_P2_U3972, new_P2_U3973, new_P2_U3974, new_P2_U3975, new_P2_U3976,
    new_P2_U3977, new_P2_U3978, new_P2_U3979, new_P2_U3980, new_P2_U3981,
    new_P2_U3982, new_P2_U3983, new_P2_U3984, new_P2_U3985, new_P2_U3986,
    new_P2_U3987, new_P2_U3988, new_P2_U3989, new_P2_U3990, new_P2_U3991,
    new_P2_U3992, new_P2_U3993, new_P2_U3994, new_P2_U3995, new_P2_U3996,
    new_P2_U3997, new_P2_U3998, new_P2_U3999, new_P2_U4000, new_P2_U4001,
    new_P2_U4002, new_P2_U4003, new_P2_U4004, new_P2_U4005, new_P2_U4006,
    new_P2_U4007, new_P2_U4008, new_P2_U4009, new_P2_U4010, new_P2_U4011,
    new_P2_U4012, new_P2_U4013, new_P2_U4014, new_P2_U4015, new_P2_U4016,
    new_P2_U4017, new_P2_U4018, new_P2_U4019, new_P2_U4020, new_P2_U4021,
    new_P2_U4022, new_P2_U4023, new_P2_U4024, new_P2_U4025, new_P2_U4026,
    new_P2_U4027, new_P2_U4028, new_P2_U4029, new_P2_U4030, new_P2_U4031,
    new_P2_U4032, new_P2_U4033, new_P2_U4034, new_P2_U4035, new_P2_U4036,
    new_P2_U4037, new_P2_U4038, new_P2_U4039, new_P2_U4040, new_P2_U4041,
    new_P2_U4042, new_P2_U4043, new_P2_U4044, new_P2_U4045, new_P2_U4046,
    new_P2_U4047, new_P2_U4048, new_P2_U4049, new_P2_U4050, new_P2_U4051,
    new_P2_U4052, new_P2_U4053, new_P2_U4054, new_P2_U4055, new_P2_U4056,
    new_P2_U4057, new_P2_U4058, new_P2_U4059, new_P2_U4060, new_P2_U4061,
    new_P2_U4062, new_P2_U4063, new_P2_U4064, new_P2_U4065, new_P2_U4066,
    new_P2_U4067, new_P2_U4068, new_P2_U4069, new_P2_U4070, new_P2_U4071,
    new_P2_U4072, new_P2_U4073, new_P2_U4074, new_P2_U4075, new_P2_U4076,
    new_P2_U4077, new_P2_U4078, new_P2_U4079, new_P2_U4080, new_P2_U4081,
    new_P2_U4082, new_P2_U4083, new_P2_U4084, new_P2_U4085, new_P2_U4086,
    new_P2_U4087, new_P2_U4088, new_P2_U4089, new_P2_U4090, new_P2_U4091,
    new_P2_U4092, new_P2_U4093, new_P2_U4094, new_P2_U4095, new_P2_U4096,
    new_P2_U4097, new_P2_U4098, new_P2_U4099, new_P2_U4100, new_P2_U4101,
    new_P2_U4102, new_P2_U4103, new_P2_U4104, new_P2_U4105, new_P2_U4106,
    new_P2_U4107, new_P2_U4108, new_P2_U4109, new_P2_U4110, new_P2_U4111,
    new_P2_U4112, new_P2_U4113, new_P2_U4114, new_P2_U4115, new_P2_U4116,
    new_P2_U4117, new_P2_U4118, new_P2_U4119, new_P2_U4120, new_P2_U4121,
    new_P2_U4122, new_P2_U4123, new_P2_U4124, new_P2_U4125, new_P2_U4126,
    new_P2_U4127, new_P2_U4128, new_P2_U4129, new_P2_U4130, new_P2_U4131,
    new_P2_U4132, new_P2_U4133, new_P2_U4134, new_P2_U4135, new_P2_U4136,
    new_P2_U4137, new_P2_U4138, new_P2_U4139, new_P2_U4140, new_P2_U4141,
    new_P2_U4142, new_P2_U4143, new_P2_U4144, new_P2_U4145, new_P2_U4146,
    new_P2_U4147, new_P2_U4148, new_P2_U4149, new_P2_U4150, new_P2_U4151,
    new_P2_U4152, new_P2_U4153, new_P2_U4154, new_P2_U4155, new_P2_U4156,
    new_P2_U4157, new_P2_U4158, new_P2_U4159, new_P2_U4160, new_P2_U4161,
    new_P2_U4162, new_P2_U4163, new_P2_U4164, new_P2_U4165, new_P2_U4166,
    new_P2_U4167, new_P2_U4168, new_P2_U4169, new_P2_U4170, new_P2_U4171,
    new_P2_U4172, new_P2_U4173, new_P2_U4174, new_P2_U4175, new_P2_U4176,
    new_P2_U4177, new_P2_U4178, new_P2_U4179, new_P2_U4180, new_P2_U4181,
    new_P2_U4182, new_P2_U4183, new_P2_U4184, new_P2_U4185, new_P2_U4186,
    new_P2_U4187, new_P2_U4188, new_P2_U4189, new_P2_U4190, new_P2_U4191,
    new_P2_U4192, new_P2_U4193, new_P2_U4194, new_P2_U4195, new_P2_U4196,
    new_P2_U4197, new_P2_U4198, new_P2_U4199, new_P2_U4200, new_P2_U4201,
    new_P2_U4202, new_P2_U4203, new_P2_U4204, new_P2_U4205, new_P2_U4206,
    new_P2_U4207, new_P2_U4208, new_P2_U4209, new_P2_U4210, new_P2_U4211,
    new_P2_U4212, new_P2_U4213, new_P2_U4214, new_P2_U4215, new_P2_U4216,
    new_P2_U4217, new_P2_U4218, new_P2_U4219, new_P2_U4220, new_P2_U4221,
    new_P2_U4222, new_P2_U4223, new_P2_U4224, new_P2_U4225, new_P2_U4226,
    new_P2_U4227, new_P2_U4228, new_P2_U4229, new_P2_U4230, new_P2_U4231,
    new_P2_U4232, new_P2_U4233, new_P2_U4234, new_P2_U4235, new_P2_U4236,
    new_P2_U4237, new_P2_U4238, new_P2_U4239, new_P2_U4240, new_P2_U4241,
    new_P2_U4242, new_P2_U4243, new_P2_U4244, new_P2_U4245, new_P2_U4246,
    new_P2_U4247, new_P2_U4248, new_P2_U4249, new_P2_U4250, new_P2_U4251,
    new_P2_U4252, new_P2_U4253, new_P2_U4254, new_P2_U4255, new_P2_U4256,
    new_P2_U4257, new_P2_U4258, new_P2_U4259, new_P2_U4260, new_P2_U4261,
    new_P2_U4262, new_P2_U4263, new_P2_U4264, new_P2_U4265, new_P2_U4266,
    new_P2_U4267, new_P2_U4268, new_P2_U4269, new_P2_U4270, new_P2_U4271,
    new_P2_U4272, new_P2_U4273, new_P2_U4274, new_P2_U4275, new_P2_U4276,
    new_P2_U4277, new_P2_U4278, new_P2_U4279, new_P2_U4280, new_P2_U4281,
    new_P2_U4282, new_P2_U4283, new_P2_U4284, new_P2_U4285, new_P2_U4286,
    new_P2_U4287, new_P2_U4288, new_P2_U4289, new_P2_U4290, new_P2_U4291,
    new_P2_U4292, new_P2_U4293, new_P2_U4294, new_P2_U4295, new_P2_U4296,
    new_P2_U4297, new_P2_U4298, new_P2_U4299, new_P2_U4300, new_P2_U4301,
    new_P2_U4302, new_P2_U4303, new_P2_U4304, new_P2_U4305, new_P2_U4306,
    new_P2_U4307, new_P2_U4308, new_P2_U4309, new_P2_U4310, new_P2_U4311,
    new_P2_U4312, new_P2_U4313, new_P2_U4314, new_P2_U4315, new_P2_U4316,
    new_P2_U4317, new_P2_U4318, new_P2_U4319, new_P2_U4320, new_P2_U4321,
    new_P2_U4322, new_P2_U4323, new_P2_U4324, new_P2_U4325, new_P2_U4326,
    new_P2_U4327, new_P2_U4328, new_P2_U4329, new_P2_U4330, new_P2_U4331,
    new_P2_U4332, new_P2_U4333, new_P2_U4334, new_P2_U4335, new_P2_U4336,
    new_P2_U4337, new_P2_U4338, new_P2_U4339, new_P2_U4340, new_P2_U4341,
    new_P2_U4342, new_P2_U4343, new_P2_U4344, new_P2_U4345, new_P2_U4346,
    new_P2_U4347, new_P2_U4348, new_P2_U4349, new_P2_U4350, new_P2_U4351,
    new_P2_U4352, new_P2_U4353, new_P2_U4354, new_P2_U4355, new_P2_U4356,
    new_P2_U4357, new_P2_U4358, new_P2_U4359, new_P2_U4360, new_P2_U4361,
    new_P2_U4362, new_P2_U4363, new_P2_U4364, new_P2_U4365, new_P2_U4366,
    new_P2_U4367, new_P2_U4368, new_P2_U4369, new_P2_U4370, new_P2_U4371,
    new_P2_U4372, new_P2_U4373, new_P2_U4374, new_P2_U4375, new_P2_U4376,
    new_P2_U4377, new_P2_U4378, new_P2_U4379, new_P2_U4380, new_P2_U4381,
    new_P2_U4382, new_P2_U4383, new_P2_U4384, new_P2_U4385, new_P2_U4386,
    new_P2_U4387, new_P2_U4388, new_P2_U4389, new_P2_U4390, new_P2_U4391,
    new_P2_U4392, new_P2_U4393, new_P2_U4394, new_P2_U4395, new_P2_U4396,
    new_P2_U4397, new_P2_U4398, new_P2_U4399, new_P2_U4400, new_P2_U4401,
    new_P2_U4402, new_P2_U4403, new_P2_U4404, new_P2_U4405, new_P2_U4406,
    new_P2_U4407, new_P2_U4408, new_P2_U4409, new_P2_U4410, new_P2_U4411,
    new_P2_U4412, new_P2_U4413, new_P2_U4414, new_P2_U4415, new_P2_U4416,
    new_P2_U4417, new_P2_U4418, new_P2_U4419, new_P2_U4420, new_P2_U4421,
    new_P2_U4422, new_P2_U4423, new_P2_U4424, new_P2_U4425, new_P2_U4426,
    new_P2_U4427, new_P2_U4428, new_P2_U4429, new_P2_U4430, new_P2_U4431,
    new_P2_U4432, new_P2_U4433, new_P2_U4434, new_P2_U4435, new_P2_U4436,
    new_P2_U4437, new_P2_U4438, new_P2_U4439, new_P2_U4440, new_P2_U4441,
    new_P2_U4442, new_P2_U4443, new_P2_U4444, new_P2_U4445, new_P2_U4446,
    new_P2_U4447, new_P2_U4448, new_P2_U4449, new_P2_U4450, new_P2_U4451,
    new_P2_U4452, new_P2_U4453, new_P2_U4454, new_P2_U4455, new_P2_U4456,
    new_P2_U4457, new_P2_U4458, new_P2_U4459, new_P2_U4460, new_P2_U4461,
    new_P2_U4462, new_P2_U4463, new_P2_U4464, new_P2_U4465, new_P2_U4466,
    new_P2_U4467, new_P2_U4468, new_P2_U4469, new_P2_U4470, new_P2_U4471,
    new_P2_U4472, new_P2_U4473, new_P2_U4474, new_P2_U4475, new_P2_U4476,
    new_P2_U4477, new_P2_U4478, new_P2_U4479, new_P2_U4480, new_P2_U4481,
    new_P2_U4482, new_P2_U4483, new_P2_U4484, new_P2_U4485, new_P2_U4486,
    new_P2_U4487, new_P2_U4488, new_P2_U4489, new_P2_U4490, new_P2_U4491,
    new_P2_U4492, new_P2_U4493, new_P2_U4494, new_P2_U4495, new_P2_U4496,
    new_P2_U4497, new_P2_U4498, new_P2_U4499, new_P2_U4500, new_P2_U4501,
    new_P2_U4502, new_P2_U4503, new_P2_U4504, new_P2_U4505, new_P2_U4506,
    new_P2_U4507, new_P2_U4508, new_P2_U4509, new_P2_U4510, new_P2_U4511,
    new_P2_U4512, new_P2_U4513, new_P2_U4514, new_P2_U4515, new_P2_U4516,
    new_P2_U4517, new_P2_U4518, new_P2_U4519, new_P2_U4520, new_P2_U4521,
    new_P2_U4522, new_P2_U4523, new_P2_U4524, new_P2_U4525, new_P2_U4526,
    new_P2_U4527, new_P2_U4528, new_P2_U4529, new_P2_U4530, new_P2_U4531,
    new_P2_U4532, new_P2_U4533, new_P2_U4534, new_P2_U4535, new_P2_U4536,
    new_P2_U4537, new_P2_U4538, new_P2_U4539, new_P2_U4540, new_P2_U4541,
    new_P2_U4542, new_P2_U4543, new_P2_U4544, new_P2_U4545, new_P2_U4546,
    new_P2_U4547, new_P2_U4548, new_P2_U4549, new_P2_U4550, new_P2_U4551,
    new_P2_U4552, new_P2_U4553, new_P2_U4554, new_P2_U4555, new_P2_U4556,
    new_P2_U4557, new_P2_U4558, new_P2_U4559, new_P2_U4560, new_P2_U4561,
    new_P2_U4562, new_P2_U4563, new_P2_U4564, new_P2_U4565, new_P2_U4566,
    new_P2_U4567, new_P2_U4568, new_P2_U4569, new_P2_U4570, new_P2_U4571,
    new_P2_U4572, new_P2_U4573, new_P2_U4574, new_P2_U4575, new_P2_U4576,
    new_P2_U4577, new_P2_U4578, new_P2_U4579, new_P2_U4580, new_P2_U4581,
    new_P2_U4582, new_P2_U4583, new_P2_U4584, new_P2_U4585, new_P2_U4586,
    new_P2_U4587, new_P2_U4588, new_P2_U4589, new_P2_U4590, new_P2_U4591,
    new_P2_U4592, new_P2_U4593, new_P2_U4594, new_P2_U4595, new_P2_U4596,
    new_P2_U4597, new_P2_U4598, new_P2_U4599, new_P2_U4600, new_P2_U4601,
    new_P2_U4602, new_P2_U4603, new_P2_U4604, new_P2_U4605, new_P2_U4606,
    new_P2_U4607, new_P2_U4608, new_P2_U4609, new_P2_U4610, new_P2_U4611,
    new_P2_U4612, new_P2_U4613, new_P2_U4614, new_P2_U4615, new_P2_U4616,
    new_P2_U4617, new_P2_U4618, new_P2_U4619, new_P2_U4620, new_P2_U4621,
    new_P2_U4622, new_P2_U4623, new_P2_U4624, new_P2_U4625, new_P2_U4626,
    new_P2_U4627, new_P2_U4628, new_P2_U4629, new_P2_U4630, new_P2_U4631,
    new_P2_U4632, new_P2_U4633, new_P2_U4634, new_P2_U4635, new_P2_U4636,
    new_P2_U4637, new_P2_U4638, new_P2_U4639, new_P2_U4640, new_P2_U4641,
    new_P2_U4642, new_P2_U4643, new_P2_U4644, new_P2_U4645, new_P2_U4646,
    new_P2_U4647, new_P2_U4648, new_P2_U4649, new_P2_U4650, new_P2_U4651,
    new_P2_U4652, new_P2_U4653, new_P2_U4654, new_P2_U4655, new_P2_U4656,
    new_P2_U4657, new_P2_U4658, new_P2_U4659, new_P2_U4660, new_P2_U4661,
    new_P2_U4662, new_P2_U4663, new_P2_U4664, new_P2_U4665, new_P2_U4666,
    new_P2_U4667, new_P2_U4668, new_P2_U4669, new_P2_U4670, new_P2_U4671,
    new_P2_U4672, new_P2_U4673, new_P2_U4674, new_P2_U4675, new_P2_U4676,
    new_P2_U4677, new_P2_U4678, new_P2_U4679, new_P2_U4680, new_P2_U4681,
    new_P2_U4682, new_P2_U4683, new_P2_U4684, new_P2_U4685, new_P2_U4686,
    new_P2_U4687, new_P2_U4688, new_P2_U4689, new_P2_U4690, new_P2_U4691,
    new_P2_U4692, new_P2_U4693, new_P2_U4694, new_P2_U4695, new_P2_U4696,
    new_P2_U4697, new_P2_U4698, new_P2_U4699, new_P2_U4700, new_P2_U4701,
    new_P2_U4702, new_P2_U4703, new_P2_U4704, new_P2_U4705, new_P2_U4706,
    new_P2_U4707, new_P2_U4708, new_P2_U4709, new_P2_U4710, new_P2_U4711,
    new_P2_U4712, new_P2_U4713, new_P2_U4714, new_P2_U4715, new_P2_U4716,
    new_P2_U4717, new_P2_U4718, new_P2_U4719, new_P2_U4720, new_P2_U4721,
    new_P2_U4722, new_P2_U4723, new_P2_U4724, new_P2_U4725, new_P2_U4726,
    new_P2_U4727, new_P2_U4728, new_P2_U4729, new_P2_U4730, new_P2_U4731,
    new_P2_U4732, new_P2_U4733, new_P2_U4734, new_P2_U4735, new_P2_U4736,
    new_P2_U4737, new_P2_U4738, new_P2_U4739, new_P2_U4740, new_P2_U4741,
    new_P2_U4742, new_P2_U4743, new_P2_U4744, new_P2_U4745, new_P2_U4746,
    new_P2_U4747, new_P2_U4748, new_P2_U4749, new_P2_U4750, new_P2_U4751,
    new_P2_U4752, new_P2_U4753, new_P2_U4754, new_P2_U4755, new_P2_U4756,
    new_P2_U4757, new_P2_U4758, new_P2_U4759, new_P2_U4760, new_P2_U4761,
    new_P2_U4762, new_P2_U4763, new_P2_U4764, new_P2_U4765, new_P2_U4766,
    new_P2_U4767, new_P2_U4768, new_P2_U4769, new_P2_U4770, new_P2_U4771,
    new_P2_U4772, new_P2_U4773, new_P2_U4774, new_P2_U4775, new_P2_U4776,
    new_P2_U4777, new_P2_U4778, new_P2_U4779, new_P2_U4780, new_P2_U4781,
    new_P2_U4782, new_P2_U4783, new_P2_U4784, new_P2_U4785, new_P2_U4786,
    new_P2_U4787, new_P2_U4788, new_P2_U4789, new_P2_U4790, new_P2_U4791,
    new_P2_U4792, new_P2_U4793, new_P2_U4794, new_P2_U4795, new_P2_U4796,
    new_P2_U4797, new_P2_U4798, new_P2_U4799, new_P2_U4800, new_P2_U4801,
    new_P2_U4802, new_P2_U4803, new_P2_U4804, new_P2_U4805, new_P2_U4806,
    new_P2_U4807, new_P2_U4808, new_P2_U4809, new_P2_U4810, new_P2_U4811,
    new_P2_U4812, new_P2_U4813, new_P2_U4814, new_P2_U4815, new_P2_U4816,
    new_P2_U4817, new_P2_U4818, new_P2_U4819, new_P2_U4820, new_P2_U4821,
    new_P2_U4822, new_P2_U4823, new_P2_U4824, new_P2_U4825, new_P2_U4826,
    new_P2_U4827, new_P2_U4828, new_P2_U4829, new_P2_U4830, new_P2_U4831,
    new_P2_U4832, new_P2_U4833, new_P2_U4834, new_P2_U4835, new_P2_U4836,
    new_P2_U4837, new_P2_U4838, new_P2_U4839, new_P2_U4840, new_P2_U4841,
    new_P2_U4842, new_P2_U4843, new_P2_U4844, new_P2_U4845, new_P2_U4846,
    new_P2_U4847, new_P2_U4848, new_P2_U4849, new_P2_U4850, new_P2_U4851,
    new_P2_U4852, new_P2_U4853, new_P2_U4854, new_P2_U4855, new_P2_U4856,
    new_P2_U4857, new_P2_U4858, new_P2_U4859, new_P2_U4860, new_P2_U4861,
    new_P2_U4862, new_P2_U4863, new_P2_U4864, new_P2_U4865, new_P2_U4866,
    new_P2_U4867, new_P2_U4868, new_P2_U4869, new_P2_U4870, new_P2_U4871,
    new_P2_U4872, new_P2_U4873, new_P2_U4874, new_P2_U4875, new_P2_U4876,
    new_P2_U4877, new_P2_U4878, new_P2_U4879, new_P2_U4880, new_P2_U4881,
    new_P2_U4882, new_P2_U4883, new_P2_U4884, new_P2_U4885, new_P2_U4886,
    new_P2_U4887, new_P2_U4888, new_P2_U4889, new_P2_U4890, new_P2_U4891,
    new_P2_U4892, new_P2_U4893, new_P2_U4894, new_P2_U4895, new_P2_U4896,
    new_P2_U4897, new_P2_U4898, new_P2_U4899, new_P2_U4900, new_P2_U4901,
    new_P2_U4902, new_P2_U4903, new_P2_U4904, new_P2_U4905, new_P2_U4906,
    new_P2_U4907, new_P2_U4908, new_P2_U4909, new_P2_U4910, new_P2_U4911,
    new_P2_U4912, new_P2_U4913, new_P2_U4914, new_P2_U4915, new_P2_U4916,
    new_P2_U4917, new_P2_U4918, new_P2_U4919, new_P2_U4920, new_P2_U4921,
    new_P2_U4922, new_P2_U4923, new_P2_U4924, new_P2_U4925, new_P2_U4926,
    new_P2_U4927, new_P2_U4928, new_P2_U4929, new_P2_U4930, new_P2_U4931,
    new_P2_U4932, new_P2_U4933, new_P2_U4934, new_P2_U4935, new_P2_U4936,
    new_P2_U4937, new_P2_U4938, new_P2_U4939, new_P2_U4940, new_P2_U4941,
    new_P2_U4942, new_P2_U4943, new_P2_U4944, new_P2_U4945, new_P2_U4946,
    new_P2_U4947, new_P2_U4948, new_P2_U4949, new_P2_U4950, new_P2_U4951,
    new_P2_U4952, new_P2_U4953, new_P2_U4954, new_P2_U4955, new_P2_U4956,
    new_P2_U4957, new_P2_U4958, new_P2_U4959, new_P2_U4960, new_P2_U4961,
    new_P2_U4962, new_P2_U4963, new_P2_U4964, new_P2_U4965, new_P2_U4966,
    new_P2_U4967, new_P2_U4968, new_P2_U4969, new_P2_U4970, new_P2_U4971,
    new_P2_U4972, new_P2_U4973, new_P2_U4974, new_P2_U4975, new_P2_U4976,
    new_P2_U4977, new_P2_U4978, new_P2_U4979, new_P2_U4980, new_P2_U4981,
    new_P2_U4982, new_P2_U4983, new_P2_U4984, new_P2_U4985, new_P2_U4986,
    new_P2_U4987, new_P2_U4988, new_P2_U4989, new_P2_U4990, new_P2_U4991,
    new_P2_U4992, new_P2_U4993, new_P2_U4994, new_P2_U4995, new_P2_U4996,
    new_P2_U4997, new_P2_U4998, new_P2_U4999, new_P2_U5000, new_P2_U5001,
    new_P2_U5002, new_P2_U5003, new_P2_U5004, new_P2_U5005, new_P2_U5006,
    new_P2_U5007, new_P2_U5008, new_P2_U5009, new_P2_U5010, new_P2_U5011,
    new_P2_U5012, new_P2_U5013, new_P2_U5014, new_P2_U5015, new_P2_U5016,
    new_P2_U5017, new_P2_U5018, new_P2_U5019, new_P2_U5020, new_P2_U5021,
    new_P2_U5022, new_P2_U5023, new_P2_U5024, new_P2_U5025, new_P2_U5026,
    new_P2_U5027, new_P2_U5028, new_P2_U5029, new_P2_U5030, new_P2_U5031,
    new_P2_U5032, new_P2_U5033, new_P2_U5034, new_P2_U5035, new_P2_U5036,
    new_P2_U5037, new_P2_U5038, new_P2_U5039, new_P2_U5040, new_P2_U5041,
    new_P2_U5042, new_P2_U5043, new_P2_U5044, new_P2_U5045, new_P2_U5046,
    new_P2_U5047, new_P2_U5048, new_P2_U5049, new_P2_U5050, new_P2_U5051,
    new_P2_U5052, new_P2_U5053, new_P2_U5054, new_P2_U5055, new_P2_U5056,
    new_P2_U5057, new_P2_U5058, new_P2_U5059, new_P2_U5060, new_P2_U5061,
    new_P2_U5062, new_P2_U5063, new_P2_U5064, new_P2_U5065, new_P2_U5066,
    new_P2_U5067, new_P2_U5068, new_P2_U5069, new_P2_U5070, new_P2_U5071,
    new_P2_U5072, new_P2_U5073, new_P2_U5074, new_P2_U5075, new_P2_U5076,
    new_P2_U5077, new_P2_U5078, new_P2_U5079, new_P2_U5080, new_P2_U5081,
    new_P2_U5082, new_P2_U5083, new_P2_U5084, new_P2_U5085, new_P2_U5086,
    new_P2_U5087, new_P2_U5088, new_P2_U5089, new_P2_U5090, new_P2_U5091,
    new_P2_U5092, new_P2_U5093, new_P2_U5094, new_P2_U5095, new_P2_U5096,
    new_P2_U5097, new_P2_U5098, new_P2_U5099, new_P2_U5100, new_P2_U5101,
    new_P2_U5102, new_P2_U5103, new_P2_U5104, new_P2_U5105, new_P2_U5106,
    new_P2_U5107, new_P2_U5108, new_P2_U5109, new_P2_U5110, new_P2_U5111,
    new_P2_U5112, new_P2_U5113, new_P2_U5114, new_P2_U5115, new_P2_U5116,
    new_P2_U5117, new_P2_U5118, new_P2_U5119, new_P2_U5120, new_P2_U5121,
    new_P2_U5122, new_P2_U5123, new_P2_U5124, new_P2_U5125, new_P2_U5126,
    new_P2_U5127, new_P2_U5128, new_P2_U5129, new_P2_U5130, new_P2_U5131,
    new_P2_U5132, new_P2_U5133, new_P2_U5134, new_P2_U5135, new_P2_U5136,
    new_P2_U5137, new_P2_U5138, new_P2_U5139, new_P2_U5140, new_P2_U5141,
    new_P2_U5142, new_P2_U5143, new_P2_U5144, new_P2_U5145, new_P2_U5146,
    new_P2_U5147, new_P2_U5148, new_P2_U5149, new_P2_U5150, new_P2_U5151,
    new_P2_U5152, new_P2_U5153, new_P2_U5154, new_P2_U5155, new_P2_U5156,
    new_P2_U5157, new_P2_U5158, new_P2_U5159, new_P2_U5160, new_P2_U5161,
    new_P2_U5162, new_P2_U5163, new_P2_U5164, new_P2_U5165, new_P2_U5166,
    new_P2_U5167, new_P2_U5168, new_P2_U5169, new_P2_U5170, new_P2_U5171,
    new_P2_U5172, new_P2_U5173, new_P2_U5174, new_P2_U5175, new_P2_U5176,
    new_P2_U5177, new_P2_U5178, new_P2_U5179, new_P2_U5180, new_P2_U5181,
    new_P2_U5182, new_P2_U5183, new_P2_U5184, new_P2_U5185, new_P2_U5186,
    new_P2_U5187, new_P2_U5188, new_P2_U5189, new_P2_U5190, new_P2_U5191,
    new_P2_U5192, new_P2_U5193, new_P2_U5194, new_P2_U5195, new_P2_U5196,
    new_P2_U5197, new_P2_U5198, new_P2_U5199, new_P2_U5200, new_P2_U5201,
    new_P2_U5202, new_P2_U5203, new_P2_U5204, new_P2_U5205, new_P2_U5206,
    new_P2_U5207, new_P2_U5208, new_P2_U5209, new_P2_U5210, new_P2_U5211,
    new_P2_U5212, new_P2_U5213, new_P2_U5214, new_P2_U5215, new_P2_U5216,
    new_P2_U5217, new_P2_U5218, new_P2_U5219, new_P2_U5220, new_P2_U5221,
    new_P2_U5222, new_P2_U5223, new_P2_U5224, new_P2_U5225, new_P2_U5226,
    new_P2_U5227, new_P2_U5228, new_P2_U5229, new_P2_U5230, new_P2_U5231,
    new_P2_U5232, new_P2_U5233, new_P2_U5234, new_P2_U5235, new_P2_U5236,
    new_P2_U5237, new_P2_U5238, new_P2_U5239, new_P2_U5240, new_P2_U5241,
    new_P2_U5242, new_P2_U5243, new_P2_U5244, new_P2_U5245, new_P2_U5246,
    new_P2_U5247, new_P2_U5248, new_P2_U5249, new_P2_U5250, new_P2_U5251,
    new_P2_U5252, new_P2_U5253, new_P2_U5254, new_P2_U5255, new_P2_U5256,
    new_P2_U5257, new_P2_U5258, new_P2_U5259, new_P2_U5260, new_P2_U5261,
    new_P2_U5262, new_P2_U5263, new_P2_U5264, new_P2_U5265, new_P2_U5266,
    new_P2_U5267, new_P2_U5268, new_P2_U5269, new_P2_U5270, new_P2_U5271,
    new_P2_U5272, new_P2_U5273, new_P2_U5274, new_P2_U5275, new_P2_U5276,
    new_P2_U5277, new_P2_U5278, new_P2_U5279, new_P2_U5280, new_P2_U5281,
    new_P2_U5282, new_P2_U5283, new_P2_U5284, new_P2_U5285, new_P2_U5286,
    new_P2_U5287, new_P2_U5288, new_P2_U5289, new_P2_U5290, new_P2_U5291,
    new_P2_U5292, new_P2_U5293, new_P2_U5294, new_P2_U5295, new_P2_U5296,
    new_P2_U5297, new_P2_U5298, new_P2_U5299, new_P2_U5300, new_P2_U5301,
    new_P2_U5302, new_P2_U5303, new_P2_U5304, new_P2_U5305, new_P2_U5306,
    new_P2_U5307, new_P2_U5308, new_P2_U5309, new_P2_U5310, new_P2_U5311,
    new_P2_U5312, new_P2_U5313, new_P2_U5314, new_P2_U5315, new_P2_U5316,
    new_P2_U5317, new_P2_U5318, new_P2_U5319, new_P2_U5320, new_P2_U5321,
    new_P2_U5322, new_P2_U5323, new_P2_U5324, new_P2_U5325, new_P2_U5326,
    new_P2_U5327, new_P2_U5328, new_P2_U5329, new_P2_U5330, new_P2_U5331,
    new_P2_U5332, new_P2_U5333, new_P2_U5334, new_P2_U5335, new_P2_U5336,
    new_P2_U5337, new_P2_U5338, new_P2_U5339, new_P2_U5340, new_P2_U5341,
    new_P2_U5342, new_P2_U5343, new_P2_U5344, new_P2_U5345, new_P2_U5346,
    new_P2_U5347, new_P2_U5348, new_P2_U5349, new_P2_U5350, new_P2_U5351,
    new_P2_U5352, new_P2_U5353, new_P2_U5354, new_P2_U5355, new_P2_U5356,
    new_P2_U5357, new_P2_U5358, new_P2_U5359, new_P2_U5360, new_P2_U5361,
    new_P2_U5362, new_P2_U5363, new_P2_U5364, new_P2_U5365, new_P2_U5366,
    new_P2_U5367, new_P2_U5368, new_P2_U5369, new_P2_U5370, new_P2_U5371,
    new_P2_U5372, new_P2_U5373, new_P2_U5374, new_P2_U5375, new_P2_U5376,
    new_P2_U5377, new_P2_U5378, new_P2_U5379, new_P2_U5380, new_P2_U5381,
    new_P2_U5382, new_P2_U5383, new_P2_U5384, new_P2_U5385, new_P2_U5386,
    new_P2_U5387, new_P2_U5388, new_P2_U5389, new_P2_U5390, new_P2_U5391,
    new_P2_U5392, new_P2_U5393, new_P2_U5394, new_P2_U5395, new_P2_U5396,
    new_P2_U5397, new_P2_U5398, new_P2_U5399, new_P2_U5400, new_P2_U5401,
    new_P2_U5402, new_P2_U5403, new_P2_U5404, new_P2_U5405, new_P2_U5406,
    new_P2_U5407, new_P2_U5408, new_P2_U5409, new_P2_U5410, new_P2_U5411,
    new_P2_U5412, new_P2_U5413, new_P2_U5414, new_P2_U5415, new_P2_U5416,
    new_P2_U5417, new_P2_U5418, new_P2_U5419, new_P2_U5420, new_P2_U5421,
    new_P2_U5422, new_P2_U5423, new_P2_U5424, new_P2_U5425, new_P2_U5426,
    new_P2_U5427, new_P2_U5428, new_P2_U5429, new_P2_U5430, new_P2_U5431,
    new_P2_U5432, new_P2_U5433, new_P2_U5434, new_P2_U5435, new_P2_U5436,
    new_P2_U5437, new_P2_U5438, new_P2_U5439, new_P2_U5440, new_P2_U5441,
    new_P2_U5442, new_P2_U5443, new_P2_U5444, new_P2_U5445, new_P2_U5446,
    new_P2_U5447, new_P2_U5448, new_P2_U5449, new_P2_U5450, new_P2_U5451,
    new_P2_U5452, new_P2_U5453, new_P2_U5454, new_P2_U5455, new_P2_U5456,
    new_P2_U5457, new_P2_U5458, new_P2_U5459, new_P2_U5460, new_P2_U5461,
    new_P2_U5462, new_P2_U5463, new_P2_U5464, new_P2_U5465, new_P2_U5466,
    new_P2_U5467, new_P2_U5468, new_P2_U5469, new_P2_U5470, new_P2_U5471,
    new_P2_U5472, new_P2_U5473, new_P2_U5474, new_P2_U5475, new_P2_U5476,
    new_P2_U5477, new_P2_U5478, new_P2_U5479, new_P2_U5480, new_P2_U5481,
    new_P2_U5482, new_P2_U5483, new_P2_U5484, new_P2_U5485, new_P2_U5486,
    new_P2_U5487, new_P2_U5488, new_P2_U5489, new_P2_U5490, new_P2_U5491,
    new_P2_U5492, new_P2_U5493, new_P2_U5494, new_P2_U5495, new_P2_U5496,
    new_P2_U5497, new_P2_U5498, new_P2_U5499, new_P2_U5500, new_P2_U5501,
    new_P2_U5502, new_P2_U5503, new_P2_U5504, new_P2_U5505, new_P2_U5506,
    new_P2_U5507, new_P2_U5508, new_P2_U5509, new_P2_U5510, new_P2_U5511,
    new_P2_U5512, new_P2_U5513, new_P2_U5514, new_P2_U5515, new_P2_U5516,
    new_P2_U5517, new_P2_U5518, new_P2_U5519, new_P2_U5520, new_P2_U5521,
    new_P2_U5522, new_P2_U5523, new_P2_U5524, new_P2_U5525, new_P2_U5526,
    new_P2_U5527, new_P2_U5528, new_P2_U5529, new_P2_U5530, new_P2_U5531,
    new_P2_U5532, new_P2_U5533, new_P2_U5534, new_P2_U5535, new_P2_U5536,
    new_P2_U5537, new_P2_U5538, new_P2_U5539, new_P2_U5540, new_P2_U5541,
    new_P2_U5542, new_P2_U5543, new_P2_U5544, new_P2_U5545, new_P2_U5546,
    new_P2_U5547, new_P2_U5548, new_P2_U5549, new_P2_U5550, new_P2_U5551,
    new_P2_U5552, new_P2_U5553, new_P2_U5554, new_P2_U5555, new_P2_U5556,
    new_P2_U5557, new_P2_U5558, new_P2_U5559, new_P2_U5560, new_P2_U5561,
    new_P2_U5562, new_P2_U5563, new_P2_U5564, new_P2_U5565, new_P2_U5566,
    new_P2_U5567, new_P2_U5568, new_P2_U5569, new_P2_U5570, new_P2_U5571,
    new_P2_U5572, new_P2_U5573, new_P2_U5574, new_P2_U5575, new_P2_U5576,
    new_P2_U5577, new_P2_U5578, new_P2_U5579, new_P2_U5580, new_P2_U5581,
    new_P2_U5582, new_P2_U5583, new_P2_U5584, new_P2_U5585, new_P2_U5586,
    new_P2_U5587, new_P2_U5588, new_P2_U5589, new_P2_U5590, new_P2_U5591,
    new_P2_U5592, new_P2_U5593, new_P2_U5594, new_P2_U5595, new_P2_U5596,
    new_P2_U5597, new_P2_U5598, new_P2_U5599, new_P2_U5600, new_P2_U5601,
    new_P2_U5602, new_P2_U5603, new_P2_U5604, new_P2_U5605, new_P2_U5606,
    new_P2_U5607, new_P2_U5608, new_P2_U5609, new_P2_U5610, new_P2_U5611,
    new_P2_U5612, new_P2_U5613, new_P2_U5614, new_P2_U5615, new_P2_U5616,
    new_P2_U5617, new_P2_U5618, new_P2_U5619, new_P2_U5620, new_P2_U5621,
    new_P2_U5622, new_P2_U5623, new_P2_U5624, new_P2_U5625, new_P2_U5626,
    new_P2_U5627, new_P2_U5628, new_P2_U5629, new_P2_U5630, new_P2_U5631,
    new_P2_U5632, new_P2_U5633, new_P2_U5634, new_P2_U5635, new_P2_U5636,
    new_P2_U5637, new_P2_U5638, new_P2_U5639, new_P2_U5640, new_P2_U5641,
    new_P2_U5642, new_P2_U5643, new_P2_U5644, new_P2_U5645, new_P2_U5646,
    new_P2_U5647, new_P2_U5648, new_P2_U5649, new_P2_U5650, new_P2_U5651,
    new_P2_U5652, new_P2_U5653, new_P2_U5654, new_P2_U5655, new_P2_U5656,
    new_P2_U5657, new_P2_U5658, new_P2_U5659, new_P2_U5660, new_P2_U5661,
    new_P2_U5662, new_P2_U5663, new_P2_U5664, new_P2_U5665, new_P2_U5666,
    new_P2_U5667, new_P2_U5668, new_P2_U5669, new_P2_U5670, new_P2_U5671,
    new_P2_U5672, new_P2_U5673, new_P2_U5674, new_P2_U5675, new_P2_U5676,
    new_P2_U5677, new_P2_U5678, new_P2_U5679, new_P2_U5680, new_P2_U5681,
    new_P2_U5682, new_P2_U5683, new_P2_U5684, new_P2_U5685, new_P2_U5686,
    new_P2_U5687, new_P2_U5688, new_P2_U5689, new_P2_U5690, new_P2_U5691,
    new_P2_U5692, new_P2_U5693, new_P2_U5694, new_P2_U5695, new_P2_U5696,
    new_P2_U5697, new_P2_U5698, new_P2_U5699, new_P2_U5700, new_P2_U5701,
    new_P2_U5702, new_P2_U5703, new_P2_U5704, new_P2_U5705, new_P2_U5706,
    new_P2_U5707, new_P2_U5708, new_P2_U5709, new_P2_U5710, new_P2_U5711,
    new_P2_U5712, new_P2_U5713, new_P2_U5714, new_P2_U5715, new_P2_U5716,
    new_P2_U5717, new_P2_U5718, new_P2_U5719, new_P2_U5720, new_P2_U5721,
    new_P2_U5722, new_P2_U5723, new_P2_U5724, new_P2_U5725, new_P2_U5726,
    new_P2_U5727, new_P2_U5728, new_P2_U5729, new_P2_U5730, new_P2_U5731,
    new_P2_U5732, new_P2_U5733, new_P2_U5734, new_P2_U5735, new_P2_U5736,
    new_P2_U5737, new_P2_U5738, new_P2_U5739, new_P2_U5740, new_P2_U5741,
    new_P2_U5742, new_P2_U5743, new_P2_U5744, new_P2_U5745, new_P2_U5746,
    new_P2_U5747, new_P2_U5748, new_P2_U5749, new_P2_U5750, new_P2_U5751,
    new_P2_U5752, new_P2_U5753, new_P2_U5754, new_P2_U5755, new_P2_U5756,
    new_P2_U5757, new_P2_U5758, new_P2_U5759, new_P2_U5760, new_P2_U5761,
    new_P2_U5762, new_P2_U5763, new_P2_U5764, new_P2_U5765, new_P2_U5766,
    new_P2_U5767, new_P2_U5768, new_P2_U5769, new_P2_U5770, new_P2_U5771,
    new_P2_U5772, new_P2_U5773, new_P2_U5774, new_P2_U5775, new_P2_U5776,
    new_P2_U5777, new_P2_U5778, new_P2_U5779, new_P2_U5780, new_P2_U5781,
    new_P2_U5782, new_P2_U5783, new_P2_U5784, new_P2_U5785, new_P2_U5786,
    new_P2_U5787, new_P2_U5788, new_P2_U5789, new_P2_U5790, new_P2_U5791,
    new_P2_U5792, new_P2_U5793, new_P2_U5794, new_P2_U5795, new_P2_U5796,
    new_P2_U5797, new_P2_U5798, new_P2_U5799, new_P2_U5800, new_P2_U5801,
    new_P2_U5802, new_P2_U5803, new_P2_U5804, new_P2_U5805, new_P2_U5806,
    new_P2_U5807, new_P2_U5808, new_P2_U5809, new_P2_U5810, new_P2_U5811,
    new_P2_U5812, new_P2_U5813, new_P2_U5814, new_P2_U5815, new_P2_U5816,
    new_P2_U5817, new_P2_U5818, new_P2_U5819, new_P2_U5820, new_P2_U5821,
    new_P2_U5822, new_P2_U5823, new_P2_U5824, new_P2_U5825, new_P2_U5826,
    new_P2_U5827, new_P2_U5828, new_P2_U5829, new_P2_U5830, new_P2_U5831,
    new_P2_U5832, new_P2_U5833, new_P2_U5834, new_P2_U5835, new_P2_U5836,
    new_P2_U5837, new_P2_U5838, new_P2_U5839, new_P2_U5840, new_P2_U5841,
    new_P2_U5842, new_P2_U5843, new_P2_U5844, new_P2_U5845, new_P2_U5846,
    new_P2_U5847, new_P2_U5848, new_P2_U5849, new_P2_U5850, new_P2_U5851,
    new_P2_U5852, new_P2_U5853, new_P2_U5854, new_P2_U5855, new_P2_U5856,
    new_P2_U5857, new_P2_U5858, new_P2_U5859, new_P2_U5860, new_P2_U5861,
    new_P2_U5862, new_P2_U5863, new_P2_U5864, new_P2_U5865, new_P2_U5866,
    new_P2_U5867, new_P2_U5868, new_P2_U5869, new_P2_U5870, new_P2_U5871,
    new_P2_U5872, new_P2_U5873, new_P2_U5874, new_P2_U5875, new_P2_U5876,
    new_P2_U5877, new_P2_U5878, new_P2_U5879, new_P2_U5880, new_P2_U5881,
    new_P2_U5882, new_P2_U5883, new_P2_U5884, new_P2_U5885, new_P2_U5886,
    new_P2_U5887, new_P2_U5888, new_P2_U5889, new_P2_U5890, new_P2_U5891,
    new_P2_U5892, new_P2_U5893, new_P2_U5894, new_P2_U5895, new_P2_U5896,
    new_P2_U5897, new_P2_U5898, new_P2_U5899, new_P2_U5900, new_P2_U5901,
    new_P2_U5902, new_P2_U5903, new_P2_U5904, new_P2_U5905, new_P2_U5906,
    new_P2_U5907, new_P2_U5908, new_P2_U5909, new_P2_U5910, new_P2_U5911,
    new_P2_U5912, new_P2_U5913, new_P2_U5914, new_P2_U5915, new_P2_U5916,
    new_P2_U5917, new_P2_U5918, new_P2_U5919, new_P2_U5920, new_P2_U5921,
    new_P2_U5922, new_P2_U5923, new_P2_U5924, new_P2_U5925, new_P2_U5926,
    new_P2_U5927, new_P2_U5928, new_P2_U5929, new_P2_U5930, new_P2_U5931,
    new_P2_U5932, new_P2_U5933, new_P2_U5934, new_P2_U5935, new_P2_U5936,
    new_P2_U5937, new_P2_U5938, new_P2_U5939, new_P2_U5940, new_P2_U5941,
    new_P2_U5942, new_P2_U5943, new_P2_U5944, new_P2_U5945, new_P2_U5946,
    new_P2_U5947, new_P2_U5948, new_P2_U5949, new_P2_U5950, new_P2_U5951,
    new_P2_U5952, new_P2_U5953, new_P2_U5954, new_P2_U5955, new_P2_U5956,
    new_P2_U5957, new_P2_U5958, new_P2_U5959, new_P2_U5960, new_P2_U5961,
    new_P2_U5962, new_P2_U5963, new_P2_U5964, new_P2_U5965, new_P2_U5966,
    new_P2_U5967, new_P2_U5968, new_P2_U5969, new_P2_U5970, new_P2_U5971,
    new_P2_U5972, new_P2_U5973, new_P2_U5974, new_P2_U5975, new_P2_U5976,
    new_P2_U5977, new_P2_U5978, new_P2_U5979, new_P2_U5980, new_P2_U5981,
    new_P2_U5982, new_P2_U5983, new_P2_U5984, new_P2_U5985, new_P2_U5986,
    new_P2_U5987, new_P2_U5988, new_P2_U5989, new_P2_U5990, new_P2_U5991,
    new_P2_U5992, new_P2_U5993, new_P2_U5994, new_P2_U5995, new_P2_U5996,
    new_P2_U5997, new_P2_U5998, new_P2_U5999, new_P2_U6000, new_P2_U6001,
    new_P2_U6002, new_P2_U6003, new_P2_U6004, new_P2_U6005, new_P2_U6006,
    new_P2_U6007, new_P2_U6008, new_P2_U6009, new_P2_U6010, new_P2_U6011,
    new_P2_U6012, new_P2_U6013, new_P2_U6014, new_P2_U6015, new_P2_U6016,
    new_P2_U6017, new_P2_U6018, new_P2_U6019, new_P2_U6020, new_P2_U6021,
    new_P2_U6022, new_P2_U6023, new_P2_U6024, new_P2_U6025, new_P2_U6026,
    new_P2_U6027, new_P2_U6028, new_P2_U6029, new_P2_U6030, new_P2_U6031,
    new_P2_U6032, new_P2_U6033, new_P2_U6034, new_P2_U6035, new_P2_U6036,
    new_P2_U6037, new_P2_U6038, new_P2_U6039, new_P2_U6040, new_P2_U6041,
    new_P2_U6042, new_P2_U6043, new_P2_U6044, new_P2_U6045, new_P2_U6046,
    new_P2_U6047, new_P2_U6048, new_P2_U6049, new_P2_U6050, new_P2_U6051,
    new_P2_U6052, new_P2_U6053, new_P2_U6054, new_P2_U6055, new_P2_U6056,
    new_P2_U6057, new_P2_U6058, new_P2_U6059, new_P2_U6060, new_P2_U6061,
    new_P2_U6062, new_P2_U6063, new_P2_U6064, new_P2_U6065, new_P2_U6066,
    new_P2_U6067, new_P2_U6068, new_P2_U6069, new_P2_U6070, new_P2_U6071,
    new_P2_U6072, new_P2_U6073, new_P2_U6074, new_P2_U6075, new_P2_U6076,
    new_P2_U6077, new_P2_U6078, new_P2_U6079, new_P2_U6080, new_P2_U6081,
    new_P2_U6082, new_P2_U6083, new_P2_U6084, new_P2_U6085, new_P2_U6086,
    new_P2_U6087, new_P2_U6088, new_P2_U6089, new_P2_U6090, new_P2_U6091,
    new_P2_U6092, new_P2_U6093, new_P2_U6094, new_P2_U6095, new_P2_U6096,
    new_P2_U6097, new_P2_U6098, new_P2_U6099, new_P2_U6100, new_P2_U6101,
    new_P2_U6102, new_P2_U6103, new_P2_U6104, new_P2_U6105, new_P2_U6106,
    new_P2_U6107, new_P2_U6108, new_P2_U6109, new_P2_U6110, new_P2_U6111,
    new_P2_U6112, new_P2_U6113, new_P2_U6114, new_P2_U6115, new_P2_U6116,
    new_P2_U6117, new_P2_U6118, new_P2_U6119, new_P2_U6120, new_P2_U6121,
    new_P2_U6122, new_P2_U6123, new_P2_U6124, new_P2_U6125, new_P2_U6126,
    new_P2_U6127, new_P2_U6128, new_P2_U6129, new_P2_U6130, new_P2_U6131,
    new_P2_U6132, new_P2_U6133, new_P2_U6134, new_P2_U6135, new_P2_U6136,
    new_P2_U6137, new_P2_U6138, new_P2_U6139, new_P2_U6140, new_P2_U6141,
    new_P2_U6142, new_P2_U6143, new_P2_U6144, new_P2_U6145, new_P2_U6146,
    new_P2_U6147, new_P2_U6148, new_P2_U6149, new_P2_U6150, new_P2_U6151,
    new_P2_U6152, new_P2_U6153, new_P2_U6154, new_P2_U6155, new_P2_U6156,
    new_P2_U6157, new_P2_U6158, new_P2_U6159, new_P2_U6160, new_P2_U6161,
    new_P2_U6162, new_P2_U6163, new_P2_U6164, new_P2_U6165, new_P2_U6166,
    new_P2_U6167, new_P2_U6168, new_P2_U6169, new_P2_U6170, new_P2_U6171,
    new_P2_U6172, new_P2_U6173, new_P2_U6174, new_P2_U6175, new_P2_U6176,
    new_P2_U6177, new_P2_U6178, new_P2_U6179, new_P2_U6180, new_P2_U6181,
    new_P2_U6182, new_P2_U6183, new_P2_U6184, new_P2_U6185, new_P2_U6186,
    new_P2_U6187, new_P2_U6188, new_P2_U6189, new_P2_U6190, new_P2_U6191,
    new_P2_U6192, new_P2_U6193, new_P2_U6194, new_P2_U6195, new_P2_U6196,
    new_P2_U6197, new_P2_U6198, new_P2_U6199, new_P2_U6200, new_P2_U6201,
    new_P2_U6202, new_P2_U6203, new_P2_U6204, new_P2_U6205, new_P2_U6206,
    new_P2_U6207, new_P2_U6208, new_P2_U6209, new_P2_U6210, new_P2_U6211,
    new_P2_U6212, new_P2_U6213, new_P2_U6214, new_P2_U6215, new_P2_U6216,
    new_P2_U6217, new_P2_U6218, new_P2_U6219, new_P2_U6220, new_P2_U6221,
    new_P2_U6222, new_P2_U6223, new_P2_U6224, new_P2_U6225, new_P2_U6226,
    new_P2_U6227, new_P2_U6228, new_P2_U6229, new_P2_U6230, new_P2_U6231,
    new_P2_U6232, new_P2_U6233, new_P2_U6234, new_P2_U6235, new_P2_U6236,
    new_P2_U6237, new_P2_U6238, new_P2_U6239, new_P2_U6240, new_P2_U6241,
    new_P2_U6242, new_P2_U6243, new_P2_U6244, new_P2_U6245, new_P2_U6246,
    new_P2_U6247, new_P2_U6248, new_P2_U6249, new_P2_U6250, new_P2_U6251,
    new_P2_U6252, new_P2_U6253, new_P2_U6254, new_P2_U6255, new_P2_U6256,
    new_P2_U6257, new_P2_U6258, new_P2_U6259, new_P2_U6260, new_P2_U6261,
    new_P2_U6262, new_P2_U6263, new_P2_U6264, new_P2_U6265, new_P2_U6266,
    new_P2_U6267, new_P2_U6268, new_P2_U6269, new_P2_U6270, new_P2_U6271,
    new_P2_U6272, new_P2_U6273, new_P2_U6274, new_P2_U6275, new_P2_U6276,
    new_P2_U6277, new_P2_U6278, new_P2_U6279, new_P2_U6280, new_P2_U6281,
    new_P2_U6282, new_P2_U6283, new_P2_U6284, new_P2_U6285, new_P2_U6286,
    new_P2_U6287, new_P2_U6288, new_P2_U6289, new_P2_U6290, new_P2_U6291,
    new_P2_U6292, new_P2_U6293, new_P2_U6294, new_P2_U6295, new_P2_U6296,
    new_P2_U6297, new_P2_U6298, new_P2_U6299, new_P2_U6300, new_P2_U6301,
    new_P2_U6302, new_P2_U6303, new_P2_U6304, new_P2_U6305, new_P2_U6306,
    new_P2_U6307, new_P2_U6308, new_P2_U6309, new_P2_U6310, new_P2_U6311,
    new_P2_U6312, new_P2_U6313, new_P2_U6314, new_P2_U6315, new_P2_U6316,
    new_P2_U6317, new_P2_U6318, new_P2_U6319, new_P2_U6320, new_P2_U6321,
    new_P2_U6322, new_P2_U6323, new_P2_U6324, new_P2_U6325, new_P2_U6326,
    new_P2_U6327, new_P2_U6328, new_P2_U6329, new_P2_U6330, new_P2_U6331,
    new_P2_U6332, new_P2_U6333, new_P2_U6334, new_P2_U6335, new_P2_U6336,
    new_P2_U6337, new_P2_U6338, new_P2_U6339, new_P2_U6340, new_P2_U6341,
    new_P2_U6342, new_P2_U6343, new_P2_U6344, new_P2_U6345, new_P2_U6346,
    new_P2_U6347, new_P2_U6348, new_P2_U6349, new_P2_U6350, new_P2_U6351,
    new_P2_U6352, new_P2_U6353, new_P2_U6354, new_P2_U6355, new_P2_U6356,
    new_P2_U6357, new_P2_U6358, new_P2_U6359, new_P2_U6360, new_P2_U6361,
    new_P2_U6362, new_P2_U6363, new_P2_U6364, new_P2_U6365, new_P2_U6366,
    new_P2_U6367, new_P2_U6368, new_P2_U6369, new_P2_U6370, new_P2_U6371,
    new_P2_U6372, new_P2_U6373, new_P2_U6374, new_P2_U6375, new_P2_U6376,
    new_P2_U6377, new_P2_U6378, new_P2_U6379, new_P2_U6380, new_P2_U6381,
    new_P2_U6382, new_P2_U6383, new_P2_U6384, new_P2_U6385, new_P2_U6386,
    new_P2_U6387, new_P2_U6388, new_P2_U6389, new_P2_U6390, new_P2_U6391,
    new_P2_U6392, new_P2_U6393, new_P2_U6394, new_P2_U6395, new_P2_U6396,
    new_P2_U6397, new_P2_U6398, new_P2_U6399, new_P2_U6400, new_P2_U6401,
    new_P2_U6402, new_P2_U6403, new_P2_U6404, new_P2_U6405, new_P2_U6406,
    new_P2_U6407, new_P2_U6408, new_P2_U6409, new_P2_U6410, new_P2_U6411,
    new_P2_U6412, new_P2_U6413, new_P2_U6414, new_P2_U6415, new_P2_U6416,
    new_P2_U6417, new_P2_U6418, new_P2_U6419, new_P2_U6420, new_P2_U6421,
    new_P2_U6422, new_P2_U6423, new_P2_U6424, new_P2_U6425, new_P2_U6426,
    new_P2_U6427, new_P2_U6428, new_P2_U6429, new_P2_U6430, new_P2_U6431,
    new_P2_U6432, new_P2_U6433, new_P2_U6434, new_P2_U6435, new_P2_U6436,
    new_P2_U6437, new_P2_U6438, new_P2_U6439, new_P2_U6440, new_P2_U6441,
    new_P2_U6442, new_P2_U6443, new_P2_U6444, new_P2_U6445, new_P2_U6446,
    new_P2_U6447, new_P2_U6448, new_P2_U6449, new_P2_U6450, new_P2_U6451,
    new_P2_U6452, new_P2_U6453, new_P2_U6454, new_P2_U6455, new_P2_U6456,
    new_P2_U6457, new_P2_U6458, new_P2_U6459, new_P2_U6460, new_P2_U6461,
    new_P2_U6462, new_P2_U6463, new_P2_U6464, new_P2_U6465, new_P2_U6466,
    new_P2_U6467, new_P2_U6468, new_P2_U6469, new_P2_U6470, new_P2_U6471,
    new_P2_U6472, new_P2_U6473, new_P2_U6474, new_P2_U6475, new_P2_U6476,
    new_P2_U6477, new_P2_U6478, new_P2_U6479, new_P2_U6480, new_P2_U6481,
    new_P2_U6482, new_P2_U6483, new_P2_U6484, new_P2_U6485, new_P2_U6486,
    new_P2_U6487, new_P2_U6488, new_P2_U6489, new_P2_U6490, new_P2_U6491,
    new_P2_U6492, new_P2_U6493, new_P2_U6494, new_P2_U6495, new_P2_U6496,
    new_P2_U6497, new_P2_U6498, new_P2_U6499, new_P2_U6500, new_P2_U6501,
    new_P2_U6502, new_P2_U6503, new_P2_U6504, new_P2_U6505, new_P2_U6506,
    new_P2_U6507, new_P2_U6508, new_P2_U6509, new_P2_U6510, new_P2_U6511,
    new_P2_U6512, new_P2_U6513, new_P2_U6514, new_P2_U6515, new_P2_U6516,
    new_P2_U6517, new_P2_U6518, new_P2_U6519, new_P2_U6520, new_P2_U6521,
    new_P2_U6522, new_P2_U6523, new_P2_U6524, new_P2_U6525, new_P2_U6526,
    new_P2_U6527, new_P2_U6528, new_P2_U6529, new_P2_U6530, new_P2_U6531,
    new_P2_U6532, new_P2_U6533, new_P2_U6534, new_P2_U6535, new_P2_U6536,
    new_P2_U6537, new_P2_U6538, new_P2_U6539, new_P2_U6540, new_P2_U6541,
    new_P2_U6542, new_P2_U6543, new_P2_U6544, new_P2_U6545, new_P2_U6546,
    new_P2_U6547, new_P2_U6548, new_P2_U6549, new_P2_U6550, new_P2_U6551,
    new_P2_U6552, new_P2_U6553, new_P2_U6554, new_P2_U6555, new_P2_U6556,
    new_P2_U6557, new_P2_U6558, new_P2_U6559, new_P2_U6560, new_P2_U6561,
    new_P2_U6562, new_P2_U6563, new_P2_U6564, new_P2_U6565, new_P2_U6566,
    new_P2_U6567, new_P2_U6568, new_P2_U6569, new_P2_U6570, new_P2_U6571,
    new_P2_U6572, new_P2_U6573, new_P2_U6574, new_P2_U6575, new_P2_U6576,
    new_P2_U6577, new_P2_U6578, new_P2_U6579, new_P2_U6580, new_P2_U6581,
    new_P2_U6582, new_P2_U6583, new_P2_U6584, new_P2_U6585, new_P2_U6586,
    new_P2_U6587, new_P2_U6588, new_P2_U6589, new_P2_U6590, new_P2_U6591,
    new_P2_U6592, new_P2_U6593, new_P2_U6594, new_P2_U6595, new_P2_U6596,
    new_P2_U6597, new_P2_U6598, new_P2_U6599, new_P2_U6600, new_P2_U6601,
    new_P2_U6602, new_P2_U6603, new_P2_U6604, new_P2_U6605, new_P2_U6606,
    new_P2_U6607, new_P2_U6608, new_P2_U6609, new_P2_U6610, new_P2_U6611,
    new_P2_U6612, new_P2_U6613, new_P2_U6614, new_P2_U6615, new_P2_U6616,
    new_P2_U6617, new_P2_U6618, new_P2_U6619, new_P2_U6620, new_P2_U6621,
    new_P2_U6622, new_P2_U6623, new_P2_U6624, new_P2_U6625, new_P2_U6626,
    new_P2_U6627, new_P2_U6628, new_P2_U6629, new_P2_U6630, new_P2_U6631,
    new_P2_U6632, new_P2_U6633, new_P2_U6634, new_P2_U6635, new_P2_U6636,
    new_P2_U6637, new_P2_U6638, new_P2_U6639, new_P2_U6640, new_P2_U6641,
    new_P2_U6642, new_P2_U6643, new_P2_U6644, new_P2_U6645, new_P2_U6646,
    new_P2_U6647, new_P2_U6648, new_P2_U6649, new_P2_U6650, new_P2_U6651,
    new_P2_U6652, new_P2_U6653, new_P2_U6654, new_P2_U6655, new_P2_U6656,
    new_P2_U6657, new_P2_U6658, new_P2_U6659, new_P2_U6660, new_P2_U6661,
    new_P2_U6662, new_P2_U6663, new_P2_U6664, new_P2_U6665, new_P2_U6666,
    new_P2_U6667, new_P2_U6668, new_P2_U6669, new_P2_U6670, new_P2_U6671,
    new_P2_U6672, new_P2_U6673, new_P2_U6674, new_P2_U6675, new_P2_U6676,
    new_P2_U6677, new_P2_U6678, new_P2_U6679, new_P2_U6680, new_P2_U6681,
    new_P2_U6682, new_P2_U6683, new_P2_U6684, new_P2_U6685, new_P2_U6686,
    new_P2_U6687, new_P2_U6688, new_P2_U6689, new_P2_U6690, new_P2_U6691,
    new_P2_U6692, new_P2_U6693, new_P2_U6694, new_P2_U6695, new_P2_U6696,
    new_P2_U6697, new_P2_U6698, new_P2_U6699, new_P2_U6700, new_P2_U6701,
    new_P2_U6702, new_P2_U6703, new_P2_U6704, new_P2_U6705, new_P2_U6706,
    new_P2_U6707, new_P2_U6708, new_P2_U6709, new_P2_U6710, new_P2_U6711,
    new_P2_U6712, new_P2_U6713, new_P2_U6714, new_P2_U6715, new_P2_U6716,
    new_P2_U6717, new_P2_U6718, new_P2_U6719, new_P2_U6720, new_P2_U6721,
    new_P2_U6722, new_P2_U6723, new_P2_U6724, new_P2_U6725, new_P2_U6726,
    new_P2_U6727, new_P2_U6728, new_P2_U6729, new_P2_U6730, new_P2_U6731,
    new_P2_U6732, new_P2_U6733, new_P2_U6734, new_P2_U6735, new_P2_U6736,
    new_P2_U6737, new_P2_U6738, new_P2_U6739, new_P2_U6740, new_P2_U6741,
    new_P2_U6742, new_P2_U6743, new_P2_U6744, new_P2_U6745, new_P2_U6746,
    new_P2_U6747, new_P2_U6748, new_P2_U6749, new_P2_U6750, new_P2_U6751,
    new_P2_U6752, new_P2_U6753, new_P2_U6754, new_P2_U6755, new_P2_U6756,
    new_P2_U6757, new_P2_U6758, new_P2_U6759, new_P2_U6760, new_P2_U6761,
    new_P2_U6762, new_P2_U6763, new_P2_U6764, new_P2_U6765, new_P2_U6766,
    new_P2_U6767, new_P2_U6768, new_P2_U6769, new_P2_U6770, new_P2_U6771,
    new_P2_U6772, new_P2_U6773, new_P2_U6774, new_P2_U6775, new_P2_U6776,
    new_P2_U6777, new_P2_U6778, new_P2_U6779, new_P2_U6780, new_P2_U6781,
    new_P2_U6782, new_P2_U6783, new_P2_U6784, new_P2_U6785, new_P2_U6786,
    new_P2_U6787, new_P2_U6788, new_P2_U6789, new_P2_U6790, new_P2_U6791,
    new_P2_U6792, new_P2_U6793, new_P2_U6794, new_P2_U6795, new_P2_U6796,
    new_P2_U6797, new_P2_U6798, new_P2_U6799, new_P2_U6800, new_P2_U6801,
    new_P2_U6802, new_P2_U6803, new_P2_U6804, new_P2_U6805, new_P2_U6806,
    new_P2_U6807, new_P2_U6808, new_P2_U6809, new_P2_U6810, new_P2_U6811,
    new_P2_U6812, new_P2_U6813, new_P2_U6814, new_P2_U6815, new_P2_U6816,
    new_P2_U6817, new_P2_U6818, new_P2_U6819, new_P2_U6820, new_P2_U6821,
    new_P2_U6822, new_P2_U6823, new_P2_U6824, new_P2_U6825, new_P2_U6826,
    new_P2_U6827, new_P2_U6828, new_P2_U6829, new_P2_U6830, new_P2_U6831,
    new_P2_U6832, new_P2_U6833, new_P2_U6834, new_P2_U6835, new_P2_U6836,
    new_P2_U6837, new_P2_U6838, new_P2_U6839, new_P2_U6840, new_P2_U6841,
    new_P2_U6842, new_P2_U6843, new_P2_U6844, new_P2_U6845, new_P2_U6846,
    new_P2_U6847, new_P2_U6848, new_P2_U6849, new_P2_U6850, new_P2_U6851,
    new_P2_U6852, new_P2_U6853, new_P2_U6854, new_P2_U6855, new_P2_U6856,
    new_P2_U6857, new_P2_U6858, new_P2_U6859, new_P2_U6860, new_P2_U6861,
    new_P2_U6862, new_P2_U6863, new_P2_U6864, new_P2_U6865, new_P2_U6866,
    new_P2_U6867, new_P2_U6868, new_P2_U6869, new_P2_U6870, new_P2_U6871,
    new_P2_U6872, new_P2_U6873, new_P2_U6874, new_P2_U6875, new_P2_U6876,
    new_P2_U6877, new_P2_U6878, new_P2_U6879, new_P2_U6880, new_P2_U6881,
    new_P2_U6882, new_P2_U6883, new_P2_U6884, new_P2_U6885, new_P2_U6886,
    new_P2_U6887, new_P2_U6888, new_P2_U6889, new_P2_U6890, new_P2_U6891,
    new_P2_U6892, new_P2_U6893, new_P2_U6894, new_P2_U6895, new_P2_U6896,
    new_P2_U6897, new_P2_U6898, new_P2_U6899, new_P2_U6900, new_P2_U6901,
    new_P2_U6902, new_P2_U6903, new_P2_U6904, new_P2_U6905, new_P2_U6906,
    new_P2_U6907, new_P2_U6908, new_P2_U6909, new_P2_U6910, new_P2_U6911,
    new_P2_U6912, new_P2_U6913, new_P2_U6914, new_P2_U6915, new_P2_U6916,
    new_P2_U6917, new_P2_U6918, new_P2_U6919, new_P2_U6920, new_P2_U6921,
    new_P2_U6922, new_P2_U6923, new_P2_U6924, new_P2_U6925, new_P2_U6926,
    new_P2_U6927, new_P2_U6928, new_P2_U6929, new_P2_U6930, new_P2_U6931,
    new_P2_U6932, new_P2_U6933, new_P2_U6934, new_P2_U6935, new_P2_U6936,
    new_P2_U6937, new_P2_U6938, new_P2_U6939, new_P2_U6940, new_P2_U6941,
    new_P2_U6942, new_P2_U6943, new_P2_U6944, new_P2_U6945, new_P2_U6946,
    new_P2_U6947, new_P2_U6948, new_P2_U6949, new_P2_U6950, new_P2_U6951,
    new_P2_U6952, new_P2_U6953, new_P2_U6954, new_P2_U6955, new_P2_U6956,
    new_P2_U6957, new_P2_U6958, new_P2_U6959, new_P2_U6960, new_P2_U6961,
    new_P2_U6962, new_P2_U6963, new_P2_U6964, new_P2_U6965, new_P2_U6966,
    new_P2_U6967, new_P2_U6968, new_P2_U6969, new_P2_U6970, new_P2_U6971,
    new_P2_U6972, new_P2_U6973, new_P2_U6974, new_P2_U6975, new_P2_U6976,
    new_P2_U6977, new_P2_U6978, new_P2_U6979, new_P2_U6980, new_P2_U6981,
    new_P2_U6982, new_P2_U6983, new_P2_U6984, new_P2_U6985, new_P2_U6986,
    new_P2_U6987, new_P2_U6988, new_P2_U6989, new_P2_U6990, new_P2_U6991,
    new_P2_U6992, new_P2_U6993, new_P2_U6994, new_P2_U6995, new_P2_U6996,
    new_P2_U6997, new_P2_U6998, new_P2_U6999, new_P2_U7000, new_P2_U7001,
    new_P2_U7002, new_P2_U7003, new_P2_U7004, new_P2_U7005, new_P2_U7006,
    new_P2_U7007, new_P2_U7008, new_P2_U7009, new_P2_U7010, new_P2_U7011,
    new_P2_U7012, new_P2_U7013, new_P2_U7014, new_P2_U7015, new_P2_U7016,
    new_P2_U7017, new_P2_U7018, new_P2_U7019, new_P2_U7020, new_P2_U7021,
    new_P2_U7022, new_P2_U7023, new_P2_U7024, new_P2_U7025, new_P2_U7026,
    new_P2_U7027, new_P2_U7028, new_P2_U7029, new_P2_U7030, new_P2_U7031,
    new_P2_U7032, new_P2_U7033, new_P2_U7034, new_P2_U7035, new_P2_U7036,
    new_P2_U7037, new_P2_U7038, new_P2_U7039, new_P2_U7040, new_P2_U7041,
    new_P2_U7042, new_P2_U7043, new_P2_U7044, new_P2_U7045, new_P2_U7046,
    new_P2_U7047, new_P2_U7048, new_P2_U7049, new_P2_U7050, new_P2_U7051,
    new_P2_U7052, new_P2_U7053, new_P2_U7054, new_P2_U7055, new_P2_U7056,
    new_P2_U7057, new_P2_U7058, new_P2_U7059, new_P2_U7060, new_P2_U7061,
    new_P2_U7062, new_P2_U7063, new_P2_U7064, new_P2_U7065, new_P2_U7066,
    new_P2_U7067, new_P2_U7068, new_P2_U7069, new_P2_U7070, new_P2_U7071,
    new_P2_U7072, new_P2_U7073, new_P2_U7074, new_P2_U7075, new_P2_U7076,
    new_P2_U7077, new_P2_U7078, new_P2_U7079, new_P2_U7080, new_P2_U7081,
    new_P2_U7082, new_P2_U7083, new_P2_U7084, new_P2_U7085, new_P2_U7086,
    new_P2_U7087, new_P2_U7088, new_P2_U7089, new_P2_U7090, new_P2_U7091,
    new_P2_U7092, new_P2_U7093, new_P2_U7094, new_P2_U7095, new_P2_U7096,
    new_P2_U7097, new_P2_U7098, new_P2_U7099, new_P2_U7100, new_P2_U7101,
    new_P2_U7102, new_P2_U7103, new_P2_U7104, new_P2_U7105, new_P2_U7106,
    new_P2_U7107, new_P2_U7108, new_P2_U7109, new_P2_U7110, new_P2_U7111,
    new_P2_U7112, new_P2_U7113, new_P2_U7114, new_P2_U7115, new_P2_U7116,
    new_P2_U7117, new_P2_U7118, new_P2_U7119, new_P2_U7120, new_P2_U7121,
    new_P2_U7122, new_P2_U7123, new_P2_U7124, new_P2_U7125, new_P2_U7126,
    new_P2_U7127, new_P2_U7128, new_P2_U7129, new_P2_U7130, new_P2_U7131,
    new_P2_U7132, new_P2_U7133, new_P2_U7134, new_P2_U7135, new_P2_U7136,
    new_P2_U7137, new_P2_U7138, new_P2_U7139, new_P2_U7140, new_P2_U7141,
    new_P2_U7142, new_P2_U7143, new_P2_U7144, new_P2_U7145, new_P2_U7146,
    new_P2_U7147, new_P2_U7148, new_P2_U7149, new_P2_U7150, new_P2_U7151,
    new_P2_U7152, new_P2_U7153, new_P2_U7154, new_P2_U7155, new_P2_U7156,
    new_P2_U7157, new_P2_U7158, new_P2_U7159, new_P2_U7160, new_P2_U7161,
    new_P2_U7162, new_P2_U7163, new_P2_U7164, new_P2_U7165, new_P2_U7166,
    new_P2_U7167, new_P2_U7168, new_P2_U7169, new_P2_U7170, new_P2_U7171,
    new_P2_U7172, new_P2_U7173, new_P2_U7174, new_P2_U7175, new_P2_U7176,
    new_P2_U7177, new_P2_U7178, new_P2_U7179, new_P2_U7180, new_P2_U7181,
    new_P2_U7182, new_P2_U7183, new_P2_U7184, new_P2_U7185, new_P2_U7186,
    new_P2_U7187, new_P2_U7188, new_P2_U7189, new_P2_U7190, new_P2_U7191,
    new_P2_U7192, new_P2_U7193, new_P2_U7194, new_P2_U7195, new_P2_U7196,
    new_P2_U7197, new_P2_U7198, new_P2_U7199, new_P2_U7200, new_P2_U7201,
    new_P2_U7202, new_P2_U7203, new_P2_U7204, new_P2_U7205, new_P2_U7206,
    new_P2_U7207, new_P2_U7208, new_P2_U7209, new_P2_U7210, new_P2_U7211,
    new_P2_U7212, new_P2_U7213, new_P2_U7214, new_P2_U7215, new_P2_U7216,
    new_P2_U7217, new_P2_U7218, new_P2_U7219, new_P2_U7220, new_P2_U7221,
    new_P2_U7222, new_P2_U7223, new_P2_U7224, new_P2_U7225, new_P2_U7226,
    new_P2_U7227, new_P2_U7228, new_P2_U7229, new_P2_U7230, new_P2_U7231,
    new_P2_U7232, new_P2_U7233, new_P2_U7234, new_P2_U7235, new_P2_U7236,
    new_P2_U7237, new_P2_U7238, new_P2_U7239, new_P2_U7240, new_P2_U7241,
    new_P2_U7242, new_P2_U7243, new_P2_U7244, new_P2_U7245, new_P2_U7246,
    new_P2_U7247, new_P2_U7248, new_P2_U7249, new_P2_U7250, new_P2_U7251,
    new_P2_U7252, new_P2_U7253, new_P2_U7254, new_P2_U7255, new_P2_U7256,
    new_P2_U7257, new_P2_U7258, new_P2_U7259, new_P2_U7260, new_P2_U7261,
    new_P2_U7262, new_P2_U7263, new_P2_U7264, new_P2_U7265, new_P2_U7266,
    new_P2_U7267, new_P2_U7268, new_P2_U7269, new_P2_U7270, new_P2_U7271,
    new_P2_U7272, new_P2_U7273, new_P2_U7274, new_P2_U7275, new_P2_U7276,
    new_P2_U7277, new_P2_U7278, new_P2_U7279, new_P2_U7280, new_P2_U7281,
    new_P2_U7282, new_P2_U7283, new_P2_U7284, new_P2_U7285, new_P2_U7286,
    new_P2_U7287, new_P2_U7288, new_P2_U7289, new_P2_U7290, new_P2_U7291,
    new_P2_U7292, new_P2_U7293, new_P2_U7294, new_P2_U7295, new_P2_U7296,
    new_P2_U7297, new_P2_U7298, new_P2_U7299, new_P2_U7300, new_P2_U7301,
    new_P2_U7302, new_P2_U7303, new_P2_U7304, new_P2_U7305, new_P2_U7306,
    new_P2_U7307, new_P2_U7308, new_P2_U7309, new_P2_U7310, new_P2_U7311,
    new_P2_U7312, new_P2_U7313, new_P2_U7314, new_P2_U7315, new_P2_U7316,
    new_P2_U7317, new_P2_U7318, new_P2_U7319, new_P2_U7320, new_P2_U7321,
    new_P2_U7322, new_P2_U7323, new_P2_U7324, new_P2_U7325, new_P2_U7326,
    new_P2_U7327, new_P2_U7328, new_P2_U7329, new_P2_U7330, new_P2_U7331,
    new_P2_U7332, new_P2_U7333, new_P2_U7334, new_P2_U7335, new_P2_U7336,
    new_P2_U7337, new_P2_U7338, new_P2_U7339, new_P2_U7340, new_P2_U7341,
    new_P2_U7342, new_P2_U7343, new_P2_U7344, new_P2_U7345, new_P2_U7346,
    new_P2_U7347, new_P2_U7348, new_P2_U7349, new_P2_U7350, new_P2_U7351,
    new_P2_U7352, new_P2_U7353, new_P2_U7354, new_P2_U7355, new_P2_U7356,
    new_P2_U7357, new_P2_U7358, new_P2_U7359, new_P2_U7360, new_P2_U7361,
    new_P2_U7362, new_P2_U7363, new_P2_U7364, new_P2_U7365, new_P2_U7366,
    new_P2_U7367, new_P2_U7368, new_P2_U7369, new_P2_U7370, new_P2_U7371,
    new_P2_U7372, new_P2_U7373, new_P2_U7374, new_P2_U7375, new_P2_U7376,
    new_P2_U7377, new_P2_U7378, new_P2_U7379, new_P2_U7380, new_P2_U7381,
    new_P2_U7382, new_P2_U7383, new_P2_U7384, new_P2_U7385, new_P2_U7386,
    new_P2_U7387, new_P2_U7388, new_P2_U7389, new_P2_U7390, new_P2_U7391,
    new_P2_U7392, new_P2_U7393, new_P2_U7394, new_P2_U7395, new_P2_U7396,
    new_P2_U7397, new_P2_U7398, new_P2_U7399, new_P2_U7400, new_P2_U7401,
    new_P2_U7402, new_P2_U7403, new_P2_U7404, new_P2_U7405, new_P2_U7406,
    new_P2_U7407, new_P2_U7408, new_P2_U7409, new_P2_U7410, new_P2_U7411,
    new_P2_U7412, new_P2_U7413, new_P2_U7414, new_P2_U7415, new_P2_U7416,
    new_P2_U7417, new_P2_U7418, new_P2_U7419, new_P2_U7420, new_P2_U7421,
    new_P2_U7422, new_P2_U7423, new_P2_U7424, new_P2_U7425, new_P2_U7426,
    new_P2_U7427, new_P2_U7428, new_P2_U7429, new_P2_U7430, new_P2_U7431,
    new_P2_U7432, new_P2_U7433, new_P2_U7434, new_P2_U7435, new_P2_U7436,
    new_P2_U7437, new_P2_U7438, new_P2_U7439, new_P2_U7440, new_P2_U7441,
    new_P2_U7442, new_P2_U7443, new_P2_U7444, new_P2_U7445, new_P2_U7446,
    new_P2_U7447, new_P2_U7448, new_P2_U7449, new_P2_U7450, new_P2_U7451,
    new_P2_U7452, new_P2_U7453, new_P2_U7454, new_P2_U7455, new_P2_U7456,
    new_P2_U7457, new_P2_U7458, new_P2_U7459, new_P2_U7460, new_P2_U7461,
    new_P2_U7462, new_P2_U7463, new_P2_U7464, new_P2_U7465, new_P2_U7466,
    new_P2_U7467, new_P2_U7468, new_P2_U7469, new_P2_U7470, new_P2_U7471,
    new_P2_U7472, new_P2_U7473, new_P2_U7474, new_P2_U7475, new_P2_U7476,
    new_P2_U7477, new_P2_U7478, new_P2_U7479, new_P2_U7480, new_P2_U7481,
    new_P2_U7482, new_P2_U7483, new_P2_U7484, new_P2_U7485, new_P2_U7486,
    new_P2_U7487, new_P2_U7488, new_P2_U7489, new_P2_U7490, new_P2_U7491,
    new_P2_U7492, new_P2_U7493, new_P2_U7494, new_P2_U7495, new_P2_U7496,
    new_P2_U7497, new_P2_U7498, new_P2_U7499, new_P2_U7500, new_P2_U7501,
    new_P2_U7502, new_P2_U7503, new_P2_U7504, new_P2_U7505, new_P2_U7506,
    new_P2_U7507, new_P2_U7508, new_P2_U7509, new_P2_U7510, new_P2_U7511,
    new_P2_U7512, new_P2_U7513, new_P2_U7514, new_P2_U7515, new_P2_U7516,
    new_P2_U7517, new_P2_U7518, new_P2_U7519, new_P2_U7520, new_P2_U7521,
    new_P2_U7522, new_P2_U7523, new_P2_U7524, new_P2_U7525, new_P2_U7526,
    new_P2_U7527, new_P2_U7528, new_P2_U7529, new_P2_U7530, new_P2_U7531,
    new_P2_U7532, new_P2_U7533, new_P2_U7534, new_P2_U7535, new_P2_U7536,
    new_P2_U7537, new_P2_U7538, new_P2_U7539, new_P2_U7540, new_P2_U7541,
    new_P2_U7542, new_P2_U7543, new_P2_U7544, new_P2_U7545, new_P2_U7546,
    new_P2_U7547, new_P2_U7548, new_P2_U7549, new_P2_U7550, new_P2_U7551,
    new_P2_U7552, new_P2_U7553, new_P2_U7554, new_P2_U7555, new_P2_U7556,
    new_P2_U7557, new_P2_U7558, new_P2_U7559, new_P2_U7560, new_P2_U7561,
    new_P2_U7562, new_P2_U7563, new_P2_U7564, new_P2_U7565, new_P2_U7566,
    new_P2_U7567, new_P2_U7568, new_P2_U7569, new_P2_U7570, new_P2_U7571,
    new_P2_U7572, new_P2_U7573, new_P2_U7574, new_P2_U7575, new_P2_U7576,
    new_P2_U7577, new_P2_U7578, new_P2_U7579, new_P2_U7580, new_P2_U7581,
    new_P2_U7582, new_P2_U7583, new_P2_U7584, new_P2_U7585, new_P2_U7586,
    new_P2_U7587, new_P2_U7588, new_P2_U7589, new_P2_U7590, new_P2_U7591,
    new_P2_U7592, new_P2_U7593, new_P2_U7594, new_P2_U7595, new_P2_U7596,
    new_P2_U7597, new_P2_U7598, new_P2_U7599, new_P2_U7600, new_P2_U7601,
    new_P2_U7602, new_P2_U7603, new_P2_U7604, new_P2_U7605, new_P2_U7606,
    new_P2_U7607, new_P2_U7608, new_P2_U7609, new_P2_U7610, new_P2_U7611,
    new_P2_U7612, new_P2_U7613, new_P2_U7614, new_P2_U7615, new_P2_U7616,
    new_P2_U7617, new_P2_U7618, new_P2_U7619, new_P2_U7620, new_P2_U7621,
    new_P2_U7622, new_P2_U7623, new_P2_U7624, new_P2_U7625, new_P2_U7626,
    new_P2_U7627, new_P2_U7628, new_P2_U7629, new_P2_U7630, new_P2_U7631,
    new_P2_U7632, new_P2_U7633, new_P2_U7634, new_P2_U7635, new_P2_U7636,
    new_P2_U7637, new_P2_U7638, new_P2_U7639, new_P2_U7640, new_P2_U7641,
    new_P2_U7642, new_P2_U7643, new_P2_U7644, new_P2_U7645, new_P2_U7646,
    new_P2_U7647, new_P2_U7648, new_P2_U7649, new_P2_U7650, new_P2_U7651,
    new_P2_U7652, new_P2_U7653, new_P2_U7654, new_P2_U7655, new_P2_U7656,
    new_P2_U7657, new_P2_U7658, new_P2_U7659, new_P2_U7660, new_P2_U7661,
    new_P2_U7662, new_P2_U7663, new_P2_U7664, new_P2_U7665, new_P2_U7666,
    new_P2_U7667, new_P2_U7668, new_P2_U7669, new_P2_U7670, new_P2_U7671,
    new_P2_U7672, new_P2_U7673, new_P2_U7674, new_P2_U7675, new_P2_U7676,
    new_P2_U7677, new_P2_U7678, new_P2_U7679, new_P2_U7680, new_P2_U7681,
    new_P2_U7682, new_P2_U7683, new_P2_U7684, new_P2_U7685, new_P2_U7686,
    new_P2_U7687, new_P2_U7688, new_P2_U7689, new_P2_U7690, new_P2_U7691,
    new_P2_U7692, new_P2_U7693, new_P2_U7694, new_P2_U7695, new_P2_U7696,
    new_P2_U7697, new_P2_U7698, new_P2_U7699, new_P2_U7700, new_P2_U7701,
    new_P2_U7702, new_P2_U7703, new_P2_U7704, new_P2_U7705, new_P2_U7706,
    new_P2_U7707, new_P2_U7708, new_P2_U7709, new_P2_U7710, new_P2_U7711,
    new_P2_U7712, new_P2_U7713, new_P2_U7714, new_P2_U7715, new_P2_U7716,
    new_P2_U7717, new_P2_U7718, new_P2_U7719, new_P2_U7720, new_P2_U7721,
    new_P2_U7722, new_P2_U7723, new_P2_U7724, new_P2_U7725, new_P2_U7726,
    new_P2_U7727, new_P2_U7728, new_P2_U7729, new_P2_U7730, new_P2_U7731,
    new_P2_U7732, new_P2_U7733, new_P2_U7734, new_P2_U7735, new_P2_U7736,
    new_P2_U7737, new_P2_U7738, new_P2_U7739, new_P2_U7740, new_P2_U7741,
    new_P2_U7742, new_P2_U7743, new_P2_U7744, new_P2_U7745, new_P2_U7746,
    new_P2_U7747, new_P2_U7748, new_P2_U7749, new_P2_U7750, new_P2_U7751,
    new_P2_U7752, new_P2_U7753, new_P2_U7754, new_P2_U7755, new_P2_U7756,
    new_P2_U7757, new_P2_U7758, new_P2_U7759, new_P2_U7760, new_P2_U7761,
    new_P2_U7762, new_P2_U7763, new_P2_U7764, new_P2_U7765, new_P2_U7766,
    new_P2_U7767, new_P2_U7768, new_P2_U7769, new_P2_U7770, new_P2_U7771,
    new_P2_U7772, new_P2_U7773, new_P2_U7774, new_P2_U7775, new_P2_U7776,
    new_P2_U7777, new_P2_U7778, new_P2_U7779, new_P2_U7780, new_P2_U7781,
    new_P2_U7782, new_P2_U7783, new_P2_U7784, new_P2_U7785, new_P2_U7786,
    new_P2_U7787, new_P2_U7788, new_P2_U7789, new_P2_U7790, new_P2_U7791,
    new_P2_U7792, new_P2_U7793, new_P2_U7794, new_P2_U7795, new_P2_U7796,
    new_P2_U7797, new_P2_U7798, new_P2_U7799, new_P2_U7800, new_P2_U7801,
    new_P2_U7802, new_P2_U7803, new_P2_U7804, new_P2_U7805, new_P2_U7806,
    new_P2_U7807, new_P2_U7808, new_P2_U7809, new_P2_U7810, new_P2_U7811,
    new_P2_U7812, new_P2_U7813, new_P2_U7814, new_P2_U7815, new_P2_U7816,
    new_P2_U7817, new_P2_U7818, new_P2_U7819, new_P2_U7820, new_P2_U7821,
    new_P2_U7822, new_P2_U7823, new_P2_U7824, new_P2_U7825, new_P2_U7826,
    new_P2_U7827, new_P2_U7828, new_P2_U7829, new_P2_U7830, new_P2_U7831,
    new_P2_U7832, new_P2_U7833, new_P2_U7834, new_P2_U7835, new_P2_U7836,
    new_P2_U7837, new_P2_U7838, new_P2_U7839, new_P2_U7840, new_P2_U7841,
    new_P2_U7842, new_P2_U7843, new_P2_U7844, new_P2_U7845, new_P2_U7846,
    new_P2_U7847, new_P2_U7848, new_P2_U7849, new_P2_U7850, new_P2_U7851,
    new_P2_U7852, new_P2_U7853, new_P2_U7854, new_P2_U7855, new_P2_U7856,
    new_P2_U7857, new_P2_U7858, new_P2_U7859, new_P2_U7860, new_P2_U7861,
    new_P2_U7862, new_P2_U7863, new_P2_U7864, new_P2_U7865, new_P2_U7866,
    new_P2_U7867, new_P2_U7868, new_P2_U7869, new_P2_U7870, new_P2_U7871,
    new_P2_U7872, new_P2_U7873, new_P2_U7874, new_P2_U7875, new_P2_U7876,
    new_P2_U7877, new_P2_U7878, new_P2_U7879, new_P2_U7880, new_P2_U7881,
    new_P2_U7882, new_P2_U7883, new_P2_U7884, new_P2_U7885, new_P2_U7886,
    new_P2_U7887, new_P2_U7888, new_P2_U7889, new_P2_U7890, new_P2_U7891,
    new_P2_U7892, new_P2_U7893, new_P2_U7894, new_P2_U7895, new_P2_U7896,
    new_P2_U7897, new_P2_U7898, new_P2_U7899, new_P2_U7900, new_P2_U7901,
    new_P2_U7902, new_P2_U7903, new_P2_U7904, new_P2_U7905, new_P2_U7906,
    new_P2_U7907, new_P2_U7908, new_P2_U7909, new_P2_U7910, new_P2_U7911,
    new_P2_U7912, new_P2_U7913, new_P2_U7914, new_P2_U7915, new_P2_U7916,
    new_P2_U7917, new_P2_U7918, new_P2_U7919, new_P2_U7920, new_P2_U7921,
    new_P2_U7922, new_P2_U7923, new_P2_U7924, new_P2_U7925, new_P2_U7926,
    new_P2_U7927, new_P2_U7928, new_P2_U7929, new_P2_U7930, new_P2_U7931,
    new_P2_U7932, new_P2_U7933, new_P2_U7934, new_P2_U7935, new_P2_U7936,
    new_P2_U7937, new_P2_U7938, new_P2_U7939, new_P2_U7940, new_P2_U7941,
    new_P2_U7942, new_P2_U7943, new_P2_U7944, new_P2_U7945, new_P2_U7946,
    new_P2_U7947, new_P2_U7948, new_P2_U7949, new_P2_U7950, new_P2_U7951,
    new_P2_U7952, new_P2_U7953, new_P2_U7954, new_P2_U7955, new_P2_U7956,
    new_P2_U7957, new_P2_U7958, new_P2_U7959, new_P2_U7960, new_P2_U7961,
    new_P2_U7962, new_P2_U7963, new_P2_U7964, new_P2_U7965, new_P2_U7966,
    new_P2_U7967, new_P2_U7968, new_P2_U7969, new_P2_U7970, new_P2_U7971,
    new_P2_U7972, new_P2_U7973, new_P2_U7974, new_P2_U7975, new_P2_U7976,
    new_P2_U7977, new_P2_U7978, new_P2_U7979, new_P2_U7980, new_P2_U7981,
    new_P2_U7982, new_P2_U7983, new_P2_U7984, new_P2_U7985, new_P2_U7986,
    new_P2_U7987, new_P2_U7988, new_P2_U7989, new_P2_U7990, new_P2_U7991,
    new_P2_U7992, new_P2_U7993, new_P2_U7994, new_P2_U7995, new_P2_U7996,
    new_P2_U7997, new_P2_U7998, new_P2_U7999, new_P2_U8000, new_P2_U8001,
    new_P2_U8002, new_P2_U8003, new_P2_U8004, new_P2_U8005, new_P2_U8006,
    new_P2_U8007, new_P2_U8008, new_P2_U8009, new_P2_U8010, new_P2_U8011,
    new_P2_U8012, new_P2_U8013, new_P2_U8014, new_P2_U8015, new_P2_U8016,
    new_P2_U8017, new_P2_U8018, new_P2_U8019, new_P2_U8020, new_P2_U8021,
    new_P2_U8022, new_P2_U8023, new_P2_U8024, new_P2_U8025, new_P2_U8026,
    new_P2_U8027, new_P2_U8028, new_P2_U8029, new_P2_U8030, new_P2_U8031,
    new_P2_U8032, new_P2_U8033, new_P2_U8034, new_P2_U8035, new_P2_U8036,
    new_P2_U8037, new_P2_U8038, new_P2_U8039, new_P2_U8040, new_P2_U8041,
    new_P2_U8042, new_P2_U8043, new_P2_U8044, new_P2_U8045, new_P2_U8046,
    new_P2_U8047, new_P2_U8048, new_P2_U8049, new_P2_U8050, new_P2_U8051,
    new_P2_U8052, new_P2_U8053, new_P2_U8054, new_P2_U8055, new_P2_U8056,
    new_P2_U8057, new_P2_U8058, new_P2_U8059, new_P2_U8060, new_P2_U8061,
    new_P2_U8062, new_P2_U8063, new_P2_U8064, new_P2_U8065, new_P2_U8066,
    new_P2_U8067, new_P2_U8068, new_P2_U8069, new_P2_U8070, new_P2_U8071,
    new_P2_U8072, new_P2_U8073, new_P2_U8074, new_P2_U8075, new_P2_U8076,
    new_P2_U8077, new_P2_U8078, new_P2_U8079, new_P2_U8080, new_P2_U8081,
    new_P2_U8082, new_P2_U8083, new_P2_U8084, new_P2_U8085, new_P2_U8086,
    new_P2_U8087, new_P2_U8088, new_P2_U8089, new_P2_U8090, new_P2_U8091,
    new_P2_U8092, new_P2_U8093, new_P2_U8094, new_P2_U8095, new_P2_U8096,
    new_P2_U8097, new_P2_U8098, new_P2_U8099, new_P2_U8100, new_P2_U8101,
    new_P2_U8102, new_P2_U8103, new_P2_U8104, new_P2_U8105, new_P2_U8106,
    new_P2_U8107, new_P2_U8108, new_P2_U8109, new_P2_U8110, new_P2_U8111,
    new_P2_U8112, new_P2_U8113, new_P2_U8114, new_P2_U8115, new_P2_U8116,
    new_P2_U8117, new_P2_U8118, new_P2_U8119, new_P2_U8120, new_P2_U8121,
    new_P2_U8122, new_P2_U8123, new_P2_U8124, new_P2_U8125, new_P2_U8126,
    new_P2_U8127, new_P2_U8128, new_P2_U8129, new_P2_U8130, new_P2_U8131,
    new_P2_U8132, new_P2_U8133, new_P2_U8134, new_P2_U8135, new_P2_U8136,
    new_P2_U8137, new_P2_U8138, new_P2_U8139, new_P2_U8140, new_P2_U8141,
    new_P2_U8142, new_P2_U8143, new_P2_U8144, new_P2_U8145, new_P2_U8146,
    new_P2_U8147, new_P2_U8148, new_P2_U8149, new_P2_U8150, new_P2_U8151,
    new_P2_U8152, new_P2_U8153, new_P2_U8154, new_P2_U8155, new_P2_U8156,
    new_P2_U8157, new_P2_U8158, new_P2_U8159, new_P2_U8160, new_P2_U8161,
    new_P2_U8162, new_P2_U8163, new_P2_U8164, new_P2_U8165, new_P2_U8166,
    new_P2_U8167, new_P2_U8168, new_P2_U8169, new_P2_U8170, new_P2_U8171,
    new_P2_U8172, new_P2_U8173, new_P2_U8174, new_P2_U8175, new_P2_U8176,
    new_P2_U8177, new_P2_U8178, new_P2_U8179, new_P2_U8180, new_P2_U8181,
    new_P2_U8182, new_P2_U8183, new_P2_U8184, new_P2_U8185, new_P2_U8186,
    new_P2_U8187, new_P2_U8188, new_P2_U8189, new_P2_U8190, new_P2_U8191,
    new_P2_U8192, new_P2_U8193, new_P2_U8194, new_P2_U8195, new_P2_U8196,
    new_P2_U8197, new_P2_U8198, new_P2_U8199, new_P2_U8200, new_P2_U8201,
    new_P2_U8202, new_P2_U8203, new_P2_U8204, new_P2_U8205, new_P2_U8206,
    new_P2_U8207, new_P2_U8208, new_P2_U8209, new_P2_U8210, new_P2_U8211,
    new_P2_U8212, new_P2_U8213, new_P2_U8214, new_P2_U8215, new_P2_U8216,
    new_P2_U8217, new_P2_U8218, new_P2_U8219, new_P2_U8220, new_P2_U8221,
    new_P2_U8222, new_P2_U8223, new_P2_U8224, new_P2_U8225, new_P2_U8226,
    new_P2_U8227, new_P2_U8228, new_P2_U8229, new_P2_U8230, new_P2_U8231,
    new_P2_U8232, new_P2_U8233, new_P2_U8234, new_P2_U8235, new_P2_U8236,
    new_P2_U8237, new_P2_U8238, new_P2_U8239, new_P2_U8240, new_P2_U8241,
    new_P2_U8242, new_P2_U8243, new_P2_U8244, new_P2_U8245, new_P2_U8246,
    new_P2_U8247, new_P2_U8248, new_P2_U8249, new_P2_U8250, new_P2_U8251,
    new_P2_U8252, new_P2_U8253, new_P2_U8254, new_P2_U8255, new_P2_U8256,
    new_P2_U8257, new_P2_U8258, new_P2_U8259, new_P2_U8260, new_P2_U8261,
    new_P2_U8262, new_P2_U8263, new_P2_U8264, new_P2_U8265, new_P2_U8266,
    new_P2_U8267, new_P2_U8268, new_P2_U8269, new_P2_U8270, new_P2_U8271,
    new_P2_U8272, new_P2_U8273, new_P2_U8274, new_P2_U8275, new_P2_U8276,
    new_P2_U8277, new_P2_U8278, new_P2_U8279, new_P2_U8280, new_P2_U8281,
    new_P2_U8282, new_P2_U8283, new_P2_U8284, new_P2_U8285, new_P2_U8286,
    new_P2_U8287, new_P2_U8288, new_P2_U8289, new_P2_U8290, new_P2_U8291,
    new_P2_U8292, new_P2_U8293, new_P2_U8294, new_P2_U8295, new_P2_U8296,
    new_P2_U8297, new_P2_U8298, new_P2_U8299, new_P2_U8300, new_P2_U8301,
    new_P2_U8302, new_P2_U8303, new_P2_U8304, new_P2_U8305, new_P2_U8306,
    new_P2_U8307, new_P2_U8308, new_P2_U8309, new_P2_U8310, new_P2_U8311,
    new_P2_U8312, new_P2_U8313, new_P2_U8314, new_P2_U8315, new_P2_U8316,
    new_P2_U8317, new_P2_U8318, new_P2_U8319, new_P2_U8320, new_P2_U8321,
    new_P2_U8322, new_P2_U8323, new_P2_U8324, new_P2_U8325, new_P2_U8326,
    new_P2_U8327, new_P2_U8328, new_P2_U8329, new_P2_U8330, new_P2_U8331,
    new_P2_U8332, new_P2_U8333, new_P2_U8334, new_P2_U8335, new_P2_U8336,
    new_P2_U8337, new_P2_U8338, new_P2_U8339, new_P2_U8340, new_P2_U8341,
    new_P2_U8342, new_P2_U8343, new_P2_U8344, new_P2_U8345, new_P2_U8346,
    new_P2_U8347, new_P2_U8348, new_P2_U8349, new_P2_U8350, new_P2_U8351,
    new_P2_U8352, new_P2_U8353, new_P2_U8354, new_P2_U8355, new_P2_U8356,
    new_P2_U8357, new_P2_U8358, new_P2_U8359, new_P2_U8360, new_P2_U8361,
    new_P2_U8362, new_P2_U8363, new_P2_U8364, new_P2_U8365, new_P2_U8366,
    new_P2_U8367, new_P2_U8368, new_P2_U8369, new_P2_U8370, new_P2_U8371,
    new_P2_U8372, new_P2_U8373, new_P2_U8374, new_P2_U8375, new_P2_U8376,
    new_P2_U8377, new_P2_U8378, new_P2_U8379, new_P2_U8380, new_P2_U8381,
    new_P2_U8382, new_P2_U8383, new_P2_U8384, new_P2_U8385, new_P2_U8386,
    new_P2_U8387, new_P2_U8388, new_P2_U8389, new_P2_U8390, new_P2_U8391,
    new_P2_U8392, new_P2_U8393, new_P2_U8394, new_P2_U8395, new_P2_U8396,
    new_P2_U8397, new_P2_U8398, new_P2_U8399, new_P2_U8400, new_P2_U8401,
    new_P2_U8402, new_P2_U8403, new_P2_U8404, new_P2_U8405, new_P2_U8406,
    new_P2_U8407, new_P2_U8408, new_P2_U8409, new_P2_U8410, new_P2_U8411,
    new_P2_U8412, new_P2_U8413, new_P2_U8414, new_P2_U8415, new_P2_U8416,
    new_P2_U8417, new_P2_U8418, new_P2_U8419, new_P2_U8420, new_P2_U8421,
    new_P2_U8422, new_P2_U8423, new_P2_U8424, new_P2_U8425, new_P2_U8426,
    new_P2_U8427, new_P2_U8428, new_P2_U8429, new_P2_U8430, new_P2_U8431,
    new_P2_U8432, new_P2_U8433, new_P2_U8434, new_P1_ADD_405_U171,
    new_P1_ADD_405_U170, new_P1_ADD_405_U169, new_P1_ADD_405_U168,
    new_P1_ADD_405_U167, new_P1_ADD_405_U166, new_P1_ADD_405_U165,
    new_P1_ADD_405_U164, new_P1_ADD_405_U163, new_P1_ADD_405_U162,
    new_P1_ADD_405_U161, new_P1_ADD_405_U160, new_P1_ADD_405_U159,
    new_P1_ADD_405_U158, new_P1_ADD_405_U157, new_P1_ADD_405_U156,
    new_P1_ADD_405_U155, new_P1_ADD_405_U154, new_P1_ADD_405_U153,
    new_P1_ADD_405_U152, new_P1_ADD_405_U151, new_P1_ADD_405_U150,
    new_P1_ADD_405_U149, new_P1_ADD_405_U148, new_P1_ADD_405_U147,
    new_P1_ADD_405_U146, new_P1_ADD_405_U145, new_P1_ADD_405_U144,
    new_P1_ADD_405_U143, new_P1_ADD_405_U142, new_P1_ADD_405_U141,
    new_P1_ADD_405_U140, new_P1_ADD_405_U139, new_P1_ADD_405_U138,
    new_P1_ADD_405_U137, new_P1_ADD_405_U136, new_P1_ADD_405_U135,
    new_P1_ADD_405_U134, new_P1_ADD_405_U133, new_P1_ADD_405_U132,
    new_P1_ADD_405_U131, new_P1_ADD_405_U130, new_P1_ADD_405_U129,
    new_P1_ADD_405_U128, new_P1_ADD_405_U127, new_P1_ADD_405_U126,
    new_P1_ADD_405_U125, new_P1_ADD_405_U124, new_P1_ADD_405_U123,
    new_P1_ADD_405_U122, new_P1_ADD_405_U121, new_P1_ADD_405_U120,
    new_P1_ADD_405_U119, new_P1_ADD_405_U118, new_P1_ADD_405_U117,
    new_P1_ADD_405_U116, new_P1_ADD_405_U115, new_P1_U2352, new_P1_U2353,
    new_P1_U2354, new_P1_U2355, new_P1_U2356, new_P1_U2357, new_P1_U2358,
    new_P1_U2359, new_P1_U2360, new_P1_U2361, new_P1_U2362, new_P1_U2363,
    new_P1_U2364, new_P1_U2365, new_P1_U2366, new_P1_U2367, new_P1_U2368,
    new_P1_U2369, new_P1_U2370, new_P1_U2371, new_P1_U2372, new_P1_U2373,
    new_P1_U2374, new_P1_U2375, new_P1_U2376, new_P1_U2377, new_P1_U2378,
    new_P1_U2379, new_P1_U2380, new_P1_U2381, new_P1_U2382, new_P1_U2383,
    new_P1_U2384, new_P1_U2385, new_P1_U2386, new_P1_U2387, new_P1_U2388,
    new_P1_U2389, new_P1_U2390, new_P1_U2391, new_P1_U2392, new_P1_U2393,
    new_P1_U2394, new_P1_U2395, new_P1_U2396, new_P1_U2397, new_P1_U2398,
    new_P1_U2399, new_P1_U2400, new_P1_U2401, new_P1_U2402, new_P1_U2403,
    new_P1_U2404, new_P1_U2405, new_P1_U2406, new_P1_U2407, new_P1_U2408,
    new_P1_U2409, new_P1_U2410, new_P1_U2411, new_P1_U2412, new_P1_U2413,
    new_P1_U2414, new_P1_U2415, new_P1_U2416, new_P1_U2417, new_P1_U2418,
    new_P1_U2419, new_P1_U2420, new_P1_U2421, new_P1_U2422, new_P1_U2423,
    new_P1_U2424, new_P1_U2425, new_P1_U2426, new_P1_U2427, new_P1_U2428,
    new_P1_U2429, new_P1_U2430, new_P1_U2431, new_P1_U2432, new_P1_U2433,
    new_P1_U2434, new_P1_U2435, new_P1_U2436, new_P1_U2437, new_P1_U2438,
    new_P1_U2439, new_P1_U2440, new_P1_U2441, new_P1_U2442, new_P1_U2443,
    new_P1_U2444, new_P1_U2445, new_P1_U2446, new_P1_U2447, new_P1_U2448,
    new_P1_U2449, new_P1_U2450, new_P1_U2451, new_P1_U2452, new_P1_U2453,
    new_P1_U2454, new_P1_U2455, new_P1_U2456, new_P1_U2457, new_P1_U2458,
    new_P1_U2459, new_P1_U2460, new_P1_U2461, new_P1_U2462, new_P1_U2463,
    new_P1_U2464, new_P1_U2465, new_P1_U2466, new_P1_U2467, new_P1_U2468,
    new_P1_U2469, new_P1_U2470, new_P1_U2471, new_P1_U2472, new_P1_U2473,
    new_P1_U2474, new_P1_U2475, new_P1_U2476, new_P1_U2477, new_P1_U2478,
    new_P1_U2479, new_P1_U2480, new_P1_U2481, new_P1_U2482, new_P1_U2483,
    new_P1_U2484, new_P1_U2485, new_P1_U2486, new_P1_U2487, new_P1_U2488,
    new_P1_U2489, new_P1_U2490, new_P1_U2491, new_P1_U2492, new_P1_U2493,
    new_P1_U2494, new_P1_U2495, new_P1_U2496, new_P1_U2497, new_P1_U2498,
    new_P1_U2499, new_P1_U2500, new_P1_U2501, new_P1_U2502, new_P1_U2503,
    new_P1_U2504, new_P1_U2505, new_P1_U2506, new_P1_U2507, new_P1_U2508,
    new_P1_U2509, new_P1_U2510, new_P1_U2511, new_P1_U2512, new_P1_U2513,
    new_P1_U2514, new_P1_U2515, new_P1_U2516, new_P1_U2517, new_P1_U2518,
    new_P1_U2519, new_P1_U2520, new_P1_U2521, new_P1_U2522, new_P1_U2523,
    new_P1_U2524, new_P1_U2525, new_P1_U2526, new_P1_U2527, new_P1_U2528,
    new_P1_U2529, new_P1_U2530, new_P1_U2531, new_P1_U2532, new_P1_U2533,
    new_P1_U2534, new_P1_U2535, new_P1_U2536, new_P1_U2537, new_P1_U2538,
    new_P1_U2539, new_P1_U2540, new_P1_U2541, new_P1_U2542, new_P1_U2543,
    new_P1_U2544, new_P1_U2545, new_P1_U2546, new_P1_U2547, new_P1_U2548,
    new_P1_U2549, new_P1_U2550, new_P1_U2551, new_P1_U2552, new_P1_U2553,
    new_P1_U2554, new_P1_U2555, new_P1_U2556, new_P1_U2557, new_P1_U2558,
    new_P1_U2559, new_P1_U2560, new_P1_U2561, new_P1_U2562, new_P1_U2563,
    new_P1_U2564, new_P1_U2565, new_P1_U2566, new_P1_U2567, new_P1_U2568,
    new_P1_U2569, new_P1_U2570, new_P1_U2571, new_P1_U2572, new_P1_U2573,
    new_P1_U2574, new_P1_U2575, new_P1_U2576, new_P1_U2577, new_P1_U2578,
    new_P1_U2579, new_P1_U2580, new_P1_U2581, new_P1_U2582, new_P1_U2583,
    new_P1_U2584, new_P1_U2585, new_P1_U2586, new_P1_U2587, new_P1_U2588,
    new_P1_U2589, new_P1_U2590, new_P1_U2591, new_P1_U2592, new_P1_U2593,
    new_P1_U2594, new_P1_U2595, new_P1_U2596, new_P1_U2597, new_P1_U2598,
    new_P1_U2599, new_P1_U2600, new_P1_U2601, new_P1_U2602, new_P1_U2603,
    new_P1_U2604, new_P1_U2605, new_P1_U2606, new_P1_U2607, new_P1_U2608,
    new_P1_U2609, new_P1_U2610, new_P1_U2611, new_P1_U2612, new_P1_U2613,
    new_P1_U2614, new_P1_U2615, new_P1_U2616, new_P1_U2617, new_P1_U2618,
    new_P1_ADD_405_U114, new_P1_U2620, new_P1_U2621, new_P1_U2622,
    new_P1_U2623, new_P1_U2624, new_P1_U2625, new_P1_U2626, new_P1_U2627,
    new_P1_U2628, new_P1_U2629, new_P1_U2630, new_P1_U2631, new_P1_U2632,
    new_P1_U2633, new_P1_U2634, new_P1_U2635, new_P1_U2636, new_P1_U2637,
    new_P1_U2638, new_P1_U2639, new_P1_U2640, new_P1_U2641, new_P1_U2642,
    new_P1_U2643, new_P1_U2644, new_P1_U2645, new_P1_U2646, new_P1_U2647,
    new_P1_U2648, new_P1_U2649, new_P1_U2650, new_P1_U2651, new_P1_U2652,
    new_P1_U2653, new_P1_U2654, new_P1_U2655, new_P1_U2656, new_P1_U2657,
    new_P1_U2658, new_P1_U2659, new_P1_U2660, new_P1_U2661, new_P1_U2662,
    new_P1_U2663, new_P1_U2664, new_P1_U2665, new_P1_U2666, new_P1_U2667,
    new_P1_U2668, new_P1_U2669, new_P1_U2670, new_P1_U2671, new_P1_U2672,
    new_P1_U2673, new_P1_U2674, new_P1_U2675, new_P1_U2676, new_P1_U2677,
    new_P1_U2678, new_P1_U2679, new_P1_U2680, new_P1_U2681, new_P1_U2682,
    new_P1_U2683, new_P1_U2684, new_P1_U2685, new_P1_U2686, new_P1_U2687,
    new_P1_U2688, new_P1_U2689, new_P1_U2690, new_P1_U2691, new_P1_U2692,
    new_P1_U2693, new_P1_U2694, new_P1_U2695, new_P1_U2696, new_P1_U2697,
    new_P1_U2698, new_P1_U2699, new_P1_U2700, new_P1_U2701, new_P1_U2702,
    new_P1_U2703, new_P1_U2704, new_P1_U2705, new_P1_U2706, new_P1_U2707,
    new_P1_U2708, new_P1_U2709, new_P1_U2710, new_P1_U2711, new_P1_U2712,
    new_P1_U2713, new_P1_U2714, new_P1_U2715, new_P1_U2716, new_P1_U2717,
    new_P1_U2718, new_P1_U2719, new_P1_U2720, new_P1_U2721, new_P1_U2722,
    new_P1_U2723, new_P1_U2724, new_P1_U2725, new_P1_U2726, new_P1_U2727,
    new_P1_U2728, new_P1_U2729, new_P1_U2730, new_P1_U2731, new_P1_U2732,
    new_P1_U2733, new_P1_U2734, new_P1_U2735, new_P1_U2736, new_P1_U2737,
    new_P1_U2738, new_P1_U2739, new_P1_U2740, new_P1_U2741, new_P1_U2742,
    new_P1_U2743, new_P1_U2744, new_P1_U2745, new_P1_U2746, new_P1_U2747,
    new_P1_U2748, new_P1_U2749, new_P1_U2750, new_P1_U2751, new_P1_U2752,
    new_P1_U2753, new_P1_U2754, new_P1_U2755, new_P1_U2756, new_P1_U2757,
    new_P1_U2758, new_P1_U2759, new_P1_U2760, new_P1_U2761, new_P1_U2762,
    new_P1_U2763, new_P1_U2764, new_P1_U2765, new_P1_U2766, new_P1_U2767,
    new_P1_U2768, new_P1_U2769, new_P1_U2770, new_P1_U2771, new_P1_U2772,
    new_P1_U2773, new_P1_U2774, new_P1_U2775, new_P1_U2776, new_P1_U2777,
    new_P1_U2778, new_P1_U2779, new_P1_U2780, new_P1_U2781, new_P1_U2782,
    new_P1_U2783, new_P1_U2784, new_P1_U2785, new_P1_U2786, new_P1_U2787,
    new_P1_U2788, new_P1_U2789, new_P1_U2790, new_P1_U2791, new_P1_U2792,
    new_P1_U2793, new_P1_U2794, new_P1_U2795, new_P1_U2796, new_P1_U2797,
    new_P1_U2798, new_P1_U2799, new_P1_U2800, new_P1_U3227, new_P1_U3228,
    new_P1_U3229, new_P1_U3230, new_P1_U3231, new_P1_U3232, new_P1_U3233,
    new_P1_U3234, new_P1_U3235, new_P1_U3236, new_P1_U3237, new_P1_U3238,
    new_P1_U3239, new_P1_U3240, new_P1_U3241, new_P1_U3242, new_P1_U3243,
    new_P1_U3244, new_P1_U3245, new_P1_U3246, new_P1_U3247, new_P1_U3248,
    new_P1_U3249, new_P1_U3250, new_P1_U3251, new_P1_U3252, new_P1_U3253,
    new_P1_U3254, new_P1_U3255, new_P1_U3256, new_P1_U3257, new_P1_U3258,
    new_P1_U3259, new_P1_U3260, new_P1_U3261, new_P1_U3262, new_P1_U3263,
    new_P1_U3264, new_P1_U3265, new_P1_U3266, new_P1_U3267, new_P1_U3268,
    new_P1_U3269, new_P1_U3270, new_P1_U3271, new_P1_U3272, new_P1_U3273,
    new_P1_U3274, new_P1_U3275, new_P1_U3276, new_P1_U3277, new_P1_U3278,
    new_P1_U3279, new_P1_U3280, new_P1_U3281, new_P1_U3282, new_P1_U3283,
    new_P1_U3284, new_P1_U3285, new_P1_U3286, new_P1_U3287, new_P1_U3288,
    new_P1_U3289, new_P1_U3290, new_P1_U3291, new_P1_U3292, new_P1_U3293,
    new_P1_U3294, new_P1_U3295, new_P1_U3296, new_P1_U3297, new_P1_U3298,
    new_P1_U3299, new_P1_U3300, new_P1_U3301, new_P1_U3302, new_P1_U3303,
    new_P1_U3304, new_P1_U3305, new_P1_U3306, new_P1_U3307, new_P1_U3308,
    new_P1_U3309, new_P1_U3310, new_P1_U3311, new_P1_U3312, new_P1_U3313,
    new_P1_U3314, new_P1_U3315, new_P1_U3316, new_P1_U3317, new_P1_U3318,
    new_P1_U3319, new_P1_U3320, new_P1_U3321, new_P1_U3322, new_P1_U3323,
    new_P1_U3324, new_P1_U3325, new_P1_U3326, new_P1_U3327, new_P1_U3328,
    new_P1_U3329, new_P1_U3330, new_P1_U3331, new_P1_U3332, new_P1_U3333,
    new_P1_U3334, new_P1_U3335, new_P1_U3336, new_P1_U3337, new_P1_U3338,
    new_P1_U3339, new_P1_U3340, new_P1_U3341, new_P1_U3342, new_P1_U3343,
    new_P1_U3344, new_P1_U3345, new_P1_U3346, new_P1_U3347, new_P1_U3348,
    new_P1_U3349, new_P1_U3350, new_P1_U3351, new_P1_U3352, new_P1_U3353,
    new_P1_U3354, new_P1_U3355, new_P1_U3356, new_P1_U3357, new_P1_U3358,
    new_P1_U3359, new_P1_U3360, new_P1_U3361, new_P1_U3362, new_P1_U3363,
    new_P1_U3364, new_P1_U3365, new_P1_U3366, new_P1_U3367, new_P1_U3368,
    new_P1_U3369, new_P1_U3370, new_P1_U3371, new_P1_U3372, new_P1_U3373,
    new_P1_U3374, new_P1_U3375, new_P1_U3376, new_P1_U3377, new_P1_U3378,
    new_P1_U3379, new_P1_U3380, new_P1_U3381, new_P1_U3382, new_P1_U3383,
    new_P1_U3384, new_P1_U3385, new_P1_U3386, new_P1_U3387, new_P1_U3388,
    new_P1_U3389, new_P1_U3390, new_P1_U3391, new_P1_U3392, new_P1_U3393,
    new_P1_U3394, new_P1_U3395, new_P1_U3396, new_P1_U3397, new_P1_U3398,
    new_P1_U3399, new_P1_U3400, new_P1_U3401, new_P1_U3402, new_P1_U3403,
    new_P1_U3404, new_P1_U3405, new_P1_U3406, new_P1_U3407, new_P1_U3408,
    new_P1_U3409, new_P1_U3410, new_P1_U3411, new_P1_U3412, new_P1_U3413,
    new_P1_U3414, new_P1_U3415, new_P1_U3416, new_P1_U3417, new_P1_U3418,
    new_P1_U3419, new_P1_U3420, new_P1_U3421, new_P1_U3422, new_P1_U3423,
    new_P1_U3424, new_P1_U3425, new_P1_U3426, new_P1_U3427, new_P1_U3428,
    new_P1_U3429, new_P1_U3430, new_P1_U3431, new_P1_U3432, new_P1_U3433,
    new_P1_U3434, new_P1_U3435, new_P1_U3436, new_P1_U3437, new_P1_U3438,
    new_P1_U3439, new_P1_U3440, new_P1_U3441, new_P1_U3442, new_P1_U3443,
    new_P1_U3444, new_P1_U3445, new_P1_U3446, new_P1_U3447, new_P1_U3448,
    new_P1_U3449, new_P1_U3450, new_P1_U3451, new_P1_U3452, new_P1_U3453,
    new_P1_U3454, new_P1_U3455, new_P1_U3456, new_P1_U3457, new_P1_U3462,
    new_P1_U3463, new_P1_U3467, new_P1_U3470, new_P1_U3471, new_P1_U3479,
    new_P1_U3480, new_P1_U3488, new_P1_U3489, new_P1_U3490, new_P1_U3491,
    new_P1_U3492, new_P1_U3493, new_P1_U3494, new_P1_U3495, new_P1_U3496,
    new_P1_U3497, new_P1_U3498, new_P1_U3499, new_P1_U3500, new_P1_U3501,
    new_P1_U3502, new_P1_U3503, new_P1_U3504, new_P1_U3505, new_P1_U3506,
    new_P1_U3507, new_P1_U3508, new_P1_U3509, new_P1_U3510, new_P1_U3511,
    new_P1_U3512, new_P1_U3513, new_P1_U3514, new_P1_U3515, new_P1_U3516,
    new_P1_U3517, new_P1_U3518, new_P1_U3519, new_P1_U3520, new_P1_U3521,
    new_P1_U3522, new_P1_U3523, new_P1_U3524, new_P1_U3525, new_P1_U3526,
    new_P1_U3527, new_P1_U3528, new_P1_U3529, new_P1_U3530, new_P1_U3531,
    new_P1_U3532, new_P1_U3533, new_P1_U3534, new_P1_U3535, new_P1_U3536,
    new_P1_U3537, new_P1_U3538, new_P1_U3539, new_P1_U3540, new_P1_U3541,
    new_P1_U3542, new_P1_U3543, new_P1_U3544, new_P1_U3545, new_P1_U3546,
    new_P1_U3547, new_P1_U3548, new_P1_U3549, new_P1_U3550, new_P1_U3551,
    new_P1_U3552, new_P1_U3553, new_P1_U3554, new_P1_U3555, new_P1_U3556,
    new_P1_U3557, new_P1_U3558, new_P1_U3559, new_P1_U3560, new_P1_U3561,
    new_P1_U3562, new_P1_U3563, new_P1_U3564, new_P1_U3565, new_P1_U3566,
    new_P1_U3567, new_P1_U3568, new_P1_U3569, new_P1_U3570, new_P1_U3571,
    new_P1_U3572, new_P1_U3573, new_P1_U3574, new_P1_U3575, new_P1_U3576,
    new_P1_U3577, new_P1_U3578, new_P1_U3579, new_P1_U3580, new_P1_U3581,
    new_P1_U3582, new_P1_U3583, new_P1_U3584, new_P1_U3585, new_P1_U3586,
    new_P1_U3587, new_P1_U3588, new_P1_U3589, new_P1_U3590, new_P1_U3591,
    new_P1_U3592, new_P1_U3593, new_P1_U3594, new_P1_U3595, new_P1_U3596,
    new_P1_U3597, new_P1_U3598, new_P1_U3599, new_P1_U3600, new_P1_U3601,
    new_P1_U3602, new_P1_U3603, new_P1_U3604, new_P1_U3605, new_P1_U3606,
    new_P1_U3607, new_P1_U3608, new_P1_U3609, new_P1_U3610, new_P1_U3611,
    new_P1_U3612, new_P1_U3613, new_P1_U3614, new_P1_U3615, new_P1_U3616,
    new_P1_U3617, new_P1_U3618, new_P1_U3619, new_P1_U3620, new_P1_U3621,
    new_P1_U3622, new_P1_U3623, new_P1_U3624, new_P1_U3625, new_P1_U3626,
    new_P1_U3627, new_P1_U3628, new_P1_U3629, new_P1_U3630, new_P1_U3631,
    new_P1_U3632, new_P1_U3633, new_P1_U3634, new_P1_U3635, new_P1_U3636,
    new_P1_U3637, new_P1_U3638, new_P1_U3639, new_P1_U3640, new_P1_U3641,
    new_P1_U3642, new_P1_U3643, new_P1_U3644, new_P1_U3645, new_P1_U3646,
    new_P1_U3647, new_P1_U3648, new_P1_U3649, new_P1_U3650, new_P1_U3651,
    new_P1_U3652, new_P1_U3653, new_P1_U3654, new_P1_U3655, new_P1_U3656,
    new_P1_U3657, new_P1_U3658, new_P1_U3659, new_P1_U3660, new_P1_U3661,
    new_P1_U3662, new_P1_U3663, new_P1_U3664, new_P1_U3665, new_P1_U3666,
    new_P1_U3667, new_P1_U3668, new_P1_U3669, new_P1_U3670, new_P1_U3671,
    new_P1_U3672, new_P1_U3673, new_P1_U3674, new_P1_U3675, new_P1_U3676,
    new_P1_U3677, new_P1_U3678, new_P1_U3679, new_P1_U3680, new_P1_U3681,
    new_P1_U3682, new_P1_U3683, new_P1_U3684, new_P1_U3685, new_P1_U3686,
    new_P1_U3687, new_P1_U3688, new_P1_U3689, new_P1_U3690, new_P1_U3691,
    new_P1_U3692, new_P1_U3693, new_P1_U3694, new_P1_U3695, new_P1_U3696,
    new_P1_U3697, new_P1_U3698, new_P1_U3699, new_P1_U3700, new_P1_U3701,
    new_P1_U3702, new_P1_U3703, new_P1_U3704, new_P1_U3705, new_P1_U3706,
    new_P1_U3707, new_P1_U3708, new_P1_U3709, new_P1_U3710, new_P1_U3711,
    new_P1_U3712, new_P1_U3713, new_P1_U3714, new_P1_U3715, new_P1_U3716,
    new_P1_U3717, new_P1_U3718, new_P1_U3719, new_P1_U3720, new_P1_U3721,
    new_P1_U3722, new_P1_U3723, new_P1_U3724, new_P1_U3725, new_P1_U3726,
    new_P1_U3727, new_P1_U3728, new_P1_U3729, new_P1_U3730, new_P1_U3731,
    new_P1_U3732, new_P1_U3733, new_P1_U3734, new_P1_U3735, new_P1_U3736,
    new_P1_U3737, new_P1_U3738, new_P1_U3739, new_P1_U3740, new_P1_U3741,
    new_P1_U3742, new_P1_U3743, new_P1_U3744, new_P1_U3745, new_P1_U3746,
    new_P1_U3747, new_P1_U3748, new_P1_U3749, new_P1_U3750, new_P1_U3751,
    new_P1_U3752, new_P1_U3753, new_P1_U3754, new_P1_U3755, new_P1_U3756,
    new_P1_U3757, new_P1_U3758, new_P1_U3759, new_P1_U3760, new_P1_U3761,
    new_P1_U3762, new_P1_U3763, new_P1_U3764, new_P1_U3765, new_P1_U3766,
    new_P1_U3767, new_P1_U3768, new_P1_U3769, new_P1_U3770, new_P1_U3771,
    new_P1_U3772, new_P1_U3773, new_P1_U3774, new_P1_U3775, new_P1_U3776,
    new_P1_U3777, new_P1_U3778, new_P1_U3779, new_P1_U3780, new_P1_U3781,
    new_P1_U3782, new_P1_U3783, new_P1_U3784, new_P1_U3785, new_P1_U3786,
    new_P1_U3787, new_P1_U3788, new_P1_U3789, new_P1_U3790, new_P1_U3791,
    new_P1_U3792, new_P1_U3793, new_P1_U3794, new_P1_U3795, new_P1_U3796,
    new_P1_U3797, new_P1_U3798, new_P1_U3799, new_P1_U3800, new_P1_U3801,
    new_P1_U3802, new_P1_U3803, new_P1_U3804, new_P1_U3805, new_P1_U3806,
    new_P1_U3807, new_P1_U3808, new_P1_U3809, new_P1_U3810, new_P1_U3811,
    new_P1_U3812, new_P1_U3813, new_P1_U3814, new_P1_U3815, new_P1_U3816,
    new_P1_U3817, new_P1_U3818, new_P1_U3819, new_P1_U3820, new_P1_U3821,
    new_P1_U3822, new_P1_U3823, new_P1_U3824, new_P1_U3825, new_P1_U3826,
    new_P1_U3827, new_P1_U3828, new_P1_U3829, new_P1_U3830, new_P1_U3831,
    new_P1_U3832, new_P1_U3833, new_P1_U3834, new_P1_U3835, new_P1_U3836,
    new_P1_U3837, new_P1_U3838, new_P1_U3839, new_P1_U3840, new_P1_U3841,
    new_P1_U3842, new_P1_U3843, new_P1_U3844, new_P1_U3845, new_P1_U3846,
    new_P1_U3847, new_P1_U3848, new_P1_U3849, new_P1_U3850, new_P1_U3851,
    new_P1_U3852, new_P1_U3853, new_P1_U3854, new_P1_U3855, new_P1_U3856,
    new_P1_U3857, new_P1_U3858, new_P1_U3859, new_P1_U3860, new_P1_U3861,
    new_P1_U3862, new_P1_U3863, new_P1_U3864, new_P1_U3865, new_P1_U3866,
    new_P1_U3867, new_P1_U3868, new_P1_U3869, new_P1_U3870, new_P1_U3871,
    new_P1_U3872, new_P1_U3873, new_P1_U3874, new_P1_U3875, new_P1_U3876,
    new_P1_U3877, new_P1_U3878, new_P1_U3879, new_P1_U3880, new_P1_U3881,
    new_P1_U3882, new_P1_U3883, new_P1_U3884, new_P1_U3885, new_P1_U3886,
    new_P1_U3887, new_P1_U3888, new_P1_U3889, new_P1_U3890, new_P1_U3891,
    new_P1_U3892, new_P1_U3893, new_P1_U3894, new_P1_U3895, new_P1_U3896,
    new_P1_U3897, new_P1_U3898, new_P1_U3899, new_P1_U3900, new_P1_U3901,
    new_P1_U3902, new_P1_U3903, new_P1_U3904, new_P1_U3905, new_P1_U3906,
    new_P1_U3907, new_P1_U3908, new_P1_U3909, new_P1_U3910, new_P1_U3911,
    new_P1_U3912, new_P1_U3913, new_P1_U3914, new_P1_U3915, new_P1_U3916,
    new_P1_U3917, new_P1_U3918, new_P1_U3919, new_P1_U3920, new_P1_U3921,
    new_P1_U3922, new_P1_U3923, new_P1_U3924, new_P1_U3925, new_P1_U3926,
    new_P1_U3927, new_P1_U3928, new_P1_U3929, new_P1_U3930, new_P1_U3931,
    new_P1_U3932, new_P1_U3933, new_P1_U3934, new_P1_U3935, new_P1_U3936,
    new_P1_U3937, new_P1_U3938, new_P1_U3939, new_P1_U3940, new_P1_U3941,
    new_P1_U3942, new_P1_U3943, new_P1_U3944, new_P1_U3945, new_P1_U3946,
    new_P1_U3947, new_P1_U3948, new_P1_U3949, new_P1_U3950, new_P1_U3951,
    new_P1_U3952, new_P1_U3953, new_P1_U3954, new_P1_U3955, new_P1_U3956,
    new_P1_U3957, new_P1_U3958, new_P1_U3959, new_P1_U3960, new_P1_U3961,
    new_P1_U3962, new_P1_U3963, new_P1_U3964, new_P1_U3965, new_P1_U3966,
    new_P1_U3967, new_P1_U3968, new_P1_U3969, new_P1_U3970, new_P1_U3971,
    new_P1_U3972, new_P1_U3973, new_P1_U3974, new_P1_U3975, new_P1_U3976,
    new_P1_U3977, new_P1_U3978, new_P1_U3979, new_P1_U3980, new_P1_U3981,
    new_P1_U3982, new_P1_U3983, new_P1_U3984, new_P1_U3985, new_P1_U3986,
    new_P1_U3987, new_P1_U3988, new_P1_U3989, new_P1_U3990, new_P1_U3991,
    new_P1_U3992, new_P1_U3993, new_P1_U3994, new_P1_U3995, new_P1_U3996,
    new_P1_U3997, new_P1_U3998, new_P1_U3999, new_P1_U4000, new_P1_U4001,
    new_P1_U4002, new_P1_U4003, new_P1_U4004, new_P1_U4005, new_P1_U4006,
    new_P1_U4007, new_P1_U4008, new_P1_U4009, new_P1_U4010, new_P1_U4011,
    new_P1_U4012, new_P1_U4013, new_P1_U4014, new_P1_U4015, new_P1_U4016,
    new_P1_U4017, new_P1_U4018, new_P1_U4019, new_P1_U4020, new_P1_U4021,
    new_P1_U4022, new_P1_U4023, new_P1_U4024, new_P1_U4025, new_P1_U4026,
    new_P1_U4027, new_P1_U4028, new_P1_U4029, new_P1_U4030, new_P1_U4031,
    new_P1_U4032, new_P1_U4033, new_P1_U4034, new_P1_U4035, new_P1_U4036,
    new_P1_U4037, new_P1_U4038, new_P1_U4039, new_P1_U4040, new_P1_U4041,
    new_P1_U4042, new_P1_U4043, new_P1_U4044, new_P1_U4045, new_P1_U4046,
    new_P1_U4047, new_P1_U4048, new_P1_U4049, new_P1_U4050, new_P1_U4051,
    new_P1_U4052, new_P1_U4053, new_P1_U4054, new_P1_U4055, new_P1_U4056,
    new_P1_U4057, new_P1_U4058, new_P1_U4059, new_P1_U4060, new_P1_U4061,
    new_P1_U4062, new_P1_U4063, new_P1_U4064, new_P1_U4065, new_P1_U4066,
    new_P1_U4067, new_P1_U4068, new_P1_U4069, new_P1_U4070, new_P1_U4071,
    new_P1_U4072, new_P1_U4073, new_P1_U4074, new_P1_U4075, new_P1_U4076,
    new_P1_U4077, new_P1_U4078, new_P1_U4079, new_P1_U4080, new_P1_U4081,
    new_P1_U4082, new_P1_U4083, new_P1_U4084, new_P1_U4085, new_P1_U4086,
    new_P1_U4087, new_P1_U4088, new_P1_U4089, new_P1_U4090, new_P1_U4091,
    new_P1_U4092, new_P1_U4093, new_P1_U4094, new_P1_U4095, new_P1_U4096,
    new_P1_U4097, new_P1_U4098, new_P1_U4099, new_P1_U4100, new_P1_U4101,
    new_P1_U4102, new_P1_U4103, new_P1_U4104, new_P1_U4105, new_P1_U4106,
    new_P1_U4107, new_P1_U4108, new_P1_U4109, new_P1_U4110, new_P1_U4111,
    new_P1_U4112, new_P1_U4113, new_P1_U4114, new_P1_U4115, new_P1_U4116,
    new_P1_U4117, new_P1_U4118, new_P1_U4119, new_P1_U4120, new_P1_U4121,
    new_P1_U4122, new_P1_U4123, new_P1_U4124, new_P1_U4125, new_P1_U4126,
    new_P1_U4127, new_P1_U4128, new_P1_U4129, new_P1_U4130, new_P1_U4131,
    new_P1_U4132, new_P1_U4133, new_P1_U4134, new_P1_U4135, new_P1_U4136,
    new_P1_U4137, new_P1_U4138, new_P1_U4139, new_P1_U4140, new_P1_U4141,
    new_P1_U4142, new_P1_U4143, new_P1_U4144, new_P1_U4145, new_P1_U4146,
    new_P1_U4147, new_P1_U4148, new_P1_U4149, new_P1_U4150, new_P1_U4151,
    new_P1_U4152, new_P1_U4153, new_P1_U4154, new_P1_U4155, new_P1_U4156,
    new_P1_U4157, new_P1_U4158, new_P1_U4159, new_P1_U4160, new_P1_U4161,
    new_P1_U4162, new_P1_U4163, new_P1_U4164, new_P1_U4165, new_P1_U4166,
    new_P1_U4167, new_P1_U4168, new_P1_U4169, new_P1_U4170, new_P1_U4171,
    new_P1_U4172, new_P1_U4173, new_P1_U4174, new_P1_U4175, new_P1_U4176,
    new_P1_U4177, new_P1_U4178, new_P1_U4179, new_P1_U4180, new_P1_U4181,
    new_P1_U4182, new_P1_U4183, new_P1_U4184, new_P1_U4185, new_P1_U4186,
    new_P1_U4187, new_P1_U4188, new_P1_U4189, new_P1_U4190, new_P1_U4191,
    new_P1_U4192, new_P1_U4193, new_P1_U4194, new_P1_U4195, new_P1_U4196,
    new_P1_U4197, new_P1_U4198, new_P1_U4199, new_P1_U4200, new_P1_U4201,
    new_P1_U4202, new_P1_U4203, new_P1_U4204, new_P1_U4205, new_P1_U4206,
    new_P1_U4207, new_P1_U4208, new_P1_U4209, new_P1_U4210, new_P1_U4211,
    new_P1_U4212, new_P1_U4213, new_P1_U4214, new_P1_U4215, new_P1_U4216,
    new_P1_U4217, new_P1_U4218, new_P1_U4219, new_P1_U4220, new_P1_U4221,
    new_P1_U4222, new_P1_U4223, new_P1_U4224, new_P1_U4225, new_P1_U4226,
    new_P1_U4227, new_P1_U4228, new_P1_U4229, new_P1_U4230, new_P1_U4231,
    new_P1_U4232, new_P1_U4233, new_P1_U4234, new_P1_U4235, new_P1_U4236,
    new_P1_U4237, new_P1_U4238, new_P1_U4239, new_P1_U4240, new_P1_U4241,
    new_P1_U4242, new_P1_U4243, new_P1_U4244, new_P1_U4245, new_P1_U4246,
    new_P1_U4247, new_P1_U4248, new_P1_U4249, new_P1_U4250, new_P1_U4251,
    new_P1_U4252, new_P1_U4253, new_P1_U4254, new_P1_U4255, new_P1_U4256,
    new_P1_U4257, new_P1_U4258, new_P1_U4259, new_P1_U4260, new_P1_U4261,
    new_P1_U4262, new_P1_U4263, new_P1_U4264, new_P1_U4265, new_P1_U4266,
    new_P1_U4267, new_P1_U4268, new_P1_U4269, new_P1_U4270, new_P1_U4271,
    new_P1_U4272, new_P1_U4273, new_P1_U4274, new_P1_U4275, new_P1_U4276,
    new_P1_U4277, new_P1_U4278, new_P1_U4279, new_P1_U4280, new_P1_U4281,
    new_P1_U4282, new_P1_U4283, new_P1_U4284, new_P1_U4285, new_P1_U4286,
    new_P1_U4287, new_P1_U4288, new_P1_U4289, new_P1_U4290, new_P1_U4291,
    new_P1_U4292, new_P1_U4293, new_P1_U4294, new_P1_U4295, new_P1_U4296,
    new_P1_U4297, new_P1_U4298, new_P1_U4299, new_P1_U4300, new_P1_U4301,
    new_P1_U4302, new_P1_U4303, new_P1_U4304, new_P1_U4305, new_P1_U4306,
    new_P1_U4307, new_P1_U4308, new_P1_U4309, new_P1_U4310, new_P1_U4311,
    new_P1_U4312, new_P1_U4313, new_P1_U4314, new_P1_U4315, new_P1_U4316,
    new_P1_U4317, new_P1_U4318, new_P1_U4319, new_P1_U4320, new_P1_U4321,
    new_P1_U4322, new_P1_U4323, new_P1_U4324, new_P1_U4325, new_P1_U4326,
    new_P1_U4327, new_P1_U4328, new_P1_U4329, new_P1_U4330, new_P1_U4331,
    new_P1_U4332, new_P1_U4333, new_P1_U4334, new_P1_U4335, new_P1_U4336,
    new_P1_U4337, new_P1_U4338, new_P1_U4339, new_P1_U4340, new_P1_U4341,
    new_P1_U4342, new_P1_U4343, new_P1_U4344, new_P1_U4345, new_P1_U4346,
    new_P1_U4347, new_P1_U4348, new_P1_U4349, new_P1_U4350, new_P1_U4351,
    new_P1_U4352, new_P1_U4353, new_P1_U4354, new_P1_U4355, new_P1_U4356,
    new_P1_U4357, new_P1_U4358, new_P1_U4359, new_P1_U4360, new_P1_U4361,
    new_P1_U4362, new_P1_U4363, new_P1_U4364, new_P1_U4365, new_P1_U4366,
    new_P1_U4367, new_P1_U4368, new_P1_U4369, new_P1_U4370, new_P1_U4371,
    new_P1_U4372, new_P1_U4373, new_P1_U4374, new_P1_U4375, new_P1_U4376,
    new_P1_U4377, new_P1_U4378, new_P1_U4379, new_P1_U4380, new_P1_U4381,
    new_P1_U4382, new_P1_U4383, new_P1_U4384, new_P1_U4385, new_P1_U4386,
    new_P1_U4387, new_P1_U4388, new_P1_U4389, new_P1_U4390, new_P1_U4391,
    new_P1_U4392, new_P1_U4393, new_P1_U4394, new_P1_U4395, new_P1_U4396,
    new_P1_U4397, new_P1_U4398, new_P1_U4399, new_P1_U4400, new_P1_U4401,
    new_P1_U4402, new_P1_U4403, new_P1_U4404, new_P1_U4405, new_P1_U4406,
    new_P1_U4407, new_P1_U4408, new_P1_U4409, new_P1_U4410, new_P1_U4411,
    new_P1_U4412, new_P1_U4413, new_P1_U4414, new_P1_U4415, new_P1_U4416,
    new_P1_U4417, new_P1_U4418, new_P1_U4419, new_P1_U4420, new_P1_U4421,
    new_P1_U4422, new_P1_U4423, new_P1_U4424, new_P1_U4425, new_P1_U4426,
    new_P1_U4427, new_P1_U4428, new_P1_U4429, new_P1_U4430, new_P1_U4431,
    new_P1_U4432, new_P1_U4433, new_P1_U4434, new_P1_U4435, new_P1_U4436,
    new_P1_U4437, new_P1_U4438, new_P1_U4439, new_P1_U4440, new_P1_U4441,
    new_P1_U4442, new_P1_U4443, new_P1_U4444, new_P1_U4445, new_P1_U4446,
    new_P1_U4447, new_P1_U4448, new_P1_U4449, new_P1_U4450, new_P1_U4451,
    new_P1_U4452, new_P1_U4453, new_P1_U4454, new_P1_U4455, new_P1_U4456,
    new_P1_U4457, new_P1_U4458, new_P1_U4459, new_P1_U4460, new_P1_U4461,
    new_P1_U4462, new_P1_U4463, new_P1_U4464, new_P1_U4465, new_P1_U4466,
    new_P1_U4467, new_P1_U4468, new_P1_U4469, new_P1_U4470, new_P1_U4471,
    new_P1_U4472, new_P1_U4473, new_P1_U4474, new_P1_U4475, new_P1_U4476,
    new_P1_U4477, new_P1_U4478, new_P1_U4479, new_P1_U4480, new_P1_U4481,
    new_P1_U4482, new_P1_U4483, new_P1_U4484, new_P1_U4485, new_P1_U4486,
    new_P1_U4487, new_P1_U4488, new_P1_U4489, new_P1_U4490, new_P1_U4491,
    new_P1_U4492, new_P1_U4493, new_P1_U4494, new_P1_U4495, new_P1_U4496,
    new_P1_U4497, new_P1_U4498, new_P1_U4499, new_P1_U4500, new_P1_U4501,
    new_P1_U4502, new_P1_U4503, new_P1_U4504, new_P1_U4505, new_P1_U4506,
    new_P1_U4507, new_P1_U4508, new_P1_U4509, new_P1_U4510, new_P1_U4511,
    new_P1_U4512, new_P1_U4513, new_P1_U4514, new_P1_U4515, new_P1_U4516,
    new_P1_U4517, new_P1_U4518, new_P1_U4519, new_P1_U4520, new_P1_U4521,
    new_P1_U4522, new_P1_U4523, new_P1_U4524, new_P1_U4525, new_P1_U4526,
    new_P1_U4527, new_P1_U4528, new_P1_U4529, new_P1_U4530, new_P1_U4531,
    new_P1_U4532, new_P1_U4533, new_P1_U4534, new_P1_U4535, new_P1_U4536,
    new_P1_U4537, new_P1_U4538, new_P1_U4539, new_P1_U4540, new_P1_U4541,
    new_P1_U4542, new_P1_U4543, new_P1_U4544, new_P1_U4545, new_P1_U4546,
    new_P1_U4547, new_P1_U4548, new_P1_U4549, new_P1_U4550, new_P1_U4551,
    new_P1_U4552, new_P1_U4553, new_P1_U4554, new_P1_U4555, new_P1_U4556,
    new_P1_U4557, new_P1_U4558, new_P1_U4559, new_P1_U4560, new_P1_U4561,
    new_P1_U4562, new_P1_U4563, new_P1_U4564, new_P1_U4565, new_P1_U4566,
    new_P1_U4567, new_P1_U4568, new_P1_U4569, new_P1_U4570, new_P1_U4571,
    new_P1_U4572, new_P1_U4573, new_P1_U4574, new_P1_U4575, new_P1_U4576,
    new_P1_U4577, new_P1_U4578, new_P1_U4579, new_P1_U4580, new_P1_U4581,
    new_P1_U4582, new_P1_U4583, new_P1_U4584, new_P1_U4585, new_P1_U4586,
    new_P1_U4587, new_P1_U4588, new_P1_U4589, new_P1_U4590, new_P1_U4591,
    new_P1_U4592, new_P1_U4593, new_P1_U4594, new_P1_U4595, new_P1_U4596,
    new_P1_U4597, new_P1_U4598, new_P1_U4599, new_P1_U4600, new_P1_U4601,
    new_P1_U4602, new_P1_U4603, new_P1_U4604, new_P1_U4605, new_P1_U4606,
    new_P1_U4607, new_P1_U4608, new_P1_U4609, new_P1_U4610, new_P1_U4611,
    new_P1_U4612, new_P1_U4613, new_P1_U4614, new_P1_U4615, new_P1_U4616,
    new_P1_U4617, new_P1_U4618, new_P1_U4619, new_P1_U4620, new_P1_U4621,
    new_P1_U4622, new_P1_U4623, new_P1_U4624, new_P1_U4625, new_P1_U4626,
    new_P1_U4627, new_P1_U4628, new_P1_U4629, new_P1_U4630, new_P1_U4631,
    new_P1_U4632, new_P1_U4633, new_P1_U4634, new_P1_U4635, new_P1_U4636,
    new_P1_U4637, new_P1_U4638, new_P1_U4639, new_P1_U4640, new_P1_U4641,
    new_P1_U4642, new_P1_U4643, new_P1_U4644, new_P1_U4645, new_P1_U4646,
    new_P1_U4647, new_P1_U4648, new_P1_U4649, new_P1_U4650, new_P1_U4651,
    new_P1_U4652, new_P1_U4653, new_P1_U4654, new_P1_U4655, new_P1_U4656,
    new_P1_U4657, new_P1_U4658, new_P1_U4659, new_P1_U4660, new_P1_U4661,
    new_P1_U4662, new_P1_U4663, new_P1_U4664, new_P1_U4665, new_P1_U4666,
    new_P1_U4667, new_P1_U4668, new_P1_U4669, new_P1_U4670, new_P1_U4671,
    new_P1_U4672, new_P1_U4673, new_P1_U4674, new_P1_U4675, new_P1_U4676,
    new_P1_U4677, new_P1_U4678, new_P1_U4679, new_P1_U4680, new_P1_U4681,
    new_P1_U4682, new_P1_U4683, new_P1_U4684, new_P1_U4685, new_P1_U4686,
    new_P1_U4687, new_P1_U4688, new_P1_U4689, new_P1_U4690, new_P1_U4691,
    new_P1_U4692, new_P1_U4693, new_P1_U4694, new_P1_U4695, new_P1_U4696,
    new_P1_U4697, new_P1_U4698, new_P1_U4699, new_P1_U4700, new_P1_U4701,
    new_P1_U4702, new_P1_U4703, new_P1_U4704, new_P1_U4705, new_P1_U4706,
    new_P1_U4707, new_P1_U4708, new_P1_U4709, new_P1_U4710, new_P1_U4711,
    new_P1_U4712, new_P1_U4713, new_P1_U4714, new_P1_U4715, new_P1_U4716,
    new_P1_U4717, new_P1_U4718, new_P1_U4719, new_P1_U4720, new_P1_U4721,
    new_P1_U4722, new_P1_U4723, new_P1_U4724, new_P1_U4725, new_P1_U4726,
    new_P1_U4727, new_P1_U4728, new_P1_U4729, new_P1_U4730, new_P1_U4731,
    new_P1_U4732, new_P1_U4733, new_P1_U4734, new_P1_U4735, new_P1_U4736,
    new_P1_U4737, new_P1_U4738, new_P1_U4739, new_P1_U4740, new_P1_U4741,
    new_P1_U4742, new_P1_U4743, new_P1_U4744, new_P1_U4745, new_P1_U4746,
    new_P1_U4747, new_P1_U4748, new_P1_U4749, new_P1_U4750, new_P1_U4751,
    new_P1_U4752, new_P1_U4753, new_P1_U4754, new_P1_U4755, new_P1_U4756,
    new_P1_U4757, new_P1_U4758, new_P1_U4759, new_P1_U4760, new_P1_U4761,
    new_P1_U4762, new_P1_U4763, new_P1_U4764, new_P1_U4765, new_P1_U4766,
    new_P1_U4767, new_P1_U4768, new_P1_U4769, new_P1_U4770, new_P1_U4771,
    new_P1_U4772, new_P1_U4773, new_P1_U4774, new_P1_U4775, new_P1_U4776,
    new_P1_U4777, new_P1_U4778, new_P1_U4779, new_P1_U4780, new_P1_U4781,
    new_P1_U4782, new_P1_U4783, new_P1_U4784, new_P1_U4785, new_P1_U4786,
    new_P1_U4787, new_P1_U4788, new_P1_U4789, new_P1_U4790, new_P1_U4791,
    new_P1_U4792, new_P1_U4793, new_P1_U4794, new_P1_U4795, new_P1_U4796,
    new_P1_U4797, new_P1_U4798, new_P1_U4799, new_P1_U4800, new_P1_U4801,
    new_P1_U4802, new_P1_U4803, new_P1_U4804, new_P1_U4805, new_P1_U4806,
    new_P1_U4807, new_P1_U4808, new_P1_U4809, new_P1_U4810, new_P1_U4811,
    new_P1_U4812, new_P1_U4813, new_P1_U4814, new_P1_U4815, new_P1_U4816,
    new_P1_U4817, new_P1_U4818, new_P1_U4819, new_P1_U4820, new_P1_U4821,
    new_P1_U4822, new_P1_U4823, new_P1_U4824, new_P1_U4825, new_P1_U4826,
    new_P1_U4827, new_P1_U4828, new_P1_U4829, new_P1_U4830, new_P1_U4831,
    new_P1_U4832, new_P1_U4833, new_P1_U4834, new_P1_U4835, new_P1_U4836,
    new_P1_U4837, new_P1_U4838, new_P1_U4839, new_P1_U4840, new_P1_U4841,
    new_P1_U4842, new_P1_U4843, new_P1_U4844, new_P1_U4845, new_P1_U4846,
    new_P1_U4847, new_P1_U4848, new_P1_U4849, new_P1_U4850, new_P1_U4851,
    new_P1_U4852, new_P1_U4853, new_P1_U4854, new_P1_U4855, new_P1_U4856,
    new_P1_U4857, new_P1_U4858, new_P1_U4859, new_P1_U4860, new_P1_U4861,
    new_P1_U4862, new_P1_U4863, new_P1_U4864, new_P1_U4865, new_P1_U4866,
    new_P1_U4867, new_P1_U4868, new_P1_U4869, new_P1_U4870, new_P1_U4871,
    new_P1_U4872, new_P1_U4873, new_P1_U4874, new_P1_U4875, new_P1_U4876,
    new_P1_U4877, new_P1_U4878, new_P1_U4879, new_P1_U4880, new_P1_U4881,
    new_P1_U4882, new_P1_U4883, new_P1_U4884, new_P1_U4885, new_P1_U4886,
    new_P1_U4887, new_P1_U4888, new_P1_U4889, new_P1_U4890, new_P1_U4891,
    new_P1_U4892, new_P1_U4893, new_P1_U4894, new_P1_U4895, new_P1_U4896,
    new_P1_U4897, new_P1_U4898, new_P1_U4899, new_P1_U4900, new_P1_U4901,
    new_P1_U4902, new_P1_U4903, new_P1_U4904, new_P1_U4905, new_P1_U4906,
    new_P1_U4907, new_P1_U4908, new_P1_U4909, new_P1_U4910, new_P1_U4911,
    new_P1_U4912, new_P1_U4913, new_P1_U4914, new_P1_U4915, new_P1_U4916,
    new_P1_U4917, new_P1_U4918, new_P1_U4919, new_P1_U4920, new_P1_U4921,
    new_P1_U4922, new_P1_U4923, new_P1_U4924, new_P1_U4925, new_P1_U4926,
    new_P1_U4927, new_P1_U4928, new_P1_U4929, new_P1_U4930, new_P1_U4931,
    new_P1_U4932, new_P1_U4933, new_P1_U4934, new_P1_U4935, new_P1_U4936,
    new_P1_U4937, new_P1_U4938, new_P1_U4939, new_P1_U4940, new_P1_U4941,
    new_P1_U4942, new_P1_U4943, new_P1_U4944, new_P1_U4945, new_P1_U4946,
    new_P1_U4947, new_P1_U4948, new_P1_U4949, new_P1_U4950, new_P1_U4951,
    new_P1_U4952, new_P1_U4953, new_P1_U4954, new_P1_U4955, new_P1_U4956,
    new_P1_U4957, new_P1_U4958, new_P1_U4959, new_P1_U4960, new_P1_U4961,
    new_P1_U4962, new_P1_U4963, new_P1_U4964, new_P1_U4965, new_P1_U4966,
    new_P1_U4967, new_P1_U4968, new_P1_U4969, new_P1_U4970, new_P1_U4971,
    new_P1_U4972, new_P1_U4973, new_P1_U4974, new_P1_U4975, new_P1_U4976,
    new_P1_U4977, new_P1_U4978, new_P1_U4979, new_P1_U4980, new_P1_U4981,
    new_P1_U4982, new_P1_U4983, new_P1_U4984, new_P1_U4985, new_P1_U4986,
    new_P1_U4987, new_P1_U4988, new_P1_U4989, new_P1_U4990, new_P1_U4991,
    new_P1_U4992, new_P1_U4993, new_P1_U4994, new_P1_U4995, new_P1_U4996,
    new_P1_U4997, new_P1_U4998, new_P1_U4999, new_P1_U5000, new_P1_U5001,
    new_P1_U5002, new_P1_U5003, new_P1_U5004, new_P1_U5005, new_P1_U5006,
    new_P1_U5007, new_P1_U5008, new_P1_U5009, new_P1_U5010, new_P1_U5011,
    new_P1_U5012, new_P1_U5013, new_P1_U5014, new_P1_U5015, new_P1_U5016,
    new_P1_U5017, new_P1_U5018, new_P1_U5019, new_P1_U5020, new_P1_U5021,
    new_P1_U5022, new_P1_U5023, new_P1_U5024, new_P1_U5025, new_P1_U5026,
    new_P1_U5027, new_P1_U5028, new_P1_U5029, new_P1_U5030, new_P1_U5031,
    new_P1_U5032, new_P1_U5033, new_P1_U5034, new_P1_U5035, new_P1_U5036,
    new_P1_U5037, new_P1_U5038, new_P1_U5039, new_P1_U5040, new_P1_U5041,
    new_P1_U5042, new_P1_U5043, new_P1_U5044, new_P1_U5045, new_P1_U5046,
    new_P1_U5047, new_P1_U5048, new_P1_U5049, new_P1_U5050, new_P1_U5051,
    new_P1_U5052, new_P1_U5053, new_P1_U5054, new_P1_U5055, new_P1_U5056,
    new_P1_U5057, new_P1_U5058, new_P1_U5059, new_P1_U5060, new_P1_U5061,
    new_P1_U5062, new_P1_U5063, new_P1_U5064, new_P1_U5065, new_P1_U5066,
    new_P1_U5067, new_P1_U5068, new_P1_U5069, new_P1_U5070, new_P1_U5071,
    new_P1_U5072, new_P1_U5073, new_P1_U5074, new_P1_U5075, new_P1_U5076,
    new_P1_U5077, new_P1_U5078, new_P1_U5079, new_P1_U5080, new_P1_U5081,
    new_P1_U5082, new_P1_U5083, new_P1_U5084, new_P1_U5085, new_P1_U5086,
    new_P1_U5087, new_P1_U5088, new_P1_U5089, new_P1_U5090, new_P1_U5091,
    new_P1_U5092, new_P1_U5093, new_P1_U5094, new_P1_U5095, new_P1_U5096,
    new_P1_U5097, new_P1_U5098, new_P1_U5099, new_P1_U5100, new_P1_U5101,
    new_P1_U5102, new_P1_U5103, new_P1_U5104, new_P1_U5105, new_P1_U5106,
    new_P1_U5107, new_P1_U5108, new_P1_U5109, new_P1_U5110, new_P1_U5111,
    new_P1_U5112, new_P1_U5113, new_P1_U5114, new_P1_U5115, new_P1_U5116,
    new_P1_U5117, new_P1_U5118, new_P1_U5119, new_P1_U5120, new_P1_U5121,
    new_P1_U5122, new_P1_U5123, new_P1_U5124, new_P1_U5125, new_P1_U5126,
    new_P1_U5127, new_P1_U5128, new_P1_U5129, new_P1_U5130, new_P1_U5131,
    new_P1_U5132, new_P1_U5133, new_P1_U5134, new_P1_U5135, new_P1_U5136,
    new_P1_U5137, new_P1_U5138, new_P1_U5139, new_P1_U5140, new_P1_U5141,
    new_P1_U5142, new_P1_U5143, new_P1_U5144, new_P1_U5145, new_P1_U5146,
    new_P1_U5147, new_P1_U5148, new_P1_U5149, new_P1_U5150, new_P1_U5151,
    new_P1_U5152, new_P1_U5153, new_P1_U5154, new_P1_U5155, new_P1_U5156,
    new_P1_U5157, new_P1_U5158, new_P1_U5159, new_P1_U5160, new_P1_U5161,
    new_P1_U5162, new_P1_U5163, new_P1_U5164, new_P1_U5165, new_P1_U5166,
    new_P1_U5167, new_P1_U5168, new_P1_U5169, new_P1_U5170, new_P1_U5171,
    new_P1_U5172, new_P1_U5173, new_P1_U5174, new_P1_U5175, new_P1_U5176,
    new_P1_U5177, new_P1_U5178, new_P1_U5179, new_P1_U5180, new_P1_U5181,
    new_P1_U5182, new_P1_U5183, new_P1_U5184, new_P1_U5185, new_P1_U5186,
    new_P1_U5187, new_P1_U5188, new_P1_U5189, new_P1_U5190, new_P1_U5191,
    new_P1_U5192, new_P1_U5193, new_P1_U5194, new_P1_U5195, new_P1_U5196,
    new_P1_U5197, new_P1_U5198, new_P1_U5199, new_P1_U5200, new_P1_U5201,
    new_P1_U5202, new_P1_U5203, new_P1_U5204, new_P1_U5205, new_P1_U5206,
    new_P1_U5207, new_P1_U5208, new_P1_U5209, new_P1_U5210, new_P1_U5211,
    new_P1_U5212, new_P1_U5213, new_P1_U5214, new_P1_U5215, new_P1_U5216,
    new_P1_U5217, new_P1_U5218, new_P1_U5219, new_P1_U5220, new_P1_U5221,
    new_P1_U5222, new_P1_U5223, new_P1_U5224, new_P1_U5225, new_P1_U5226,
    new_P1_U5227, new_P1_U5228, new_P1_U5229, new_P1_U5230, new_P1_U5231,
    new_P1_U5232, new_P1_U5233, new_P1_U5234, new_P1_U5235, new_P1_U5236,
    new_P1_U5237, new_P1_U5238, new_P1_U5239, new_P1_U5240, new_P1_U5241,
    new_P1_U5242, new_P1_U5243, new_P1_U5244, new_P1_U5245, new_P1_U5246,
    new_P1_U5247, new_P1_U5248, new_P1_U5249, new_P1_U5250, new_P1_U5251,
    new_P1_U5252, new_P1_U5253, new_P1_U5254, new_P1_U5255, new_P1_U5256,
    new_P1_U5257, new_P1_U5258, new_P1_U5259, new_P1_U5260, new_P1_U5261,
    new_P1_U5262, new_P1_U5263, new_P1_U5264, new_P1_U5265, new_P1_U5266,
    new_P1_U5267, new_P1_U5268, new_P1_U5269, new_P1_U5270, new_P1_U5271,
    new_P1_U5272, new_P1_U5273, new_P1_U5274, new_P1_U5275, new_P1_U5276,
    new_P1_U5277, new_P1_U5278, new_P1_U5279, new_P1_U5280, new_P1_U5281,
    new_P1_U5282, new_P1_U5283, new_P1_U5284, new_P1_U5285, new_P1_U5286,
    new_P1_U5287, new_P1_U5288, new_P1_U5289, new_P1_U5290, new_P1_U5291,
    new_P1_U5292, new_P1_U5293, new_P1_U5294, new_P1_U5295, new_P1_U5296,
    new_P1_U5297, new_P1_U5298, new_P1_U5299, new_P1_U5300, new_P1_U5301,
    new_P1_U5302, new_P1_U5303, new_P1_U5304, new_P1_U5305, new_P1_U5306,
    new_P1_U5307, new_P1_U5308, new_P1_U5309, new_P1_U5310, new_P1_U5311,
    new_P1_U5312, new_P1_U5313, new_P1_U5314, new_P1_U5315, new_P1_U5316,
    new_P1_U5317, new_P1_U5318, new_P1_U5319, new_P1_U5320, new_P1_U5321,
    new_P1_U5322, new_P1_U5323, new_P1_U5324, new_P1_U5325, new_P1_U5326,
    new_P1_U5327, new_P1_U5328, new_P1_U5329, new_P1_U5330, new_P1_U5331,
    new_P1_U5332, new_P1_U5333, new_P1_U5334, new_P1_U5335, new_P1_U5336,
    new_P1_U5337, new_P1_U5338, new_P1_U5339, new_P1_U5340, new_P1_U5341,
    new_P1_U5342, new_P1_U5343, new_P1_U5344, new_P1_U5345, new_P1_U5346,
    new_P1_U5347, new_P1_U5348, new_P1_U5349, new_P1_U5350, new_P1_U5351,
    new_P1_U5352, new_P1_U5353, new_P1_U5354, new_P1_U5355, new_P1_U5356,
    new_P1_U5357, new_P1_U5358, new_P1_U5359, new_P1_U5360, new_P1_U5361,
    new_P1_U5362, new_P1_U5363, new_P1_U5364, new_P1_U5365, new_P1_U5366,
    new_P1_U5367, new_P1_U5368, new_P1_U5369, new_P1_U5370, new_P1_U5371,
    new_P1_U5372, new_P1_U5373, new_P1_U5374, new_P1_U5375, new_P1_U5376,
    new_P1_U5377, new_P1_U5378, new_P1_U5379, new_P1_U5380, new_P1_U5381,
    new_P1_U5382, new_P1_U5383, new_P1_U5384, new_P1_U5385, new_P1_U5386,
    new_P1_U5387, new_P1_U5388, new_P1_U5389, new_P1_U5390, new_P1_U5391,
    new_P1_U5392, new_P1_U5393, new_P1_U5394, new_P1_U5395, new_P1_U5396,
    new_P1_U5397, new_P1_U5398, new_P1_U5399, new_P1_U5400, new_P1_U5401,
    new_P1_U5402, new_P1_U5403, new_P1_U5404, new_P1_U5405, new_P1_U5406,
    new_P1_U5407, new_P1_U5408, new_P1_U5409, new_P1_U5410, new_P1_U5411,
    new_P1_U5412, new_P1_U5413, new_P1_U5414, new_P1_U5415, new_P1_U5416,
    new_P1_U5417, new_P1_U5418, new_P1_U5419, new_P1_U5420, new_P1_U5421,
    new_P1_U5422, new_P1_U5423, new_P1_U5424, new_P1_U5425, new_P1_U5426,
    new_P1_U5427, new_P1_U5428, new_P1_U5429, new_P1_U5430, new_P1_U5431,
    new_P1_U5432, new_P1_U5433, new_P1_U5434, new_P1_U5435, new_P1_U5436,
    new_P1_U5437, new_P1_U5438, new_P1_U5439, new_P1_U5440, new_P1_U5441,
    new_P1_U5442, new_P1_U5443, new_P1_U5444, new_P1_U5445, new_P1_U5446,
    new_P1_U5447, new_P1_U5448, new_P1_U5449, new_P1_U5450, new_P1_U5451,
    new_P1_U5452, new_P1_U5453, new_P1_U5454, new_P1_U5455, new_P1_U5456,
    new_P1_U5457, new_P1_U5458, new_P1_U5459, new_P1_U5460, new_P1_U5461,
    new_P1_U5462, new_P1_U5463, new_P1_U5464, new_P1_U5465, new_P1_U5466,
    new_P1_U5467, new_P1_U5468, new_P1_U5469, new_P1_U5470, new_P1_U5471,
    new_P1_U5472, new_P1_U5473, new_P1_U5474, new_P1_U5475, new_P1_U5476,
    new_P1_U5477, new_P1_U5478, new_P1_U5479, new_P1_U5480, new_P1_U5481,
    new_P1_U5482, new_P1_U5483, new_P1_U5484, new_P1_U5485, new_P1_U5486,
    new_P1_U5487, new_P1_U5488, new_P1_U5489, new_P1_U5490, new_P1_U5491,
    new_P1_U5492, new_P1_U5493, new_P1_U5494, new_P1_U5495, new_P1_U5496,
    new_P1_U5497, new_P1_U5498, new_P1_U5499, new_P1_U5500, new_P1_U5501,
    new_P1_U5502, new_P1_U5503, new_P1_U5504, new_P1_U5505, new_P1_U5506,
    new_P1_U5507, new_P1_U5508, new_P1_U5509, new_P1_U5510, new_P1_U5511,
    new_P1_U5512, new_P1_U5513, new_P1_U5514, new_P1_U5515, new_P1_U5516,
    new_P1_U5517, new_P1_U5518, new_P1_U5519, new_P1_U5520, new_P1_U5521,
    new_P1_U5522, new_P1_U5523, new_P1_U5524, new_P1_U5525, new_P1_U5526,
    new_P1_U5527, new_P1_U5528, new_P1_U5529, new_P1_U5530, new_P1_U5531,
    new_P1_U5532, new_P1_U5533, new_P1_U5534, new_P1_U5535, new_P1_U5536,
    new_P1_U5537, new_P1_U5538, new_P1_U5539, new_P1_U5540, new_P1_U5541,
    new_P1_U5542, new_P1_U5543, new_P1_U5544, new_P1_U5545, new_P1_U5546,
    new_P1_U5547, new_P1_U5548, new_P1_U5549, new_P1_U5550, new_P1_U5551,
    new_P1_U5552, new_P1_U5553, new_P1_U5554, new_P1_U5555, new_P1_U5556,
    new_P1_U5557, new_P1_U5558, new_P1_U5559, new_P1_U5560, new_P1_U5561,
    new_P1_U5562, new_P1_U5563, new_P1_U5564, new_P1_U5565, new_P1_U5566,
    new_P1_U5567, new_P1_U5568, new_P1_U5569, new_P1_U5570, new_P1_U5571,
    new_P1_U5572, new_P1_U5573, new_P1_U5574, new_P1_U5575, new_P1_U5576,
    new_P1_U5577, new_P1_U5578, new_P1_U5579, new_P1_U5580, new_P1_U5581,
    new_P1_U5582, new_P1_U5583, new_P1_U5584, new_P1_U5585, new_P1_U5586,
    new_P1_U5587, new_P1_U5588, new_P1_U5589, new_P1_U5590, new_P1_U5591,
    new_P1_U5592, new_P1_U5593, new_P1_U5594, new_P1_U5595, new_P1_U5596,
    new_P1_U5597, new_P1_U5598, new_P1_U5599, new_P1_U5600, new_P1_U5601,
    new_P1_U5602, new_P1_U5603, new_P1_U5604, new_P1_U5605, new_P1_U5606,
    new_P1_U5607, new_P1_U5608, new_P1_U5609, new_P1_U5610, new_P1_U5611,
    new_P1_U5612, new_P1_U5613, new_P1_U5614, new_P1_U5615, new_P1_U5616,
    new_P1_U5617, new_P1_U5618, new_P1_U5619, new_P1_U5620, new_P1_U5621,
    new_P1_U5622, new_P1_U5623, new_P1_U5624, new_P1_U5625, new_P1_U5626,
    new_P1_U5627, new_P1_U5628, new_P1_U5629, new_P1_U5630, new_P1_U5631,
    new_P1_U5632, new_P1_U5633, new_P1_U5634, new_P1_U5635, new_P1_U5636,
    new_P1_U5637, new_P1_U5638, new_P1_U5639, new_P1_U5640, new_P1_U5641,
    new_P1_U5642, new_P1_U5643, new_P1_U5644, new_P1_U5645, new_P1_U5646,
    new_P1_U5647, new_P1_U5648, new_P1_U5649, new_P1_U5650, new_P1_U5651,
    new_P1_U5652, new_P1_U5653, new_P1_U5654, new_P1_U5655, new_P1_U5656,
    new_P1_U5657, new_P1_U5658, new_P1_U5659, new_P1_U5660, new_P1_U5661,
    new_P1_U5662, new_P1_U5663, new_P1_U5664, new_P1_U5665, new_P1_U5666,
    new_P1_U5667, new_P1_U5668, new_P1_U5669, new_P1_U5670, new_P1_U5671,
    new_P1_U5672, new_P1_U5673, new_P1_U5674, new_P1_U5675, new_P1_U5676,
    new_P1_U5677, new_P1_U5678, new_P1_U5679, new_P1_U5680, new_P1_U5681,
    new_P1_U5682, new_P1_U5683, new_P1_U5684, new_P1_U5685, new_P1_U5686,
    new_P1_U5687, new_P1_U5688, new_P1_U5689, new_P1_U5690, new_P1_U5691,
    new_P1_U5692, new_P1_U5693, new_P1_U5694, new_P1_U5695, new_P1_U5696,
    new_P1_U5697, new_P1_U5698, new_P1_U5699, new_P1_U5700, new_P1_U5701,
    new_P1_U5702, new_P1_U5703, new_P1_U5704, new_P1_U5705, new_P1_U5706,
    new_P1_U5707, new_P1_U5708, new_P1_U5709, new_P1_U5710, new_P1_U5711,
    new_P1_U5712, new_P1_U5713, new_P1_U5714, new_P1_U5715, new_P1_U5716,
    new_P1_U5717, new_P1_U5718, new_P1_U5719, new_P1_U5720, new_P1_U5721,
    new_P1_U5722, new_P1_U5723, new_P1_U5724, new_P1_U5725, new_P1_U5726,
    new_P1_U5727, new_P1_U5728, new_P1_U5729, new_P1_U5730, new_P1_U5731,
    new_P1_U5732, new_P1_U5733, new_P1_U5734, new_P1_U5735, new_P1_U5736,
    new_P1_U5737, new_P1_U5738, new_P1_U5739, new_P1_U5740, new_P1_U5741,
    new_P1_U5742, new_P1_U5743, new_P1_U5744, new_P1_U5745, new_P1_U5746,
    new_P1_U5747, new_P1_U5748, new_P1_U5749, new_P1_U5750, new_P1_U5751,
    new_P1_U5752, new_P1_U5753, new_P1_U5754, new_P1_U5755, new_P1_U5756,
    new_P1_U5757, new_P1_U5758, new_P1_U5759, new_P1_U5760, new_P1_U5761,
    new_P1_U5762, new_P1_U5763, new_P1_U5764, new_P1_U5765, new_P1_U5766,
    new_P1_U5767, new_P1_U5768, new_P1_U5769, new_P1_U5770, new_P1_U5771,
    new_P1_U5772, new_P1_U5773, new_P1_U5774, new_P1_U5775, new_P1_U5776,
    new_P1_U5777, new_P1_U5778, new_P1_U5779, new_P1_U5780, new_P1_U5781,
    new_P1_U5782, new_P1_U5783, new_P1_U5784, new_P1_U5785, new_P1_U5786,
    new_P1_U5787, new_P1_U5788, new_P1_U5789, new_P1_U5790, new_P1_U5791,
    new_P1_U5792, new_P1_U5793, new_P1_U5794, new_P1_U5795, new_P1_U5796,
    new_P1_U5797, new_P1_U5798, new_P1_U5799, new_P1_U5800, new_P1_U5801,
    new_P1_U5802, new_P1_U5803, new_P1_U5804, new_P1_U5805, new_P1_U5806,
    new_P1_U5807, new_P1_U5808, new_P1_U5809, new_P1_U5810, new_P1_U5811,
    new_P1_U5812, new_P1_U5813, new_P1_U5814, new_P1_U5815, new_P1_U5816,
    new_P1_U5817, new_P1_U5818, new_P1_U5819, new_P1_U5820, new_P1_U5821,
    new_P1_U5822, new_P1_U5823, new_P1_U5824, new_P1_U5825, new_P1_U5826,
    new_P1_U5827, new_P1_U5828, new_P1_U5829, new_P1_U5830, new_P1_U5831,
    new_P1_U5832, new_P1_U5833, new_P1_U5834, new_P1_U5835, new_P1_U5836,
    new_P1_U5837, new_P1_U5838, new_P1_U5839, new_P1_U5840, new_P1_U5841,
    new_P1_U5842, new_P1_U5843, new_P1_U5844, new_P1_U5845, new_P1_U5846,
    new_P1_U5847, new_P1_U5848, new_P1_U5849, new_P1_U5850, new_P1_U5851,
    new_P1_U5852, new_P1_U5853, new_P1_U5854, new_P1_U5855, new_P1_U5856,
    new_P1_U5857, new_P1_U5858, new_P1_U5859, new_P1_U5860, new_P1_U5861,
    new_P1_U5862, new_P1_U5863, new_P1_U5864, new_P1_U5865, new_P1_U5866,
    new_P1_U5867, new_P1_U5868, new_P1_U5869, new_P1_U5870, new_P1_U5871,
    new_P1_U5872, new_P1_U5873, new_P1_U5874, new_P1_U5875, new_P1_U5876,
    new_P1_U5877, new_P1_U5878, new_P1_U5879, new_P1_U5880, new_P1_U5881,
    new_P1_U5882, new_P1_U5883, new_P1_U5884, new_P1_U5885, new_P1_U5886,
    new_P1_U5887, new_P1_U5888, new_P1_U5889, new_P1_U5890, new_P1_U5891,
    new_P1_U5892, new_P1_U5893, new_P1_U5894, new_P1_U5895, new_P1_U5896,
    new_P1_U5897, new_P1_U5898, new_P1_U5899, new_P1_U5900, new_P1_U5901,
    new_P1_U5902, new_P1_U5903, new_P1_U5904, new_P1_U5905, new_P1_U5906,
    new_P1_U5907, new_P1_U5908, new_P1_U5909, new_P1_U5910, new_P1_U5911,
    new_P1_U5912, new_P1_U5913, new_P1_U5914, new_P1_U5915, new_P1_U5916,
    new_P1_U5917, new_P1_U5918, new_P1_U5919, new_P1_U5920, new_P1_U5921,
    new_P1_U5922, new_P1_U5923, new_P1_U5924, new_P1_U5925, new_P1_U5926,
    new_P1_U5927, new_P1_U5928, new_P1_U5929, new_P1_U5930, new_P1_U5931,
    new_P1_U5932, new_P1_U5933, new_P1_U5934, new_P1_U5935, new_P1_U5936,
    new_P1_U5937, new_P1_U5938, new_P1_U5939, new_P1_U5940, new_P1_U5941,
    new_P1_U5942, new_P1_U5943, new_P1_U5944, new_P1_U5945, new_P1_U5946,
    new_P1_U5947, new_P1_U5948, new_P1_U5949, new_P1_U5950, new_P1_U5951,
    new_P1_U5952, new_P1_U5953, new_P1_U5954, new_P1_U5955, new_P1_U5956,
    new_P1_U5957, new_P1_U5958, new_P1_U5959, new_P1_U5960, new_P1_U5961,
    new_P1_U5962, new_P1_U5963, new_P1_U5964, new_P1_U5965, new_P1_U5966,
    new_P1_U5967, new_P1_U5968, new_P1_U5969, new_P1_U5970, new_P1_U5971,
    new_P1_U5972, new_P1_U5973, new_P1_U5974, new_P1_U5975, new_P1_U5976,
    new_P1_U5977, new_P1_U5978, new_P1_U5979, new_P1_U5980, new_P1_U5981,
    new_P1_U5982, new_P1_U5983, new_P1_U5984, new_P1_U5985, new_P1_U5986,
    new_P1_U5987, new_P1_U5988, new_P1_U5989, new_P1_U5990, new_P1_U5991,
    new_P1_U5992, new_P1_U5993, new_P1_U5994, new_P1_U5995, new_P1_U5996,
    new_P1_U5997, new_P1_U5998, new_P1_U5999, new_P1_U6000, new_P1_U6001,
    new_P1_U6002, new_P1_U6003, new_P1_U6004, new_P1_U6005, new_P1_U6006,
    new_P1_U6007, new_P1_U6008, new_P1_U6009, new_P1_U6010, new_P1_U6011,
    new_P1_U6012, new_P1_U6013, new_P1_U6014, new_P1_U6015, new_P1_U6016,
    new_P1_U6017, new_P1_U6018, new_P1_U6019, new_P1_U6020, new_P1_U6021,
    new_P1_U6022, new_P1_U6023, new_P1_U6024, new_P1_U6025, new_P1_U6026,
    new_P1_U6027, new_P1_U6028, new_P1_U6029, new_P1_U6030, new_P1_U6031,
    new_P1_U6032, new_P1_U6033, new_P1_U6034, new_P1_U6035, new_P1_U6036,
    new_P1_U6037, new_P1_U6038, new_P1_U6039, new_P1_U6040, new_P1_U6041,
    new_P1_U6042, new_P1_U6043, new_P1_U6044, new_P1_U6045, new_P1_U6046,
    new_P1_U6047, new_P1_U6048, new_P1_U6049, new_P1_U6050, new_P1_U6051,
    new_P1_U6052, new_P1_U6053, new_P1_U6054, new_P1_U6055, new_P1_U6056,
    new_P1_U6057, new_P1_U6058, new_P1_U6059, new_P1_U6060, new_P1_U6061,
    new_P1_U6062, new_P1_U6063, new_P1_U6064, new_P1_U6065, new_P1_U6066,
    new_P1_U6067, new_P1_U6068, new_P1_U6069, new_P1_U6070, new_P1_U6071,
    new_P1_U6072, new_P1_U6073, new_P1_U6074, new_P1_U6075, new_P1_U6076,
    new_P1_U6077, new_P1_U6078, new_P1_U6079, new_P1_U6080, new_P1_U6081,
    new_P1_U6082, new_P1_U6083, new_P1_U6084, new_P1_U6085, new_P1_U6086,
    new_P1_U6087, new_P1_U6088, new_P1_U6089, new_P1_U6090, new_P1_U6091,
    new_P1_U6092, new_P1_U6093, new_P1_U6094, new_P1_U6095, new_P1_U6096,
    new_P1_U6097, new_P1_U6098, new_P1_U6099, new_P1_U6100, new_P1_U6101,
    new_P1_U6102, new_P1_U6103, new_P1_U6104, new_P1_U6105, new_P1_U6106,
    new_P1_U6107, new_P1_U6108, new_P1_U6109, new_P1_U6110, new_P1_U6111,
    new_P1_U6112, new_P1_U6113, new_P1_U6114, new_P1_U6115, new_P1_U6116,
    new_P1_U6117, new_P1_U6118, new_P1_U6119, new_P1_U6120, new_P1_U6121,
    new_P1_U6122, new_P1_U6123, new_P1_U6124, new_P1_U6125, new_P1_U6126,
    new_P1_U6127, new_P1_U6128, new_P1_U6129, new_P1_U6130, new_P1_U6131,
    new_P1_U6132, new_P1_U6133, new_P1_U6134, new_P1_U6135, new_P1_U6136,
    new_P1_U6137, new_P1_U6138, new_P1_U6139, new_P1_U6140, new_P1_U6141,
    new_P1_U6142, new_P1_U6143, new_P1_U6144, new_P1_U6145, new_P1_U6146,
    new_P1_U6147, new_P1_U6148, new_P1_U6149, new_P1_U6150, new_P1_U6151,
    new_P1_U6152, new_P1_U6153, new_P1_U6154, new_P1_U6155, new_P1_U6156,
    new_P1_U6157, new_P1_U6158, new_P1_U6159, new_P1_U6160, new_P1_U6161,
    new_P1_U6162, new_P1_U6163, new_P1_U6164, new_P1_U6165, new_P1_U6166,
    new_P1_U6167, new_P1_U6168, new_P1_U6169, new_P1_U6170, new_P1_U6171,
    new_P1_U6172, new_P1_U6173, new_P1_U6174, new_P1_U6175, new_P1_U6176,
    new_P1_U6177, new_P1_U6178, new_P1_U6179, new_P1_U6180, new_P1_U6181,
    new_P1_U6182, new_P1_U6183, new_P1_U6184, new_P1_U6185, new_P1_U6186,
    new_P1_U6187, new_P1_U6188, new_P1_U6189, new_P1_U6190, new_P1_U6191,
    new_P1_U6192, new_P1_U6193, new_P1_U6194, new_P1_U6195, new_P1_U6196,
    new_P1_U6197, new_P1_U6198, new_P1_U6199, new_P1_U6200, new_P1_U6201,
    new_P1_U6202, new_P1_U6203, new_P1_U6204, new_P1_U6205, new_P1_U6206,
    new_P1_U6207, new_P1_U6208, new_P1_U6209, new_P1_U6210, new_P1_U6211,
    new_P1_U6212, new_P1_U6213, new_P1_U6214, new_P1_U6215, new_P1_U6216,
    new_P1_U6217, new_P1_U6218, new_P1_U6219, new_P1_U6220, new_P1_U6221,
    new_P1_U6222, new_P1_U6223, new_P1_U6224, new_P1_U6225, new_P1_U6226,
    new_P1_U6227, new_P1_U6228, new_P1_U6229, new_P1_U6230, new_P1_U6231,
    new_P1_U6232, new_P1_U6233, new_P1_U6234, new_P1_U6235, new_P1_U6236,
    new_P1_U6237, new_P1_U6238, new_P1_U6239, new_P1_U6240, new_P1_U6241,
    new_P1_U6242, new_P1_U6243, new_P1_U6244, new_P1_U6245, new_P1_U6246,
    new_P1_U6247, new_P1_U6248, new_P1_U6249, new_P1_U6250, new_P1_U6251,
    new_P1_U6252, new_P1_U6253, new_P1_U6254, new_P1_U6255, new_P1_U6256,
    new_P1_U6257, new_P1_U6258, new_P1_U6259, new_P1_U6260, new_P1_U6261,
    new_P1_U6262, new_P1_U6263, new_P1_U6264, new_P1_U6265, new_P1_U6266,
    new_P1_U6267, new_P1_U6268, new_P1_U6269, new_P1_U6270, new_P1_U6271,
    new_P1_U6272, new_P1_U6273, new_P1_U6274, new_P1_U6275, new_P1_U6276,
    new_P1_U6277, new_P1_U6278, new_P1_U6279, new_P1_U6280, new_P1_U6281,
    new_P1_U6282, new_P1_U6283, new_P1_U6284, new_P1_U6285, new_P1_U6286,
    new_P1_U6287, new_P1_U6288, new_P1_U6289, new_P1_U6290, new_P1_U6291,
    new_P1_U6292, new_P1_U6293, new_P1_U6294, new_P1_U6295, new_P1_U6296,
    new_P1_U6297, new_P1_U6298, new_P1_U6299, new_P1_U6300, new_P1_U6301,
    new_P1_U6302, new_P1_U6303, new_P1_U6304, new_P1_U6305, new_P1_U6306,
    new_P1_U6307, new_P1_U6308, new_P1_U6309, new_P1_U6310, new_P1_U6311,
    new_P1_U6312, new_P1_U6313, new_P1_U6314, new_P1_U6315, new_P1_U6316,
    new_P1_U6317, new_P1_U6318, new_P1_U6319, new_P1_U6320, new_P1_U6321,
    new_P1_U6322, new_P1_U6323, new_P1_U6324, new_P1_U6325, new_P1_U6326,
    new_P1_U6327, new_P1_U6328, new_P1_U6329, new_P1_U6330, new_P1_U6331,
    new_P1_U6332, new_P1_U6333, new_P1_U6334, new_P1_U6335, new_P1_U6336,
    new_P1_U6337, new_P1_U6338, new_P1_U6339, new_P1_U6340, new_P1_U6341,
    new_P1_U6342, new_P1_U6343, new_P1_U6344, new_P1_U6345, new_P1_U6346,
    new_P1_U6347, new_P1_U6348, new_P1_U6349, new_P1_U6350, new_P1_U6351,
    new_P1_U6352, new_P1_U6353, new_P1_U6354, new_P1_U6355, new_P1_U6356,
    new_P1_U6357, new_P1_U6358, new_P1_U6359, new_P1_U6360, new_P1_U6361,
    new_P1_U6362, new_P1_U6363, new_P1_U6364, new_P1_U6365, new_P1_U6366,
    new_P1_U6367, new_P1_U6368, new_P1_U6369, new_P1_U6370, new_P1_U6371,
    new_P1_U6372, new_P1_U6373, new_P1_U6374, new_P1_U6375, new_P1_U6376,
    new_P1_U6377, new_P1_U6378, new_P1_U6379, new_P1_U6380, new_P1_U6381,
    new_P1_U6382, new_P1_U6383, new_P1_U6384, new_P1_U6385, new_P1_U6386,
    new_P1_U6387, new_P1_U6388, new_P1_U6389, new_P1_U6390, new_P1_U6391,
    new_P1_U6392, new_P1_U6393, new_P1_U6394, new_P1_U6395, new_P1_U6396,
    new_P1_U6397, new_P1_U6398, new_P1_U6399, new_P1_U6400, new_P1_U6401,
    new_P1_U6402, new_P1_U6403, new_P1_U6404, new_P1_U6405, new_P1_U6406,
    new_P1_U6407, new_P1_U6408, new_P1_U6409, new_P1_U6410, new_P1_U6411,
    new_P1_U6412, new_P1_U6413, new_P1_U6414, new_P1_U6415, new_P1_U6416,
    new_P1_U6417, new_P1_U6418, new_P1_U6419, new_P1_U6420, new_P1_U6421,
    new_P1_U6422, new_P1_U6423, new_P1_U6424, new_P1_U6425, new_P1_U6426,
    new_P1_U6427, new_P1_U6428, new_P1_U6429, new_P1_U6430, new_P1_U6431,
    new_P1_U6432, new_P1_U6433, new_P1_U6434, new_P1_U6435, new_P1_U6436,
    new_P1_U6437, new_P1_U6438, new_P1_U6439, new_P1_U6440, new_P1_U6441,
    new_P1_U6442, new_P1_U6443, new_P1_U6444, new_P1_U6445, new_P1_U6446,
    new_P1_U6447, new_P1_U6448, new_P1_U6449, new_P1_U6450, new_P1_U6451,
    new_P1_U6452, new_P1_U6453, new_P1_U6454, new_P1_U6455, new_P1_U6456,
    new_P1_U6457, new_P1_U6458, new_P1_U6459, new_P1_U6460, new_P1_U6461,
    new_P1_U6462, new_P1_U6463, new_P1_U6464, new_P1_U6465, new_P1_U6466,
    new_P1_U6467, new_P1_U6468, new_P1_U6469, new_P1_U6470, new_P1_U6471,
    new_P1_U6472, new_P1_U6473, new_P1_U6474, new_P1_U6475, new_P1_U6476,
    new_P1_U6477, new_P1_U6478, new_P1_U6479, new_P1_U6480, new_P1_U6481,
    new_P1_U6482, new_P1_U6483, new_P1_U6484, new_P1_U6485, new_P1_U6486,
    new_P1_U6487, new_P1_U6488, new_P1_U6489, new_P1_U6490, new_P1_U6491,
    new_P1_U6492, new_P1_U6493, new_P1_U6494, new_P1_U6495, new_P1_U6496,
    new_P1_U6497, new_P1_U6498, new_P1_U6499, new_P1_U6500, new_P1_U6501,
    new_P1_U6502, new_P1_U6503, new_P1_U6504, new_P1_U6505, new_P1_U6506,
    new_P1_U6507, new_P1_U6508, new_P1_U6509, new_P1_U6510, new_P1_U6511,
    new_P1_U6512, new_P1_U6513, new_P1_U6514, new_P1_U6515, new_P1_U6516,
    new_P1_U6517, new_P1_U6518, new_P1_U6519, new_P1_U6520, new_P1_U6521,
    new_P1_U6522, new_P1_U6523, new_P1_U6524, new_P1_U6525, new_P1_U6526,
    new_P1_U6527, new_P1_U6528, new_P1_U6529, new_P1_U6530, new_P1_U6531,
    new_P1_U6532, new_P1_U6533, new_P1_U6534, new_P1_U6535, new_P1_U6536,
    new_P1_U6537, new_P1_U6538, new_P1_U6539, new_P1_U6540, new_P1_U6541,
    new_P1_U6542, new_P1_U6543, new_P1_U6544, new_P1_U6545, new_P1_U6546,
    new_P1_U6547, new_P1_U6548, new_P1_U6549, new_P1_U6550, new_P1_U6551,
    new_P1_U6552, new_P1_U6553, new_P1_U6554, new_P1_U6555, new_P1_U6556,
    new_P1_U6557, new_P1_U6558, new_P1_U6559, new_P1_U6560, new_P1_U6561,
    new_P1_U6562, new_P1_U6563, new_P1_U6564, new_P1_U6565, new_P1_U6566,
    new_P1_U6567, new_P1_U6568, new_P1_U6569, new_P1_U6570, new_P1_U6571,
    new_P1_U6572, new_P1_U6573, new_P1_U6574, new_P1_U6575, new_P1_U6576,
    new_P1_U6577, new_P1_U6578, new_P1_U6579, new_P1_U6580, new_P1_U6581,
    new_P1_U6582, new_P1_U6583, new_P1_U6584, new_P1_U6585, new_P1_U6586,
    new_P1_U6587, new_P1_U6588, new_P1_U6589, new_P1_U6590, new_P1_U6591,
    new_P1_U6592, new_P1_U6593, new_P1_U6594, new_P1_U6595, new_P1_U6596,
    new_P1_U6597, new_P1_U6598, new_P1_U6599, new_P1_U6600, new_P1_U6601,
    new_P1_U6602, new_P1_U6603, new_P1_U6604, new_P1_U6605, new_P1_U6606,
    new_P1_U6607, new_P1_U6608, new_P1_U6609, new_P1_U6610, new_P1_U6611,
    new_P1_U6612, new_P1_U6613, new_P1_U6614, new_P1_U6615, new_P1_U6616,
    new_P1_U6617, new_P1_U6618, new_P1_U6619, new_P1_U6620, new_P1_U6621,
    new_P1_U6622, new_P1_U6623, new_P1_U6624, new_P1_U6625, new_P1_U6626,
    new_P1_U6627, new_P1_U6628, new_P1_U6629, new_P1_U6630, new_P1_U6631,
    new_P1_U6632, new_P1_U6633, new_P1_U6634, new_P1_U6635, new_P1_U6636,
    new_P1_U6637, new_P1_U6638, new_P1_U6639, new_P1_U6640, new_P1_U6641,
    new_P1_U6642, new_P1_U6643, new_P1_U6644, new_P1_U6645, new_P1_U6646,
    new_P1_U6647, new_P1_U6648, new_P1_U6649, new_P1_U6650, new_P1_U6651,
    new_P1_U6652, new_P1_U6653, new_P1_U6654, new_P1_U6655, new_P1_U6656,
    new_P1_U6657, new_P1_U6658, new_P1_U6659, new_P1_U6660, new_P1_U6661,
    new_P1_U6662, new_P1_U6663, new_P1_U6664, new_P1_U6665, new_P1_U6666,
    new_P1_U6667, new_P1_U6668, new_P1_U6669, new_P1_U6670, new_P1_U6671,
    new_P1_U6672, new_P1_U6673, new_P1_U6674, new_P1_U6675, new_P1_U6676,
    new_P1_U6677, new_P1_U6678, new_P1_U6679, new_P1_U6680, new_P1_U6681,
    new_P1_U6682, new_P1_U6683, new_P1_U6684, new_P1_U6685, new_P1_U6686,
    new_P1_U6687, new_P1_U6688, new_P1_U6689, new_P1_U6690, new_P1_U6691,
    new_P1_U6692, new_P1_U6693, new_P1_U6694, new_P1_U6695, new_P1_U6696,
    new_P1_U6697, new_P1_U6698, new_P1_U6699, new_P1_U6700, new_P1_U6701,
    new_P1_U6702, new_P1_U6703, new_P1_U6704, new_P1_U6705, new_P1_U6706,
    new_P1_U6707, new_P1_U6708, new_P1_U6709, new_P1_U6710, new_P1_U6711,
    new_P1_U6712, new_P1_U6713, new_P1_U6714, new_P1_U6715, new_P1_U6716,
    new_P1_U6717, new_P1_U6718, new_P1_U6719, new_P1_U6720, new_P1_U6721,
    new_P1_U6722, new_P1_U6723, new_P1_U6724, new_P1_U6725, new_P1_U6726,
    new_P1_U6727, new_P1_U6728, new_P1_U6729, new_P1_U6730, new_P1_U6731,
    new_P1_U6732, new_P1_U6733, new_P1_U6734, new_P1_U6735, new_P1_U6736,
    new_P1_U6737, new_P1_U6738, new_P1_U6739, new_P1_U6740, new_P1_U6741,
    new_P1_U6742, new_P1_U6743, new_P1_U6744, new_P1_U6745, new_P1_U6746,
    new_P1_U6747, new_P1_U6748, new_P1_U6749, new_P1_U6750, new_P1_U6751,
    new_P1_U6752, new_P1_U6753, new_P1_U6754, new_P1_U6755, new_P1_U6756,
    new_P1_U6757, new_P1_U6758, new_P1_U6759, new_P1_U6760, new_P1_U6761,
    new_P1_U6762, new_P1_U6763, new_P1_U6764, new_P1_U6765, new_P1_U6766,
    new_P1_U6767, new_P1_U6768, new_P1_U6769, new_P1_U6770, new_P1_U6771,
    new_P1_U6772, new_P1_U6773, new_P1_U6774, new_P1_U6775, new_P1_U6776,
    new_P1_U6777, new_P1_U6778, new_P1_U6779, new_P1_U6780, new_P1_U6781,
    new_P1_U6782, new_P1_U6783, new_P1_U6784, new_P1_U6785, new_P1_U6786,
    new_P1_U6787, new_P1_U6788, new_P1_U6789, new_P1_U6790, new_P1_U6791,
    new_P1_U6792, new_P1_U6793, new_P1_U6794, new_P1_U6795, new_P1_U6796,
    new_P1_U6797, new_P1_U6798, new_P1_U6799, new_P1_U6800, new_P1_U6801,
    new_P1_U6802, new_P1_U6803, new_P1_U6804, new_P1_U6805, new_P1_U6806,
    new_P1_U6807, new_P1_U6808, new_P1_U6809, new_P1_U6810, new_P1_U6811,
    new_P1_U6812, new_P1_U6813, new_P1_U6814, new_P1_U6815, new_P1_U6816,
    new_P1_U6817, new_P1_U6818, new_P1_U6819, new_P1_U6820, new_P1_U6821,
    new_P1_U6822, new_P1_U6823, new_P1_U6824, new_P1_U6825, new_P1_U6826,
    new_P1_U6827, new_P1_U6828, new_P1_U6829, new_P1_U6830, new_P1_U6831,
    new_P1_U6832, new_P1_U6833, new_P1_U6834, new_P1_U6835, new_P1_U6836,
    new_P1_U6837, new_P1_U6838, new_P1_U6839, new_P1_U6840, new_P1_U6841,
    new_P1_U6842, new_P1_U6843, new_P1_U6844, new_P1_U6845, new_P1_U6846,
    new_P1_U6847, new_P1_U6848, new_P1_U6849, new_P1_U6850, new_P1_U6851,
    new_P1_U6852, new_P1_U6853, new_P1_U6854, new_P1_U6855, new_P1_U6856,
    new_P1_U6857, new_P1_U6858, new_P1_U6859, new_P1_U6860, new_P1_U6861,
    new_P1_U6862, new_P1_U6863, new_P1_U6864, new_P1_U6865, new_P1_U6866,
    new_P1_U6867, new_P1_U6868, new_P1_U6869, new_P1_U6870, new_P1_U6871,
    new_P1_U6872, new_P1_U6873, new_P1_U6874, new_P1_U6875, new_P1_U6876,
    new_P1_U6877, new_P1_U6878, new_P1_U6879, new_P1_U6880, new_P1_U6881,
    new_P1_U6882, new_P1_U6883, new_P1_U6884, new_P1_U6885, new_P1_U6886,
    new_P1_U6887, new_P1_U6888, new_P1_U6889, new_P1_U6890, new_P1_U6891,
    new_P1_U6892, new_P1_U6893, new_P1_U6894, new_P1_U6895, new_P1_U6896,
    new_P1_U6897, new_P1_U6898, new_P1_U6899, new_P1_U6900, new_P1_U6901,
    new_P1_U6902, new_P1_U6903, new_P1_U6904, new_P1_U6905, new_P1_U6906,
    new_P1_U6907, new_P1_U6908, new_P1_U6909, new_P1_U6910, new_P1_U6911,
    new_P1_U6912, new_P1_U6913, new_P1_U6914, new_P1_U6915, new_P1_U6916,
    new_P1_U6917, new_P1_U6918, new_P1_U6919, new_P1_U6920, new_P1_U6921,
    new_P1_U6922, new_P1_U6923, new_P1_U6924, new_P1_U6925, new_P1_U6926,
    new_P1_U6927, new_P1_U6928, new_P1_U6929, new_P1_U6930, new_P1_U6931,
    new_P1_U6932, new_P1_U6933, new_P1_U6934, new_P1_U6935, new_P1_U6936,
    new_P1_U6937, new_P1_U6938, new_P1_U6939, new_P1_U6940, new_P1_U6941,
    new_P1_U6942, new_P1_U6943, new_P1_U6944, new_P1_U6945, new_P1_U6946,
    new_P1_U6947, new_P1_U6948, new_P1_U6949, new_P1_U6950, new_P1_U6951,
    new_P1_U6952, new_P1_U6953, new_P1_U6954, new_P1_U6955, new_P1_U6956,
    new_P1_U6957, new_P1_U6958, new_P1_U6959, new_P1_U6960, new_P1_U6961,
    new_P1_U6962, new_P1_U6963, new_P1_U6964, new_P1_U6965, new_P1_U6966,
    new_P1_U6967, new_P1_U6968, new_P1_U6969, new_P1_U6970, new_P1_U6971,
    new_P1_U6972, new_P1_U6973, new_P1_U6974, new_P1_U6975, new_P1_U6976,
    new_P1_U6977, new_P1_U6978, new_P1_U6979, new_P1_U6980, new_P1_U6981,
    new_P1_U6982, new_P1_U6983, new_P1_U6984, new_P1_U6985, new_P1_U6986,
    new_P1_U6987, new_P1_U6988, new_P1_U6989, new_P1_U6990, new_P1_U6991,
    new_P1_U6992, new_P1_U6993, new_P1_U6994, new_P1_U6995, new_P1_U6996,
    new_P1_U6997, new_P1_U6998, new_P1_U6999, new_P1_U7000, new_P1_U7001,
    new_P1_U7002, new_P1_U7003, new_P1_U7004, new_P1_U7005, new_P1_U7006,
    new_P1_U7007, new_P1_U7008, new_P1_U7009, new_P1_U7010, new_P1_U7011,
    new_P1_U7012, new_P1_U7013, new_P1_U7014, new_P1_U7015, new_P1_U7016,
    new_P1_U7017, new_P1_U7018, new_P1_U7019, new_P1_U7020, new_P1_U7021,
    new_P1_U7022, new_P1_U7023, new_P1_U7024, new_P1_U7025, new_P1_U7026,
    new_P1_U7027, new_P1_U7028, new_P1_U7029, new_P1_U7030, new_P1_U7031,
    new_P1_U7032, new_P1_U7033, new_P1_U7034, new_P1_U7035, new_P1_U7036,
    new_P1_U7037, new_P1_U7038, new_P1_U7039, new_P1_U7040, new_P1_U7041,
    new_P1_U7042, new_P1_U7043, new_P1_U7044, new_P1_U7045, new_P1_U7046,
    new_P1_U7047, new_P1_U7048, new_P1_U7049, new_P1_U7050, new_P1_U7051,
    new_P1_U7052, new_P1_U7053, new_P1_U7054, new_P1_U7055, new_P1_U7056,
    new_P1_U7057, new_P1_U7058, new_P1_U7059, new_P1_U7060, new_P1_U7061,
    new_P1_U7062, new_P1_U7063, new_P1_U7064, new_P1_U7065, new_P1_U7066,
    new_P1_U7067, new_P1_U7068, new_P1_U7069, new_P1_U7070, new_P1_U7071,
    new_P1_U7072, new_P1_U7073, new_P1_U7074, new_P1_U7075, new_P1_U7076,
    new_P1_U7077, new_P1_U7078, new_P1_U7079, new_P1_U7080, new_P1_U7081,
    new_P1_U7082, new_P1_U7083, new_P1_U7084, new_P1_U7085, new_P1_U7086,
    new_P1_U7087, new_P1_U7088, new_P1_U7089, new_P1_U7090, new_P1_U7091,
    new_P1_U7092, new_P1_U7093, new_P1_U7094, new_P1_U7095, new_P1_U7096,
    new_P1_U7097, new_P1_U7098, new_P1_U7099, new_P1_U7100, new_P1_U7101,
    new_P1_U7102, new_P1_U7103, new_P1_U7104, new_P1_U7105, new_P1_U7106,
    new_P1_U7107, new_P1_U7108, new_P1_U7109, new_P1_U7110, new_P1_U7111,
    new_P1_U7112, new_P1_U7113, new_P1_U7114, new_P1_U7115, new_P1_U7116,
    new_P1_U7117, new_P1_U7118, new_P1_U7119, new_P1_U7120, new_P1_U7121,
    new_P1_U7122, new_P1_U7123, new_P1_U7124, new_P1_U7125, new_P1_U7126,
    new_P1_U7127, new_P1_U7128, new_P1_U7129, new_P1_U7130, new_P1_U7131,
    new_P1_U7132, new_P1_U7133, new_P1_U7134, new_P1_U7135, new_P1_U7136,
    new_P1_U7137, new_P1_U7138, new_P1_U7139, new_P1_U7140, new_P1_U7141,
    new_P1_U7142, new_P1_U7143, new_P1_U7144, new_P1_U7145, new_P1_U7146,
    new_P1_U7147, new_P1_U7148, new_P1_U7149, new_P1_U7150, new_P1_U7151,
    new_P1_U7152, new_P1_U7153, new_P1_U7154, new_P1_U7155, new_P1_U7156,
    new_P1_U7157, new_P1_U7158, new_P1_U7159, new_P1_U7160, new_P1_U7161,
    new_P1_U7162, new_P1_U7163, new_P1_U7164, new_P1_U7165, new_P1_U7166,
    new_P1_U7167, new_P1_U7168, new_P1_U7169, new_P1_U7170, new_P1_U7171,
    new_P1_U7172, new_P1_U7173, new_P1_U7174, new_P1_U7175, new_P1_U7176,
    new_P1_U7177, new_P1_U7178, new_P1_U7179, new_P1_U7180, new_P1_U7181,
    new_P1_U7182, new_P1_U7183, new_P1_U7184, new_P1_U7185, new_P1_U7186,
    new_P1_U7187, new_P1_U7188, new_P1_U7189, new_P1_U7190, new_P1_U7191,
    new_P1_U7192, new_P1_U7193, new_P1_U7194, new_P1_U7195, new_P1_U7196,
    new_P1_U7197, new_P1_U7198, new_P1_U7199, new_P1_U7200, new_P1_U7201,
    new_P1_U7202, new_P1_U7203, new_P1_U7204, new_P1_U7205, new_P1_U7206,
    new_P1_U7207, new_P1_U7208, new_P1_U7209, new_P1_U7210, new_P1_U7211,
    new_P1_U7212, new_P1_U7213, new_P1_U7214, new_P1_U7215, new_P1_U7216,
    new_P1_U7217, new_P1_U7218, new_P1_U7219, new_P1_U7220, new_P1_U7221,
    new_P1_U7222, new_P1_U7223, new_P1_U7224, new_P1_U7225, new_P1_U7226,
    new_P1_U7227, new_P1_U7228, new_P1_U7229, new_P1_U7230, new_P1_U7231,
    new_P1_U7232, new_P1_U7233, new_P1_U7234, new_P1_U7235, new_P1_U7236,
    new_P1_U7237, new_P1_U7238, new_P1_U7239, new_P1_U7240, new_P1_U7241,
    new_P1_U7242, new_P1_U7243, new_P1_U7244, new_P1_U7245, new_P1_U7246,
    new_P1_U7247, new_P1_U7248, new_P1_U7249, new_P1_U7250, new_P1_U7251,
    new_P1_U7252, new_P1_U7253, new_P1_U7254, new_P1_U7255, new_P1_U7256,
    new_P1_U7257, new_P1_U7258, new_P1_U7259, new_P1_U7260, new_P1_U7261,
    new_P1_U7262, new_P1_U7263, new_P1_U7264, new_P1_U7265, new_P1_U7266,
    new_P1_U7267, new_P1_U7268, new_P1_U7269, new_P1_U7270, new_P1_U7271,
    new_P1_U7272, new_P1_U7273, new_P1_U7274, new_P1_U7275, new_P1_U7276,
    new_P1_U7277, new_P1_U7278, new_P1_U7279, new_P1_U7280, new_P1_U7281,
    new_P1_U7282, new_P1_U7283, new_P1_U7284, new_P1_U7285, new_P1_U7286,
    new_P1_U7287, new_P1_U7288, new_P1_U7289, new_P1_U7290, new_P1_U7291,
    new_P1_U7292, new_P1_U7293, new_P1_U7294, new_P1_U7295, new_P1_U7296,
    new_P1_U7297, new_P1_U7298, new_P1_U7299, new_P1_U7300, new_P1_U7301,
    new_P1_U7302, new_P1_U7303, new_P1_U7304, new_P1_U7305, new_P1_U7306,
    new_P1_U7307, new_P1_U7308, new_P1_U7309, new_P1_U7310, new_P1_U7311,
    new_P1_U7312, new_P1_U7313, new_P1_U7314, new_P1_U7315, new_P1_U7316,
    new_P1_U7317, new_P1_U7318, new_P1_U7319, new_P1_U7320, new_P1_U7321,
    new_P1_U7322, new_P1_U7323, new_P1_U7324, new_P1_U7325, new_P1_U7326,
    new_P1_U7327, new_P1_U7328, new_P1_U7329, new_P1_U7330, new_P1_U7331,
    new_P1_U7332, new_P1_U7333, new_P1_U7334, new_P1_U7335, new_P1_U7336,
    new_P1_U7337, new_P1_U7338, new_P1_U7339, new_P1_U7340, new_P1_U7341,
    new_P1_U7342, new_P1_U7343, new_P1_U7344, new_P1_U7345, new_P1_U7346,
    new_P1_U7347, new_P1_U7348, new_P1_U7349, new_P1_U7350, new_P1_U7351,
    new_P1_U7352, new_P1_U7353, new_P1_U7354, new_P1_U7355, new_P1_U7356,
    new_P1_U7357, new_P1_U7358, new_P1_U7359, new_P1_U7360, new_P1_U7361,
    new_P1_U7362, new_P1_U7363, new_P1_U7364, new_P1_U7365, new_P1_U7366,
    new_P1_U7367, new_P1_U7368, new_P1_U7369, new_P1_U7370, new_P1_U7371,
    new_P1_U7372, new_P1_U7373, new_P1_U7374, new_P1_U7375, new_P1_U7376,
    new_P1_U7377, new_P1_U7378, new_P1_U7379, new_P1_U7380, new_P1_U7381,
    new_P1_U7382, new_P1_U7383, new_P1_U7384, new_P1_U7385, new_P1_U7386,
    new_P1_U7387, new_P1_U7388, new_P1_U7389, new_P1_U7390, new_P1_U7391,
    new_P1_U7392, new_P1_U7393, new_P1_U7394, new_P1_U7395, new_P1_U7396,
    new_P1_U7397, new_P1_U7398, new_P1_U7399, new_P1_U7400, new_P1_U7401,
    new_P1_U7402, new_P1_U7403, new_P1_U7404, new_P1_U7405, new_P1_U7406,
    new_P1_U7407, new_P1_U7408, new_P1_U7409, new_P1_U7410, new_P1_U7411,
    new_P1_U7412, new_P1_U7413, new_P1_U7414, new_P1_U7415, new_P1_U7416,
    new_P1_U7417, new_P1_U7418, new_P1_U7419, new_P1_U7420, new_P1_U7421,
    new_P1_U7422, new_P1_U7423, new_P1_U7424, new_P1_U7425, new_P1_U7426,
    new_P1_U7427, new_P1_U7428, new_P1_U7429, new_P1_U7430, new_P1_U7431,
    new_P1_U7432, new_P1_U7433, new_P1_U7434, new_P1_U7435, new_P1_U7436,
    new_P1_U7437, new_P1_U7438, new_P1_U7439, new_P1_U7440, new_P1_U7441,
    new_P1_U7442, new_P1_U7443, new_P1_U7444, new_P1_U7445, new_P1_U7446,
    new_P1_U7447, new_P1_U7448, new_P1_U7449, new_P1_U7450, new_P1_U7451,
    new_P1_U7452, new_P1_U7453, new_P1_U7454, new_P1_U7455, new_P1_U7456,
    new_P1_U7457, new_P1_U7458, new_P1_U7459, new_P1_U7460, new_P1_U7461,
    new_P1_U7462, new_P1_U7463, new_P1_U7464, new_P1_U7465, new_P1_U7466,
    new_P1_U7467, new_P1_U7468, new_P1_U7469, new_P1_U7470, new_P1_U7471,
    new_P1_U7472, new_P1_U7473, new_P1_U7474, new_P1_U7475, new_P1_U7476,
    new_P1_U7477, new_P1_U7478, new_P1_U7479, new_P1_U7480, new_P1_U7481,
    new_P1_U7482, new_P1_U7483, new_P1_U7484, new_P1_U7485, new_P1_U7486,
    new_P1_U7487, new_P1_U7488, new_P1_U7489, new_P1_U7490, new_P1_U7491,
    new_P1_U7492, new_P1_U7493, new_P1_U7494, new_P1_U7495, new_P1_U7496,
    new_P1_U7497, new_P1_U7498, new_P1_U7499, new_P1_U7500, new_P1_U7501,
    new_P1_U7502, new_P1_U7503, new_P1_U7504, new_P1_U7505, new_P1_U7506,
    new_P1_U7507, new_P1_U7508, new_P1_U7509, new_P1_U7510, new_P1_U7511,
    new_P1_U7512, new_P1_U7513, new_P1_U7514, new_P1_U7515, new_P1_U7516,
    new_P1_U7517, new_P1_U7518, new_P1_U7519, new_P1_U7520, new_P1_U7521,
    new_P1_U7522, new_P1_U7523, new_P1_U7524, new_P1_U7525, new_P1_U7526,
    new_P1_U7527, new_P1_U7528, new_P1_U7529, new_P1_U7530, new_P1_U7531,
    new_P1_U7532, new_P1_U7533, new_P1_U7534, new_P1_U7535, new_P1_U7536,
    new_P1_U7537, new_P1_U7538, new_P1_U7539, new_P1_U7540, new_P1_U7541,
    new_P1_U7542, new_P1_U7543, new_P1_U7544, new_P1_U7545, new_P1_U7546,
    new_P1_U7547, new_P1_U7548, new_P1_U7549, new_P1_U7550, new_P1_U7551,
    new_P1_U7552, new_P1_U7553, new_P1_U7554, new_P1_U7555, new_P1_U7556,
    new_P1_U7557, new_P1_U7558, new_P1_U7559, new_P1_U7560, new_P1_U7561,
    new_P1_U7562, new_P1_U7563, new_P1_U7564, new_P1_U7565, new_P1_U7566,
    new_P1_U7567, new_P1_U7568, new_P1_U7569, new_P1_U7570, new_P1_U7571,
    new_P1_U7572, new_P1_U7573, new_P1_U7574, new_P1_U7575, new_P1_U7576,
    new_P1_U7577, new_P1_U7578, new_P1_U7579, new_P1_U7580, new_P1_U7581,
    new_P1_U7582, new_P1_U7583, new_P1_U7584, new_P1_U7585, new_P1_U7586,
    new_P1_U7587, new_P1_U7588, new_P1_U7589, new_P1_U7590, new_P1_U7591,
    new_P1_U7592, new_P1_U7593, new_P1_U7594, new_P1_U7595, new_P1_U7596,
    new_P1_U7597, new_P1_U7598, new_P1_U7599, new_P1_U7600, new_P1_U7601,
    new_P1_U7602, new_P1_U7603, new_P1_U7604, new_P1_U7605, new_P1_U7606,
    new_P1_U7607, new_P1_U7608, new_P1_U7609, new_P1_U7610, new_P1_U7611,
    new_P1_U7612, new_P1_U7613, new_P1_U7614, new_P1_U7615, new_P1_U7616,
    new_P1_U7617, new_P1_U7618, new_P1_U7619, new_P1_U7620, new_P1_U7621,
    new_P1_U7622, new_P1_U7623, new_P1_U7624, new_P1_U7625, new_P1_U7626,
    new_P1_U7627, new_P1_U7628, new_P1_U7629, new_P1_U7630, new_P1_U7631,
    new_P1_U7632, new_P1_U7633, new_P1_U7634, new_P1_U7635, new_P1_U7636,
    new_P1_U7637, new_P1_U7638, new_P1_U7639, new_P1_U7640, new_P1_U7641,
    new_P1_U7642, new_P1_U7643, new_P1_U7644, new_P1_U7645, new_P1_U7646,
    new_P1_U7647, new_P1_U7648, new_P1_U7649, new_P1_U7650, new_P1_U7651,
    new_P1_U7652, new_P1_U7653, new_P1_U7654, new_P1_U7655, new_P1_U7656,
    new_P1_U7657, new_P1_U7658, new_P1_U7659, new_P1_U7660, new_P1_U7661,
    new_P1_U7662, new_P1_U7663, new_P1_U7664, new_P1_U7665, new_P1_U7666,
    new_P1_U7667, new_P1_U7668, new_P1_U7669, new_P1_U7670, new_P1_U7671,
    new_P1_U7672, new_P1_U7673, new_P1_U7674, new_P1_U7675, new_P1_U7676,
    new_P1_U7677, new_P1_U7678, new_P1_U7679, new_P1_U7680, new_P1_U7681,
    new_P1_U7682, new_P1_U7683, new_P1_U7684, new_P1_U7685, new_P1_U7686,
    new_P1_U7687, new_P1_U7688, new_P1_U7689, new_P1_U7690, new_P1_U7691,
    new_P1_U7692, new_P1_U7693, new_P1_U7694, new_P1_U7695, new_P1_U7696,
    new_P1_U7697, new_P1_U7698, new_P1_U7699, new_P1_U7700, new_P1_U7701,
    new_P1_U7702, new_P1_U7703, new_P1_U7704, new_P1_U7705, new_P1_U7706,
    new_P1_U7707, new_P1_U7708, new_P1_U7709, new_P1_U7710, new_P1_U7711,
    new_P1_U7712, new_P1_U7713, new_P1_U7714, new_P1_U7715, new_P1_U7716,
    new_P1_U7717, new_P1_U7718, new_P1_U7719, new_P1_U7720, new_P1_U7721,
    new_P1_U7722, new_P1_U7723, new_P1_U7724, new_P1_U7725, new_P1_U7726,
    new_P1_U7727, new_P1_U7728, new_P1_U7729, new_P1_U7730, new_P1_U7731,
    new_P1_U7732, new_P1_U7733, new_P1_U7734, new_P1_U7735, new_P1_U7736,
    new_P1_U7737, new_P1_U7738, new_P1_U7739, new_P1_U7740, new_P1_U7741,
    new_P1_U7742, new_P1_U7743, new_P1_U7744, new_P1_U7745, new_P1_U7746,
    new_P1_U7747, new_P1_U7748, new_P1_U7749, new_P1_U7750, new_P1_U7751,
    new_P1_U7752, new_P1_U7753, new_P1_U7754, new_P1_U7755, new_P1_U7756,
    new_P1_U7757, new_P1_U7758, new_P1_U7759, new_P1_U7760, new_P1_U7761,
    new_P1_U7762, new_P1_U7763, new_P1_U7764, new_P1_U7765, new_P1_U7766,
    new_P1_U7767, new_P1_U7768, new_P1_U7769, new_P1_U7770, new_P1_U7771,
    new_P1_U7772, new_P1_U7773, new_P1_U7774, new_P1_U7775, new_P1_U7776,
    new_P1_U7777, new_P1_U7778, new_P1_U7779, new_P1_U7780, new_P1_U7781,
    new_P1_U7782, new_P1_U7783, new_P1_U7784, new_P1_U7785, new_P1_U7786,
    new_P1_U7787, new_P1_U7788, new_P1_U7789, new_P1_U7790, new_P1_U7791,
    new_P1_U7792, new_P1_U7793, new_P1_U7794, new_P1_ADD_405_U113,
    new_P1_ADD_405_U112, new_P1_ADD_405_U111, new_P1_ADD_405_U110,
    new_P1_ADD_405_U109, new_P1_ADD_405_U108, new_P1_ADD_405_U107,
    new_P1_ADD_405_U106, new_P1_ADD_405_U105, new_P1_ADD_405_U104,
    new_P1_ADD_405_U103, new_P1_ADD_405_U102, new_P1_ADD_405_U101,
    new_P1_ADD_405_U100, new_P1_ADD_405_U99, new_P1_ADD_405_U98,
    new_P1_ADD_405_U97, new_P1_ADD_405_U96, new_P1_ADD_405_U95,
    new_P1_ADD_405_U94, new_P1_ADD_405_U93, new_P1_ADD_405_U92,
    new_P1_ADD_405_U91, new_P1_ADD_405_U90, new_P1_ADD_405_U89,
    new_P1_ADD_405_U88, new_P1_ADD_405_U87, new_LT_782_120_U6,
    new_LT_782_120_U7, new_LT_782_U6, new_LT_782_U7, new_LT_748_U6,
    new_R170_U6, new_R170_U7, new_R170_U8, new_R170_U9, new_R170_U10,
    new_R170_U11, new_R170_U12, new_R170_U13, new_R170_U14, new_R170_U15,
    new_R165_U6, new_R165_U7, new_R165_U8, new_R165_U9, new_R165_U10,
    new_R165_U11, new_R165_U12, new_R165_U13, new_R165_U14, new_R165_U15,
    new_LT_782_119_U6, new_LT_782_119_U7, new_P3_ADD_526_U5,
    new_P3_ADD_526_U6, new_P3_ADD_526_U7, new_P3_ADD_526_U8,
    new_P3_ADD_526_U9, new_P3_ADD_526_U10, new_P3_ADD_526_U11,
    new_P3_ADD_526_U12, new_P3_ADD_526_U13, new_P3_ADD_526_U14,
    new_P3_ADD_526_U15, new_P3_ADD_526_U16, new_P3_ADD_526_U17,
    new_P3_ADD_526_U18, new_P3_ADD_526_U19, new_P3_ADD_526_U20,
    new_P3_ADD_526_U21, new_P3_ADD_526_U22, new_P3_ADD_526_U23,
    new_P3_ADD_526_U24, new_P3_ADD_526_U25, new_P3_ADD_526_U26,
    new_P3_ADD_526_U27, new_P3_ADD_526_U28, new_P3_ADD_526_U29,
    new_P3_ADD_526_U30, new_P3_ADD_526_U31, new_P3_ADD_526_U32,
    new_P3_ADD_526_U33, new_P3_ADD_526_U34, new_P3_ADD_526_U35,
    new_P3_ADD_526_U36, new_P3_ADD_526_U37, new_P3_ADD_526_U38,
    new_P3_ADD_526_U39, new_P3_ADD_526_U40, new_P3_ADD_526_U41,
    new_P3_ADD_526_U42, new_P3_ADD_526_U43, new_P3_ADD_526_U44,
    new_P3_ADD_526_U45, new_P3_ADD_526_U46, new_P3_ADD_526_U47,
    new_P3_ADD_526_U48, new_P3_ADD_526_U49, new_P3_ADD_526_U50,
    new_P3_ADD_526_U51, new_P3_ADD_526_U52, new_P3_ADD_526_U53,
    new_P3_ADD_526_U54, new_P3_ADD_526_U55, new_P3_ADD_526_U56,
    new_P3_ADD_526_U57, new_P3_ADD_526_U58, new_P3_ADD_526_U59,
    new_P3_ADD_526_U60, new_P3_ADD_526_U61, new_P3_ADD_526_U62,
    new_P3_ADD_526_U63, new_P3_ADD_526_U64, new_P3_ADD_526_U65,
    new_P3_ADD_526_U66, new_P3_ADD_526_U67, new_P3_ADD_526_U68,
    new_P3_ADD_526_U69, new_P3_ADD_526_U70, new_P3_ADD_526_U71,
    new_P3_ADD_526_U72, new_P3_ADD_526_U73, new_P3_ADD_526_U74,
    new_P3_ADD_526_U75, new_P3_ADD_526_U76, new_P3_ADD_526_U77,
    new_P3_ADD_526_U78, new_P3_ADD_526_U79, new_P3_ADD_526_U80,
    new_P3_ADD_526_U81, new_P3_ADD_526_U82, new_P3_ADD_526_U83,
    new_P3_ADD_526_U84, new_P3_ADD_526_U85, new_P3_ADD_526_U86,
    new_P3_ADD_526_U87, new_P3_ADD_526_U88, new_P3_ADD_526_U89,
    new_P3_ADD_526_U90, new_P3_ADD_526_U91, new_P3_ADD_526_U92,
    new_P3_ADD_526_U93, new_P3_ADD_526_U94, new_P3_ADD_526_U95,
    new_P3_ADD_526_U96, new_P3_ADD_526_U97, new_P3_ADD_526_U98,
    new_P3_ADD_526_U99, new_P3_ADD_526_U100, new_P3_ADD_526_U101,
    new_P3_ADD_526_U102, new_P3_ADD_526_U103, new_P3_ADD_526_U104,
    new_P3_ADD_526_U105, new_P3_ADD_526_U106, new_P3_ADD_526_U107,
    new_P3_ADD_526_U108, new_P3_ADD_526_U109, new_P3_ADD_526_U110,
    new_P3_ADD_526_U111, new_P3_ADD_526_U112, new_P3_ADD_526_U113,
    new_P3_ADD_526_U114, new_P3_ADD_526_U115, new_P3_ADD_526_U116,
    new_P3_ADD_526_U117, new_P3_ADD_526_U118, new_P3_ADD_526_U119,
    new_P3_ADD_526_U120, new_P3_ADD_526_U121, new_P3_ADD_526_U122,
    new_P3_ADD_526_U123, new_P3_ADD_526_U124, new_P3_ADD_526_U125,
    new_P3_ADD_526_U126, new_P3_ADD_526_U127, new_P3_ADD_526_U128,
    new_P3_ADD_526_U129, new_P3_ADD_526_U130, new_P3_ADD_526_U131,
    new_P3_ADD_526_U132, new_P3_ADD_526_U133, new_P3_ADD_526_U134,
    new_P3_ADD_526_U135, new_P3_ADD_526_U136, new_P3_ADD_526_U137,
    new_P3_ADD_526_U138, new_P3_ADD_526_U139, new_P3_ADD_526_U140,
    new_P3_ADD_526_U141, new_P3_ADD_526_U142, new_P3_ADD_526_U143,
    new_P3_ADD_526_U144, new_P3_ADD_526_U145, new_P3_ADD_526_U146,
    new_P3_ADD_526_U147, new_P3_ADD_526_U148, new_P3_ADD_526_U149,
    new_P3_ADD_526_U150, new_P3_ADD_526_U151, new_P3_ADD_526_U152,
    new_P3_ADD_526_U153, new_P3_ADD_526_U154, new_P3_ADD_526_U155,
    new_P3_ADD_526_U156, new_P3_ADD_526_U157, new_P3_ADD_526_U158,
    new_P3_ADD_526_U159, new_P3_ADD_526_U160, new_P3_ADD_526_U161,
    new_P3_ADD_526_U162, new_P3_ADD_526_U163, new_P3_ADD_526_U164,
    new_P3_ADD_526_U165, new_P3_ADD_526_U166, new_P3_ADD_526_U167,
    new_P3_ADD_526_U168, new_P3_ADD_526_U169, new_P3_ADD_526_U170,
    new_P3_ADD_526_U171, new_P3_ADD_526_U172, new_P3_ADD_526_U173,
    new_P3_ADD_526_U174, new_P3_ADD_526_U175, new_P3_ADD_526_U176,
    new_P3_ADD_526_U177, new_P3_ADD_526_U178, new_P3_ADD_526_U179,
    new_P3_ADD_526_U180, new_P3_ADD_526_U181, new_P3_ADD_526_U182,
    new_P3_ADD_526_U183, new_P3_ADD_526_U184, new_P3_ADD_526_U185,
    new_P3_ADD_526_U186, new_P3_ADD_526_U187, new_P3_ADD_526_U188,
    new_P3_ADD_526_U189, new_P3_ADD_526_U190, new_P3_ADD_526_U191,
    new_P3_ADD_526_U192, new_P3_ADD_526_U193, new_P3_ADD_526_U194,
    new_P3_ADD_526_U195, new_P3_ADD_526_U196, new_P3_ADD_526_U197,
    new_P3_ADD_526_U198, new_P3_ADD_526_U199, new_P3_ADD_526_U200,
    new_P3_ADD_526_U201, new_P3_ADD_526_U202, new_P3_ADD_552_U5,
    new_P3_ADD_552_U6, new_P3_ADD_552_U7, new_P3_ADD_552_U8,
    new_P3_ADD_552_U9, new_P3_ADD_552_U10, new_P3_ADD_552_U11,
    new_P3_ADD_552_U12, new_P3_ADD_552_U13, new_P3_ADD_552_U14,
    new_P3_ADD_552_U15, new_P3_ADD_552_U16, new_P3_ADD_552_U17,
    new_P3_ADD_552_U18, new_P3_ADD_552_U19, new_P3_ADD_552_U20,
    new_P3_ADD_552_U21, new_P3_ADD_552_U22, new_P3_ADD_552_U23,
    new_P3_ADD_552_U24, new_P3_ADD_552_U25, new_P3_ADD_552_U26,
    new_P3_ADD_552_U27, new_P3_ADD_552_U28, new_P3_ADD_552_U29,
    new_P3_ADD_552_U30, new_P3_ADD_552_U31, new_P3_ADD_552_U32,
    new_P3_ADD_552_U33, new_P3_ADD_552_U34, new_P3_ADD_552_U35,
    new_P3_ADD_552_U36, new_P3_ADD_552_U37, new_P3_ADD_552_U38,
    new_P3_ADD_552_U39, new_P3_ADD_552_U40, new_P3_ADD_552_U41,
    new_P3_ADD_552_U42, new_P3_ADD_552_U43, new_P3_ADD_552_U44,
    new_P3_ADD_552_U45, new_P3_ADD_552_U46, new_P3_ADD_552_U47,
    new_P3_ADD_552_U48, new_P3_ADD_552_U49, new_P3_ADD_552_U50,
    new_P3_ADD_552_U51, new_P3_ADD_552_U52, new_P3_ADD_552_U53,
    new_P3_ADD_552_U54, new_P3_ADD_552_U55, new_P3_ADD_552_U56,
    new_P3_ADD_552_U57, new_P3_ADD_552_U58, new_P3_ADD_552_U59,
    new_P3_ADD_552_U60, new_P3_ADD_552_U61, new_P3_ADD_552_U62,
    new_P3_ADD_552_U63, new_P3_ADD_552_U64, new_P3_ADD_552_U65,
    new_P3_ADD_552_U66, new_P3_ADD_552_U67, new_P3_ADD_552_U68,
    new_P3_ADD_552_U69, new_P3_ADD_552_U70, new_P3_ADD_552_U71,
    new_P3_ADD_552_U72, new_P3_ADD_552_U73, new_P3_ADD_552_U74,
    new_P3_ADD_552_U75, new_P3_ADD_552_U76, new_P3_ADD_552_U77,
    new_P3_ADD_552_U78, new_P3_ADD_552_U79, new_P3_ADD_552_U80,
    new_P3_ADD_552_U81, new_P3_ADD_552_U82, new_P3_ADD_552_U83,
    new_P3_ADD_552_U84, new_P3_ADD_552_U85, new_P3_ADD_552_U86,
    new_P3_ADD_552_U87, new_P3_ADD_552_U88, new_P3_ADD_552_U89,
    new_P3_ADD_552_U90, new_P3_ADD_552_U91, new_P3_ADD_552_U92,
    new_P3_ADD_552_U93, new_P3_ADD_552_U94, new_P3_ADD_552_U95,
    new_P3_ADD_552_U96, new_P3_ADD_552_U97, new_P3_ADD_552_U98,
    new_P3_ADD_552_U99, new_P3_ADD_552_U100, new_P3_ADD_552_U101,
    new_P3_ADD_552_U102, new_P3_ADD_552_U103, new_P3_ADD_552_U104,
    new_P3_ADD_552_U105, new_P3_ADD_552_U106, new_P3_ADD_552_U107,
    new_P3_ADD_552_U108, new_P3_ADD_552_U109, new_P3_ADD_552_U110,
    new_P3_ADD_552_U111, new_P3_ADD_552_U112, new_P3_ADD_552_U113,
    new_P3_ADD_552_U114, new_P3_ADD_552_U115, new_P3_ADD_552_U116,
    new_P3_ADD_552_U117, new_P3_ADD_552_U118, new_P3_ADD_552_U119,
    new_P3_ADD_552_U120, new_P3_ADD_552_U121, new_P3_ADD_552_U122,
    new_P3_ADD_552_U123, new_P3_ADD_552_U124, new_P3_ADD_552_U125,
    new_P3_ADD_552_U126, new_P3_ADD_552_U127, new_P3_ADD_552_U128,
    new_P3_ADD_552_U129, new_P3_ADD_552_U130, new_P3_ADD_552_U131,
    new_P3_ADD_552_U132, new_P3_ADD_552_U133, new_P3_ADD_552_U134,
    new_P3_ADD_552_U135, new_P3_ADD_552_U136, new_P3_ADD_552_U137,
    new_P3_ADD_552_U138, new_P3_ADD_552_U139, new_P3_ADD_552_U140,
    new_P3_ADD_552_U141, new_P3_ADD_552_U142, new_P3_ADD_552_U143,
    new_P3_ADD_552_U144, new_P3_ADD_552_U145, new_P3_ADD_552_U146,
    new_P3_ADD_552_U147, new_P3_ADD_552_U148, new_P3_ADD_552_U149,
    new_P3_ADD_552_U150, new_P3_ADD_552_U151, new_P3_ADD_552_U152,
    new_P3_ADD_552_U153, new_P3_ADD_552_U154, new_P3_ADD_552_U155,
    new_P3_ADD_552_U156, new_P3_ADD_552_U157, new_P3_ADD_552_U158,
    new_P3_ADD_552_U159, new_P3_ADD_552_U160, new_P3_ADD_552_U161,
    new_P3_ADD_552_U162, new_P3_ADD_552_U163, new_P3_ADD_552_U164,
    new_P3_ADD_552_U165, new_P3_ADD_552_U166, new_P3_ADD_552_U167,
    new_P3_ADD_552_U168, new_P3_ADD_552_U169, new_P3_ADD_552_U170,
    new_P3_ADD_552_U171, new_P3_ADD_552_U172, new_P3_ADD_552_U173,
    new_P3_ADD_552_U174, new_P3_ADD_552_U175, new_P3_ADD_552_U176,
    new_P3_ADD_552_U177, new_P3_ADD_552_U178, new_P3_ADD_552_U179,
    new_P3_ADD_552_U180, new_P3_ADD_552_U181, new_P3_ADD_552_U182,
    new_P3_ADD_552_U183, new_P3_ADD_552_U184, new_P3_ADD_552_U185,
    new_P3_ADD_552_U186, new_P3_ADD_552_U187, new_P3_ADD_552_U188,
    new_P3_ADD_552_U189, new_P3_ADD_552_U190, new_P3_ADD_552_U191,
    new_P3_ADD_552_U192, new_P3_ADD_552_U193, new_P3_ADD_552_U194,
    new_P3_ADD_552_U195, new_P3_ADD_552_U196, new_P3_ADD_552_U197,
    new_P3_ADD_552_U198, new_P3_ADD_552_U199, new_P3_ADD_552_U200,
    new_P3_ADD_552_U201, new_P3_ADD_552_U202, new_P3_ADD_546_U5,
    new_P3_ADD_546_U6, new_P3_ADD_546_U7, new_P3_ADD_546_U8,
    new_P3_ADD_546_U9, new_P3_ADD_546_U10, new_P3_ADD_546_U11,
    new_P3_ADD_546_U12, new_P3_ADD_546_U13, new_P3_ADD_546_U14,
    new_P3_ADD_546_U15, new_P3_ADD_546_U16, new_P3_ADD_546_U17,
    new_P3_ADD_546_U18, new_P3_ADD_546_U19, new_P3_ADD_546_U20,
    new_P3_ADD_546_U21, new_P3_ADD_546_U22, new_P3_ADD_546_U23,
    new_P3_ADD_546_U24, new_P3_ADD_546_U25, new_P3_ADD_546_U26,
    new_P3_ADD_546_U27, new_P3_ADD_546_U28, new_P3_ADD_546_U29,
    new_P3_ADD_546_U30, new_P3_ADD_546_U31, new_P3_ADD_546_U32,
    new_P3_ADD_546_U33, new_P3_ADD_546_U34, new_P3_ADD_546_U35,
    new_P3_ADD_546_U36, new_P3_ADD_546_U37, new_P3_ADD_546_U38,
    new_P3_ADD_546_U39, new_P3_ADD_546_U40, new_P3_ADD_546_U41,
    new_P3_ADD_546_U42, new_P3_ADD_546_U43, new_P3_ADD_546_U44,
    new_P3_ADD_546_U45, new_P3_ADD_546_U46, new_P3_ADD_546_U47,
    new_P3_ADD_546_U48, new_P3_ADD_546_U49, new_P3_ADD_546_U50,
    new_P3_ADD_546_U51, new_P3_ADD_546_U52, new_P3_ADD_546_U53,
    new_P3_ADD_546_U54, new_P3_ADD_546_U55, new_P3_ADD_546_U56,
    new_P3_ADD_546_U57, new_P3_ADD_546_U58, new_P3_ADD_546_U59,
    new_P3_ADD_546_U60, new_P3_ADD_546_U61, new_P3_ADD_546_U62,
    new_P3_ADD_546_U63, new_P3_ADD_546_U64, new_P3_ADD_546_U65,
    new_P3_ADD_546_U66, new_P3_ADD_546_U67, new_P3_ADD_546_U68,
    new_P3_ADD_546_U69, new_P3_ADD_546_U70, new_P3_ADD_546_U71,
    new_P3_ADD_546_U72, new_P3_ADD_546_U73, new_P3_ADD_546_U74,
    new_P3_ADD_546_U75, new_P3_ADD_546_U76, new_P3_ADD_546_U77,
    new_P3_ADD_546_U78, new_P3_ADD_546_U79, new_P3_ADD_546_U80,
    new_P3_ADD_546_U81, new_P3_ADD_546_U82, new_P3_ADD_546_U83,
    new_P3_ADD_546_U84, new_P3_ADD_546_U85, new_P3_ADD_546_U86,
    new_P3_ADD_546_U87, new_P3_ADD_546_U88, new_P3_ADD_546_U89,
    new_P3_ADD_546_U90, new_P3_ADD_546_U91, new_P3_ADD_546_U92,
    new_P3_ADD_546_U93, new_P3_ADD_546_U94, new_P3_ADD_546_U95,
    new_P3_ADD_546_U96, new_P3_ADD_546_U97, new_P3_ADD_546_U98,
    new_P3_ADD_546_U99, new_P3_ADD_546_U100, new_P3_ADD_546_U101,
    new_P3_ADD_546_U102, new_P3_ADD_546_U103, new_P3_ADD_546_U104,
    new_P3_ADD_546_U105, new_P3_ADD_546_U106, new_P3_ADD_546_U107,
    new_P3_ADD_546_U108, new_P3_ADD_546_U109, new_P3_ADD_546_U110,
    new_P3_ADD_546_U111, new_P3_ADD_546_U112, new_P3_ADD_546_U113,
    new_P3_ADD_546_U114, new_P3_ADD_546_U115, new_P3_ADD_546_U116,
    new_P3_ADD_546_U117, new_P3_ADD_546_U118, new_P3_ADD_546_U119,
    new_P3_ADD_546_U120, new_P3_ADD_546_U121, new_P3_ADD_546_U122,
    new_P3_ADD_546_U123, new_P3_ADD_546_U124, new_P3_ADD_546_U125,
    new_P3_ADD_546_U126, new_P3_ADD_546_U127, new_P3_ADD_546_U128,
    new_P3_ADD_546_U129, new_P3_ADD_546_U130, new_P3_ADD_546_U131,
    new_P3_ADD_546_U132, new_P3_ADD_546_U133, new_P3_ADD_546_U134,
    new_P3_ADD_546_U135, new_P3_ADD_546_U136, new_P3_ADD_546_U137,
    new_P3_ADD_546_U138, new_P3_ADD_546_U139, new_P3_ADD_546_U140,
    new_P3_ADD_546_U141, new_P3_ADD_546_U142, new_P3_ADD_546_U143,
    new_P3_ADD_546_U144, new_P3_ADD_546_U145, new_P3_ADD_546_U146,
    new_P3_ADD_546_U147, new_P3_ADD_546_U148, new_P3_ADD_546_U149,
    new_P3_ADD_546_U150, new_P3_ADD_546_U151, new_P3_ADD_546_U152,
    new_P3_ADD_546_U153, new_P3_ADD_546_U154, new_P3_ADD_546_U155,
    new_P3_ADD_546_U156, new_P3_ADD_546_U157, new_P3_ADD_546_U158,
    new_P3_ADD_546_U159, new_P3_ADD_546_U160, new_P3_ADD_546_U161,
    new_P3_ADD_546_U162, new_P3_ADD_546_U163, new_P3_ADD_546_U164,
    new_P3_ADD_546_U165, new_P3_ADD_546_U166, new_P3_ADD_546_U167,
    new_P3_ADD_546_U168, new_P3_ADD_546_U169, new_P3_ADD_546_U170,
    new_P3_ADD_546_U171, new_P3_ADD_546_U172, new_P3_ADD_546_U173,
    new_P3_ADD_546_U174, new_P3_ADD_546_U175, new_P3_ADD_546_U176,
    new_P3_ADD_546_U177, new_P3_ADD_546_U178, new_P3_ADD_546_U179,
    new_P3_ADD_546_U180, new_P3_ADD_546_U181, new_P3_ADD_546_U182,
    new_P3_ADD_546_U183, new_P3_ADD_546_U184, new_P3_ADD_546_U185,
    new_P3_ADD_546_U186, new_P3_ADD_546_U187, new_P3_ADD_546_U188,
    new_P3_ADD_546_U189, new_P3_ADD_546_U190, new_P3_ADD_546_U191,
    new_P3_ADD_546_U192, new_P3_ADD_546_U193, new_P3_ADD_546_U194,
    new_P3_ADD_546_U195, new_P3_ADD_546_U196, new_P3_ADD_546_U197,
    new_P3_ADD_546_U198, new_P3_ADD_546_U199, new_P3_ADD_546_U200,
    new_P3_ADD_546_U201, new_P3_ADD_546_U202, new_P3_GTE_401_U6,
    new_P3_GTE_401_U7, new_P3_GTE_401_U8, new_P3_GTE_401_U9,
    new_P3_ADD_391_1180_U4, new_P3_ADD_391_1180_U5, new_P3_ADD_391_1180_U6,
    new_P3_ADD_391_1180_U7, new_P3_ADD_391_1180_U8, new_P3_ADD_391_1180_U9,
    new_P3_ADD_391_1180_U10, new_P3_ADD_391_1180_U11,
    new_P3_ADD_391_1180_U12, new_P3_ADD_391_1180_U13,
    new_P3_ADD_391_1180_U14, new_P3_ADD_391_1180_U15,
    new_P3_ADD_391_1180_U16, new_P3_ADD_391_1180_U17,
    new_P3_ADD_391_1180_U18, new_P3_ADD_391_1180_U19,
    new_P3_ADD_391_1180_U20, new_P3_ADD_391_1180_U21,
    new_P3_ADD_391_1180_U22, new_P3_ADD_391_1180_U23,
    new_P3_ADD_391_1180_U24, new_P3_ADD_391_1180_U25,
    new_P3_ADD_391_1180_U26, new_P3_ADD_391_1180_U27,
    new_P3_ADD_391_1180_U28, new_P3_ADD_391_1180_U29,
    new_P3_ADD_391_1180_U30, new_P3_ADD_391_1180_U31,
    new_P3_ADD_391_1180_U32, new_P3_ADD_391_1180_U33,
    new_P3_ADD_391_1180_U34, new_P3_ADD_391_1180_U35,
    new_P3_ADD_391_1180_U36, new_P3_ADD_391_1180_U37,
    new_P3_ADD_391_1180_U38, new_P3_ADD_391_1180_U39,
    new_P3_ADD_391_1180_U40, new_P3_ADD_391_1180_U41,
    new_P3_ADD_391_1180_U42, new_P3_ADD_391_1180_U43,
    new_P3_ADD_391_1180_U44, new_P3_ADD_391_1180_U45,
    new_P3_ADD_391_1180_U46, new_P3_ADD_391_1180_U47,
    new_P3_ADD_391_1180_U48, new_P3_ADD_391_1180_U49,
    new_P3_ADD_391_1180_U50, new_P3_ADD_476_U4, new_P3_ADD_476_U5,
    new_P3_ADD_476_U6, new_P3_ADD_476_U7, new_P3_ADD_476_U8,
    new_P3_ADD_476_U9, new_P3_ADD_476_U10, new_P3_ADD_476_U11,
    new_P3_ADD_476_U12, new_P3_ADD_476_U13, new_P3_ADD_476_U14,
    new_P3_ADD_476_U15, new_P3_ADD_476_U16, new_P3_ADD_476_U17,
    new_P3_ADD_476_U18, new_P3_ADD_476_U19, new_P3_ADD_476_U20,
    new_P3_ADD_476_U21, new_P3_ADD_476_U22, new_P3_ADD_476_U23,
    new_P3_ADD_476_U24, new_P3_ADD_476_U25, new_P3_ADD_476_U26,
    new_P3_ADD_476_U27, new_P3_ADD_476_U28, new_P3_ADD_476_U29,
    new_P3_ADD_476_U30, new_P3_ADD_476_U31, new_P3_ADD_476_U32,
    new_P3_ADD_476_U33, new_P3_ADD_476_U34, new_P3_ADD_476_U35,
    new_P3_ADD_476_U36, new_P3_ADD_476_U37, new_P3_ADD_476_U38,
    new_P3_ADD_476_U39, new_P3_ADD_476_U40, new_P3_ADD_476_U41,
    new_P3_ADD_476_U42, new_P3_ADD_476_U43, new_P3_ADD_476_U44,
    new_P3_ADD_476_U45, new_P3_ADD_476_U46, new_P3_ADD_476_U47,
    new_P3_ADD_476_U48, new_P3_ADD_476_U49, new_P3_ADD_476_U50,
    new_P3_ADD_476_U51, new_P3_ADD_476_U52, new_P3_ADD_476_U53,
    new_P3_ADD_476_U54, new_P3_ADD_476_U55, new_P3_ADD_476_U56,
    new_P3_ADD_476_U57, new_P3_ADD_476_U58, new_P3_ADD_476_U59,
    new_P3_ADD_476_U60, new_P3_ADD_476_U61, new_P3_ADD_476_U62,
    new_P3_ADD_476_U63, new_P3_ADD_476_U64, new_P3_ADD_476_U65,
    new_P3_ADD_476_U66, new_P3_ADD_476_U67, new_P3_ADD_476_U68,
    new_P3_ADD_476_U69, new_P3_ADD_476_U70, new_P3_ADD_476_U71,
    new_P3_ADD_476_U72, new_P3_ADD_476_U73, new_P3_ADD_476_U74,
    new_P3_ADD_476_U75, new_P3_ADD_476_U76, new_P3_ADD_476_U77,
    new_P3_ADD_476_U78, new_P3_ADD_476_U79, new_P3_ADD_476_U80,
    new_P3_ADD_476_U81, new_P3_ADD_476_U82, new_P3_ADD_476_U83,
    new_P3_ADD_476_U84, new_P3_ADD_476_U85, new_P3_ADD_476_U86,
    new_P3_ADD_476_U87, new_P3_ADD_476_U88, new_P3_ADD_476_U89,
    new_P3_ADD_476_U90, new_P3_ADD_476_U91, new_P3_ADD_476_U92,
    new_P3_ADD_476_U93, new_P3_ADD_476_U94, new_P3_ADD_476_U95,
    new_P3_ADD_476_U96, new_P3_ADD_476_U97, new_P3_ADD_476_U98,
    new_P3_ADD_476_U99, new_P3_ADD_476_U100, new_P3_ADD_476_U101,
    new_P3_ADD_476_U102, new_P3_ADD_476_U103, new_P3_ADD_476_U104,
    new_P3_ADD_476_U105, new_P3_ADD_476_U106, new_P3_ADD_476_U107,
    new_P3_ADD_476_U108, new_P3_ADD_476_U109, new_P3_ADD_476_U110,
    new_P3_ADD_476_U111, new_P3_ADD_476_U112, new_P3_ADD_476_U113,
    new_P3_ADD_476_U114, new_P3_ADD_476_U115, new_P3_ADD_476_U116,
    new_P3_ADD_476_U117, new_P3_ADD_476_U118, new_P3_ADD_476_U119,
    new_P3_ADD_476_U120, new_P3_ADD_476_U121, new_P3_ADD_476_U122,
    new_P3_ADD_476_U123, new_P3_ADD_476_U124, new_P3_ADD_476_U125,
    new_P3_ADD_476_U126, new_P3_ADD_476_U127, new_P3_ADD_476_U128,
    new_P3_ADD_476_U129, new_P3_ADD_476_U130, new_P3_ADD_476_U131,
    new_P3_ADD_476_U132, new_P3_ADD_476_U133, new_P3_ADD_476_U134,
    new_P3_ADD_476_U135, new_P3_ADD_476_U136, new_P3_ADD_476_U137,
    new_P3_ADD_476_U138, new_P3_ADD_476_U139, new_P3_ADD_476_U140,
    new_P3_ADD_476_U141, new_P3_ADD_476_U142, new_P3_ADD_476_U143,
    new_P3_ADD_476_U144, new_P3_ADD_476_U145, new_P3_ADD_476_U146,
    new_P3_ADD_476_U147, new_P3_ADD_476_U148, new_P3_ADD_476_U149,
    new_P3_ADD_476_U150, new_P3_ADD_476_U151, new_P3_ADD_476_U152,
    new_P3_ADD_476_U153, new_P3_ADD_476_U154, new_P3_ADD_476_U155,
    new_P3_ADD_476_U156, new_P3_ADD_476_U157, new_P3_ADD_476_U158,
    new_P3_ADD_476_U159, new_P3_ADD_476_U160, new_P3_ADD_476_U161,
    new_P3_ADD_476_U162, new_P3_ADD_476_U163, new_P3_ADD_476_U164,
    new_P3_ADD_476_U165, new_P3_ADD_476_U166, new_P3_ADD_476_U167,
    new_P3_ADD_476_U168, new_P3_ADD_476_U169, new_P3_ADD_476_U170,
    new_P3_ADD_476_U171, new_P3_ADD_476_U172, new_P3_ADD_476_U173,
    new_P3_ADD_476_U174, new_P3_ADD_476_U175, new_P3_ADD_476_U176,
    new_P3_ADD_476_U177, new_P3_ADD_476_U178, new_P3_ADD_476_U179,
    new_P3_ADD_476_U180, new_P3_ADD_476_U181, new_P3_ADD_476_U182,
    new_P3_GTE_390_U6, new_P3_GTE_390_U7, new_P3_GTE_390_U8,
    new_P3_GTE_390_U9, new_P3_ADD_531_U5, new_P3_ADD_531_U6,
    new_P3_ADD_531_U7, new_P3_ADD_531_U8, new_P3_ADD_531_U9,
    new_P3_ADD_531_U10, new_P3_ADD_531_U11, new_P3_ADD_531_U12,
    new_P3_ADD_531_U13, new_P3_ADD_531_U14, new_P3_ADD_531_U15,
    new_P3_ADD_531_U16, new_P3_ADD_531_U17, new_P3_ADD_531_U18,
    new_P3_ADD_531_U19, new_P3_ADD_531_U20, new_P3_ADD_531_U21,
    new_P3_ADD_531_U22, new_P3_ADD_531_U23, new_P3_ADD_531_U24,
    new_P3_ADD_531_U25, new_P3_ADD_531_U26, new_P3_ADD_531_U27,
    new_P3_ADD_531_U28, new_P3_ADD_531_U29, new_P3_ADD_531_U30,
    new_P3_ADD_531_U31, new_P3_ADD_531_U32, new_P3_ADD_531_U33,
    new_P3_ADD_531_U34, new_P3_ADD_531_U35, new_P3_ADD_531_U36,
    new_P3_ADD_531_U37, new_P3_ADD_531_U38, new_P3_ADD_531_U39,
    new_P3_ADD_531_U40, new_P3_ADD_531_U41, new_P3_ADD_531_U42,
    new_P3_ADD_531_U43, new_P3_ADD_531_U44, new_P3_ADD_531_U45,
    new_P3_ADD_531_U46, new_P3_ADD_531_U47, new_P3_ADD_531_U48,
    new_P3_ADD_531_U49, new_P3_ADD_531_U50, new_P3_ADD_531_U51,
    new_P3_ADD_531_U52, new_P3_ADD_531_U53, new_P3_ADD_531_U54,
    new_P3_ADD_531_U55, new_P3_ADD_531_U56, new_P3_ADD_531_U57,
    new_P3_ADD_531_U58, new_P3_ADD_531_U59, new_P3_ADD_531_U60,
    new_P3_ADD_531_U61, new_P3_ADD_531_U62, new_P3_ADD_531_U63,
    new_P3_ADD_531_U64, new_P3_ADD_531_U65, new_P3_ADD_531_U66,
    new_P3_ADD_531_U67, new_P3_ADD_531_U68, new_P3_ADD_531_U69,
    new_P3_ADD_531_U70, new_P3_ADD_531_U71, new_P3_ADD_531_U72,
    new_P3_ADD_531_U73, new_P3_ADD_531_U74, new_P3_ADD_531_U75,
    new_P3_ADD_531_U76, new_P3_ADD_531_U77, new_P3_ADD_531_U78,
    new_P3_ADD_531_U79, new_P3_ADD_531_U80, new_P3_ADD_531_U81,
    new_P3_ADD_531_U82, new_P3_ADD_531_U83, new_P3_ADD_531_U84,
    new_P3_ADD_531_U85, new_P3_ADD_531_U86, new_P3_ADD_531_U87,
    new_P3_ADD_531_U88, new_P3_ADD_531_U89, new_P3_ADD_531_U90,
    new_P3_ADD_531_U91, new_P3_ADD_531_U92, new_P3_ADD_531_U93,
    new_P3_ADD_531_U94, new_P3_ADD_531_U95, new_P3_ADD_531_U96,
    new_P3_ADD_531_U97, new_P3_ADD_531_U98, new_P3_ADD_531_U99,
    new_P3_ADD_531_U100, new_P3_ADD_531_U101, new_P3_ADD_531_U102,
    new_P3_ADD_531_U103, new_P3_ADD_531_U104, new_P3_ADD_531_U105,
    new_P3_ADD_531_U106, new_P3_ADD_531_U107, new_P3_ADD_531_U108,
    new_P3_ADD_531_U109, new_P3_ADD_531_U110, new_P3_ADD_531_U111,
    new_P3_ADD_531_U112, new_P3_ADD_531_U113, new_P3_ADD_531_U114,
    new_P3_ADD_531_U115, new_P3_ADD_531_U116, new_P3_ADD_531_U117,
    new_P3_ADD_531_U118, new_P3_ADD_531_U119, new_P3_ADD_531_U120,
    new_P3_ADD_531_U121, new_P3_ADD_531_U122, new_P3_ADD_531_U123,
    new_P3_ADD_531_U124, new_P3_ADD_531_U125, new_P3_ADD_531_U126,
    new_P3_ADD_531_U127, new_P3_ADD_531_U128, new_P3_ADD_531_U129,
    new_P3_ADD_531_U130, new_P3_ADD_531_U131, new_P3_ADD_531_U132,
    new_P3_ADD_531_U133, new_P3_ADD_531_U134, new_P3_ADD_531_U135,
    new_P3_ADD_531_U136, new_P3_ADD_531_U137, new_P3_ADD_531_U138,
    new_P3_ADD_531_U139, new_P3_ADD_531_U140, new_P3_ADD_531_U141,
    new_P3_ADD_531_U142, new_P3_ADD_531_U143, new_P3_ADD_531_U144,
    new_P3_ADD_531_U145, new_P3_ADD_531_U146, new_P3_ADD_531_U147,
    new_P3_ADD_531_U148, new_P3_ADD_531_U149, new_P3_ADD_531_U150,
    new_P3_ADD_531_U151, new_P3_ADD_531_U152, new_P3_ADD_531_U153,
    new_P3_ADD_531_U154, new_P3_ADD_531_U155, new_P3_ADD_531_U156,
    new_P3_ADD_531_U157, new_P3_ADD_531_U158, new_P3_ADD_531_U159,
    new_P3_ADD_531_U160, new_P3_ADD_531_U161, new_P3_ADD_531_U162,
    new_P3_ADD_531_U163, new_P3_ADD_531_U164, new_P3_ADD_531_U165,
    new_P3_ADD_531_U166, new_P3_ADD_531_U167, new_P3_ADD_531_U168,
    new_P3_ADD_531_U169, new_P3_ADD_531_U170, new_P3_ADD_531_U171,
    new_P3_ADD_531_U172, new_P3_ADD_531_U173, new_P3_ADD_531_U174,
    new_P3_ADD_531_U175, new_P3_ADD_531_U176, new_P3_ADD_531_U177,
    new_P3_ADD_531_U178, new_P3_ADD_531_U179, new_P3_ADD_531_U180,
    new_P3_ADD_531_U181, new_P3_ADD_531_U182, new_P3_ADD_531_U183,
    new_P3_ADD_531_U184, new_P3_ADD_531_U185, new_P3_ADD_531_U186,
    new_P3_ADD_531_U187, new_P3_ADD_531_U188, new_P3_ADD_531_U189,
    new_P3_SUB_320_U6, new_P3_SUB_320_U7, new_P3_SUB_320_U8,
    new_P3_SUB_320_U9, new_P3_SUB_320_U10, new_P3_SUB_320_U11,
    new_P3_SUB_320_U12, new_P3_SUB_320_U13, new_P3_SUB_320_U14,
    new_P3_SUB_320_U15, new_P3_SUB_320_U16, new_P3_SUB_320_U17,
    new_P3_SUB_320_U18, new_P3_SUB_320_U19, new_P3_SUB_320_U20,
    new_P3_SUB_320_U21, new_P3_SUB_320_U22, new_P3_SUB_320_U23,
    new_P3_SUB_320_U24, new_P3_SUB_320_U25, new_P3_SUB_320_U26,
    new_P3_SUB_320_U27, new_P3_SUB_320_U28, new_P3_SUB_320_U29,
    new_P3_SUB_320_U30, new_P3_SUB_320_U31, new_P3_SUB_320_U32,
    new_P3_SUB_320_U33, new_P3_SUB_320_U34, new_P3_SUB_320_U35,
    new_P3_SUB_320_U36, new_P3_SUB_320_U37, new_P3_SUB_320_U38,
    new_P3_SUB_320_U39, new_P3_SUB_320_U40, new_P3_SUB_320_U41,
    new_P3_SUB_320_U42, new_P3_SUB_320_U43, new_P3_SUB_320_U44,
    new_P3_SUB_320_U45, new_P3_SUB_320_U46, new_P3_SUB_320_U47,
    new_P3_SUB_320_U48, new_P3_SUB_320_U49, new_P3_SUB_320_U50,
    new_P3_SUB_320_U51, new_P3_SUB_320_U52, new_P3_SUB_320_U53,
    new_P3_SUB_320_U54, new_P3_SUB_320_U55, new_P3_SUB_320_U56,
    new_P3_SUB_320_U57, new_P3_SUB_320_U58, new_P3_SUB_320_U59,
    new_P3_SUB_320_U60, new_P3_SUB_320_U61, new_P3_SUB_320_U62,
    new_P3_SUB_320_U63, new_P3_SUB_320_U64, new_P3_SUB_320_U65,
    new_P3_SUB_320_U66, new_P3_SUB_320_U67, new_P3_SUB_320_U68,
    new_P3_SUB_320_U69, new_P3_SUB_320_U70, new_P3_SUB_320_U71,
    new_P3_SUB_320_U72, new_P3_SUB_320_U73, new_P3_SUB_320_U74,
    new_P3_SUB_320_U75, new_P3_SUB_320_U76, new_P3_SUB_320_U77,
    new_P3_SUB_320_U78, new_P3_SUB_320_U79, new_P3_SUB_320_U80,
    new_P3_SUB_320_U81, new_P3_SUB_320_U82, new_P3_SUB_320_U83,
    new_P3_SUB_320_U84, new_P3_SUB_320_U85, new_P3_SUB_320_U86,
    new_P3_SUB_320_U87, new_P3_SUB_320_U88, new_P3_SUB_320_U89,
    new_P3_SUB_320_U90, new_P3_SUB_320_U91, new_P3_SUB_320_U92,
    new_P3_SUB_320_U93, new_P3_SUB_320_U94, new_P3_SUB_320_U95,
    new_P3_SUB_320_U96, new_P3_SUB_320_U97, new_P3_SUB_320_U98,
    new_P3_SUB_320_U99, new_P3_SUB_320_U100, new_P3_SUB_320_U101,
    new_P3_SUB_320_U102, new_P3_SUB_320_U103, new_P3_SUB_320_U104,
    new_P3_SUB_320_U105, new_P3_SUB_320_U106, new_P3_SUB_320_U107,
    new_P3_SUB_320_U108, new_P3_SUB_320_U109, new_P3_SUB_320_U110,
    new_P3_SUB_320_U111, new_P3_SUB_320_U112, new_P3_SUB_320_U113,
    new_P3_SUB_320_U114, new_P3_SUB_320_U115, new_P3_SUB_320_U116,
    new_P3_SUB_320_U117, new_P3_SUB_320_U118, new_P3_SUB_320_U119,
    new_P3_SUB_320_U120, new_P3_SUB_320_U121, new_P3_SUB_320_U122,
    new_P3_SUB_320_U123, new_P3_SUB_320_U124, new_P3_SUB_320_U125,
    new_P3_SUB_320_U126, new_P3_SUB_320_U127, new_P3_SUB_320_U128,
    new_P3_SUB_320_U129, new_P3_SUB_320_U130, new_P3_SUB_320_U131,
    new_P3_SUB_320_U132, new_P3_SUB_320_U133, new_P3_SUB_320_U134,
    new_P3_SUB_320_U135, new_P3_SUB_320_U136, new_P3_SUB_320_U137,
    new_P3_SUB_320_U138, new_P3_SUB_320_U139, new_P3_SUB_320_U140,
    new_P3_SUB_320_U141, new_P3_SUB_320_U142, new_P3_SUB_320_U143,
    new_P3_SUB_320_U144, new_P3_SUB_320_U145, new_P3_SUB_320_U146,
    new_P3_SUB_320_U147, new_P3_SUB_320_U148, new_P3_SUB_320_U149,
    new_P3_SUB_320_U150, new_P3_SUB_320_U151, new_P3_SUB_320_U152,
    new_P3_SUB_320_U153, new_P3_SUB_320_U154, new_P3_SUB_320_U155,
    new_P3_SUB_320_U156, new_P3_SUB_320_U157, new_P3_SUB_320_U158,
    new_P3_SUB_320_U159, new_P3_ADD_505_U5, new_P3_ADD_505_U6,
    new_P3_ADD_505_U7, new_P3_ADD_505_U8, new_P3_ADD_505_U9,
    new_P3_ADD_505_U10, new_P3_ADD_505_U11, new_P3_ADD_505_U12,
    new_P3_ADD_505_U13, new_P3_ADD_505_U14, new_P3_ADD_505_U15,
    new_P3_ADD_505_U16, new_P3_ADD_505_U17, new_P3_ADD_505_U18,
    new_P3_ADD_505_U19, new_P3_ADD_505_U20, new_P3_ADD_505_U21,
    new_P3_ADD_505_U22, new_P3_ADD_505_U23, new_P3_ADD_505_U24,
    new_P3_ADD_505_U25, new_P3_ADD_505_U26, new_P3_ADD_505_U27,
    new_P3_ADD_505_U28, new_P3_GTE_485_U6, new_P3_GTE_485_U7,
    new_P3_ADD_318_U4, new_P3_ADD_318_U5, new_P3_ADD_318_U6,
    new_P3_ADD_318_U7, new_P3_ADD_318_U8, new_P3_ADD_318_U9,
    new_P3_ADD_318_U10, new_P3_ADD_318_U11, new_P3_ADD_318_U12,
    new_P3_ADD_318_U13, new_P3_ADD_318_U14, new_P3_ADD_318_U15,
    new_P3_ADD_318_U16, new_P3_ADD_318_U17, new_P3_ADD_318_U18,
    new_P3_ADD_318_U19, new_P3_ADD_318_U20, new_P3_ADD_318_U21,
    new_P3_ADD_318_U22, new_P3_ADD_318_U23, new_P3_ADD_318_U24,
    new_P3_ADD_318_U25, new_P3_ADD_318_U26, new_P3_ADD_318_U27,
    new_P3_ADD_318_U28, new_P3_ADD_318_U29, new_P3_ADD_318_U30,
    new_P3_ADD_318_U31, new_P3_ADD_318_U32, new_P3_ADD_318_U33,
    new_P3_ADD_318_U34, new_P3_ADD_318_U35, new_P3_ADD_318_U36,
    new_P3_ADD_318_U37, new_P3_ADD_318_U38, new_P3_ADD_318_U39,
    new_P3_ADD_318_U40, new_P3_ADD_318_U41, new_P3_ADD_318_U42,
    new_P3_ADD_318_U43, new_P3_ADD_318_U44, new_P3_ADD_318_U45,
    new_P3_ADD_318_U46, new_P3_ADD_318_U47, new_P3_ADD_318_U48,
    new_P3_ADD_318_U49, new_P3_ADD_318_U50, new_P3_ADD_318_U51,
    new_P3_ADD_318_U52, new_P3_ADD_318_U53, new_P3_ADD_318_U54,
    new_P3_ADD_318_U55, new_P3_ADD_318_U56, new_P3_ADD_318_U57,
    new_P3_ADD_318_U58, new_P3_ADD_318_U59, new_P3_ADD_318_U60,
    new_P3_ADD_318_U61, new_P3_ADD_318_U62, new_P3_ADD_318_U63,
    new_P3_ADD_318_U64, new_P3_ADD_318_U65, new_P3_ADD_318_U66,
    new_P3_ADD_318_U67, new_P3_ADD_318_U68, new_P3_ADD_318_U69,
    new_P3_ADD_318_U70, new_P3_ADD_318_U71, new_P3_ADD_318_U72,
    new_P3_ADD_318_U73, new_P3_ADD_318_U74, new_P3_ADD_318_U75,
    new_P3_ADD_318_U76, new_P3_ADD_318_U77, new_P3_ADD_318_U78,
    new_P3_ADD_318_U79, new_P3_ADD_318_U80, new_P3_ADD_318_U81,
    new_P3_ADD_318_U82, new_P3_ADD_318_U83, new_P3_ADD_318_U84,
    new_P3_ADD_318_U85, new_P3_ADD_318_U86, new_P3_ADD_318_U87,
    new_P3_ADD_318_U88, new_P3_ADD_318_U89, new_P3_ADD_318_U90,
    new_P3_ADD_318_U91, new_P3_ADD_318_U92, new_P3_ADD_318_U93,
    new_P3_ADD_318_U94, new_P3_ADD_318_U95, new_P3_ADD_318_U96,
    new_P3_ADD_318_U97, new_P3_ADD_318_U98, new_P3_ADD_318_U99,
    new_P3_ADD_318_U100, new_P3_ADD_318_U101, new_P3_ADD_318_U102,
    new_P3_ADD_318_U103, new_P3_ADD_318_U104, new_P3_ADD_318_U105,
    new_P3_ADD_318_U106, new_P3_ADD_318_U107, new_P3_ADD_318_U108,
    new_P3_ADD_318_U109, new_P3_ADD_318_U110, new_P3_ADD_318_U111,
    new_P3_ADD_318_U112, new_P3_ADD_318_U113, new_P3_ADD_318_U114,
    new_P3_ADD_318_U115, new_P3_ADD_318_U116, new_P3_ADD_318_U117,
    new_P3_ADD_318_U118, new_P3_ADD_318_U119, new_P3_ADD_318_U120,
    new_P3_ADD_318_U121, new_P3_ADD_318_U122, new_P3_ADD_318_U123,
    new_P3_ADD_318_U124, new_P3_ADD_318_U125, new_P3_ADD_318_U126,
    new_P3_ADD_318_U127, new_P3_ADD_318_U128, new_P3_ADD_318_U129,
    new_P3_ADD_318_U130, new_P3_ADD_318_U131, new_P3_ADD_318_U132,
    new_P3_ADD_318_U133, new_P3_ADD_318_U134, new_P3_ADD_318_U135,
    new_P3_ADD_318_U136, new_P3_ADD_318_U137, new_P3_ADD_318_U138,
    new_P3_ADD_318_U139, new_P3_ADD_318_U140, new_P3_ADD_318_U141,
    new_P3_ADD_318_U142, new_P3_ADD_318_U143, new_P3_ADD_318_U144,
    new_P3_ADD_318_U145, new_P3_ADD_318_U146, new_P3_ADD_318_U147,
    new_P3_ADD_318_U148, new_P3_ADD_318_U149, new_P3_ADD_318_U150,
    new_P3_ADD_318_U151, new_P3_ADD_318_U152, new_P3_ADD_318_U153,
    new_P3_ADD_318_U154, new_P3_ADD_318_U155, new_P3_ADD_318_U156,
    new_P3_ADD_318_U157, new_P3_ADD_318_U158, new_P3_ADD_318_U159,
    new_P3_ADD_318_U160, new_P3_ADD_318_U161, new_P3_ADD_318_U162,
    new_P3_ADD_318_U163, new_P3_ADD_318_U164, new_P3_ADD_318_U165,
    new_P3_ADD_318_U166, new_P3_ADD_318_U167, new_P3_ADD_318_U168,
    new_P3_ADD_318_U169, new_P3_ADD_318_U170, new_P3_ADD_318_U171,
    new_P3_ADD_318_U172, new_P3_ADD_318_U173, new_P3_ADD_318_U174,
    new_P3_ADD_318_U175, new_P3_ADD_318_U176, new_P3_ADD_318_U177,
    new_P3_ADD_318_U178, new_P3_ADD_318_U179, new_P3_ADD_318_U180,
    new_P3_ADD_318_U181, new_P3_ADD_318_U182, new_P3_SUB_370_U6,
    new_P3_SUB_370_U7, new_P3_SUB_370_U8, new_P3_SUB_370_U9,
    new_P3_SUB_370_U10, new_P3_SUB_370_U11, new_P3_SUB_370_U12,
    new_P3_SUB_370_U13, new_P3_SUB_370_U14, new_P3_SUB_370_U15,
    new_P3_SUB_370_U16, new_P3_SUB_370_U17, new_P3_SUB_370_U18,
    new_P3_SUB_370_U19, new_P3_SUB_370_U20, new_P3_SUB_370_U21,
    new_P3_SUB_370_U22, new_P3_SUB_370_U23, new_P3_SUB_370_U24,
    new_P3_SUB_370_U25, new_P3_SUB_370_U26, new_P3_SUB_370_U27,
    new_P3_SUB_370_U28, new_P3_SUB_370_U29, new_P3_SUB_370_U30,
    new_P3_SUB_370_U31, new_P3_SUB_370_U32, new_P3_SUB_370_U33,
    new_P3_SUB_370_U34, new_P3_SUB_370_U35, new_P3_SUB_370_U36,
    new_P3_SUB_370_U37, new_P3_SUB_370_U38, new_P3_SUB_370_U39,
    new_P3_SUB_370_U40, new_P3_SUB_370_U41, new_P3_SUB_370_U42,
    new_P3_SUB_370_U43, new_P3_SUB_370_U44, new_P3_SUB_370_U45,
    new_P3_SUB_370_U46, new_P3_SUB_370_U47, new_P3_SUB_370_U48,
    new_P3_SUB_370_U49, new_P3_SUB_370_U50, new_P3_SUB_370_U51,
    new_P3_SUB_370_U52, new_P3_SUB_370_U53, new_P3_SUB_370_U54,
    new_P3_SUB_370_U55, new_P3_SUB_370_U56, new_P3_SUB_370_U57,
    new_P3_SUB_370_U58, new_P3_SUB_370_U59, new_P3_SUB_370_U60,
    new_P3_SUB_370_U61, new_P3_SUB_370_U62, new_P3_SUB_370_U63,
    new_P3_SUB_370_U64, new_P3_SUB_370_U65, new_P3_SUB_370_U66,
    new_P3_ADD_315_U4, new_P3_ADD_315_U5, new_P3_ADD_315_U6,
    new_P3_ADD_315_U7, new_P3_ADD_315_U8, new_P3_ADD_315_U9,
    new_P3_ADD_315_U10, new_P3_ADD_315_U11, new_P3_ADD_315_U12,
    new_P3_ADD_315_U13, new_P3_ADD_315_U14, new_P3_ADD_315_U15,
    new_P3_ADD_315_U16, new_P3_ADD_315_U17, new_P3_ADD_315_U18,
    new_P3_ADD_315_U19, new_P3_ADD_315_U20, new_P3_ADD_315_U21,
    new_P3_ADD_315_U22, new_P3_ADD_315_U23, new_P3_ADD_315_U24,
    new_P3_ADD_315_U25, new_P3_ADD_315_U26, new_P3_ADD_315_U27,
    new_P3_ADD_315_U28, new_P3_ADD_315_U29, new_P3_ADD_315_U30,
    new_P3_ADD_315_U31, new_P3_ADD_315_U32, new_P3_ADD_315_U33,
    new_P3_ADD_315_U34, new_P3_ADD_315_U35, new_P3_ADD_315_U36,
    new_P3_ADD_315_U37, new_P3_ADD_315_U38, new_P3_ADD_315_U39,
    new_P3_ADD_315_U40, new_P3_ADD_315_U41, new_P3_ADD_315_U42,
    new_P3_ADD_315_U43, new_P3_ADD_315_U44, new_P3_ADD_315_U45,
    new_P3_ADD_315_U46, new_P3_ADD_315_U47, new_P3_ADD_315_U48,
    new_P3_ADD_315_U49, new_P3_ADD_315_U50, new_P3_ADD_315_U51,
    new_P3_ADD_315_U52, new_P3_ADD_315_U53, new_P3_ADD_315_U54,
    new_P3_ADD_315_U55, new_P3_ADD_315_U56, new_P3_ADD_315_U57,
    new_P3_ADD_315_U58, new_P3_ADD_315_U59, new_P3_ADD_315_U60,
    new_P3_ADD_315_U61, new_P3_ADD_315_U62, new_P3_ADD_315_U63,
    new_P3_ADD_315_U64, new_P3_ADD_315_U65, new_P3_ADD_315_U66,
    new_P3_ADD_315_U67, new_P3_ADD_315_U68, new_P3_ADD_315_U69,
    new_P3_ADD_315_U70, new_P3_ADD_315_U71, new_P3_ADD_315_U72,
    new_P3_ADD_315_U73, new_P3_ADD_315_U74, new_P3_ADD_315_U75,
    new_P3_ADD_315_U76, new_P3_ADD_315_U77, new_P3_ADD_315_U78,
    new_P3_ADD_315_U79, new_P3_ADD_315_U80, new_P3_ADD_315_U81,
    new_P3_ADD_315_U82, new_P3_ADD_315_U83, new_P3_ADD_315_U84,
    new_P3_ADD_315_U85, new_P3_ADD_315_U86, new_P3_ADD_315_U87,
    new_P3_ADD_315_U88, new_P3_ADD_315_U89, new_P3_ADD_315_U90,
    new_P3_ADD_315_U91, new_P3_ADD_315_U92, new_P3_ADD_315_U93,
    new_P3_ADD_315_U94, new_P3_ADD_315_U95, new_P3_ADD_315_U96,
    new_P3_ADD_315_U97, new_P3_ADD_315_U98, new_P3_ADD_315_U99,
    new_P3_ADD_315_U100, new_P3_ADD_315_U101, new_P3_ADD_315_U102,
    new_P3_ADD_315_U103, new_P3_ADD_315_U104, new_P3_ADD_315_U105,
    new_P3_ADD_315_U106, new_P3_ADD_315_U107, new_P3_ADD_315_U108,
    new_P3_ADD_315_U109, new_P3_ADD_315_U110, new_P3_ADD_315_U111,
    new_P3_ADD_315_U112, new_P3_ADD_315_U113, new_P3_ADD_315_U114,
    new_P3_ADD_315_U115, new_P3_ADD_315_U116, new_P3_ADD_315_U117,
    new_P3_ADD_315_U118, new_P3_ADD_315_U119, new_P3_ADD_315_U120,
    new_P3_ADD_315_U121, new_P3_ADD_315_U122, new_P3_ADD_315_U123,
    new_P3_ADD_315_U124, new_P3_ADD_315_U125, new_P3_ADD_315_U126,
    new_P3_ADD_315_U127, new_P3_ADD_315_U128, new_P3_ADD_315_U129,
    new_P3_ADD_315_U130, new_P3_ADD_315_U131, new_P3_ADD_315_U132,
    new_P3_ADD_315_U133, new_P3_ADD_315_U134, new_P3_ADD_315_U135,
    new_P3_ADD_315_U136, new_P3_ADD_315_U137, new_P3_ADD_315_U138,
    new_P3_ADD_315_U139, new_P3_ADD_315_U140, new_P3_ADD_315_U141,
    new_P3_ADD_315_U142, new_P3_ADD_315_U143, new_P3_ADD_315_U144,
    new_P3_ADD_315_U145, new_P3_ADD_315_U146, new_P3_ADD_315_U147,
    new_P3_ADD_315_U148, new_P3_ADD_315_U149, new_P3_ADD_315_U150,
    new_P3_ADD_315_U151, new_P3_ADD_315_U152, new_P3_ADD_315_U153,
    new_P3_ADD_315_U154, new_P3_ADD_315_U155, new_P3_ADD_315_U156,
    new_P3_ADD_315_U157, new_P3_ADD_315_U158, new_P3_ADD_315_U159,
    new_P3_ADD_315_U160, new_P3_ADD_315_U161, new_P3_ADD_315_U162,
    new_P3_ADD_315_U163, new_P3_ADD_315_U164, new_P3_ADD_315_U165,
    new_P3_ADD_315_U166, new_P3_ADD_315_U167, new_P3_ADD_315_U168,
    new_P3_ADD_315_U169, new_P3_ADD_315_U170, new_P3_ADD_315_U171,
    new_P3_ADD_315_U172, new_P3_ADD_315_U173, new_P3_ADD_315_U174,
    new_P3_ADD_315_U175, new_P3_ADD_315_U176, new_P3_GTE_355_U6,
    new_P3_GTE_355_U7, new_P3_GTE_355_U8, new_P3_ADD_360_1242_U4,
    new_P3_ADD_360_1242_U5, new_P3_ADD_360_1242_U6, new_P3_ADD_360_1242_U7,
    new_P3_ADD_360_1242_U8, new_P3_ADD_360_1242_U9,
    new_P3_ADD_360_1242_U10, new_P3_ADD_360_1242_U11,
    new_P3_ADD_360_1242_U12, new_P3_ADD_360_1242_U13,
    new_P3_ADD_360_1242_U14, new_P3_ADD_360_1242_U15,
    new_P3_ADD_360_1242_U16, new_P3_ADD_360_1242_U17,
    new_P3_ADD_360_1242_U18, new_P3_ADD_360_1242_U19,
    new_P3_ADD_360_1242_U20, new_P3_ADD_360_1242_U21,
    new_P3_ADD_360_1242_U22, new_P3_ADD_360_1242_U23,
    new_P3_ADD_360_1242_U24, new_P3_ADD_360_1242_U25,
    new_P3_ADD_360_1242_U26, new_P3_ADD_360_1242_U27,
    new_P3_ADD_360_1242_U28, new_P3_ADD_360_1242_U29,
    new_P3_ADD_360_1242_U30, new_P3_ADD_360_1242_U31,
    new_P3_ADD_360_1242_U32, new_P3_ADD_360_1242_U33,
    new_P3_ADD_360_1242_U34, new_P3_ADD_360_1242_U35,
    new_P3_ADD_360_1242_U36, new_P3_ADD_360_1242_U37,
    new_P3_ADD_360_1242_U38, new_P3_ADD_360_1242_U39,
    new_P3_ADD_360_1242_U40, new_P3_ADD_360_1242_U41,
    new_P3_ADD_360_1242_U42, new_P3_ADD_360_1242_U43,
    new_P3_ADD_360_1242_U44, new_P3_ADD_360_1242_U45,
    new_P3_ADD_360_1242_U46, new_P3_ADD_360_1242_U47,
    new_P3_ADD_360_1242_U48, new_P3_ADD_360_1242_U49,
    new_P3_ADD_360_1242_U50, new_P3_ADD_360_1242_U51,
    new_P3_ADD_360_1242_U52, new_P3_ADD_360_1242_U53,
    new_P3_ADD_360_1242_U54, new_P3_ADD_360_1242_U55,
    new_P3_ADD_360_1242_U56, new_P3_ADD_360_1242_U57,
    new_P3_ADD_360_1242_U58, new_P3_ADD_360_1242_U59,
    new_P3_ADD_360_1242_U60, new_P3_ADD_360_1242_U61,
    new_P3_ADD_360_1242_U62, new_P3_ADD_360_1242_U63,
    new_P3_ADD_360_1242_U64, new_P3_ADD_360_1242_U65,
    new_P3_ADD_360_1242_U66, new_P3_ADD_360_1242_U67,
    new_P3_ADD_360_1242_U68, new_P3_ADD_360_1242_U69,
    new_P3_ADD_360_1242_U70, new_P3_ADD_360_1242_U71,
    new_P3_ADD_360_1242_U72, new_P3_ADD_360_1242_U73,
    new_P3_ADD_360_1242_U74, new_P3_ADD_360_1242_U75,
    new_P3_ADD_360_1242_U76, new_P3_ADD_360_1242_U77,
    new_P3_ADD_360_1242_U78, new_P3_ADD_360_1242_U79,
    new_P3_ADD_360_1242_U80, new_P3_ADD_360_1242_U81,
    new_P3_ADD_360_1242_U82, new_P3_ADD_360_1242_U83,
    new_P3_ADD_360_1242_U84, new_P3_ADD_360_1242_U85,
    new_P3_ADD_360_1242_U86, new_P3_ADD_360_1242_U87,
    new_P3_ADD_360_1242_U88, new_P3_ADD_360_1242_U89,
    new_P3_ADD_360_1242_U90, new_P3_ADD_360_1242_U91,
    new_P3_ADD_360_1242_U92, new_P3_ADD_360_1242_U93,
    new_P3_ADD_360_1242_U94, new_P3_ADD_360_1242_U95,
    new_P3_ADD_360_1242_U96, new_P3_ADD_360_1242_U97,
    new_P3_ADD_360_1242_U98, new_P3_ADD_360_1242_U99,
    new_P3_ADD_360_1242_U100, new_P3_ADD_360_1242_U101,
    new_P3_ADD_360_1242_U102, new_P3_ADD_360_1242_U103,
    new_P3_ADD_360_1242_U104, new_P3_ADD_360_1242_U105,
    new_P3_ADD_360_1242_U106, new_P3_ADD_360_1242_U107,
    new_P3_ADD_360_1242_U108, new_P3_ADD_360_1242_U109,
    new_P3_ADD_360_1242_U110, new_P3_ADD_360_1242_U111,
    new_P3_ADD_360_1242_U112, new_P3_ADD_360_1242_U113,
    new_P3_ADD_360_1242_U114, new_P3_ADD_360_1242_U115,
    new_P3_ADD_360_1242_U116, new_P3_ADD_360_1242_U117,
    new_P3_ADD_360_1242_U118, new_P3_ADD_360_1242_U119,
    new_P3_ADD_360_1242_U120, new_P3_ADD_360_1242_U121,
    new_P3_ADD_360_1242_U122, new_P3_ADD_360_1242_U123,
    new_P3_ADD_360_1242_U124, new_P3_ADD_360_1242_U125,
    new_P3_ADD_360_1242_U126, new_P3_ADD_360_1242_U127,
    new_P3_ADD_360_1242_U128, new_P3_ADD_360_1242_U129,
    new_P3_ADD_360_1242_U130, new_P3_ADD_360_1242_U131,
    new_P3_ADD_360_1242_U132, new_P3_ADD_360_1242_U133,
    new_P3_ADD_360_1242_U134, new_P3_ADD_360_1242_U135,
    new_P3_ADD_360_1242_U136, new_P3_ADD_360_1242_U137,
    new_P3_ADD_360_1242_U138, new_P3_ADD_360_1242_U139,
    new_P3_ADD_360_1242_U140, new_P3_ADD_360_1242_U141,
    new_P3_ADD_360_1242_U142, new_P3_ADD_360_1242_U143,
    new_P3_ADD_360_1242_U144, new_P3_ADD_360_1242_U145,
    new_P3_ADD_360_1242_U146, new_P3_ADD_360_1242_U147,
    new_P3_ADD_360_1242_U148, new_P3_ADD_360_1242_U149,
    new_P3_ADD_360_1242_U150, new_P3_ADD_360_1242_U151,
    new_P3_ADD_360_1242_U152, new_P3_ADD_360_1242_U153,
    new_P3_ADD_360_1242_U154, new_P3_ADD_360_1242_U155,
    new_P3_ADD_360_1242_U156, new_P3_ADD_360_1242_U157,
    new_P3_ADD_360_1242_U158, new_P3_ADD_360_1242_U159,
    new_P3_ADD_360_1242_U160, new_P3_ADD_360_1242_U161,
    new_P3_ADD_360_1242_U162, new_P3_ADD_360_1242_U163,
    new_P3_ADD_360_1242_U164, new_P3_ADD_360_1242_U165,
    new_P3_ADD_360_1242_U166, new_P3_ADD_360_1242_U167,
    new_P3_ADD_360_1242_U168, new_P3_ADD_360_1242_U169,
    new_P3_ADD_360_1242_U170, new_P3_ADD_360_1242_U171,
    new_P3_ADD_360_1242_U172, new_P3_ADD_360_1242_U173,
    new_P3_ADD_360_1242_U174, new_P3_ADD_360_1242_U175,
    new_P3_ADD_360_1242_U176, new_P3_ADD_360_1242_U177,
    new_P3_ADD_360_1242_U178, new_P3_ADD_360_1242_U179,
    new_P3_ADD_360_1242_U180, new_P3_ADD_360_1242_U181,
    new_P3_ADD_360_1242_U182, new_P3_ADD_360_1242_U183,
    new_P3_ADD_360_1242_U184, new_P3_ADD_360_1242_U185,
    new_P3_ADD_360_1242_U186, new_P3_ADD_360_1242_U187,
    new_P3_ADD_360_1242_U188, new_P3_ADD_360_1242_U189,
    new_P3_ADD_360_1242_U190, new_P3_ADD_360_1242_U191,
    new_P3_ADD_360_1242_U192, new_P3_ADD_360_1242_U193,
    new_P3_ADD_360_1242_U194, new_P3_ADD_360_1242_U195,
    new_P3_ADD_360_1242_U196, new_P3_ADD_360_1242_U197,
    new_P3_ADD_360_1242_U198, new_P3_ADD_360_1242_U199,
    new_P3_ADD_360_1242_U200, new_P3_ADD_360_1242_U201,
    new_P3_ADD_360_1242_U202, new_P3_ADD_360_1242_U203,
    new_P3_ADD_360_1242_U204, new_P3_ADD_360_1242_U205,
    new_P3_ADD_360_1242_U206, new_P3_ADD_360_1242_U207,
    new_P3_ADD_360_1242_U208, new_P3_ADD_360_1242_U209,
    new_P3_ADD_360_1242_U210, new_P3_ADD_360_1242_U211,
    new_P3_ADD_360_1242_U212, new_P3_ADD_360_1242_U213,
    new_P3_ADD_360_1242_U214, new_P3_ADD_360_1242_U215,
    new_P3_ADD_360_1242_U216, new_P3_ADD_360_1242_U217,
    new_P3_ADD_360_1242_U218, new_P3_ADD_360_1242_U219,
    new_P3_ADD_360_1242_U220, new_P3_ADD_360_1242_U221,
    new_P3_ADD_360_1242_U222, new_P3_ADD_360_1242_U223,
    new_P3_ADD_360_1242_U224, new_P3_ADD_360_1242_U225,
    new_P3_ADD_360_1242_U226, new_P3_ADD_360_1242_U227,
    new_P3_ADD_360_1242_U228, new_P3_ADD_360_1242_U229,
    new_P3_ADD_360_1242_U230, new_P3_ADD_360_1242_U231,
    new_P3_ADD_360_1242_U232, new_P3_ADD_360_1242_U233,
    new_P3_ADD_360_1242_U234, new_P3_ADD_360_1242_U235,
    new_P3_ADD_360_1242_U236, new_P3_ADD_360_1242_U237,
    new_P3_ADD_360_1242_U238, new_P3_ADD_360_1242_U239,
    new_P3_ADD_360_1242_U240, new_P3_ADD_360_1242_U241,
    new_P3_ADD_360_1242_U242, new_P3_ADD_360_1242_U243,
    new_P3_ADD_360_1242_U244, new_P3_ADD_360_1242_U245,
    new_P3_ADD_360_1242_U246, new_P3_ADD_360_1242_U247,
    new_P3_ADD_360_1242_U248, new_P3_ADD_360_1242_U249,
    new_P3_ADD_360_1242_U250, new_P3_ADD_360_1242_U251,
    new_P3_ADD_360_1242_U252, new_P3_ADD_360_1242_U253,
    new_P3_ADD_360_1242_U254, new_P3_ADD_360_1242_U255,
    new_P3_ADD_360_1242_U256, new_P3_ADD_360_1242_U257,
    new_P3_ADD_360_1242_U258, new_P3_LT_563_1260_U6, new_P3_LT_563_1260_U7,
    new_P3_SUB_589_U6, new_P3_SUB_589_U7, new_P3_SUB_589_U8,
    new_P3_SUB_589_U9, new_P3_ADD_467_U4, new_P3_ADD_467_U5,
    new_P3_ADD_467_U6, new_P3_ADD_467_U7, new_P3_ADD_467_U8,
    new_P3_ADD_467_U9, new_P3_ADD_467_U10, new_P3_ADD_467_U11,
    new_P3_ADD_467_U12, new_P3_ADD_467_U13, new_P3_ADD_467_U14,
    new_P3_ADD_467_U15, new_P3_ADD_467_U16, new_P3_ADD_467_U17,
    new_P3_ADD_467_U18, new_P3_ADD_467_U19, new_P3_ADD_467_U20,
    new_P3_ADD_467_U21, new_P3_ADD_467_U22, new_P3_ADD_467_U23,
    new_P3_ADD_467_U24, new_P3_ADD_467_U25, new_P3_ADD_467_U26,
    new_P3_ADD_467_U27, new_P3_ADD_467_U28, new_P3_ADD_467_U29,
    new_P3_ADD_467_U30, new_P3_ADD_467_U31, new_P3_ADD_467_U32,
    new_P3_ADD_467_U33, new_P3_ADD_467_U34, new_P3_ADD_467_U35,
    new_P3_ADD_467_U36, new_P3_ADD_467_U37, new_P3_ADD_467_U38,
    new_P3_ADD_467_U39, new_P3_ADD_467_U40, new_P3_ADD_467_U41,
    new_P3_ADD_467_U42, new_P3_ADD_467_U43, new_P3_ADD_467_U44,
    new_P3_ADD_467_U45, new_P3_ADD_467_U46, new_P3_ADD_467_U47,
    new_P3_ADD_467_U48, new_P3_ADD_467_U49, new_P3_ADD_467_U50,
    new_P3_ADD_467_U51, new_P3_ADD_467_U52, new_P3_ADD_467_U53,
    new_P3_ADD_467_U54, new_P3_ADD_467_U55, new_P3_ADD_467_U56,
    new_P3_ADD_467_U57, new_P3_ADD_467_U58, new_P3_ADD_467_U59,
    new_P3_ADD_467_U60, new_P3_ADD_467_U61, new_P3_ADD_467_U62,
    new_P3_ADD_467_U63, new_P3_ADD_467_U64, new_P3_ADD_467_U65,
    new_P3_ADD_467_U66, new_P3_ADD_467_U67, new_P3_ADD_467_U68,
    new_P3_ADD_467_U69, new_P3_ADD_467_U70, new_P3_ADD_467_U71,
    new_P3_ADD_467_U72, new_P3_ADD_467_U73, new_P3_ADD_467_U74,
    new_P3_ADD_467_U75, new_P3_ADD_467_U76, new_P3_ADD_467_U77,
    new_P3_ADD_467_U78, new_P3_ADD_467_U79, new_P3_ADD_467_U80,
    new_P3_ADD_467_U81, new_P3_ADD_467_U82, new_P3_ADD_467_U83,
    new_P3_ADD_467_U84, new_P3_ADD_467_U85, new_P3_ADD_467_U86,
    new_P3_ADD_467_U87, new_P3_ADD_467_U88, new_P3_ADD_467_U89,
    new_P3_ADD_467_U90, new_P3_ADD_467_U91, new_P3_ADD_467_U92,
    new_P3_ADD_467_U93, new_P3_ADD_467_U94, new_P3_ADD_467_U95,
    new_P3_ADD_467_U96, new_P3_ADD_467_U97, new_P3_ADD_467_U98,
    new_P3_ADD_467_U99, new_P3_ADD_467_U100, new_P3_ADD_467_U101,
    new_P3_ADD_467_U102, new_P3_ADD_467_U103, new_P3_ADD_467_U104,
    new_P3_ADD_467_U105, new_P3_ADD_467_U106, new_P3_ADD_467_U107,
    new_P3_ADD_467_U108, new_P3_ADD_467_U109, new_P3_ADD_467_U110,
    new_P3_ADD_467_U111, new_P3_ADD_467_U112, new_P3_ADD_467_U113,
    new_P3_ADD_467_U114, new_P3_ADD_467_U115, new_P3_ADD_467_U116,
    new_P3_ADD_467_U117, new_P3_ADD_467_U118, new_P3_ADD_467_U119,
    new_P3_ADD_467_U120, new_P3_ADD_467_U121, new_P3_ADD_467_U122,
    new_P3_ADD_467_U123, new_P3_ADD_467_U124, new_P3_ADD_467_U125,
    new_P3_ADD_467_U126, new_P3_ADD_467_U127, new_P3_ADD_467_U128,
    new_P3_ADD_467_U129, new_P3_ADD_467_U130, new_P3_ADD_467_U131,
    new_P3_ADD_467_U132, new_P3_ADD_467_U133, new_P3_ADD_467_U134,
    new_P3_ADD_467_U135, new_P3_ADD_467_U136, new_P3_ADD_467_U137,
    new_P3_ADD_467_U138, new_P3_ADD_467_U139, new_P3_ADD_467_U140,
    new_P3_ADD_467_U141, new_P3_ADD_467_U142, new_P3_ADD_467_U143,
    new_P3_ADD_467_U144, new_P3_ADD_467_U145, new_P3_ADD_467_U146,
    new_P3_ADD_467_U147, new_P3_ADD_467_U148, new_P3_ADD_467_U149,
    new_P3_ADD_467_U150, new_P3_ADD_467_U151, new_P3_ADD_467_U152,
    new_P3_ADD_467_U153, new_P3_ADD_467_U154, new_P3_ADD_467_U155,
    new_P3_ADD_467_U156, new_P3_ADD_467_U157, new_P3_ADD_467_U158,
    new_P3_ADD_467_U159, new_P3_ADD_467_U160, new_P3_ADD_467_U161,
    new_P3_ADD_467_U162, new_P3_ADD_467_U163, new_P3_ADD_467_U164,
    new_P3_ADD_467_U165, new_P3_ADD_467_U166, new_P3_ADD_467_U167,
    new_P3_ADD_467_U168, new_P3_ADD_467_U169, new_P3_ADD_467_U170,
    new_P3_ADD_467_U171, new_P3_ADD_467_U172, new_P3_ADD_467_U173,
    new_P3_ADD_467_U174, new_P3_ADD_467_U175, new_P3_ADD_467_U176,
    new_P3_ADD_467_U177, new_P3_ADD_467_U178, new_P3_ADD_467_U179,
    new_P3_ADD_467_U180, new_P3_ADD_467_U181, new_P3_ADD_467_U182,
    new_P3_ADD_430_U4, new_P3_ADD_430_U5, new_P3_ADD_430_U6,
    new_P3_ADD_430_U7, new_P3_ADD_430_U8, new_P3_ADD_430_U9,
    new_P3_ADD_430_U10, new_P3_ADD_430_U11, new_P3_ADD_430_U12,
    new_P3_ADD_430_U13, new_P3_ADD_430_U14, new_P3_ADD_430_U15,
    new_P3_ADD_430_U16, new_P3_ADD_430_U17, new_P3_ADD_430_U18,
    new_P3_ADD_430_U19, new_P3_ADD_430_U20, new_P3_ADD_430_U21,
    new_P3_ADD_430_U22, new_P3_ADD_430_U23, new_P3_ADD_430_U24,
    new_P3_ADD_430_U25, new_P3_ADD_430_U26, new_P3_ADD_430_U27,
    new_P3_ADD_430_U28, new_P3_ADD_430_U29, new_P3_ADD_430_U30,
    new_P3_ADD_430_U31, new_P3_ADD_430_U32, new_P3_ADD_430_U33,
    new_P3_ADD_430_U34, new_P3_ADD_430_U35, new_P3_ADD_430_U36,
    new_P3_ADD_430_U37, new_P3_ADD_430_U38, new_P3_ADD_430_U39,
    new_P3_ADD_430_U40, new_P3_ADD_430_U41, new_P3_ADD_430_U42,
    new_P3_ADD_430_U43, new_P3_ADD_430_U44, new_P3_ADD_430_U45,
    new_P3_ADD_430_U46, new_P3_ADD_430_U47, new_P3_ADD_430_U48,
    new_P3_ADD_430_U49, new_P3_ADD_430_U50, new_P3_ADD_430_U51,
    new_P3_ADD_430_U52, new_P3_ADD_430_U53, new_P3_ADD_430_U54,
    new_P3_ADD_430_U55, new_P3_ADD_430_U56, new_P3_ADD_430_U57,
    new_P3_ADD_430_U58, new_P3_ADD_430_U59, new_P3_ADD_430_U60,
    new_P3_ADD_430_U61, new_P3_ADD_430_U62, new_P3_ADD_430_U63,
    new_P3_ADD_430_U64, new_P3_ADD_430_U65, new_P3_ADD_430_U66,
    new_P3_ADD_430_U67, new_P3_ADD_430_U68, new_P3_ADD_430_U69,
    new_P3_ADD_430_U70, new_P3_ADD_430_U71, new_P3_ADD_430_U72,
    new_P3_ADD_430_U73, new_P3_ADD_430_U74, new_P3_ADD_430_U75,
    new_P3_ADD_430_U76, new_P3_ADD_430_U77, new_P3_ADD_430_U78,
    new_P3_ADD_430_U79, new_P3_ADD_430_U80, new_P3_ADD_430_U81,
    new_P3_ADD_430_U82, new_P3_ADD_430_U83, new_P3_ADD_430_U84,
    new_P3_ADD_430_U85, new_P3_ADD_430_U86, new_P3_ADD_430_U87,
    new_P3_ADD_430_U88, new_P3_ADD_430_U89, new_P3_ADD_430_U90,
    new_P3_ADD_430_U91, new_P3_ADD_430_U92, new_P3_ADD_430_U93,
    new_P3_ADD_430_U94, new_P3_ADD_430_U95, new_P3_ADD_430_U96,
    new_P3_ADD_430_U97, new_P3_ADD_430_U98, new_P3_ADD_430_U99,
    new_P3_ADD_430_U100, new_P3_ADD_430_U101, new_P3_ADD_430_U102,
    new_P3_ADD_430_U103, new_P3_ADD_430_U104, new_P3_ADD_430_U105,
    new_P3_ADD_430_U106, new_P3_ADD_430_U107, new_P3_ADD_430_U108,
    new_P3_ADD_430_U109, new_P3_ADD_430_U110, new_P3_ADD_430_U111,
    new_P3_ADD_430_U112, new_P3_ADD_430_U113, new_P3_ADD_430_U114,
    new_P3_ADD_430_U115, new_P3_ADD_430_U116, new_P3_ADD_430_U117,
    new_P3_ADD_430_U118, new_P3_ADD_430_U119, new_P3_ADD_430_U120,
    new_P3_ADD_430_U121, new_P3_ADD_430_U122, new_P3_ADD_430_U123,
    new_P3_ADD_430_U124, new_P3_ADD_430_U125, new_P3_ADD_430_U126,
    new_P3_ADD_430_U127, new_P3_ADD_430_U128, new_P3_ADD_430_U129,
    new_P3_ADD_430_U130, new_P3_ADD_430_U131, new_P3_ADD_430_U132,
    new_P3_ADD_430_U133, new_P3_ADD_430_U134, new_P3_ADD_430_U135,
    new_P3_ADD_430_U136, new_P3_ADD_430_U137, new_P3_ADD_430_U138,
    new_P3_ADD_430_U139, new_P3_ADD_430_U140, new_P3_ADD_430_U141,
    new_P3_ADD_430_U142, new_P3_ADD_430_U143, new_P3_ADD_430_U144,
    new_P3_ADD_430_U145, new_P3_ADD_430_U146, new_P3_ADD_430_U147,
    new_P3_ADD_430_U148, new_P3_ADD_430_U149, new_P3_ADD_430_U150,
    new_P3_ADD_430_U151, new_P3_ADD_430_U152, new_P3_ADD_430_U153,
    new_P3_ADD_430_U154, new_P3_ADD_430_U155, new_P3_ADD_430_U156,
    new_P3_ADD_430_U157, new_P3_ADD_430_U158, new_P3_ADD_430_U159,
    new_P3_ADD_430_U160, new_P3_ADD_430_U161, new_P3_ADD_430_U162,
    new_P3_ADD_430_U163, new_P3_ADD_430_U164, new_P3_ADD_430_U165,
    new_P3_ADD_430_U166, new_P3_ADD_430_U167, new_P3_ADD_430_U168,
    new_P3_ADD_430_U169, new_P3_ADD_430_U170, new_P3_ADD_430_U171,
    new_P3_ADD_430_U172, new_P3_ADD_430_U173, new_P3_ADD_430_U174,
    new_P3_ADD_430_U175, new_P3_ADD_430_U176, new_P3_ADD_430_U177,
    new_P3_ADD_430_U178, new_P3_ADD_430_U179, new_P3_ADD_430_U180,
    new_P3_ADD_430_U181, new_P3_ADD_430_U182, new_P3_ADD_380_U5,
    new_P3_ADD_380_U6, new_P3_ADD_380_U7, new_P3_ADD_380_U8,
    new_P3_ADD_380_U9, new_P3_ADD_380_U10, new_P3_ADD_380_U11,
    new_P3_ADD_380_U12, new_P3_ADD_380_U13, new_P3_ADD_380_U14,
    new_P3_ADD_380_U15, new_P3_ADD_380_U16, new_P3_ADD_380_U17,
    new_P3_ADD_380_U18, new_P3_ADD_380_U19, new_P3_ADD_380_U20,
    new_P3_ADD_380_U21, new_P3_ADD_380_U22, new_P3_ADD_380_U23,
    new_P3_ADD_380_U24, new_P3_ADD_380_U25, new_P3_ADD_380_U26,
    new_P3_ADD_380_U27, new_P3_ADD_380_U28, new_P3_ADD_380_U29,
    new_P3_ADD_380_U30, new_P3_ADD_380_U31, new_P3_ADD_380_U32,
    new_P3_ADD_380_U33, new_P3_ADD_380_U34, new_P3_ADD_380_U35,
    new_P3_ADD_380_U36, new_P3_ADD_380_U37, new_P3_ADD_380_U38,
    new_P3_ADD_380_U39, new_P3_ADD_380_U40, new_P3_ADD_380_U41,
    new_P3_ADD_380_U42, new_P3_ADD_380_U43, new_P3_ADD_380_U44,
    new_P3_ADD_380_U45, new_P3_ADD_380_U46, new_P3_ADD_380_U47,
    new_P3_ADD_380_U48, new_P3_ADD_380_U49, new_P3_ADD_380_U50,
    new_P3_ADD_380_U51, new_P3_ADD_380_U52, new_P3_ADD_380_U53,
    new_P3_ADD_380_U54, new_P3_ADD_380_U55, new_P3_ADD_380_U56,
    new_P3_ADD_380_U57, new_P3_ADD_380_U58, new_P3_ADD_380_U59,
    new_P3_ADD_380_U60, new_P3_ADD_380_U61, new_P3_ADD_380_U62,
    new_P3_ADD_380_U63, new_P3_ADD_380_U64, new_P3_ADD_380_U65,
    new_P3_ADD_380_U66, new_P3_ADD_380_U67, new_P3_ADD_380_U68,
    new_P3_ADD_380_U69, new_P3_ADD_380_U70, new_P3_ADD_380_U71,
    new_P3_ADD_380_U72, new_P3_ADD_380_U73, new_P3_ADD_380_U74,
    new_P3_ADD_380_U75, new_P3_ADD_380_U76, new_P3_ADD_380_U77,
    new_P3_ADD_380_U78, new_P3_ADD_380_U79, new_P3_ADD_380_U80,
    new_P3_ADD_380_U81, new_P3_ADD_380_U82, new_P3_ADD_380_U83,
    new_P3_ADD_380_U84, new_P3_ADD_380_U85, new_P3_ADD_380_U86,
    new_P3_ADD_380_U87, new_P3_ADD_380_U88, new_P3_ADD_380_U89,
    new_P3_ADD_380_U90, new_P3_ADD_380_U91, new_P3_ADD_380_U92,
    new_P3_ADD_380_U93, new_P3_ADD_380_U94, new_P3_ADD_380_U95,
    new_P3_ADD_380_U96, new_P3_ADD_380_U97, new_P3_ADD_380_U98,
    new_P3_ADD_380_U99, new_P3_ADD_380_U100, new_P3_ADD_380_U101,
    new_P3_ADD_380_U102, new_P3_ADD_380_U103, new_P3_ADD_380_U104,
    new_P3_ADD_380_U105, new_P3_ADD_380_U106, new_P3_ADD_380_U107,
    new_P3_ADD_380_U108, new_P3_ADD_380_U109, new_P3_ADD_380_U110,
    new_P3_ADD_380_U111, new_P3_ADD_380_U112, new_P3_ADD_380_U113,
    new_P3_ADD_380_U114, new_P3_ADD_380_U115, new_P3_ADD_380_U116,
    new_P3_ADD_380_U117, new_P3_ADD_380_U118, new_P3_ADD_380_U119,
    new_P3_ADD_380_U120, new_P3_ADD_380_U121, new_P3_ADD_380_U122,
    new_P3_ADD_380_U123, new_P3_ADD_380_U124, new_P3_ADD_380_U125,
    new_P3_ADD_380_U126, new_P3_ADD_380_U127, new_P3_ADD_380_U128,
    new_P3_ADD_380_U129, new_P3_ADD_380_U130, new_P3_ADD_380_U131,
    new_P3_ADD_380_U132, new_P3_ADD_380_U133, new_P3_ADD_380_U134,
    new_P3_ADD_380_U135, new_P3_ADD_380_U136, new_P3_ADD_380_U137,
    new_P3_ADD_380_U138, new_P3_ADD_380_U139, new_P3_ADD_380_U140,
    new_P3_ADD_380_U141, new_P3_ADD_380_U142, new_P3_ADD_380_U143,
    new_P3_ADD_380_U144, new_P3_ADD_380_U145, new_P3_ADD_380_U146,
    new_P3_ADD_380_U147, new_P3_ADD_380_U148, new_P3_ADD_380_U149,
    new_P3_ADD_380_U150, new_P3_ADD_380_U151, new_P3_ADD_380_U152,
    new_P3_ADD_380_U153, new_P3_ADD_380_U154, new_P3_ADD_380_U155,
    new_P3_ADD_380_U156, new_P3_ADD_380_U157, new_P3_ADD_380_U158,
    new_P3_ADD_380_U159, new_P3_ADD_380_U160, new_P3_ADD_380_U161,
    new_P3_ADD_380_U162, new_P3_ADD_380_U163, new_P3_ADD_380_U164,
    new_P3_ADD_380_U165, new_P3_ADD_380_U166, new_P3_ADD_380_U167,
    new_P3_ADD_380_U168, new_P3_ADD_380_U169, new_P3_ADD_380_U170,
    new_P3_ADD_380_U171, new_P3_ADD_380_U172, new_P3_ADD_380_U173,
    new_P3_ADD_380_U174, new_P3_ADD_380_U175, new_P3_ADD_380_U176,
    new_P3_ADD_380_U177, new_P3_ADD_380_U178, new_P3_ADD_380_U179,
    new_P3_ADD_380_U180, new_P3_ADD_380_U181, new_P3_ADD_380_U182,
    new_P3_ADD_380_U183, new_P3_ADD_380_U184, new_P3_ADD_380_U185,
    new_P3_ADD_380_U186, new_P3_ADD_380_U187, new_P3_ADD_380_U188,
    new_P3_ADD_380_U189, new_P3_GTE_370_U6, new_P3_GTE_370_U7,
    new_P3_GTE_370_U8, new_P3_GTE_370_U9, new_P3_ADD_344_U5,
    new_P3_ADD_344_U6, new_P3_ADD_344_U7, new_P3_ADD_344_U8,
    new_P3_ADD_344_U9, new_P3_ADD_344_U10, new_P3_ADD_344_U11,
    new_P3_ADD_344_U12, new_P3_ADD_344_U13, new_P3_ADD_344_U14,
    new_P3_ADD_344_U15, new_P3_ADD_344_U16, new_P3_ADD_344_U17,
    new_P3_ADD_344_U18, new_P3_ADD_344_U19, new_P3_ADD_344_U20,
    new_P3_ADD_344_U21, new_P3_ADD_344_U22, new_P3_ADD_344_U23,
    new_P3_ADD_344_U24, new_P3_ADD_344_U25, new_P3_ADD_344_U26,
    new_P3_ADD_344_U27, new_P3_ADD_344_U28, new_P3_ADD_344_U29,
    new_P3_ADD_344_U30, new_P3_ADD_344_U31, new_P3_ADD_344_U32,
    new_P3_ADD_344_U33, new_P3_ADD_344_U34, new_P3_ADD_344_U35,
    new_P3_ADD_344_U36, new_P3_ADD_344_U37, new_P3_ADD_344_U38,
    new_P3_ADD_344_U39, new_P3_ADD_344_U40, new_P3_ADD_344_U41,
    new_P3_ADD_344_U42, new_P3_ADD_344_U43, new_P3_ADD_344_U44,
    new_P3_ADD_344_U45, new_P3_ADD_344_U46, new_P3_ADD_344_U47,
    new_P3_ADD_344_U48, new_P3_ADD_344_U49, new_P3_ADD_344_U50,
    new_P3_ADD_344_U51, new_P3_ADD_344_U52, new_P3_ADD_344_U53,
    new_P3_ADD_344_U54, new_P3_ADD_344_U55, new_P3_ADD_344_U56,
    new_P3_ADD_344_U57, new_P3_ADD_344_U58, new_P3_ADD_344_U59,
    new_P3_ADD_344_U60, new_P3_ADD_344_U61, new_P3_ADD_344_U62,
    new_P3_ADD_344_U63, new_P3_ADD_344_U64, new_P3_ADD_344_U65,
    new_P3_ADD_344_U66, new_P3_ADD_344_U67, new_P3_ADD_344_U68,
    new_P3_ADD_344_U69, new_P3_ADD_344_U70, new_P3_ADD_344_U71,
    new_P3_ADD_344_U72, new_P3_ADD_344_U73, new_P3_ADD_344_U74,
    new_P3_ADD_344_U75, new_P3_ADD_344_U76, new_P3_ADD_344_U77,
    new_P3_ADD_344_U78, new_P3_ADD_344_U79, new_P3_ADD_344_U80,
    new_P3_ADD_344_U81, new_P3_ADD_344_U82, new_P3_ADD_344_U83,
    new_P3_ADD_344_U84, new_P3_ADD_344_U85, new_P3_ADD_344_U86,
    new_P3_ADD_344_U87, new_P3_ADD_344_U88, new_P3_ADD_344_U89,
    new_P3_ADD_344_U90, new_P3_ADD_344_U91, new_P3_ADD_344_U92,
    new_P3_ADD_344_U93, new_P3_ADD_344_U94, new_P3_ADD_344_U95,
    new_P3_ADD_344_U96, new_P3_ADD_344_U97, new_P3_ADD_344_U98,
    new_P3_ADD_344_U99, new_P3_ADD_344_U100, new_P3_ADD_344_U101,
    new_P3_ADD_344_U102, new_P3_ADD_344_U103, new_P3_ADD_344_U104,
    new_P3_ADD_344_U105, new_P3_ADD_344_U106, new_P3_ADD_344_U107,
    new_P3_ADD_344_U108, new_P3_ADD_344_U109, new_P3_ADD_344_U110,
    new_P3_ADD_344_U111, new_P3_ADD_344_U112, new_P3_ADD_344_U113,
    new_P3_ADD_344_U114, new_P3_ADD_344_U115, new_P3_ADD_344_U116,
    new_P3_ADD_344_U117, new_P3_ADD_344_U118, new_P3_ADD_344_U119,
    new_P3_ADD_344_U120, new_P3_ADD_344_U121, new_P3_ADD_344_U122,
    new_P3_ADD_344_U123, new_P3_ADD_344_U124, new_P3_ADD_344_U125,
    new_P3_ADD_344_U126, new_P3_ADD_344_U127, new_P3_ADD_344_U128,
    new_P3_ADD_344_U129, new_P3_ADD_344_U130, new_P3_ADD_344_U131,
    new_P3_ADD_344_U132, new_P3_ADD_344_U133, new_P3_ADD_344_U134,
    new_P3_ADD_344_U135, new_P3_ADD_344_U136, new_P3_ADD_344_U137,
    new_P3_ADD_344_U138, new_P3_ADD_344_U139, new_P3_ADD_344_U140,
    new_P3_ADD_344_U141, new_P3_ADD_344_U142, new_P3_ADD_344_U143,
    new_P3_ADD_344_U144, new_P3_ADD_344_U145, new_P3_ADD_344_U146,
    new_P3_ADD_344_U147, new_P3_ADD_344_U148, new_P3_ADD_344_U149,
    new_P3_ADD_344_U150, new_P3_ADD_344_U151, new_P3_ADD_344_U152,
    new_P3_ADD_344_U153, new_P3_ADD_344_U154, new_P3_ADD_344_U155,
    new_P3_ADD_344_U156, new_P3_ADD_344_U157, new_P3_ADD_344_U158,
    new_P3_ADD_344_U159, new_P3_ADD_344_U160, new_P3_ADD_344_U161,
    new_P3_ADD_344_U162, new_P3_ADD_344_U163, new_P3_ADD_344_U164,
    new_P3_ADD_344_U165, new_P3_ADD_344_U166, new_P3_ADD_344_U167,
    new_P3_ADD_344_U168, new_P3_ADD_344_U169, new_P3_ADD_344_U170,
    new_P3_ADD_344_U171, new_P3_ADD_344_U172, new_P3_ADD_344_U173,
    new_P3_ADD_344_U174, new_P3_ADD_344_U175, new_P3_ADD_344_U176,
    new_P3_ADD_344_U177, new_P3_ADD_344_U178, new_P3_ADD_344_U179,
    new_P3_ADD_344_U180, new_P3_ADD_344_U181, new_P3_ADD_344_U182,
    new_P3_ADD_344_U183, new_P3_ADD_344_U184, new_P3_ADD_344_U185,
    new_P3_ADD_344_U186, new_P3_ADD_344_U187, new_P3_ADD_344_U188,
    new_P3_ADD_344_U189, new_P3_LT_563_U6, new_P3_LT_563_U7,
    new_P3_LT_563_U8, new_P3_LT_563_U9, new_P3_LT_563_U10,
    new_P3_LT_563_U11, new_P3_LT_563_U12, new_P3_LT_563_U13,
    new_P3_LT_563_U14, new_P3_LT_563_U15, new_P3_LT_563_U16,
    new_P3_LT_563_U17, new_P3_LT_563_U18, new_P3_LT_563_U19,
    new_P3_LT_563_U20, new_P3_LT_563_U21, new_P3_LT_563_U22,
    new_P3_LT_563_U23, new_P3_LT_563_U24, new_P3_LT_563_U25,
    new_P3_LT_563_U26, new_P3_LT_563_U27, new_P3_LT_563_U28,
    new_P3_ADD_339_U4, new_P3_ADD_339_U5, new_P3_ADD_339_U6,
    new_P3_ADD_339_U7, new_P3_ADD_339_U8, new_P3_ADD_339_U9,
    new_P3_ADD_339_U10, new_P3_ADD_339_U11, new_P3_ADD_339_U12,
    new_P3_ADD_339_U13, new_P3_ADD_339_U14, new_P3_ADD_339_U15,
    new_P3_ADD_339_U16, new_P3_ADD_339_U17, new_P3_ADD_339_U18,
    new_P3_ADD_339_U19, new_P3_ADD_339_U20, new_P3_ADD_339_U21,
    new_P3_ADD_339_U22, new_P3_ADD_339_U23, new_P3_ADD_339_U24,
    new_P3_ADD_339_U25, new_P3_ADD_339_U26, new_P3_ADD_339_U27,
    new_P3_ADD_339_U28, new_P3_ADD_339_U29, new_P3_ADD_339_U30,
    new_P3_ADD_339_U31, new_P3_ADD_339_U32, new_P3_ADD_339_U33,
    new_P3_ADD_339_U34, new_P3_ADD_339_U35, new_P3_ADD_339_U36,
    new_P3_ADD_339_U37, new_P3_ADD_339_U38, new_P3_ADD_339_U39,
    new_P3_ADD_339_U40, new_P3_ADD_339_U41, new_P3_ADD_339_U42,
    new_P3_ADD_339_U43, new_P3_ADD_339_U44, new_P3_ADD_339_U45,
    new_P3_ADD_339_U46, new_P3_ADD_339_U47, new_P3_ADD_339_U48,
    new_P3_ADD_339_U49, new_P3_ADD_339_U50, new_P3_ADD_339_U51,
    new_P3_ADD_339_U52, new_P3_ADD_339_U53, new_P3_ADD_339_U54,
    new_P3_ADD_339_U55, new_P3_ADD_339_U56, new_P3_ADD_339_U57,
    new_P3_ADD_339_U58, new_P3_ADD_339_U59, new_P3_ADD_339_U60,
    new_P3_ADD_339_U61, new_P3_ADD_339_U62, new_P3_ADD_339_U63,
    new_P3_ADD_339_U64, new_P3_ADD_339_U65, new_P3_ADD_339_U66,
    new_P3_ADD_339_U67, new_P3_ADD_339_U68, new_P3_ADD_339_U69,
    new_P3_ADD_339_U70, new_P3_ADD_339_U71, new_P3_ADD_339_U72,
    new_P3_ADD_339_U73, new_P3_ADD_339_U74, new_P3_ADD_339_U75,
    new_P3_ADD_339_U76, new_P3_ADD_339_U77, new_P3_ADD_339_U78,
    new_P3_ADD_339_U79, new_P3_ADD_339_U80, new_P3_ADD_339_U81,
    new_P3_ADD_339_U82, new_P3_ADD_339_U83, new_P3_ADD_339_U84,
    new_P3_ADD_339_U85, new_P3_ADD_339_U86, new_P3_ADD_339_U87,
    new_P3_ADD_339_U88, new_P3_ADD_339_U89, new_P3_ADD_339_U90,
    new_P3_ADD_339_U91, new_P3_ADD_339_U92, new_P3_ADD_339_U93,
    new_P3_ADD_339_U94, new_P3_ADD_339_U95, new_P3_ADD_339_U96,
    new_P3_ADD_339_U97, new_P3_ADD_339_U98, new_P3_ADD_339_U99,
    new_P3_ADD_339_U100, new_P3_ADD_339_U101, new_P3_ADD_339_U102,
    new_P3_ADD_339_U103, new_P3_ADD_339_U104, new_P3_ADD_339_U105,
    new_P3_ADD_339_U106, new_P3_ADD_339_U107, new_P3_ADD_339_U108,
    new_P3_ADD_339_U109, new_P3_ADD_339_U110, new_P3_ADD_339_U111,
    new_P3_ADD_339_U112, new_P3_ADD_339_U113, new_P3_ADD_339_U114,
    new_P3_ADD_339_U115, new_P3_ADD_339_U116, new_P3_ADD_339_U117,
    new_P3_ADD_339_U118, new_P3_ADD_339_U119, new_P3_ADD_339_U120,
    new_P3_ADD_339_U121, new_P3_ADD_339_U122, new_P3_ADD_339_U123,
    new_P3_ADD_339_U124, new_P3_ADD_339_U125, new_P3_ADD_339_U126,
    new_P3_ADD_339_U127, new_P3_ADD_339_U128, new_P3_ADD_339_U129,
    new_P3_ADD_339_U130, new_P3_ADD_339_U131, new_P3_ADD_339_U132,
    new_P3_ADD_339_U133, new_P3_ADD_339_U134, new_P3_ADD_339_U135,
    new_P3_ADD_339_U136, new_P3_ADD_339_U137, new_P3_ADD_339_U138,
    new_P3_ADD_339_U139, new_P3_ADD_339_U140, new_P3_ADD_339_U141,
    new_P3_ADD_339_U142, new_P3_ADD_339_U143, new_P3_ADD_339_U144,
    new_P3_ADD_339_U145, new_P3_ADD_339_U146, new_P3_ADD_339_U147,
    new_P3_ADD_339_U148, new_P3_ADD_339_U149, new_P3_ADD_339_U150,
    new_P3_ADD_339_U151, new_P3_ADD_339_U152, new_P3_ADD_339_U153,
    new_P3_ADD_339_U154, new_P3_ADD_339_U155, new_P3_ADD_339_U156,
    new_P3_ADD_339_U157, new_P3_ADD_339_U158, new_P3_ADD_339_U159,
    new_P3_ADD_339_U160, new_P3_ADD_339_U161, new_P3_ADD_339_U162,
    new_P3_ADD_339_U163, new_P3_ADD_339_U164, new_P3_ADD_339_U165,
    new_P3_ADD_339_U166, new_P3_ADD_339_U167, new_P3_ADD_339_U168,
    new_P3_ADD_339_U169, new_P3_ADD_339_U170, new_P3_ADD_339_U171,
    new_P3_ADD_339_U172, new_P3_ADD_339_U173, new_P3_ADD_339_U174,
    new_P3_ADD_339_U175, new_P3_ADD_339_U176, new_P3_ADD_339_U177,
    new_P3_ADD_339_U178, new_P3_ADD_339_U179, new_P3_ADD_339_U180,
    new_P3_ADD_339_U181, new_P3_ADD_339_U182, new_P3_ADD_360_U4,
    new_P3_ADD_360_U5, new_P3_ADD_360_U6, new_P3_ADD_360_U7,
    new_P3_ADD_360_U8, new_P3_ADD_360_U9, new_P3_ADD_360_U10,
    new_P3_ADD_360_U11, new_P3_ADD_360_U12, new_P3_ADD_360_U13,
    new_P3_ADD_360_U14, new_P3_ADD_360_U15, new_P3_ADD_360_U16,
    new_P3_ADD_360_U17, new_P3_ADD_360_U18, new_P3_ADD_360_U19,
    new_P3_ADD_360_U20, new_P3_ADD_360_U21, new_P3_ADD_360_U22,
    new_P3_ADD_360_U23, new_P3_ADD_360_U24, new_P3_ADD_360_U25,
    new_P3_ADD_360_U26, new_P3_ADD_360_U27, new_P3_ADD_360_U28,
    new_P3_ADD_360_U29, new_P3_ADD_360_U30, new_P3_ADD_360_U31,
    new_P3_ADD_360_U32, new_P3_ADD_360_U33, new_P3_ADD_360_U34,
    new_P3_ADD_360_U35, new_P3_ADD_360_U36, new_P3_ADD_360_U37,
    new_P3_ADD_360_U38, new_P3_ADD_360_U39, new_P3_ADD_360_U40,
    new_P3_LTE_597_U6, new_P3_SUB_580_U6, new_P3_SUB_580_U7,
    new_P3_SUB_580_U8, new_P3_SUB_580_U9, new_P3_SUB_580_U10,
    new_P3_LT_589_U6, new_P3_LT_589_U7, new_P3_LT_589_U8,
    new_P3_ADD_541_U4, new_P3_ADD_541_U5, new_P3_ADD_541_U6,
    new_P3_ADD_541_U7, new_P3_ADD_541_U8, new_P3_ADD_541_U9,
    new_P3_ADD_541_U10, new_P3_ADD_541_U11, new_P3_ADD_541_U12,
    new_P3_ADD_541_U13, new_P3_ADD_541_U14, new_P3_ADD_541_U15,
    new_P3_ADD_541_U16, new_P3_ADD_541_U17, new_P3_ADD_541_U18,
    new_P3_ADD_541_U19, new_P3_ADD_541_U20, new_P3_ADD_541_U21,
    new_P3_ADD_541_U22, new_P3_ADD_541_U23, new_P3_ADD_541_U24,
    new_P3_ADD_541_U25, new_P3_ADD_541_U26, new_P3_ADD_541_U27,
    new_P3_ADD_541_U28, new_P3_ADD_541_U29, new_P3_ADD_541_U30,
    new_P3_ADD_541_U31, new_P3_ADD_541_U32, new_P3_ADD_541_U33,
    new_P3_ADD_541_U34, new_P3_ADD_541_U35, new_P3_ADD_541_U36,
    new_P3_ADD_541_U37, new_P3_ADD_541_U38, new_P3_ADD_541_U39,
    new_P3_ADD_541_U40, new_P3_ADD_541_U41, new_P3_ADD_541_U42,
    new_P3_ADD_541_U43, new_P3_ADD_541_U44, new_P3_ADD_541_U45,
    new_P3_ADD_541_U46, new_P3_ADD_541_U47, new_P3_ADD_541_U48,
    new_P3_ADD_541_U49, new_P3_ADD_541_U50, new_P3_ADD_541_U51,
    new_P3_ADD_541_U52, new_P3_ADD_541_U53, new_P3_ADD_541_U54,
    new_P3_ADD_541_U55, new_P3_ADD_541_U56, new_P3_ADD_541_U57,
    new_P3_ADD_541_U58, new_P3_ADD_541_U59, new_P3_ADD_541_U60,
    new_P3_ADD_541_U61, new_P3_ADD_541_U62, new_P3_ADD_541_U63,
    new_P3_ADD_541_U64, new_P3_ADD_541_U65, new_P3_ADD_541_U66,
    new_P3_ADD_541_U67, new_P3_ADD_541_U68, new_P3_ADD_541_U69,
    new_P3_ADD_541_U70, new_P3_ADD_541_U71, new_P3_ADD_541_U72,
    new_P3_ADD_541_U73, new_P3_ADD_541_U74, new_P3_ADD_541_U75,
    new_P3_ADD_541_U76, new_P3_ADD_541_U77, new_P3_ADD_541_U78,
    new_P3_ADD_541_U79, new_P3_ADD_541_U80, new_P3_ADD_541_U81,
    new_P3_ADD_541_U82, new_P3_ADD_541_U83, new_P3_ADD_541_U84,
    new_P3_ADD_541_U85, new_P3_ADD_541_U86, new_P3_ADD_541_U87,
    new_P3_ADD_541_U88, new_P3_ADD_541_U89, new_P3_ADD_541_U90,
    new_P3_ADD_541_U91, new_P3_ADD_541_U92, new_P3_ADD_541_U93,
    new_P3_ADD_541_U94, new_P3_ADD_541_U95, new_P3_ADD_541_U96,
    new_P3_ADD_541_U97, new_P3_ADD_541_U98, new_P3_ADD_541_U99,
    new_P3_ADD_541_U100, new_P3_ADD_541_U101, new_P3_ADD_541_U102,
    new_P3_ADD_541_U103, new_P3_ADD_541_U104, new_P3_ADD_541_U105,
    new_P3_ADD_541_U106, new_P3_ADD_541_U107, new_P3_ADD_541_U108,
    new_P3_ADD_541_U109, new_P3_ADD_541_U110, new_P3_ADD_541_U111,
    new_P3_ADD_541_U112, new_P3_ADD_541_U113, new_P3_ADD_541_U114,
    new_P3_ADD_541_U115, new_P3_ADD_541_U116, new_P3_ADD_541_U117,
    new_P3_ADD_541_U118, new_P3_ADD_541_U119, new_P3_ADD_541_U120,
    new_P3_ADD_541_U121, new_P3_ADD_541_U122, new_P3_ADD_541_U123,
    new_P3_ADD_541_U124, new_P3_ADD_541_U125, new_P3_ADD_541_U126,
    new_P3_ADD_541_U127, new_P3_ADD_541_U128, new_P3_ADD_541_U129,
    new_P3_ADD_541_U130, new_P3_ADD_541_U131, new_P3_ADD_541_U132,
    new_P3_ADD_541_U133, new_P3_ADD_541_U134, new_P3_ADD_541_U135,
    new_P3_ADD_541_U136, new_P3_ADD_541_U137, new_P3_ADD_541_U138,
    new_P3_ADD_541_U139, new_P3_ADD_541_U140, new_P3_ADD_541_U141,
    new_P3_ADD_541_U142, new_P3_ADD_541_U143, new_P3_ADD_541_U144,
    new_P3_ADD_541_U145, new_P3_ADD_541_U146, new_P3_ADD_541_U147,
    new_P3_ADD_541_U148, new_P3_ADD_541_U149, new_P3_ADD_541_U150,
    new_P3_ADD_541_U151, new_P3_ADD_541_U152, new_P3_ADD_541_U153,
    new_P3_ADD_541_U154, new_P3_ADD_541_U155, new_P3_ADD_541_U156,
    new_P3_ADD_541_U157, new_P3_ADD_541_U158, new_P3_ADD_541_U159,
    new_P3_ADD_541_U160, new_P3_ADD_541_U161, new_P3_ADD_541_U162,
    new_P3_ADD_541_U163, new_P3_ADD_541_U164, new_P3_ADD_541_U165,
    new_P3_ADD_541_U166, new_P3_ADD_541_U167, new_P3_ADD_541_U168,
    new_P3_ADD_541_U169, new_P3_ADD_541_U170, new_P3_ADD_541_U171,
    new_P3_ADD_541_U172, new_P3_ADD_541_U173, new_P3_ADD_541_U174,
    new_P3_ADD_541_U175, new_P3_ADD_541_U176, new_P3_ADD_541_U177,
    new_P3_ADD_541_U178, new_P3_ADD_541_U179, new_P3_ADD_541_U180,
    new_P3_ADD_541_U181, new_P3_ADD_541_U182, new_P3_SUB_355_U6,
    new_P3_SUB_355_U7, new_P3_SUB_355_U8, new_P3_SUB_355_U9,
    new_P3_SUB_355_U10, new_P3_SUB_355_U11, new_P3_SUB_355_U12,
    new_P3_SUB_355_U13, new_P3_SUB_355_U14, new_P3_SUB_355_U15,
    new_P3_SUB_355_U16, new_P3_SUB_355_U17, new_P3_SUB_355_U18,
    new_P3_SUB_355_U19, new_P3_SUB_355_U20, new_P3_SUB_355_U21,
    new_P3_SUB_355_U22, new_P3_SUB_355_U23, new_P3_SUB_355_U24,
    new_P3_SUB_355_U25, new_P3_SUB_355_U26, new_P3_SUB_355_U27,
    new_P3_SUB_355_U28, new_P3_SUB_355_U29, new_P3_SUB_355_U30,
    new_P3_SUB_355_U31, new_P3_SUB_355_U32, new_P3_SUB_355_U33,
    new_P3_SUB_355_U34, new_P3_SUB_355_U35, new_P3_SUB_355_U36,
    new_P3_SUB_355_U37, new_P3_SUB_355_U38, new_P3_SUB_355_U39,
    new_P3_SUB_355_U40, new_P3_SUB_355_U41, new_P3_SUB_355_U42,
    new_P3_SUB_355_U43, new_P3_SUB_355_U44, new_P3_SUB_355_U45,
    new_P3_SUB_355_U46, new_P3_SUB_355_U47, new_P3_SUB_355_U48,
    new_P3_SUB_355_U49, new_P3_SUB_355_U50, new_P3_SUB_355_U51,
    new_P3_SUB_355_U52, new_P3_SUB_355_U53, new_P3_SUB_355_U54,
    new_P3_SUB_355_U55, new_P3_SUB_355_U56, new_P3_SUB_355_U57,
    new_P3_SUB_355_U58, new_P3_SUB_355_U59, new_P3_SUB_355_U60,
    new_P3_SUB_355_U61, new_P3_SUB_355_U62, new_P3_SUB_355_U63,
    new_P3_SUB_355_U64, new_P3_SUB_355_U65, new_P3_SUB_355_U66,
    new_P3_SUB_450_U6, new_P3_SUB_450_U7, new_P3_SUB_450_U8,
    new_P3_SUB_450_U9, new_P3_SUB_450_U10, new_P3_SUB_450_U11,
    new_P3_SUB_450_U12, new_P3_SUB_450_U13, new_P3_SUB_450_U14,
    new_P3_SUB_450_U15, new_P3_SUB_450_U16, new_P3_SUB_450_U17,
    new_P3_SUB_450_U18, new_P3_SUB_450_U19, new_P3_SUB_450_U20,
    new_P3_SUB_450_U21, new_P3_SUB_450_U22, new_P3_SUB_450_U23,
    new_P3_SUB_450_U24, new_P3_SUB_450_U25, new_P3_SUB_450_U26,
    new_P3_SUB_450_U27, new_P3_SUB_450_U28, new_P3_SUB_450_U29,
    new_P3_SUB_450_U30, new_P3_SUB_450_U31, new_P3_SUB_450_U32,
    new_P3_SUB_450_U33, new_P3_SUB_450_U34, new_P3_SUB_450_U35,
    new_P3_SUB_450_U36, new_P3_SUB_450_U37, new_P3_SUB_450_U38,
    new_P3_SUB_450_U39, new_P3_SUB_450_U40, new_P3_SUB_450_U41,
    new_P3_SUB_450_U42, new_P3_SUB_450_U43, new_P3_SUB_450_U44,
    new_P3_SUB_450_U45, new_P3_SUB_450_U46, new_P3_SUB_450_U47,
    new_P3_SUB_450_U48, new_P3_SUB_450_U49, new_P3_SUB_450_U50,
    new_P3_SUB_450_U51, new_P3_SUB_450_U52, new_P3_SUB_450_U53,
    new_P3_SUB_450_U54, new_P3_SUB_450_U55, new_P3_SUB_450_U56,
    new_P3_SUB_450_U57, new_P3_SUB_450_U58, new_P3_SUB_450_U59,
    new_P3_SUB_450_U60, new_P3_SUB_450_U61, new_P3_SUB_450_U62,
    new_P3_SUB_450_U63, new_P3_SUB_357_1258_U4, new_P3_SUB_357_1258_U5,
    new_P3_SUB_357_1258_U6, new_P3_SUB_357_1258_U7, new_P3_SUB_357_1258_U8,
    new_P3_SUB_357_1258_U9, new_P3_SUB_357_1258_U10,
    new_P3_SUB_357_1258_U11, new_P3_SUB_357_1258_U12,
    new_P3_SUB_357_1258_U13, new_P3_SUB_357_1258_U14,
    new_P3_SUB_357_1258_U15, new_P3_SUB_357_1258_U16,
    new_P3_SUB_357_1258_U17, new_P3_SUB_357_1258_U18,
    new_P3_SUB_357_1258_U19, new_P3_SUB_357_1258_U20,
    new_P3_SUB_357_1258_U21, new_P3_SUB_357_1258_U22,
    new_P3_SUB_357_1258_U23, new_P3_SUB_357_1258_U24,
    new_P3_SUB_357_1258_U25, new_P3_SUB_357_1258_U26,
    new_P3_SUB_357_1258_U27, new_P3_SUB_357_1258_U28,
    new_P3_SUB_357_1258_U29, new_P3_SUB_357_1258_U30,
    new_P3_SUB_357_1258_U31, new_P3_SUB_357_1258_U32,
    new_P3_SUB_357_1258_U33, new_P3_SUB_357_1258_U34,
    new_P3_SUB_357_1258_U35, new_P3_SUB_357_1258_U36,
    new_P3_SUB_357_1258_U37, new_P3_SUB_357_1258_U38,
    new_P3_SUB_357_1258_U39, new_P3_SUB_357_1258_U40,
    new_P3_SUB_357_1258_U41, new_P3_SUB_357_1258_U42,
    new_P3_SUB_357_1258_U43, new_P3_SUB_357_1258_U44,
    new_P3_SUB_357_1258_U45, new_P3_SUB_357_1258_U46,
    new_P3_SUB_357_1258_U47, new_P3_SUB_357_1258_U48,
    new_P3_SUB_357_1258_U49, new_P3_SUB_357_1258_U50,
    new_P3_SUB_357_1258_U51, new_P3_SUB_357_1258_U52,
    new_P3_SUB_357_1258_U53, new_P3_SUB_357_1258_U54,
    new_P3_SUB_357_1258_U55, new_P3_SUB_357_1258_U56,
    new_P3_SUB_357_1258_U57, new_P3_SUB_357_1258_U58,
    new_P3_SUB_357_1258_U59, new_P3_SUB_357_1258_U60,
    new_P3_SUB_357_1258_U61, new_P3_SUB_357_1258_U62,
    new_P3_SUB_357_1258_U63, new_P3_SUB_357_1258_U64,
    new_P3_SUB_357_1258_U65, new_P3_SUB_357_1258_U66,
    new_P3_SUB_357_1258_U67, new_P3_SUB_357_1258_U68,
    new_P3_SUB_357_1258_U69, new_P3_SUB_357_1258_U70,
    new_P3_SUB_357_1258_U71, new_P3_SUB_357_1258_U72,
    new_P3_SUB_357_1258_U73, new_P3_SUB_357_1258_U74,
    new_P3_SUB_357_1258_U75, new_P3_SUB_357_1258_U76,
    new_P3_SUB_357_1258_U77, new_P3_SUB_357_1258_U78,
    new_P3_SUB_357_1258_U79, new_P3_SUB_357_1258_U80,
    new_P3_SUB_357_1258_U81, new_P3_SUB_357_1258_U82,
    new_P3_SUB_357_1258_U83, new_P3_SUB_357_1258_U84,
    new_P3_SUB_357_1258_U85, new_P3_SUB_357_1258_U86,
    new_P3_SUB_357_1258_U87, new_P3_SUB_357_1258_U88,
    new_P3_SUB_357_1258_U89, new_P3_SUB_357_1258_U90,
    new_P3_SUB_357_1258_U91, new_P3_SUB_357_1258_U92,
    new_P3_SUB_357_1258_U93, new_P3_SUB_357_1258_U94,
    new_P3_SUB_357_1258_U95, new_P3_SUB_357_1258_U96,
    new_P3_SUB_357_1258_U97, new_P3_SUB_357_1258_U98,
    new_P3_SUB_357_1258_U99, new_P3_SUB_357_1258_U100,
    new_P3_SUB_357_1258_U101, new_P3_SUB_357_1258_U102,
    new_P3_SUB_357_1258_U103, new_P3_SUB_357_1258_U104,
    new_P3_SUB_357_1258_U105, new_P3_SUB_357_1258_U106,
    new_P3_SUB_357_1258_U107, new_P3_SUB_357_1258_U108,
    new_P3_SUB_357_1258_U109, new_P3_SUB_357_1258_U110,
    new_P3_SUB_357_1258_U111, new_P3_SUB_357_1258_U112,
    new_P3_SUB_357_1258_U113, new_P3_SUB_357_1258_U114,
    new_P3_SUB_357_1258_U115, new_P3_SUB_357_1258_U116,
    new_P3_SUB_357_1258_U117, new_P3_SUB_357_1258_U118,
    new_P3_SUB_357_1258_U119, new_P3_SUB_357_1258_U120,
    new_P3_SUB_357_1258_U121, new_P3_SUB_357_1258_U122,
    new_P3_SUB_357_1258_U123, new_P3_SUB_357_1258_U124,
    new_P3_SUB_357_1258_U125, new_P3_SUB_357_1258_U126,
    new_P3_SUB_357_1258_U127, new_P3_SUB_357_1258_U128,
    new_P3_SUB_357_1258_U129, new_P3_SUB_357_1258_U130,
    new_P3_SUB_357_1258_U131, new_P3_SUB_357_1258_U132,
    new_P3_SUB_357_1258_U133, new_P3_SUB_357_1258_U134,
    new_P3_SUB_357_1258_U135, new_P3_SUB_357_1258_U136,
    new_P3_SUB_357_1258_U137, new_P3_SUB_357_1258_U138,
    new_P3_SUB_357_1258_U139, new_P3_SUB_357_1258_U140,
    new_P3_SUB_357_1258_U141, new_P3_SUB_357_1258_U142,
    new_P3_SUB_357_1258_U143, new_P3_SUB_357_1258_U144,
    new_P3_SUB_357_1258_U145, new_P3_SUB_357_1258_U146,
    new_P3_SUB_357_1258_U147, new_P3_SUB_357_1258_U148,
    new_P3_SUB_357_1258_U149, new_P3_SUB_357_1258_U150,
    new_P3_SUB_357_1258_U151, new_P3_SUB_357_1258_U152,
    new_P3_SUB_357_1258_U153, new_P3_SUB_357_1258_U154,
    new_P3_SUB_357_1258_U155, new_P3_SUB_357_1258_U156,
    new_P3_SUB_357_1258_U157, new_P3_SUB_357_1258_U158,
    new_P3_SUB_357_1258_U159, new_P3_SUB_357_1258_U160,
    new_P3_SUB_357_1258_U161, new_P3_SUB_357_1258_U162,
    new_P3_SUB_357_1258_U163, new_P3_SUB_357_1258_U164,
    new_P3_SUB_357_1258_U165, new_P3_SUB_357_1258_U166,
    new_P3_SUB_357_1258_U167, new_P3_SUB_357_1258_U168,
    new_P3_SUB_357_1258_U169, new_P3_SUB_357_1258_U170,
    new_P3_SUB_357_1258_U171, new_P3_SUB_357_1258_U172,
    new_P3_SUB_357_1258_U173, new_P3_SUB_357_1258_U174,
    new_P3_SUB_357_1258_U175, new_P3_SUB_357_1258_U176,
    new_P3_SUB_357_1258_U177, new_P3_SUB_357_1258_U178,
    new_P3_SUB_357_1258_U179, new_P3_SUB_357_1258_U180,
    new_P3_SUB_357_1258_U181, new_P3_SUB_357_1258_U182,
    new_P3_SUB_357_1258_U183, new_P3_SUB_357_1258_U184,
    new_P3_SUB_357_1258_U185, new_P3_SUB_357_1258_U186,
    new_P3_SUB_357_1258_U187, new_P3_SUB_357_1258_U188,
    new_P3_SUB_357_1258_U189, new_P3_SUB_357_1258_U190,
    new_P3_SUB_357_1258_U191, new_P3_SUB_357_1258_U192,
    new_P3_SUB_357_1258_U193, new_P3_SUB_357_1258_U194,
    new_P3_SUB_357_1258_U195, new_P3_SUB_357_1258_U196,
    new_P3_SUB_357_1258_U197, new_P3_SUB_357_1258_U198,
    new_P3_SUB_357_1258_U199, new_P3_SUB_357_1258_U200,
    new_P3_SUB_357_1258_U201, new_P3_SUB_357_1258_U202,
    new_P3_SUB_357_1258_U203, new_P3_SUB_357_1258_U204,
    new_P3_SUB_357_1258_U205, new_P3_SUB_357_1258_U206,
    new_P3_SUB_357_1258_U207, new_P3_SUB_357_1258_U208,
    new_P3_SUB_357_1258_U209, new_P3_SUB_357_1258_U210,
    new_P3_SUB_357_1258_U211, new_P3_SUB_357_1258_U212,
    new_P3_SUB_357_1258_U213, new_P3_SUB_357_1258_U214,
    new_P3_SUB_357_1258_U215, new_P3_SUB_357_1258_U216,
    new_P3_SUB_357_1258_U217, new_P3_SUB_357_1258_U218,
    new_P3_SUB_357_1258_U219, new_P3_SUB_357_1258_U220,
    new_P3_SUB_357_1258_U221, new_P3_SUB_357_1258_U222,
    new_P3_SUB_357_1258_U223, new_P3_SUB_357_1258_U224,
    new_P3_SUB_357_1258_U225, new_P3_SUB_357_1258_U226,
    new_P3_SUB_357_1258_U227, new_P3_SUB_357_1258_U228,
    new_P3_SUB_357_1258_U229, new_P3_SUB_357_1258_U230,
    new_P3_SUB_357_1258_U231, new_P3_SUB_357_1258_U232,
    new_P3_SUB_357_1258_U233, new_P3_SUB_357_1258_U234,
    new_P3_SUB_357_1258_U235, new_P3_SUB_357_1258_U236,
    new_P3_SUB_357_1258_U237, new_P3_SUB_357_1258_U238,
    new_P3_SUB_357_1258_U239, new_P3_SUB_357_1258_U240,
    new_P3_SUB_357_1258_U241, new_P3_SUB_357_1258_U242,
    new_P3_SUB_357_1258_U243, new_P3_SUB_357_1258_U244,
    new_P3_SUB_357_1258_U245, new_P3_SUB_357_1258_U246,
    new_P3_SUB_357_1258_U247, new_P3_SUB_357_1258_U248,
    new_P3_SUB_357_1258_U249, new_P3_SUB_357_1258_U250,
    new_P3_SUB_357_1258_U251, new_P3_SUB_357_1258_U252,
    new_P3_SUB_357_1258_U253, new_P3_SUB_357_1258_U254,
    new_P3_SUB_357_1258_U255, new_P3_SUB_357_1258_U256,
    new_P3_SUB_357_1258_U257, new_P3_SUB_357_1258_U258,
    new_P3_SUB_357_1258_U259, new_P3_SUB_357_1258_U260,
    new_P3_SUB_357_1258_U261, new_P3_SUB_357_1258_U262,
    new_P3_SUB_357_1258_U263, new_P3_SUB_357_1258_U264,
    new_P3_SUB_357_1258_U265, new_P3_SUB_357_1258_U266,
    new_P3_SUB_357_1258_U267, new_P3_SUB_357_1258_U268,
    new_P3_SUB_357_1258_U269, new_P3_SUB_357_1258_U270,
    new_P3_SUB_357_1258_U271, new_P3_SUB_357_1258_U272,
    new_P3_SUB_357_1258_U273, new_P3_SUB_357_1258_U274,
    new_P3_SUB_357_1258_U275, new_P3_SUB_357_1258_U276,
    new_P3_SUB_357_1258_U277, new_P3_SUB_357_1258_U278,
    new_P3_SUB_357_1258_U279, new_P3_SUB_357_1258_U280,
    new_P3_SUB_357_1258_U281, new_P3_SUB_357_1258_U282,
    new_P3_SUB_357_1258_U283, new_P3_SUB_357_1258_U284,
    new_P3_SUB_357_1258_U285, new_P3_SUB_357_1258_U286,
    new_P3_SUB_357_1258_U287, new_P3_SUB_357_1258_U288,
    new_P3_SUB_357_1258_U289, new_P3_SUB_357_1258_U290,
    new_P3_SUB_357_1258_U291, new_P3_SUB_357_1258_U292,
    new_P3_SUB_357_1258_U293, new_P3_SUB_357_1258_U294,
    new_P3_SUB_357_1258_U295, new_P3_SUB_357_1258_U296,
    new_P3_SUB_357_1258_U297, new_P3_SUB_357_1258_U298,
    new_P3_SUB_357_1258_U299, new_P3_SUB_357_1258_U300,
    new_P3_SUB_357_1258_U301, new_P3_SUB_357_1258_U302,
    new_P3_SUB_357_1258_U303, new_P3_SUB_357_1258_U304,
    new_P3_SUB_357_1258_U305, new_P3_SUB_357_1258_U306,
    new_P3_SUB_357_1258_U307, new_P3_SUB_357_1258_U308,
    new_P3_SUB_357_1258_U309, new_P3_SUB_357_1258_U310,
    new_P3_SUB_357_1258_U311, new_P3_SUB_357_1258_U312,
    new_P3_SUB_357_1258_U313, new_P3_SUB_357_1258_U314,
    new_P3_SUB_357_1258_U315, new_P3_SUB_357_1258_U316,
    new_P3_SUB_357_1258_U317, new_P3_SUB_357_1258_U318,
    new_P3_SUB_357_1258_U319, new_P3_SUB_357_1258_U320,
    new_P3_SUB_357_1258_U321, new_P3_SUB_357_1258_U322,
    new_P3_SUB_357_1258_U323, new_P3_SUB_357_1258_U324,
    new_P3_SUB_357_1258_U325, new_P3_SUB_357_1258_U326,
    new_P3_SUB_357_1258_U327, new_P3_SUB_357_1258_U328,
    new_P3_SUB_357_1258_U329, new_P3_SUB_357_1258_U330,
    new_P3_SUB_357_1258_U331, new_P3_SUB_357_1258_U332,
    new_P3_SUB_357_1258_U333, new_P3_SUB_357_1258_U334,
    new_P3_SUB_357_1258_U335, new_P3_SUB_357_1258_U336,
    new_P3_SUB_357_1258_U337, new_P3_SUB_357_1258_U338,
    new_P3_SUB_357_1258_U339, new_P3_SUB_357_1258_U340,
    new_P3_SUB_357_1258_U341, new_P3_SUB_357_1258_U342,
    new_P3_SUB_357_1258_U343, new_P3_SUB_357_1258_U344,
    new_P3_SUB_357_1258_U345, new_P3_SUB_357_1258_U346,
    new_P3_SUB_357_1258_U347, new_P3_SUB_357_1258_U348,
    new_P3_SUB_357_1258_U349, new_P3_SUB_357_1258_U350,
    new_P3_SUB_357_1258_U351, new_P3_SUB_357_1258_U352,
    new_P3_SUB_357_1258_U353, new_P3_SUB_357_1258_U354,
    new_P3_SUB_357_1258_U355, new_P3_SUB_357_1258_U356,
    new_P3_SUB_357_1258_U357, new_P3_SUB_357_1258_U358,
    new_P3_SUB_357_1258_U359, new_P3_SUB_357_1258_U360,
    new_P3_SUB_357_1258_U361, new_P3_SUB_357_1258_U362,
    new_P3_SUB_357_1258_U363, new_P3_SUB_357_1258_U364,
    new_P3_SUB_357_1258_U365, new_P3_SUB_357_1258_U366,
    new_P3_SUB_357_1258_U367, new_P3_SUB_357_1258_U368,
    new_P3_SUB_357_1258_U369, new_P3_SUB_357_1258_U370,
    new_P3_SUB_357_1258_U371, new_P3_SUB_357_1258_U372,
    new_P3_SUB_357_1258_U373, new_P3_SUB_357_1258_U374,
    new_P3_SUB_357_1258_U375, new_P3_SUB_357_1258_U376,
    new_P3_SUB_357_1258_U377, new_P3_SUB_357_1258_U378,
    new_P3_SUB_357_1258_U379, new_P3_SUB_357_1258_U380,
    new_P3_SUB_357_1258_U381, new_P3_SUB_357_1258_U382,
    new_P3_SUB_357_1258_U383, new_P3_SUB_357_1258_U384,
    new_P3_SUB_357_1258_U385, new_P3_SUB_357_1258_U386,
    new_P3_SUB_357_1258_U387, new_P3_SUB_357_1258_U388,
    new_P3_SUB_357_1258_U389, new_P3_SUB_357_1258_U390,
    new_P3_SUB_357_1258_U391, new_P3_SUB_357_1258_U392,
    new_P3_SUB_357_1258_U393, new_P3_SUB_357_1258_U394,
    new_P3_SUB_357_1258_U395, new_P3_SUB_357_1258_U396,
    new_P3_SUB_357_1258_U397, new_P3_SUB_357_1258_U398,
    new_P3_SUB_357_1258_U399, new_P3_SUB_357_1258_U400,
    new_P3_SUB_357_1258_U401, new_P3_SUB_357_1258_U402,
    new_P3_SUB_357_1258_U403, new_P3_SUB_357_1258_U404,
    new_P3_SUB_357_1258_U405, new_P3_SUB_357_1258_U406,
    new_P3_SUB_357_1258_U407, new_P3_SUB_357_1258_U408,
    new_P3_SUB_357_1258_U409, new_P3_SUB_357_1258_U410,
    new_P3_SUB_357_1258_U411, new_P3_SUB_357_1258_U412,
    new_P3_SUB_357_1258_U413, new_P3_SUB_357_1258_U414,
    new_P3_SUB_357_1258_U415, new_P3_SUB_357_1258_U416,
    new_P3_SUB_357_1258_U417, new_P3_SUB_357_1258_U418,
    new_P3_SUB_357_1258_U419, new_P3_SUB_357_1258_U420,
    new_P3_SUB_357_1258_U421, new_P3_SUB_357_1258_U422,
    new_P3_SUB_357_1258_U423, new_P3_SUB_357_1258_U424,
    new_P3_SUB_357_1258_U425, new_P3_SUB_357_1258_U426,
    new_P3_SUB_357_1258_U427, new_P3_SUB_357_1258_U428,
    new_P3_SUB_357_1258_U429, new_P3_SUB_357_1258_U430,
    new_P3_SUB_357_1258_U431, new_P3_SUB_357_1258_U432,
    new_P3_SUB_357_1258_U433, new_P3_SUB_357_1258_U434,
    new_P3_SUB_357_1258_U435, new_P3_SUB_357_1258_U436,
    new_P3_SUB_357_1258_U437, new_P3_SUB_357_1258_U438,
    new_P3_SUB_357_1258_U439, new_P3_SUB_357_1258_U440,
    new_P3_SUB_357_1258_U441, new_P3_SUB_357_1258_U442,
    new_P3_SUB_357_1258_U443, new_P3_SUB_357_1258_U444,
    new_P3_SUB_357_1258_U445, new_P3_SUB_357_1258_U446,
    new_P3_SUB_357_1258_U447, new_P3_SUB_357_1258_U448,
    new_P3_SUB_357_1258_U449, new_P3_SUB_357_1258_U450,
    new_P3_SUB_357_1258_U451, new_P3_SUB_357_1258_U452,
    new_P3_SUB_357_1258_U453, new_P3_SUB_357_1258_U454,
    new_P3_SUB_357_1258_U455, new_P3_SUB_357_1258_U456,
    new_P3_SUB_357_1258_U457, new_P3_SUB_357_1258_U458,
    new_P3_SUB_357_1258_U459, new_P3_SUB_357_1258_U460,
    new_P3_SUB_357_1258_U461, new_P3_SUB_357_1258_U462,
    new_P3_SUB_357_1258_U463, new_P3_SUB_357_1258_U464,
    new_P3_SUB_357_1258_U465, new_P3_SUB_357_1258_U466,
    new_P3_SUB_357_1258_U467, new_P3_SUB_357_1258_U468,
    new_P3_SUB_357_1258_U469, new_P3_SUB_357_1258_U470,
    new_P3_SUB_357_1258_U471, new_P3_SUB_357_1258_U472,
    new_P3_SUB_357_1258_U473, new_P3_SUB_357_1258_U474,
    new_P3_SUB_357_1258_U475, new_P3_SUB_357_1258_U476,
    new_P3_SUB_357_1258_U477, new_P3_SUB_357_1258_U478,
    new_P3_SUB_357_1258_U479, new_P3_SUB_357_1258_U480,
    new_P3_SUB_357_1258_U481, new_P3_SUB_357_1258_U482,
    new_P3_SUB_357_1258_U483, new_P3_SUB_357_1258_U484, new_P3_ADD_486_U5,
    new_P3_ADD_486_U6, new_P3_ADD_486_U7, new_P3_ADD_486_U8,
    new_P3_ADD_486_U9, new_P3_ADD_486_U10, new_P3_ADD_486_U11,
    new_P3_ADD_486_U12, new_P3_ADD_486_U13, new_P3_ADD_486_U14,
    new_P3_ADD_486_U15, new_P3_ADD_486_U16, new_P3_ADD_486_U17,
    new_P3_ADD_486_U18, new_P3_ADD_486_U19, new_P3_ADD_486_U20,
    new_P3_ADD_486_U21, new_P3_ADD_486_U22, new_P3_ADD_486_U23,
    new_P3_ADD_486_U24, new_P3_ADD_486_U25, new_P3_ADD_486_U26,
    new_P3_ADD_486_U27, new_P3_ADD_486_U28, new_P3_SUB_485_U6,
    new_P3_SUB_485_U7, new_P3_SUB_485_U8, new_P3_SUB_485_U9,
    new_P3_SUB_485_U10, new_P3_SUB_485_U11, new_P3_SUB_485_U12,
    new_P3_SUB_485_U13, new_P3_SUB_485_U14, new_P3_SUB_485_U15,
    new_P3_SUB_485_U16, new_P3_SUB_485_U17, new_P3_SUB_485_U18,
    new_P3_SUB_485_U19, new_P3_SUB_485_U20, new_P3_SUB_485_U21,
    new_P3_SUB_485_U22, new_P3_SUB_485_U23, new_P3_SUB_485_U24,
    new_P3_SUB_485_U25, new_P3_SUB_485_U26, new_P3_SUB_485_U27,
    new_P3_SUB_485_U28, new_P3_SUB_485_U29, new_P3_SUB_485_U30,
    new_P3_SUB_485_U31, new_P3_SUB_485_U32, new_P3_SUB_485_U33,
    new_P3_SUB_485_U34, new_P3_SUB_485_U35, new_P3_SUB_485_U36,
    new_P3_SUB_485_U37, new_P3_SUB_485_U38, new_P3_SUB_485_U39,
    new_P3_SUB_485_U40, new_P3_SUB_485_U41, new_P3_SUB_485_U42,
    new_P3_SUB_485_U43, new_P3_SUB_485_U44, new_P3_SUB_485_U45,
    new_P3_SUB_485_U46, new_P3_SUB_485_U47, new_P3_SUB_485_U48,
    new_P3_SUB_485_U49, new_P3_SUB_485_U50, new_P3_SUB_485_U51,
    new_P3_SUB_485_U52, new_P3_SUB_485_U53, new_P3_SUB_485_U54,
    new_P3_SUB_485_U55, new_P3_SUB_485_U56, new_P3_SUB_485_U57,
    new_P3_SUB_485_U58, new_P3_SUB_485_U59, new_P3_SUB_485_U60,
    new_P3_SUB_485_U61, new_P3_SUB_485_U62, new_P3_SUB_485_U63,
    new_P3_SUB_563_U6, new_P3_SUB_563_U7, new_P3_ADD_515_U4,
    new_P3_ADD_515_U5, new_P3_ADD_515_U6, new_P3_ADD_515_U7,
    new_P3_ADD_515_U8, new_P3_ADD_515_U9, new_P3_ADD_515_U10,
    new_P3_ADD_515_U11, new_P3_ADD_515_U12, new_P3_ADD_515_U13,
    new_P3_ADD_515_U14, new_P3_ADD_515_U15, new_P3_ADD_515_U16,
    new_P3_ADD_515_U17, new_P3_ADD_515_U18, new_P3_ADD_515_U19,
    new_P3_ADD_515_U20, new_P3_ADD_515_U21, new_P3_ADD_515_U22,
    new_P3_ADD_515_U23, new_P3_ADD_515_U24, new_P3_ADD_515_U25,
    new_P3_ADD_515_U26, new_P3_ADD_515_U27, new_P3_ADD_515_U28,
    new_P3_ADD_515_U29, new_P3_ADD_515_U30, new_P3_ADD_515_U31,
    new_P3_ADD_515_U32, new_P3_ADD_515_U33, new_P3_ADD_515_U34,
    new_P3_ADD_515_U35, new_P3_ADD_515_U36, new_P3_ADD_515_U37,
    new_P3_ADD_515_U38, new_P3_ADD_515_U39, new_P3_ADD_515_U40,
    new_P3_ADD_515_U41, new_P3_ADD_515_U42, new_P3_ADD_515_U43,
    new_P3_ADD_515_U44, new_P3_ADD_515_U45, new_P3_ADD_515_U46,
    new_P3_ADD_515_U47, new_P3_ADD_515_U48, new_P3_ADD_515_U49,
    new_P3_ADD_515_U50, new_P3_ADD_515_U51, new_P3_ADD_515_U52,
    new_P3_ADD_515_U53, new_P3_ADD_515_U54, new_P3_ADD_515_U55,
    new_P3_ADD_515_U56, new_P3_ADD_515_U57, new_P3_ADD_515_U58,
    new_P3_ADD_515_U59, new_P3_ADD_515_U60, new_P3_ADD_515_U61,
    new_P3_ADD_515_U62, new_P3_ADD_515_U63, new_P3_ADD_515_U64,
    new_P3_ADD_515_U65, new_P3_ADD_515_U66, new_P3_ADD_515_U67,
    new_P3_ADD_515_U68, new_P3_ADD_515_U69, new_P3_ADD_515_U70,
    new_P3_ADD_515_U71, new_P3_ADD_515_U72, new_P3_ADD_515_U73,
    new_P3_ADD_515_U74, new_P3_ADD_515_U75, new_P3_ADD_515_U76,
    new_P3_ADD_515_U77, new_P3_ADD_515_U78, new_P3_ADD_515_U79,
    new_P3_ADD_515_U80, new_P3_ADD_515_U81, new_P3_ADD_515_U82,
    new_P3_ADD_515_U83, new_P3_ADD_515_U84, new_P3_ADD_515_U85,
    new_P3_ADD_515_U86, new_P3_ADD_515_U87, new_P3_ADD_515_U88,
    new_P3_ADD_515_U89, new_P3_ADD_515_U90, new_P3_ADD_515_U91,
    new_P3_ADD_515_U92, new_P3_ADD_515_U93, new_P3_ADD_515_U94,
    new_P3_ADD_515_U95, new_P3_ADD_515_U96, new_P3_ADD_515_U97,
    new_P3_ADD_515_U98, new_P3_ADD_515_U99, new_P3_ADD_515_U100,
    new_P3_ADD_515_U101, new_P3_ADD_515_U102, new_P3_ADD_515_U103,
    new_P3_ADD_515_U104, new_P3_ADD_515_U105, new_P3_ADD_515_U106,
    new_P3_ADD_515_U107, new_P3_ADD_515_U108, new_P3_ADD_515_U109,
    new_P3_ADD_515_U110, new_P3_ADD_515_U111, new_P3_ADD_515_U112,
    new_P3_ADD_515_U113, new_P3_ADD_515_U114, new_P3_ADD_515_U115,
    new_P3_ADD_515_U116, new_P3_ADD_515_U117, new_P3_ADD_515_U118,
    new_P3_ADD_515_U119, new_P3_ADD_515_U120, new_P3_ADD_515_U121,
    new_P3_ADD_515_U122, new_P3_ADD_515_U123, new_P3_ADD_515_U124,
    new_P3_ADD_515_U125, new_P3_ADD_515_U126, new_P3_ADD_515_U127,
    new_P3_ADD_515_U128, new_P3_ADD_515_U129, new_P3_ADD_515_U130,
    new_P3_ADD_515_U131, new_P3_ADD_515_U132, new_P3_ADD_515_U133,
    new_P3_ADD_515_U134, new_P3_ADD_515_U135, new_P3_ADD_515_U136,
    new_P3_ADD_515_U137, new_P3_ADD_515_U138, new_P3_ADD_515_U139,
    new_P3_ADD_515_U140, new_P3_ADD_515_U141, new_P3_ADD_515_U142,
    new_P3_ADD_515_U143, new_P3_ADD_515_U144, new_P3_ADD_515_U145,
    new_P3_ADD_515_U146, new_P3_ADD_515_U147, new_P3_ADD_515_U148,
    new_P3_ADD_515_U149, new_P3_ADD_515_U150, new_P3_ADD_515_U151,
    new_P3_ADD_515_U152, new_P3_ADD_515_U153, new_P3_ADD_515_U154,
    new_P3_ADD_515_U155, new_P3_ADD_515_U156, new_P3_ADD_515_U157,
    new_P3_ADD_515_U158, new_P3_ADD_515_U159, new_P3_ADD_515_U160,
    new_P3_ADD_515_U161, new_P3_ADD_515_U162, new_P3_ADD_515_U163,
    new_P3_ADD_515_U164, new_P3_ADD_515_U165, new_P3_ADD_515_U166,
    new_P3_ADD_515_U167, new_P3_ADD_515_U168, new_P3_ADD_515_U169,
    new_P3_ADD_515_U170, new_P3_ADD_515_U171, new_P3_ADD_515_U172,
    new_P3_ADD_515_U173, new_P3_ADD_515_U174, new_P3_ADD_515_U175,
    new_P3_ADD_515_U176, new_P3_ADD_515_U177, new_P3_ADD_515_U178,
    new_P3_ADD_515_U179, new_P3_ADD_515_U180, new_P3_ADD_515_U181,
    new_P3_ADD_515_U182, new_P3_ADD_394_U4, new_P3_ADD_394_U5,
    new_P3_ADD_394_U6, new_P3_ADD_394_U7, new_P3_ADD_394_U8,
    new_P3_ADD_394_U9, new_P3_ADD_394_U10, new_P3_ADD_394_U11,
    new_P3_ADD_394_U12, new_P3_ADD_394_U13, new_P3_ADD_394_U14,
    new_P3_ADD_394_U15, new_P3_ADD_394_U16, new_P3_ADD_394_U17,
    new_P3_ADD_394_U18, new_P3_ADD_394_U19, new_P3_ADD_394_U20,
    new_P3_ADD_394_U21, new_P3_ADD_394_U22, new_P3_ADD_394_U23,
    new_P3_ADD_394_U24, new_P3_ADD_394_U25, new_P3_ADD_394_U26,
    new_P3_ADD_394_U27, new_P3_ADD_394_U28, new_P3_ADD_394_U29,
    new_P3_ADD_394_U30, new_P3_ADD_394_U31, new_P3_ADD_394_U32,
    new_P3_ADD_394_U33, new_P3_ADD_394_U34, new_P3_ADD_394_U35,
    new_P3_ADD_394_U36, new_P3_ADD_394_U37, new_P3_ADD_394_U38,
    new_P3_ADD_394_U39, new_P3_ADD_394_U40, new_P3_ADD_394_U41,
    new_P3_ADD_394_U42, new_P3_ADD_394_U43, new_P3_ADD_394_U44,
    new_P3_ADD_394_U45, new_P3_ADD_394_U46, new_P3_ADD_394_U47,
    new_P3_ADD_394_U48, new_P3_ADD_394_U49, new_P3_ADD_394_U50,
    new_P3_ADD_394_U51, new_P3_ADD_394_U52, new_P3_ADD_394_U53,
    new_P3_ADD_394_U54, new_P3_ADD_394_U55, new_P3_ADD_394_U56,
    new_P3_ADD_394_U57, new_P3_ADD_394_U58, new_P3_ADD_394_U59,
    new_P3_ADD_394_U60, new_P3_ADD_394_U61, new_P3_ADD_394_U62,
    new_P3_ADD_394_U63, new_P3_ADD_394_U64, new_P3_ADD_394_U65,
    new_P3_ADD_394_U66, new_P3_ADD_394_U67, new_P3_ADD_394_U68,
    new_P3_ADD_394_U69, new_P3_ADD_394_U70, new_P3_ADD_394_U71,
    new_P3_ADD_394_U72, new_P3_ADD_394_U73, new_P3_ADD_394_U74,
    new_P3_ADD_394_U75, new_P3_ADD_394_U76, new_P3_ADD_394_U77,
    new_P3_ADD_394_U78, new_P3_ADD_394_U79, new_P3_ADD_394_U80,
    new_P3_ADD_394_U81, new_P3_ADD_394_U82, new_P3_ADD_394_U83,
    new_P3_ADD_394_U84, new_P3_ADD_394_U85, new_P3_ADD_394_U86,
    new_P3_ADD_394_U87, new_P3_ADD_394_U88, new_P3_ADD_394_U89,
    new_P3_ADD_394_U90, new_P3_ADD_394_U91, new_P3_ADD_394_U92,
    new_P3_ADD_394_U93, new_P3_ADD_394_U94, new_P3_ADD_394_U95,
    new_P3_ADD_394_U96, new_P3_ADD_394_U97, new_P3_ADD_394_U98,
    new_P3_ADD_394_U99, new_P3_ADD_394_U100, new_P3_ADD_394_U101,
    new_P3_ADD_394_U102, new_P3_ADD_394_U103, new_P3_ADD_394_U104,
    new_P3_ADD_394_U105, new_P3_ADD_394_U106, new_P3_ADD_394_U107,
    new_P3_ADD_394_U108, new_P3_ADD_394_U109, new_P3_ADD_394_U110,
    new_P3_ADD_394_U111, new_P3_ADD_394_U112, new_P3_ADD_394_U113,
    new_P3_ADD_394_U114, new_P3_ADD_394_U115, new_P3_ADD_394_U116,
    new_P3_ADD_394_U117, new_P3_ADD_394_U118, new_P3_ADD_394_U119,
    new_P3_ADD_394_U120, new_P3_ADD_394_U121, new_P3_ADD_394_U122,
    new_P3_ADD_394_U123, new_P3_ADD_394_U124, new_P3_ADD_394_U125,
    new_P3_ADD_394_U126, new_P3_ADD_394_U127, new_P3_ADD_394_U128,
    new_P3_ADD_394_U129, new_P3_ADD_394_U130, new_P3_ADD_394_U131,
    new_P3_ADD_394_U132, new_P3_ADD_394_U133, new_P3_ADD_394_U134,
    new_P3_ADD_394_U135, new_P3_ADD_394_U136, new_P3_ADD_394_U137,
    new_P3_ADD_394_U138, new_P3_ADD_394_U139, new_P3_ADD_394_U140,
    new_P3_ADD_394_U141, new_P3_ADD_394_U142, new_P3_ADD_394_U143,
    new_P3_ADD_394_U144, new_P3_ADD_394_U145, new_P3_ADD_394_U146,
    new_P3_ADD_394_U147, new_P3_ADD_394_U148, new_P3_ADD_394_U149,
    new_P3_ADD_394_U150, new_P3_ADD_394_U151, new_P3_ADD_394_U152,
    new_P3_ADD_394_U153, new_P3_ADD_394_U154, new_P3_ADD_394_U155,
    new_P3_ADD_394_U156, new_P3_ADD_394_U157, new_P3_ADD_394_U158,
    new_P3_ADD_394_U159, new_P3_ADD_394_U160, new_P3_ADD_394_U161,
    new_P3_ADD_394_U162, new_P3_ADD_394_U163, new_P3_ADD_394_U164,
    new_P3_ADD_394_U165, new_P3_ADD_394_U166, new_P3_ADD_394_U167,
    new_P3_ADD_394_U168, new_P3_ADD_394_U169, new_P3_ADD_394_U170,
    new_P3_ADD_394_U171, new_P3_ADD_394_U172, new_P3_ADD_394_U173,
    new_P3_ADD_394_U174, new_P3_ADD_394_U175, new_P3_ADD_394_U176,
    new_P3_ADD_394_U177, new_P3_ADD_394_U178, new_P3_ADD_394_U179,
    new_P3_ADD_394_U180, new_P3_ADD_394_U181, new_P3_ADD_394_U182,
    new_P3_ADD_394_U183, new_P3_ADD_394_U184, new_P3_ADD_394_U185,
    new_P3_ADD_394_U186, new_P3_GTE_450_U6, new_P3_GTE_450_U7,
    new_P3_SUB_414_U6, new_P3_SUB_414_U7, new_P3_SUB_414_U8,
    new_P3_SUB_414_U9, new_P3_SUB_414_U10, new_P3_SUB_414_U11,
    new_P3_SUB_414_U12, new_P3_SUB_414_U13, new_P3_SUB_414_U14,
    new_P3_SUB_414_U15, new_P3_SUB_414_U16, new_P3_SUB_414_U17,
    new_P3_SUB_414_U18, new_P3_SUB_414_U19, new_P3_SUB_414_U20,
    new_P3_SUB_414_U21, new_P3_SUB_414_U22, new_P3_SUB_414_U23,
    new_P3_SUB_414_U24, new_P3_SUB_414_U25, new_P3_SUB_414_U26,
    new_P3_SUB_414_U27, new_P3_SUB_414_U28, new_P3_SUB_414_U29,
    new_P3_SUB_414_U30, new_P3_SUB_414_U31, new_P3_SUB_414_U32,
    new_P3_SUB_414_U33, new_P3_SUB_414_U34, new_P3_SUB_414_U35,
    new_P3_SUB_414_U36, new_P3_SUB_414_U37, new_P3_SUB_414_U38,
    new_P3_SUB_414_U39, new_P3_SUB_414_U40, new_P3_SUB_414_U41,
    new_P3_SUB_414_U42, new_P3_SUB_414_U43, new_P3_SUB_414_U44,
    new_P3_SUB_414_U45, new_P3_SUB_414_U46, new_P3_SUB_414_U47,
    new_P3_SUB_414_U48, new_P3_SUB_414_U49, new_P3_SUB_414_U50,
    new_P3_SUB_414_U51, new_P3_SUB_414_U52, new_P3_SUB_414_U53,
    new_P3_SUB_414_U54, new_P3_SUB_414_U55, new_P3_SUB_414_U56,
    new_P3_SUB_414_U57, new_P3_SUB_414_U58, new_P3_SUB_414_U59,
    new_P3_SUB_414_U60, new_P3_SUB_414_U61, new_P3_SUB_414_U62,
    new_P3_SUB_414_U63, new_P3_SUB_414_U64, new_P3_SUB_414_U65,
    new_P3_SUB_414_U66, new_P3_SUB_414_U67, new_P3_SUB_414_U68,
    new_P3_SUB_414_U69, new_P3_SUB_414_U70, new_P3_SUB_414_U71,
    new_P3_SUB_414_U72, new_P3_SUB_414_U73, new_P3_SUB_414_U74,
    new_P3_SUB_414_U75, new_P3_SUB_414_U76, new_P3_SUB_414_U77,
    new_P3_SUB_414_U78, new_P3_SUB_414_U79, new_P3_SUB_414_U80,
    new_P3_SUB_414_U81, new_P3_SUB_414_U82, new_P3_SUB_414_U83,
    new_P3_SUB_414_U84, new_P3_SUB_414_U85, new_P3_SUB_414_U86,
    new_P3_SUB_414_U87, new_P3_SUB_414_U88, new_P3_SUB_414_U89,
    new_P3_SUB_414_U90, new_P3_SUB_414_U91, new_P3_SUB_414_U92,
    new_P3_SUB_414_U93, new_P3_SUB_414_U94, new_P3_SUB_414_U95,
    new_P3_SUB_414_U96, new_P3_SUB_414_U97, new_P3_SUB_414_U98,
    new_P3_SUB_414_U99, new_P3_SUB_414_U100, new_P3_SUB_414_U101,
    new_P3_SUB_414_U102, new_P3_SUB_414_U103, new_P3_SUB_414_U104,
    new_P3_SUB_414_U105, new_P3_SUB_414_U106, new_P3_SUB_414_U107,
    new_P3_SUB_414_U108, new_P3_SUB_414_U109, new_P3_SUB_414_U110,
    new_P3_SUB_414_U111, new_P3_SUB_414_U112, new_P3_SUB_414_U113,
    new_P3_SUB_414_U114, new_P3_SUB_414_U115, new_P3_SUB_414_U116,
    new_P3_SUB_414_U117, new_P3_SUB_414_U118, new_P3_SUB_414_U119,
    new_P3_SUB_414_U120, new_P3_SUB_414_U121, new_P3_SUB_414_U122,
    new_P3_SUB_414_U123, new_P3_SUB_414_U124, new_P3_SUB_414_U125,
    new_P3_SUB_414_U126, new_P3_SUB_414_U127, new_P3_SUB_414_U128,
    new_P3_SUB_414_U129, new_P3_SUB_414_U130, new_P3_SUB_414_U131,
    new_P3_SUB_414_U132, new_P3_SUB_414_U133, new_P3_SUB_414_U134,
    new_P3_SUB_414_U135, new_P3_SUB_414_U136, new_P3_SUB_414_U137,
    new_P3_SUB_414_U138, new_P3_SUB_414_U139, new_P3_SUB_414_U140,
    new_P3_SUB_414_U141, new_P3_SUB_414_U142, new_P3_SUB_414_U143,
    new_P3_SUB_414_U144, new_P3_SUB_414_U145, new_P3_SUB_414_U146,
    new_P3_SUB_414_U147, new_P3_SUB_414_U148, new_P3_SUB_414_U149,
    new_P3_SUB_414_U150, new_P3_SUB_414_U151, new_P3_SUB_414_U152,
    new_P3_SUB_414_U153, new_P3_SUB_414_U154, new_P3_SUB_414_U155,
    new_P3_SUB_414_U156, new_P3_SUB_414_U157, new_P3_SUB_414_U158,
    new_P3_SUB_414_U159, new_P3_ADD_441_U4, new_P3_ADD_441_U5,
    new_P3_ADD_441_U6, new_P3_ADD_441_U7, new_P3_ADD_441_U8,
    new_P3_ADD_441_U9, new_P3_ADD_441_U10, new_P3_ADD_441_U11,
    new_P3_ADD_441_U12, new_P3_ADD_441_U13, new_P3_ADD_441_U14,
    new_P3_ADD_441_U15, new_P3_ADD_441_U16, new_P3_ADD_441_U17,
    new_P3_ADD_441_U18, new_P3_ADD_441_U19, new_P3_ADD_441_U20,
    new_P3_ADD_441_U21, new_P3_ADD_441_U22, new_P3_ADD_441_U23,
    new_P3_ADD_441_U24, new_P3_ADD_441_U25, new_P3_ADD_441_U26,
    new_P3_ADD_441_U27, new_P3_ADD_441_U28, new_P3_ADD_441_U29,
    new_P3_ADD_441_U30, new_P3_ADD_441_U31, new_P3_ADD_441_U32,
    new_P3_ADD_441_U33, new_P3_ADD_441_U34, new_P3_ADD_441_U35,
    new_P3_ADD_441_U36, new_P3_ADD_441_U37, new_P3_ADD_441_U38,
    new_P3_ADD_441_U39, new_P3_ADD_441_U40, new_P3_ADD_441_U41,
    new_P3_ADD_441_U42, new_P3_ADD_441_U43, new_P3_ADD_441_U44,
    new_P3_ADD_441_U45, new_P3_ADD_441_U46, new_P3_ADD_441_U47,
    new_P3_ADD_441_U48, new_P3_ADD_441_U49, new_P3_ADD_441_U50,
    new_P3_ADD_441_U51, new_P3_ADD_441_U52, new_P3_ADD_441_U53,
    new_P3_ADD_441_U54, new_P3_ADD_441_U55, new_P3_ADD_441_U56,
    new_P3_ADD_441_U57, new_P3_ADD_441_U58, new_P3_ADD_441_U59,
    new_P3_ADD_441_U60, new_P3_ADD_441_U61, new_P3_ADD_441_U62,
    new_P3_ADD_441_U63, new_P3_ADD_441_U64, new_P3_ADD_441_U65,
    new_P3_ADD_441_U66, new_P3_ADD_441_U67, new_P3_ADD_441_U68,
    new_P3_ADD_441_U69, new_P3_ADD_441_U70, new_P3_ADD_441_U71,
    new_P3_ADD_441_U72, new_P3_ADD_441_U73, new_P3_ADD_441_U74,
    new_P3_ADD_441_U75, new_P3_ADD_441_U76, new_P3_ADD_441_U77,
    new_P3_ADD_441_U78, new_P3_ADD_441_U79, new_P3_ADD_441_U80,
    new_P3_ADD_441_U81, new_P3_ADD_441_U82, new_P3_ADD_441_U83,
    new_P3_ADD_441_U84, new_P3_ADD_441_U85, new_P3_ADD_441_U86,
    new_P3_ADD_441_U87, new_P3_ADD_441_U88, new_P3_ADD_441_U89,
    new_P3_ADD_441_U90, new_P3_ADD_441_U91, new_P3_ADD_441_U92,
    new_P3_ADD_441_U93, new_P3_ADD_441_U94, new_P3_ADD_441_U95,
    new_P3_ADD_441_U96, new_P3_ADD_441_U97, new_P3_ADD_441_U98,
    new_P3_ADD_441_U99, new_P3_ADD_441_U100, new_P3_ADD_441_U101,
    new_P3_ADD_441_U102, new_P3_ADD_441_U103, new_P3_ADD_441_U104,
    new_P3_ADD_441_U105, new_P3_ADD_441_U106, new_P3_ADD_441_U107,
    new_P3_ADD_441_U108, new_P3_ADD_441_U109, new_P3_ADD_441_U110,
    new_P3_ADD_441_U111, new_P3_ADD_441_U112, new_P3_ADD_441_U113,
    new_P3_ADD_441_U114, new_P3_ADD_441_U115, new_P3_ADD_441_U116,
    new_P3_ADD_441_U117, new_P3_ADD_441_U118, new_P3_ADD_441_U119,
    new_P3_ADD_441_U120, new_P3_ADD_441_U121, new_P3_ADD_441_U122,
    new_P3_ADD_441_U123, new_P3_ADD_441_U124, new_P3_ADD_441_U125,
    new_P3_ADD_441_U126, new_P3_ADD_441_U127, new_P3_ADD_441_U128,
    new_P3_ADD_441_U129, new_P3_ADD_441_U130, new_P3_ADD_441_U131,
    new_P3_ADD_441_U132, new_P3_ADD_441_U133, new_P3_ADD_441_U134,
    new_P3_ADD_441_U135, new_P3_ADD_441_U136, new_P3_ADD_441_U137,
    new_P3_ADD_441_U138, new_P3_ADD_441_U139, new_P3_ADD_441_U140,
    new_P3_ADD_441_U141, new_P3_ADD_441_U142, new_P3_ADD_441_U143,
    new_P3_ADD_441_U144, new_P3_ADD_441_U145, new_P3_ADD_441_U146,
    new_P3_ADD_441_U147, new_P3_ADD_441_U148, new_P3_ADD_441_U149,
    new_P3_ADD_441_U150, new_P3_ADD_441_U151, new_P3_ADD_441_U152,
    new_P3_ADD_441_U153, new_P3_ADD_441_U154, new_P3_ADD_441_U155,
    new_P3_ADD_441_U156, new_P3_ADD_441_U157, new_P3_ADD_441_U158,
    new_P3_ADD_441_U159, new_P3_ADD_441_U160, new_P3_ADD_441_U161,
    new_P3_ADD_441_U162, new_P3_ADD_441_U163, new_P3_ADD_441_U164,
    new_P3_ADD_441_U165, new_P3_ADD_441_U166, new_P3_ADD_441_U167,
    new_P3_ADD_441_U168, new_P3_ADD_441_U169, new_P3_ADD_441_U170,
    new_P3_ADD_441_U171, new_P3_ADD_441_U172, new_P3_ADD_441_U173,
    new_P3_ADD_441_U174, new_P3_ADD_441_U175, new_P3_ADD_441_U176,
    new_P3_ADD_441_U177, new_P3_ADD_441_U178, new_P3_ADD_441_U179,
    new_P3_ADD_441_U180, new_P3_ADD_441_U181, new_P3_ADD_441_U182,
    new_P3_ADD_349_U5, new_P3_ADD_349_U6, new_P3_ADD_349_U7,
    new_P3_ADD_349_U8, new_P3_ADD_349_U9, new_P3_ADD_349_U10,
    new_P3_ADD_349_U11, new_P3_ADD_349_U12, new_P3_ADD_349_U13,
    new_P3_ADD_349_U14, new_P3_ADD_349_U15, new_P3_ADD_349_U16,
    new_P3_ADD_349_U17, new_P3_ADD_349_U18, new_P3_ADD_349_U19,
    new_P3_ADD_349_U20, new_P3_ADD_349_U21, new_P3_ADD_349_U22,
    new_P3_ADD_349_U23, new_P3_ADD_349_U24, new_P3_ADD_349_U25,
    new_P3_ADD_349_U26, new_P3_ADD_349_U27, new_P3_ADD_349_U28,
    new_P3_ADD_349_U29, new_P3_ADD_349_U30, new_P3_ADD_349_U31,
    new_P3_ADD_349_U32, new_P3_ADD_349_U33, new_P3_ADD_349_U34,
    new_P3_ADD_349_U35, new_P3_ADD_349_U36, new_P3_ADD_349_U37,
    new_P3_ADD_349_U38, new_P3_ADD_349_U39, new_P3_ADD_349_U40,
    new_P3_ADD_349_U41, new_P3_ADD_349_U42, new_P3_ADD_349_U43,
    new_P3_ADD_349_U44, new_P3_ADD_349_U45, new_P3_ADD_349_U46,
    new_P3_ADD_349_U47, new_P3_ADD_349_U48, new_P3_ADD_349_U49,
    new_P3_ADD_349_U50, new_P3_ADD_349_U51, new_P3_ADD_349_U52,
    new_P3_ADD_349_U53, new_P3_ADD_349_U54, new_P3_ADD_349_U55,
    new_P3_ADD_349_U56, new_P3_ADD_349_U57, new_P3_ADD_349_U58,
    new_P3_ADD_349_U59, new_P3_ADD_349_U60, new_P3_ADD_349_U61,
    new_P3_ADD_349_U62, new_P3_ADD_349_U63, new_P3_ADD_349_U64,
    new_P3_ADD_349_U65, new_P3_ADD_349_U66, new_P3_ADD_349_U67,
    new_P3_ADD_349_U68, new_P3_ADD_349_U69, new_P3_ADD_349_U70,
    new_P3_ADD_349_U71, new_P3_ADD_349_U72, new_P3_ADD_349_U73,
    new_P3_ADD_349_U74, new_P3_ADD_349_U75, new_P3_ADD_349_U76,
    new_P3_ADD_349_U77, new_P3_ADD_349_U78, new_P3_ADD_349_U79,
    new_P3_ADD_349_U80, new_P3_ADD_349_U81, new_P3_ADD_349_U82,
    new_P3_ADD_349_U83, new_P3_ADD_349_U84, new_P3_ADD_349_U85,
    new_P3_ADD_349_U86, new_P3_ADD_349_U87, new_P3_ADD_349_U88,
    new_P3_ADD_349_U89, new_P3_ADD_349_U90, new_P3_ADD_349_U91,
    new_P3_ADD_349_U92, new_P3_ADD_349_U93, new_P3_ADD_349_U94,
    new_P3_ADD_349_U95, new_P3_ADD_349_U96, new_P3_ADD_349_U97,
    new_P3_ADD_349_U98, new_P3_ADD_349_U99, new_P3_ADD_349_U100,
    new_P3_ADD_349_U101, new_P3_ADD_349_U102, new_P3_ADD_349_U103,
    new_P3_ADD_349_U104, new_P3_ADD_349_U105, new_P3_ADD_349_U106,
    new_P3_ADD_349_U107, new_P3_ADD_349_U108, new_P3_ADD_349_U109,
    new_P3_ADD_349_U110, new_P3_ADD_349_U111, new_P3_ADD_349_U112,
    new_P3_ADD_349_U113, new_P3_ADD_349_U114, new_P3_ADD_349_U115,
    new_P3_ADD_349_U116, new_P3_ADD_349_U117, new_P3_ADD_349_U118,
    new_P3_ADD_349_U119, new_P3_ADD_349_U120, new_P3_ADD_349_U121,
    new_P3_ADD_349_U122, new_P3_ADD_349_U123, new_P3_ADD_349_U124,
    new_P3_ADD_349_U125, new_P3_ADD_349_U126, new_P3_ADD_349_U127,
    new_P3_ADD_349_U128, new_P3_ADD_349_U129, new_P3_ADD_349_U130,
    new_P3_ADD_349_U131, new_P3_ADD_349_U132, new_P3_ADD_349_U133,
    new_P3_ADD_349_U134, new_P3_ADD_349_U135, new_P3_ADD_349_U136,
    new_P3_ADD_349_U137, new_P3_ADD_349_U138, new_P3_ADD_349_U139,
    new_P3_ADD_349_U140, new_P3_ADD_349_U141, new_P3_ADD_349_U142,
    new_P3_ADD_349_U143, new_P3_ADD_349_U144, new_P3_ADD_349_U145,
    new_P3_ADD_349_U146, new_P3_ADD_349_U147, new_P3_ADD_349_U148,
    new_P3_ADD_349_U149, new_P3_ADD_349_U150, new_P3_ADD_349_U151,
    new_P3_ADD_349_U152, new_P3_ADD_349_U153, new_P3_ADD_349_U154,
    new_P3_ADD_349_U155, new_P3_ADD_349_U156, new_P3_ADD_349_U157,
    new_P3_ADD_349_U158, new_P3_ADD_349_U159, new_P3_ADD_349_U160,
    new_P3_ADD_349_U161, new_P3_ADD_349_U162, new_P3_ADD_349_U163,
    new_P3_ADD_349_U164, new_P3_ADD_349_U165, new_P3_ADD_349_U166,
    new_P3_ADD_349_U167, new_P3_ADD_349_U168, new_P3_ADD_349_U169,
    new_P3_ADD_349_U170, new_P3_ADD_349_U171, new_P3_ADD_349_U172,
    new_P3_ADD_349_U173, new_P3_ADD_349_U174, new_P3_ADD_349_U175,
    new_P3_ADD_349_U176, new_P3_ADD_349_U177, new_P3_ADD_349_U178,
    new_P3_ADD_349_U179, new_P3_ADD_349_U180, new_P3_ADD_349_U181,
    new_P3_ADD_349_U182, new_P3_ADD_349_U183, new_P3_ADD_349_U184,
    new_P3_ADD_349_U185, new_P3_ADD_349_U186, new_P3_ADD_349_U187,
    new_P3_ADD_349_U188, new_P3_ADD_349_U189, new_P3_ADD_405_U4,
    new_P3_ADD_405_U5, new_P3_ADD_405_U6, new_P3_ADD_405_U7,
    new_P3_ADD_405_U8, new_P3_ADD_405_U9, new_P3_ADD_405_U10,
    new_P3_ADD_405_U11, new_P3_ADD_405_U12, new_P3_ADD_405_U13,
    new_P3_ADD_405_U14, new_P3_ADD_405_U15, new_P3_ADD_405_U16,
    new_P3_ADD_405_U17, new_P3_ADD_405_U18, new_P3_ADD_405_U19,
    new_P3_ADD_405_U20, new_P3_ADD_405_U21, new_P3_ADD_405_U22,
    new_P3_ADD_405_U23, new_P3_ADD_405_U24, new_P3_ADD_405_U25,
    new_P3_ADD_405_U26, new_P3_ADD_405_U27, new_P3_ADD_405_U28,
    new_P3_ADD_405_U29, new_P3_ADD_405_U30, new_P3_ADD_405_U31,
    new_P3_ADD_405_U32, new_P3_ADD_405_U33, new_P3_ADD_405_U34,
    new_P3_ADD_405_U35, new_P3_ADD_405_U36, new_P3_ADD_405_U37,
    new_P3_ADD_405_U38, new_P3_ADD_405_U39, new_P3_ADD_405_U40,
    new_P3_ADD_405_U41, new_P3_ADD_405_U42, new_P3_ADD_405_U43,
    new_P3_ADD_405_U44, new_P3_ADD_405_U45, new_P3_ADD_405_U46,
    new_P3_ADD_405_U47, new_P3_ADD_405_U48, new_P3_ADD_405_U49,
    new_P3_ADD_405_U50, new_P3_ADD_405_U51, new_P3_ADD_405_U52,
    new_P3_ADD_405_U53, new_P3_ADD_405_U54, new_P3_ADD_405_U55,
    new_P3_ADD_405_U56, new_P3_ADD_405_U57, new_P3_ADD_405_U58,
    new_P3_ADD_405_U59, new_P3_ADD_405_U60, new_P3_ADD_405_U61,
    new_P3_ADD_405_U62, new_P3_ADD_405_U63, new_P3_ADD_405_U64,
    new_P3_ADD_405_U65, new_P3_ADD_405_U66, new_P3_ADD_405_U67,
    new_P3_ADD_405_U68, new_P3_ADD_405_U69, new_P3_ADD_405_U70,
    new_P3_ADD_405_U71, new_P3_ADD_405_U72, new_P3_ADD_405_U73,
    new_P3_ADD_405_U74, new_P3_ADD_405_U75, new_P3_ADD_405_U76,
    new_P3_ADD_405_U77, new_P3_ADD_405_U78, new_P3_ADD_405_U79,
    new_P3_ADD_405_U80, new_P3_ADD_405_U81, new_P3_ADD_405_U82,
    new_P3_ADD_405_U83, new_P3_ADD_405_U84, new_P3_ADD_405_U85,
    new_P3_ADD_405_U86, new_P3_ADD_405_U87, new_P3_ADD_405_U88,
    new_P3_ADD_405_U89, new_P3_ADD_405_U90, new_P3_ADD_405_U91,
    new_P3_ADD_405_U92, new_P3_ADD_405_U93, new_P3_ADD_405_U94,
    new_P3_ADD_405_U95, new_P3_ADD_405_U96, new_P3_ADD_405_U97,
    new_P3_ADD_405_U98, new_P3_ADD_405_U99, new_P3_ADD_405_U100,
    new_P3_ADD_405_U101, new_P3_ADD_405_U102, new_P3_ADD_405_U103,
    new_P3_ADD_405_U104, new_P3_ADD_405_U105, new_P3_ADD_405_U106,
    new_P3_ADD_405_U107, new_P3_ADD_405_U108, new_P3_ADD_405_U109,
    new_P3_ADD_405_U110, new_P3_ADD_405_U111, new_P3_ADD_405_U112,
    new_P3_ADD_405_U113, new_P3_ADD_405_U114, new_P3_ADD_405_U115,
    new_P3_ADD_405_U116, new_P3_ADD_405_U117, new_P3_ADD_405_U118,
    new_P3_ADD_405_U119, new_P3_ADD_405_U120, new_P3_ADD_405_U121,
    new_P3_ADD_405_U122, new_P3_ADD_405_U123, new_P3_ADD_405_U124,
    new_P3_ADD_405_U125, new_P3_ADD_405_U126, new_P3_ADD_405_U127,
    new_P3_ADD_405_U128, new_P3_ADD_405_U129, new_P3_ADD_405_U130,
    new_P3_ADD_405_U131, new_P3_ADD_405_U132, new_P3_ADD_405_U133,
    new_P3_ADD_405_U134, new_P3_ADD_405_U135, new_P3_ADD_405_U136,
    new_P3_ADD_405_U137, new_P3_ADD_405_U138, new_P3_ADD_405_U139,
    new_P3_ADD_405_U140, new_P3_ADD_405_U141, new_P3_ADD_405_U142,
    new_P3_ADD_405_U143, new_P3_ADD_405_U144, new_P3_ADD_405_U145,
    new_P3_ADD_405_U146, new_P3_ADD_405_U147, new_P3_ADD_405_U148,
    new_P3_ADD_405_U149, new_P3_ADD_405_U150, new_P3_ADD_405_U151,
    new_P3_ADD_405_U152, new_P3_ADD_405_U153, new_P3_ADD_405_U154,
    new_P3_ADD_405_U155, new_P3_ADD_405_U156, new_P3_ADD_405_U157,
    new_P3_ADD_405_U158, new_P3_ADD_405_U159, new_P3_ADD_405_U160,
    new_P3_ADD_405_U161, new_P3_ADD_405_U162, new_P3_ADD_405_U163,
    new_P3_ADD_405_U164, new_P3_ADD_405_U165, new_P3_ADD_405_U166,
    new_P3_ADD_405_U167, new_P3_ADD_405_U168, new_P3_ADD_405_U169,
    new_P3_ADD_405_U170, new_P3_ADD_405_U171, new_P3_ADD_405_U172,
    new_P3_ADD_405_U173, new_P3_ADD_405_U174, new_P3_ADD_405_U175,
    new_P3_ADD_405_U176, new_P3_ADD_405_U177, new_P3_ADD_405_U178,
    new_P3_ADD_405_U179, new_P3_ADD_405_U180, new_P3_ADD_405_U181,
    new_P3_ADD_405_U182, new_P3_ADD_405_U183, new_P3_ADD_405_U184,
    new_P3_ADD_405_U185, new_P3_ADD_405_U186, new_P3_ADD_553_U5,
    new_P3_ADD_553_U6, new_P3_ADD_553_U7, new_P3_ADD_553_U8,
    new_P3_ADD_553_U9, new_P3_ADD_553_U10, new_P3_ADD_553_U11,
    new_P3_ADD_553_U12, new_P3_ADD_553_U13, new_P3_ADD_553_U14,
    new_P3_ADD_553_U15, new_P3_ADD_553_U16, new_P3_ADD_553_U17,
    new_P3_ADD_553_U18, new_P3_ADD_553_U19, new_P3_ADD_553_U20,
    new_P3_ADD_553_U21, new_P3_ADD_553_U22, new_P3_ADD_553_U23,
    new_P3_ADD_553_U24, new_P3_ADD_553_U25, new_P3_ADD_553_U26,
    new_P3_ADD_553_U27, new_P3_ADD_553_U28, new_P3_ADD_553_U29,
    new_P3_ADD_553_U30, new_P3_ADD_553_U31, new_P3_ADD_553_U32,
    new_P3_ADD_553_U33, new_P3_ADD_553_U34, new_P3_ADD_553_U35,
    new_P3_ADD_553_U36, new_P3_ADD_553_U37, new_P3_ADD_553_U38,
    new_P3_ADD_553_U39, new_P3_ADD_553_U40, new_P3_ADD_553_U41,
    new_P3_ADD_553_U42, new_P3_ADD_553_U43, new_P3_ADD_553_U44,
    new_P3_ADD_553_U45, new_P3_ADD_553_U46, new_P3_ADD_553_U47,
    new_P3_ADD_553_U48, new_P3_ADD_553_U49, new_P3_ADD_553_U50,
    new_P3_ADD_553_U51, new_P3_ADD_553_U52, new_P3_ADD_553_U53,
    new_P3_ADD_553_U54, new_P3_ADD_553_U55, new_P3_ADD_553_U56,
    new_P3_ADD_553_U57, new_P3_ADD_553_U58, new_P3_ADD_553_U59,
    new_P3_ADD_553_U60, new_P3_ADD_553_U61, new_P3_ADD_553_U62,
    new_P3_ADD_553_U63, new_P3_ADD_553_U64, new_P3_ADD_553_U65,
    new_P3_ADD_553_U66, new_P3_ADD_553_U67, new_P3_ADD_553_U68,
    new_P3_ADD_553_U69, new_P3_ADD_553_U70, new_P3_ADD_553_U71,
    new_P3_ADD_553_U72, new_P3_ADD_553_U73, new_P3_ADD_553_U74,
    new_P3_ADD_553_U75, new_P3_ADD_553_U76, new_P3_ADD_553_U77,
    new_P3_ADD_553_U78, new_P3_ADD_553_U79, new_P3_ADD_553_U80,
    new_P3_ADD_553_U81, new_P3_ADD_553_U82, new_P3_ADD_553_U83,
    new_P3_ADD_553_U84, new_P3_ADD_553_U85, new_P3_ADD_553_U86,
    new_P3_ADD_553_U87, new_P3_ADD_553_U88, new_P3_ADD_553_U89,
    new_P3_ADD_553_U90, new_P3_ADD_553_U91, new_P3_ADD_553_U92,
    new_P3_ADD_553_U93, new_P3_ADD_553_U94, new_P3_ADD_553_U95,
    new_P3_ADD_553_U96, new_P3_ADD_553_U97, new_P3_ADD_553_U98,
    new_P3_ADD_553_U99, new_P3_ADD_553_U100, new_P3_ADD_553_U101,
    new_P3_ADD_553_U102, new_P3_ADD_553_U103, new_P3_ADD_553_U104,
    new_P3_ADD_553_U105, new_P3_ADD_553_U106, new_P3_ADD_553_U107,
    new_P3_ADD_553_U108, new_P3_ADD_553_U109, new_P3_ADD_553_U110,
    new_P3_ADD_553_U111, new_P3_ADD_553_U112, new_P3_ADD_553_U113,
    new_P3_ADD_553_U114, new_P3_ADD_553_U115, new_P3_ADD_553_U116,
    new_P3_ADD_553_U117, new_P3_ADD_553_U118, new_P3_ADD_553_U119,
    new_P3_ADD_553_U120, new_P3_ADD_553_U121, new_P3_ADD_553_U122,
    new_P3_ADD_553_U123, new_P3_ADD_553_U124, new_P3_ADD_553_U125,
    new_P3_ADD_553_U126, new_P3_ADD_553_U127, new_P3_ADD_553_U128,
    new_P3_ADD_553_U129, new_P3_ADD_553_U130, new_P3_ADD_553_U131,
    new_P3_ADD_553_U132, new_P3_ADD_553_U133, new_P3_ADD_553_U134,
    new_P3_ADD_553_U135, new_P3_ADD_553_U136, new_P3_ADD_553_U137,
    new_P3_ADD_553_U138, new_P3_ADD_553_U139, new_P3_ADD_553_U140,
    new_P3_ADD_553_U141, new_P3_ADD_553_U142, new_P3_ADD_553_U143,
    new_P3_ADD_553_U144, new_P3_ADD_553_U145, new_P3_ADD_553_U146,
    new_P3_ADD_553_U147, new_P3_ADD_553_U148, new_P3_ADD_553_U149,
    new_P3_ADD_553_U150, new_P3_ADD_553_U151, new_P3_ADD_553_U152,
    new_P3_ADD_553_U153, new_P3_ADD_553_U154, new_P3_ADD_553_U155,
    new_P3_ADD_553_U156, new_P3_ADD_553_U157, new_P3_ADD_553_U158,
    new_P3_ADD_553_U159, new_P3_ADD_553_U160, new_P3_ADD_553_U161,
    new_P3_ADD_553_U162, new_P3_ADD_553_U163, new_P3_ADD_553_U164,
    new_P3_ADD_553_U165, new_P3_ADD_553_U166, new_P3_ADD_553_U167,
    new_P3_ADD_553_U168, new_P3_ADD_553_U169, new_P3_ADD_553_U170,
    new_P3_ADD_553_U171, new_P3_ADD_553_U172, new_P3_ADD_553_U173,
    new_P3_ADD_553_U174, new_P3_ADD_553_U175, new_P3_ADD_553_U176,
    new_P3_ADD_553_U177, new_P3_ADD_553_U178, new_P3_ADD_553_U179,
    new_P3_ADD_553_U180, new_P3_ADD_553_U181, new_P3_ADD_553_U182,
    new_P3_ADD_553_U183, new_P3_ADD_553_U184, new_P3_ADD_553_U185,
    new_P3_ADD_553_U186, new_P3_ADD_553_U187, new_P3_ADD_553_U188,
    new_P3_ADD_553_U189, new_P3_ADD_558_U5, new_P3_ADD_558_U6,
    new_P3_ADD_558_U7, new_P3_ADD_558_U8, new_P3_ADD_558_U9,
    new_P3_ADD_558_U10, new_P3_ADD_558_U11, new_P3_ADD_558_U12,
    new_P3_ADD_558_U13, new_P3_ADD_558_U14, new_P3_ADD_558_U15,
    new_P3_ADD_558_U16, new_P3_ADD_558_U17, new_P3_ADD_558_U18,
    new_P3_ADD_558_U19, new_P3_ADD_558_U20, new_P3_ADD_558_U21,
    new_P3_ADD_558_U22, new_P3_ADD_558_U23, new_P3_ADD_558_U24,
    new_P3_ADD_558_U25, new_P3_ADD_558_U26, new_P3_ADD_558_U27,
    new_P3_ADD_558_U28, new_P3_ADD_558_U29, new_P3_ADD_558_U30,
    new_P3_ADD_558_U31, new_P3_ADD_558_U32, new_P3_ADD_558_U33,
    new_P3_ADD_558_U34, new_P3_ADD_558_U35, new_P3_ADD_558_U36,
    new_P3_ADD_558_U37, new_P3_ADD_558_U38, new_P3_ADD_558_U39,
    new_P3_ADD_558_U40, new_P3_ADD_558_U41, new_P3_ADD_558_U42,
    new_P3_ADD_558_U43, new_P3_ADD_558_U44, new_P3_ADD_558_U45,
    new_P3_ADD_558_U46, new_P3_ADD_558_U47, new_P3_ADD_558_U48,
    new_P3_ADD_558_U49, new_P3_ADD_558_U50, new_P3_ADD_558_U51,
    new_P3_ADD_558_U52, new_P3_ADD_558_U53, new_P3_ADD_558_U54,
    new_P3_ADD_558_U55, new_P3_ADD_558_U56, new_P3_ADD_558_U57,
    new_P3_ADD_558_U58, new_P3_ADD_558_U59, new_P3_ADD_558_U60,
    new_P3_ADD_558_U61, new_P3_ADD_558_U62, new_P3_ADD_558_U63,
    new_P3_ADD_558_U64, new_P3_ADD_558_U65, new_P3_ADD_558_U66,
    new_P3_ADD_558_U67, new_P3_ADD_558_U68, new_P3_ADD_558_U69,
    new_P3_ADD_558_U70, new_P3_ADD_558_U71, new_P3_ADD_558_U72,
    new_P3_ADD_558_U73, new_P3_ADD_558_U74, new_P3_ADD_558_U75,
    new_P3_ADD_558_U76, new_P3_ADD_558_U77, new_P3_ADD_558_U78,
    new_P3_ADD_558_U79, new_P3_ADD_558_U80, new_P3_ADD_558_U81,
    new_P3_ADD_558_U82, new_P3_ADD_558_U83, new_P3_ADD_558_U84,
    new_P3_ADD_558_U85, new_P3_ADD_558_U86, new_P3_ADD_558_U87,
    new_P3_ADD_558_U88, new_P3_ADD_558_U89, new_P3_ADD_558_U90,
    new_P3_ADD_558_U91, new_P3_ADD_558_U92, new_P3_ADD_558_U93,
    new_P3_ADD_558_U94, new_P3_ADD_558_U95, new_P3_ADD_558_U96,
    new_P3_ADD_558_U97, new_P3_ADD_558_U98, new_P3_ADD_558_U99,
    new_P3_ADD_558_U100, new_P3_ADD_558_U101, new_P3_ADD_558_U102,
    new_P3_ADD_558_U103, new_P3_ADD_558_U104, new_P3_ADD_558_U105,
    new_P3_ADD_558_U106, new_P3_ADD_558_U107, new_P3_ADD_558_U108,
    new_P3_ADD_558_U109, new_P3_ADD_558_U110, new_P3_ADD_558_U111,
    new_P3_ADD_558_U112, new_P3_ADD_558_U113, new_P3_ADD_558_U114,
    new_P3_ADD_558_U115, new_P3_ADD_558_U116, new_P3_ADD_558_U117,
    new_P3_ADD_558_U118, new_P3_ADD_558_U119, new_P3_ADD_558_U120,
    new_P3_ADD_558_U121, new_P3_ADD_558_U122, new_P3_ADD_558_U123,
    new_P3_ADD_558_U124, new_P3_ADD_558_U125, new_P3_ADD_558_U126,
    new_P3_ADD_558_U127, new_P3_ADD_558_U128, new_P3_ADD_558_U129,
    new_P3_ADD_558_U130, new_P3_ADD_558_U131, new_P3_ADD_558_U132,
    new_P3_ADD_558_U133, new_P3_ADD_558_U134, new_P3_ADD_558_U135,
    new_P3_ADD_558_U136, new_P3_ADD_558_U137, new_P3_ADD_558_U138,
    new_P3_ADD_558_U139, new_P3_ADD_558_U140, new_P3_ADD_558_U141,
    new_P3_ADD_558_U142, new_P3_ADD_558_U143, new_P3_ADD_558_U144,
    new_P3_ADD_558_U145, new_P3_ADD_558_U146, new_P3_ADD_558_U147,
    new_P3_ADD_558_U148, new_P3_ADD_558_U149, new_P3_ADD_558_U150,
    new_P3_ADD_558_U151, new_P3_ADD_558_U152, new_P3_ADD_558_U153,
    new_P3_ADD_558_U154, new_P3_ADD_558_U155, new_P3_ADD_558_U156,
    new_P3_ADD_558_U157, new_P3_ADD_558_U158, new_P3_ADD_558_U159,
    new_P3_ADD_558_U160, new_P3_ADD_558_U161, new_P3_ADD_558_U162,
    new_P3_ADD_558_U163, new_P3_ADD_558_U164, new_P3_ADD_558_U165,
    new_P3_ADD_558_U166, new_P3_ADD_558_U167, new_P3_ADD_558_U168,
    new_P3_ADD_558_U169, new_P3_ADD_558_U170, new_P3_ADD_558_U171,
    new_P3_ADD_558_U172, new_P3_ADD_558_U173, new_P3_ADD_558_U174,
    new_P3_ADD_558_U175, new_P3_ADD_558_U176, new_P3_ADD_558_U177,
    new_P3_ADD_558_U178, new_P3_ADD_558_U179, new_P3_ADD_558_U180,
    new_P3_ADD_558_U181, new_P3_ADD_558_U182, new_P3_ADD_558_U183,
    new_P3_ADD_558_U184, new_P3_ADD_558_U185, new_P3_ADD_558_U186,
    new_P3_ADD_558_U187, new_P3_ADD_558_U188, new_P3_ADD_558_U189,
    new_P3_ADD_385_U5, new_P3_ADD_385_U6, new_P3_ADD_385_U7,
    new_P3_ADD_385_U8, new_P3_ADD_385_U9, new_P3_ADD_385_U10,
    new_P3_ADD_385_U11, new_P3_ADD_385_U12, new_P3_ADD_385_U13,
    new_P3_ADD_385_U14, new_P3_ADD_385_U15, new_P3_ADD_385_U16,
    new_P3_ADD_385_U17, new_P3_ADD_385_U18, new_P3_ADD_385_U19,
    new_P3_ADD_385_U20, new_P3_ADD_385_U21, new_P3_ADD_385_U22,
    new_P3_ADD_385_U23, new_P3_ADD_385_U24, new_P3_ADD_385_U25,
    new_P3_ADD_385_U26, new_P3_ADD_385_U27, new_P3_ADD_385_U28,
    new_P3_ADD_385_U29, new_P3_ADD_385_U30, new_P3_ADD_385_U31,
    new_P3_ADD_385_U32, new_P3_ADD_385_U33, new_P3_ADD_385_U34,
    new_P3_ADD_385_U35, new_P3_ADD_385_U36, new_P3_ADD_385_U37,
    new_P3_ADD_385_U38, new_P3_ADD_385_U39, new_P3_ADD_385_U40,
    new_P3_ADD_385_U41, new_P3_ADD_385_U42, new_P3_ADD_385_U43,
    new_P3_ADD_385_U44, new_P3_ADD_385_U45, new_P3_ADD_385_U46,
    new_P3_ADD_385_U47, new_P3_ADD_385_U48, new_P3_ADD_385_U49,
    new_P3_ADD_385_U50, new_P3_ADD_385_U51, new_P3_ADD_385_U52,
    new_P3_ADD_385_U53, new_P3_ADD_385_U54, new_P3_ADD_385_U55,
    new_P3_ADD_385_U56, new_P3_ADD_385_U57, new_P3_ADD_385_U58,
    new_P3_ADD_385_U59, new_P3_ADD_385_U60, new_P3_ADD_385_U61,
    new_P3_ADD_385_U62, new_P3_ADD_385_U63, new_P3_ADD_385_U64,
    new_P3_ADD_385_U65, new_P3_ADD_385_U66, new_P3_ADD_385_U67,
    new_P3_ADD_385_U68, new_P3_ADD_385_U69, new_P3_ADD_385_U70,
    new_P3_ADD_385_U71, new_P3_ADD_385_U72, new_P3_ADD_385_U73,
    new_P3_ADD_385_U74, new_P3_ADD_385_U75, new_P3_ADD_385_U76,
    new_P3_ADD_385_U77, new_P3_ADD_385_U78, new_P3_ADD_385_U79,
    new_P3_ADD_385_U80, new_P3_ADD_385_U81, new_P3_ADD_385_U82,
    new_P3_ADD_385_U83, new_P3_ADD_385_U84, new_P3_ADD_385_U85,
    new_P3_ADD_385_U86, new_P3_ADD_385_U87, new_P3_ADD_385_U88,
    new_P3_ADD_385_U89, new_P3_ADD_385_U90, new_P3_ADD_385_U91,
    new_P3_ADD_385_U92, new_P3_ADD_385_U93, new_P3_ADD_385_U94,
    new_P3_ADD_385_U95, new_P3_ADD_385_U96, new_P3_ADD_385_U97,
    new_P3_ADD_385_U98, new_P3_ADD_385_U99, new_P3_ADD_385_U100,
    new_P3_ADD_385_U101, new_P3_ADD_385_U102, new_P3_ADD_385_U103,
    new_P3_ADD_385_U104, new_P3_ADD_385_U105, new_P3_ADD_385_U106,
    new_P3_ADD_385_U107, new_P3_ADD_385_U108, new_P3_ADD_385_U109,
    new_P3_ADD_385_U110, new_P3_ADD_385_U111, new_P3_ADD_385_U112,
    new_P3_ADD_385_U113, new_P3_ADD_385_U114, new_P3_ADD_385_U115,
    new_P3_ADD_385_U116, new_P3_ADD_385_U117, new_P3_ADD_385_U118,
    new_P3_ADD_385_U119, new_P3_ADD_385_U120, new_P3_ADD_385_U121,
    new_P3_ADD_385_U122, new_P3_ADD_385_U123, new_P3_ADD_385_U124,
    new_P3_ADD_385_U125, new_P3_ADD_385_U126, new_P3_ADD_385_U127,
    new_P3_ADD_385_U128, new_P3_ADD_385_U129, new_P3_ADD_385_U130,
    new_P3_ADD_385_U131, new_P3_ADD_385_U132, new_P3_ADD_385_U133,
    new_P3_ADD_385_U134, new_P3_ADD_385_U135, new_P3_ADD_385_U136,
    new_P3_ADD_385_U137, new_P3_ADD_385_U138, new_P3_ADD_385_U139,
    new_P3_ADD_385_U140, new_P3_ADD_385_U141, new_P3_ADD_385_U142,
    new_P3_ADD_385_U143, new_P3_ADD_385_U144, new_P3_ADD_385_U145,
    new_P3_ADD_385_U146, new_P3_ADD_385_U147, new_P3_ADD_385_U148,
    new_P3_ADD_385_U149, new_P3_ADD_385_U150, new_P3_ADD_385_U151,
    new_P3_ADD_385_U152, new_P3_ADD_385_U153, new_P3_ADD_385_U154,
    new_P3_ADD_385_U155, new_P3_ADD_385_U156, new_P3_ADD_385_U157,
    new_P3_ADD_385_U158, new_P3_ADD_385_U159, new_P3_ADD_385_U160,
    new_P3_ADD_385_U161, new_P3_ADD_385_U162, new_P3_ADD_385_U163,
    new_P3_ADD_385_U164, new_P3_ADD_385_U165, new_P3_ADD_385_U166,
    new_P3_ADD_385_U167, new_P3_ADD_385_U168, new_P3_ADD_385_U169,
    new_P3_ADD_385_U170, new_P3_ADD_385_U171, new_P3_ADD_385_U172,
    new_P3_ADD_385_U173, new_P3_ADD_385_U174, new_P3_ADD_385_U175,
    new_P3_ADD_385_U176, new_P3_ADD_385_U177, new_P3_ADD_385_U178,
    new_P3_ADD_385_U179, new_P3_ADD_385_U180, new_P3_ADD_385_U181,
    new_P3_ADD_385_U182, new_P3_ADD_385_U183, new_P3_ADD_385_U184,
    new_P3_ADD_385_U185, new_P3_ADD_385_U186, new_P3_ADD_385_U187,
    new_P3_ADD_385_U188, new_P3_ADD_385_U189, new_P3_ADD_357_U6,
    new_P3_ADD_357_U7, new_P3_ADD_357_U8, new_P3_ADD_357_U9,
    new_P3_ADD_357_U10, new_P3_ADD_357_U11, new_P3_ADD_357_U12,
    new_P3_ADD_357_U13, new_P3_ADD_357_U14, new_P3_ADD_357_U15,
    new_P3_ADD_357_U16, new_P3_ADD_357_U17, new_P3_ADD_357_U18,
    new_P3_ADD_357_U19, new_P3_ADD_357_U20, new_P3_ADD_357_U21,
    new_P3_ADD_357_U22, new_P3_ADD_357_U23, new_P3_ADD_357_U24,
    new_P3_ADD_357_U25, new_P3_ADD_357_U26, new_P3_ADD_357_U27,
    new_P3_ADD_357_U28, new_P3_ADD_357_U29, new_P3_ADD_357_U30,
    new_P3_ADD_357_U31, new_P3_ADD_357_U32, new_P3_ADD_357_U33,
    new_P3_ADD_357_U34, new_P3_ADD_357_U35, new_P3_ADD_547_U5,
    new_P3_ADD_547_U6, new_P3_ADD_547_U7, new_P3_ADD_547_U8,
    new_P3_ADD_547_U9, new_P3_ADD_547_U10, new_P3_ADD_547_U11,
    new_P3_ADD_547_U12, new_P3_ADD_547_U13, new_P3_ADD_547_U14,
    new_P3_ADD_547_U15, new_P3_ADD_547_U16, new_P3_ADD_547_U17,
    new_P3_ADD_547_U18, new_P3_ADD_547_U19, new_P3_ADD_547_U20,
    new_P3_ADD_547_U21, new_P3_ADD_547_U22, new_P3_ADD_547_U23,
    new_P3_ADD_547_U24, new_P3_ADD_547_U25, new_P3_ADD_547_U26,
    new_P3_ADD_547_U27, new_P3_ADD_547_U28, new_P3_ADD_547_U29,
    new_P3_ADD_547_U30, new_P3_ADD_547_U31, new_P3_ADD_547_U32,
    new_P3_ADD_547_U33, new_P3_ADD_547_U34, new_P3_ADD_547_U35,
    new_P3_ADD_547_U36, new_P3_ADD_547_U37, new_P3_ADD_547_U38,
    new_P3_ADD_547_U39, new_P3_ADD_547_U40, new_P3_ADD_547_U41,
    new_P3_ADD_547_U42, new_P3_ADD_547_U43, new_P3_ADD_547_U44,
    new_P3_ADD_547_U45, new_P3_ADD_547_U46, new_P3_ADD_547_U47,
    new_P3_ADD_547_U48, new_P3_ADD_547_U49, new_P3_ADD_547_U50,
    new_P3_ADD_547_U51, new_P3_ADD_547_U52, new_P3_ADD_547_U53,
    new_P3_ADD_547_U54, new_P3_ADD_547_U55, new_P3_ADD_547_U56,
    new_P3_ADD_547_U57, new_P3_ADD_547_U58, new_P3_ADD_547_U59,
    new_P3_ADD_547_U60, new_P3_ADD_547_U61, new_P3_ADD_547_U62,
    new_P3_ADD_547_U63, new_P3_ADD_547_U64, new_P3_ADD_547_U65,
    new_P3_ADD_547_U66, new_P3_ADD_547_U67, new_P3_ADD_547_U68,
    new_P3_ADD_547_U69, new_P3_ADD_547_U70, new_P3_ADD_547_U71,
    new_P3_ADD_547_U72, new_P3_ADD_547_U73, new_P3_ADD_547_U74,
    new_P3_ADD_547_U75, new_P3_ADD_547_U76, new_P3_ADD_547_U77,
    new_P3_ADD_547_U78, new_P3_ADD_547_U79, new_P3_ADD_547_U80,
    new_P3_ADD_547_U81, new_P3_ADD_547_U82, new_P3_ADD_547_U83,
    new_P3_ADD_547_U84, new_P3_ADD_547_U85, new_P3_ADD_547_U86,
    new_P3_ADD_547_U87, new_P3_ADD_547_U88, new_P3_ADD_547_U89,
    new_P3_ADD_547_U90, new_P3_ADD_547_U91, new_P3_ADD_547_U92,
    new_P3_ADD_547_U93, new_P3_ADD_547_U94, new_P3_ADD_547_U95,
    new_P3_ADD_547_U96, new_P3_ADD_547_U97, new_P3_ADD_547_U98,
    new_P3_ADD_547_U99, new_P3_ADD_547_U100, new_P3_ADD_547_U101,
    new_P3_ADD_547_U102, new_P3_ADD_547_U103, new_P3_ADD_547_U104,
    new_P3_ADD_547_U105, new_P3_ADD_547_U106, new_P3_ADD_547_U107,
    new_P3_ADD_547_U108, new_P3_ADD_547_U109, new_P3_ADD_547_U110,
    new_P3_ADD_547_U111, new_P3_ADD_547_U112, new_P3_ADD_547_U113,
    new_P3_ADD_547_U114, new_P3_ADD_547_U115, new_P3_ADD_547_U116,
    new_P3_ADD_547_U117, new_P3_ADD_547_U118, new_P3_ADD_547_U119,
    new_P3_ADD_547_U120, new_P3_ADD_547_U121, new_P3_ADD_547_U122,
    new_P3_ADD_547_U123, new_P3_ADD_547_U124, new_P3_ADD_547_U125,
    new_P3_ADD_547_U126, new_P3_ADD_547_U127, new_P3_ADD_547_U128,
    new_P3_ADD_547_U129, new_P3_ADD_547_U130, new_P3_ADD_547_U131,
    new_P3_ADD_547_U132, new_P3_ADD_547_U133, new_P3_ADD_547_U134,
    new_P3_ADD_547_U135, new_P3_ADD_547_U136, new_P3_ADD_547_U137,
    new_P3_ADD_547_U138, new_P3_ADD_547_U139, new_P3_ADD_547_U140,
    new_P3_ADD_547_U141, new_P3_ADD_547_U142, new_P3_ADD_547_U143,
    new_P3_ADD_547_U144, new_P3_ADD_547_U145, new_P3_ADD_547_U146,
    new_P3_ADD_547_U147, new_P3_ADD_547_U148, new_P3_ADD_547_U149,
    new_P3_ADD_547_U150, new_P3_ADD_547_U151, new_P3_ADD_547_U152,
    new_P3_ADD_547_U153, new_P3_ADD_547_U154, new_P3_ADD_547_U155,
    new_P3_ADD_547_U156, new_P3_ADD_547_U157, new_P3_ADD_547_U158,
    new_P3_ADD_547_U159, new_P3_ADD_547_U160, new_P3_ADD_547_U161,
    new_P3_ADD_547_U162, new_P3_ADD_547_U163, new_P3_ADD_547_U164,
    new_P3_ADD_547_U165, new_P3_ADD_547_U166, new_P3_ADD_547_U167,
    new_P3_ADD_547_U168, new_P3_ADD_547_U169, new_P3_ADD_547_U170,
    new_P3_ADD_547_U171, new_P3_ADD_547_U172, new_P3_ADD_547_U173,
    new_P3_ADD_547_U174, new_P3_ADD_547_U175, new_P3_ADD_547_U176,
    new_P3_ADD_547_U177, new_P3_ADD_547_U178, new_P3_ADD_547_U179,
    new_P3_ADD_547_U180, new_P3_ADD_547_U181, new_P3_ADD_547_U182,
    new_P3_ADD_547_U183, new_P3_ADD_547_U184, new_P3_ADD_547_U185,
    new_P3_ADD_547_U186, new_P3_ADD_547_U187, new_P3_ADD_547_U188,
    new_P3_ADD_547_U189, new_P3_SUB_412_U6, new_P3_SUB_412_U7,
    new_P3_SUB_412_U8, new_P3_SUB_412_U9, new_P3_SUB_412_U10,
    new_P3_SUB_412_U11, new_P3_SUB_412_U12, new_P3_SUB_412_U13,
    new_P3_SUB_412_U14, new_P3_SUB_412_U15, new_P3_SUB_412_U16,
    new_P3_SUB_412_U17, new_P3_SUB_412_U18, new_P3_SUB_412_U19,
    new_P3_SUB_412_U20, new_P3_SUB_412_U21, new_P3_SUB_412_U22,
    new_P3_SUB_412_U23, new_P3_SUB_412_U24, new_P3_SUB_412_U25,
    new_P3_SUB_412_U26, new_P3_SUB_412_U27, new_P3_SUB_412_U28,
    new_P3_SUB_412_U29, new_P3_SUB_412_U30, new_P3_SUB_412_U31,
    new_P3_SUB_412_U32, new_P3_SUB_412_U33, new_P3_SUB_412_U34,
    new_P3_SUB_412_U35, new_P3_SUB_412_U36, new_P3_SUB_412_U37,
    new_P3_SUB_412_U38, new_P3_SUB_412_U39, new_P3_SUB_412_U40,
    new_P3_SUB_412_U41, new_P3_SUB_412_U42, new_P3_SUB_412_U43,
    new_P3_SUB_412_U44, new_P3_SUB_412_U45, new_P3_SUB_412_U46,
    new_P3_SUB_412_U47, new_P3_SUB_412_U48, new_P3_SUB_412_U49,
    new_P3_SUB_412_U50, new_P3_SUB_412_U51, new_P3_SUB_412_U52,
    new_P3_SUB_412_U53, new_P3_SUB_412_U54, new_P3_SUB_412_U55,
    new_P3_SUB_412_U56, new_P3_SUB_412_U57, new_P3_SUB_412_U58,
    new_P3_SUB_412_U59, new_P3_SUB_412_U60, new_P3_SUB_412_U61,
    new_P3_SUB_412_U62, new_P3_SUB_412_U63, new_P3_ADD_371_1212_U4,
    new_P3_ADD_371_1212_U5, new_P3_ADD_371_1212_U6, new_P3_ADD_371_1212_U7,
    new_P3_ADD_371_1212_U8, new_P3_ADD_371_1212_U9,
    new_P3_ADD_371_1212_U10, new_P3_ADD_371_1212_U11,
    new_P3_ADD_371_1212_U12, new_P3_ADD_371_1212_U13,
    new_P3_ADD_371_1212_U14, new_P3_ADD_371_1212_U15,
    new_P3_ADD_371_1212_U16, new_P3_ADD_371_1212_U17,
    new_P3_ADD_371_1212_U18, new_P3_ADD_371_1212_U19,
    new_P3_ADD_371_1212_U20, new_P3_ADD_371_1212_U21,
    new_P3_ADD_371_1212_U22, new_P3_ADD_371_1212_U23,
    new_P3_ADD_371_1212_U24, new_P3_ADD_371_1212_U25,
    new_P3_ADD_371_1212_U26, new_P3_ADD_371_1212_U27,
    new_P3_ADD_371_1212_U28, new_P3_ADD_371_1212_U29,
    new_P3_ADD_371_1212_U30, new_P3_ADD_371_1212_U31,
    new_P3_ADD_371_1212_U32, new_P3_ADD_371_1212_U33,
    new_P3_ADD_371_1212_U34, new_P3_ADD_371_1212_U35,
    new_P3_ADD_371_1212_U36, new_P3_ADD_371_1212_U37,
    new_P3_ADD_371_1212_U38, new_P3_ADD_371_1212_U39,
    new_P3_ADD_371_1212_U40, new_P3_ADD_371_1212_U41,
    new_P3_ADD_371_1212_U42, new_P3_ADD_371_1212_U43,
    new_P3_ADD_371_1212_U44, new_P3_ADD_371_1212_U45,
    new_P3_ADD_371_1212_U46, new_P3_ADD_371_1212_U47,
    new_P3_ADD_371_1212_U48, new_P3_ADD_371_1212_U49,
    new_P3_ADD_371_1212_U50, new_P3_ADD_371_1212_U51,
    new_P3_ADD_371_1212_U52, new_P3_ADD_371_1212_U53,
    new_P3_ADD_371_1212_U54, new_P3_ADD_371_1212_U55,
    new_P3_ADD_371_1212_U56, new_P3_ADD_371_1212_U57,
    new_P3_ADD_371_1212_U58, new_P3_ADD_371_1212_U59,
    new_P3_ADD_371_1212_U60, new_P3_ADD_371_1212_U61,
    new_P3_ADD_371_1212_U62, new_P3_ADD_371_1212_U63,
    new_P3_ADD_371_1212_U64, new_P3_ADD_371_1212_U65,
    new_P3_ADD_371_1212_U66, new_P3_ADD_371_1212_U67,
    new_P3_ADD_371_1212_U68, new_P3_ADD_371_1212_U69,
    new_P3_ADD_371_1212_U70, new_P3_ADD_371_1212_U71,
    new_P3_ADD_371_1212_U72, new_P3_ADD_371_1212_U73,
    new_P3_ADD_371_1212_U74, new_P3_ADD_371_1212_U75,
    new_P3_ADD_371_1212_U76, new_P3_ADD_371_1212_U77,
    new_P3_ADD_371_1212_U78, new_P3_ADD_371_1212_U79,
    new_P3_ADD_371_1212_U80, new_P3_ADD_371_1212_U81,
    new_P3_ADD_371_1212_U82, new_P3_ADD_371_1212_U83,
    new_P3_ADD_371_1212_U84, new_P3_ADD_371_1212_U85,
    new_P3_ADD_371_1212_U86, new_P3_ADD_371_1212_U87,
    new_P3_ADD_371_1212_U88, new_P3_ADD_371_1212_U89,
    new_P3_ADD_371_1212_U90, new_P3_ADD_371_1212_U91,
    new_P3_ADD_371_1212_U92, new_P3_ADD_371_1212_U93,
    new_P3_ADD_371_1212_U94, new_P3_ADD_371_1212_U95,
    new_P3_ADD_371_1212_U96, new_P3_ADD_371_1212_U97,
    new_P3_ADD_371_1212_U98, new_P3_ADD_371_1212_U99,
    new_P3_ADD_371_1212_U100, new_P3_ADD_371_1212_U101,
    new_P3_ADD_371_1212_U102, new_P3_ADD_371_1212_U103,
    new_P3_ADD_371_1212_U104, new_P3_ADD_371_1212_U105,
    new_P3_ADD_371_1212_U106, new_P3_ADD_371_1212_U107,
    new_P3_ADD_371_1212_U108, new_P3_ADD_371_1212_U109,
    new_P3_ADD_371_1212_U110, new_P3_ADD_371_1212_U111,
    new_P3_ADD_371_1212_U112, new_P3_ADD_371_1212_U113,
    new_P3_ADD_371_1212_U114, new_P3_ADD_371_1212_U115,
    new_P3_ADD_371_1212_U116, new_P3_ADD_371_1212_U117,
    new_P3_ADD_371_1212_U118, new_P3_ADD_371_1212_U119,
    new_P3_ADD_371_1212_U120, new_P3_ADD_371_1212_U121,
    new_P3_ADD_371_1212_U122, new_P3_ADD_371_1212_U123,
    new_P3_ADD_371_1212_U124, new_P3_ADD_371_1212_U125,
    new_P3_ADD_371_1212_U126, new_P3_ADD_371_1212_U127,
    new_P3_ADD_371_1212_U128, new_P3_ADD_371_1212_U129,
    new_P3_ADD_371_1212_U130, new_P3_ADD_371_1212_U131,
    new_P3_ADD_371_1212_U132, new_P3_ADD_371_1212_U133,
    new_P3_ADD_371_1212_U134, new_P3_ADD_371_1212_U135,
    new_P3_ADD_371_1212_U136, new_P3_ADD_371_1212_U137,
    new_P3_ADD_371_1212_U138, new_P3_ADD_371_1212_U139,
    new_P3_ADD_371_1212_U140, new_P3_ADD_371_1212_U141,
    new_P3_ADD_371_1212_U142, new_P3_ADD_371_1212_U143,
    new_P3_ADD_371_1212_U144, new_P3_ADD_371_1212_U145,
    new_P3_ADD_371_1212_U146, new_P3_ADD_371_1212_U147,
    new_P3_ADD_371_1212_U148, new_P3_ADD_371_1212_U149,
    new_P3_ADD_371_1212_U150, new_P3_ADD_371_1212_U151,
    new_P3_ADD_371_1212_U152, new_P3_ADD_371_1212_U153,
    new_P3_ADD_371_1212_U154, new_P3_ADD_371_1212_U155,
    new_P3_ADD_371_1212_U156, new_P3_ADD_371_1212_U157,
    new_P3_ADD_371_1212_U158, new_P3_ADD_371_1212_U159,
    new_P3_ADD_371_1212_U160, new_P3_ADD_371_1212_U161,
    new_P3_ADD_371_1212_U162, new_P3_ADD_371_1212_U163,
    new_P3_ADD_371_1212_U164, new_P3_ADD_371_1212_U165,
    new_P3_ADD_371_1212_U166, new_P3_ADD_371_1212_U167,
    new_P3_ADD_371_1212_U168, new_P3_ADD_371_1212_U169,
    new_P3_ADD_371_1212_U170, new_P3_ADD_371_1212_U171,
    new_P3_ADD_371_1212_U172, new_P3_ADD_371_1212_U173,
    new_P3_ADD_371_1212_U174, new_P3_ADD_371_1212_U175,
    new_P3_ADD_371_1212_U176, new_P3_ADD_371_1212_U177,
    new_P3_ADD_371_1212_U178, new_P3_ADD_371_1212_U179,
    new_P3_ADD_371_1212_U180, new_P3_ADD_371_1212_U181,
    new_P3_ADD_371_1212_U182, new_P3_ADD_371_1212_U183,
    new_P3_ADD_371_1212_U184, new_P3_ADD_371_1212_U185,
    new_P3_ADD_371_1212_U186, new_P3_ADD_371_1212_U187,
    new_P3_ADD_371_1212_U188, new_P3_ADD_371_1212_U189,
    new_P3_ADD_371_1212_U190, new_P3_ADD_371_1212_U191,
    new_P3_ADD_371_1212_U192, new_P3_ADD_371_1212_U193,
    new_P3_ADD_371_1212_U194, new_P3_ADD_371_1212_U195,
    new_P3_ADD_371_1212_U196, new_P3_ADD_371_1212_U197,
    new_P3_ADD_371_1212_U198, new_P3_ADD_371_1212_U199,
    new_P3_ADD_371_1212_U200, new_P3_ADD_371_1212_U201,
    new_P3_ADD_371_1212_U202, new_P3_ADD_371_1212_U203,
    new_P3_ADD_371_1212_U204, new_P3_ADD_371_1212_U205,
    new_P3_ADD_371_1212_U206, new_P3_ADD_371_1212_U207,
    new_P3_ADD_371_1212_U208, new_P3_ADD_371_1212_U209,
    new_P3_ADD_371_1212_U210, new_P3_ADD_371_1212_U211,
    new_P3_ADD_371_1212_U212, new_P3_ADD_371_1212_U213,
    new_P3_ADD_371_1212_U214, new_P3_ADD_371_1212_U215,
    new_P3_ADD_371_1212_U216, new_P3_ADD_371_1212_U217,
    new_P3_ADD_371_1212_U218, new_P3_ADD_371_1212_U219,
    new_P3_ADD_371_1212_U220, new_P3_ADD_371_1212_U221,
    new_P3_ADD_371_1212_U222, new_P3_ADD_371_1212_U223,
    new_P3_ADD_371_1212_U224, new_P3_ADD_371_1212_U225,
    new_P3_ADD_371_1212_U226, new_P3_ADD_371_1212_U227,
    new_P3_ADD_371_1212_U228, new_P3_ADD_371_1212_U229,
    new_P3_ADD_371_1212_U230, new_P3_ADD_371_1212_U231,
    new_P3_ADD_371_1212_U232, new_P3_ADD_371_1212_U233,
    new_P3_ADD_371_1212_U234, new_P3_ADD_371_1212_U235,
    new_P3_ADD_371_1212_U236, new_P3_ADD_371_1212_U237,
    new_P3_ADD_371_1212_U238, new_P3_ADD_371_1212_U239,
    new_P3_ADD_371_1212_U240, new_P3_ADD_371_1212_U241,
    new_P3_ADD_371_1212_U242, new_P3_ADD_371_1212_U243,
    new_P3_ADD_371_1212_U244, new_P3_ADD_371_1212_U245,
    new_P3_ADD_371_1212_U246, new_P3_ADD_371_1212_U247,
    new_P3_ADD_371_1212_U248, new_P3_ADD_371_1212_U249,
    new_P3_ADD_371_1212_U250, new_P3_ADD_371_1212_U251,
    new_P3_ADD_371_1212_U252, new_P3_ADD_371_1212_U253,
    new_P3_ADD_371_1212_U254, new_P3_ADD_371_1212_U255,
    new_P3_ADD_371_1212_U256, new_P3_ADD_371_1212_U257,
    new_P3_ADD_371_1212_U258, new_P3_ADD_371_1212_U259,
    new_P3_ADD_371_1212_U260, new_P3_ADD_371_1212_U261,
    new_P3_ADD_371_1212_U262, new_P3_ADD_371_1212_U263,
    new_P3_ADD_371_1212_U264, new_P3_ADD_371_1212_U265, new_P3_SUB_504_U6,
    new_P3_SUB_504_U7, new_P3_SUB_504_U8, new_P3_SUB_504_U9,
    new_P3_SUB_504_U10, new_P3_SUB_504_U11, new_P3_SUB_504_U12,
    new_P3_SUB_504_U13, new_P3_SUB_504_U14, new_P3_SUB_504_U15,
    new_P3_SUB_504_U16, new_P3_SUB_504_U17, new_P3_SUB_504_U18,
    new_P3_SUB_504_U19, new_P3_SUB_504_U20, new_P3_SUB_504_U21,
    new_P3_SUB_504_U22, new_P3_SUB_504_U23, new_P3_SUB_504_U24,
    new_P3_SUB_504_U25, new_P3_SUB_504_U26, new_P3_SUB_504_U27,
    new_P3_SUB_504_U28, new_P3_SUB_504_U29, new_P3_SUB_504_U30,
    new_P3_SUB_504_U31, new_P3_SUB_504_U32, new_P3_SUB_504_U33,
    new_P3_SUB_504_U34, new_P3_SUB_504_U35, new_P3_SUB_504_U36,
    new_P3_SUB_504_U37, new_P3_SUB_504_U38, new_P3_SUB_504_U39,
    new_P3_SUB_504_U40, new_P3_SUB_504_U41, new_P3_SUB_504_U42,
    new_P3_SUB_504_U43, new_P3_SUB_504_U44, new_P3_SUB_504_U45,
    new_P3_SUB_504_U46, new_P3_SUB_504_U47, new_P3_SUB_504_U48,
    new_P3_SUB_504_U49, new_P3_SUB_504_U50, new_P3_SUB_504_U51,
    new_P3_SUB_504_U52, new_P3_SUB_504_U53, new_P3_SUB_504_U54,
    new_P3_SUB_504_U55, new_P3_SUB_504_U56, new_P3_SUB_504_U57,
    new_P3_SUB_504_U58, new_P3_SUB_504_U59, new_P3_SUB_504_U60,
    new_P3_SUB_504_U61, new_P3_SUB_504_U62, new_P3_SUB_504_U63,
    new_P3_SUB_401_U6, new_P3_SUB_401_U7, new_P3_SUB_401_U8,
    new_P3_SUB_401_U9, new_P3_SUB_401_U10, new_P3_SUB_401_U11,
    new_P3_SUB_401_U12, new_P3_SUB_401_U13, new_P3_SUB_401_U14,
    new_P3_SUB_401_U15, new_P3_SUB_401_U16, new_P3_SUB_401_U17,
    new_P3_SUB_401_U18, new_P3_SUB_401_U19, new_P3_SUB_401_U20,
    new_P3_SUB_401_U21, new_P3_SUB_401_U22, new_P3_SUB_401_U23,
    new_P3_SUB_401_U24, new_P3_SUB_401_U25, new_P3_SUB_401_U26,
    new_P3_SUB_401_U27, new_P3_SUB_401_U28, new_P3_SUB_401_U29,
    new_P3_SUB_401_U30, new_P3_SUB_401_U31, new_P3_SUB_401_U32,
    new_P3_SUB_401_U33, new_P3_SUB_401_U34, new_P3_SUB_401_U35,
    new_P3_SUB_401_U36, new_P3_SUB_401_U37, new_P3_SUB_401_U38,
    new_P3_SUB_401_U39, new_P3_SUB_401_U40, new_P3_SUB_401_U41,
    new_P3_SUB_401_U42, new_P3_SUB_401_U43, new_P3_SUB_401_U44,
    new_P3_SUB_401_U45, new_P3_SUB_401_U46, new_P3_SUB_401_U47,
    new_P3_SUB_401_U48, new_P3_SUB_401_U49, new_P3_SUB_401_U50,
    new_P3_SUB_401_U51, new_P3_SUB_401_U52, new_P3_SUB_401_U53,
    new_P3_SUB_401_U54, new_P3_SUB_401_U55, new_P3_SUB_401_U56,
    new_P3_SUB_401_U57, new_P3_SUB_401_U58, new_P3_SUB_401_U59,
    new_P3_SUB_401_U60, new_P3_SUB_401_U61, new_P3_SUB_401_U62,
    new_P3_SUB_401_U63, new_P3_SUB_401_U64, new_P3_SUB_401_U65,
    new_P3_SUB_401_U66, new_P3_ADD_371_U4, new_P3_ADD_371_U5,
    new_P3_ADD_371_U6, new_P3_ADD_371_U7, new_P3_ADD_371_U8,
    new_P3_ADD_371_U9, new_P3_ADD_371_U10, new_P3_ADD_371_U11,
    new_P3_ADD_371_U12, new_P3_ADD_371_U13, new_P3_ADD_371_U14,
    new_P3_ADD_371_U15, new_P3_ADD_371_U16, new_P3_ADD_371_U17,
    new_P3_ADD_371_U18, new_P3_ADD_371_U19, new_P3_ADD_371_U20,
    new_P3_ADD_371_U21, new_P3_ADD_371_U22, new_P3_ADD_371_U23,
    new_P3_ADD_371_U24, new_P3_ADD_371_U25, new_P3_ADD_371_U26,
    new_P3_ADD_371_U27, new_P3_ADD_371_U28, new_P3_ADD_371_U29,
    new_P3_ADD_371_U30, new_P3_ADD_371_U31, new_P3_ADD_371_U32,
    new_P3_ADD_371_U33, new_P3_ADD_371_U34, new_P3_ADD_371_U35,
    new_P3_ADD_371_U36, new_P3_ADD_371_U37, new_P3_ADD_371_U38,
    new_P3_ADD_371_U39, new_P3_ADD_371_U40, new_P3_ADD_371_U41,
    new_P3_ADD_371_U42, new_P3_ADD_371_U43, new_P3_ADD_371_U44,
    new_P3_SUB_390_U6, new_P3_SUB_390_U7, new_P3_SUB_390_U8,
    new_P3_SUB_390_U9, new_P3_SUB_390_U10, new_P3_SUB_390_U11,
    new_P3_SUB_390_U12, new_P3_SUB_390_U13, new_P3_SUB_390_U14,
    new_P3_SUB_390_U15, new_P3_SUB_390_U16, new_P3_SUB_390_U17,
    new_P3_SUB_390_U18, new_P3_SUB_390_U19, new_P3_SUB_390_U20,
    new_P3_SUB_390_U21, new_P3_SUB_390_U22, new_P3_SUB_390_U23,
    new_P3_SUB_390_U24, new_P3_SUB_390_U25, new_P3_SUB_390_U26,
    new_P3_SUB_390_U27, new_P3_SUB_390_U28, new_P3_SUB_390_U29,
    new_P3_SUB_390_U30, new_P3_SUB_390_U31, new_P3_SUB_390_U32,
    new_P3_SUB_390_U33, new_P3_SUB_390_U34, new_P3_SUB_390_U35,
    new_P3_SUB_390_U36, new_P3_SUB_390_U37, new_P3_SUB_390_U38,
    new_P3_SUB_390_U39, new_P3_SUB_390_U40, new_P3_SUB_390_U41,
    new_P3_SUB_390_U42, new_P3_SUB_390_U43, new_P3_SUB_390_U44,
    new_P3_SUB_390_U45, new_P3_SUB_390_U46, new_P3_SUB_390_U47,
    new_P3_SUB_390_U48, new_P3_SUB_390_U49, new_P3_SUB_390_U50,
    new_P3_SUB_390_U51, new_P3_SUB_390_U52, new_P3_SUB_390_U53,
    new_P3_SUB_390_U54, new_P3_SUB_390_U55, new_P3_SUB_390_U56,
    new_P3_SUB_390_U57, new_P3_SUB_390_U58, new_P3_SUB_390_U59,
    new_P3_SUB_390_U60, new_P3_SUB_390_U61, new_P3_SUB_390_U62,
    new_P3_SUB_390_U63, new_P3_SUB_390_U64, new_P3_SUB_390_U65,
    new_P3_SUB_390_U66, new_P3_SUB_357_U6, new_P3_SUB_357_U7,
    new_P3_SUB_357_U8, new_P3_SUB_357_U9, new_P3_SUB_357_U10,
    new_P3_SUB_357_U11, new_P3_SUB_357_U12, new_P3_SUB_357_U13,
    new_P3_ADD_495_U4, new_P3_ADD_495_U5, new_P3_ADD_495_U6,
    new_P3_ADD_495_U7, new_P3_ADD_495_U8, new_P3_ADD_495_U9,
    new_P3_ADD_495_U10, new_P3_ADD_495_U11, new_P3_ADD_495_U12,
    new_P3_ADD_495_U13, new_P3_ADD_495_U14, new_P3_ADD_495_U15,
    new_P3_ADD_495_U16, new_P3_ADD_495_U17, new_P3_ADD_495_U18,
    new_P3_ADD_495_U19, new_P3_ADD_495_U20, new_P3_GTE_412_U6,
    new_P3_GTE_412_U7, new_P3_GTE_504_U6, new_P3_GTE_504_U7,
    new_P3_ADD_494_U4, new_P3_ADD_494_U5, new_P3_ADD_494_U6,
    new_P3_ADD_494_U7, new_P3_ADD_494_U8, new_P3_ADD_494_U9,
    new_P3_ADD_494_U10, new_P3_ADD_494_U11, new_P3_ADD_494_U12,
    new_P3_ADD_494_U13, new_P3_ADD_494_U14, new_P3_ADD_494_U15,
    new_P3_ADD_494_U16, new_P3_ADD_494_U17, new_P3_ADD_494_U18,
    new_P3_ADD_494_U19, new_P3_ADD_494_U20, new_P3_ADD_494_U21,
    new_P3_ADD_494_U22, new_P3_ADD_494_U23, new_P3_ADD_494_U24,
    new_P3_ADD_494_U25, new_P3_ADD_494_U26, new_P3_ADD_494_U27,
    new_P3_ADD_494_U28, new_P3_ADD_494_U29, new_P3_ADD_494_U30,
    new_P3_ADD_494_U31, new_P3_ADD_494_U32, new_P3_ADD_494_U33,
    new_P3_ADD_494_U34, new_P3_ADD_494_U35, new_P3_ADD_494_U36,
    new_P3_ADD_494_U37, new_P3_ADD_494_U38, new_P3_ADD_494_U39,
    new_P3_ADD_494_U40, new_P3_ADD_494_U41, new_P3_ADD_494_U42,
    new_P3_ADD_494_U43, new_P3_ADD_494_U44, new_P3_ADD_494_U45,
    new_P3_ADD_494_U46, new_P3_ADD_494_U47, new_P3_ADD_494_U48,
    new_P3_ADD_494_U49, new_P3_ADD_494_U50, new_P3_ADD_494_U51,
    new_P3_ADD_494_U52, new_P3_ADD_494_U53, new_P3_ADD_494_U54,
    new_P3_ADD_494_U55, new_P3_ADD_494_U56, new_P3_ADD_494_U57,
    new_P3_ADD_494_U58, new_P3_ADD_494_U59, new_P3_ADD_494_U60,
    new_P3_ADD_494_U61, new_P3_ADD_494_U62, new_P3_ADD_494_U63,
    new_P3_ADD_494_U64, new_P3_ADD_494_U65, new_P3_ADD_494_U66,
    new_P3_ADD_494_U67, new_P3_ADD_494_U68, new_P3_ADD_494_U69,
    new_P3_ADD_494_U70, new_P3_ADD_494_U71, new_P3_ADD_494_U72,
    new_P3_ADD_494_U73, new_P3_ADD_494_U74, new_P3_ADD_494_U75,
    new_P3_ADD_494_U76, new_P3_ADD_494_U77, new_P3_ADD_494_U78,
    new_P3_ADD_494_U79, new_P3_ADD_494_U80, new_P3_ADD_494_U81,
    new_P3_ADD_494_U82, new_P3_ADD_494_U83, new_P3_ADD_494_U84,
    new_P3_ADD_494_U85, new_P3_ADD_494_U86, new_P3_ADD_494_U87,
    new_P3_ADD_494_U88, new_P3_ADD_494_U89, new_P3_ADD_494_U90,
    new_P3_ADD_494_U91, new_P3_ADD_494_U92, new_P3_ADD_494_U93,
    new_P3_ADD_494_U94, new_P3_ADD_494_U95, new_P3_ADD_494_U96,
    new_P3_ADD_494_U97, new_P3_ADD_494_U98, new_P3_ADD_494_U99,
    new_P3_ADD_494_U100, new_P3_ADD_494_U101, new_P3_ADD_494_U102,
    new_P3_ADD_494_U103, new_P3_ADD_494_U104, new_P3_ADD_494_U105,
    new_P3_ADD_494_U106, new_P3_ADD_494_U107, new_P3_ADD_494_U108,
    new_P3_ADD_494_U109, new_P3_ADD_494_U110, new_P3_ADD_494_U111,
    new_P3_ADD_494_U112, new_P3_ADD_494_U113, new_P3_ADD_494_U114,
    new_P3_ADD_494_U115, new_P3_ADD_494_U116, new_P3_ADD_494_U117,
    new_P3_ADD_494_U118, new_P3_ADD_494_U119, new_P3_ADD_494_U120,
    new_P3_ADD_494_U121, new_P3_ADD_494_U122, new_P3_ADD_494_U123,
    new_P3_ADD_494_U124, new_P3_ADD_494_U125, new_P3_ADD_494_U126,
    new_P3_ADD_494_U127, new_P3_ADD_494_U128, new_P3_ADD_494_U129,
    new_P3_ADD_494_U130, new_P3_ADD_494_U131, new_P3_ADD_494_U132,
    new_P3_ADD_494_U133, new_P3_ADD_494_U134, new_P3_ADD_494_U135,
    new_P3_ADD_494_U136, new_P3_ADD_494_U137, new_P3_ADD_494_U138,
    new_P3_ADD_494_U139, new_P3_ADD_494_U140, new_P3_ADD_494_U141,
    new_P3_ADD_494_U142, new_P3_ADD_494_U143, new_P3_ADD_494_U144,
    new_P3_ADD_494_U145, new_P3_ADD_494_U146, new_P3_ADD_494_U147,
    new_P3_ADD_494_U148, new_P3_ADD_494_U149, new_P3_ADD_494_U150,
    new_P3_ADD_494_U151, new_P3_ADD_494_U152, new_P3_ADD_494_U153,
    new_P3_ADD_494_U154, new_P3_ADD_494_U155, new_P3_ADD_494_U156,
    new_P3_ADD_494_U157, new_P3_ADD_494_U158, new_P3_ADD_494_U159,
    new_P3_ADD_494_U160, new_P3_ADD_494_U161, new_P3_ADD_494_U162,
    new_P3_ADD_494_U163, new_P3_ADD_494_U164, new_P3_ADD_494_U165,
    new_P3_ADD_494_U166, new_P3_ADD_494_U167, new_P3_ADD_494_U168,
    new_P3_ADD_494_U169, new_P3_ADD_494_U170, new_P3_ADD_494_U171,
    new_P3_ADD_494_U172, new_P3_ADD_494_U173, new_P3_ADD_494_U174,
    new_P3_ADD_494_U175, new_P3_ADD_494_U176, new_P3_ADD_494_U177,
    new_P3_ADD_494_U178, new_P3_ADD_494_U179, new_P3_ADD_494_U180,
    new_P3_ADD_494_U181, new_P3_ADD_494_U182, new_P3_ADD_536_U4,
    new_P3_ADD_536_U5, new_P3_ADD_536_U6, new_P3_ADD_536_U7,
    new_P3_ADD_536_U8, new_P3_ADD_536_U9, new_P3_ADD_536_U10,
    new_P3_ADD_536_U11, new_P3_ADD_536_U12, new_P3_ADD_536_U13,
    new_P3_ADD_536_U14, new_P3_ADD_536_U15, new_P3_ADD_536_U16,
    new_P3_ADD_536_U17, new_P3_ADD_536_U18, new_P3_ADD_536_U19,
    new_P3_ADD_536_U20, new_P3_ADD_536_U21, new_P3_ADD_536_U22,
    new_P3_ADD_536_U23, new_P3_ADD_536_U24, new_P3_ADD_536_U25,
    new_P3_ADD_536_U26, new_P3_ADD_536_U27, new_P3_ADD_536_U28,
    new_P3_ADD_536_U29, new_P3_ADD_536_U30, new_P3_ADD_536_U31,
    new_P3_ADD_536_U32, new_P3_ADD_536_U33, new_P3_ADD_536_U34,
    new_P3_ADD_536_U35, new_P3_ADD_536_U36, new_P3_ADD_536_U37,
    new_P3_ADD_536_U38, new_P3_ADD_536_U39, new_P3_ADD_536_U40,
    new_P3_ADD_536_U41, new_P3_ADD_536_U42, new_P3_ADD_536_U43,
    new_P3_ADD_536_U44, new_P3_ADD_536_U45, new_P3_ADD_536_U46,
    new_P3_ADD_536_U47, new_P3_ADD_536_U48, new_P3_ADD_536_U49,
    new_P3_ADD_536_U50, new_P3_ADD_536_U51, new_P3_ADD_536_U52,
    new_P3_ADD_536_U53, new_P3_ADD_536_U54, new_P3_ADD_536_U55,
    new_P3_ADD_536_U56, new_P3_ADD_536_U57, new_P3_ADD_536_U58,
    new_P3_ADD_536_U59, new_P3_ADD_536_U60, new_P3_ADD_536_U61,
    new_P3_ADD_536_U62, new_P3_ADD_536_U63, new_P3_ADD_536_U64,
    new_P3_ADD_536_U65, new_P3_ADD_536_U66, new_P3_ADD_536_U67,
    new_P3_ADD_536_U68, new_P3_ADD_536_U69, new_P3_ADD_536_U70,
    new_P3_ADD_536_U71, new_P3_ADD_536_U72, new_P3_ADD_536_U73,
    new_P3_ADD_536_U74, new_P3_ADD_536_U75, new_P3_ADD_536_U76,
    new_P3_ADD_536_U77, new_P3_ADD_536_U78, new_P3_ADD_536_U79,
    new_P3_ADD_536_U80, new_P3_ADD_536_U81, new_P3_ADD_536_U82,
    new_P3_ADD_536_U83, new_P3_ADD_536_U84, new_P3_ADD_536_U85,
    new_P3_ADD_536_U86, new_P3_ADD_536_U87, new_P3_ADD_536_U88,
    new_P3_ADD_536_U89, new_P3_ADD_536_U90, new_P3_ADD_536_U91,
    new_P3_ADD_536_U92, new_P3_ADD_536_U93, new_P3_ADD_536_U94,
    new_P3_ADD_536_U95, new_P3_ADD_536_U96, new_P3_ADD_536_U97,
    new_P3_ADD_536_U98, new_P3_ADD_536_U99, new_P3_ADD_536_U100,
    new_P3_ADD_536_U101, new_P3_ADD_536_U102, new_P3_ADD_536_U103,
    new_P3_ADD_536_U104, new_P3_ADD_536_U105, new_P3_ADD_536_U106,
    new_P3_ADD_536_U107, new_P3_ADD_536_U108, new_P3_ADD_536_U109,
    new_P3_ADD_536_U110, new_P3_ADD_536_U111, new_P3_ADD_536_U112,
    new_P3_ADD_536_U113, new_P3_ADD_536_U114, new_P3_ADD_536_U115,
    new_P3_ADD_536_U116, new_P3_ADD_536_U117, new_P3_ADD_536_U118,
    new_P3_ADD_536_U119, new_P3_ADD_536_U120, new_P3_ADD_536_U121,
    new_P3_ADD_536_U122, new_P3_ADD_536_U123, new_P3_ADD_536_U124,
    new_P3_ADD_536_U125, new_P3_ADD_536_U126, new_P3_ADD_536_U127,
    new_P3_ADD_536_U128, new_P3_ADD_536_U129, new_P3_ADD_536_U130,
    new_P3_ADD_536_U131, new_P3_ADD_536_U132, new_P3_ADD_536_U133,
    new_P3_ADD_536_U134, new_P3_ADD_536_U135, new_P3_ADD_536_U136,
    new_P3_ADD_536_U137, new_P3_ADD_536_U138, new_P3_ADD_536_U139,
    new_P3_ADD_536_U140, new_P3_ADD_536_U141, new_P3_ADD_536_U142,
    new_P3_ADD_536_U143, new_P3_ADD_536_U144, new_P3_ADD_536_U145,
    new_P3_ADD_536_U146, new_P3_ADD_536_U147, new_P3_ADD_536_U148,
    new_P3_ADD_536_U149, new_P3_ADD_536_U150, new_P3_ADD_536_U151,
    new_P3_ADD_536_U152, new_P3_ADD_536_U153, new_P3_ADD_536_U154,
    new_P3_ADD_536_U155, new_P3_ADD_536_U156, new_P3_ADD_536_U157,
    new_P3_ADD_536_U158, new_P3_ADD_536_U159, new_P3_ADD_536_U160,
    new_P3_ADD_536_U161, new_P3_ADD_536_U162, new_P3_ADD_536_U163,
    new_P3_ADD_536_U164, new_P3_ADD_536_U165, new_P3_ADD_536_U166,
    new_P3_ADD_536_U167, new_P3_ADD_536_U168, new_P3_ADD_536_U169,
    new_P3_ADD_536_U170, new_P3_ADD_536_U171, new_P3_ADD_536_U172,
    new_P3_ADD_536_U173, new_P3_ADD_536_U174, new_P3_ADD_536_U175,
    new_P3_ADD_536_U176, new_P3_ADD_536_U177, new_P3_ADD_536_U178,
    new_P3_ADD_536_U179, new_P3_ADD_536_U180, new_P3_ADD_536_U181,
    new_P3_ADD_536_U182, new_P3_ADD_402_1132_U4, new_P3_ADD_402_1132_U5,
    new_P3_ADD_402_1132_U6, new_P3_ADD_402_1132_U7, new_P3_ADD_402_1132_U8,
    new_P3_ADD_402_1132_U9, new_P3_ADD_402_1132_U10,
    new_P3_ADD_402_1132_U11, new_P3_ADD_402_1132_U12,
    new_P3_ADD_402_1132_U13, new_P3_ADD_402_1132_U14,
    new_P3_ADD_402_1132_U15, new_P3_ADD_402_1132_U16,
    new_P3_ADD_402_1132_U17, new_P3_ADD_402_1132_U18,
    new_P3_ADD_402_1132_U19, new_P3_ADD_402_1132_U20,
    new_P3_ADD_402_1132_U21, new_P3_ADD_402_1132_U22,
    new_P3_ADD_402_1132_U23, new_P3_ADD_402_1132_U24,
    new_P3_ADD_402_1132_U25, new_P3_ADD_402_1132_U26,
    new_P3_ADD_402_1132_U27, new_P3_ADD_402_1132_U28,
    new_P3_ADD_402_1132_U29, new_P3_ADD_402_1132_U30,
    new_P3_ADD_402_1132_U31, new_P3_ADD_402_1132_U32,
    new_P3_ADD_402_1132_U33, new_P3_ADD_402_1132_U34,
    new_P3_ADD_402_1132_U35, new_P3_ADD_402_1132_U36,
    new_P3_ADD_402_1132_U37, new_P3_ADD_402_1132_U38,
    new_P3_ADD_402_1132_U39, new_P3_ADD_402_1132_U40,
    new_P3_ADD_402_1132_U41, new_P3_ADD_402_1132_U42,
    new_P3_ADD_402_1132_U43, new_P3_ADD_402_1132_U44,
    new_P3_ADD_402_1132_U45, new_P3_ADD_402_1132_U46,
    new_P3_ADD_402_1132_U47, new_P3_ADD_402_1132_U48,
    new_P3_ADD_402_1132_U49, new_P3_ADD_402_1132_U50, new_P2_R2099_U5,
    new_P2_R2099_U6, new_P2_R2099_U7, new_P2_R2099_U8, new_P2_R2099_U9,
    new_P2_R2099_U10, new_P2_R2099_U11, new_P2_R2099_U12, new_P2_R2099_U13,
    new_P2_R2099_U14, new_P2_R2099_U15, new_P2_R2099_U16, new_P2_R2099_U17,
    new_P2_R2099_U18, new_P2_R2099_U19, new_P2_R2099_U20, new_P2_R2099_U21,
    new_P2_R2099_U22, new_P2_R2099_U23, new_P2_R2099_U24, new_P2_R2099_U25,
    new_P2_R2099_U26, new_P2_R2099_U27, new_P2_R2099_U28, new_P2_R2099_U29,
    new_P2_R2099_U30, new_P2_R2099_U31, new_P2_R2099_U32, new_P2_R2099_U33,
    new_P2_R2099_U34, new_P2_R2099_U35, new_P2_R2099_U36, new_P2_R2099_U37,
    new_P2_R2099_U38, new_P2_R2099_U39, new_P2_R2099_U40, new_P2_R2099_U41,
    new_P2_R2099_U42, new_P2_R2099_U43, new_P2_R2099_U44, new_P2_R2099_U45,
    new_P2_R2099_U46, new_P2_R2099_U47, new_P2_R2099_U48, new_P2_R2099_U49,
    new_P2_R2099_U50, new_P2_R2099_U51, new_P2_R2099_U52, new_P2_R2099_U53,
    new_P2_R2099_U54, new_P2_R2099_U55, new_P2_R2099_U56, new_P2_R2099_U57,
    new_P2_R2099_U58, new_P2_R2099_U59, new_P2_R2099_U60, new_P2_R2099_U61,
    new_P2_R2099_U62, new_P2_R2099_U63, new_P2_R2099_U64, new_P2_R2099_U65,
    new_P2_R2099_U66, new_P2_R2099_U67, new_P2_R2099_U68, new_P2_R2099_U69,
    new_P2_R2099_U70, new_P2_R2099_U71, new_P2_R2099_U72, new_P2_R2099_U73,
    new_P2_R2099_U74, new_P2_R2099_U75, new_P2_R2099_U76, new_P2_R2099_U77,
    new_P2_R2099_U78, new_P2_R2099_U79, new_P2_R2099_U80, new_P2_R2099_U81,
    new_P2_R2099_U82, new_P2_R2099_U83, new_P2_R2099_U84, new_P2_R2099_U85,
    new_P2_R2099_U86, new_P2_R2099_U87, new_P2_R2099_U88, new_P2_R2099_U89,
    new_P2_R2099_U90, new_P2_R2099_U91, new_P2_R2099_U92, new_P2_R2099_U93,
    new_P2_R2099_U94, new_P2_R2099_U95, new_P2_R2099_U96, new_P2_R2099_U97,
    new_P2_R2099_U98, new_P2_R2099_U99, new_P2_R2099_U100,
    new_P2_R2099_U101, new_P2_R2099_U102, new_P2_R2099_U103,
    new_P2_R2099_U104, new_P2_R2099_U105, new_P2_R2099_U106,
    new_P2_R2099_U107, new_P2_R2099_U108, new_P2_R2099_U109,
    new_P2_R2099_U110, new_P2_R2099_U111, new_P2_R2099_U112,
    new_P2_R2099_U113, new_P2_R2099_U114, new_P2_R2099_U115,
    new_P2_R2099_U116, new_P2_R2099_U117, new_P2_R2099_U118,
    new_P2_R2099_U119, new_P2_R2099_U120, new_P2_R2099_U121,
    new_P2_R2099_U122, new_P2_R2099_U123, new_P2_R2099_U124,
    new_P2_R2099_U125, new_P2_R2099_U126, new_P2_R2099_U127,
    new_P2_R2099_U128, new_P2_R2099_U129, new_P2_R2099_U130,
    new_P2_R2099_U131, new_P2_R2099_U132, new_P2_R2099_U133,
    new_P2_R2099_U134, new_P2_R2099_U135, new_P2_R2099_U136,
    new_P2_R2099_U137, new_P2_R2099_U138, new_P2_R2099_U139,
    new_P2_R2099_U140, new_P2_R2099_U141, new_P2_R2099_U142,
    new_P2_R2099_U143, new_P2_R2099_U144, new_P2_R2099_U145,
    new_P2_R2099_U146, new_P2_R2099_U147, new_P2_R2099_U148,
    new_P2_R2099_U149, new_P2_R2099_U150, new_P2_R2099_U151,
    new_P2_R2099_U152, new_P2_R2099_U153, new_P2_R2099_U154,
    new_P2_R2099_U155, new_P2_R2099_U156, new_P2_R2099_U157,
    new_P2_R2099_U158, new_P2_R2099_U159, new_P2_R2099_U160,
    new_P2_R2099_U161, new_P2_R2099_U162, new_P2_R2099_U163,
    new_P2_R2099_U164, new_P2_R2099_U165, new_P2_R2099_U166,
    new_P2_R2099_U167, new_P2_R2099_U168, new_P2_R2099_U169,
    new_P2_R2099_U170, new_P2_R2099_U171, new_P2_R2099_U172,
    new_P2_R2099_U173, new_P2_R2099_U174, new_P2_R2099_U175,
    new_P2_R2099_U176, new_P2_R2099_U177, new_P2_R2099_U178,
    new_P2_R2099_U179, new_P2_R2099_U180, new_P2_R2099_U181,
    new_P2_R2099_U182, new_P2_R2099_U183, new_P2_R2099_U184,
    new_P2_R2099_U185, new_P2_R2099_U186, new_P2_R2099_U187,
    new_P2_R2099_U188, new_P2_R2099_U189, new_P2_R2099_U190,
    new_P2_R2099_U191, new_P2_R2099_U192, new_P2_R2099_U193,
    new_P2_R2099_U194, new_P2_R2099_U195, new_P2_R2099_U196,
    new_P2_R2099_U197, new_P2_R2099_U198, new_P2_R2099_U199,
    new_P2_R2099_U200, new_P2_R2099_U201, new_P2_R2099_U202,
    new_P2_R2099_U203, new_P2_R2099_U204, new_P2_R2099_U205,
    new_P2_R2099_U206, new_P2_R2099_U207, new_P2_R2099_U208,
    new_P2_R2099_U209, new_P2_R2099_U210, new_P2_R2099_U211,
    new_P2_R2099_U212, new_P2_R2099_U213, new_P2_R2099_U214,
    new_P2_R2099_U215, new_P2_R2099_U216, new_P2_R2099_U217,
    new_P2_R2099_U218, new_P2_R2099_U219, new_P2_R2099_U220,
    new_P2_R2099_U221, new_P2_R2099_U222, new_P2_R2099_U223,
    new_P2_R2099_U224, new_P2_R2099_U225, new_P2_ADD_391_1196_U5,
    new_P2_ADD_391_1196_U6, new_P2_ADD_391_1196_U7, new_P2_ADD_391_1196_U8,
    new_P2_ADD_391_1196_U9, new_P2_ADD_391_1196_U10,
    new_P2_ADD_391_1196_U11, new_P2_ADD_391_1196_U12,
    new_P2_ADD_391_1196_U13, new_P2_ADD_391_1196_U14,
    new_P2_ADD_391_1196_U15, new_P2_ADD_391_1196_U16,
    new_P2_ADD_391_1196_U17, new_P2_ADD_391_1196_U18,
    new_P2_ADD_391_1196_U19, new_P2_ADD_391_1196_U20,
    new_P2_ADD_391_1196_U21, new_P2_ADD_391_1196_U22,
    new_P2_ADD_391_1196_U23, new_P2_ADD_391_1196_U24,
    new_P2_ADD_391_1196_U25, new_P2_ADD_391_1196_U26,
    new_P2_ADD_391_1196_U27, new_P2_ADD_391_1196_U28,
    new_P2_ADD_391_1196_U29, new_P2_ADD_391_1196_U30,
    new_P2_ADD_391_1196_U31, new_P2_ADD_391_1196_U32,
    new_P2_ADD_391_1196_U33, new_P2_ADD_391_1196_U34,
    new_P2_ADD_391_1196_U35, new_P2_ADD_391_1196_U36,
    new_P2_ADD_391_1196_U37, new_P2_ADD_391_1196_U38,
    new_P2_ADD_391_1196_U39, new_P2_ADD_391_1196_U40,
    new_P2_ADD_391_1196_U41, new_P2_ADD_391_1196_U42,
    new_P2_ADD_391_1196_U43, new_P2_ADD_391_1196_U44,
    new_P2_ADD_391_1196_U45, new_P2_ADD_391_1196_U46,
    new_P2_ADD_391_1196_U47, new_P2_ADD_391_1196_U48,
    new_P2_ADD_391_1196_U49, new_P2_ADD_391_1196_U50,
    new_P2_ADD_391_1196_U51, new_P2_ADD_391_1196_U52,
    new_P2_ADD_391_1196_U53, new_P2_ADD_391_1196_U54,
    new_P2_ADD_391_1196_U55, new_P2_ADD_391_1196_U56,
    new_P2_ADD_391_1196_U57, new_P2_ADD_391_1196_U58,
    new_P2_ADD_391_1196_U59, new_P2_ADD_391_1196_U60,
    new_P2_ADD_391_1196_U61, new_P2_ADD_391_1196_U62,
    new_P2_ADD_391_1196_U63, new_P2_ADD_391_1196_U64,
    new_P2_ADD_391_1196_U65, new_P2_ADD_391_1196_U66,
    new_P2_ADD_391_1196_U67, new_P2_ADD_391_1196_U68,
    new_P2_ADD_391_1196_U69, new_P2_ADD_391_1196_U70,
    new_P2_ADD_391_1196_U71, new_P2_ADD_391_1196_U72,
    new_P2_ADD_391_1196_U73, new_P2_ADD_391_1196_U74,
    new_P2_ADD_391_1196_U75, new_P2_ADD_391_1196_U76,
    new_P2_ADD_391_1196_U77, new_P2_ADD_391_1196_U78,
    new_P2_ADD_391_1196_U79, new_P2_ADD_391_1196_U80,
    new_P2_ADD_391_1196_U81, new_P2_ADD_391_1196_U82,
    new_P2_ADD_391_1196_U83, new_P2_ADD_391_1196_U84,
    new_P2_ADD_391_1196_U85, new_P2_ADD_391_1196_U86,
    new_P2_ADD_391_1196_U87, new_P2_ADD_391_1196_U88,
    new_P2_ADD_391_1196_U89, new_P2_ADD_391_1196_U90,
    new_P2_ADD_391_1196_U91, new_P2_ADD_391_1196_U92,
    new_P2_ADD_391_1196_U93, new_P2_ADD_391_1196_U94,
    new_P2_ADD_391_1196_U95, new_P2_ADD_391_1196_U96,
    new_P2_ADD_391_1196_U97, new_P2_ADD_391_1196_U98,
    new_P2_ADD_391_1196_U99, new_P2_ADD_391_1196_U100,
    new_P2_ADD_391_1196_U101, new_P2_ADD_391_1196_U102,
    new_P2_ADD_391_1196_U103, new_P2_ADD_391_1196_U104,
    new_P2_ADD_391_1196_U105, new_P2_ADD_391_1196_U106,
    new_P2_ADD_391_1196_U107, new_P2_ADD_391_1196_U108,
    new_P2_ADD_391_1196_U109, new_P2_ADD_391_1196_U110,
    new_P2_ADD_391_1196_U111, new_P2_ADD_391_1196_U112,
    new_P2_ADD_391_1196_U113, new_P2_ADD_391_1196_U114,
    new_P2_ADD_391_1196_U115, new_P2_ADD_391_1196_U116,
    new_P2_ADD_391_1196_U117, new_P2_ADD_391_1196_U118,
    new_P2_ADD_391_1196_U119, new_P2_ADD_391_1196_U120,
    new_P2_ADD_391_1196_U121, new_P2_ADD_391_1196_U122,
    new_P2_ADD_391_1196_U123, new_P2_ADD_391_1196_U124,
    new_P2_ADD_391_1196_U125, new_P2_ADD_391_1196_U126,
    new_P2_ADD_391_1196_U127, new_P2_ADD_391_1196_U128,
    new_P2_ADD_391_1196_U129, new_P2_ADD_391_1196_U130,
    new_P2_ADD_391_1196_U131, new_P2_ADD_391_1196_U132,
    new_P2_ADD_391_1196_U133, new_P2_ADD_391_1196_U134,
    new_P2_ADD_391_1196_U135, new_P2_ADD_391_1196_U136,
    new_P2_ADD_391_1196_U137, new_P2_ADD_391_1196_U138,
    new_P2_ADD_391_1196_U139, new_P2_ADD_391_1196_U140,
    new_P2_ADD_391_1196_U141, new_P2_ADD_391_1196_U142,
    new_P2_ADD_391_1196_U143, new_P2_ADD_391_1196_U144,
    new_P2_ADD_391_1196_U145, new_P2_ADD_391_1196_U146,
    new_P2_ADD_391_1196_U147, new_P2_ADD_391_1196_U148,
    new_P2_ADD_391_1196_U149, new_P2_ADD_391_1196_U150,
    new_P2_ADD_391_1196_U151, new_P2_ADD_391_1196_U152,
    new_P2_ADD_391_1196_U153, new_P2_ADD_391_1196_U154,
    new_P2_ADD_391_1196_U155, new_P2_ADD_391_1196_U156,
    new_P2_ADD_391_1196_U157, new_P2_ADD_391_1196_U158,
    new_P2_ADD_391_1196_U159, new_P2_ADD_391_1196_U160,
    new_P2_ADD_391_1196_U161, new_P2_ADD_391_1196_U162,
    new_P2_ADD_391_1196_U163, new_P2_ADD_391_1196_U164,
    new_P2_ADD_391_1196_U165, new_P2_ADD_391_1196_U166,
    new_P2_ADD_391_1196_U167, new_P2_ADD_391_1196_U168,
    new_P2_ADD_391_1196_U169, new_P2_ADD_391_1196_U170,
    new_P2_ADD_391_1196_U171, new_P2_ADD_391_1196_U172,
    new_P2_ADD_391_1196_U173, new_P2_ADD_391_1196_U174,
    new_P2_ADD_391_1196_U175, new_P2_ADD_391_1196_U176,
    new_P2_ADD_391_1196_U177, new_P2_ADD_391_1196_U178,
    new_P2_ADD_391_1196_U179, new_P2_ADD_391_1196_U180,
    new_P2_ADD_391_1196_U181, new_P2_ADD_391_1196_U182,
    new_P2_ADD_391_1196_U183, new_P2_ADD_391_1196_U184,
    new_P2_ADD_391_1196_U185, new_P2_ADD_391_1196_U186,
    new_P2_ADD_391_1196_U187, new_P2_ADD_391_1196_U188,
    new_P2_ADD_391_1196_U189, new_P2_ADD_391_1196_U190,
    new_P2_ADD_391_1196_U191, new_P2_ADD_391_1196_U192,
    new_P2_ADD_391_1196_U193, new_P2_ADD_391_1196_U194,
    new_P2_ADD_391_1196_U195, new_P2_ADD_391_1196_U196,
    new_P2_ADD_391_1196_U197, new_P2_ADD_391_1196_U198,
    new_P2_ADD_391_1196_U199, new_P2_ADD_391_1196_U200,
    new_P2_ADD_391_1196_U201, new_P2_ADD_391_1196_U202,
    new_P2_ADD_391_1196_U203, new_P2_ADD_391_1196_U204,
    new_P2_ADD_391_1196_U205, new_P2_ADD_391_1196_U206,
    new_P2_ADD_391_1196_U207, new_P2_ADD_391_1196_U208,
    new_P2_ADD_391_1196_U209, new_P2_ADD_391_1196_U210,
    new_P2_ADD_391_1196_U211, new_P2_ADD_391_1196_U212,
    new_P2_ADD_391_1196_U213, new_P2_ADD_391_1196_U214,
    new_P2_ADD_391_1196_U215, new_P2_ADD_391_1196_U216,
    new_P2_ADD_391_1196_U217, new_P2_ADD_391_1196_U218,
    new_P2_ADD_391_1196_U219, new_P2_ADD_391_1196_U220,
    new_P2_ADD_391_1196_U221, new_P2_ADD_391_1196_U222,
    new_P2_ADD_391_1196_U223, new_P2_ADD_391_1196_U224,
    new_P2_ADD_391_1196_U225, new_P2_ADD_391_1196_U226,
    new_P2_ADD_391_1196_U227, new_P2_ADD_391_1196_U228,
    new_P2_ADD_391_1196_U229, new_P2_ADD_391_1196_U230,
    new_P2_ADD_391_1196_U231, new_P2_ADD_391_1196_U232,
    new_P2_ADD_391_1196_U233, new_P2_ADD_391_1196_U234,
    new_P2_ADD_391_1196_U235, new_P2_ADD_391_1196_U236,
    new_P2_ADD_391_1196_U237, new_P2_ADD_391_1196_U238,
    new_P2_ADD_391_1196_U239, new_P2_ADD_391_1196_U240,
    new_P2_ADD_391_1196_U241, new_P2_ADD_391_1196_U242,
    new_P2_ADD_391_1196_U243, new_P2_ADD_391_1196_U244,
    new_P2_ADD_391_1196_U245, new_P2_ADD_391_1196_U246,
    new_P2_ADD_391_1196_U247, new_P2_ADD_391_1196_U248,
    new_P2_ADD_391_1196_U249, new_P2_ADD_391_1196_U250,
    new_P2_ADD_391_1196_U251, new_P2_ADD_391_1196_U252,
    new_P2_ADD_391_1196_U253, new_P2_ADD_391_1196_U254,
    new_P2_ADD_391_1196_U255, new_P2_ADD_391_1196_U256,
    new_P2_ADD_391_1196_U257, new_P2_ADD_391_1196_U258,
    new_P2_ADD_391_1196_U259, new_P2_ADD_391_1196_U260,
    new_P2_ADD_391_1196_U261, new_P2_ADD_391_1196_U262,
    new_P2_ADD_391_1196_U263, new_P2_ADD_391_1196_U264,
    new_P2_ADD_391_1196_U265, new_P2_ADD_391_1196_U266,
    new_P2_ADD_391_1196_U267, new_P2_ADD_391_1196_U268,
    new_P2_ADD_391_1196_U269, new_P2_ADD_391_1196_U270,
    new_P2_ADD_391_1196_U271, new_P2_ADD_391_1196_U272,
    new_P2_ADD_391_1196_U273, new_P2_ADD_391_1196_U274,
    new_P2_ADD_391_1196_U275, new_P2_ADD_391_1196_U276,
    new_P2_ADD_391_1196_U277, new_P2_ADD_391_1196_U278,
    new_P2_ADD_391_1196_U279, new_P2_ADD_391_1196_U280,
    new_P2_ADD_391_1196_U281, new_P2_ADD_391_1196_U282,
    new_P2_ADD_391_1196_U283, new_P2_ADD_391_1196_U284,
    new_P2_ADD_391_1196_U285, new_P2_ADD_391_1196_U286,
    new_P2_ADD_391_1196_U287, new_P2_ADD_391_1196_U288,
    new_P2_ADD_391_1196_U289, new_P2_ADD_391_1196_U290,
    new_P2_ADD_391_1196_U291, new_P2_ADD_391_1196_U292,
    new_P2_ADD_391_1196_U293, new_P2_ADD_391_1196_U294,
    new_P2_ADD_391_1196_U295, new_P2_ADD_391_1196_U296,
    new_P2_ADD_391_1196_U297, new_P2_ADD_391_1196_U298,
    new_P2_ADD_391_1196_U299, new_P2_ADD_391_1196_U300,
    new_P2_ADD_391_1196_U301, new_P2_ADD_391_1196_U302,
    new_P2_ADD_391_1196_U303, new_P2_ADD_391_1196_U304,
    new_P2_ADD_391_1196_U305, new_P2_ADD_391_1196_U306,
    new_P2_ADD_391_1196_U307, new_P2_ADD_391_1196_U308,
    new_P2_ADD_391_1196_U309, new_P2_ADD_391_1196_U310,
    new_P2_ADD_391_1196_U311, new_P2_ADD_391_1196_U312,
    new_P2_ADD_391_1196_U313, new_P2_ADD_391_1196_U314,
    new_P2_ADD_391_1196_U315, new_P2_ADD_391_1196_U316,
    new_P2_ADD_391_1196_U317, new_P2_ADD_391_1196_U318,
    new_P2_ADD_391_1196_U319, new_P2_ADD_391_1196_U320,
    new_P2_ADD_391_1196_U321, new_P2_ADD_391_1196_U322,
    new_P2_ADD_391_1196_U323, new_P2_ADD_391_1196_U324,
    new_P2_ADD_391_1196_U325, new_P2_ADD_391_1196_U326,
    new_P2_ADD_391_1196_U327, new_P2_ADD_391_1196_U328,
    new_P2_ADD_391_1196_U329, new_P2_ADD_391_1196_U330,
    new_P2_ADD_391_1196_U331, new_P2_ADD_391_1196_U332,
    new_P2_ADD_391_1196_U333, new_P2_ADD_391_1196_U334,
    new_P2_ADD_391_1196_U335, new_P2_ADD_391_1196_U336,
    new_P2_ADD_391_1196_U337, new_P2_ADD_391_1196_U338,
    new_P2_ADD_391_1196_U339, new_P2_ADD_391_1196_U340,
    new_P2_ADD_391_1196_U341, new_P2_ADD_391_1196_U342,
    new_P2_ADD_391_1196_U343, new_P2_ADD_391_1196_U344,
    new_P2_ADD_391_1196_U345, new_P2_ADD_391_1196_U346,
    new_P2_ADD_391_1196_U347, new_P2_ADD_391_1196_U348,
    new_P2_ADD_391_1196_U349, new_P2_ADD_391_1196_U350,
    new_P2_ADD_391_1196_U351, new_P2_ADD_391_1196_U352,
    new_P2_ADD_391_1196_U353, new_P2_ADD_391_1196_U354,
    new_P2_ADD_391_1196_U355, new_P2_ADD_391_1196_U356,
    new_P2_ADD_391_1196_U357, new_P2_ADD_391_1196_U358,
    new_P2_ADD_391_1196_U359, new_P2_ADD_391_1196_U360,
    new_P2_ADD_391_1196_U361, new_P2_ADD_391_1196_U362,
    new_P2_ADD_391_1196_U363, new_P2_ADD_391_1196_U364,
    new_P2_ADD_391_1196_U365, new_P2_ADD_391_1196_U366,
    new_P2_ADD_391_1196_U367, new_P2_ADD_391_1196_U368,
    new_P2_ADD_391_1196_U369, new_P2_ADD_391_1196_U370,
    new_P2_ADD_391_1196_U371, new_P2_ADD_391_1196_U372,
    new_P2_ADD_391_1196_U373, new_P2_ADD_391_1196_U374,
    new_P2_ADD_391_1196_U375, new_P2_ADD_391_1196_U376,
    new_P2_ADD_391_1196_U377, new_P2_ADD_391_1196_U378,
    new_P2_ADD_391_1196_U379, new_P2_ADD_391_1196_U380,
    new_P2_ADD_391_1196_U381, new_P2_ADD_391_1196_U382,
    new_P2_ADD_391_1196_U383, new_P2_ADD_391_1196_U384,
    new_P2_ADD_391_1196_U385, new_P2_ADD_391_1196_U386,
    new_P2_ADD_391_1196_U387, new_P2_ADD_391_1196_U388,
    new_P2_ADD_391_1196_U389, new_P2_ADD_391_1196_U390,
    new_P2_ADD_391_1196_U391, new_P2_ADD_391_1196_U392,
    new_P2_ADD_391_1196_U393, new_P2_ADD_391_1196_U394,
    new_P2_ADD_391_1196_U395, new_P2_ADD_391_1196_U396,
    new_P2_ADD_391_1196_U397, new_P2_ADD_391_1196_U398,
    new_P2_ADD_391_1196_U399, new_P2_ADD_391_1196_U400,
    new_P2_ADD_391_1196_U401, new_P2_ADD_391_1196_U402,
    new_P2_ADD_391_1196_U403, new_P2_ADD_391_1196_U404,
    new_P2_ADD_391_1196_U405, new_P2_ADD_391_1196_U406,
    new_P2_ADD_391_1196_U407, new_P2_ADD_391_1196_U408,
    new_P2_ADD_391_1196_U409, new_P2_ADD_391_1196_U410,
    new_P2_ADD_391_1196_U411, new_P2_ADD_391_1196_U412,
    new_P2_ADD_391_1196_U413, new_P2_ADD_391_1196_U414,
    new_P2_ADD_391_1196_U415, new_P2_ADD_391_1196_U416,
    new_P2_ADD_391_1196_U417, new_P2_ADD_391_1196_U418,
    new_P2_ADD_391_1196_U419, new_P2_ADD_391_1196_U420,
    new_P2_ADD_391_1196_U421, new_P2_ADD_391_1196_U422,
    new_P2_ADD_391_1196_U423, new_P2_ADD_391_1196_U424,
    new_P2_ADD_391_1196_U425, new_P2_ADD_391_1196_U426,
    new_P2_ADD_391_1196_U427, new_P2_ADD_391_1196_U428,
    new_P2_ADD_391_1196_U429, new_P2_ADD_391_1196_U430,
    new_P2_ADD_391_1196_U431, new_P2_ADD_391_1196_U432,
    new_P2_ADD_391_1196_U433, new_P2_ADD_391_1196_U434,
    new_P2_ADD_391_1196_U435, new_P2_ADD_391_1196_U436,
    new_P2_ADD_391_1196_U437, new_P2_ADD_391_1196_U438,
    new_P2_ADD_391_1196_U439, new_P2_ADD_391_1196_U440,
    new_P2_ADD_391_1196_U441, new_P2_ADD_391_1196_U442,
    new_P2_ADD_391_1196_U443, new_P2_ADD_391_1196_U444,
    new_P2_ADD_391_1196_U445, new_P2_ADD_391_1196_U446,
    new_P2_ADD_391_1196_U447, new_P2_ADD_391_1196_U448,
    new_P2_ADD_391_1196_U449, new_P2_ADD_391_1196_U450,
    new_P2_ADD_391_1196_U451, new_P2_ADD_391_1196_U452,
    new_P2_ADD_391_1196_U453, new_P2_ADD_391_1196_U454,
    new_P2_ADD_391_1196_U455, new_P2_ADD_391_1196_U456,
    new_P2_ADD_391_1196_U457, new_P2_ADD_391_1196_U458,
    new_P2_ADD_391_1196_U459, new_P2_ADD_391_1196_U460,
    new_P2_ADD_391_1196_U461, new_P2_ADD_391_1196_U462,
    new_P2_ADD_391_1196_U463, new_P2_ADD_391_1196_U464,
    new_P2_ADD_391_1196_U465, new_P2_ADD_391_1196_U466,
    new_P2_ADD_391_1196_U467, new_P2_ADD_391_1196_U468,
    new_P2_ADD_391_1196_U469, new_P2_ADD_391_1196_U470,
    new_P2_ADD_391_1196_U471, new_P2_ADD_391_1196_U472,
    new_P2_ADD_391_1196_U473, new_P2_ADD_391_1196_U474,
    new_P2_ADD_391_1196_U475, new_P2_ADD_391_1196_U476,
    new_P2_ADD_391_1196_U477, new_P2_ADD_391_1196_U478,
    new_P2_ADD_402_1132_U4, new_P2_ADD_402_1132_U5, new_P2_ADD_402_1132_U6,
    new_P2_ADD_402_1132_U7, new_P2_ADD_402_1132_U8, new_P2_ADD_402_1132_U9,
    new_P2_ADD_402_1132_U10, new_P2_ADD_402_1132_U11,
    new_P2_ADD_402_1132_U12, new_P2_ADD_402_1132_U13,
    new_P2_ADD_402_1132_U14, new_P2_ADD_402_1132_U15,
    new_P2_ADD_402_1132_U16, new_P2_ADD_402_1132_U17,
    new_P2_ADD_402_1132_U18, new_P2_ADD_402_1132_U19,
    new_P2_ADD_402_1132_U20, new_P2_ADD_402_1132_U21,
    new_P2_ADD_402_1132_U22, new_P2_ADD_402_1132_U23,
    new_P2_ADD_402_1132_U24, new_P2_ADD_402_1132_U25,
    new_P2_ADD_402_1132_U26, new_P2_ADD_402_1132_U27,
    new_P2_ADD_402_1132_U28, new_P2_ADD_402_1132_U29,
    new_P2_ADD_402_1132_U30, new_P2_ADD_402_1132_U31,
    new_P2_ADD_402_1132_U32, new_P2_ADD_402_1132_U33,
    new_P2_ADD_402_1132_U34, new_P2_ADD_402_1132_U35,
    new_P2_ADD_402_1132_U36, new_P2_ADD_402_1132_U37,
    new_P2_ADD_402_1132_U38, new_P2_ADD_402_1132_U39,
    new_P2_ADD_402_1132_U40, new_P2_ADD_402_1132_U41,
    new_P2_ADD_402_1132_U42, new_P2_ADD_402_1132_U43,
    new_P2_ADD_402_1132_U44, new_P2_ADD_402_1132_U45,
    new_P2_ADD_402_1132_U46, new_P2_ADD_402_1132_U47,
    new_P2_ADD_402_1132_U48, new_P2_ADD_402_1132_U49,
    new_P2_ADD_402_1132_U50, new_P2_SUB_563_U6, new_P2_SUB_563_U7,
    new_P2_R2182_U4, new_P2_R2182_U5, new_P2_R2182_U6, new_P2_R2182_U7,
    new_P2_R2182_U8, new_P2_R2182_U9, new_P2_R2182_U10, new_P2_R2182_U11,
    new_P2_R2182_U12, new_P2_R2182_U13, new_P2_R2182_U14, new_P2_R2182_U15,
    new_P2_R2182_U16, new_P2_R2182_U17, new_P2_R2182_U18, new_P2_R2182_U19,
    new_P2_R2182_U20, new_P2_R2182_U21, new_P2_R2182_U22, new_P2_R2182_U23,
    new_P2_R2182_U24, new_P2_R2182_U25, new_P2_R2182_U26, new_P2_R2182_U27,
    new_P2_R2182_U28, new_P2_R2182_U29, new_P2_R2182_U30, new_P2_R2182_U31,
    new_P2_R2182_U32, new_P2_R2182_U33, new_P2_R2182_U34, new_P2_R2182_U35,
    new_P2_R2182_U36, new_P2_R2182_U37, new_P2_R2182_U38, new_P2_R2182_U39,
    new_P2_R2182_U40, new_P2_R2182_U41, new_P2_R2182_U42, new_P2_R2182_U43,
    new_P2_R2182_U44, new_P2_R2182_U45, new_P2_R2182_U46, new_P2_R2182_U47,
    new_P2_R2182_U48, new_P2_R2182_U49, new_P2_R2182_U50, new_P2_R2182_U51,
    new_P2_R2182_U52, new_P2_R2182_U53, new_P2_R2182_U54, new_P2_R2182_U55,
    new_P2_R2182_U56, new_P2_R2182_U57, new_P2_R2182_U58, new_P2_R2182_U59,
    new_P2_R2182_U60, new_P2_R2182_U61, new_P2_R2182_U62, new_P2_R2182_U63,
    new_P2_R2182_U64, new_P2_R2182_U65, new_P2_R2182_U66, new_P2_R2182_U67,
    new_P2_R2182_U68, new_P2_R2182_U69, new_P2_R2182_U70, new_P2_R2182_U71,
    new_P2_R2182_U72, new_P2_R2182_U73, new_P2_R2182_U74, new_P2_R2182_U75,
    new_P2_R2182_U76, new_P2_R2182_U77, new_P2_R2182_U78, new_P2_R2182_U79,
    new_P2_R2182_U80, new_P2_R2182_U81, new_P2_R2182_U82, new_P2_R2182_U83,
    new_P2_R2182_U84, new_P2_R2182_U85, new_P2_R2182_U86, new_P2_R2182_U87,
    new_P2_R2182_U88, new_P2_R2182_U89, new_P2_R2182_U90, new_P2_R2182_U91,
    new_P2_R2182_U92, new_P2_R2182_U93, new_P2_R2182_U94, new_P2_R2182_U95,
    new_P2_R2182_U96, new_P2_R2182_U97, new_P2_R2182_U98, new_P2_R2182_U99,
    new_P2_R2182_U100, new_P2_R2182_U101, new_P2_R2182_U102,
    new_P2_R2182_U103, new_P2_R2182_U104, new_P2_R2182_U105,
    new_P2_R2182_U106, new_P2_R2182_U107, new_P2_R2182_U108,
    new_P2_R2182_U109, new_P2_R2182_U110, new_P2_R2182_U111,
    new_P2_R2182_U112, new_P2_R2182_U113, new_P2_R2182_U114,
    new_P2_R2182_U115, new_P2_R2182_U116, new_P2_R2182_U117,
    new_P2_R2182_U118, new_P2_R2182_U119, new_P2_R2182_U120,
    new_P2_R2182_U121, new_P2_R2182_U122, new_P2_R2182_U123,
    new_P2_R2182_U124, new_P2_R2182_U125, new_P2_R2182_U126,
    new_P2_R2182_U127, new_P2_R2182_U128, new_P2_R2182_U129,
    new_P2_R2182_U130, new_P2_R2182_U131, new_P2_R2182_U132,
    new_P2_R2182_U133, new_P2_R2182_U134, new_P2_R2182_U135,
    new_P2_R2182_U136, new_P2_R2182_U137, new_P2_R2182_U138,
    new_P2_R2182_U139, new_P2_R2182_U140, new_P2_R2182_U141,
    new_P2_R2182_U142, new_P2_R2182_U143, new_P2_R2182_U144,
    new_P2_R2182_U145, new_P2_R2182_U146, new_P2_R2182_U147,
    new_P2_R2182_U148, new_P2_R2182_U149, new_P2_R2182_U150,
    new_P2_R2182_U151, new_P2_R2182_U152, new_P2_R2182_U153,
    new_P2_R2182_U154, new_P2_R2182_U155, new_P2_R2182_U156,
    new_P2_R2182_U157, new_P2_R2182_U158, new_P2_R2182_U159,
    new_P2_R2182_U160, new_P2_R2182_U161, new_P2_R2182_U162,
    new_P2_R2182_U163, new_P2_R2182_U164, new_P2_R2182_U165,
    new_P2_R2182_U166, new_P2_R2182_U167, new_P2_R2182_U168,
    new_P2_R2182_U169, new_P2_R2182_U170, new_P2_R2182_U171,
    new_P2_R2182_U172, new_P2_R2182_U173, new_P2_R2182_U174,
    new_P2_R2182_U175, new_P2_R2182_U176, new_P2_R2182_U177,
    new_P2_R2182_U178, new_P2_R2182_U179, new_P2_R2182_U180,
    new_P2_R2182_U181, new_P2_R2182_U182, new_P2_R2182_U183,
    new_P2_R2182_U184, new_P2_R2182_U185, new_P2_R2182_U186,
    new_P2_R2182_U187, new_P2_R2182_U188, new_P2_R2182_U189,
    new_P2_R2182_U190, new_P2_R2182_U191, new_P2_R2182_U192,
    new_P2_R2182_U193, new_P2_R2182_U194, new_P2_R2182_U195,
    new_P2_R2182_U196, new_P2_R2182_U197, new_P2_R2182_U198,
    new_P2_R2182_U199, new_P2_R2182_U200, new_P2_R2182_U201,
    new_P2_R2182_U202, new_P2_R2182_U203, new_P2_R2182_U204,
    new_P2_R2182_U205, new_P2_R2182_U206, new_P2_R2182_U207,
    new_P2_R2182_U208, new_P2_R2182_U209, new_P2_R2182_U210,
    new_P2_R2182_U211, new_P2_R2182_U212, new_P2_R2182_U213,
    new_P2_R2182_U214, new_P2_R2182_U215, new_P2_R2182_U216,
    new_P2_R2182_U217, new_P2_R2182_U218, new_P2_R2182_U219,
    new_P2_R2182_U220, new_P2_R2182_U221, new_P2_R2182_U222,
    new_P2_R2182_U223, new_P2_R2182_U224, new_P2_R2182_U225,
    new_P2_R2182_U226, new_P2_R2182_U227, new_P2_R2182_U228,
    new_P2_R2182_U229, new_P2_R2182_U230, new_P2_R2182_U231,
    new_P2_R2182_U232, new_P2_R2182_U233, new_P2_R2182_U234,
    new_P2_R2182_U235, new_P2_R2182_U236, new_P2_R2182_U237,
    new_P2_R2182_U238, new_P2_R2182_U239, new_P2_R2182_U240,
    new_P2_R2182_U241, new_P2_R2182_U242, new_P2_R2182_U243,
    new_P2_R2182_U244, new_P2_R2182_U245, new_P2_R2182_U246,
    new_P2_R2182_U247, new_P2_R2182_U248, new_P2_R2182_U249,
    new_P2_R2182_U250, new_P2_R2182_U251, new_P2_R2182_U252,
    new_P2_R2182_U253, new_P2_R2182_U254, new_P2_R2182_U255,
    new_P2_R2182_U256, new_P2_R2182_U257, new_P2_R2182_U258,
    new_P2_R2182_U259, new_P2_R2182_U260, new_P2_R2182_U261,
    new_P2_R2182_U262, new_P2_R2182_U263, new_P2_R2182_U264,
    new_P2_R2182_U265, new_P2_R2182_U266, new_P2_R2182_U267,
    new_P2_R2182_U268, new_P2_R2182_U269, new_P2_R2182_U270,
    new_P2_R2182_U271, new_P2_R2182_U272, new_P2_R2182_U273,
    new_P2_R2182_U274, new_P2_R2182_U275, new_P2_R2182_U276,
    new_P2_R2182_U277, new_P2_R2182_U278, new_P2_R2182_U279,
    new_P2_R2182_U280, new_P2_R2182_U281, new_P2_R2182_U282,
    new_P2_R2182_U283, new_P2_R2182_U284, new_P2_R2182_U285,
    new_P2_R2182_U286, new_P2_R2182_U287, new_P2_R2182_U288,
    new_P2_R2182_U289, new_P2_R2182_U290, new_P2_R2182_U291,
    new_P2_R2182_U292, new_P2_R2182_U293, new_P2_R2182_U294,
    new_P2_R2182_U295, new_P2_R2182_U296, new_P2_R2182_U297,
    new_P2_R2182_U298, new_P2_R2182_U299, new_P2_R2182_U300,
    new_P2_R2182_U301, new_P2_R2182_U302, new_P2_R2182_U303,
    new_P2_R2182_U304, new_P2_R2182_U305, new_P2_R2167_U6, new_P2_R2167_U7,
    new_P2_R2167_U8, new_P2_R2167_U9, new_P2_R2167_U10, new_P2_R2167_U11,
    new_P2_R2167_U12, new_P2_R2167_U13, new_P2_R2167_U14, new_P2_R2167_U15,
    new_P2_R2167_U16, new_P2_R2167_U17, new_P2_R2167_U18, new_P2_R2167_U19,
    new_P2_R2167_U20, new_P2_R2167_U21, new_P2_R2167_U22, new_P2_R2167_U23,
    new_P2_R2167_U24, new_P2_R2167_U25, new_P2_R2167_U26, new_P2_R2167_U27,
    new_P2_R2167_U28, new_P2_R2167_U29, new_P2_R2167_U30, new_P2_R2167_U31,
    new_P2_R2167_U32, new_P2_R2167_U33, new_P2_R2167_U34, new_P2_R2167_U35,
    new_P2_R2167_U36, new_P2_R2167_U37, new_P2_R2167_U38, new_P2_R2167_U39,
    new_P2_R2167_U40, new_P2_R2167_U41, new_P2_R2167_U42, new_P2_R2027_U5,
    new_P2_R2027_U6, new_P2_R2027_U7, new_P2_R2027_U8, new_P2_R2027_U9,
    new_P2_R2027_U10, new_P2_R2027_U11, new_P2_R2027_U12, new_P2_R2027_U13,
    new_P2_R2027_U14, new_P2_R2027_U15, new_P2_R2027_U16, new_P2_R2027_U17,
    new_P2_R2027_U18, new_P2_R2027_U19, new_P2_R2027_U20, new_P2_R2027_U21,
    new_P2_R2027_U22, new_P2_R2027_U23, new_P2_R2027_U24, new_P2_R2027_U25,
    new_P2_R2027_U26, new_P2_R2027_U27, new_P2_R2027_U28, new_P2_R2027_U29,
    new_P2_R2027_U30, new_P2_R2027_U31, new_P2_R2027_U32, new_P2_R2027_U33,
    new_P2_R2027_U34, new_P2_R2027_U35, new_P2_R2027_U36, new_P2_R2027_U37,
    new_P2_R2027_U38, new_P2_R2027_U39, new_P2_R2027_U40, new_P2_R2027_U41,
    new_P2_R2027_U42, new_P2_R2027_U43, new_P2_R2027_U44, new_P2_R2027_U45,
    new_P2_R2027_U46, new_P2_R2027_U47, new_P2_R2027_U48, new_P2_R2027_U49,
    new_P2_R2027_U50, new_P2_R2027_U51, new_P2_R2027_U52, new_P2_R2027_U53,
    new_P2_R2027_U54, new_P2_R2027_U55, new_P2_R2027_U56, new_P2_R2027_U57,
    new_P2_R2027_U58, new_P2_R2027_U59, new_P2_R2027_U60, new_P2_R2027_U61,
    new_P2_R2027_U62, new_P2_R2027_U63, new_P2_R2027_U64, new_P2_R2027_U65,
    new_P2_R2027_U66, new_P2_R2027_U67, new_P2_R2027_U68, new_P2_R2027_U69,
    new_P2_R2027_U70, new_P2_R2027_U71, new_P2_R2027_U72, new_P2_R2027_U73,
    new_P2_R2027_U74, new_P2_R2027_U75, new_P2_R2027_U76, new_P2_R2027_U77,
    new_P2_R2027_U78, new_P2_R2027_U79, new_P2_R2027_U80, new_P2_R2027_U81,
    new_P2_R2027_U82, new_P2_R2027_U83, new_P2_R2027_U84, new_P2_R2027_U85,
    new_P2_R2027_U86, new_P2_R2027_U87, new_P2_R2027_U88, new_P2_R2027_U89,
    new_P2_R2027_U90, new_P2_R2027_U91, new_P2_R2027_U92, new_P2_R2027_U93,
    new_P2_R2027_U94, new_P2_R2027_U95, new_P2_R2027_U96, new_P2_R2027_U97,
    new_P2_R2027_U98, new_P2_R2027_U99, new_P2_R2027_U100,
    new_P2_R2027_U101, new_P2_R2027_U102, new_P2_R2027_U103,
    new_P2_R2027_U104, new_P2_R2027_U105, new_P2_R2027_U106,
    new_P2_R2027_U107, new_P2_R2027_U108, new_P2_R2027_U109,
    new_P2_R2027_U110, new_P2_R2027_U111, new_P2_R2027_U112,
    new_P2_R2027_U113, new_P2_R2027_U114, new_P2_R2027_U115,
    new_P2_R2027_U116, new_P2_R2027_U117, new_P2_R2027_U118,
    new_P2_R2027_U119, new_P2_R2027_U120, new_P2_R2027_U121,
    new_P2_R2027_U122, new_P2_R2027_U123, new_P2_R2027_U124,
    new_P2_R2027_U125, new_P2_R2027_U126, new_P2_R2027_U127,
    new_P2_R2027_U128, new_P2_R2027_U129, new_P2_R2027_U130,
    new_P2_R2027_U131, new_P2_R2027_U132, new_P2_R2027_U133,
    new_P2_R2027_U134, new_P2_R2027_U135, new_P2_R2027_U136,
    new_P2_R2027_U137, new_P2_R2027_U138, new_P2_R2027_U139,
    new_P2_R2027_U140, new_P2_R2027_U141, new_P2_R2027_U142,
    new_P2_R2027_U143, new_P2_R2027_U144, new_P2_R2027_U145,
    new_P2_R2027_U146, new_P2_R2027_U147, new_P2_R2027_U148,
    new_P2_R2027_U149, new_P2_R2027_U150, new_P2_R2027_U151,
    new_P2_R2027_U152, new_P2_R2027_U153, new_P2_R2027_U154,
    new_P2_R2027_U155, new_P2_R2027_U156, new_P2_R2027_U157,
    new_P2_R2027_U158, new_P2_R2027_U159, new_P2_R2027_U160,
    new_P2_R2027_U161, new_P2_R2027_U162, new_P2_R2027_U163,
    new_P2_R2027_U164, new_P2_R2027_U165, new_P2_R2027_U166,
    new_P2_R2027_U167, new_P2_R2027_U168, new_P2_R2027_U169,
    new_P2_R2027_U170, new_P2_R2027_U171, new_P2_R2027_U172,
    new_P2_R2027_U173, new_P2_R2027_U174, new_P2_R2027_U175,
    new_P2_R2027_U176, new_P2_R2027_U177, new_P2_R2027_U178,
    new_P2_R2027_U179, new_P2_R2027_U180, new_P2_R2027_U181,
    new_P2_R2027_U182, new_P2_R2027_U183, new_P2_R2027_U184,
    new_P2_R2027_U185, new_P2_R2027_U186, new_P2_R2027_U187,
    new_P2_R2027_U188, new_P2_R2027_U189, new_P2_LT_563_1260_U6,
    new_P2_LT_563_1260_U7, new_P2_R2337_U4, new_P2_R2337_U5,
    new_P2_R2337_U6, new_P2_R2337_U7, new_P2_R2337_U8, new_P2_R2337_U9,
    new_P2_R2337_U10, new_P2_R2337_U11, new_P2_R2337_U12, new_P2_R2337_U13,
    new_P2_R2337_U14, new_P2_R2337_U15, new_P2_R2337_U16, new_P2_R2337_U17,
    new_P2_R2337_U18, new_P2_R2337_U19, new_P2_R2337_U20, new_P2_R2337_U21,
    new_P2_R2337_U22, new_P2_R2337_U23, new_P2_R2337_U24, new_P2_R2337_U25,
    new_P2_R2337_U26, new_P2_R2337_U27, new_P2_R2337_U28, new_P2_R2337_U29,
    new_P2_R2337_U30, new_P2_R2337_U31, new_P2_R2337_U32, new_P2_R2337_U33,
    new_P2_R2337_U34, new_P2_R2337_U35, new_P2_R2337_U36, new_P2_R2337_U37,
    new_P2_R2337_U38, new_P2_R2337_U39, new_P2_R2337_U40, new_P2_R2337_U41,
    new_P2_R2337_U42, new_P2_R2337_U43, new_P2_R2337_U44, new_P2_R2337_U45,
    new_P2_R2337_U46, new_P2_R2337_U47, new_P2_R2337_U48, new_P2_R2337_U49,
    new_P2_R2337_U50, new_P2_R2337_U51, new_P2_R2337_U52, new_P2_R2337_U53,
    new_P2_R2337_U54, new_P2_R2337_U55, new_P2_R2337_U56, new_P2_R2337_U57,
    new_P2_R2337_U58, new_P2_R2337_U59, new_P2_R2337_U60, new_P2_R2337_U61,
    new_P2_R2337_U62, new_P2_R2337_U63, new_P2_R2337_U64, new_P2_R2337_U65,
    new_P2_R2337_U66, new_P2_R2337_U67, new_P2_R2337_U68, new_P2_R2337_U69,
    new_P2_R2337_U70, new_P2_R2337_U71, new_P2_R2337_U72, new_P2_R2337_U73,
    new_P2_R2337_U74, new_P2_R2337_U75, new_P2_R2337_U76, new_P2_R2337_U77,
    new_P2_R2337_U78, new_P2_R2337_U79, new_P2_R2337_U80, new_P2_R2337_U81,
    new_P2_R2337_U82, new_P2_R2337_U83, new_P2_R2337_U84, new_P2_R2337_U85,
    new_P2_R2337_U86, new_P2_R2337_U87, new_P2_R2337_U88, new_P2_R2337_U89,
    new_P2_R2337_U90, new_P2_R2337_U91, new_P2_R2337_U92, new_P2_R2337_U93,
    new_P2_R2337_U94, new_P2_R2337_U95, new_P2_R2337_U96, new_P2_R2337_U97,
    new_P2_R2337_U98, new_P2_R2337_U99, new_P2_R2337_U100,
    new_P2_R2337_U101, new_P2_R2337_U102, new_P2_R2337_U103,
    new_P2_R2337_U104, new_P2_R2337_U105, new_P2_R2337_U106,
    new_P2_R2337_U107, new_P2_R2337_U108, new_P2_R2337_U109,
    new_P2_R2337_U110, new_P2_R2337_U111, new_P2_R2337_U112,
    new_P2_R2337_U113, new_P2_R2337_U114, new_P2_R2337_U115,
    new_P2_R2337_U116, new_P2_R2337_U117, new_P2_R2337_U118,
    new_P2_R2337_U119, new_P2_R2337_U120, new_P2_R2337_U121,
    new_P2_R2337_U122, new_P2_R2337_U123, new_P2_R2337_U124,
    new_P2_R2337_U125, new_P2_R2337_U126, new_P2_R2337_U127,
    new_P2_R2337_U128, new_P2_R2337_U129, new_P2_R2337_U130,
    new_P2_R2337_U131, new_P2_R2337_U132, new_P2_R2337_U133,
    new_P2_R2337_U134, new_P2_R2337_U135, new_P2_R2337_U136,
    new_P2_R2337_U137, new_P2_R2337_U138, new_P2_R2337_U139,
    new_P2_R2337_U140, new_P2_R2337_U141, new_P2_R2337_U142,
    new_P2_R2337_U143, new_P2_R2337_U144, new_P2_R2337_U145,
    new_P2_R2337_U146, new_P2_R2337_U147, new_P2_R2337_U148,
    new_P2_R2337_U149, new_P2_R2337_U150, new_P2_R2337_U151,
    new_P2_R2337_U152, new_P2_R2337_U153, new_P2_R2337_U154,
    new_P2_R2337_U155, new_P2_R2337_U156, new_P2_R2337_U157,
    new_P2_R2337_U158, new_P2_R2337_U159, new_P2_R2337_U160,
    new_P2_R2337_U161, new_P2_R2337_U162, new_P2_R2337_U163,
    new_P2_R2337_U164, new_P2_R2337_U165, new_P2_R2337_U166,
    new_P2_R2337_U167, new_P2_R2337_U168, new_P2_R2337_U169,
    new_P2_R2337_U170, new_P2_R2337_U171, new_P2_R2337_U172,
    new_P2_R2337_U173, new_P2_R2337_U174, new_P2_R2337_U175,
    new_P2_R2337_U176, new_P2_R2337_U177, new_P2_R2337_U178,
    new_P2_R2337_U179, new_P2_R2337_U180, new_P2_R2337_U181,
    new_P2_R2337_U182, new_P2_R2147_U4, new_P2_R2147_U5, new_P2_R2147_U6,
    new_P2_R2147_U7, new_P2_R2147_U8, new_P2_R2147_U9, new_P2_R2147_U10,
    new_P2_R2147_U11, new_P2_R2147_U12, new_P2_R2147_U13, new_P2_R2147_U14,
    new_P2_R2147_U15, new_P2_R2147_U16, new_P2_R2147_U17, new_P2_R2147_U18,
    new_P2_R2147_U19, new_P2_R2147_U20, new_P2_R2219_U6, new_P2_R2219_U7,
    new_P2_R2219_U8, new_P2_R2219_U9, new_P2_R2219_U10, new_P2_R2219_U11,
    new_P2_R2219_U12, new_P2_R2219_U13, new_P2_R2219_U14, new_P2_R2219_U15,
    new_P2_R2219_U16, new_P2_R2219_U17, new_P2_R2219_U18, new_P2_R2219_U19,
    new_P2_R2219_U20, new_P2_R2219_U21, new_P2_R2219_U22, new_P2_R2219_U23,
    new_P2_R2219_U24, new_P2_R2219_U25, new_P2_R2219_U26, new_P2_R2219_U27,
    new_P2_R2219_U28, new_P2_R2219_U29, new_P2_R2219_U30, new_P2_R2219_U31,
    new_P2_R2219_U32, new_P2_R2219_U33, new_P2_R2219_U34, new_P2_R2219_U35,
    new_P2_R2219_U36, new_P2_R2219_U37, new_P2_R2219_U38, new_P2_R2219_U39,
    new_P2_R2219_U40, new_P2_R2219_U41, new_P2_R2219_U42, new_P2_R2219_U43,
    new_P2_R2219_U44, new_P2_R2219_U45, new_P2_R2219_U46, new_P2_R2219_U47,
    new_P2_R2219_U48, new_P2_R2219_U49, new_P2_R2219_U50, new_P2_R2219_U51,
    new_P2_R2219_U52, new_P2_R2219_U53, new_P2_R2219_U54, new_P2_R2219_U55,
    new_P2_R2219_U56, new_P2_R2219_U57, new_P2_R2219_U58, new_P2_R2219_U59,
    new_P2_R2219_U60, new_P2_R2219_U61, new_P2_R2219_U62, new_P2_R2219_U63,
    new_P2_R2219_U64, new_P2_R2219_U65, new_P2_R2219_U66, new_P2_R2219_U67,
    new_P2_R2219_U68, new_P2_R2219_U69, new_P2_R2219_U70, new_P2_R2219_U71,
    new_P2_R2219_U72, new_P2_R2219_U73, new_P2_R2219_U74, new_P2_R2219_U75,
    new_P2_R2219_U76, new_P2_R2219_U77, new_P2_R2219_U78, new_P2_R2219_U79,
    new_P2_R2219_U80, new_P2_R2219_U81, new_P2_R2219_U82, new_P2_R2219_U83,
    new_P2_R2219_U84, new_P2_R2219_U85, new_P2_R2219_U86, new_P2_R2219_U87,
    new_P2_R2219_U88, new_P2_R2219_U89, new_P2_R2219_U90, new_P2_R2219_U91,
    new_P2_R2219_U92, new_P2_R2219_U93, new_P2_R2219_U94, new_P2_R2219_U95,
    new_P2_R2219_U96, new_P2_R2219_U97, new_P2_R2219_U98, new_P2_R2219_U99,
    new_P2_R2219_U100, new_P2_R2219_U101, new_P2_R2219_U102,
    new_P2_R2219_U103, new_P2_R2219_U104, new_P2_R2219_U105,
    new_P2_R2219_U106, new_P2_R2219_U107, new_P2_R2219_U108,
    new_P2_R2219_U109, new_P2_R2219_U110, new_P2_R2219_U111,
    new_P2_R2219_U112, new_P2_R2219_U113, new_P2_R2219_U114,
    new_P2_R2219_U115, new_P2_R2219_U116, new_P2_R2243_U6, new_P2_R2243_U7,
    new_P2_R2243_U8, new_P2_R2243_U9, new_P2_R2243_U10, new_P2_R2243_U11,
    new_P2_SUB_589_U6, new_P2_SUB_589_U7, new_P2_SUB_589_U8,
    new_P2_SUB_589_U9, new_P2_R2096_U4, new_P2_R2096_U5, new_P2_R2096_U6,
    new_P2_R2096_U7, new_P2_R2096_U8, new_P2_R2096_U9, new_P2_R2096_U10,
    new_P2_R2096_U11, new_P2_R2096_U12, new_P2_R2096_U13, new_P2_R2096_U14,
    new_P2_R2096_U15, new_P2_R2096_U16, new_P2_R2096_U17, new_P2_R2096_U18,
    new_P2_R2096_U19, new_P2_R2096_U20, new_P2_R2096_U21, new_P2_R2096_U22,
    new_P2_R2096_U23, new_P2_R2096_U24, new_P2_R2096_U25, new_P2_R2096_U26,
    new_P2_R2096_U27, new_P2_R2096_U28, new_P2_R2096_U29, new_P2_R2096_U30,
    new_P2_R2096_U31, new_P2_R2096_U32, new_P2_R2096_U33, new_P2_R2096_U34,
    new_P2_R2096_U35, new_P2_R2096_U36, new_P2_R2096_U37, new_P2_R2096_U38,
    new_P2_R2096_U39, new_P2_R2096_U40, new_P2_R2096_U41, new_P2_R2096_U42,
    new_P2_R2096_U43, new_P2_R2096_U44, new_P2_R2096_U45, new_P2_R2096_U46,
    new_P2_R2096_U47, new_P2_R2096_U48, new_P2_R2096_U49, new_P2_R2096_U50,
    new_P2_R2096_U51, new_P2_R2096_U52, new_P2_R2096_U53, new_P2_R2096_U54,
    new_P2_R2096_U55, new_P2_R2096_U56, new_P2_R2096_U57, new_P2_R2096_U58,
    new_P2_R2096_U59, new_P2_R2096_U60, new_P2_R2096_U61, new_P2_R2096_U62,
    new_P2_R2096_U63, new_P2_R2096_U64, new_P2_R2096_U65, new_P2_R2096_U66,
    new_P2_R2096_U67, new_P2_R2096_U68, new_P2_R2096_U69, new_P2_R2096_U70,
    new_P2_R2096_U71, new_P2_R2096_U72, new_P2_R2096_U73, new_P2_R2096_U74,
    new_P2_R2096_U75, new_P2_R2096_U76, new_P2_R2096_U77, new_P2_R2096_U78,
    new_P2_R2096_U79, new_P2_R2096_U80, new_P2_R2096_U81, new_P2_R2096_U82,
    new_P2_R2096_U83, new_P2_R2096_U84, new_P2_R2096_U85, new_P2_R2096_U86,
    new_P2_R2096_U87, new_P2_R2096_U88, new_P2_R2096_U89, new_P2_R2096_U90,
    new_P2_R2096_U91, new_P2_R2096_U92, new_P2_R2096_U93, new_P2_R2096_U94,
    new_P2_R2096_U95, new_P2_R2096_U96, new_P2_R2096_U97, new_P2_R2096_U98,
    new_P2_R2096_U99, new_P2_R2096_U100, new_P2_R2096_U101,
    new_P2_R2096_U102, new_P2_R2096_U103, new_P2_R2096_U104,
    new_P2_R2096_U105, new_P2_R2096_U106, new_P2_R2096_U107,
    new_P2_R2096_U108, new_P2_R2096_U109, new_P2_R2096_U110,
    new_P2_R2096_U111, new_P2_R2096_U112, new_P2_R2096_U113,
    new_P2_R2096_U114, new_P2_R2096_U115, new_P2_R2096_U116,
    new_P2_R2096_U117, new_P2_R2096_U118, new_P2_R2096_U119,
    new_P2_R2096_U120, new_P2_R2096_U121, new_P2_R2096_U122,
    new_P2_R2096_U123, new_P2_R2096_U124, new_P2_R2096_U125,
    new_P2_R2096_U126, new_P2_R2096_U127, new_P2_R2096_U128,
    new_P2_R2096_U129, new_P2_R2096_U130, new_P2_R2096_U131,
    new_P2_R2096_U132, new_P2_R2096_U133, new_P2_R2096_U134,
    new_P2_R2096_U135, new_P2_R2096_U136, new_P2_R2096_U137,
    new_P2_R2096_U138, new_P2_R2096_U139, new_P2_R2096_U140,
    new_P2_R2096_U141, new_P2_R2096_U142, new_P2_R2096_U143,
    new_P2_R2096_U144, new_P2_R2096_U145, new_P2_R2096_U146,
    new_P2_R2096_U147, new_P2_R2096_U148, new_P2_R2096_U149,
    new_P2_R2096_U150, new_P2_R2096_U151, new_P2_R2096_U152,
    new_P2_R2096_U153, new_P2_R2096_U154, new_P2_R2096_U155,
    new_P2_R2096_U156, new_P2_R2096_U157, new_P2_R2096_U158,
    new_P2_R2096_U159, new_P2_R2096_U160, new_P2_R2096_U161,
    new_P2_R2096_U162, new_P2_R2096_U163, new_P2_R2096_U164,
    new_P2_R2096_U165, new_P2_R2096_U166, new_P2_R2096_U167,
    new_P2_R2096_U168, new_P2_R2096_U169, new_P2_R2096_U170,
    new_P2_R2096_U171, new_P2_R2096_U172, new_P2_R2096_U173,
    new_P2_R2096_U174, new_P2_R2096_U175, new_P2_R2096_U176,
    new_P2_R2096_U177, new_P2_R2096_U178, new_P2_R2096_U179,
    new_P2_R2096_U180, new_P2_R2096_U181, new_P2_R2096_U182,
    new_P2_R2096_U183, new_P2_R2096_U184, new_P2_R2096_U185,
    new_P2_R2096_U186, new_P2_R2096_U187, new_P2_R2096_U188,
    new_P2_R2096_U189, new_P2_R2096_U190, new_P2_R2096_U191,
    new_P2_R2096_U192, new_P2_R2096_U193, new_P2_R2096_U194,
    new_P2_R2096_U195, new_P2_R2096_U196, new_P2_R2096_U197,
    new_P2_R2096_U198, new_P2_R2096_U199, new_P2_R2096_U200,
    new_P2_R2096_U201, new_P2_R2096_U202, new_P2_R2096_U203,
    new_P2_R2096_U204, new_P2_R2096_U205, new_P2_R2096_U206,
    new_P2_R2096_U207, new_P2_R2096_U208, new_P2_R2096_U209,
    new_P2_R2096_U210, new_P2_R2096_U211, new_P2_R2096_U212,
    new_P2_R2096_U213, new_P2_R2096_U214, new_P2_R2096_U215,
    new_P2_R2096_U216, new_P2_R2096_U217, new_P2_R2096_U218,
    new_P2_R2096_U219, new_P2_R2096_U220, new_P2_R2096_U221,
    new_P2_R2096_U222, new_P2_R2096_U223, new_P2_R2096_U224,
    new_P2_R2096_U225, new_P2_R2096_U226, new_P2_R2096_U227,
    new_P2_R2096_U228, new_P2_R2096_U229, new_P2_R2096_U230,
    new_P2_R2096_U231, new_P2_R2096_U232, new_P2_R2096_U233,
    new_P2_R2096_U234, new_P2_R2096_U235, new_P2_R2096_U236,
    new_P2_R2096_U237, new_P2_R2096_U238, new_P2_R2096_U239,
    new_P2_R2096_U240, new_P2_R2096_U241, new_P2_R2096_U242,
    new_P2_R2096_U243, new_P2_R2096_U244, new_P2_R2096_U245,
    new_P2_R2096_U246, new_P2_R2096_U247, new_P2_R2096_U248,
    new_P2_R2096_U249, new_P2_R2096_U250, new_P2_R2096_U251,
    new_P2_R2096_U252, new_P2_R2096_U253, new_P2_R2096_U254,
    new_P2_R2096_U255, new_P2_R2096_U256, new_P2_R2096_U257,
    new_P2_R2096_U258, new_P2_R2096_U259, new_P2_R2096_U260,
    new_P2_R2096_U261, new_P2_R2096_U262, new_P2_R2096_U263,
    new_P2_R2096_U264, new_P2_R2096_U265, new_P2_GTE_370_U6,
    new_P2_GTE_370_U7, new_P2_GTE_370_U8, new_P2_GTE_370_U9,
    new_P2_LT_563_U6, new_P2_LT_563_U7, new_P2_LT_563_U8, new_P2_LT_563_U9,
    new_P2_LT_563_U10, new_P2_LT_563_U11, new_P2_LT_563_U12,
    new_P2_LT_563_U13, new_P2_LT_563_U14, new_P2_LT_563_U15,
    new_P2_LT_563_U16, new_P2_LT_563_U17, new_P2_LT_563_U18,
    new_P2_LT_563_U19, new_P2_LT_563_U20, new_P2_LT_563_U21,
    new_P2_LT_563_U22, new_P2_LT_563_U23, new_P2_LT_563_U24,
    new_P2_LT_563_U25, new_P2_LT_563_U26, new_P2_LT_563_U27,
    new_P2_R2256_U4, new_P2_R2256_U5, new_P2_R2256_U6, new_P2_R2256_U7,
    new_P2_R2256_U8, new_P2_R2256_U9, new_P2_R2256_U10, new_P2_R2256_U11,
    new_P2_R2256_U12, new_P2_R2256_U13, new_P2_R2256_U14, new_P2_R2256_U15,
    new_P2_R2256_U16, new_P2_R2256_U17, new_P2_R2256_U18, new_P2_R2256_U19,
    new_P2_R2256_U20, new_P2_R2256_U21, new_P2_R2256_U22, new_P2_R2256_U23,
    new_P2_R2256_U24, new_P2_R2256_U25, new_P2_R2256_U26, new_P2_R2256_U27,
    new_P2_R2256_U28, new_P2_R2256_U29, new_P2_R2256_U30, new_P2_R2256_U31,
    new_P2_R2256_U32, new_P2_R2256_U33, new_P2_R2256_U34, new_P2_R2256_U35,
    new_P2_R2256_U36, new_P2_R2256_U37, new_P2_R2256_U38, new_P2_R2256_U39,
    new_P2_R2256_U40, new_P2_R2256_U41, new_P2_R2256_U42, new_P2_R2256_U43,
    new_P2_R2256_U44, new_P2_R2256_U45, new_P2_R2256_U46, new_P2_R2256_U47,
    new_P2_R2256_U48, new_P2_R2256_U49, new_P2_R2256_U50, new_P2_R2256_U51,
    new_P2_R2256_U52, new_P2_R2256_U53, new_P2_R2256_U54, new_P2_R2256_U55,
    new_P2_R2256_U56, new_P2_R2256_U57, new_P2_R2256_U58, new_P2_R2256_U59,
    new_P2_R2256_U60, new_P2_R2256_U61, new_P2_R2256_U62, new_P2_R2256_U63,
    new_P2_R2256_U64, new_P2_R2256_U65, new_P2_R2256_U66, new_P2_R2256_U67,
    new_P2_R2256_U68, new_P2_R2256_U69, new_P2_R2256_U70, new_P2_R2238_U6,
    new_P2_R2238_U7, new_P2_R2238_U8, new_P2_R2238_U9, new_P2_R2238_U10,
    new_P2_R2238_U11, new_P2_R2238_U12, new_P2_R2238_U13, new_P2_R2238_U14,
    new_P2_R2238_U15, new_P2_R2238_U16, new_P2_R2238_U17, new_P2_R2238_U18,
    new_P2_R2238_U19, new_P2_R2238_U20, new_P2_R2238_U21, new_P2_R2238_U22,
    new_P2_R2238_U23, new_P2_R2238_U24, new_P2_R2238_U25, new_P2_R2238_U26,
    new_P2_R2238_U27, new_P2_R2238_U28, new_P2_R2238_U29, new_P2_R2238_U30,
    new_P2_R2238_U31, new_P2_R2238_U32, new_P2_R2238_U33, new_P2_R2238_U34,
    new_P2_R2238_U35, new_P2_R2238_U36, new_P2_R2238_U37, new_P2_R2238_U38,
    new_P2_R2238_U39, new_P2_R2238_U40, new_P2_R2238_U41, new_P2_R2238_U42,
    new_P2_R2238_U43, new_P2_R2238_U44, new_P2_R2238_U45, new_P2_R2238_U46,
    new_P2_R2238_U47, new_P2_R2238_U48, new_P2_R2238_U49, new_P2_R2238_U50,
    new_P2_R2238_U51, new_P2_R2238_U52, new_P2_R2238_U53, new_P2_R2238_U54,
    new_P2_R2238_U55, new_P2_R2238_U56, new_P2_R2238_U57, new_P2_R2238_U58,
    new_P2_R2238_U59, new_P2_R2238_U60, new_P2_R2238_U61, new_P2_R2238_U62,
    new_P2_R2238_U63, new_P2_R2238_U64, new_P2_R2238_U65, new_P2_R2238_U66,
    new_P2_R1957_U6, new_P2_R1957_U7, new_P2_R1957_U8, new_P2_R1957_U9,
    new_P2_R1957_U10, new_P2_R1957_U11, new_P2_R1957_U12, new_P2_R1957_U13,
    new_P2_R1957_U14, new_P2_R1957_U15, new_P2_R1957_U16, new_P2_R1957_U17,
    new_P2_R1957_U18, new_P2_R1957_U19, new_P2_R1957_U20, new_P2_R1957_U21,
    new_P2_R1957_U22, new_P2_R1957_U23, new_P2_R1957_U24, new_P2_R1957_U25,
    new_P2_R1957_U26, new_P2_R1957_U27, new_P2_R1957_U28, new_P2_R1957_U29,
    new_P2_R1957_U30, new_P2_R1957_U31, new_P2_R1957_U32, new_P2_R1957_U33,
    new_P2_R1957_U34, new_P2_R1957_U35, new_P2_R1957_U36, new_P2_R1957_U37,
    new_P2_R1957_U38, new_P2_R1957_U39, new_P2_R1957_U40, new_P2_R1957_U41,
    new_P2_R1957_U42, new_P2_R1957_U43, new_P2_R1957_U44, new_P2_R1957_U45,
    new_P2_R1957_U46, new_P2_R1957_U47, new_P2_R1957_U48, new_P2_R1957_U49,
    new_P2_R1957_U50, new_P2_R1957_U51, new_P2_R1957_U52, new_P2_R1957_U53,
    new_P2_R1957_U54, new_P2_R1957_U55, new_P2_R1957_U56, new_P2_R1957_U57,
    new_P2_R1957_U58, new_P2_R1957_U59, new_P2_R1957_U60, new_P2_R1957_U61,
    new_P2_R1957_U62, new_P2_R1957_U63, new_P2_R1957_U64, new_P2_R1957_U65,
    new_P2_R1957_U66, new_P2_R1957_U67, new_P2_R1957_U68, new_P2_R1957_U69,
    new_P2_R1957_U70, new_P2_R1957_U71, new_P2_R1957_U72, new_P2_R1957_U73,
    new_P2_R1957_U74, new_P2_R1957_U75, new_P2_R1957_U76, new_P2_R1957_U77,
    new_P2_R1957_U78, new_P2_R1957_U79, new_P2_R1957_U80, new_P2_R1957_U81,
    new_P2_R1957_U82, new_P2_R1957_U83, new_P2_R1957_U84, new_P2_R1957_U85,
    new_P2_R1957_U86, new_P2_R1957_U87, new_P2_R1957_U88, new_P2_R1957_U89,
    new_P2_R1957_U90, new_P2_R1957_U91, new_P2_R1957_U92, new_P2_R1957_U93,
    new_P2_R1957_U94, new_P2_R1957_U95, new_P2_R1957_U96, new_P2_R1957_U97,
    new_P2_R1957_U98, new_P2_R1957_U99, new_P2_R1957_U100,
    new_P2_R1957_U101, new_P2_R1957_U102, new_P2_R1957_U103,
    new_P2_R1957_U104, new_P2_R1957_U105, new_P2_R1957_U106,
    new_P2_R1957_U107, new_P2_R1957_U108, new_P2_R1957_U109,
    new_P2_R1957_U110, new_P2_R1957_U111, new_P2_R1957_U112,
    new_P2_R1957_U113, new_P2_R1957_U114, new_P2_R1957_U115,
    new_P2_R1957_U116, new_P2_R1957_U117, new_P2_R1957_U118,
    new_P2_R1957_U119, new_P2_R1957_U120, new_P2_R1957_U121,
    new_P2_R1957_U122, new_P2_R1957_U123, new_P2_R1957_U124,
    new_P2_R1957_U125, new_P2_R1957_U126, new_P2_R1957_U127,
    new_P2_R1957_U128, new_P2_R1957_U129, new_P2_R1957_U130,
    new_P2_R1957_U131, new_P2_R1957_U132, new_P2_R1957_U133,
    new_P2_R1957_U134, new_P2_R1957_U135, new_P2_R1957_U136,
    new_P2_R1957_U137, new_P2_R1957_U138, new_P2_R1957_U139,
    new_P2_R1957_U140, new_P2_R1957_U141, new_P2_R1957_U142,
    new_P2_R1957_U143, new_P2_R1957_U144, new_P2_R1957_U145,
    new_P2_R1957_U146, new_P2_R1957_U147, new_P2_R1957_U148,
    new_P2_R1957_U149, new_P2_R1957_U150, new_P2_R1957_U151,
    new_P2_R1957_U152, new_P2_R1957_U153, new_P2_R1957_U154,
    new_P2_R1957_U155, new_P2_R1957_U156, new_P2_R1957_U157,
    new_P2_R1957_U158, new_P2_R1957_U159, new_P2_R2278_U4, new_P2_R2278_U5,
    new_P2_R2278_U6, new_P2_R2278_U7, new_P2_R2278_U8, new_P2_R2278_U9,
    new_P2_R2278_U10, new_P2_R2278_U11, new_P2_R2278_U12, new_P2_R2278_U13,
    new_P2_R2278_U14, new_P2_R2278_U15, new_P2_R2278_U16, new_P2_R2278_U17,
    new_P2_R2278_U18, new_P2_R2278_U19, new_P2_R2278_U20, new_P2_R2278_U21,
    new_P2_R2278_U22, new_P2_R2278_U23, new_P2_R2278_U24, new_P2_R2278_U25,
    new_P2_R2278_U26, new_P2_R2278_U27, new_P2_R2278_U28, new_P2_R2278_U29,
    new_P2_R2278_U30, new_P2_R2278_U31, new_P2_R2278_U32, new_P2_R2278_U33,
    new_P2_R2278_U34, new_P2_R2278_U35, new_P2_R2278_U36, new_P2_R2278_U37,
    new_P2_R2278_U38, new_P2_R2278_U39, new_P2_R2278_U40, new_P2_R2278_U41,
    new_P2_R2278_U42, new_P2_R2278_U43, new_P2_R2278_U44, new_P2_R2278_U45,
    new_P2_R2278_U46, new_P2_R2278_U47, new_P2_R2278_U48, new_P2_R2278_U49,
    new_P2_R2278_U50, new_P2_R2278_U51, new_P2_R2278_U52, new_P2_R2278_U53,
    new_P2_R2278_U54, new_P2_R2278_U55, new_P2_R2278_U56, new_P2_R2278_U57,
    new_P2_R2278_U58, new_P2_R2278_U59, new_P2_R2278_U60, new_P2_R2278_U61,
    new_P2_R2278_U62, new_P2_R2278_U63, new_P2_R2278_U64, new_P2_R2278_U65,
    new_P2_R2278_U66, new_P2_R2278_U67, new_P2_R2278_U68, new_P2_R2278_U69,
    new_P2_R2278_U70, new_P2_R2278_U71, new_P2_R2278_U72, new_P2_R2278_U73,
    new_P2_R2278_U74, new_P2_R2278_U75, new_P2_R2278_U76, new_P2_R2278_U77,
    new_P2_R2278_U78, new_P2_R2278_U79, new_P2_R2278_U80, new_P2_R2278_U81,
    new_P2_R2278_U82, new_P2_R2278_U83, new_P2_R2278_U84, new_P2_R2278_U85,
    new_P2_R2278_U86, new_P2_R2278_U87, new_P2_R2278_U88, new_P2_R2278_U89,
    new_P2_R2278_U90, new_P2_R2278_U91, new_P2_R2278_U92, new_P2_R2278_U93,
    new_P2_R2278_U94, new_P2_R2278_U95, new_P2_R2278_U96, new_P2_R2278_U97,
    new_P2_R2278_U98, new_P2_R2278_U99, new_P2_R2278_U100,
    new_P2_R2278_U101, new_P2_R2278_U102, new_P2_R2278_U103,
    new_P2_R2278_U104, new_P2_R2278_U105, new_P2_R2278_U106,
    new_P2_R2278_U107, new_P2_R2278_U108, new_P2_R2278_U109,
    new_P2_R2278_U110, new_P2_R2278_U111, new_P2_R2278_U112,
    new_P2_R2278_U113, new_P2_R2278_U114, new_P2_R2278_U115,
    new_P2_R2278_U116, new_P2_R2278_U117, new_P2_R2278_U118,
    new_P2_R2278_U119, new_P2_R2278_U120, new_P2_R2278_U121,
    new_P2_R2278_U122, new_P2_R2278_U123, new_P2_R2278_U124,
    new_P2_R2278_U125, new_P2_R2278_U126, new_P2_R2278_U127,
    new_P2_R2278_U128, new_P2_R2278_U129, new_P2_R2278_U130,
    new_P2_R2278_U131, new_P2_R2278_U132, new_P2_R2278_U133,
    new_P2_R2278_U134, new_P2_R2278_U135, new_P2_R2278_U136,
    new_P2_R2278_U137, new_P2_R2278_U138, new_P2_R2278_U139,
    new_P2_R2278_U140, new_P2_R2278_U141, new_P2_R2278_U142,
    new_P2_R2278_U143, new_P2_R2278_U144, new_P2_R2278_U145,
    new_P2_R2278_U146, new_P2_R2278_U147, new_P2_R2278_U148,
    new_P2_R2278_U149, new_P2_R2278_U150, new_P2_R2278_U151,
    new_P2_R2278_U152, new_P2_R2278_U153, new_P2_R2278_U154,
    new_P2_R2278_U155, new_P2_R2278_U156, new_P2_R2278_U157,
    new_P2_R2278_U158, new_P2_R2278_U159, new_P2_R2278_U160,
    new_P2_R2278_U161, new_P2_R2278_U162, new_P2_R2278_U163,
    new_P2_R2278_U164, new_P2_R2278_U165, new_P2_R2278_U166,
    new_P2_R2278_U167, new_P2_R2278_U168, new_P2_R2278_U169,
    new_P2_R2278_U170, new_P2_R2278_U171, new_P2_R2278_U172,
    new_P2_R2278_U173, new_P2_R2278_U174, new_P2_R2278_U175,
    new_P2_R2278_U176, new_P2_R2278_U177, new_P2_R2278_U178,
    new_P2_R2278_U179, new_P2_R2278_U180, new_P2_R2278_U181,
    new_P2_R2278_U182, new_P2_R2278_U183, new_P2_R2278_U184,
    new_P2_R2278_U185, new_P2_R2278_U186, new_P2_R2278_U187,
    new_P2_R2278_U188, new_P2_R2278_U189, new_P2_R2278_U190,
    new_P2_R2278_U191, new_P2_R2278_U192, new_P2_R2278_U193,
    new_P2_R2278_U194, new_P2_R2278_U195, new_P2_R2278_U196,
    new_P2_R2278_U197, new_P2_R2278_U198, new_P2_R2278_U199,
    new_P2_R2278_U200, new_P2_R2278_U201, new_P2_R2278_U202,
    new_P2_R2278_U203, new_P2_R2278_U204, new_P2_R2278_U205,
    new_P2_R2278_U206, new_P2_R2278_U207, new_P2_R2278_U208,
    new_P2_R2278_U209, new_P2_R2278_U210, new_P2_R2278_U211,
    new_P2_R2278_U212, new_P2_R2278_U213, new_P2_R2278_U214,
    new_P2_R2278_U215, new_P2_R2278_U216, new_P2_R2278_U217,
    new_P2_R2278_U218, new_P2_R2278_U219, new_P2_R2278_U220,
    new_P2_R2278_U221, new_P2_R2278_U222, new_P2_R2278_U223,
    new_P2_R2278_U224, new_P2_R2278_U225, new_P2_R2278_U226,
    new_P2_R2278_U227, new_P2_R2278_U228, new_P2_R2278_U229,
    new_P2_R2278_U230, new_P2_R2278_U231, new_P2_R2278_U232,
    new_P2_R2278_U233, new_P2_R2278_U234, new_P2_R2278_U235,
    new_P2_R2278_U236, new_P2_R2278_U237, new_P2_R2278_U238,
    new_P2_R2278_U239, new_P2_R2278_U240, new_P2_R2278_U241,
    new_P2_R2278_U242, new_P2_R2278_U243, new_P2_R2278_U244,
    new_P2_R2278_U245, new_P2_R2278_U246, new_P2_R2278_U247,
    new_P2_R2278_U248, new_P2_R2278_U249, new_P2_R2278_U250,
    new_P2_R2278_U251, new_P2_R2278_U252, new_P2_R2278_U253,
    new_P2_R2278_U254, new_P2_R2278_U255, new_P2_R2278_U256,
    new_P2_R2278_U257, new_P2_R2278_U258, new_P2_R2278_U259,
    new_P2_R2278_U260, new_P2_R2278_U261, new_P2_R2278_U262,
    new_P2_R2278_U263, new_P2_R2278_U264, new_P2_R2278_U265,
    new_P2_R2278_U266, new_P2_R2278_U267, new_P2_R2278_U268,
    new_P2_R2278_U269, new_P2_R2278_U270, new_P2_R2278_U271,
    new_P2_R2278_U272, new_P2_R2278_U273, new_P2_R2278_U274,
    new_P2_R2278_U275, new_P2_R2278_U276, new_P2_R2278_U277,
    new_P2_R2278_U278, new_P2_R2278_U279, new_P2_R2278_U280,
    new_P2_R2278_U281, new_P2_R2278_U282, new_P2_R2278_U283,
    new_P2_R2278_U284, new_P2_R2278_U285, new_P2_R2278_U286,
    new_P2_R2278_U287, new_P2_R2278_U288, new_P2_R2278_U289,
    new_P2_R2278_U290, new_P2_R2278_U291, new_P2_R2278_U292,
    new_P2_R2278_U293, new_P2_R2278_U294, new_P2_R2278_U295,
    new_P2_R2278_U296, new_P2_R2278_U297, new_P2_R2278_U298,
    new_P2_R2278_U299, new_P2_R2278_U300, new_P2_R2278_U301,
    new_P2_R2278_U302, new_P2_R2278_U303, new_P2_R2278_U304,
    new_P2_R2278_U305, new_P2_R2278_U306, new_P2_R2278_U307,
    new_P2_R2278_U308, new_P2_R2278_U309, new_P2_R2278_U310,
    new_P2_R2278_U311, new_P2_R2278_U312, new_P2_R2278_U313,
    new_P2_R2278_U314, new_P2_R2278_U315, new_P2_R2278_U316,
    new_P2_R2278_U317, new_P2_R2278_U318, new_P2_R2278_U319,
    new_P2_R2278_U320, new_P2_R2278_U321, new_P2_R2278_U322,
    new_P2_R2278_U323, new_P2_R2278_U324, new_P2_R2278_U325,
    new_P2_R2278_U326, new_P2_R2278_U327, new_P2_R2278_U328,
    new_P2_R2278_U329, new_P2_R2278_U330, new_P2_R2278_U331,
    new_P2_R2278_U332, new_P2_R2278_U333, new_P2_R2278_U334,
    new_P2_R2278_U335, new_P2_R2278_U336, new_P2_R2278_U337,
    new_P2_R2278_U338, new_P2_R2278_U339, new_P2_R2278_U340,
    new_P2_R2278_U341, new_P2_R2278_U342, new_P2_R2278_U343,
    new_P2_R2278_U344, new_P2_R2278_U345, new_P2_R2278_U346,
    new_P2_R2278_U347, new_P2_R2278_U348, new_P2_R2278_U349,
    new_P2_R2278_U350, new_P2_R2278_U351, new_P2_R2278_U352,
    new_P2_R2278_U353, new_P2_R2278_U354, new_P2_R2278_U355,
    new_P2_R2278_U356, new_P2_R2278_U357, new_P2_R2278_U358,
    new_P2_R2278_U359, new_P2_R2278_U360, new_P2_R2278_U361,
    new_P2_R2278_U362, new_P2_R2278_U363, new_P2_R2278_U364,
    new_P2_R2278_U365, new_P2_R2278_U366, new_P2_R2278_U367,
    new_P2_R2278_U368, new_P2_R2278_U369, new_P2_R2278_U370,
    new_P2_R2278_U371, new_P2_R2278_U372, new_P2_R2278_U373,
    new_P2_R2278_U374, new_P2_R2278_U375, new_P2_R2278_U376,
    new_P2_R2278_U377, new_P2_R2278_U378, new_P2_R2278_U379,
    new_P2_R2278_U380, new_P2_R2278_U381, new_P2_R2278_U382,
    new_P2_R2278_U383, new_P2_R2278_U384, new_P2_R2278_U385,
    new_P2_R2278_U386, new_P2_R2278_U387, new_P2_R2278_U388,
    new_P2_R2278_U389, new_P2_R2278_U390, new_P2_R2278_U391,
    new_P2_R2278_U392, new_P2_R2278_U393, new_P2_R2278_U394,
    new_P2_R2278_U395, new_P2_R2278_U396, new_P2_R2278_U397,
    new_P2_R2278_U398, new_P2_R2278_U399, new_P2_R2278_U400,
    new_P2_R2278_U401, new_P2_R2278_U402, new_P2_R2278_U403,
    new_P2_R2278_U404, new_P2_R2278_U405, new_P2_R2278_U406,
    new_P2_R2278_U407, new_P2_R2278_U408, new_P2_R2278_U409,
    new_P2_R2278_U410, new_P2_R2278_U411, new_P2_R2278_U412,
    new_P2_R2278_U413, new_P2_R2278_U414, new_P2_R2278_U415,
    new_P2_R2278_U416, new_P2_R2278_U417, new_P2_R2278_U418,
    new_P2_R2278_U419, new_P2_R2278_U420, new_P2_R2278_U421,
    new_P2_R2278_U422, new_P2_R2278_U423, new_P2_R2278_U424,
    new_P2_R2278_U425, new_P2_R2278_U426, new_P2_R2278_U427,
    new_P2_R2278_U428, new_P2_R2278_U429, new_P2_R2278_U430,
    new_P2_R2278_U431, new_P2_R2278_U432, new_P2_R2278_U433,
    new_P2_R2278_U434, new_P2_R2278_U435, new_P2_R2278_U436,
    new_P2_R2278_U437, new_P2_R2278_U438, new_P2_R2278_U439,
    new_P2_R2278_U440, new_P2_R2278_U441, new_P2_R2278_U442,
    new_P2_R2278_U443, new_P2_R2278_U444, new_P2_R2278_U445,
    new_P2_R2278_U446, new_P2_R2278_U447, new_P2_R2278_U448,
    new_P2_R2278_U449, new_P2_R2278_U450, new_P2_R2278_U451,
    new_P2_R2278_U452, new_P2_R2278_U453, new_P2_R2278_U454,
    new_P2_R2278_U455, new_P2_R2278_U456, new_P2_R2278_U457,
    new_P2_R2278_U458, new_P2_R2278_U459, new_P2_R2278_U460,
    new_P2_R2278_U461, new_P2_R2278_U462, new_P2_R2278_U463,
    new_P2_R2278_U464, new_P2_R2278_U465, new_P2_R2278_U466,
    new_P2_R2278_U467, new_P2_R2278_U468, new_P2_R2278_U469,
    new_P2_R2278_U470, new_P2_R2278_U471, new_P2_R2278_U472,
    new_P2_R2278_U473, new_P2_R2278_U474, new_P2_R2278_U475,
    new_P2_R2278_U476, new_P2_R2278_U477, new_P2_R2278_U478,
    new_P2_R2278_U479, new_P2_R2278_U480, new_P2_R2278_U481,
    new_P2_R2278_U482, new_P2_R2278_U483, new_P2_R2278_U484,
    new_P2_R2278_U485, new_P2_R2278_U486, new_P2_R2278_U487,
    new_P2_R2278_U488, new_P2_R2278_U489, new_P2_R2278_U490,
    new_P2_R2278_U491, new_P2_R2278_U492, new_P2_R2278_U493,
    new_P2_R2278_U494, new_P2_R2278_U495, new_P2_R2278_U496,
    new_P2_R2278_U497, new_P2_R2278_U498, new_P2_R2278_U499,
    new_P2_R2278_U500, new_P2_R2278_U501, new_P2_R2278_U502,
    new_P2_R2278_U503, new_P2_R2278_U504, new_P2_R2278_U505,
    new_P2_R2278_U506, new_P2_R2278_U507, new_P2_R2278_U508,
    new_P2_R2278_U509, new_P2_R2278_U510, new_P2_R2278_U511,
    new_P2_R2278_U512, new_P2_R2278_U513, new_P2_R2278_U514,
    new_P2_R2278_U515, new_P2_R2278_U516, new_P2_R2278_U517,
    new_P2_R2278_U518, new_P2_R2278_U519, new_P2_R2278_U520,
    new_P2_R2278_U521, new_P2_R2278_U522, new_P2_R2278_U523,
    new_P2_R2278_U524, new_P2_R2278_U525, new_P2_R2278_U526,
    new_P2_R2278_U527, new_P2_R2278_U528, new_P2_R2278_U529,
    new_P2_R2278_U530, new_P2_R2278_U531, new_P2_R2278_U532,
    new_P2_R2278_U533, new_P2_R2278_U534, new_P2_R2278_U535,
    new_P2_R2278_U536, new_P2_R2278_U537, new_P2_R2278_U538,
    new_P2_R2278_U539, new_P2_R2278_U540, new_P2_R2278_U541,
    new_P2_R2278_U542, new_P2_R2278_U543, new_P2_R2278_U544,
    new_P2_R2278_U545, new_P2_R2278_U546, new_P2_R2278_U547,
    new_P2_R2278_U548, new_P2_R2278_U549, new_P2_R2278_U550,
    new_P2_R2278_U551, new_P2_R2278_U552, new_P2_R2278_U553,
    new_P2_R2278_U554, new_P2_R2278_U555, new_P2_R2278_U556,
    new_P2_R2278_U557, new_P2_R2278_U558, new_P2_R2278_U559,
    new_P2_R2278_U560, new_P2_R2278_U561, new_P2_R2278_U562,
    new_P2_SUB_450_U6, new_P2_SUB_450_U7, new_P2_SUB_450_U8,
    new_P2_SUB_450_U9, new_P2_SUB_450_U10, new_P2_SUB_450_U11,
    new_P2_SUB_450_U12, new_P2_SUB_450_U13, new_P2_SUB_450_U14,
    new_P2_SUB_450_U15, new_P2_SUB_450_U16, new_P2_SUB_450_U17,
    new_P2_SUB_450_U18, new_P2_SUB_450_U19, new_P2_SUB_450_U20,
    new_P2_SUB_450_U21, new_P2_SUB_450_U22, new_P2_SUB_450_U23,
    new_P2_SUB_450_U24, new_P2_SUB_450_U25, new_P2_SUB_450_U26,
    new_P2_SUB_450_U27, new_P2_SUB_450_U28, new_P2_SUB_450_U29,
    new_P2_SUB_450_U30, new_P2_SUB_450_U31, new_P2_SUB_450_U32,
    new_P2_SUB_450_U33, new_P2_SUB_450_U34, new_P2_SUB_450_U35,
    new_P2_SUB_450_U36, new_P2_SUB_450_U37, new_P2_SUB_450_U38,
    new_P2_SUB_450_U39, new_P2_SUB_450_U40, new_P2_SUB_450_U41,
    new_P2_SUB_450_U42, new_P2_SUB_450_U43, new_P2_SUB_450_U44,
    new_P2_SUB_450_U45, new_P2_SUB_450_U46, new_P2_SUB_450_U47,
    new_P2_SUB_450_U48, new_P2_SUB_450_U49, new_P2_SUB_450_U50,
    new_P2_SUB_450_U51, new_P2_SUB_450_U52, new_P2_SUB_450_U53,
    new_P2_SUB_450_U54, new_P2_SUB_450_U55, new_P2_SUB_450_U56,
    new_P2_SUB_450_U57, new_P2_SUB_450_U58, new_P2_SUB_450_U59,
    new_P2_SUB_450_U60, new_P2_SUB_450_U61, new_P2_SUB_450_U62,
    new_P2_SUB_450_U63, new_P2_R2088_U6, new_P2_R2088_U7,
    new_P2_ADD_394_U4, new_P2_ADD_394_U5, new_P2_ADD_394_U6,
    new_P2_ADD_394_U7, new_P2_ADD_394_U8, new_P2_ADD_394_U9,
    new_P2_ADD_394_U10, new_P2_ADD_394_U11, new_P2_ADD_394_U12,
    new_P2_ADD_394_U13, new_P2_ADD_394_U14, new_P2_ADD_394_U15,
    new_P2_ADD_394_U16, new_P2_ADD_394_U17, new_P2_ADD_394_U18,
    new_P2_ADD_394_U19, new_P2_ADD_394_U20, new_P2_ADD_394_U21,
    new_P2_ADD_394_U22, new_P2_ADD_394_U23, new_P2_ADD_394_U24,
    new_P2_ADD_394_U25, new_P2_ADD_394_U26, new_P2_ADD_394_U27,
    new_P2_ADD_394_U28, new_P2_ADD_394_U29, new_P2_ADD_394_U30,
    new_P2_ADD_394_U31, new_P2_ADD_394_U32, new_P2_ADD_394_U33,
    new_P2_ADD_394_U34, new_P2_ADD_394_U35, new_P2_ADD_394_U36,
    new_P2_ADD_394_U37, new_P2_ADD_394_U38, new_P2_ADD_394_U39,
    new_P2_ADD_394_U40, new_P2_ADD_394_U41, new_P2_ADD_394_U42,
    new_P2_ADD_394_U43, new_P2_ADD_394_U44, new_P2_ADD_394_U45,
    new_P2_ADD_394_U46, new_P2_ADD_394_U47, new_P2_ADD_394_U48,
    new_P2_ADD_394_U49, new_P2_ADD_394_U50, new_P2_ADD_394_U51,
    new_P2_ADD_394_U52, new_P2_ADD_394_U53, new_P2_ADD_394_U54,
    new_P2_ADD_394_U55, new_P2_ADD_394_U56, new_P2_ADD_394_U57,
    new_P2_ADD_394_U58, new_P2_ADD_394_U59, new_P2_ADD_394_U60,
    new_P2_ADD_394_U61, new_P2_ADD_394_U62, new_P2_ADD_394_U63,
    new_P2_ADD_394_U64, new_P2_ADD_394_U65, new_P2_ADD_394_U66,
    new_P2_ADD_394_U67, new_P2_ADD_394_U68, new_P2_ADD_394_U69,
    new_P2_ADD_394_U70, new_P2_ADD_394_U71, new_P2_ADD_394_U72,
    new_P2_ADD_394_U73, new_P2_ADD_394_U74, new_P2_ADD_394_U75,
    new_P2_ADD_394_U76, new_P2_ADD_394_U77, new_P2_ADD_394_U78,
    new_P2_ADD_394_U79, new_P2_ADD_394_U80, new_P2_ADD_394_U81,
    new_P2_ADD_394_U82, new_P2_ADD_394_U83, new_P2_ADD_394_U84,
    new_P2_ADD_394_U85, new_P2_ADD_394_U86, new_P2_ADD_394_U87,
    new_P2_ADD_394_U88, new_P2_ADD_394_U89, new_P2_ADD_394_U90,
    new_P2_ADD_394_U91, new_P2_ADD_394_U92, new_P2_ADD_394_U93,
    new_P2_ADD_394_U94, new_P2_ADD_394_U95, new_P2_ADD_394_U96,
    new_P2_ADD_394_U97, new_P2_ADD_394_U98, new_P2_ADD_394_U99,
    new_P2_ADD_394_U100, new_P2_ADD_394_U101, new_P2_ADD_394_U102,
    new_P2_ADD_394_U103, new_P2_ADD_394_U104, new_P2_ADD_394_U105,
    new_P2_ADD_394_U106, new_P2_ADD_394_U107, new_P2_ADD_394_U108,
    new_P2_ADD_394_U109, new_P2_ADD_394_U110, new_P2_ADD_394_U111,
    new_P2_ADD_394_U112, new_P2_ADD_394_U113, new_P2_ADD_394_U114,
    new_P2_ADD_394_U115, new_P2_ADD_394_U116, new_P2_ADD_394_U117,
    new_P2_ADD_394_U118, new_P2_ADD_394_U119, new_P2_ADD_394_U120,
    new_P2_ADD_394_U121, new_P2_ADD_394_U122, new_P2_ADD_394_U123,
    new_P2_ADD_394_U124, new_P2_ADD_394_U125, new_P2_ADD_394_U126,
    new_P2_ADD_394_U127, new_P2_ADD_394_U128, new_P2_ADD_394_U129,
    new_P2_ADD_394_U130, new_P2_ADD_394_U131, new_P2_ADD_394_U132,
    new_P2_ADD_394_U133, new_P2_ADD_394_U134, new_P2_ADD_394_U135,
    new_P2_ADD_394_U136, new_P2_ADD_394_U137, new_P2_ADD_394_U138,
    new_P2_ADD_394_U139, new_P2_ADD_394_U140, new_P2_ADD_394_U141,
    new_P2_ADD_394_U142, new_P2_ADD_394_U143, new_P2_ADD_394_U144,
    new_P2_ADD_394_U145, new_P2_ADD_394_U146, new_P2_ADD_394_U147,
    new_P2_ADD_394_U148, new_P2_ADD_394_U149, new_P2_ADD_394_U150,
    new_P2_ADD_394_U151, new_P2_ADD_394_U152, new_P2_ADD_394_U153,
    new_P2_ADD_394_U154, new_P2_ADD_394_U155, new_P2_ADD_394_U156,
    new_P2_ADD_394_U157, new_P2_ADD_394_U158, new_P2_ADD_394_U159,
    new_P2_ADD_394_U160, new_P2_ADD_394_U161, new_P2_ADD_394_U162,
    new_P2_ADD_394_U163, new_P2_ADD_394_U164, new_P2_ADD_394_U165,
    new_P2_ADD_394_U166, new_P2_ADD_394_U167, new_P2_ADD_394_U168,
    new_P2_ADD_394_U169, new_P2_ADD_394_U170, new_P2_ADD_394_U171,
    new_P2_ADD_394_U172, new_P2_ADD_394_U173, new_P2_ADD_394_U174,
    new_P2_ADD_394_U175, new_P2_ADD_394_U176, new_P2_ADD_394_U177,
    new_P2_ADD_394_U178, new_P2_ADD_394_U179, new_P2_ADD_394_U180,
    new_P2_ADD_394_U181, new_P2_ADD_394_U182, new_P2_ADD_394_U183,
    new_P2_ADD_394_U184, new_P2_ADD_394_U185, new_P2_ADD_394_U186,
    new_P2_R2267_U6, new_P2_R2267_U7, new_P2_R2267_U8, new_P2_R2267_U9,
    new_P2_R2267_U10, new_P2_R2267_U11, new_P2_R2267_U12, new_P2_R2267_U13,
    new_P2_R2267_U14, new_P2_R2267_U15, new_P2_R2267_U16, new_P2_R2267_U17,
    new_P2_R2267_U18, new_P2_R2267_U19, new_P2_R2267_U20, new_P2_R2267_U21,
    new_P2_R2267_U22, new_P2_R2267_U23, new_P2_R2267_U24, new_P2_R2267_U25,
    new_P2_R2267_U26, new_P2_R2267_U27, new_P2_R2267_U28, new_P2_R2267_U29,
    new_P2_R2267_U30, new_P2_R2267_U31, new_P2_R2267_U32, new_P2_R2267_U33,
    new_P2_R2267_U34, new_P2_R2267_U35, new_P2_R2267_U36, new_P2_R2267_U37,
    new_P2_R2267_U38, new_P2_R2267_U39, new_P2_R2267_U40, new_P2_R2267_U41,
    new_P2_R2267_U42, new_P2_R2267_U43, new_P2_R2267_U44, new_P2_R2267_U45,
    new_P2_R2267_U46, new_P2_R2267_U47, new_P2_R2267_U48, new_P2_R2267_U49,
    new_P2_R2267_U50, new_P2_R2267_U51, new_P2_R2267_U52, new_P2_R2267_U53,
    new_P2_R2267_U54, new_P2_R2267_U55, new_P2_R2267_U56, new_P2_R2267_U57,
    new_P2_R2267_U58, new_P2_R2267_U59, new_P2_R2267_U60, new_P2_R2267_U61,
    new_P2_R2267_U62, new_P2_R2267_U63, new_P2_R2267_U64, new_P2_R2267_U65,
    new_P2_R2267_U66, new_P2_R2267_U67, new_P2_R2267_U68, new_P2_R2267_U69,
    new_P2_R2267_U70, new_P2_R2267_U71, new_P2_R2267_U72, new_P2_R2267_U73,
    new_P2_R2267_U74, new_P2_R2267_U75, new_P2_R2267_U76, new_P2_R2267_U77,
    new_P2_R2267_U78, new_P2_R2267_U79, new_P2_R2267_U80, new_P2_R2267_U81,
    new_P2_R2267_U82, new_P2_R2267_U83, new_P2_R2267_U84, new_P2_R2267_U85,
    new_P2_R2267_U86, new_P2_R2267_U87, new_P2_R2267_U88, new_P2_R2267_U89,
    new_P2_R2267_U90, new_P2_R2267_U91, new_P2_R2267_U92, new_P2_R2267_U93,
    new_P2_R2267_U94, new_P2_R2267_U95, new_P2_R2267_U96, new_P2_R2267_U97,
    new_P2_R2267_U98, new_P2_R2267_U99, new_P2_R2267_U100,
    new_P2_R2267_U101, new_P2_R2267_U102, new_P2_R2267_U103,
    new_P2_R2267_U104, new_P2_R2267_U105, new_P2_R2267_U106,
    new_P2_R2267_U107, new_P2_R2267_U108, new_P2_R2267_U109,
    new_P2_R2267_U110, new_P2_R2267_U111, new_P2_R2267_U112,
    new_P2_R2267_U113, new_P2_R2267_U114, new_P2_R2267_U115,
    new_P2_R2267_U116, new_P2_R2267_U117, new_P2_R2267_U118,
    new_P2_R2267_U119, new_P2_R2267_U120, new_P2_R2267_U121,
    new_P2_R2267_U122, new_P2_R2267_U123, new_P2_R2267_U124,
    new_P2_R2267_U125, new_P2_R2267_U126, new_P2_R2267_U127,
    new_P2_R2267_U128, new_P2_R2267_U129, new_P2_R2267_U130,
    new_P2_R2267_U131, new_P2_R2267_U132, new_P2_R2267_U133,
    new_P2_R2267_U134, new_P2_R2267_U135, new_P2_R2267_U136,
    new_P2_R2267_U137, new_P2_R2267_U138, new_P2_R2267_U139,
    new_P2_R2267_U140, new_P2_R2267_U141, new_P2_R2267_U142,
    new_P2_R2267_U143, new_P2_R2267_U144, new_P2_R2267_U145,
    new_P2_R2267_U146, new_P2_R2267_U147, new_P2_R2267_U148,
    new_P2_R2267_U149, new_P2_R2267_U150, new_P2_R2267_U151,
    new_P2_R2267_U152, new_P2_R2267_U153, new_P2_R2267_U154,
    new_P2_R2267_U155, new_P2_R2267_U156, new_P2_R2267_U157,
    new_P2_R2267_U158, new_P2_R2267_U159, new_P2_R2267_U160,
    new_P2_R2267_U161, new_P2_R2267_U162, new_P2_R2267_U163,
    new_P2_R2267_U164, new_P2_R2267_U165, new_P2_R2267_U166,
    new_P2_ADD_371_1212_U4, new_P2_ADD_371_1212_U5, new_P2_ADD_371_1212_U6,
    new_P2_ADD_371_1212_U7, new_P2_ADD_371_1212_U8, new_P2_ADD_371_1212_U9,
    new_P2_ADD_371_1212_U10, new_P2_ADD_371_1212_U11,
    new_P2_ADD_371_1212_U12, new_P2_ADD_371_1212_U13,
    new_P2_ADD_371_1212_U14, new_P2_ADD_371_1212_U15,
    new_P2_ADD_371_1212_U16, new_P2_ADD_371_1212_U17,
    new_P2_ADD_371_1212_U18, new_P2_ADD_371_1212_U19,
    new_P2_ADD_371_1212_U20, new_P2_ADD_371_1212_U21,
    new_P2_ADD_371_1212_U22, new_P2_ADD_371_1212_U23,
    new_P2_ADD_371_1212_U24, new_P2_ADD_371_1212_U25,
    new_P2_ADD_371_1212_U26, new_P2_ADD_371_1212_U27,
    new_P2_ADD_371_1212_U28, new_P2_ADD_371_1212_U29,
    new_P2_ADD_371_1212_U30, new_P2_ADD_371_1212_U31,
    new_P2_ADD_371_1212_U32, new_P2_ADD_371_1212_U33,
    new_P2_ADD_371_1212_U34, new_P2_ADD_371_1212_U35,
    new_P2_ADD_371_1212_U36, new_P2_ADD_371_1212_U37,
    new_P2_ADD_371_1212_U38, new_P2_ADD_371_1212_U39,
    new_P2_ADD_371_1212_U40, new_P2_ADD_371_1212_U41,
    new_P2_ADD_371_1212_U42, new_P2_ADD_371_1212_U43,
    new_P2_ADD_371_1212_U44, new_P2_ADD_371_1212_U45,
    new_P2_ADD_371_1212_U46, new_P2_ADD_371_1212_U47,
    new_P2_ADD_371_1212_U48, new_P2_ADD_371_1212_U49,
    new_P2_ADD_371_1212_U50, new_P2_ADD_371_1212_U51,
    new_P2_ADD_371_1212_U52, new_P2_ADD_371_1212_U53,
    new_P2_ADD_371_1212_U54, new_P2_ADD_371_1212_U55,
    new_P2_ADD_371_1212_U56, new_P2_ADD_371_1212_U57,
    new_P2_ADD_371_1212_U58, new_P2_ADD_371_1212_U59,
    new_P2_ADD_371_1212_U60, new_P2_ADD_371_1212_U61,
    new_P2_ADD_371_1212_U62, new_P2_ADD_371_1212_U63,
    new_P2_ADD_371_1212_U64, new_P2_ADD_371_1212_U65,
    new_P2_ADD_371_1212_U66, new_P2_ADD_371_1212_U67,
    new_P2_ADD_371_1212_U68, new_P2_ADD_371_1212_U69,
    new_P2_ADD_371_1212_U70, new_P2_ADD_371_1212_U71,
    new_P2_ADD_371_1212_U72, new_P2_ADD_371_1212_U73,
    new_P2_ADD_371_1212_U74, new_P2_ADD_371_1212_U75,
    new_P2_ADD_371_1212_U76, new_P2_ADD_371_1212_U77,
    new_P2_ADD_371_1212_U78, new_P2_ADD_371_1212_U79,
    new_P2_ADD_371_1212_U80, new_P2_ADD_371_1212_U81,
    new_P2_ADD_371_1212_U82, new_P2_ADD_371_1212_U83,
    new_P2_ADD_371_1212_U84, new_P2_ADD_371_1212_U85,
    new_P2_ADD_371_1212_U86, new_P2_ADD_371_1212_U87,
    new_P2_ADD_371_1212_U88, new_P2_ADD_371_1212_U89,
    new_P2_ADD_371_1212_U90, new_P2_ADD_371_1212_U91,
    new_P2_ADD_371_1212_U92, new_P2_ADD_371_1212_U93,
    new_P2_ADD_371_1212_U94, new_P2_ADD_371_1212_U95,
    new_P2_ADD_371_1212_U96, new_P2_ADD_371_1212_U97,
    new_P2_ADD_371_1212_U98, new_P2_ADD_371_1212_U99,
    new_P2_ADD_371_1212_U100, new_P2_ADD_371_1212_U101,
    new_P2_ADD_371_1212_U102, new_P2_ADD_371_1212_U103,
    new_P2_ADD_371_1212_U104, new_P2_ADD_371_1212_U105,
    new_P2_ADD_371_1212_U106, new_P2_ADD_371_1212_U107,
    new_P2_ADD_371_1212_U108, new_P2_ADD_371_1212_U109,
    new_P2_ADD_371_1212_U110, new_P2_ADD_371_1212_U111,
    new_P2_ADD_371_1212_U112, new_P2_ADD_371_1212_U113,
    new_P2_ADD_371_1212_U114, new_P2_ADD_371_1212_U115,
    new_P2_ADD_371_1212_U116, new_P2_ADD_371_1212_U117,
    new_P2_ADD_371_1212_U118, new_P2_ADD_371_1212_U119,
    new_P2_ADD_371_1212_U120, new_P2_ADD_371_1212_U121,
    new_P2_ADD_371_1212_U122, new_P2_ADD_371_1212_U123,
    new_P2_ADD_371_1212_U124, new_P2_ADD_371_1212_U125,
    new_P2_ADD_371_1212_U126, new_P2_ADD_371_1212_U127,
    new_P2_ADD_371_1212_U128, new_P2_ADD_371_1212_U129,
    new_P2_ADD_371_1212_U130, new_P2_ADD_371_1212_U131,
    new_P2_ADD_371_1212_U132, new_P2_ADD_371_1212_U133,
    new_P2_ADD_371_1212_U134, new_P2_ADD_371_1212_U135,
    new_P2_ADD_371_1212_U136, new_P2_ADD_371_1212_U137,
    new_P2_ADD_371_1212_U138, new_P2_ADD_371_1212_U139,
    new_P2_ADD_371_1212_U140, new_P2_ADD_371_1212_U141,
    new_P2_ADD_371_1212_U142, new_P2_ADD_371_1212_U143,
    new_P2_ADD_371_1212_U144, new_P2_ADD_371_1212_U145,
    new_P2_ADD_371_1212_U146, new_P2_ADD_371_1212_U147,
    new_P2_ADD_371_1212_U148, new_P2_ADD_371_1212_U149,
    new_P2_ADD_371_1212_U150, new_P2_ADD_371_1212_U151,
    new_P2_ADD_371_1212_U152, new_P2_ADD_371_1212_U153,
    new_P2_ADD_371_1212_U154, new_P2_ADD_371_1212_U155,
    new_P2_ADD_371_1212_U156, new_P2_ADD_371_1212_U157,
    new_P2_ADD_371_1212_U158, new_P2_ADD_371_1212_U159,
    new_P2_ADD_371_1212_U160, new_P2_ADD_371_1212_U161,
    new_P2_ADD_371_1212_U162, new_P2_ADD_371_1212_U163,
    new_P2_ADD_371_1212_U164, new_P2_ADD_371_1212_U165,
    new_P2_ADD_371_1212_U166, new_P2_ADD_371_1212_U167,
    new_P2_ADD_371_1212_U168, new_P2_ADD_371_1212_U169,
    new_P2_ADD_371_1212_U170, new_P2_ADD_371_1212_U171,
    new_P2_ADD_371_1212_U172, new_P2_ADD_371_1212_U173,
    new_P2_ADD_371_1212_U174, new_P2_ADD_371_1212_U175,
    new_P2_ADD_371_1212_U176, new_P2_ADD_371_1212_U177,
    new_P2_ADD_371_1212_U178, new_P2_ADD_371_1212_U179,
    new_P2_ADD_371_1212_U180, new_P2_ADD_371_1212_U181,
    new_P2_ADD_371_1212_U182, new_P2_ADD_371_1212_U183,
    new_P2_ADD_371_1212_U184, new_P2_ADD_371_1212_U185,
    new_P2_ADD_371_1212_U186, new_P2_ADD_371_1212_U187,
    new_P2_ADD_371_1212_U188, new_P2_ADD_371_1212_U189,
    new_P2_ADD_371_1212_U190, new_P2_ADD_371_1212_U191,
    new_P2_ADD_371_1212_U192, new_P2_ADD_371_1212_U193,
    new_P2_ADD_371_1212_U194, new_P2_ADD_371_1212_U195,
    new_P2_ADD_371_1212_U196, new_P2_ADD_371_1212_U197,
    new_P2_ADD_371_1212_U198, new_P2_ADD_371_1212_U199,
    new_P2_ADD_371_1212_U200, new_P2_ADD_371_1212_U201,
    new_P2_ADD_371_1212_U202, new_P2_ADD_371_1212_U203,
    new_P2_ADD_371_1212_U204, new_P2_ADD_371_1212_U205,
    new_P2_ADD_371_1212_U206, new_P2_ADD_371_1212_U207,
    new_P2_ADD_371_1212_U208, new_P2_ADD_371_1212_U209,
    new_P2_ADD_371_1212_U210, new_P2_ADD_371_1212_U211,
    new_P2_ADD_371_1212_U212, new_P2_ADD_371_1212_U213,
    new_P2_ADD_371_1212_U214, new_P2_ADD_371_1212_U215,
    new_P2_ADD_371_1212_U216, new_P2_ADD_371_1212_U217,
    new_P2_ADD_371_1212_U218, new_P2_ADD_371_1212_U219,
    new_P2_ADD_371_1212_U220, new_P2_ADD_371_1212_U221,
    new_P2_ADD_371_1212_U222, new_P2_ADD_371_1212_U223,
    new_P2_ADD_371_1212_U224, new_P2_ADD_371_1212_U225,
    new_P2_ADD_371_1212_U226, new_P2_ADD_371_1212_U227,
    new_P2_ADD_371_1212_U228, new_P2_ADD_371_1212_U229,
    new_P2_ADD_371_1212_U230, new_P2_ADD_371_1212_U231,
    new_P2_ADD_371_1212_U232, new_P2_ADD_371_1212_U233,
    new_P2_ADD_371_1212_U234, new_P2_ADD_371_1212_U235,
    new_P2_ADD_371_1212_U236, new_P2_ADD_371_1212_U237,
    new_P2_ADD_371_1212_U238, new_P2_ADD_371_1212_U239,
    new_P2_ADD_371_1212_U240, new_P2_ADD_371_1212_U241,
    new_P2_ADD_371_1212_U242, new_P2_ADD_371_1212_U243,
    new_P2_ADD_371_1212_U244, new_P2_ADD_371_1212_U245,
    new_P2_ADD_371_1212_U246, new_P2_ADD_371_1212_U247,
    new_P2_ADD_371_1212_U248, new_P2_ADD_371_1212_U249,
    new_P2_ADD_371_1212_U250, new_P2_ADD_371_1212_U251,
    new_P2_ADD_371_1212_U252, new_P2_ADD_371_1212_U253,
    new_P2_ADD_371_1212_U254, new_P2_ADD_371_1212_U255,
    new_P2_ADD_371_1212_U256, new_P2_ADD_371_1212_U257,
    new_P2_ADD_371_1212_U258, new_P2_ADD_371_1212_U259,
    new_P2_ADD_371_1212_U260, new_P2_ADD_371_1212_U261,
    new_P2_ADD_371_1212_U262, new_P2_ADD_371_1212_U263,
    new_P2_ADD_371_1212_U264, new_P2_ADD_371_1212_U265,
    new_P2_ADD_371_1212_U266, new_P2_ADD_371_1212_U267,
    new_P2_ADD_371_1212_U268, new_P2_ADD_371_1212_U269,
    new_P2_ADD_371_1212_U270, new_P2_ADD_371_1212_U271,
    new_P2_ADD_371_1212_U272, new_P2_ADD_371_1212_U273,
    new_P2_ADD_371_1212_U274, new_P2_ADD_371_1212_U275,
    new_P2_ADD_371_1212_U276, new_P2_ADD_371_1212_U277,
    new_P2_ADD_371_1212_U278, new_P2_ADD_371_1212_U279,
    new_P2_ADD_371_1212_U280, new_P2_ADD_371_1212_U281,
    new_P2_ADD_371_1212_U282, new_P1_R2027_U5, new_P1_R2027_U6,
    new_P1_R2027_U7, new_P1_R2027_U8, new_P1_R2027_U9, new_P1_R2027_U10,
    new_P1_R2027_U11, new_P1_R2027_U12, new_P1_R2027_U13, new_P1_R2027_U14,
    new_P1_R2027_U15, new_P1_R2027_U16, new_P1_R2027_U17, new_P1_R2027_U18,
    new_P1_R2027_U19, new_P1_R2027_U20, new_P1_R2027_U21, new_P1_R2027_U22,
    new_P1_R2027_U23, new_P1_R2027_U24, new_P1_R2027_U25, new_P1_R2027_U26,
    new_P1_R2027_U27, new_P1_R2027_U28, new_P1_R2027_U29, new_P1_R2027_U30,
    new_P1_R2027_U31, new_P1_R2027_U32, new_P1_R2027_U33, new_P1_R2027_U34,
    new_P1_R2027_U35, new_P1_R2027_U36, new_P1_R2027_U37, new_P1_R2027_U38,
    new_P1_R2027_U39, new_P1_R2027_U40, new_P1_R2027_U41, new_P1_R2027_U42,
    new_P1_R2027_U43, new_P1_R2027_U44, new_P1_R2027_U45, new_P1_R2027_U46,
    new_P1_R2027_U47, new_P1_R2027_U48, new_P1_R2027_U49, new_P1_R2027_U50,
    new_P1_R2027_U51, new_P1_R2027_U52, new_P1_R2027_U53, new_P1_R2027_U54,
    new_P1_R2027_U55, new_P1_R2027_U56, new_P1_R2027_U57, new_P1_R2027_U58,
    new_P1_R2027_U59, new_P1_R2027_U60, new_P1_R2027_U61, new_P1_R2027_U62,
    new_P1_R2027_U63, new_P1_R2027_U64, new_P1_R2027_U65, new_P1_R2027_U66,
    new_P1_R2027_U67, new_P1_R2027_U68, new_P1_R2027_U69, new_P1_R2027_U70,
    new_P1_R2027_U71, new_P1_R2027_U72, new_P1_R2027_U73, new_P1_R2027_U74,
    new_P1_R2027_U75, new_P1_R2027_U76, new_P1_R2027_U77, new_P1_R2027_U78,
    new_P1_R2027_U79, new_P1_R2027_U80, new_P1_R2027_U81, new_P1_R2027_U82,
    new_P1_R2027_U83, new_P1_R2027_U84, new_P1_R2027_U85, new_P1_R2027_U86,
    new_P1_R2027_U87, new_P1_R2027_U88, new_P1_R2027_U89, new_P1_R2027_U90,
    new_P1_R2027_U91, new_P1_R2027_U92, new_P1_R2027_U93, new_P1_R2027_U94,
    new_P1_R2027_U95, new_P1_R2027_U96, new_P1_R2027_U97, new_P1_R2027_U98,
    new_P1_R2027_U99, new_P1_R2027_U100, new_P1_R2027_U101,
    new_P1_R2027_U102, new_P1_R2027_U103, new_P1_R2027_U104,
    new_P1_R2027_U105, new_P1_R2027_U106, new_P1_R2027_U107,
    new_P1_R2027_U108, new_P1_R2027_U109, new_P1_R2027_U110,
    new_P1_R2027_U111, new_P1_R2027_U112, new_P1_R2027_U113,
    new_P1_R2027_U114, new_P1_R2027_U115, new_P1_R2027_U116,
    new_P1_R2027_U117, new_P1_R2027_U118, new_P1_R2027_U119,
    new_P1_R2027_U120, new_P1_R2027_U121, new_P1_R2027_U122,
    new_P1_R2027_U123, new_P1_R2027_U124, new_P1_R2027_U125,
    new_P1_R2027_U126, new_P1_R2027_U127, new_P1_R2027_U128,
    new_P1_R2027_U129, new_P1_R2027_U130, new_P1_R2027_U131,
    new_P1_R2027_U132, new_P1_R2027_U133, new_P1_R2027_U134,
    new_P1_R2027_U135, new_P1_R2027_U136, new_P1_R2027_U137,
    new_P1_R2027_U138, new_P1_R2027_U139, new_P1_R2027_U140,
    new_P1_R2027_U141, new_P1_R2027_U142, new_P1_R2027_U143,
    new_P1_R2027_U144, new_P1_R2027_U145, new_P1_R2027_U146,
    new_P1_R2027_U147, new_P1_R2027_U148, new_P1_R2027_U149,
    new_P1_R2027_U150, new_P1_R2027_U151, new_P1_R2027_U152,
    new_P1_R2027_U153, new_P1_R2027_U154, new_P1_R2027_U155,
    new_P1_R2027_U156, new_P1_R2027_U157, new_P1_R2027_U158,
    new_P1_R2027_U159, new_P1_R2027_U160, new_P1_R2027_U161,
    new_P1_R2027_U162, new_P1_R2027_U163, new_P1_R2027_U164,
    new_P1_R2027_U165, new_P1_R2027_U166, new_P1_R2027_U167,
    new_P1_R2027_U168, new_P1_R2027_U169, new_P1_R2027_U170,
    new_P1_R2027_U171, new_P1_R2027_U172, new_P1_R2027_U173,
    new_P1_R2027_U174, new_P1_R2027_U175, new_P1_R2027_U176,
    new_P1_R2027_U177, new_P1_R2027_U178, new_P1_R2027_U179,
    new_P1_R2027_U180, new_P1_R2027_U181, new_P1_R2027_U182,
    new_P1_R2027_U183, new_P1_R2027_U184, new_P1_R2027_U185,
    new_P1_R2027_U186, new_P1_R2027_U187, new_P1_R2027_U188,
    new_P1_R2027_U189, new_P1_R2027_U190, new_P1_R2027_U191,
    new_P1_R2027_U192, new_P1_R2027_U193, new_P1_R2027_U194,
    new_P1_R2027_U195, new_P1_R2027_U196, new_P1_R2027_U197,
    new_P1_R2027_U198, new_P1_R2027_U199, new_P1_R2027_U200,
    new_P1_R2027_U201, new_P1_R2027_U202, new_P1_R2182_U5, new_P1_R2182_U6,
    new_P1_R2182_U7, new_P1_R2182_U8, new_P1_R2182_U9, new_P1_R2182_U10,
    new_P1_R2182_U11, new_P1_R2182_U12, new_P1_R2182_U13, new_P1_R2182_U14,
    new_P1_R2182_U15, new_P1_R2182_U16, new_P1_R2182_U17, new_P1_R2182_U18,
    new_P1_R2182_U19, new_P1_R2182_U20, new_P1_R2182_U21, new_P1_R2182_U22,
    new_P1_R2182_U23, new_P1_R2182_U24, new_P1_R2182_U25, new_P1_R2182_U26,
    new_P1_R2182_U27, new_P1_R2182_U28, new_P1_R2182_U29, new_P1_R2182_U30,
    new_P1_R2182_U31, new_P1_R2182_U32, new_P1_R2182_U33, new_P1_R2182_U34,
    new_P1_R2182_U35, new_P1_R2182_U36, new_P1_R2182_U37, new_P1_R2182_U38,
    new_P1_R2182_U39, new_P1_R2182_U40, new_P1_R2182_U41, new_P1_R2182_U42,
    new_P1_R2182_U43, new_P1_R2182_U44, new_P1_R2182_U45, new_P1_R2182_U46,
    new_P1_R2182_U47, new_P1_R2182_U48, new_P1_R2182_U49, new_P1_R2182_U50,
    new_P1_R2182_U51, new_P1_R2182_U52, new_P1_R2182_U53, new_P1_R2182_U54,
    new_P1_R2182_U55, new_P1_R2182_U56, new_P1_R2182_U57, new_P1_R2182_U58,
    new_P1_R2182_U59, new_P1_R2182_U60, new_P1_R2182_U61, new_P1_R2182_U62,
    new_P1_R2182_U63, new_P1_R2182_U64, new_P1_R2182_U65, new_P1_R2182_U66,
    new_P1_R2182_U67, new_P1_R2182_U68, new_P1_R2182_U69, new_P1_R2182_U70,
    new_P1_R2182_U71, new_P1_R2182_U72, new_P1_R2182_U73, new_P1_R2182_U74,
    new_P1_R2182_U75, new_P1_R2182_U76, new_P1_R2182_U77, new_P1_R2182_U78,
    new_P1_R2182_U79, new_P1_R2182_U80, new_P1_R2182_U81, new_P1_R2182_U82,
    new_P1_R2182_U83, new_P1_R2182_U84, new_P1_R2182_U85, new_P1_R2182_U86,
    new_P1_R2144_U5, new_P1_R2144_U6, new_P1_R2144_U7, new_P1_R2144_U8,
    new_P1_R2144_U9, new_P1_R2144_U10, new_P1_R2144_U11, new_P1_R2144_U12,
    new_P1_R2144_U13, new_P1_R2144_U14, new_P1_R2144_U15, new_P1_R2144_U16,
    new_P1_R2144_U17, new_P1_R2144_U18, new_P1_R2144_U19, new_P1_R2144_U20,
    new_P1_R2144_U21, new_P1_R2144_U22, new_P1_R2144_U23, new_P1_R2144_U24,
    new_P1_R2144_U25, new_P1_R2144_U26, new_P1_R2144_U27, new_P1_R2144_U28,
    new_P1_R2144_U29, new_P1_R2144_U30, new_P1_R2144_U31, new_P1_R2144_U32,
    new_P1_R2144_U33, new_P1_R2144_U34, new_P1_R2144_U35, new_P1_R2144_U36,
    new_P1_R2144_U37, new_P1_R2144_U38, new_P1_R2144_U39, new_P1_R2144_U40,
    new_P1_R2144_U41, new_P1_R2144_U42, new_P1_R2144_U43, new_P1_R2144_U44,
    new_P1_R2144_U45, new_P1_R2144_U46, new_P1_R2144_U47, new_P1_R2144_U48,
    new_P1_R2144_U49, new_P1_R2144_U50, new_P1_R2144_U51, new_P1_R2144_U52,
    new_P1_R2144_U53, new_P1_R2144_U54, new_P1_R2144_U55, new_P1_R2144_U56,
    new_P1_R2144_U57, new_P1_R2144_U58, new_P1_R2144_U59, new_P1_R2144_U60,
    new_P1_R2144_U61, new_P1_R2144_U62, new_P1_R2144_U63, new_P1_R2144_U64,
    new_P1_R2144_U65, new_P1_R2144_U66, new_P1_R2144_U67, new_P1_R2144_U68,
    new_P1_R2144_U69, new_P1_R2144_U70, new_P1_R2144_U71, new_P1_R2144_U72,
    new_P1_R2144_U73, new_P1_R2144_U74, new_P1_R2144_U75, new_P1_R2144_U76,
    new_P1_R2144_U77, new_P1_R2144_U78, new_P1_R2144_U79, new_P1_R2144_U80,
    new_P1_R2144_U81, new_P1_R2144_U82, new_P1_R2144_U83, new_P1_R2144_U84,
    new_P1_R2144_U85, new_P1_R2144_U86, new_P1_R2144_U87, new_P1_R2144_U88,
    new_P1_R2144_U89, new_P1_R2144_U90, new_P1_R2144_U91, new_P1_R2144_U92,
    new_P1_R2144_U93, new_P1_R2144_U94, new_P1_R2144_U95, new_P1_R2144_U96,
    new_P1_R2144_U97, new_P1_R2144_U98, new_P1_R2144_U99,
    new_P1_R2144_U100, new_P1_R2144_U101, new_P1_R2144_U102,
    new_P1_R2144_U103, new_P1_R2144_U104, new_P1_R2144_U105,
    new_P1_R2144_U106, new_P1_R2144_U107, new_P1_R2144_U108,
    new_P1_R2144_U109, new_P1_R2144_U110, new_P1_R2144_U111,
    new_P1_R2144_U112, new_P1_R2144_U113, new_P1_R2144_U114,
    new_P1_R2144_U115, new_P1_R2144_U116, new_P1_R2144_U117,
    new_P1_R2144_U118, new_P1_R2144_U119, new_P1_R2144_U120,
    new_P1_R2144_U121, new_P1_R2144_U122, new_P1_R2144_U123,
    new_P1_R2144_U124, new_P1_R2144_U125, new_P1_R2144_U126,
    new_P1_R2144_U127, new_P1_R2144_U128, new_P1_R2144_U129,
    new_P1_R2144_U130, new_P1_R2144_U131, new_P1_R2144_U132,
    new_P1_R2144_U133, new_P1_R2144_U134, new_P1_R2144_U135,
    new_P1_R2144_U136, new_P1_R2144_U137, new_P1_R2144_U138,
    new_P1_R2144_U139, new_P1_R2144_U140, new_P1_R2144_U141,
    new_P1_R2144_U142, new_P1_R2144_U143, new_P1_R2144_U144,
    new_P1_R2144_U145, new_P1_R2144_U146, new_P1_R2144_U147,
    new_P1_R2144_U148, new_P1_R2144_U149, new_P1_R2144_U150,
    new_P1_R2144_U151, new_P1_R2144_U152, new_P1_R2144_U153,
    new_P1_R2144_U154, new_P1_R2144_U155, new_P1_R2144_U156,
    new_P1_R2144_U157, new_P1_R2144_U158, new_P1_R2144_U159,
    new_P1_R2144_U160, new_P1_R2144_U161, new_P1_R2144_U162,
    new_P1_R2144_U163, new_P1_R2144_U164, new_P1_R2144_U165,
    new_P1_R2144_U166, new_P1_R2144_U167, new_P1_R2144_U168,
    new_P1_R2144_U169, new_P1_R2144_U170, new_P1_R2144_U171,
    new_P1_R2144_U172, new_P1_R2144_U173, new_P1_R2144_U174,
    new_P1_R2144_U175, new_P1_R2144_U176, new_P1_R2144_U177,
    new_P1_R2144_U178, new_P1_R2144_U179, new_P1_R2144_U180,
    new_P1_R2144_U181, new_P1_R2144_U182, new_P1_R2144_U183,
    new_P1_R2144_U184, new_P1_R2144_U185, new_P1_R2144_U186,
    new_P1_R2144_U187, new_P1_R2144_U188, new_P1_R2144_U189,
    new_P1_R2144_U190, new_P1_R2144_U191, new_P1_R2144_U192,
    new_P1_R2144_U193, new_P1_R2144_U194, new_P1_R2144_U195,
    new_P1_R2144_U196, new_P1_R2144_U197, new_P1_R2144_U198,
    new_P1_R2144_U199, new_P1_R2144_U200, new_P1_R2144_U201,
    new_P1_R2144_U202, new_P1_R2144_U203, new_P1_R2144_U204,
    new_P1_R2144_U205, new_P1_R2144_U206, new_P1_R2144_U207,
    new_P1_R2144_U208, new_P1_R2144_U209, new_P1_R2144_U210,
    new_P1_R2144_U211, new_P1_R2144_U212, new_P1_R2144_U213,
    new_P1_R2144_U214, new_P1_R2144_U215, new_P1_R2144_U216,
    new_P1_R2144_U217, new_P1_R2144_U218, new_P1_R2144_U219,
    new_P1_R2144_U220, new_P1_R2144_U221, new_P1_R2144_U222,
    new_P1_R2144_U223, new_P1_R2144_U224, new_P1_R2144_U225,
    new_P1_R2144_U226, new_P1_R2144_U227, new_P1_R2144_U228,
    new_P1_R2144_U229, new_P1_R2144_U230, new_P1_R2144_U231,
    new_P1_R2144_U232, new_P1_R2144_U233, new_P1_R2144_U234,
    new_P1_R2144_U235, new_P1_R2144_U236, new_P1_R2144_U237,
    new_P1_R2144_U238, new_P1_R2144_U239, new_P1_R2144_U240,
    new_P1_R2144_U241, new_P1_R2144_U242, new_P1_R2144_U243,
    new_P1_R2144_U244, new_P1_R2144_U245, new_P1_R2144_U246,
    new_P1_R2144_U247, new_P1_R2144_U248, new_P1_R2144_U249,
    new_P1_R2144_U250, new_P1_R2144_U251, new_P1_R2144_U252,
    new_P1_R2144_U253, new_P1_R2144_U254, new_P1_R2144_U255,
    new_P1_R2144_U256, new_P1_R2144_U257, new_P1_R2144_U258,
    new_P1_R2144_U259, new_P1_R2144_U260, new_P1_R2278_U5, new_P1_R2278_U6,
    new_P1_R2278_U7, new_P1_R2278_U8, new_P1_R2278_U9, new_P1_R2278_U10,
    new_P1_R2278_U11, new_P1_R2278_U12, new_P1_R2278_U13, new_P1_R2278_U14,
    new_P1_R2278_U15, new_P1_R2278_U16, new_P1_R2278_U17, new_P1_R2278_U18,
    new_P1_R2278_U19, new_P1_R2278_U20, new_P1_R2278_U21, new_P1_R2278_U22,
    new_P1_R2278_U23, new_P1_R2278_U24, new_P1_R2278_U25, new_P1_R2278_U26,
    new_P1_R2278_U27, new_P1_R2278_U28, new_P1_R2278_U29, new_P1_R2278_U30,
    new_P1_R2278_U31, new_P1_R2278_U32, new_P1_R2278_U33, new_P1_R2278_U34,
    new_P1_R2278_U35, new_P1_R2278_U36, new_P1_R2278_U37, new_P1_R2278_U38,
    new_P1_R2278_U39, new_P1_R2278_U40, new_P1_R2278_U41, new_P1_R2278_U42,
    new_P1_R2278_U43, new_P1_R2278_U44, new_P1_R2278_U45, new_P1_R2278_U46,
    new_P1_R2278_U47, new_P1_R2278_U48, new_P1_R2278_U49, new_P1_R2278_U50,
    new_P1_R2278_U51, new_P1_R2278_U52, new_P1_R2278_U53, new_P1_R2278_U54,
    new_P1_R2278_U55, new_P1_R2278_U56, new_P1_R2278_U57, new_P1_R2278_U58,
    new_P1_R2278_U59, new_P1_R2278_U60, new_P1_R2278_U61, new_P1_R2278_U62,
    new_P1_R2278_U63, new_P1_R2278_U64, new_P1_R2278_U65, new_P1_R2278_U66,
    new_P1_R2278_U67, new_P1_R2278_U68, new_P1_R2278_U69, new_P1_R2278_U70,
    new_P1_R2278_U71, new_P1_R2278_U72, new_P1_R2278_U73, new_P1_R2278_U74,
    new_P1_R2278_U75, new_P1_R2278_U76, new_P1_R2278_U77, new_P1_R2278_U78,
    new_P1_R2278_U79, new_P1_R2278_U80, new_P1_R2278_U81, new_P1_R2278_U82,
    new_P1_R2278_U83, new_P1_R2278_U84, new_P1_R2278_U85, new_P1_R2278_U86,
    new_P1_R2278_U87, new_P1_R2278_U88, new_P1_R2278_U89, new_P1_R2278_U90,
    new_P1_R2278_U91, new_P1_R2278_U92, new_P1_R2278_U93, new_P1_R2278_U94,
    new_P1_R2278_U95, new_P1_R2278_U96, new_P1_R2278_U97, new_P1_R2278_U98,
    new_P1_R2278_U99, new_P1_R2278_U100, new_P1_R2278_U101,
    new_P1_R2278_U102, new_P1_R2278_U103, new_P1_R2278_U104,
    new_P1_R2278_U105, new_P1_R2278_U106, new_P1_R2278_U107,
    new_P1_R2278_U108, new_P1_R2278_U109, new_P1_R2278_U110,
    new_P1_R2278_U111, new_P1_R2278_U112, new_P1_R2278_U113,
    new_P1_R2278_U114, new_P1_R2278_U115, new_P1_R2278_U116,
    new_P1_R2278_U117, new_P1_R2278_U118, new_P1_R2278_U119,
    new_P1_R2278_U120, new_P1_R2278_U121, new_P1_R2278_U122,
    new_P1_R2278_U123, new_P1_R2278_U124, new_P1_R2278_U125,
    new_P1_R2278_U126, new_P1_R2278_U127, new_P1_R2278_U128,
    new_P1_R2278_U129, new_P1_R2278_U130, new_P1_R2278_U131,
    new_P1_R2278_U132, new_P1_R2278_U133, new_P1_R2278_U134,
    new_P1_R2278_U135, new_P1_R2278_U136, new_P1_R2278_U137,
    new_P1_R2278_U138, new_P1_R2278_U139, new_P1_R2278_U140,
    new_P1_R2278_U141, new_P1_R2278_U142, new_P1_R2278_U143,
    new_P1_R2278_U144, new_P1_R2278_U145, new_P1_R2278_U146,
    new_P1_R2278_U147, new_P1_R2278_U148, new_P1_R2278_U149,
    new_P1_R2278_U150, new_P1_R2278_U151, new_P1_R2278_U152,
    new_P1_R2278_U153, new_P1_R2278_U154, new_P1_R2278_U155,
    new_P1_R2278_U156, new_P1_R2278_U157, new_P1_R2278_U158,
    new_P1_R2278_U159, new_P1_R2278_U160, new_P1_R2278_U161,
    new_P1_R2278_U162, new_P1_R2278_U163, new_P1_R2278_U164,
    new_P1_R2278_U165, new_P1_R2278_U166, new_P1_R2278_U167,
    new_P1_R2278_U168, new_P1_R2278_U169, new_P1_R2278_U170,
    new_P1_R2278_U171, new_P1_R2278_U172, new_P1_R2278_U173,
    new_P1_R2278_U174, new_P1_R2278_U175, new_P1_R2278_U176,
    new_P1_R2278_U177, new_P1_R2278_U178, new_P1_R2278_U179,
    new_P1_R2278_U180, new_P1_R2278_U181, new_P1_R2278_U182,
    new_P1_R2278_U183, new_P1_R2278_U184, new_P1_R2278_U185,
    new_P1_R2278_U186, new_P1_R2278_U187, new_P1_R2278_U188,
    new_P1_R2278_U189, new_P1_R2278_U190, new_P1_R2278_U191,
    new_P1_R2278_U192, new_P1_R2278_U193, new_P1_R2278_U194,
    new_P1_R2278_U195, new_P1_R2278_U196, new_P1_R2278_U197,
    new_P1_R2278_U198, new_P1_R2278_U199, new_P1_R2278_U200,
    new_P1_R2278_U201, new_P1_R2278_U202, new_P1_R2278_U203,
    new_P1_R2278_U204, new_P1_R2278_U205, new_P1_R2278_U206,
    new_P1_R2278_U207, new_P1_R2278_U208, new_P1_R2278_U209,
    new_P1_R2278_U210, new_P1_R2278_U211, new_P1_R2278_U212,
    new_P1_R2278_U213, new_P1_R2278_U214, new_P1_R2278_U215,
    new_P1_R2278_U216, new_P1_R2278_U217, new_P1_R2278_U218,
    new_P1_R2278_U219, new_P1_R2278_U220, new_P1_R2278_U221,
    new_P1_R2278_U222, new_P1_R2278_U223, new_P1_R2278_U224,
    new_P1_R2278_U225, new_P1_R2278_U226, new_P1_R2278_U227,
    new_P1_R2278_U228, new_P1_R2278_U229, new_P1_R2278_U230,
    new_P1_R2278_U231, new_P1_R2278_U232, new_P1_R2278_U233,
    new_P1_R2278_U234, new_P1_R2278_U235, new_P1_R2278_U236,
    new_P1_R2278_U237, new_P1_R2278_U238, new_P1_R2278_U239,
    new_P1_R2278_U240, new_P1_R2278_U241, new_P1_R2278_U242,
    new_P1_R2278_U243, new_P1_R2278_U244, new_P1_R2278_U245,
    new_P1_R2278_U246, new_P1_R2278_U247, new_P1_R2278_U248,
    new_P1_R2278_U249, new_P1_R2278_U250, new_P1_R2278_U251,
    new_P1_R2278_U252, new_P1_R2278_U253, new_P1_R2278_U254,
    new_P1_R2278_U255, new_P1_R2278_U256, new_P1_R2278_U257,
    new_P1_R2278_U258, new_P1_R2278_U259, new_P1_R2278_U260,
    new_P1_R2278_U261, new_P1_R2278_U262, new_P1_R2278_U263,
    new_P1_R2278_U264, new_P1_R2278_U265, new_P1_R2278_U266,
    new_P1_R2278_U267, new_P1_R2278_U268, new_P1_R2278_U269,
    new_P1_R2278_U270, new_P1_R2278_U271, new_P1_R2278_U272,
    new_P1_R2278_U273, new_P1_R2278_U274, new_P1_R2278_U275,
    new_P1_R2278_U276, new_P1_R2278_U277, new_P1_R2278_U278,
    new_P1_R2278_U279, new_P1_R2278_U280, new_P1_R2278_U281,
    new_P1_R2278_U282, new_P1_R2278_U283, new_P1_R2278_U284,
    new_P1_R2278_U285, new_P1_R2278_U286, new_P1_R2278_U287,
    new_P1_R2278_U288, new_P1_R2278_U289, new_P1_R2278_U290,
    new_P1_R2278_U291, new_P1_R2278_U292, new_P1_R2278_U293,
    new_P1_R2278_U294, new_P1_R2278_U295, new_P1_R2278_U296,
    new_P1_R2278_U297, new_P1_R2278_U298, new_P1_R2278_U299,
    new_P1_R2278_U300, new_P1_R2278_U301, new_P1_R2278_U302,
    new_P1_R2278_U303, new_P1_R2278_U304, new_P1_R2278_U305,
    new_P1_R2278_U306, new_P1_R2278_U307, new_P1_R2278_U308,
    new_P1_R2278_U309, new_P1_R2278_U310, new_P1_R2278_U311,
    new_P1_R2278_U312, new_P1_R2278_U313, new_P1_R2278_U314,
    new_P1_R2278_U315, new_P1_R2278_U316, new_P1_R2278_U317,
    new_P1_R2278_U318, new_P1_R2278_U319, new_P1_R2278_U320,
    new_P1_R2278_U321, new_P1_R2278_U322, new_P1_R2278_U323,
    new_P1_R2278_U324, new_P1_R2278_U325, new_P1_R2278_U326,
    new_P1_R2278_U327, new_P1_R2278_U328, new_P1_R2278_U329,
    new_P1_R2278_U330, new_P1_R2278_U331, new_P1_R2278_U332,
    new_P1_R2278_U333, new_P1_R2278_U334, new_P1_R2278_U335,
    new_P1_R2278_U336, new_P1_R2278_U337, new_P1_R2278_U338,
    new_P1_R2278_U339, new_P1_R2278_U340, new_P1_R2278_U341,
    new_P1_R2278_U342, new_P1_R2278_U343, new_P1_R2278_U344,
    new_P1_R2278_U345, new_P1_R2278_U346, new_P1_R2278_U347,
    new_P1_R2278_U348, new_P1_R2278_U349, new_P1_R2278_U350,
    new_P1_R2278_U351, new_P1_R2278_U352, new_P1_R2278_U353,
    new_P1_R2278_U354, new_P1_R2278_U355, new_P1_R2278_U356,
    new_P1_R2278_U357, new_P1_R2278_U358, new_P1_R2278_U359,
    new_P1_R2278_U360, new_P1_R2278_U361, new_P1_R2278_U362,
    new_P1_R2278_U363, new_P1_R2278_U364, new_P1_R2278_U365,
    new_P1_R2278_U366, new_P1_R2278_U367, new_P1_R2278_U368,
    new_P1_R2278_U369, new_P1_R2278_U370, new_P1_R2278_U371,
    new_P1_R2278_U372, new_P1_R2278_U373, new_P1_R2278_U374,
    new_P1_R2278_U375, new_P1_R2278_U376, new_P1_R2278_U377,
    new_P1_R2278_U378, new_P1_R2278_U379, new_P1_R2278_U380,
    new_P1_R2278_U381, new_P1_R2278_U382, new_P1_R2278_U383,
    new_P1_R2278_U384, new_P1_R2278_U385, new_P1_R2278_U386,
    new_P1_R2278_U387, new_P1_R2278_U388, new_P1_R2278_U389,
    new_P1_R2278_U390, new_P1_R2278_U391, new_P1_R2278_U392,
    new_P1_R2278_U393, new_P1_R2278_U394, new_P1_R2278_U395,
    new_P1_R2278_U396, new_P1_R2278_U397, new_P1_R2278_U398,
    new_P1_R2278_U399, new_P1_R2278_U400, new_P1_R2278_U401,
    new_P1_R2278_U402, new_P1_R2278_U403, new_P1_R2278_U404,
    new_P1_R2278_U405, new_P1_R2278_U406, new_P1_R2278_U407,
    new_P1_R2278_U408, new_P1_R2278_U409, new_P1_R2278_U410,
    new_P1_R2278_U411, new_P1_R2278_U412, new_P1_R2278_U413,
    new_P1_R2278_U414, new_P1_R2278_U415, new_P1_R2278_U416,
    new_P1_R2278_U417, new_P1_R2278_U418, new_P1_R2278_U419,
    new_P1_R2278_U420, new_P1_R2278_U421, new_P1_R2278_U422,
    new_P1_R2278_U423, new_P1_R2278_U424, new_P1_R2278_U425,
    new_P1_R2278_U426, new_P1_R2278_U427, new_P1_R2278_U428,
    new_P1_R2278_U429, new_P1_R2278_U430, new_P1_R2278_U431,
    new_P1_R2278_U432, new_P1_R2278_U433, new_P1_R2278_U434,
    new_P1_R2278_U435, new_P1_R2278_U436, new_P1_R2278_U437,
    new_P1_R2278_U438, new_P1_R2278_U439, new_P1_R2278_U440,
    new_P1_R2278_U441, new_P1_R2278_U442, new_P1_R2278_U443,
    new_P1_R2278_U444, new_P1_R2278_U445, new_P1_R2278_U446,
    new_P1_R2278_U447, new_P1_R2278_U448, new_P1_R2278_U449,
    new_P1_R2278_U450, new_P1_R2278_U451, new_P1_R2278_U452,
    new_P1_R2278_U453, new_P1_R2278_U454, new_P1_R2278_U455,
    new_P1_R2278_U456, new_P1_R2278_U457, new_P1_R2278_U458,
    new_P1_R2278_U459, new_P1_R2278_U460, new_P1_R2278_U461,
    new_P1_R2278_U462, new_P1_R2278_U463, new_P1_R2278_U464,
    new_P1_R2278_U465, new_P1_R2278_U466, new_P1_R2278_U467,
    new_P1_R2278_U468, new_P1_R2278_U469, new_P1_R2278_U470,
    new_P1_R2278_U471, new_P1_R2278_U472, new_P1_R2278_U473,
    new_P1_R2278_U474, new_P1_R2278_U475, new_P1_R2278_U476,
    new_P1_R2278_U477, new_P1_R2278_U478, new_P1_R2278_U479,
    new_P1_R2278_U480, new_P1_R2278_U481, new_P1_R2278_U482,
    new_P1_R2278_U483, new_P1_R2278_U484, new_P1_R2278_U485,
    new_P1_R2278_U486, new_P1_R2278_U487, new_P1_R2278_U488,
    new_P1_R2278_U489, new_P1_R2278_U490, new_P1_R2278_U491,
    new_P1_R2278_U492, new_P1_R2278_U493, new_P1_R2278_U494,
    new_P1_R2278_U495, new_P1_R2278_U496, new_P1_R2278_U497,
    new_P1_R2278_U498, new_P1_R2278_U499, new_P1_R2278_U500,
    new_P1_R2278_U501, new_P1_R2278_U502, new_P1_R2278_U503,
    new_P1_R2278_U504, new_P1_R2278_U505, new_P1_R2278_U506,
    new_P1_R2278_U507, new_P1_R2278_U508, new_P1_R2278_U509,
    new_P1_R2278_U510, new_P1_R2278_U511, new_P1_R2278_U512,
    new_P1_R2278_U513, new_P1_R2278_U514, new_P1_R2278_U515,
    new_P1_R2278_U516, new_P1_R2278_U517, new_P1_R2278_U518,
    new_P1_R2278_U519, new_P1_R2278_U520, new_P1_R2278_U521,
    new_P1_R2278_U522, new_P1_R2278_U523, new_P1_R2278_U524,
    new_P1_R2278_U525, new_P1_R2278_U526, new_P1_R2278_U527,
    new_P1_R2278_U528, new_P1_R2278_U529, new_P1_R2278_U530,
    new_P1_R2278_U531, new_P1_R2278_U532, new_P1_R2278_U533,
    new_P1_R2278_U534, new_P1_R2278_U535, new_P1_R2278_U536,
    new_P1_R2278_U537, new_P1_R2278_U538, new_P1_R2278_U539,
    new_P1_R2278_U540, new_P1_R2278_U541, new_P1_R2278_U542,
    new_P1_R2278_U543, new_P1_R2278_U544, new_P1_R2278_U545,
    new_P1_R2278_U546, new_P1_R2278_U547, new_P1_R2278_U548,
    new_P1_R2278_U549, new_P1_R2278_U550, new_P1_R2278_U551,
    new_P1_R2278_U552, new_P1_R2278_U553, new_P1_R2278_U554,
    new_P1_R2278_U555, new_P1_R2278_U556, new_P1_R2278_U557,
    new_P1_R2278_U558, new_P1_R2278_U559, new_P1_R2278_U560,
    new_P1_R2278_U561, new_P1_R2278_U562, new_P1_R2278_U563,
    new_P1_R2278_U564, new_P1_R2278_U565, new_P1_R2278_U566,
    new_P1_R2278_U567, new_P1_R2278_U568, new_P1_R2278_U569,
    new_P1_R2278_U570, new_P1_R2278_U571, new_P1_R2278_U572,
    new_P1_R2278_U573, new_P1_R2278_U574, new_P1_R2278_U575,
    new_P1_R2278_U576, new_P1_R2278_U577, new_P1_R2278_U578,
    new_P1_R2278_U579, new_P1_R2278_U580, new_P1_R2278_U581,
    new_P1_R2278_U582, new_P1_R2278_U583, new_P1_R2278_U584,
    new_P1_R2278_U585, new_P1_R2278_U586, new_P1_R2278_U587,
    new_P1_R2278_U588, new_P1_R2278_U589, new_P1_R2278_U590,
    new_P1_R2278_U591, new_P1_R2278_U592, new_P1_R2278_U593,
    new_P1_R2278_U594, new_P1_R2278_U595, new_P1_R2278_U596,
    new_P1_R2278_U597, new_P1_R2278_U598, new_P1_R2278_U599,
    new_P1_R2278_U600, new_P1_R2278_U601, new_P1_R2278_U602,
    new_P1_R2278_U603, new_P1_R2278_U604, new_P1_R2278_U605,
    new_P1_R2278_U606, new_P1_R2278_U607, new_P1_R2278_U608,
    new_P1_R2278_U609, new_P1_R2278_U610, new_P1_R2358_U5, new_P1_R2358_U6,
    new_P1_R2358_U7, new_P1_R2358_U8, new_P1_R2358_U9, new_P1_R2358_U10,
    new_P1_R2358_U11, new_P1_R2358_U12, new_P1_R2358_U13, new_P1_R2358_U14,
    new_P1_R2358_U15, new_P1_R2358_U16, new_P1_R2358_U17, new_P1_R2358_U18,
    new_P1_R2358_U19, new_P1_R2358_U20, new_P1_R2358_U21, new_P1_R2358_U22,
    new_P1_R2358_U23, new_P1_R2358_U24, new_P1_R2358_U25, new_P1_R2358_U26,
    new_P1_R2358_U27, new_P1_R2358_U28, new_P1_R2358_U29, new_P1_R2358_U30,
    new_P1_R2358_U31, new_P1_R2358_U32, new_P1_R2358_U33, new_P1_R2358_U34,
    new_P1_R2358_U35, new_P1_R2358_U36, new_P1_R2358_U37, new_P1_R2358_U38,
    new_P1_R2358_U39, new_P1_R2358_U40, new_P1_R2358_U41, new_P1_R2358_U42,
    new_P1_R2358_U43, new_P1_R2358_U44, new_P1_R2358_U45, new_P1_R2358_U46,
    new_P1_R2358_U47, new_P1_R2358_U48, new_P1_R2358_U49, new_P1_R2358_U50,
    new_P1_R2358_U51, new_P1_R2358_U52, new_P1_R2358_U53, new_P1_R2358_U54,
    new_P1_R2358_U55, new_P1_R2358_U56, new_P1_R2358_U57, new_P1_R2358_U58,
    new_P1_R2358_U59, new_P1_R2358_U60, new_P1_R2358_U61, new_P1_R2358_U62,
    new_P1_R2358_U63, new_P1_R2358_U64, new_P1_R2358_U65, new_P1_R2358_U66,
    new_P1_R2358_U67, new_P1_R2358_U68, new_P1_R2358_U69, new_P1_R2358_U70,
    new_P1_R2358_U71, new_P1_R2358_U72, new_P1_R2358_U73, new_P1_R2358_U74,
    new_P1_R2358_U75, new_P1_R2358_U76, new_P1_R2358_U77, new_P1_R2358_U78,
    new_P1_R2358_U79, new_P1_R2358_U80, new_P1_R2358_U81, new_P1_R2358_U82,
    new_P1_R2358_U83, new_P1_R2358_U84, new_P1_R2358_U85, new_P1_R2358_U86,
    new_P1_R2358_U87, new_P1_R2358_U88, new_P1_R2358_U89, new_P1_R2358_U90,
    new_P1_R2358_U91, new_P1_R2358_U92, new_P1_R2358_U93, new_P1_R2358_U94,
    new_P1_R2358_U95, new_P1_R2358_U96, new_P1_R2358_U97, new_P1_R2358_U98,
    new_P1_R2358_U99, new_P1_R2358_U100, new_P1_R2358_U101,
    new_P1_R2358_U102, new_P1_R2358_U103, new_P1_R2358_U104,
    new_P1_R2358_U105, new_P1_R2358_U106, new_P1_R2358_U107,
    new_P1_R2358_U108, new_P1_R2358_U109, new_P1_R2358_U110,
    new_P1_R2358_U111, new_P1_R2358_U112, new_P1_R2358_U113,
    new_P1_R2358_U114, new_P1_R2358_U115, new_P1_R2358_U116,
    new_P1_R2358_U117, new_P1_R2358_U118, new_P1_R2358_U119,
    new_P1_R2358_U120, new_P1_R2358_U121, new_P1_R2358_U122,
    new_P1_R2358_U123, new_P1_R2358_U124, new_P1_R2358_U125,
    new_P1_R2358_U126, new_P1_R2358_U127, new_P1_R2358_U128,
    new_P1_R2358_U129, new_P1_R2358_U130, new_P1_R2358_U131,
    new_P1_R2358_U132, new_P1_R2358_U133, new_P1_R2358_U134,
    new_P1_R2358_U135, new_P1_R2358_U136, new_P1_R2358_U137,
    new_P1_R2358_U138, new_P1_R2358_U139, new_P1_R2358_U140,
    new_P1_R2358_U141, new_P1_R2358_U142, new_P1_R2358_U143,
    new_P1_R2358_U144, new_P1_R2358_U145, new_P1_R2358_U146,
    new_P1_R2358_U147, new_P1_R2358_U148, new_P1_R2358_U149,
    new_P1_R2358_U150, new_P1_R2358_U151, new_P1_R2358_U152,
    new_P1_R2358_U153, new_P1_R2358_U154, new_P1_R2358_U155,
    new_P1_R2358_U156, new_P1_R2358_U157, new_P1_R2358_U158,
    new_P1_R2358_U159, new_P1_R2358_U160, new_P1_R2358_U161,
    new_P1_R2358_U162, new_P1_R2358_U163, new_P1_R2358_U164,
    new_P1_R2358_U165, new_P1_R2358_U166, new_P1_R2358_U167,
    new_P1_R2358_U168, new_P1_R2358_U169, new_P1_R2358_U170,
    new_P1_R2358_U171, new_P1_R2358_U172, new_P1_R2358_U173,
    new_P1_R2358_U174, new_P1_R2358_U175, new_P1_R2358_U176,
    new_P1_R2358_U177, new_P1_R2358_U178, new_P1_R2358_U179,
    new_P1_R2358_U180, new_P1_R2358_U181, new_P1_R2358_U182,
    new_P1_R2358_U183, new_P1_R2358_U184, new_P1_R2358_U185,
    new_P1_R2358_U186, new_P1_R2358_U187, new_P1_R2358_U188,
    new_P1_R2358_U189, new_P1_R2358_U190, new_P1_R2358_U191,
    new_P1_R2358_U192, new_P1_R2358_U193, new_P1_R2358_U194,
    new_P1_R2358_U195, new_P1_R2358_U196, new_P1_R2358_U197,
    new_P1_R2358_U198, new_P1_R2358_U199, new_P1_R2358_U200,
    new_P1_R2358_U201, new_P1_R2358_U202, new_P1_R2358_U203,
    new_P1_R2358_U204, new_P1_R2358_U205, new_P1_R2358_U206,
    new_P1_R2358_U207, new_P1_R2358_U208, new_P1_R2358_U209,
    new_P1_R2358_U210, new_P1_R2358_U211, new_P1_R2358_U212,
    new_P1_R2358_U213, new_P1_R2358_U214, new_P1_R2358_U215,
    new_P1_R2358_U216, new_P1_R2358_U217, new_P1_R2358_U218,
    new_P1_R2358_U219, new_P1_R2358_U220, new_P1_R2358_U221,
    new_P1_R2358_U222, new_P1_R2358_U223, new_P1_R2358_U224,
    new_P1_R2358_U225, new_P1_R2358_U226, new_P1_R2358_U227,
    new_P1_R2358_U228, new_P1_R2358_U229, new_P1_R2358_U230,
    new_P1_R2358_U231, new_P1_R2358_U232, new_P1_R2358_U233,
    new_P1_R2358_U234, new_P1_R2358_U235, new_P1_R2358_U236,
    new_P1_R2358_U237, new_P1_R2358_U238, new_P1_R2358_U239,
    new_P1_R2358_U240, new_P1_R2358_U241, new_P1_R2358_U242,
    new_P1_R2358_U243, new_P1_R2358_U244, new_P1_R2358_U245,
    new_P1_R2358_U246, new_P1_R2358_U247, new_P1_R2358_U248,
    new_P1_R2358_U249, new_P1_R2358_U250, new_P1_R2358_U251,
    new_P1_R2358_U252, new_P1_R2358_U253, new_P1_R2358_U254,
    new_P1_R2358_U255, new_P1_R2358_U256, new_P1_R2358_U257,
    new_P1_R2358_U258, new_P1_R2358_U259, new_P1_R2358_U260,
    new_P1_R2358_U261, new_P1_R2358_U262, new_P1_R2358_U263,
    new_P1_R2358_U264, new_P1_R2358_U265, new_P1_R2358_U266,
    new_P1_R2358_U267, new_P1_R2358_U268, new_P1_R2358_U269,
    new_P1_R2358_U270, new_P1_R2358_U271, new_P1_R2358_U272,
    new_P1_R2358_U273, new_P1_R2358_U274, new_P1_R2358_U275,
    new_P1_R2358_U276, new_P1_R2358_U277, new_P1_R2358_U278,
    new_P1_R2358_U279, new_P1_R2358_U280, new_P1_R2358_U281,
    new_P1_R2358_U282, new_P1_R2358_U283, new_P1_R2358_U284,
    new_P1_R2358_U285, new_P1_R2358_U286, new_P1_R2358_U287,
    new_P1_R2358_U288, new_P1_R2358_U289, new_P1_R2358_U290,
    new_P1_R2358_U291, new_P1_R2358_U292, new_P1_R2358_U293,
    new_P1_R2358_U294, new_P1_R2358_U295, new_P1_R2358_U296,
    new_P1_R2358_U297, new_P1_R2358_U298, new_P1_R2358_U299,
    new_P1_R2358_U300, new_P1_R2358_U301, new_P1_R2358_U302,
    new_P1_R2358_U303, new_P1_R2358_U304, new_P1_R2358_U305,
    new_P1_R2358_U306, new_P1_R2358_U307, new_P1_R2358_U308,
    new_P1_R2358_U309, new_P1_R2358_U310, new_P1_R2358_U311,
    new_P1_R2358_U312, new_P1_R2358_U313, new_P1_R2358_U314,
    new_P1_R2358_U315, new_P1_R2358_U316, new_P1_R2358_U317,
    new_P1_R2358_U318, new_P1_R2358_U319, new_P1_R2358_U320,
    new_P1_R2358_U321, new_P1_R2358_U322, new_P1_R2358_U323,
    new_P1_R2358_U324, new_P1_R2358_U325, new_P1_R2358_U326,
    new_P1_R2358_U327, new_P1_R2358_U328, new_P1_R2358_U329,
    new_P1_R2358_U330, new_P1_R2358_U331, new_P1_R2358_U332,
    new_P1_R2358_U333, new_P1_R2358_U334, new_P1_R2358_U335,
    new_P1_R2358_U336, new_P1_R2358_U337, new_P1_R2358_U338,
    new_P1_R2358_U339, new_P1_R2358_U340, new_P1_R2358_U341,
    new_P1_R2358_U342, new_P1_R2358_U343, new_P1_R2358_U344,
    new_P1_R2358_U345, new_P1_R2358_U346, new_P1_R2358_U347,
    new_P1_R2358_U348, new_P1_R2358_U349, new_P1_R2358_U350,
    new_P1_R2358_U351, new_P1_R2358_U352, new_P1_R2358_U353,
    new_P1_R2358_U354, new_P1_R2358_U355, new_P1_R2358_U356,
    new_P1_R2358_U357, new_P1_R2358_U358, new_P1_R2358_U359,
    new_P1_R2358_U360, new_P1_R2358_U361, new_P1_R2358_U362,
    new_P1_R2358_U363, new_P1_R2358_U364, new_P1_R2358_U365,
    new_P1_R2358_U366, new_P1_R2358_U367, new_P1_R2358_U368,
    new_P1_R2358_U369, new_P1_R2358_U370, new_P1_R2358_U371,
    new_P1_R2358_U372, new_P1_R2358_U373, new_P1_R2358_U374,
    new_P1_R2358_U375, new_P1_R2358_U376, new_P1_R2358_U377,
    new_P1_R2358_U378, new_P1_R2358_U379, new_P1_R2358_U380,
    new_P1_R2358_U381, new_P1_R2358_U382, new_P1_R2358_U383,
    new_P1_R2358_U384, new_P1_R2358_U385, new_P1_R2358_U386,
    new_P1_R2358_U387, new_P1_R2358_U388, new_P1_R2358_U389,
    new_P1_R2358_U390, new_P1_R2358_U391, new_P1_R2358_U392,
    new_P1_R2358_U393, new_P1_R2358_U394, new_P1_R2358_U395,
    new_P1_R2358_U396, new_P1_R2358_U397, new_P1_R2358_U398,
    new_P1_R2358_U399, new_P1_R2358_U400, new_P1_R2358_U401,
    new_P1_R2358_U402, new_P1_R2358_U403, new_P1_R2358_U404,
    new_P1_R2358_U405, new_P1_R2358_U406, new_P1_R2358_U407,
    new_P1_R2358_U408, new_P1_R2358_U409, new_P1_R2358_U410,
    new_P1_R2358_U411, new_P1_R2358_U412, new_P1_R2358_U413,
    new_P1_R2358_U414, new_P1_R2358_U415, new_P1_R2358_U416,
    new_P1_R2358_U417, new_P1_R2358_U418, new_P1_R2358_U419,
    new_P1_R2358_U420, new_P1_R2358_U421, new_P1_R2358_U422,
    new_P1_R2358_U423, new_P1_R2358_U424, new_P1_R2358_U425,
    new_P1_R2358_U426, new_P1_R2358_U427, new_P1_R2358_U428,
    new_P1_R2358_U429, new_P1_R2358_U430, new_P1_R2358_U431,
    new_P1_R2358_U432, new_P1_R2358_U433, new_P1_R2358_U434,
    new_P1_R2358_U435, new_P1_R2358_U436, new_P1_R2358_U437,
    new_P1_R2358_U438, new_P1_R2358_U439, new_P1_R2358_U440,
    new_P1_R2358_U441, new_P1_R2358_U442, new_P1_R2358_U443,
    new_P1_R2358_U444, new_P1_R2358_U445, new_P1_R2358_U446,
    new_P1_R2358_U447, new_P1_R2358_U448, new_P1_R2358_U449,
    new_P1_R2358_U450, new_P1_R2358_U451, new_P1_R2358_U452,
    new_P1_R2358_U453, new_P1_R2358_U454, new_P1_R2358_U455,
    new_P1_R2358_U456, new_P1_R2358_U457, new_P1_R2358_U458,
    new_P1_R2358_U459, new_P1_R2358_U460, new_P1_R2358_U461,
    new_P1_R2358_U462, new_P1_R2358_U463, new_P1_R2358_U464,
    new_P1_R2358_U465, new_P1_R2358_U466, new_P1_R2358_U467,
    new_P1_R2358_U468, new_P1_R2358_U469, new_P1_R2358_U470,
    new_P1_R2358_U471, new_P1_R2358_U472, new_P1_R2358_U473,
    new_P1_R2358_U474, new_P1_R2358_U475, new_P1_R2358_U476,
    new_P1_R2358_U477, new_P1_R2358_U478, new_P1_R2358_U479,
    new_P1_R2358_U480, new_P1_R2358_U481, new_P1_R2358_U482,
    new_P1_R2358_U483, new_P1_R2358_U484, new_P1_R2358_U485,
    new_P1_R2358_U486, new_P1_R2358_U487, new_P1_R2358_U488,
    new_P1_R2358_U489, new_P1_R2358_U490, new_P1_R2358_U491,
    new_P1_R2358_U492, new_P1_R2358_U493, new_P1_R2358_U494,
    new_P1_R2358_U495, new_P1_R2358_U496, new_P1_R2358_U497,
    new_P1_R2358_U498, new_P1_R2358_U499, new_P1_R2358_U500,
    new_P1_R2358_U501, new_P1_R2358_U502, new_P1_R2358_U503,
    new_P1_R2358_U504, new_P1_R2358_U505, new_P1_R2358_U506,
    new_P1_R2358_U507, new_P1_R2358_U508, new_P1_R2358_U509,
    new_P1_R2358_U510, new_P1_R2358_U511, new_P1_R2358_U512,
    new_P1_R2358_U513, new_P1_R2358_U514, new_P1_R2358_U515,
    new_P1_R2358_U516, new_P1_R2358_U517, new_P1_R2358_U518,
    new_P1_R2358_U519, new_P1_R2358_U520, new_P1_R2358_U521,
    new_P1_R2358_U522, new_P1_R2358_U523, new_P1_R2358_U524,
    new_P1_R2358_U525, new_P1_R2358_U526, new_P1_R2358_U527,
    new_P1_R2358_U528, new_P1_R2358_U529, new_P1_R2358_U530,
    new_P1_R2358_U531, new_P1_R2358_U532, new_P1_R2358_U533,
    new_P1_R2358_U534, new_P1_R2358_U535, new_P1_R2358_U536,
    new_P1_R2358_U537, new_P1_R2358_U538, new_P1_R2358_U539,
    new_P1_R2358_U540, new_P1_R2358_U541, new_P1_R2358_U542,
    new_P1_R2358_U543, new_P1_R2358_U544, new_P1_R2358_U545,
    new_P1_R2358_U546, new_P1_R2358_U547, new_P1_R2358_U548,
    new_P1_R2358_U549, new_P1_R2358_U550, new_P1_R2358_U551,
    new_P1_R2358_U552, new_P1_R2358_U553, new_P1_R2358_U554,
    new_P1_R2358_U555, new_P1_R2358_U556, new_P1_R2358_U557,
    new_P1_R2358_U558, new_P1_R2358_U559, new_P1_R2358_U560,
    new_P1_R2358_U561, new_P1_R2358_U562, new_P1_R2358_U563,
    new_P1_R2358_U564, new_P1_R2358_U565, new_P1_R2358_U566,
    new_P1_R2358_U567, new_P1_R2358_U568, new_P1_R2358_U569,
    new_P1_R2358_U570, new_P1_R2358_U571, new_P1_R2358_U572,
    new_P1_R2358_U573, new_P1_R2358_U574, new_P1_R2358_U575,
    new_P1_R2358_U576, new_P1_R2358_U577, new_P1_R2358_U578,
    new_P1_R2358_U579, new_P1_R2358_U580, new_P1_R2358_U581,
    new_P1_R2358_U582, new_P1_R2358_U583, new_P1_R2358_U584,
    new_P1_R2358_U585, new_P1_R2358_U586, new_P1_R2358_U587,
    new_P1_R2358_U588, new_P1_R2358_U589, new_P1_R2358_U590,
    new_P1_R2358_U591, new_P1_R2358_U592, new_P1_R2358_U593,
    new_P1_R2358_U594, new_P1_R2358_U595, new_P1_R2358_U596,
    new_P1_R2358_U597, new_P1_R2358_U598, new_P1_R2358_U599,
    new_P1_R2358_U600, new_P1_R2358_U601, new_P1_R2358_U602,
    new_P1_R2358_U603, new_P1_R2358_U604, new_P1_R2358_U605,
    new_P1_R2358_U606, new_P1_R2358_U607, new_P1_R2358_U608,
    new_P1_R2358_U609, new_P1_R2358_U610, new_P1_R2358_U611,
    new_P1_LT_589_U6, new_P1_LT_589_U7, new_P1_LT_589_U8, new_P1_R584_U6,
    new_P1_R584_U7, new_P1_R584_U8, new_P1_R584_U9, new_P1_R2099_U4,
    new_P1_R2099_U5, new_P1_R2099_U6, new_P1_R2099_U7, new_P1_R2099_U8,
    new_P1_R2099_U9, new_P1_R2099_U10, new_P1_R2099_U11, new_P1_R2099_U12,
    new_P1_R2099_U13, new_P1_R2099_U14, new_P1_R2099_U15, new_P1_R2099_U16,
    new_P1_R2099_U17, new_P1_R2099_U18, new_P1_R2099_U19, new_P1_R2099_U20,
    new_P1_R2099_U21, new_P1_R2099_U22, new_P1_R2099_U23, new_P1_R2099_U24,
    new_P1_R2099_U25, new_P1_R2099_U26, new_P1_R2099_U27, new_P1_R2099_U28,
    new_P1_R2099_U29, new_P1_R2099_U30, new_P1_R2099_U31, new_P1_R2099_U32,
    new_P1_R2099_U33, new_P1_R2099_U34, new_P1_R2099_U35, new_P1_R2099_U36,
    new_P1_R2099_U37, new_P1_R2099_U38, new_P1_R2099_U39, new_P1_R2099_U40,
    new_P1_R2099_U41, new_P1_R2099_U42, new_P1_R2099_U43, new_P1_R2099_U44,
    new_P1_R2099_U45, new_P1_R2099_U46, new_P1_R2099_U47, new_P1_R2099_U48,
    new_P1_R2099_U49, new_P1_R2099_U50, new_P1_R2099_U51, new_P1_R2099_U52,
    new_P1_R2099_U53, new_P1_R2099_U54, new_P1_R2099_U55, new_P1_R2099_U56,
    new_P1_R2099_U57, new_P1_R2099_U58, new_P1_R2099_U59, new_P1_R2099_U60,
    new_P1_R2099_U61, new_P1_R2099_U62, new_P1_R2099_U63, new_P1_R2099_U64,
    new_P1_R2099_U65, new_P1_R2099_U66, new_P1_R2099_U67, new_P1_R2099_U68,
    new_P1_R2099_U69, new_P1_R2099_U70, new_P1_R2099_U71, new_P1_R2099_U72,
    new_P1_R2099_U73, new_P1_R2099_U74, new_P1_R2099_U75, new_P1_R2099_U76,
    new_P1_R2099_U77, new_P1_R2099_U78, new_P1_R2099_U79, new_P1_R2099_U80,
    new_P1_R2099_U81, new_P1_R2099_U82, new_P1_R2099_U83, new_P1_R2099_U84,
    new_P1_R2099_U85, new_P1_R2099_U86, new_P1_R2099_U87, new_P1_R2099_U88,
    new_P1_R2099_U89, new_P1_R2099_U90, new_P1_R2099_U91, new_P1_R2099_U92,
    new_P1_R2099_U93, new_P1_R2099_U94, new_P1_R2099_U95, new_P1_R2099_U96,
    new_P1_R2099_U97, new_P1_R2099_U98, new_P1_R2099_U99,
    new_P1_R2099_U100, new_P1_R2099_U101, new_P1_R2099_U102,
    new_P1_R2099_U103, new_P1_R2099_U104, new_P1_R2099_U105,
    new_P1_R2099_U106, new_P1_R2099_U107, new_P1_R2099_U108,
    new_P1_R2099_U109, new_P1_R2099_U110, new_P1_R2099_U111,
    new_P1_R2099_U112, new_P1_R2099_U113, new_P1_R2099_U114,
    new_P1_R2099_U115, new_P1_R2099_U116, new_P1_R2099_U117,
    new_P1_R2099_U118, new_P1_R2099_U119, new_P1_R2099_U120,
    new_P1_R2099_U121, new_P1_R2099_U122, new_P1_R2099_U123,
    new_P1_R2099_U124, new_P1_R2099_U125, new_P1_R2099_U126,
    new_P1_R2099_U127, new_P1_R2099_U128, new_P1_R2099_U129,
    new_P1_R2099_U130, new_P1_R2099_U131, new_P1_R2099_U132,
    new_P1_R2099_U133, new_P1_R2099_U134, new_P1_R2099_U135,
    new_P1_R2099_U136, new_P1_R2099_U137, new_P1_R2099_U138,
    new_P1_R2099_U139, new_P1_R2099_U140, new_P1_R2099_U141,
    new_P1_R2099_U142, new_P1_R2099_U143, new_P1_R2099_U144,
    new_P1_R2099_U145, new_P1_R2099_U146, new_P1_R2099_U147,
    new_P1_R2099_U148, new_P1_R2099_U149, new_P1_R2099_U150,
    new_P1_R2099_U151, new_P1_R2099_U152, new_P1_R2099_U153,
    new_P1_R2099_U154, new_P1_R2099_U155, new_P1_R2099_U156,
    new_P1_R2099_U157, new_P1_R2099_U158, new_P1_R2099_U159,
    new_P1_R2099_U160, new_P1_R2099_U161, new_P1_R2099_U162,
    new_P1_R2099_U163, new_P1_R2099_U164, new_P1_R2099_U165,
    new_P1_R2099_U166, new_P1_R2099_U167, new_P1_R2099_U168,
    new_P1_R2099_U169, new_P1_R2099_U170, new_P1_R2099_U171,
    new_P1_R2099_U172, new_P1_R2099_U173, new_P1_R2099_U174,
    new_P1_R2099_U175, new_P1_R2099_U176, new_P1_R2099_U177,
    new_P1_R2099_U178, new_P1_R2099_U179, new_P1_R2099_U180,
    new_P1_R2099_U181, new_P1_R2099_U182, new_P1_R2099_U183,
    new_P1_R2099_U184, new_P1_R2099_U185, new_P1_R2099_U186,
    new_P1_R2099_U187, new_P1_R2099_U188, new_P1_R2099_U189,
    new_P1_R2099_U190, new_P1_R2099_U191, new_P1_R2099_U192,
    new_P1_R2099_U193, new_P1_R2099_U194, new_P1_R2099_U195,
    new_P1_R2099_U196, new_P1_R2099_U197, new_P1_R2099_U198,
    new_P1_R2099_U199, new_P1_R2099_U200, new_P1_R2099_U201,
    new_P1_R2099_U202, new_P1_R2099_U203, new_P1_R2099_U204,
    new_P1_R2099_U205, new_P1_R2099_U206, new_P1_R2099_U207,
    new_P1_R2099_U208, new_P1_R2099_U209, new_P1_R2099_U210,
    new_P1_R2099_U211, new_P1_R2099_U212, new_P1_R2099_U213,
    new_P1_R2099_U214, new_P1_R2099_U215, new_P1_R2099_U216,
    new_P1_R2099_U217, new_P1_R2099_U218, new_P1_R2099_U219,
    new_P1_R2099_U220, new_P1_R2099_U221, new_P1_R2099_U222,
    new_P1_R2099_U223, new_P1_R2099_U224, new_P1_R2099_U225,
    new_P1_R2099_U226, new_P1_R2099_U227, new_P1_R2099_U228,
    new_P1_R2099_U229, new_P1_R2099_U230, new_P1_R2099_U231,
    new_P1_R2099_U232, new_P1_R2099_U233, new_P1_R2099_U234,
    new_P1_R2099_U235, new_P1_R2099_U236, new_P1_R2099_U237,
    new_P1_R2099_U238, new_P1_R2099_U239, new_P1_R2099_U240,
    new_P1_R2099_U241, new_P1_R2099_U242, new_P1_R2099_U243,
    new_P1_R2099_U244, new_P1_R2099_U245, new_P1_R2099_U246,
    new_P1_R2099_U247, new_P1_R2099_U248, new_P1_R2099_U249,
    new_P1_R2099_U250, new_P1_R2099_U251, new_P1_R2099_U252,
    new_P1_R2099_U253, new_P1_R2099_U254, new_P1_R2099_U255,
    new_P1_R2099_U256, new_P1_R2099_U257, new_P1_R2099_U258,
    new_P1_R2099_U259, new_P1_R2099_U260, new_P1_R2099_U261,
    new_P1_R2099_U262, new_P1_R2099_U263, new_P1_R2099_U264,
    new_P1_R2099_U265, new_P1_R2099_U266, new_P1_R2099_U267,
    new_P1_R2099_U268, new_P1_R2099_U269, new_P1_R2099_U270,
    new_P1_R2099_U271, new_P1_R2099_U272, new_P1_R2099_U273,
    new_P1_R2099_U274, new_P1_R2099_U275, new_P1_R2099_U276,
    new_P1_R2099_U277, new_P1_R2099_U278, new_P1_R2099_U279,
    new_P1_R2099_U280, new_P1_R2099_U281, new_P1_R2099_U282,
    new_P1_R2099_U283, new_P1_R2099_U284, new_P1_R2099_U285,
    new_P1_R2099_U286, new_P1_R2099_U287, new_P1_R2099_U288,
    new_P1_R2099_U289, new_P1_R2099_U290, new_P1_R2099_U291,
    new_P1_R2099_U292, new_P1_R2099_U293, new_P1_R2099_U294,
    new_P1_R2099_U295, new_P1_R2099_U296, new_P1_R2099_U297,
    new_P1_R2099_U298, new_P1_R2099_U299, new_P1_R2099_U300,
    new_P1_R2099_U301, new_P1_R2099_U302, new_P1_R2099_U303,
    new_P1_R2099_U304, new_P1_R2099_U305, new_P1_R2099_U306,
    new_P1_R2099_U307, new_P1_R2099_U308, new_P1_R2099_U309,
    new_P1_R2099_U310, new_P1_R2099_U311, new_P1_R2099_U312,
    new_P1_R2099_U313, new_P1_R2099_U314, new_P1_R2099_U315,
    new_P1_R2099_U316, new_P1_R2099_U317, new_P1_R2099_U318,
    new_P1_R2099_U319, new_P1_R2099_U320, new_P1_R2099_U321,
    new_P1_R2099_U322, new_P1_R2099_U323, new_P1_R2099_U324,
    new_P1_R2099_U325, new_P1_R2099_U326, new_P1_R2099_U327,
    new_P1_R2099_U328, new_P1_R2099_U329, new_P1_R2099_U330,
    new_P1_R2099_U331, new_P1_R2099_U332, new_P1_R2099_U333,
    new_P1_R2099_U334, new_P1_R2099_U335, new_P1_R2099_U336,
    new_P1_R2099_U337, new_P1_R2099_U338, new_P1_R2099_U339,
    new_P1_R2099_U340, new_P1_R2099_U341, new_P1_R2099_U342,
    new_P1_R2099_U343, new_P1_R2099_U344, new_P1_R2099_U345,
    new_P1_R2099_U346, new_P1_R2099_U347, new_P1_R2099_U348,
    new_P1_R2099_U349, new_P1_R2167_U6, new_P1_R2167_U7, new_P1_R2167_U8,
    new_P1_R2167_U9, new_P1_R2167_U10, new_P1_R2167_U11, new_P1_R2167_U12,
    new_P1_R2167_U13, new_P1_R2167_U14, new_P1_R2167_U15, new_P1_R2167_U16,
    new_P1_R2167_U17, new_P1_R2167_U18, new_P1_R2167_U19, new_P1_R2167_U20,
    new_P1_R2167_U21, new_P1_R2167_U22, new_P1_R2167_U23, new_P1_R2167_U24,
    new_P1_R2167_U25, new_P1_R2167_U26, new_P1_R2167_U27, new_P1_R2167_U28,
    new_P1_R2167_U29, new_P1_R2167_U30, new_P1_R2167_U31, new_P1_R2167_U32,
    new_P1_R2167_U33, new_P1_R2167_U34, new_P1_R2167_U35, new_P1_R2167_U36,
    new_P1_R2167_U37, new_P1_R2167_U38, new_P1_R2167_U39, new_P1_R2167_U40,
    new_P1_R2167_U41, new_P1_R2167_U42, new_P1_R2167_U43, new_P1_R2167_U44,
    new_P1_R2167_U45, new_P1_R2167_U46, new_P1_R2167_U47, new_P1_R2167_U48,
    new_P1_R2167_U49, new_P1_R2167_U50, new_P1_R2337_U4, new_P1_R2337_U5,
    new_P1_R2337_U6, new_P1_R2337_U7, new_P1_R2337_U8, new_P1_R2337_U9,
    new_P1_R2337_U10, new_P1_R2337_U11, new_P1_R2337_U12, new_P1_R2337_U13,
    new_P1_R2337_U14, new_P1_R2337_U15, new_P1_R2337_U16, new_P1_R2337_U17,
    new_P1_R2337_U18, new_P1_R2337_U19, new_P1_R2337_U20, new_P1_R2337_U21,
    new_P1_R2337_U22, new_P1_R2337_U23, new_P1_R2337_U24, new_P1_R2337_U25,
    new_P1_R2337_U26, new_P1_R2337_U27, new_P1_R2337_U28, new_P1_R2337_U29,
    new_P1_R2337_U30, new_P1_R2337_U31, new_P1_R2337_U32, new_P1_R2337_U33,
    new_P1_R2337_U34, new_P1_R2337_U35, new_P1_R2337_U36, new_P1_R2337_U37,
    new_P1_R2337_U38, new_P1_R2337_U39, new_P1_R2337_U40, new_P1_R2337_U41,
    new_P1_R2337_U42, new_P1_R2337_U43, new_P1_R2337_U44, new_P1_R2337_U45,
    new_P1_R2337_U46, new_P1_R2337_U47, new_P1_R2337_U48, new_P1_R2337_U49,
    new_P1_R2337_U50, new_P1_R2337_U51, new_P1_R2337_U52, new_P1_R2337_U53,
    new_P1_R2337_U54, new_P1_R2337_U55, new_P1_R2337_U56, new_P1_R2337_U57,
    new_P1_R2337_U58, new_P1_R2337_U59, new_P1_R2337_U60, new_P1_R2337_U61,
    new_P1_R2337_U62, new_P1_R2337_U63, new_P1_R2337_U64, new_P1_R2337_U65,
    new_P1_R2337_U66, new_P1_R2337_U67, new_P1_R2337_U68, new_P1_R2337_U69,
    new_P1_R2337_U70, new_P1_R2337_U71, new_P1_R2337_U72, new_P1_R2337_U73,
    new_P1_R2337_U74, new_P1_R2337_U75, new_P1_R2337_U76, new_P1_R2337_U77,
    new_P1_R2337_U78, new_P1_R2337_U79, new_P1_R2337_U80, new_P1_R2337_U81,
    new_P1_R2337_U82, new_P1_R2337_U83, new_P1_R2337_U84, new_P1_R2337_U85,
    new_P1_R2337_U86, new_P1_R2337_U87, new_P1_R2337_U88, new_P1_R2337_U89,
    new_P1_R2337_U90, new_P1_R2337_U91, new_P1_R2337_U92, new_P1_R2337_U93,
    new_P1_R2337_U94, new_P1_R2337_U95, new_P1_R2337_U96, new_P1_R2337_U97,
    new_P1_R2337_U98, new_P1_R2337_U99, new_P1_R2337_U100,
    new_P1_R2337_U101, new_P1_R2337_U102, new_P1_R2337_U103,
    new_P1_R2337_U104, new_P1_R2337_U105, new_P1_R2337_U106,
    new_P1_R2337_U107, new_P1_R2337_U108, new_P1_R2337_U109,
    new_P1_R2337_U110, new_P1_R2337_U111, new_P1_R2337_U112,
    new_P1_R2337_U113, new_P1_R2337_U114, new_P1_R2337_U115,
    new_P1_R2337_U116, new_P1_R2337_U117, new_P1_R2337_U118,
    new_P1_R2337_U119, new_P1_R2337_U120, new_P1_R2337_U121,
    new_P1_R2337_U122, new_P1_R2337_U123, new_P1_R2337_U124,
    new_P1_R2337_U125, new_P1_R2337_U126, new_P1_R2337_U127,
    new_P1_R2337_U128, new_P1_R2337_U129, new_P1_R2337_U130,
    new_P1_R2337_U131, new_P1_R2337_U132, new_P1_R2337_U133,
    new_P1_R2337_U134, new_P1_R2337_U135, new_P1_R2337_U136,
    new_P1_R2337_U137, new_P1_R2337_U138, new_P1_R2337_U139,
    new_P1_R2337_U140, new_P1_R2337_U141, new_P1_R2337_U142,
    new_P1_R2337_U143, new_P1_R2337_U144, new_P1_R2337_U145,
    new_P1_R2337_U146, new_P1_R2337_U147, new_P1_R2337_U148,
    new_P1_R2337_U149, new_P1_R2337_U150, new_P1_R2337_U151,
    new_P1_R2337_U152, new_P1_R2337_U153, new_P1_R2337_U154,
    new_P1_R2337_U155, new_P1_R2337_U156, new_P1_R2337_U157,
    new_P1_R2337_U158, new_P1_R2337_U159, new_P1_R2337_U160,
    new_P1_R2337_U161, new_P1_R2337_U162, new_P1_R2337_U163,
    new_P1_R2337_U164, new_P1_R2337_U165, new_P1_R2337_U166,
    new_P1_R2337_U167, new_P1_R2337_U168, new_P1_R2337_U169,
    new_P1_R2337_U170, new_P1_R2337_U171, new_P1_R2337_U172,
    new_P1_R2337_U173, new_P1_R2337_U174, new_P1_R2337_U175,
    new_P1_R2337_U176, new_P1_R2337_U177, new_P1_R2337_U178,
    new_P1_R2337_U179, new_P1_R2337_U180, new_P1_R2337_U181,
    new_P1_R2337_U182, new_P1_SUB_357_U6, new_P1_SUB_357_U7,
    new_P1_SUB_357_U8, new_P1_SUB_357_U9, new_P1_SUB_357_U10,
    new_P1_SUB_357_U11, new_P1_SUB_357_U12, new_P1_SUB_357_U13,
    new_P1_LT_563_1260_U6, new_P1_LT_563_1260_U7, new_P1_LT_563_1260_U8,
    new_P1_LT_563_1260_U9, new_P1_SUB_580_U6, new_P1_SUB_580_U7,
    new_P1_SUB_580_U8, new_P1_SUB_580_U9, new_P1_SUB_580_U10,
    new_P1_R2096_U4, new_P1_R2096_U5, new_P1_R2096_U6, new_P1_R2096_U7,
    new_P1_R2096_U8, new_P1_R2096_U9, new_P1_R2096_U10, new_P1_R2096_U11,
    new_P1_R2096_U12, new_P1_R2096_U13, new_P1_R2096_U14, new_P1_R2096_U15,
    new_P1_R2096_U16, new_P1_R2096_U17, new_P1_R2096_U18, new_P1_R2096_U19,
    new_P1_R2096_U20, new_P1_R2096_U21, new_P1_R2096_U22, new_P1_R2096_U23,
    new_P1_R2096_U24, new_P1_R2096_U25, new_P1_R2096_U26, new_P1_R2096_U27,
    new_P1_R2096_U28, new_P1_R2096_U29, new_P1_R2096_U30, new_P1_R2096_U31,
    new_P1_R2096_U32, new_P1_R2096_U33, new_P1_R2096_U34, new_P1_R2096_U35,
    new_P1_R2096_U36, new_P1_R2096_U37, new_P1_R2096_U38, new_P1_R2096_U39,
    new_P1_R2096_U40, new_P1_R2096_U41, new_P1_R2096_U42, new_P1_R2096_U43,
    new_P1_R2096_U44, new_P1_R2096_U45, new_P1_R2096_U46, new_P1_R2096_U47,
    new_P1_R2096_U48, new_P1_R2096_U49, new_P1_R2096_U50, new_P1_R2096_U51,
    new_P1_R2096_U52, new_P1_R2096_U53, new_P1_R2096_U54, new_P1_R2096_U55,
    new_P1_R2096_U56, new_P1_R2096_U57, new_P1_R2096_U58, new_P1_R2096_U59,
    new_P1_R2096_U60, new_P1_R2096_U61, new_P1_R2096_U62, new_P1_R2096_U63,
    new_P1_R2096_U64, new_P1_R2096_U65, new_P1_R2096_U66, new_P1_R2096_U67,
    new_P1_R2096_U68, new_P1_R2096_U69, new_P1_R2096_U70, new_P1_R2096_U71,
    new_P1_R2096_U72, new_P1_R2096_U73, new_P1_R2096_U74, new_P1_R2096_U75,
    new_P1_R2096_U76, new_P1_R2096_U77, new_P1_R2096_U78, new_P1_R2096_U79,
    new_P1_R2096_U80, new_P1_R2096_U81, new_P1_R2096_U82, new_P1_R2096_U83,
    new_P1_R2096_U84, new_P1_R2096_U85, new_P1_R2096_U86, new_P1_R2096_U87,
    new_P1_R2096_U88, new_P1_R2096_U89, new_P1_R2096_U90, new_P1_R2096_U91,
    new_P1_R2096_U92, new_P1_R2096_U93, new_P1_R2096_U94, new_P1_R2096_U95,
    new_P1_R2096_U96, new_P1_R2096_U97, new_P1_R2096_U98, new_P1_R2096_U99,
    new_P1_R2096_U100, new_P1_R2096_U101, new_P1_R2096_U102,
    new_P1_R2096_U103, new_P1_R2096_U104, new_P1_R2096_U105,
    new_P1_R2096_U106, new_P1_R2096_U107, new_P1_R2096_U108,
    new_P1_R2096_U109, new_P1_R2096_U110, new_P1_R2096_U111,
    new_P1_R2096_U112, new_P1_R2096_U113, new_P1_R2096_U114,
    new_P1_R2096_U115, new_P1_R2096_U116, new_P1_R2096_U117,
    new_P1_R2096_U118, new_P1_R2096_U119, new_P1_R2096_U120,
    new_P1_R2096_U121, new_P1_R2096_U122, new_P1_R2096_U123,
    new_P1_R2096_U124, new_P1_R2096_U125, new_P1_R2096_U126,
    new_P1_R2096_U127, new_P1_R2096_U128, new_P1_R2096_U129,
    new_P1_R2096_U130, new_P1_R2096_U131, new_P1_R2096_U132,
    new_P1_R2096_U133, new_P1_R2096_U134, new_P1_R2096_U135,
    new_P1_R2096_U136, new_P1_R2096_U137, new_P1_R2096_U138,
    new_P1_R2096_U139, new_P1_R2096_U140, new_P1_R2096_U141,
    new_P1_R2096_U142, new_P1_R2096_U143, new_P1_R2096_U144,
    new_P1_R2096_U145, new_P1_R2096_U146, new_P1_R2096_U147,
    new_P1_R2096_U148, new_P1_R2096_U149, new_P1_R2096_U150,
    new_P1_R2096_U151, new_P1_R2096_U152, new_P1_R2096_U153,
    new_P1_R2096_U154, new_P1_R2096_U155, new_P1_R2096_U156,
    new_P1_R2096_U157, new_P1_R2096_U158, new_P1_R2096_U159,
    new_P1_R2096_U160, new_P1_R2096_U161, new_P1_R2096_U162,
    new_P1_R2096_U163, new_P1_R2096_U164, new_P1_R2096_U165,
    new_P1_R2096_U166, new_P1_R2096_U167, new_P1_R2096_U168,
    new_P1_R2096_U169, new_P1_R2096_U170, new_P1_R2096_U171,
    new_P1_R2096_U172, new_P1_R2096_U173, new_P1_R2096_U174,
    new_P1_R2096_U175, new_P1_R2096_U176, new_P1_R2096_U177,
    new_P1_R2096_U178, new_P1_R2096_U179, new_P1_R2096_U180,
    new_P1_R2096_U181, new_P1_R2096_U182, new_P1_LT_563_U6,
    new_P1_LT_563_U7, new_P1_LT_563_U8, new_P1_LT_563_U9,
    new_P1_LT_563_U10, new_P1_LT_563_U11, new_P1_LT_563_U12,
    new_P1_LT_563_U13, new_P1_LT_563_U14, new_P1_LT_563_U15,
    new_P1_LT_563_U16, new_P1_LT_563_U17, new_P1_LT_563_U18,
    new_P1_LT_563_U19, new_P1_LT_563_U20, new_P1_LT_563_U21,
    new_P1_LT_563_U22, new_P1_LT_563_U23, new_P1_LT_563_U24,
    new_P1_LT_563_U25, new_P1_LT_563_U26, new_P1_LT_563_U27,
    new_P1_LT_563_U28, new_P1_R2238_U6, new_P1_R2238_U7, new_P1_R2238_U8,
    new_P1_R2238_U9, new_P1_R2238_U10, new_P1_R2238_U11, new_P1_R2238_U12,
    new_P1_R2238_U13, new_P1_R2238_U14, new_P1_R2238_U15, new_P1_R2238_U16,
    new_P1_R2238_U17, new_P1_R2238_U18, new_P1_R2238_U19, new_P1_R2238_U20,
    new_P1_R2238_U21, new_P1_R2238_U22, new_P1_R2238_U23, new_P1_R2238_U24,
    new_P1_R2238_U25, new_P1_R2238_U26, new_P1_R2238_U27, new_P1_R2238_U28,
    new_P1_R2238_U29, new_P1_R2238_U30, new_P1_R2238_U31, new_P1_R2238_U32,
    new_P1_R2238_U33, new_P1_R2238_U34, new_P1_R2238_U35, new_P1_R2238_U36,
    new_P1_R2238_U37, new_P1_R2238_U38, new_P1_R2238_U39, new_P1_R2238_U40,
    new_P1_R2238_U41, new_P1_R2238_U42, new_P1_R2238_U43, new_P1_R2238_U44,
    new_P1_R2238_U45, new_P1_R2238_U46, new_P1_R2238_U47, new_P1_R2238_U48,
    new_P1_R2238_U49, new_P1_R2238_U50, new_P1_R2238_U51, new_P1_R2238_U52,
    new_P1_R2238_U53, new_P1_R2238_U54, new_P1_R2238_U55, new_P1_R2238_U56,
    new_P1_R2238_U57, new_P1_R2238_U58, new_P1_R2238_U59, new_P1_R2238_U60,
    new_P1_R2238_U61, new_P1_R2238_U62, new_P1_R2238_U63, new_P1_R2238_U64,
    new_P1_R2238_U65, new_P1_R2238_U66, new_P1_SUB_450_U6,
    new_P1_SUB_450_U7, new_P1_SUB_450_U8, new_P1_SUB_450_U9,
    new_P1_SUB_450_U10, new_P1_SUB_450_U11, new_P1_SUB_450_U12,
    new_P1_SUB_450_U13, new_P1_SUB_450_U14, new_P1_SUB_450_U15,
    new_P1_SUB_450_U16, new_P1_SUB_450_U17, new_P1_SUB_450_U18,
    new_P1_SUB_450_U19, new_P1_SUB_450_U20, new_P1_SUB_450_U21,
    new_P1_SUB_450_U22, new_P1_SUB_450_U23, new_P1_SUB_450_U24,
    new_P1_SUB_450_U25, new_P1_SUB_450_U26, new_P1_SUB_450_U27,
    new_P1_SUB_450_U28, new_P1_SUB_450_U29, new_P1_SUB_450_U30,
    new_P1_SUB_450_U31, new_P1_SUB_450_U32, new_P1_SUB_450_U33,
    new_P1_SUB_450_U34, new_P1_SUB_450_U35, new_P1_SUB_450_U36,
    new_P1_SUB_450_U37, new_P1_SUB_450_U38, new_P1_SUB_450_U39,
    new_P1_SUB_450_U40, new_P1_SUB_450_U41, new_P1_SUB_450_U42,
    new_P1_SUB_450_U43, new_P1_SUB_450_U44, new_P1_SUB_450_U45,
    new_P1_SUB_450_U46, new_P1_SUB_450_U47, new_P1_SUB_450_U48,
    new_P1_SUB_450_U49, new_P1_SUB_450_U50, new_P1_SUB_450_U51,
    new_P1_SUB_450_U52, new_P1_SUB_450_U53, new_P1_SUB_450_U54,
    new_P1_SUB_450_U55, new_P1_SUB_450_U56, new_P1_SUB_450_U57,
    new_P1_SUB_450_U58, new_P1_SUB_450_U59, new_P1_SUB_450_U60,
    new_P1_SUB_450_U61, new_P1_SUB_450_U62, new_P1_SUB_450_U63,
    new_P1_SUB_450_U64, new_P1_SUB_450_U65, new_P1_SUB_450_U66,
    new_P1_ADD_371_U4, new_P1_ADD_371_U5, new_P1_ADD_371_U6,
    new_P1_ADD_371_U7, new_P1_ADD_371_U8, new_P1_ADD_371_U9,
    new_P1_ADD_371_U10, new_P1_ADD_371_U11, new_P1_ADD_371_U12,
    new_P1_ADD_371_U13, new_P1_ADD_371_U14, new_P1_ADD_371_U15,
    new_P1_ADD_371_U16, new_P1_ADD_371_U17, new_P1_ADD_371_U18,
    new_P1_ADD_371_U19, new_P1_ADD_371_U20, new_P1_ADD_371_U21,
    new_P1_ADD_371_U22, new_P1_ADD_371_U23, new_P1_ADD_371_U24,
    new_P1_ADD_371_U25, new_P1_ADD_371_U26, new_P1_ADD_371_U27,
    new_P1_ADD_371_U28, new_P1_ADD_371_U29, new_P1_ADD_371_U30,
    new_P1_ADD_371_U31, new_P1_ADD_371_U32, new_P1_ADD_371_U33,
    new_P1_ADD_371_U34, new_P1_ADD_371_U35, new_P1_ADD_371_U36,
    new_P1_ADD_371_U37, new_P1_ADD_371_U38, new_P1_ADD_371_U39,
    new_P1_ADD_371_U40, new_P1_ADD_371_U41, new_P1_ADD_371_U42,
    new_P1_ADD_371_U43, new_P1_ADD_371_U44, new_P1_ADD_405_U4,
    new_P1_ADD_405_U5, new_P1_ADD_405_U6, new_P1_ADD_405_U7,
    new_P1_ADD_405_U8, new_P1_ADD_405_U9, new_P1_ADD_405_U10,
    new_P1_ADD_405_U11, new_P1_ADD_405_U12, new_P1_ADD_405_U13,
    new_P1_ADD_405_U14, new_P1_ADD_405_U15, new_P1_ADD_405_U16,
    new_P1_ADD_405_U17, new_P1_ADD_405_U18, new_P1_ADD_405_U19,
    new_P1_ADD_405_U20, new_P1_ADD_405_U21, new_P1_ADD_405_U22,
    new_P1_ADD_405_U23, new_P1_ADD_405_U24, new_P1_ADD_405_U25,
    new_P1_ADD_405_U26, new_P1_ADD_405_U27, new_P1_ADD_405_U28,
    new_P1_ADD_405_U29, new_P1_ADD_405_U30, new_P1_ADD_405_U31,
    new_P1_ADD_405_U32, new_P1_ADD_405_U33, new_P1_ADD_405_U34,
    new_P1_ADD_405_U35, new_P1_ADD_405_U36, new_P1_ADD_405_U37,
    new_P1_ADD_405_U38, new_P1_ADD_405_U39, new_P1_ADD_405_U40,
    new_P1_ADD_405_U41, new_P1_ADD_405_U42, new_P1_ADD_405_U43,
    new_P1_ADD_405_U44, new_P1_ADD_405_U45, new_P1_ADD_405_U46,
    new_P1_ADD_405_U47, new_P1_ADD_405_U48, new_P1_ADD_405_U49,
    new_P1_ADD_405_U50, new_P1_ADD_405_U51, new_P1_ADD_405_U52,
    new_P1_ADD_405_U53, new_P1_ADD_405_U54, new_P1_ADD_405_U55,
    new_P1_ADD_405_U56, new_P1_ADD_405_U57, new_P1_ADD_405_U58,
    new_P1_ADD_405_U59, new_P1_ADD_405_U60, new_P1_ADD_405_U61,
    new_P1_ADD_405_U62, new_P1_ADD_405_U63, new_P1_ADD_405_U64,
    new_P1_ADD_405_U65, new_P1_ADD_405_U66, new_P1_ADD_405_U67,
    new_P1_ADD_405_U68, new_P1_ADD_405_U69, new_P1_ADD_405_U70,
    new_P1_ADD_405_U71, new_P1_ADD_405_U72, new_P1_ADD_405_U73,
    new_P1_ADD_405_U74, new_P1_ADD_405_U75, new_P1_ADD_405_U76,
    new_P1_ADD_405_U77, new_P1_ADD_405_U78, new_P1_ADD_405_U79,
    new_P1_ADD_405_U80, new_P1_ADD_405_U81, new_P1_ADD_405_U82,
    new_P1_ADD_405_U83, new_P1_ADD_405_U84, new_P1_ADD_405_U85,
    new_P1_ADD_405_U86, new_not_keyinput0, new_not_keyinput1,
    new_not_keyinput2, new_not_keyinput3, new_not_keyinput4, new_not_0,
    new_and_1, new_not_2, new_and_3, new_not_4, new_and_5, new_not_6,
    new_and_7, new_not_9, new_and_10, new_not_11, new_and_12, new_not_13,
    new_and_14, new_not_16, new_and_17, new_not_18, new_and_19,
    new_not_Q_0, new_not_Q_1, new_not_Q_2, new_not_Q_3, new_count_state_1,
    new_count_state_2, new_count_state_3, new_count_state_4,
    new_count_state_5, new_count_state_6, new_count_state_7,
    new_count_state_8, new_count_state_9, new_count_state_10,
    new_count_state_11, new_count_state_12, new_count_state_13,
    new_count_state_14, new_count_state_15, new_y_mux_key0_and_0,
    new_y_mux_key0_and_1, new_y_mux_key0, new_y_mux_key1_and_0,
    new_y_mux_key1_and_1, new_y_mux_key1, new_y_mux_key2_and_0,
    new_y_mux_key2_and_1, new_y_mux_key2, new_y_mux_key3_and_0,
    new_y_mux_key3_and_1, new_y_mux_key3, new_y_mux_key4_and_0,
    new_y_mux_key4_and_1, new_y_mux_key4, new_y_mux_key5_and_0,
    new_y_mux_key5_and_1, new_y_mux_key5, new_y_mux_key6_and_0,
    new_y_mux_key6_and_1, new_y_mux_key6, new_y_mux_key7_and_0,
    new_y_mux_key7_and_1, new_y_mux_key7, new_y_mux_key8_and_0,
    new_y_mux_key8_and_1, new_y_mux_key8, new_y_mux_key9_and_0,
    new_y_mux_key9_and_1, new_y_mux_key9, new_y_mux_key10_and_0,
    new_y_mux_key10_and_1, new_y_mux_key10, new_y_mux_key11_and_0,
    new_y_mux_key11_and_1, new_y_mux_key11, new_y_mux_key12_and_0,
    new_y_mux_key12_and_1, new_y_mux_key12, new_y_mux_key13_and_0,
    new_y_mux_key13_and_1, new_y_mux_key13, new_y_mux_key14_and_0,
    new_y_mux_key14_and_1, new_y_mux_key14, new_y_mux_key15_and_0,
    new_y_mux_key15_and_1, new_y_mux_key15, new__state_1, new__state_2,
    new__state_3, new__state_4, new__state_5, new__state_6, new__state_7,
    new__state_8, new__state_9, new__state_10, new__state_11,
    new__state_12, new__state_13, new__state_14, new__state_15,
    new__state_17, new__state_18, new__state_19, new__state_20,
    new__state_21, new__state_22, new__state_23, new__state_25,
    new__state_26, new__state_27, new__state_29, new_s__state_1,
    new_not_s__state_1, new_I0__state_1, new_I1__state_1,
    new_and_mux__state_1, new_and_mux__state_1_2, new_y_mux_16,
    new_s__state_3, new_not_s__state_3, new_I0__state_3, new_I1__state_3,
    new_and_mux__state_3, new_and_mux__state_3_2, new_y_mux_17,
    new_s__state_5, new_not_s__state_5, new_I0__state_5, new_I1__state_5,
    new_and_mux__state_5, new_and_mux__state_5_2, new_y_mux_18,
    new_s__state_7, new_not_s__state_7, new_I0__state_7, new_I1__state_7,
    new_and_mux__state_7, new_and_mux__state_7_2, new_y_mux_19,
    new_s__state_9, new_not_s__state_9, new_I0__state_9, new_I1__state_9,
    new_and_mux__state_9, new_and_mux__state_9_2, new_y_mux_20,
    new_s__state_11, new_not_s__state_11, new_I0__state_11,
    new_I1__state_11, new_and_mux__state_11, new_and_mux__state_11_2,
    new_y_mux_21, new_s__state_13, new_not_s__state_13, new_I0__state_13,
    new_I1__state_13, new_and_mux__state_13, new_and_mux__state_13_2,
    new_y_mux_22, new_s__state_15, new_not_s__state_15, new_I0__state_15,
    new_I1__state_15, new_and_mux__state_15, new_and_mux__state_15_2,
    new_y_mux_23, new_s__state_17, new_not_s__state_17, new_I0__state_17,
    new_I1__state_17, new_and_mux__state_17, new_and_mux__state_17_2,
    new_y_mux_24, new_s__state_19, new_not_s__state_19, new_I0__state_19,
    new_I1__state_19, new_and_mux__state_19, new_and_mux__state_19_2,
    new_y_mux_25, new_s__state_21, new_not_s__state_21, new_I0__state_21,
    new_I1__state_21, new_and_mux__state_21, new_and_mux__state_21_2,
    new_y_mux_26, new_s__state_23, new_not_s__state_23, new_I0__state_23,
    new_I1__state_23, new_and_mux__state_23, new_and_mux__state_23_2,
    new_y_mux_27, new_s__state_25, new_not_s__state_25, new_I0__state_25,
    new_I1__state_25, new_and_mux__state_25, new_and_mux__state_25_2,
    new_y_mux_28, new_s__state_27, new_not_s__state_27, new_I0__state_27,
    new_I1__state_27, new_and_mux__state_27, new_and_mux__state_27_2,
    new_y_mux_29, new_s__state_29, new_not_s__state_29, new_I0__state_29,
    new_I1__state_29, new_and_mux__state_29, new_and_mux__state_29_2, n280,
    n285, n290, n295, n300, n305, n310, n315, n320, n325, n330, n335, n340,
    n345, n350, n355, n360, n365, n370, n375, n380, n385, n390, n395, n400,
    n405, n410, n415, n420, n425, n430, n435, n440, n445, n450, n455, n460,
    n465, n470, n475, n480, n485, n490, n495, n500, n505, n510, n515, n520,
    n525, n530, n535, n540, n545, n550, n555, n560, n565, n570, n575, n580,
    n585, n590, n595, n600, n605, n610, n615, n620, n625, n630, n635, n640,
    n645, n650, n655, n660, n665, n670, n675, n680, n685, n690, n695, n700,
    n705, n710, n715, n720, n725, n730, n735, n740, n745, n750, n755, n760,
    n765, n770, n775, n780, n785, n790, n795, n800, n805, n810, n815, n820,
    n825, n830, n835, n840, n845, n850, n855, n860, n865, n870, n875, n880,
    n885, n890, n895, n900, n905, n910, n915, n920, n925, n930, n935, n940,
    n945, n950, n955, n960, n965, n970, n975, n980, n985, n990, n995,
    n1000, n1005, n1010, n1015, n1020, n1025, n1030, n1035, n1040, n1045,
    n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085, n1090, n1095,
    n1100, n1105, n1110, n1115, n1120, n1125, n1130, n1135, n1140, n1145,
    n1150, n1155, n1160, n1165, n1170, n1175, n1180, n1185, n1190, n1195,
    n1200, n1205, n1210, n1215, n1220, n1225, n1230, n1235, n1240, n1245,
    n1250, n1255, n1260, n1265, n1270, n1275, n1280, n1285, n1290, n1295,
    n1300, n1305, n1310, n1315, n1320, n1325, n1330, n1335, n1340, n1345,
    n1350, n1355, n1360, n1365, n1370, n1375, n1380, n1385, n1390, n1395,
    n1400, n1405, n1410, n1415, n1420, n1425, n1430, n1435, n1440, n1445,
    n1450, n1455, n1460, n1465, n1470, n1475, n1480, n1485, n1490, n1495,
    n1500, n1505, n1510, n1515, n1520, n1525, n1530, n1535, n1540, n1545,
    n1550, n1555, n1560, n1565, n1570, n1575, n1580, n1585, n1590, n1595,
    n1600, n1605, n1610, n1615, n1620, n1625, n1630, n1635, n1640, n1645,
    n1650, n1655, n1660, n1665, n1670, n1675, n1680, n1685, n1690, n1695,
    n1700, n1705, n1710, n1715, n1720, n1725, n1730, n1735, n1740, n1745,
    n1750, n1755, n1760, n1765, n1770, n1775, n1780, n1785, n1790, n1795,
    n1800, n1805, n1810, n1815, n1820, n1825, n1830, n1835, n1840, n1845,
    n1850, n1855, n1860, n1865, n1870, n1875, n1880, n1885, n1890, n1895,
    n1900, n1905, n1910, n1915, n1920, n1925, n1930, n1935, n1940, n1945,
    n1950, n1955, n1960, n1965, n1970, n1975, n1980, n1985, n1990, n1995,
    n2000, n2005, n2010, n2015, n2020, n2025, n2030, n2035, n2040, n2045,
    n2050, n2055, n2060, n2065, n2070, n2075, n2080, n2085, n2090, n2095,
    n2100, n2105, n2110, n2115, n2120, n2125, n2130, n2135, n2140, n2145,
    n2150, n2154, n2158, n2162, n2166, n2170, n2174, n2178, n2182, n2186,
    n2190, n2194, n2198, n2202, n2206, n2210, n2214, n2218, n2222, n2226,
    n2230, n2234, n2238, n2242, n2246, n2250, n2254, n2258, n2262, n2266,
    n2270, n2274, n2278, n2283, n2288, n2293, n2298, n2303, n2308, n2313,
    n2318, n2323, n2328, n2333, n2338, n2343, n2348, n2353, n2358, n2363,
    n2368, n2373, n2378, n2383, n2388, n2393, n2398, n2403, n2408, n2413,
    n2418, n2423, n2428, n2433, n2438, n2443, n2448, n2453, n2458, n2463,
    n2468, n2473, n2478, n2483, n2488, n2493, n2498, n2503, n2508, n2513,
    n2518, n2523, n2528, n2533, n2538, n2543, n2548, n2553, n2558, n2563,
    n2568, n2573, n2578, n2583, n2588, n2593, n2598, n2603, n2608, n2613,
    n2618, n2623, n2628, n2633, n2638, n2643, n2648, n2653, n2658, n2663,
    n2668, n2673, n2678, n2683, n2688, n2693, n2698, n2703, n2708, n2713,
    n2718, n2723, n2728, n2733, n2738, n2743, n2748, n2753, n2758, n2763,
    n2768, n2773, n2778, n2782, n2787, n2792, n2797, n2802, n2806, n2810,
    n2815, n2819, n2824, n2829, n2834, n2839, n2844, n2849, n2854, n2859,
    n2864, n2869, n2874, n2879, n2884, n2889, n2894, n2899, n2904, n2909,
    n2914, n2919, n2924, n2929, n2934, n2939, n2944, n2949, n2954, n2959,
    n2964, n2969, n2974, n2979, n2984, n2989, n2994, n2999, n3004, n3009,
    n3014, n3019, n3024, n3029, n3034, n3039, n3044, n3049, n3054, n3059,
    n3064, n3069, n3074, n3079, n3084, n3089, n3094, n3099, n3104, n3109,
    n3114, n3119, n3124, n3129, n3134, n3139, n3144, n3149, n3154, n3159,
    n3164, n3169, n3174, n3179, n3184, n3189, n3194, n3199, n3204, n3209,
    n3214, n3219, n3224, n3229, n3234, n3239, n3244, n3249, n3254, n3259,
    n3264, n3269, n3274, n3279, n3284, n3289, n3294, n3299, n3304, n3309,
    n3314, n3319, n3324, n3329, n3334, n3339, n3344, n3349, n3354, n3359,
    n3364, n3369, n3374, n3379, n3384, n3389, n3394, n3399, n3404, n3409,
    n3414, n3419, n3424, n3429, n3434, n3439, n3444, n3449, n3454, n3459,
    n3464, n3469, n3474, n3479, n3484, n3489, n3494, n3499, n3504, n3509,
    n3514, n3519, n3524, n3529, n3534, n3539, n3544, n3549, n3554, n3559,
    n3564, n3569, n3574, n3579, n3584, n3589, n3594, n3599, n3604, n3609,
    n3614, n3619, n3624, n3629, n3634, n3639, n3644, n3649, n3654, n3659,
    n3664, n3669, n3674, n3679, n3684, n3689, n3694, n3699, n3704, n3709,
    n3714, n3719, n3724, n3729, n3734, n3739, n3744, n3749, n3754, n3759,
    n3764, n3769, n3774, n3779, n3784, n3789, n3794, n3799, n3804, n3809,
    n3814, n3819, n3824, n3829, n3834, n3839, n3844, n3849, n3854, n3859,
    n3864, n3869, n3874, n3879, n3884, n3889, n3894, n3899, n3904, n3909,
    n3914, n3919, n3924, n3929, n3934, n3939, n3944, n3949, n3954, n3959,
    n3964, n3969, n3974, n3979, n3984, n3989, n3994, n3999, n4004, n4009,
    n4014, n4019, n4024, n4029, n4034, n4039, n4044, n4049, n4054, n4059,
    n4064, n4069, n4074, n4079, n4084, n4089, n4094, n4099, n4104, n4109,
    n4114, n4119, n4124, n4129, n4134, n4139, n4144, n4149, n4154, n4159,
    n4164, n4169, n4174, n4179, n4184, n4189, n4194, n4199, n4204, n4209,
    n4214, n4219, n4224, n4229, n4234, n4239, n4244, n4249, n4254, n4259,
    n4264, n4269, n4274, n4279, n4284, n4289, n4294, n4299, n4304, n4309,
    n4314, n4319, n4324, n4329, n4334, n4339, n4344, n4349, n4354, n4359,
    n4364, n4369, n4374, n4379, n4384, n4389, n4394, n4399, n4404, n4409,
    n4414, n4419, n4424, n4429, n4434, n4439, n4444, n4449, n4454, n4459,
    n4464, n4469, n4474, n4479, n4484, n4489, n4494, n4499, n4504, n4509,
    n4514, n4519, n4524, n4529, n4534, n4539, n4544, n4549, n4554, n4559,
    n4564, n4569, n4574, n4579, n4584, n4589, n4594, n4599, n4604, n4609,
    n4614, n4619, n4624, n4629, n4634, n4639, n4644, n4649, n4654, n4659,
    n4664, n4669, n4674, n4679, n4684, n4689, n4694, n4699, n4704, n4709,
    n4714, n4719, n4724, n4729, n4734, n4739, n4744, n4749, n4754, n4759,
    n4764, n4769, n4774, n4779, n4784, n4789, n4794, n4799, n4804, n4809,
    n4814, n4819, n4824, n4829, n4834, n4839, n4844, n4849, n4854, n4859,
    n4864, n4869, n4874, n4879, n4884, n4889, n4894, n4899, n4904, n4909,
    n4914, n4919, n4924, n4929, n4934, n4939, n4944, n4949, n4954, n4959,
    n4964, n4969, n4974, n4979, n4984, n4989, n4994, n4999, n5004, n5009,
    n5014, n5019, n5024, n5029, n5034, n5039, n5044, n5049, n5054, n5059,
    n5064, n5069, n5074, n5079, n5084, n5089, n5094, n5098, n5102, n5106,
    n5110, n5114, n5118, n5122, n5126, n5130, n5134, n5138, n5142, n5146,
    n5150, n5154, n5158, n5162, n5166, n5170, n5174, n5178, n5182, n5186,
    n5190, n5194, n5198, n5202, n5206, n5210, n5214, n5219, n5224, n5229,
    n5234, n5239, n5244, n5249, n5254, n5259, n5264, n5269, n5274, n5279,
    n5284, n5289, n5294, n5299, n5304, n5309, n5314, n5319, n5324, n5329,
    n5334, n5339, n5344, n5349, n5354, n5359, n5364, n5369, n5374, n5379,
    n5384, n5389, n5394, n5399, n5404, n5409, n5414, n5419, n5424, n5429,
    n5434, n5439, n5444, n5449, n5454, n5459, n5464, n5469, n5474, n5479,
    n5484, n5489, n5494, n5499, n5504, n5509, n5514, n5519, n5524, n5529,
    n5534, n5539, n5544, n5549, n5554, n5559, n5564, n5569, n5574, n5579,
    n5584, n5589, n5594, n5599, n5604, n5609, n5614, n5619, n5624, n5629,
    n5634, n5639, n5644, n5649, n5654, n5659, n5664, n5669, n5674, n5679,
    n5684, n5689, n5694, n5699, n5704, n5709, n5714, n5719, n5724, n5729,
    n5734, n5739, n5744, n5749, n5754, n5759, n5764, n5769, n5774, n5779,
    n5784, n5789, n5794, n5799, n5804, n5809, n5814, n5819, n5824, n5829,
    n5834, n5839, n5844, n5849, n5854, n5859, n5864, n5869, n5874, n5879,
    n5884, n5889, n5894, n5899, n5904, n5909, n5914, n5919, n5924, n5929,
    n5934, n5939, n5944, n5949, n5954, n5959, n5964, n5969, n5974, n5979,
    n5984, n5989, n5994, n5999, n6004, n6009, n6014, n6019, n6024, n6029,
    n6034, n6039, n6044, n6049, n6054, n6059, n6064, n6069, n6074, n6079,
    n6084, n6089, n6094, n6099, n6104, n6109, n6114, n6119, n6124, n6129,
    n6134, n6139, n6144, n6149, n6154, n6159, n6164, n6169, n6174, n6179,
    n6184, n6189, n6194, n6199, n6204, n6209, n6214, n6219, n6224, n6229,
    n6234, n6239, n6244, n6249, n6254, n6259, n6264, n6269, n6274, n6279,
    n6284, n6289, n6294, n6299, n6304, n6309, n6314, n6319, n6324, n6329,
    n6334, n6339, n6344, n6349, n6354, n6359, n6364, n6369, n6374, n6379,
    n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429,
    n6434, n6439, n6444, n6449, n6454, n6459, n6464, n6469, n6474, n6479,
    n6484, n6489, n6494, n6499, n6504, n6509, n6514, n6519, n6524, n6529,
    n6534, n6539, n6544, n6549, n6554, n6559, n6564, n6569, n6574, n6579,
    n6584, n6589, n6594, n6599, n6604, n6609, n6614, n6619, n6624, n6629,
    n6634, n6639, n6644, n6649, n6654, n6659, n6664, n6669, n6674, n6679,
    n6684, n6689, n6694, n6699, n6704, n6709, n6714, n6719, n6724, n6729,
    n6734, n6739, n6744, n6749, n6754, n6759, n6764, n6769, n6774, n6779,
    n6784, n6789, n6794, n6799, n6804, n6809, n6814, n6819, n6824, n6829,
    n6834, n6839, n6844, n6849, n6854, n6859, n6864, n6869, n6874, n6879,
    n6884, n6889, n6894, n6899, n6904, n6909, n6914, n6919, n6924, n6929,
    n6934, n6939, n6944, n6949, n6954, n6959, n6964, n6969, n6974, n6979,
    n6984, n6989, n6994, n6999, n7004, n7009, n7014, n7019, n7024, n7029,
    n7034, n7039, n7044, n7049, n7054, n7059, n7064, n7069, n7074, n7079,
    n7084, n7089, n7094, n7099, n7104, n7109, n7114, n7119, n7124, n7129,
    n7134, n7139, n7144, n7149, n7154, n7159, n7164, n7169, n7174, n7179,
    n7184, n7189, n7194, n7199, n7204, n7209, n7214, n7219, n7224, n7229,
    n7234, n7239, n7244, n7249, n7254, n7259, n7264, n7269, n7274, n7278,
    n7283, n67455, n67458, n67461, n67464;
  assign new_P1_ADD_515_U182 = ~new_P1_ADD_515_U107 | ~new_P1_ADD_515_U33;
  assign new_P1_ADD_515_U181 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_ADD_515_U32;
  assign new_P1_ADD_515_U180 = ~new_P1_ADD_515_U116 | ~new_P1_ADD_515_U51;
  assign new_U207 = new_U250 & n615;
  assign new_U208 = new_U377 & new_U378 & P2_W_R_N_REG & P2_M_IO_N_REG;
  assign new_U209 = READY22_REG & READY2;
  assign new_U210 = READY11_REG & READY1;
  assign new_U211 = READY12_REG & READY21_REG;
  assign n600 = ~n615 | ~new_U208 | ~new_R170_U6;
  assign n610 = ~n605 | ~new_U379 | ~P3_M_IO_N_REG | ~new_U380;
  assign n615 = ~new_R165_U6 | ~new_U381 | ~P1_W_R_N_REG | ~P1_M_IO_N_REG | ~new_U383;
  assign n605 = ~new_LT_748_U6 | ~new_U208;
  assign n435 = ~new_U482 | ~new_U483 | ~new_U484;
  assign n430 = ~new_U479 | ~new_U480 | ~new_U481;
  assign n425 = ~new_U476 | ~new_U477 | ~new_U478;
  assign n420 = ~new_U473 | ~new_U474 | ~new_U475;
  assign n415 = ~new_U470 | ~new_U471 | ~new_U472;
  assign n410 = ~new_U467 | ~new_U468 | ~new_U469;
  assign n405 = ~new_U464 | ~new_U465 | ~new_U466;
  assign n400 = ~new_U461 | ~new_U462 | ~new_U463;
  assign n395 = ~new_U458 | ~new_U459 | ~new_U460;
  assign n390 = ~new_U455 | ~new_U456 | ~new_U457;
  assign n385 = ~new_U452 | ~new_U453 | ~new_U454;
  assign n380 = ~new_U449 | ~new_U450 | ~new_U451;
  assign n375 = ~new_U446 | ~new_U447 | ~new_U448;
  assign n370 = ~new_U443 | ~new_U444 | ~new_U445;
  assign n365 = ~new_U440 | ~new_U441 | ~new_U442;
  assign n360 = ~new_U437 | ~new_U438 | ~new_U439;
  assign n355 = ~new_U434 | ~new_U435 | ~new_U436;
  assign n350 = ~new_U431 | ~new_U432 | ~new_U433;
  assign n345 = ~new_U428 | ~new_U429 | ~new_U430;
  assign n340 = ~new_U425 | ~new_U426 | ~new_U427;
  assign n335 = ~new_U422 | ~new_U423 | ~new_U424;
  assign n330 = ~new_U419 | ~new_U420 | ~new_U421;
  assign n325 = ~new_U416 | ~new_U417 | ~new_U418;
  assign n320 = ~new_U413 | ~new_U414 | ~new_U415;
  assign n315 = ~new_U410 | ~new_U411 | ~new_U412;
  assign n310 = ~new_U407 | ~new_U408 | ~new_U409;
  assign n305 = ~new_U404 | ~new_U405 | ~new_U406;
  assign n300 = ~new_U401 | ~new_U402 | ~new_U403;
  assign n295 = ~new_U398 | ~new_U399 | ~new_U400;
  assign n290 = ~new_U395 | ~new_U396 | ~new_U397;
  assign n285 = ~new_U392 | ~new_U393 | ~new_U394;
  assign new_U247 = ~new_U389 | ~new_U390 | ~new_U391;
  assign new_U248 = ~new_R165_U6;
  assign new_U249 = ~new_R170_U6;
  assign new_U250 = ~n615 | ~new_U387;
  assign n440 = ~new_U486 | ~new_U485;
  assign n445 = ~new_U488 | ~new_U487;
  assign n450 = ~new_U490 | ~new_U489;
  assign n455 = ~new_U492 | ~new_U491;
  assign n460 = ~new_U494 | ~new_U493;
  assign n465 = ~new_U496 | ~new_U495;
  assign n470 = ~new_U498 | ~new_U497;
  assign n475 = ~new_U500 | ~new_U499;
  assign n480 = ~new_U502 | ~new_U501;
  assign n485 = ~new_U504 | ~new_U503;
  assign n490 = ~new_U506 | ~new_U505;
  assign n495 = ~new_U508 | ~new_U507;
  assign n500 = ~new_U510 | ~new_U509;
  assign n505 = ~new_U512 | ~new_U511;
  assign n510 = ~new_U514 | ~new_U513;
  assign n515 = ~new_U516 | ~new_U515;
  assign n520 = ~new_U518 | ~new_U517;
  assign n525 = ~new_U520 | ~new_U519;
  assign n530 = ~new_U522 | ~new_U521;
  assign n535 = ~new_U524 | ~new_U523;
  assign n540 = ~new_U526 | ~new_U525;
  assign n545 = ~new_U528 | ~new_U527;
  assign n550 = ~new_U530 | ~new_U529;
  assign n555 = ~new_U532 | ~new_U531;
  assign n560 = ~new_U534 | ~new_U533;
  assign n565 = ~new_U536 | ~new_U535;
  assign n570 = ~new_U538 | ~new_U537;
  assign n575 = ~new_U540 | ~new_U539;
  assign n580 = ~new_U542 | ~new_U541;
  assign n585 = ~new_U544 | ~new_U543;
  assign n590 = ~new_U546 | ~new_U545;
  assign n595 = ~new_U548 | ~new_U547;
  assign new_U283 = ~new_U550 | ~new_U549;
  assign new_U284 = ~new_U552 | ~new_U551;
  assign new_U285 = ~new_U554 | ~new_U553;
  assign new_U286 = ~new_U556 | ~new_U555;
  assign new_U287 = ~new_U558 | ~new_U557;
  assign new_U288 = ~new_U560 | ~new_U559;
  assign new_U289 = ~new_U562 | ~new_U561;
  assign new_U290 = ~new_U564 | ~new_U563;
  assign new_U291 = ~new_U566 | ~new_U565;
  assign new_U292 = ~new_U568 | ~new_U567;
  assign new_U293 = ~new_U570 | ~new_U569;
  assign new_U294 = ~new_U572 | ~new_U571;
  assign new_U295 = ~new_U574 | ~new_U573;
  assign new_U296 = ~new_U576 | ~new_U575;
  assign new_U297 = ~new_U578 | ~new_U577;
  assign new_U298 = ~new_U580 | ~new_U579;
  assign new_U299 = ~new_U582 | ~new_U581;
  assign new_U300 = ~new_U584 | ~new_U583;
  assign new_U301 = ~new_U586 | ~new_U585;
  assign new_U302 = ~new_U588 | ~new_U587;
  assign new_U303 = ~new_U590 | ~new_U589;
  assign new_U304 = ~new_U592 | ~new_U591;
  assign new_U305 = ~new_U594 | ~new_U593;
  assign new_U306 = ~new_U596 | ~new_U595;
  assign new_U307 = ~new_U598 | ~new_U597;
  assign new_U308 = ~new_U600 | ~new_U599;
  assign new_U309 = ~new_U602 | ~new_U601;
  assign new_U310 = ~new_U604 | ~new_U603;
  assign new_U311 = ~new_U606 | ~new_U605;
  assign new_U312 = ~new_U608 | ~new_U607;
  assign new_U313 = ~new_U610 | ~new_U609;
  assign new_U314 = ~new_U612 | ~new_U611;
  assign new_U315 = ~new_U614 | ~new_U613;
  assign new_U316 = ~new_U616 | ~new_U615;
  assign new_U317 = ~new_U618 | ~new_U617;
  assign new_U318 = ~new_U620 | ~new_U619;
  assign new_U319 = ~new_U622 | ~new_U621;
  assign new_U320 = ~new_U624 | ~new_U623;
  assign new_U321 = ~new_U626 | ~new_U625;
  assign new_U322 = ~new_U628 | ~new_U627;
  assign new_U323 = ~new_U630 | ~new_U629;
  assign new_U324 = ~new_U632 | ~new_U631;
  assign new_U325 = ~new_U634 | ~new_U633;
  assign new_U326 = ~new_U636 | ~new_U635;
  assign new_U327 = ~new_U638 | ~new_U637;
  assign new_U328 = ~new_U640 | ~new_U639;
  assign new_U329 = ~new_U642 | ~new_U641;
  assign new_U330 = ~new_U644 | ~new_U643;
  assign new_U331 = ~new_U646 | ~new_U645;
  assign new_U332 = ~new_U648 | ~new_U647;
  assign new_U333 = ~new_U650 | ~new_U649;
  assign new_U334 = ~new_U652 | ~new_U651;
  assign new_U335 = ~new_U654 | ~new_U653;
  assign new_U336 = ~new_U656 | ~new_U655;
  assign new_U337 = ~new_U658 | ~new_U657;
  assign new_U338 = ~new_U660 | ~new_U659;
  assign new_U339 = ~new_U662 | ~new_U661;
  assign new_U340 = ~new_U664 | ~new_U663;
  assign new_U341 = ~new_U666 | ~new_U665;
  assign new_U342 = ~new_U668 | ~new_U667;
  assign new_U343 = ~new_U670 | ~new_U669;
  assign new_U344 = ~new_U672 | ~new_U671;
  assign new_U345 = ~new_U674 | ~new_U673;
  assign new_U346 = ~new_U676 | ~new_U675;
  assign U347 = ~new_U678 | ~new_U677;
  assign U348 = ~new_U680 | ~new_U679;
  assign U349 = ~new_U682 | ~new_U681;
  assign U350 = ~new_U684 | ~new_U683;
  assign U351 = ~new_U686 | ~new_U685;
  assign U352 = ~new_U688 | ~new_U687;
  assign U353 = ~new_U690 | ~new_U689;
  assign U354 = ~new_U692 | ~new_U691;
  assign U355 = ~new_U694 | ~new_U693;
  assign U356 = ~new_U696 | ~new_U695;
  assign U357 = ~new_U698 | ~new_U697;
  assign U358 = ~new_U700 | ~new_U699;
  assign U359 = ~new_U702 | ~new_U701;
  assign U360 = ~new_U704 | ~new_U703;
  assign U361 = ~new_U706 | ~new_U705;
  assign U362 = ~new_U708 | ~new_U707;
  assign U363 = ~new_U710 | ~new_U709;
  assign U364 = ~new_U712 | ~new_U711;
  assign U365 = ~new_U714 | ~new_U713;
  assign U366 = ~new_U716 | ~new_U715;
  assign U367 = ~new_U718 | ~new_U717;
  assign U368 = ~new_U720 | ~new_U719;
  assign U369 = ~new_U722 | ~new_U721;
  assign U370 = ~new_U724 | ~new_U723;
  assign U371 = ~new_U726 | ~new_U725;
  assign U372 = ~new_U728 | ~new_U727;
  assign U373 = ~new_U730 | ~new_U729;
  assign U374 = ~new_U732 | ~new_U731;
  assign U375 = ~new_U734 | ~new_U733;
  assign U376 = ~new_U736 | ~new_U735;
  assign new_U377 = ~P2_BE_N_REG_1_ & ~P2_BE_N_REG_2_ & ~P2_BE_N_REG_0_ & ~P2_ADS_N_REG;
  assign new_U378 = ~P2_D_C_N_REG & ~P2_BE_N_REG_3_;
  assign new_U379 = ~P3_W_R_N_REG & ~P3_D_C_N_REG & ~P3_ADS_N_REG & ~P3_BE_N_REG_1_ & ~P3_BE_N_REG_0_;
  assign new_U380 = ~P3_BE_N_REG_3_ & ~P3_BE_N_REG_2_;
  assign new_U381 = ~P1_BE_N_REG_0_ & ~P1_ADS_N_REG & ~P1_D_C_N_REG & ~P1_BE_N_REG_1_ & ~P1_BE_N_REG_3_;
  assign new_U382 = ~new_LT_782_119_U6 | ~new_LT_782_120_U6 | ~new_LT_782_U6;
  assign new_U383 = ~P1_BE_N_REG_2_;
  assign new_U384 = ~new_U382;
  assign new_U385 = ~n615;
  assign new_U386 = ~n605;
  assign new_U387 = ~new_R170_U6 | ~new_U208;
  assign new_U388 = ~new_U250;
  assign new_U389 = ~P2_DATAO_REG_0_ | ~new_U207;
  assign new_U390 = ~P1_DATAO_REG_0_ | ~new_U385;
  assign new_U391 = ~BUF1_REG_0_ | ~new_U388;
  assign new_U392 = ~P2_DATAO_REG_1_ | ~new_U207;
  assign new_U393 = ~P1_DATAO_REG_1_ | ~new_U385;
  assign new_U394 = ~BUF1_REG_1_ | ~new_U388;
  assign new_U395 = ~P2_DATAO_REG_2_ | ~new_U207;
  assign new_U396 = ~P1_DATAO_REG_2_ | ~new_U385;
  assign new_U397 = ~BUF1_REG_2_ | ~new_U388;
  assign new_U398 = ~P2_DATAO_REG_3_ | ~new_U207;
  assign new_U399 = ~P1_DATAO_REG_3_ | ~new_U385;
  assign new_U400 = ~BUF1_REG_3_ | ~new_U388;
  assign new_U401 = ~P2_DATAO_REG_4_ | ~new_U207;
  assign new_U402 = ~P1_DATAO_REG_4_ | ~new_U385;
  assign new_U403 = ~BUF1_REG_4_ | ~new_U388;
  assign new_U404 = ~P2_DATAO_REG_5_ | ~new_U207;
  assign new_U405 = ~P1_DATAO_REG_5_ | ~new_U385;
  assign new_U406 = ~BUF1_REG_5_ | ~new_U388;
  assign new_U407 = ~P2_DATAO_REG_6_ | ~new_U207;
  assign new_U408 = ~P1_DATAO_REG_6_ | ~new_U385;
  assign new_U409 = ~BUF1_REG_6_ | ~new_U388;
  assign new_U410 = ~P2_DATAO_REG_7_ | ~new_U207;
  assign new_U411 = ~P1_DATAO_REG_7_ | ~new_U385;
  assign new_U412 = ~BUF1_REG_7_ | ~new_U388;
  assign new_U413 = ~P2_DATAO_REG_8_ | ~new_U207;
  assign new_U414 = ~P1_DATAO_REG_8_ | ~new_U385;
  assign new_U415 = ~BUF1_REG_8_ | ~new_U388;
  assign new_U416 = ~P2_DATAO_REG_9_ | ~new_U207;
  assign new_U417 = ~P1_DATAO_REG_9_ | ~new_U385;
  assign new_U418 = ~BUF1_REG_9_ | ~new_U388;
  assign new_U419 = ~P2_DATAO_REG_10_ | ~new_U207;
  assign new_U420 = ~P1_DATAO_REG_10_ | ~new_U385;
  assign new_U421 = ~BUF1_REG_10_ | ~new_U388;
  assign new_U422 = ~P2_DATAO_REG_11_ | ~new_U207;
  assign new_U423 = ~P1_DATAO_REG_11_ | ~new_U385;
  assign new_U424 = ~BUF1_REG_11_ | ~new_U388;
  assign new_U425 = ~P2_DATAO_REG_12_ | ~new_U207;
  assign new_U426 = ~P1_DATAO_REG_12_ | ~new_U385;
  assign new_U427 = ~BUF1_REG_12_ | ~new_U388;
  assign new_U428 = ~P2_DATAO_REG_13_ | ~new_U207;
  assign new_U429 = ~P1_DATAO_REG_13_ | ~new_U385;
  assign new_U430 = ~BUF1_REG_13_ | ~new_U388;
  assign new_U431 = ~P2_DATAO_REG_14_ | ~new_U207;
  assign new_U432 = ~P1_DATAO_REG_14_ | ~new_U385;
  assign new_U433 = ~BUF1_REG_14_ | ~new_U388;
  assign new_U434 = ~P2_DATAO_REG_15_ | ~new_U207;
  assign new_U435 = ~P1_DATAO_REG_15_ | ~new_U385;
  assign new_U436 = ~BUF1_REG_15_ | ~new_U388;
  assign new_U437 = ~P2_DATAO_REG_16_ | ~new_U207;
  assign new_U438 = ~P1_DATAO_REG_16_ | ~new_U385;
  assign new_U439 = ~BUF1_REG_16_ | ~new_U388;
  assign new_U440 = ~P2_DATAO_REG_17_ | ~new_U207;
  assign new_U441 = ~P1_DATAO_REG_17_ | ~new_U385;
  assign new_U442 = ~BUF1_REG_17_ | ~new_U388;
  assign new_U443 = ~P2_DATAO_REG_18_ | ~new_U207;
  assign new_U444 = ~P1_DATAO_REG_18_ | ~new_U385;
  assign new_U445 = ~BUF1_REG_18_ | ~new_U388;
  assign new_U446 = ~P2_DATAO_REG_19_ | ~new_U207;
  assign new_U447 = ~P1_DATAO_REG_19_ | ~new_U385;
  assign new_U448 = ~BUF1_REG_19_ | ~new_U388;
  assign new_U449 = ~P2_DATAO_REG_20_ | ~new_U207;
  assign new_U450 = ~P1_DATAO_REG_20_ | ~new_U385;
  assign new_U451 = ~BUF1_REG_20_ | ~new_U388;
  assign new_U452 = ~P2_DATAO_REG_21_ | ~new_U207;
  assign new_U453 = ~P1_DATAO_REG_21_ | ~new_U385;
  assign new_U454 = ~BUF1_REG_21_ | ~new_U388;
  assign new_U455 = ~P2_DATAO_REG_22_ | ~new_U207;
  assign new_U456 = ~P1_DATAO_REG_22_ | ~new_U385;
  assign new_U457 = ~BUF1_REG_22_ | ~new_U388;
  assign new_U458 = ~P2_DATAO_REG_23_ | ~new_U207;
  assign new_U459 = ~P1_DATAO_REG_23_ | ~new_U385;
  assign new_U460 = ~BUF1_REG_23_ | ~new_U388;
  assign new_U461 = ~P2_DATAO_REG_24_ | ~new_U207;
  assign new_U462 = ~P1_DATAO_REG_24_ | ~new_U385;
  assign new_U463 = ~BUF1_REG_24_ | ~new_U388;
  assign new_U464 = ~P2_DATAO_REG_25_ | ~new_U207;
  assign new_U465 = ~P1_DATAO_REG_25_ | ~new_U385;
  assign new_U466 = ~BUF1_REG_25_ | ~new_U388;
  assign new_U467 = ~P2_DATAO_REG_26_ | ~new_U207;
  assign new_U468 = ~P1_DATAO_REG_26_ | ~new_U385;
  assign new_U469 = ~BUF1_REG_26_ | ~new_U388;
  assign new_U470 = ~P2_DATAO_REG_27_ | ~new_U207;
  assign new_U471 = ~P1_DATAO_REG_27_ | ~new_U385;
  assign new_U472 = ~BUF1_REG_27_ | ~new_U388;
  assign new_U473 = ~P2_DATAO_REG_28_ | ~new_U207;
  assign new_U474 = ~P1_DATAO_REG_28_ | ~new_U385;
  assign new_U475 = ~BUF1_REG_28_ | ~new_U388;
  assign new_U476 = ~P2_DATAO_REG_29_ | ~new_U207;
  assign new_U477 = ~P1_DATAO_REG_29_ | ~new_U385;
  assign new_U478 = ~BUF1_REG_29_ | ~new_U388;
  assign new_U479 = ~P2_DATAO_REG_30_ | ~new_U207;
  assign new_U480 = ~P1_DATAO_REG_30_ | ~new_U385;
  assign new_U481 = ~BUF1_REG_30_ | ~new_U388;
  assign new_U482 = ~P2_DATAO_REG_31_ | ~new_U207;
  assign new_U483 = ~P1_DATAO_REG_31_ | ~new_U385;
  assign new_U484 = ~BUF1_REG_31_ | ~new_U388;
  assign new_U485 = ~BUF2_REG_0_ | ~n605;
  assign new_U486 = ~P2_DATAO_REG_0_ | ~new_U386;
  assign new_U487 = ~BUF2_REG_1_ | ~n605;
  assign new_U488 = ~P2_DATAO_REG_1_ | ~new_U386;
  assign new_U489 = ~BUF2_REG_2_ | ~n605;
  assign new_U490 = ~P2_DATAO_REG_2_ | ~new_U386;
  assign new_U491 = ~BUF2_REG_3_ | ~n605;
  assign new_U492 = ~P2_DATAO_REG_3_ | ~new_U386;
  assign new_U493 = ~BUF2_REG_4_ | ~n605;
  assign new_U494 = ~P2_DATAO_REG_4_ | ~new_U386;
  assign new_U495 = ~BUF2_REG_5_ | ~n605;
  assign new_U496 = ~P2_DATAO_REG_5_ | ~new_U386;
  assign new_U497 = ~BUF2_REG_6_ | ~n605;
  assign new_U498 = ~P2_DATAO_REG_6_ | ~new_U386;
  assign new_U499 = ~BUF2_REG_7_ | ~n605;
  assign new_U500 = ~P2_DATAO_REG_7_ | ~new_U386;
  assign new_U501 = ~BUF2_REG_8_ | ~n605;
  assign new_U502 = ~P2_DATAO_REG_8_ | ~new_U386;
  assign new_U503 = ~BUF2_REG_9_ | ~n605;
  assign new_U504 = ~P2_DATAO_REG_9_ | ~new_U386;
  assign new_U505 = ~BUF2_REG_10_ | ~n605;
  assign new_U506 = ~P2_DATAO_REG_10_ | ~new_U386;
  assign new_U507 = ~BUF2_REG_11_ | ~n605;
  assign new_U508 = ~P2_DATAO_REG_11_ | ~new_U386;
  assign new_U509 = ~BUF2_REG_12_ | ~n605;
  assign new_U510 = ~P2_DATAO_REG_12_ | ~new_U386;
  assign new_U511 = ~BUF2_REG_13_ | ~n605;
  assign new_U512 = ~P2_DATAO_REG_13_ | ~new_U386;
  assign new_U513 = ~BUF2_REG_14_ | ~n605;
  assign new_U514 = ~P2_DATAO_REG_14_ | ~new_U386;
  assign new_U515 = ~BUF2_REG_15_ | ~n605;
  assign new_U516 = ~P2_DATAO_REG_15_ | ~new_U386;
  assign new_U517 = ~BUF2_REG_16_ | ~n605;
  assign new_U518 = ~P2_DATAO_REG_16_ | ~new_U386;
  assign new_U519 = ~BUF2_REG_17_ | ~n605;
  assign new_U520 = ~P2_DATAO_REG_17_ | ~new_U386;
  assign new_U521 = ~BUF2_REG_18_ | ~n605;
  assign new_U522 = ~P2_DATAO_REG_18_ | ~new_U386;
  assign new_U523 = ~BUF2_REG_19_ | ~n605;
  assign new_U524 = ~P2_DATAO_REG_19_ | ~new_U386;
  assign new_U525 = ~BUF2_REG_20_ | ~n605;
  assign new_U526 = ~P2_DATAO_REG_20_ | ~new_U386;
  assign new_U527 = ~BUF2_REG_21_ | ~n605;
  assign new_U528 = ~P2_DATAO_REG_21_ | ~new_U386;
  assign new_U529 = ~BUF2_REG_22_ | ~n605;
  assign new_U530 = ~P2_DATAO_REG_22_ | ~new_U386;
  assign new_U531 = ~BUF2_REG_23_ | ~n605;
  assign new_U532 = ~P2_DATAO_REG_23_ | ~new_U386;
  assign new_U533 = ~BUF2_REG_24_ | ~n605;
  assign new_U534 = ~P2_DATAO_REG_24_ | ~new_U386;
  assign new_U535 = ~BUF2_REG_25_ | ~n605;
  assign new_U536 = ~P2_DATAO_REG_25_ | ~new_U386;
  assign new_U537 = ~BUF2_REG_26_ | ~n605;
  assign new_U538 = ~P2_DATAO_REG_26_ | ~new_U386;
  assign new_U539 = ~BUF2_REG_27_ | ~n605;
  assign new_U540 = ~P2_DATAO_REG_27_ | ~new_U386;
  assign new_U541 = ~BUF2_REG_28_ | ~n605;
  assign new_U542 = ~P2_DATAO_REG_28_ | ~new_U386;
  assign new_U543 = ~BUF2_REG_29_ | ~n605;
  assign new_U544 = ~P2_DATAO_REG_29_ | ~new_U386;
  assign new_U545 = ~BUF2_REG_30_ | ~n605;
  assign new_U546 = ~P2_DATAO_REG_30_ | ~new_U386;
  assign new_U547 = ~BUF2_REG_31_ | ~n605;
  assign new_U548 = ~P2_DATAO_REG_31_ | ~new_U386;
  assign new_U549 = ~BUF2_REG_9_ | ~new_U249;
  assign new_U550 = ~BUF1_REG_9_ | ~new_R170_U6;
  assign new_U551 = ~BUF2_REG_8_ | ~new_U249;
  assign new_U552 = ~BUF1_REG_8_ | ~new_R170_U6;
  assign new_U553 = ~BUF2_REG_7_ | ~new_U249;
  assign new_U554 = ~BUF1_REG_7_ | ~new_R170_U6;
  assign new_U555 = ~BUF2_REG_6_ | ~new_U249;
  assign new_U556 = ~BUF1_REG_6_ | ~new_R170_U6;
  assign new_U557 = ~BUF2_REG_5_ | ~new_U249;
  assign new_U558 = ~BUF1_REG_5_ | ~new_R170_U6;
  assign new_U559 = ~BUF2_REG_4_ | ~new_U249;
  assign new_U560 = ~BUF1_REG_4_ | ~new_R170_U6;
  assign new_U561 = ~BUF2_REG_3_ | ~new_U249;
  assign new_U562 = ~BUF1_REG_3_ | ~new_R170_U6;
  assign new_U563 = ~BUF2_REG_31_ | ~new_U249;
  assign new_U564 = ~BUF1_REG_31_ | ~new_R170_U6;
  assign new_U565 = ~BUF2_REG_30_ | ~new_U249;
  assign new_U566 = ~BUF1_REG_30_ | ~new_R170_U6;
  assign new_U567 = ~BUF2_REG_2_ | ~new_U249;
  assign new_U568 = ~BUF1_REG_2_ | ~new_R170_U6;
  assign new_U569 = ~BUF2_REG_29_ | ~new_U249;
  assign new_U570 = ~BUF1_REG_29_ | ~new_R170_U6;
  assign new_U571 = ~BUF2_REG_28_ | ~new_U249;
  assign new_U572 = ~BUF1_REG_28_ | ~new_R170_U6;
  assign new_U573 = ~BUF2_REG_27_ | ~new_U249;
  assign new_U574 = ~BUF1_REG_27_ | ~new_R170_U6;
  assign new_U575 = ~BUF2_REG_26_ | ~new_U249;
  assign new_U576 = ~BUF1_REG_26_ | ~new_R170_U6;
  assign new_U577 = ~BUF2_REG_25_ | ~new_U249;
  assign new_U578 = ~BUF1_REG_25_ | ~new_R170_U6;
  assign new_U579 = ~BUF2_REG_24_ | ~new_U249;
  assign new_U580 = ~BUF1_REG_24_ | ~new_R170_U6;
  assign new_U581 = ~BUF2_REG_23_ | ~new_U249;
  assign new_U582 = ~BUF1_REG_23_ | ~new_R170_U6;
  assign new_U583 = ~BUF2_REG_22_ | ~new_U249;
  assign new_U584 = ~BUF1_REG_22_ | ~new_R170_U6;
  assign new_U585 = ~BUF2_REG_21_ | ~new_U249;
  assign new_U586 = ~BUF1_REG_21_ | ~new_R170_U6;
  assign new_U587 = ~BUF2_REG_20_ | ~new_U249;
  assign new_U588 = ~BUF1_REG_20_ | ~new_R170_U6;
  assign new_U589 = ~BUF2_REG_1_ | ~new_U249;
  assign new_U590 = ~BUF1_REG_1_ | ~new_R170_U6;
  assign new_U591 = ~BUF2_REG_19_ | ~new_U249;
  assign new_U592 = ~BUF1_REG_19_ | ~new_R170_U6;
  assign new_U593 = ~BUF2_REG_18_ | ~new_U249;
  assign new_U594 = ~BUF1_REG_18_ | ~new_R170_U6;
  assign new_U595 = ~BUF2_REG_17_ | ~new_U249;
  assign new_U596 = ~BUF1_REG_17_ | ~new_R170_U6;
  assign new_U597 = ~BUF2_REG_16_ | ~new_U249;
  assign new_U598 = ~BUF1_REG_16_ | ~new_R170_U6;
  assign new_U599 = ~BUF2_REG_15_ | ~new_U249;
  assign new_U600 = ~BUF1_REG_15_ | ~new_R170_U6;
  assign new_U601 = ~BUF2_REG_14_ | ~new_U249;
  assign new_U602 = ~BUF1_REG_14_ | ~new_R170_U6;
  assign new_U603 = ~BUF2_REG_13_ | ~new_U249;
  assign new_U604 = ~BUF1_REG_13_ | ~new_R170_U6;
  assign new_U605 = ~BUF2_REG_12_ | ~new_U249;
  assign new_U606 = ~BUF1_REG_12_ | ~new_R170_U6;
  assign new_U607 = ~BUF2_REG_11_ | ~new_U249;
  assign new_U608 = ~BUF1_REG_11_ | ~new_R170_U6;
  assign new_U609 = ~BUF2_REG_10_ | ~new_U249;
  assign new_U610 = ~BUF1_REG_10_ | ~new_R170_U6;
  assign new_U611 = ~BUF2_REG_0_ | ~new_U249;
  assign new_U612 = ~BUF1_REG_0_ | ~new_R170_U6;
  assign new_U613 = ~DATAI_9_ | ~new_U248;
  assign new_U614 = ~BUF1_REG_9_ | ~new_R165_U6;
  assign new_U615 = ~DATAI_8_ | ~new_U248;
  assign new_U616 = ~BUF1_REG_8_ | ~new_R165_U6;
  assign new_U617 = ~DATAI_7_ | ~new_U248;
  assign new_U618 = ~BUF1_REG_7_ | ~new_R165_U6;
  assign new_U619 = ~DATAI_6_ | ~new_U248;
  assign new_U620 = ~BUF1_REG_6_ | ~new_R165_U6;
  assign new_U621 = ~DATAI_5_ | ~new_U248;
  assign new_U622 = ~BUF1_REG_5_ | ~new_R165_U6;
  assign new_U623 = ~DATAI_4_ | ~new_U248;
  assign new_U624 = ~BUF1_REG_4_ | ~new_R165_U6;
  assign new_U625 = ~DATAI_3_ | ~new_U248;
  assign new_U626 = ~BUF1_REG_3_ | ~new_R165_U6;
  assign new_U627 = ~DATAI_31_ | ~new_U248;
  assign new_U628 = ~BUF1_REG_31_ | ~new_R165_U6;
  assign new_U629 = ~DATAI_30_ | ~new_U248;
  assign new_U630 = ~BUF1_REG_30_ | ~new_R165_U6;
  assign new_U631 = ~DATAI_2_ | ~new_U248;
  assign new_U632 = ~BUF1_REG_2_ | ~new_R165_U6;
  assign new_U633 = ~DATAI_29_ | ~new_U248;
  assign new_U634 = ~BUF1_REG_29_ | ~new_R165_U6;
  assign new_U635 = ~DATAI_28_ | ~new_U248;
  assign new_U636 = ~BUF1_REG_28_ | ~new_R165_U6;
  assign new_U637 = ~DATAI_27_ | ~new_U248;
  assign new_U638 = ~BUF1_REG_27_ | ~new_R165_U6;
  assign new_U639 = ~DATAI_26_ | ~new_U248;
  assign new_U640 = ~BUF1_REG_26_ | ~new_R165_U6;
  assign new_U641 = ~DATAI_25_ | ~new_U248;
  assign new_U642 = ~BUF1_REG_25_ | ~new_R165_U6;
  assign new_U643 = ~DATAI_24_ | ~new_U248;
  assign new_U644 = ~BUF1_REG_24_ | ~new_R165_U6;
  assign new_U645 = ~DATAI_23_ | ~new_U248;
  assign new_U646 = ~BUF1_REG_23_ | ~new_R165_U6;
  assign new_U647 = ~DATAI_22_ | ~new_U248;
  assign new_U648 = ~BUF1_REG_22_ | ~new_R165_U6;
  assign new_U649 = ~DATAI_21_ | ~new_U248;
  assign new_U650 = ~BUF1_REG_21_ | ~new_R165_U6;
  assign new_U651 = ~DATAI_20_ | ~new_U248;
  assign new_U652 = ~BUF1_REG_20_ | ~new_R165_U6;
  assign new_U653 = ~DATAI_1_ | ~new_U248;
  assign new_U654 = ~BUF1_REG_1_ | ~new_R165_U6;
  assign new_U655 = ~DATAI_19_ | ~new_U248;
  assign new_U656 = ~BUF1_REG_19_ | ~new_R165_U6;
  assign new_U657 = ~DATAI_18_ | ~new_U248;
  assign new_U658 = ~BUF1_REG_18_ | ~new_R165_U6;
  assign new_U659 = ~DATAI_17_ | ~new_U248;
  assign new_U660 = ~BUF1_REG_17_ | ~new_R165_U6;
  assign new_U661 = ~DATAI_16_ | ~new_U248;
  assign new_U662 = ~BUF1_REG_16_ | ~new_R165_U6;
  assign new_U663 = ~DATAI_15_ | ~new_U248;
  assign new_U664 = ~BUF1_REG_15_ | ~new_R165_U6;
  assign new_U665 = ~DATAI_14_ | ~new_U248;
  assign new_U666 = ~BUF1_REG_14_ | ~new_R165_U6;
  assign new_U667 = ~DATAI_13_ | ~new_U248;
  assign new_U668 = ~BUF1_REG_13_ | ~new_R165_U6;
  assign new_U669 = ~DATAI_12_ | ~new_U248;
  assign new_U670 = ~BUF1_REG_12_ | ~new_R165_U6;
  assign new_U671 = ~DATAI_11_ | ~new_U248;
  assign new_U672 = ~BUF1_REG_11_ | ~new_R165_U6;
  assign new_U673 = ~DATAI_10_ | ~new_U248;
  assign new_U674 = ~BUF1_REG_10_ | ~new_R165_U6;
  assign new_U675 = ~DATAI_0_ | ~new_U248;
  assign new_U676 = ~BUF1_REG_0_ | ~new_R165_U6;
  assign new_U677 = ~P2_ADDRESS_REG_9_ | ~new_U382;
  assign new_U678 = ~P3_ADDRESS_REG_9_ | ~new_U384;
  assign new_U679 = ~P2_ADDRESS_REG_8_ | ~new_U382;
  assign new_U680 = ~P3_ADDRESS_REG_8_ | ~new_U384;
  assign new_U681 = ~P2_ADDRESS_REG_7_ | ~new_U382;
  assign new_U682 = ~P3_ADDRESS_REG_7_ | ~new_U384;
  assign new_U683 = ~P2_ADDRESS_REG_6_ | ~new_U382;
  assign new_U684 = ~P3_ADDRESS_REG_6_ | ~new_U384;
  assign new_U685 = ~P2_ADDRESS_REG_5_ | ~new_U382;
  assign new_U686 = ~P3_ADDRESS_REG_5_ | ~new_U384;
  assign new_U687 = ~P2_ADDRESS_REG_4_ | ~new_U382;
  assign new_U688 = ~P3_ADDRESS_REG_4_ | ~new_U384;
  assign new_U689 = ~P2_ADDRESS_REG_3_ | ~new_U382;
  assign new_U690 = ~P3_ADDRESS_REG_3_ | ~new_U384;
  assign new_U691 = ~P2_ADDRESS_REG_2_ | ~new_U382;
  assign new_U692 = ~P3_ADDRESS_REG_2_ | ~new_U384;
  assign new_U693 = ~P2_ADDRESS_REG_29_ | ~new_U382;
  assign new_U694 = ~P3_ADDRESS_REG_29_ | ~new_U384;
  assign new_U695 = ~P2_ADDRESS_REG_28_ | ~new_U382;
  assign new_U696 = ~P3_ADDRESS_REG_28_ | ~new_U384;
  assign new_U697 = ~P2_ADDRESS_REG_27_ | ~new_U382;
  assign new_U698 = ~P3_ADDRESS_REG_27_ | ~new_U384;
  assign new_U699 = ~P2_ADDRESS_REG_26_ | ~new_U382;
  assign new_U700 = ~P3_ADDRESS_REG_26_ | ~new_U384;
  assign new_U701 = ~P2_ADDRESS_REG_25_ | ~new_U382;
  assign new_U702 = ~P3_ADDRESS_REG_25_ | ~new_U384;
  assign new_U703 = ~P2_ADDRESS_REG_24_ | ~new_U382;
  assign new_U704 = ~P3_ADDRESS_REG_24_ | ~new_U384;
  assign new_U705 = ~P2_ADDRESS_REG_23_ | ~new_U382;
  assign new_U706 = ~P3_ADDRESS_REG_23_ | ~new_U384;
  assign new_U707 = ~P2_ADDRESS_REG_22_ | ~new_U382;
  assign new_U708 = ~P3_ADDRESS_REG_22_ | ~new_U384;
  assign new_U709 = ~P2_ADDRESS_REG_21_ | ~new_U382;
  assign new_U710 = ~P3_ADDRESS_REG_21_ | ~new_U384;
  assign new_U711 = ~P2_ADDRESS_REG_20_ | ~new_U382;
  assign new_U712 = ~P3_ADDRESS_REG_20_ | ~new_U384;
  assign new_U713 = ~P2_ADDRESS_REG_1_ | ~new_U382;
  assign new_U714 = ~P3_ADDRESS_REG_1_ | ~new_U384;
  assign new_U715 = ~P2_ADDRESS_REG_19_ | ~new_U382;
  assign new_U716 = ~P3_ADDRESS_REG_19_ | ~new_U384;
  assign new_U717 = ~P2_ADDRESS_REG_18_ | ~new_U382;
  assign new_U718 = ~P3_ADDRESS_REG_18_ | ~new_U384;
  assign new_U719 = ~P2_ADDRESS_REG_17_ | ~new_U382;
  assign new_U720 = ~P3_ADDRESS_REG_17_ | ~new_U384;
  assign new_U721 = ~P2_ADDRESS_REG_16_ | ~new_U382;
  assign new_U722 = ~P3_ADDRESS_REG_16_ | ~new_U384;
  assign new_U723 = ~P2_ADDRESS_REG_15_ | ~new_U382;
  assign new_U724 = ~P3_ADDRESS_REG_15_ | ~new_U384;
  assign new_U725 = ~P2_ADDRESS_REG_14_ | ~new_U382;
  assign new_U726 = ~P3_ADDRESS_REG_14_ | ~new_U384;
  assign new_U727 = ~P2_ADDRESS_REG_13_ | ~new_U382;
  assign new_U728 = ~P3_ADDRESS_REG_13_ | ~new_U384;
  assign new_U729 = ~P2_ADDRESS_REG_12_ | ~new_U382;
  assign new_U730 = ~P3_ADDRESS_REG_12_ | ~new_U384;
  assign new_U731 = ~P2_ADDRESS_REG_11_ | ~new_U382;
  assign new_U732 = ~P3_ADDRESS_REG_11_ | ~new_U384;
  assign new_U733 = ~P2_ADDRESS_REG_10_ | ~new_U382;
  assign new_U734 = ~P3_ADDRESS_REG_10_ | ~new_U384;
  assign new_U735 = ~P2_ADDRESS_REG_0_ | ~new_U382;
  assign new_U736 = ~P3_ADDRESS_REG_0_ | ~new_U384;
  assign new_P1_ADD_515_U179 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_ADD_515_U50;
  assign new_P1_ADD_515_U178 = ~new_P1_ADD_515_U98 | ~new_P1_ADD_515_U15;
  assign new_P1_ADD_515_U177 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_ADD_515_U14;
  assign new_P1_ADD_515_U176 = ~new_P1_ADD_515_U103 | ~new_P1_ADD_515_U25;
  assign new_P1_ADD_515_U175 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_ADD_515_U24;
  assign new_P1_ADD_515_U174 = ~new_P1_ADD_515_U112 | ~new_P1_ADD_515_U43;
  assign new_P1_ADD_515_U173 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_ADD_515_U42;
  assign new_P1_ADD_515_U172 = ~new_P1_ADD_515_U119 | ~new_P1_ADD_515_U57;
  assign new_P1_ADD_515_U171 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_ADD_515_U56;
  assign new_P3_U2352 = ~new_U209 & ~P3_STATEBS16_REG;
  assign new_P3_U2353 = new_P3_U3354 & new_P3_U2449;
  assign new_P3_U2354 = new_P3_U3688 & new_P3_U4325;
  assign new_P3_U2355 = new_P3_U3689 & new_P3_U4325;
  assign new_P3_U2356 = new_P3_U3355 & new_P3_U2353;
  assign new_P3_U2357 = new_P3_U4323 & new_P3_U2451;
  assign new_P3_U2358 = new_P3_U3690 & new_P3_U4341;
  assign new_P3_U2359 = new_P3_U4324 & new_P3_U2462;
  assign new_P3_U2360 = new_P3_U4296 & new_P3_U2462;
  assign new_P3_U2361 = new_P3_U4297 & new_P3_U2462;
  assign new_P3_U2362 = new_P3_U3691 & new_P3_U4341;
  assign new_P3_U2363 = new_P3_U5442 & new_P3_U5435;
  assign new_P3_U2364 = new_P3_U5392 & new_P3_U3204;
  assign new_P3_U2365 = new_P3_U5341 & new_P3_U3201;
  assign new_P3_U2366 = new_P3_U5290 & new_P3_U3198;
  assign new_P3_U2367 = new_P3_U5239 & new_P3_U5232;
  assign new_P3_U2368 = new_P3_U5189 & new_P3_U3193;
  assign new_P3_U2369 = new_P3_U5137 & new_P3_U3189;
  assign new_P3_U2370 = new_P3_U5085 & new_P3_U3185;
  assign new_P3_U2371 = new_P3_U5036 & new_P3_U5028;
  assign new_P3_U2372 = new_P3_U4985 & new_P3_U3176;
  assign new_P3_U2373 = new_P3_U4933 & new_P3_U3172;
  assign new_P3_U2374 = new_P3_U4881 & new_P3_U3168;
  assign new_P3_U2375 = new_P3_U4829 & new_P3_U4821;
  assign new_P3_U2376 = new_P3_U4778 & new_P3_U3160;
  assign new_P3_U2377 = new_P3_U4726 & new_P3_U3152;
  assign new_P3_U2378 = new_P3_U4674 & new_P3_U3146;
  assign new_P3_U2379 = new_P3_U4322 & new_P3_U4312;
  assign new_P3_U2380 = P3_STATE2_REG_2_ & new_P3_U3260;
  assign new_P3_U2381 = new_P3_U4312 & P3_STATE2_REG_3_;
  assign new_P3_U2382 = new_P3_U3951 & new_P3_U3249;
  assign new_P3_U2383 = new_P3_U2380 & new_P3_U4296;
  assign new_P3_U2384 = new_P3_U2380 & new_P3_U4297;
  assign new_P3_U2385 = P3_STATE2_REG_1_ & new_P3_U3260;
  assign new_P3_U2386 = P3_STATE2_REG_1_ & new_P3_U3249;
  assign new_P3_U2387 = new_P3_U3953 & new_P3_U3249;
  assign new_P3_U2388 = new_P3_U3952 & new_P3_U3249;
  assign new_P3_U2389 = new_P3_U4354 & new_P3_U3249;
  assign new_P3_U2390 = new_P3_U4353 & P3_STATE2_REG_0_;
  assign new_P3_U2391 = new_P3_U4310 & new_P3_U3218;
  assign new_P3_U2392 = new_P3_U2383 & new_P3_U4293;
  assign new_P3_U2393 = new_P3_U2628 & new_P3_U2361;
  assign new_P3_U2394 = new_P3_U2382 & new_P3_U2628;
  assign new_P3_U2395 = new_P3_U2361 & new_P3_U3241;
  assign new_P3_U2396 = new_P3_U2382 & new_P3_U3241;
  assign new_P3_U2397 = new_P3_U2386 & P3_STATEBS16_REG;
  assign new_P3_U2398 = new_P3_U2386 & new_P3_U2631;
  assign new_P3_U2399 = new_P3_U4309 & new_P3_U4573;
  assign new_P3_U2400 = new_P3_U4310 & new_P3_U4573;
  assign new_P3_U2401 = P3_STATE2_REG_3_ & new_P3_U3260;
  assign new_P3_U2402 = new_P3_U3248 & new_P3_U3090;
  assign new_P3_U2403 = new_P3_U2385 & new_P3_U3258;
  assign new_P3_U2404 = new_P3_U2384 & new_P3_U3257;
  assign new_P3_U2405 = new_P3_U7095 & new_P3_U2384;
  assign new_P3_U2406 = new_P3_U4311 & new_P3_U3104;
  assign new_P3_U2407 = new_P3_U4311 & new_P3_U4505;
  assign new_P3_U2408 = new_P3_U4309 & new_P3_U3218;
  assign new_P3_U2409 = P3_STATE2_REG_0_ & new_P3_U3251;
  assign new_P3_U2410 = new_P3_U3251 & new_P3_U3121;
  assign new_P3_U2411 = new_P3_U4310 & new_P3_U4608;
  assign new_P3_U2412 = new_P3_U4539 & new_P3_U3218 & new_P3_U3107;
  assign new_P3_U2413 = BUF2_REG_0_ & new_P3_U4312;
  assign new_P3_U2414 = BUF2_REG_1_ & new_P3_U4312;
  assign new_P3_U2415 = BUF2_REG_2_ & new_P3_U4312;
  assign new_P3_U2416 = BUF2_REG_3_ & new_P3_U4312;
  assign new_P3_U2417 = BUF2_REG_4_ & new_P3_U4312;
  assign new_P3_U2418 = BUF2_REG_5_ & new_P3_U4312;
  assign new_P3_U2419 = BUF2_REG_6_ & new_P3_U4312;
  assign new_P3_U2420 = BUF2_REG_7_ & new_P3_U4312;
  assign new_P3_U2421 = BUF2_REG_24_ & new_P3_U2379;
  assign new_P3_U2422 = BUF2_REG_16_ & new_P3_U2379;
  assign new_P3_U2423 = BUF2_REG_25_ & new_P3_U2379;
  assign new_P3_U2424 = BUF2_REG_17_ & new_P3_U2379;
  assign new_P3_U2425 = BUF2_REG_26_ & new_P3_U2379;
  assign new_P3_U2426 = BUF2_REG_18_ & new_P3_U2379;
  assign new_P3_U2427 = BUF2_REG_27_ & new_P3_U2379;
  assign new_P3_U2428 = BUF2_REG_19_ & new_P3_U2379;
  assign new_P3_U2429 = BUF2_REG_28_ & new_P3_U2379;
  assign new_P3_U2430 = BUF2_REG_20_ & new_P3_U2379;
  assign new_P3_U2431 = BUF2_REG_29_ & new_P3_U2379;
  assign new_P3_U2432 = BUF2_REG_21_ & new_P3_U2379;
  assign new_P3_U2433 = BUF2_REG_30_ & new_P3_U2379;
  assign new_P3_U2434 = BUF2_REG_22_ & new_P3_U2379;
  assign new_P3_U2435 = BUF2_REG_31_ & new_P3_U2379;
  assign new_P3_U2436 = BUF2_REG_23_ & new_P3_U2379;
  assign new_P3_U2437 = new_P3_U2381 & new_P3_U3108;
  assign new_P3_U2438 = new_P3_U2381 & new_P3_U3104;
  assign new_P3_U2439 = new_P3_U2381 & new_P3_U3101;
  assign new_P3_U2440 = new_P3_U2381 & new_P3_U3107;
  assign new_P3_U2441 = new_P3_U2381 & new_P3_U3102;
  assign new_P3_U2442 = new_P3_U2381 & new_P3_U3110;
  assign new_P3_U2443 = new_P3_U2381 & new_P3_U3074;
  assign new_P3_U2444 = new_P3_U2391 & new_P3_U3074;
  assign new_P3_U2445 = new_P3_U2381 & new_P3_U3218;
  assign new_P3_U2446 = new_P3_U2391 & new_P3_U3113;
  assign new_P3_U2447 = new_P3_U2409 & new_P3_U3108;
  assign new_P3_U2448 = new_P3_U2391 & new_P3_U4590;
  assign new_P3_U2449 = new_P3_U4344 & new_P3_U4522;
  assign new_P3_U2450 = new_P3_U3660 & new_P3_U4351;
  assign new_P3_U2451 = new_P3_U2412 & new_P3_U4608 & new_P3_U3102;
  assign new_P3_U2452 = new_P3_U2412 & new_P3_U2463 & new_P3_U4522;
  assign new_P3_U2453 = P3_STATE2_REG_2_ & P3_STATE2_REG_1_;
  assign new_P3_U2454 = new_P3_U2380 & new_P3_U4323;
  assign new_P3_U2455 = new_P3_U2380 & new_P3_U4324;
  assign new_P3_U2456 = new_P3_U4556 & new_P3_U4607;
  assign new_P3_U2457 = new_P3_U3269 & new_P3_U3139;
  assign new_P3_U2458 = new_P3_U4652 & new_P3_U3269;
  assign new_P3_U2459 = new_P3_U7962 & new_P3_U3139;
  assign new_P3_U2460 = new_P3_U7962 & new_P3_U4652;
  assign new_P3_U2461 = new_P3_U4573 & new_P3_U4522;
  assign new_P3_U2462 = new_P3_U2412 & new_P3_U2449;
  assign new_P3_U2463 = new_P3_U4590 & new_P3_U4607;
  assign new_P3_U2464 = P3_INSTQUEUERD_ADDR_REG_3_ & P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_U2465 = new_P3_U2464 & new_P3_U4332;
  assign new_P3_U2466 = P3_INSTQUEUERD_ADDR_REG_1_ & new_P3_U3093;
  assign new_P3_U2467 = new_P3_U2464 & new_P3_U2466;
  assign new_P3_U2468 = P3_INSTQUEUERD_ADDR_REG_0_ & new_P3_U3094;
  assign new_P3_U2469 = new_P3_U2464 & new_P3_U2468;
  assign new_P3_U2470 = new_P3_U2464 & new_P3_U4467;
  assign new_P3_U2471 = P3_INSTQUEUERD_ADDR_REG_3_ & new_P3_U4468;
  assign new_P3_U2472 = new_P3_U2466 & new_P3_U3097;
  assign new_P3_U2473 = new_P3_U2472 & P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_U2474 = new_P3_U2468 & new_P3_U3097;
  assign new_P3_U2475 = new_P3_U2474 & P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_U2476 = P3_INSTQUEUERD_ADDR_REG_3_ & new_P3_U4469;
  assign new_P3_U2477 = new_P3_U4470 & new_P3_U2466;
  assign new_P3_U2478 = new_P3_U4470 & new_P3_U2468;
  assign new_P3_U2479 = new_P3_U4470 & new_P3_U4467;
  assign new_P3_U2480 = new_P3_U4468 & new_P3_U3100;
  assign new_P3_U2481 = ~P3_INSTQUEUERD_ADDR_REG_3_ & ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_U2482 = new_P3_U2466 & new_P3_U2481;
  assign new_P3_U2483 = new_P3_U2468 & new_P3_U2481;
  assign new_P3_U2484 = new_P3_U4469 & new_P3_U3100;
  assign new_P3_U2485 = new_P3_U4656 & new_P3_U3270;
  assign new_P3_U2486 = new_P3_U3271 & new_P3_U3182;
  assign new_P3_U2487 = new_P3_U3270 & new_P3_U3142;
  assign new_P3_U2488 = new_P3_U4657 & new_P3_U2487;
  assign new_P3_U2489 = new_P3_U3090 & new_P3_U4315;
  assign new_P3_U2490 = P3_INSTQUEUEWR_ADDR_REG_0_ & new_P3_U3156;
  assign new_P3_U2491 = new_P3_U4644 & new_P3_U2487;
  assign new_P3_U2492 = P3_INSTQUEUEWR_ADDR_REG_2_ & new_P3_U3128;
  assign new_P3_U2493 = new_P3_U4646 & new_P3_U3128;
  assign new_P3_U2494 = new_P3_U4645 & new_P3_U2487;
  assign new_P3_U2495 = new_P3_U4646 & P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_U2496 = new_P3_U4643 & new_P3_U3128;
  assign new_P3_U2497 = new_P3_U2496 & new_P3_U2487;
  assign new_P3_U2498 = new_P3_U7968 & new_P3_U3182;
  assign new_P3_U2499 = new_P3_U4658 & new_P3_U4657;
  assign new_P3_U2500 = new_P3_U4658 & new_P3_U4644;
  assign new_P3_U2501 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_U2502 = new_P3_U4658 & new_P3_U4645;
  assign new_P3_U2503 = new_P3_U4658 & new_P3_U2496;
  assign new_P3_U2504 = new_P3_U4660 & new_P3_U3271;
  assign new_P3_U2505 = new_P3_U4644 & new_P3_U2485;
  assign new_P3_U2506 = new_P3_U4645 & new_P3_U2485;
  assign new_P3_U2507 = new_P3_U2496 & new_P3_U2485;
  assign new_P3_U2508 = new_P3_U4660 & new_P3_U7968;
  assign new_P3_U2509 = new_P3_U7965 & new_P3_U4656;
  assign new_P3_U2510 = new_P3_U2509 & new_P3_U4657;
  assign new_P3_U2511 = new_P3_U2509 & new_P3_U4644;
  assign new_P3_U2512 = new_P3_U2509 & new_P3_U4645;
  assign new_P3_U2513 = new_P3_U2509 & new_P3_U2496;
  assign new_P3_U2514 = new_P3_U3218 & new_P3_U3216;
  assign new_P3_U2515 = new_P3_U5485 & new_P3_U7970 & new_P3_U7969;
  assign new_P3_U2516 = new_P3_U5493 & new_P3_U5492;
  assign new_P3_U2517 = new_P3_U3246 & new_P3_U5526;
  assign new_P3_U2518 = new_P3_U3668 & new_P3_U5522;
  assign new_P3_U2519 = P3_INSTQUEUERD_ADDR_REG_0_ & new_P3_U3228;
  assign new_P3_U2520 = new_P3_U5543 & new_P3_U5548;
  assign new_P3_U2521 = new_P3_U2520 & new_P3_U2519;
  assign new_P3_U2522 = new_P3_U3093 & new_P3_U3228;
  assign new_P3_U2523 = new_P3_U2520 & new_P3_U2522;
  assign new_P3_U2524 = new_P3_U5558 & P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_U2525 = new_P3_U2520 & new_P3_U2524;
  assign new_P3_U2526 = new_P3_U5558 & new_P3_U3093;
  assign new_P3_U2527 = new_P3_U2520 & new_P3_U2526;
  assign new_P3_U2528 = new_P3_U5543 & new_P3_U3225;
  assign new_P3_U2529 = new_P3_U2528 & new_P3_U2519;
  assign new_P3_U2530 = new_P3_U2528 & new_P3_U2522;
  assign new_P3_U2531 = new_P3_U2528 & new_P3_U2524;
  assign new_P3_U2532 = new_P3_U2528 & new_P3_U2526;
  assign new_P3_U2533 = new_P3_U5548 & new_P3_U3265;
  assign new_P3_U2534 = new_P3_U2533 & new_P3_U2519;
  assign new_P3_U2535 = new_P3_U2533 & new_P3_U2522;
  assign new_P3_U2536 = new_P3_U2533 & new_P3_U2524;
  assign new_P3_U2537 = new_P3_U2533 & new_P3_U2526;
  assign new_P3_U2538 = new_P3_U3265 & new_P3_U3225;
  assign new_P3_U2539 = new_P3_U2519 & new_P3_U2538;
  assign new_P3_U2540 = new_P3_U2522 & new_P3_U2538;
  assign new_P3_U2541 = new_P3_U2524 & new_P3_U2538;
  assign new_P3_U2542 = new_P3_U2526 & new_P3_U2538;
  assign new_P3_U2543 = new_P3_U3272 & new_P3_U3266;
  assign new_P3_U2544 = new_P3_U2543 & new_P3_U2468;
  assign new_P3_U2545 = new_P3_U2543 & new_P3_U4467;
  assign new_P3_U2546 = new_P3_U2543 & new_P3_U4332;
  assign new_P3_U2547 = new_P3_U2543 & new_P3_U2466;
  assign new_P3_U2548 = new_P3_U8034 & new_P3_U3266;
  assign new_P3_U2549 = new_P3_U2548 & new_P3_U2468;
  assign new_P3_U2550 = new_P3_U2548 & new_P3_U4467;
  assign new_P3_U2551 = new_P3_U2548 & new_P3_U4332;
  assign new_P3_U2552 = new_P3_U2548 & new_P3_U2466;
  assign new_P3_U2553 = new_P3_U7516 & new_P3_U3272;
  assign new_P3_U2554 = new_P3_U2553 & new_P3_U2468;
  assign new_P3_U2555 = new_P3_U2553 & new_P3_U4467;
  assign new_P3_U2556 = new_P3_U2553 & new_P3_U4332;
  assign new_P3_U2557 = new_P3_U2553 & new_P3_U2466;
  assign new_P3_U2558 = new_P3_U7516 & new_P3_U8034;
  assign new_P3_U2559 = new_P3_U2558 & new_P3_U2468;
  assign new_P3_U2560 = new_P3_U2558 & new_P3_U4467;
  assign new_P3_U2561 = new_P3_U2558 & new_P3_U4332;
  assign new_P3_U2562 = new_P3_U2558 & new_P3_U2466;
  assign new_P3_U2563 = new_P3_U8037 & new_P3_U4291;
  assign new_P3_U2564 = new_P3_U2563 & new_P3_U2522;
  assign new_P3_U2565 = new_P3_U2563 & new_P3_U2519;
  assign new_P3_U2566 = new_P3_U2563 & new_P3_U2526;
  assign new_P3_U2567 = new_P3_U2563 & new_P3_U2524;
  assign new_P3_U2568 = new_P3_U8037 & new_P3_U3267;
  assign new_P3_U2569 = new_P3_U2568 & new_P3_U2522;
  assign new_P3_U2570 = new_P3_U2568 & new_P3_U2519;
  assign new_P3_U2571 = new_P3_U2568 & new_P3_U2526;
  assign new_P3_U2572 = new_P3_U2568 & new_P3_U2524;
  assign new_P3_U2573 = new_P3_U4291 & new_P3_U3273;
  assign new_P3_U2574 = new_P3_U2573 & new_P3_U2522;
  assign new_P3_U2575 = new_P3_U2573 & new_P3_U2519;
  assign new_P3_U2576 = new_P3_U2573 & new_P3_U2526;
  assign new_P3_U2577 = new_P3_U2573 & new_P3_U2524;
  assign new_P3_U2578 = new_P3_U3273 & new_P3_U3267;
  assign new_P3_U2579 = new_P3_U2578 & new_P3_U2522;
  assign new_P3_U2580 = new_P3_U2578 & new_P3_U2519;
  assign new_P3_U2581 = new_P3_U2578 & new_P3_U2526;
  assign new_P3_U2582 = new_P3_U2578 & new_P3_U2524;
  assign new_P3_U2583 = new_P3_U7775 & new_P3_U4468;
  assign new_P3_U2584 = new_P3_U7775 & new_P3_U2472;
  assign new_P3_U2585 = new_P3_U7775 & new_P3_U2474;
  assign new_P3_U2586 = new_P3_U7775 & new_P3_U4469;
  assign new_P3_U2587 = new_P3_U7775 & P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_U2588 = new_P3_U2587 & new_P3_U4332;
  assign new_P3_U2589 = new_P3_U2587 & new_P3_U2466;
  assign new_P3_U2590 = new_P3_U2587 & new_P3_U2468;
  assign new_P3_U2591 = new_P3_U2587 & new_P3_U4467;
  assign new_P3_U2592 = new_P3_U4468 & new_P3_U3268;
  assign new_P3_U2593 = new_P3_U2472 & new_P3_U3268;
  assign new_P3_U2594 = new_P3_U2474 & new_P3_U3268;
  assign new_P3_U2595 = new_P3_U4469 & new_P3_U3268;
  assign new_P3_U2596 = P3_INSTQUEUERD_ADDR_REG_2_ & new_P3_U3268;
  assign new_P3_U2597 = new_P3_U2596 & new_P3_U4332;
  assign new_P3_U2598 = new_P3_U2596 & new_P3_U2466;
  assign new_P3_U2599 = new_P3_U2596 & new_P3_U2468;
  assign new_P3_U2600 = new_P3_U2596 & new_P3_U4467;
  assign new_P3_U2601 = new_P3_U2392 & new_P3_U2352;
  assign new_P3_U2602 = P3_EBX_REG_31_ & new_P3_U2404;
  assign new_P3_U2603 = new_P3_U4133 & new_P3_U7359 & new_P3_U7360 & new_P3_U7358;
  assign new_P3_U2604 = new_P3_U7947 & new_P3_U7946;
  assign new_P3_U2605 = ~new_P3_U4212 | ~new_P3_U4213 | ~new_P3_U4215 | ~new_P3_U4214;
  assign new_P3_U2606 = ~new_P3_U4208 | ~new_P3_U4209 | ~new_P3_U4211 | ~new_P3_U4210;
  assign new_P3_U2607 = ~new_P3_U4204 | ~new_P3_U4205 | ~new_P3_U4207 | ~new_P3_U4206;
  assign new_P3_U2608 = ~new_P3_U4200 | ~new_P3_U4201 | ~new_P3_U4203 | ~new_P3_U4202;
  assign new_P3_U2609 = ~new_P3_U4196 | ~new_P3_U4197 | ~new_P3_U4199 | ~new_P3_U4198;
  assign new_P3_U2610 = ~new_P3_U4192 | ~new_P3_U4193 | ~new_P3_U4195 | ~new_P3_U4194;
  assign new_P3_U2611 = ~new_P3_U4188 | ~new_P3_U4189 | ~new_P3_U4191 | ~new_P3_U4190;
  assign new_P3_U2612 = ~new_P3_U4184 | ~new_P3_U4185 | ~new_P3_U4187 | ~new_P3_U4186;
  assign new_P3_U2613 = ~new_P3_U4276 | ~new_P3_U4277 | ~new_P3_U4279 | ~new_P3_U4278;
  assign new_P3_U2614 = ~new_P3_U4272 | ~new_P3_U4273 | ~new_P3_U4275 | ~new_P3_U4274;
  assign new_P3_U2615 = ~new_P3_U4268 | ~new_P3_U4269 | ~new_P3_U4271 | ~new_P3_U4270;
  assign new_P3_U2616 = ~new_P3_U4264 | ~new_P3_U4265 | ~new_P3_U4267 | ~new_P3_U4266;
  assign new_P3_U2617 = ~new_P3_U4260 | ~new_P3_U4261 | ~new_P3_U4263 | ~new_P3_U4262;
  assign new_P3_U2618 = ~new_P3_U4256 | ~new_P3_U4257 | ~new_P3_U4259 | ~new_P3_U4258;
  assign new_P3_U2619 = ~new_P3_U4252 | ~new_P3_U4253 | ~new_P3_U4255 | ~new_P3_U4254;
  assign new_P3_U2620 = ~new_P3_U4248 | ~new_P3_U4249 | ~new_P3_U4251 | ~new_P3_U4250;
  assign new_P3_U2621 = ~new_P3_U4180 | ~new_P3_U4181 | ~new_P3_U4183 | ~new_P3_U4182;
  assign new_P3_U2622 = ~new_P3_U4176 | ~new_P3_U4177 | ~new_P3_U4179 | ~new_P3_U4178;
  assign new_P3_U2623 = ~new_P3_U4172 | ~new_P3_U4173 | ~new_P3_U4175 | ~new_P3_U4174;
  assign new_P3_U2624 = ~new_P3_U4168 | ~new_P3_U4169 | ~new_P3_U4171 | ~new_P3_U4170;
  assign new_P3_U2625 = ~new_P3_U4164 | ~new_P3_U4165 | ~new_P3_U4167 | ~new_P3_U4166;
  assign new_P3_U2626 = ~new_P3_U4160 | ~new_P3_U4161 | ~new_P3_U4163 | ~new_P3_U4162;
  assign new_P3_U2627 = ~new_P3_U4156 | ~new_P3_U4157 | ~new_P3_U4159 | ~new_P3_U4158;
  assign new_P3_U2628 = ~new_P3_U4152 | ~new_P3_U4153 | ~new_P3_U4155 | ~new_P3_U4154;
  assign new_P3_U2629 = P3_INSTQUEUERD_ADDR_REG_4_ & new_P3_U3207;
  assign new_P3_U2630 = ~new_U209;
  assign new_P3_U2631 = ~P3_STATEBS16_REG;
  assign new_P3_U2632 = P3_INSTQUEUERD_ADDR_REG_3_ & new_P3_U3207;
  assign n2815 = ~new_P3_U7937 | ~new_P3_U7383;
  assign n2810 = ~new_P3_U7382 | ~new_P3_U7381;
  assign n2802 = ~new_P3_U4335 | ~new_P3_U8025 | ~new_P3_U8024;
  assign n2792 = ~new_P3_U4335 | ~new_P3_U8021 | ~new_P3_U8020;
  assign n2782 = ~new_P3_U7370 | ~new_P3_U7369;
  assign n2768 = ~new_P3_U4327 | ~new_P3_U8013 | ~new_P3_U8012;
  assign n2758 = ~new_P3_U4327 | ~new_P3_U8003 | ~new_P3_U8002;
  assign n2753 = new_P3_U7357 & new_P3_U7907;
  assign n2748 = ~new_P3_U4130 | ~new_P3_U7354 | ~new_P3_U4129 | ~new_P3_U7352 | ~new_P3_U7351;
  assign n2743 = ~new_P3_U4127 | ~new_P3_U7346 | ~new_P3_U4126 | ~new_P3_U7344 | ~new_P3_U7343;
  assign n2738 = ~new_P3_U4124 | ~new_P3_U7338 | ~new_P3_U4123 | ~new_P3_U7336 | ~new_P3_U7335;
  assign n2733 = ~new_P3_U4121 | ~new_P3_U7330 | ~new_P3_U4120 | ~new_P3_U7328 | ~new_P3_U7327;
  assign n2728 = ~new_P3_U4118 | ~new_P3_U7322 | ~new_P3_U4117 | ~new_P3_U7320 | ~new_P3_U7319;
  assign n2723 = ~new_P3_U4115 | ~new_P3_U7314 | ~new_P3_U4114 | ~new_P3_U7312 | ~new_P3_U7311;
  assign n2718 = ~new_P3_U4112 | ~new_P3_U7306 | ~new_P3_U4111 | ~new_P3_U7304 | ~new_P3_U7303;
  assign n2713 = ~new_P3_U4109 | ~new_P3_U7298 | ~new_P3_U4108 | ~new_P3_U7296 | ~new_P3_U7295;
  assign n2708 = ~new_P3_U4106 | ~new_P3_U7290 | ~new_P3_U4105 | ~new_P3_U7288 | ~new_P3_U7287;
  assign n2703 = ~new_P3_U4103 | ~new_P3_U7282 | ~new_P3_U4102 | ~new_P3_U7280 | ~new_P3_U7279;
  assign n2698 = ~new_P3_U4100 | ~new_P3_U7274 | ~new_P3_U4099 | ~new_P3_U7272 | ~new_P3_U7271;
  assign n2693 = ~new_P3_U4097 | ~new_P3_U7266 | ~new_P3_U4096 | ~new_P3_U7264 | ~new_P3_U7263;
  assign n2688 = ~new_P3_U4094 | ~new_P3_U7258 | ~new_P3_U4093 | ~new_P3_U7256 | ~new_P3_U7255;
  assign n2683 = ~new_P3_U4091 | ~new_P3_U7250 | ~new_P3_U4090 | ~new_P3_U7248 | ~new_P3_U7247;
  assign n2678 = ~new_P3_U4088 | ~new_P3_U7242 | ~new_P3_U4087 | ~new_P3_U7240 | ~new_P3_U7239;
  assign n2673 = ~new_P3_U4085 | ~new_P3_U7234 | ~new_P3_U4084 | ~new_P3_U7232 | ~new_P3_U7231;
  assign n2668 = ~new_P3_U4082 | ~new_P3_U7226 | ~new_P3_U4081 | ~new_P3_U7224 | ~new_P3_U7223;
  assign n2663 = ~new_P3_U4079 | ~new_P3_U7218 | ~new_P3_U4078 | ~new_P3_U7216 | ~new_P3_U7215;
  assign n2658 = ~new_P3_U4076 | ~new_P3_U7210 | ~new_P3_U4075 | ~new_P3_U7208 | ~new_P3_U7207;
  assign n2653 = ~new_P3_U4073 | ~new_P3_U7202 | ~new_P3_U4072 | ~new_P3_U7200 | ~new_P3_U7199;
  assign n2648 = ~new_P3_U4070 | ~new_P3_U7194 | ~new_P3_U4069 | ~new_P3_U7192 | ~new_P3_U7191;
  assign n2643 = ~new_P3_U4067 | ~new_P3_U7186 | ~new_P3_U4066 | ~new_P3_U7184 | ~new_P3_U7183;
  assign n2638 = ~new_P3_U4064 | ~new_P3_U7178 | ~new_P3_U4063 | ~new_P3_U7176 | ~new_P3_U7175;
  assign n2633 = ~new_P3_U4061 | ~new_P3_U7170 | ~new_P3_U4060 | ~new_P3_U7168 | ~new_P3_U7167;
  assign n2628 = ~new_P3_U4058 | ~new_P3_U7162 | ~new_P3_U4057 | ~new_P3_U7160 | ~new_P3_U7159;
  assign n2623 = ~new_P3_U4056 | ~new_P3_U4054;
  assign n2618 = ~new_P3_U4051 | ~new_P3_U4049;
  assign n2613 = ~new_P3_U4045 | ~new_P3_U7133 | ~new_P3_U7132 | ~new_P3_U7129 | ~new_P3_U4043;
  assign n2608 = ~new_P3_U4041 | ~new_P3_U7123 | ~new_P3_U7122 | ~new_P3_U7119 | ~new_P3_U4039;
  assign n2603 = ~new_P3_U4037 | ~new_P3_U7113 | ~new_P3_U7112 | ~new_P3_U7109 | ~new_P3_U4035;
  assign n2598 = ~new_P3_U4033 | ~new_P3_U7103 | ~new_P3_U7102 | ~new_P3_U7099 | ~new_P3_U4031;
  assign n2593 = ~new_P3_U7092 | ~new_P3_U7091;
  assign n2588 = ~new_P3_U7089 | ~new_P3_U7090 | ~new_P3_U7088;
  assign n2583 = ~new_P3_U7086 | ~new_P3_U7087 | ~new_P3_U7085;
  assign n2578 = ~new_P3_U7083 | ~new_P3_U7084 | ~new_P3_U7082;
  assign n2573 = ~new_P3_U7080 | ~new_P3_U7081 | ~new_P3_U7079;
  assign n2568 = ~new_P3_U7077 | ~new_P3_U7078 | ~new_P3_U7076;
  assign n2563 = ~new_P3_U7074 | ~new_P3_U7075 | ~new_P3_U7073;
  assign n2558 = ~new_P3_U7071 | ~new_P3_U7072 | ~new_P3_U7070;
  assign n2553 = ~new_P3_U7068 | ~new_P3_U7069 | ~new_P3_U7067;
  assign n2548 = ~new_P3_U7065 | ~new_P3_U7066 | ~new_P3_U7064;
  assign n2543 = ~new_P3_U7062 | ~new_P3_U7063 | ~new_P3_U7061;
  assign n2538 = ~new_P3_U7059 | ~new_P3_U7060 | ~new_P3_U7058;
  assign n2533 = ~new_P3_U7056 | ~new_P3_U7057 | ~new_P3_U7055;
  assign n2528 = ~new_P3_U7053 | ~new_P3_U7054 | ~new_P3_U7052;
  assign n2523 = ~new_P3_U7050 | ~new_P3_U7051 | ~new_P3_U7049;
  assign n2518 = ~new_P3_U7047 | ~new_P3_U7048 | ~new_P3_U7046;
  assign n2513 = ~new_P3_U7044 | ~new_P3_U7045 | ~new_P3_U7043;
  assign n2508 = ~new_P3_U7041 | ~new_P3_U7042 | ~new_P3_U7040;
  assign n2503 = ~new_P3_U7038 | ~new_P3_U7039 | ~new_P3_U7037;
  assign n2498 = ~new_P3_U7035 | ~new_P3_U7036 | ~new_P3_U7034;
  assign n2493 = ~new_P3_U7032 | ~new_P3_U7033 | ~new_P3_U7031;
  assign n2488 = ~new_P3_U7029 | ~new_P3_U7030 | ~new_P3_U7028;
  assign n2483 = ~new_P3_U7027 | ~new_P3_U7026 | ~new_P3_U7025;
  assign n2478 = ~new_P3_U7024 | ~new_P3_U7023 | ~new_P3_U7022;
  assign n2473 = ~new_P3_U7021 | ~new_P3_U7020 | ~new_P3_U7019;
  assign n2468 = ~new_P3_U7018 | ~new_P3_U7017 | ~new_P3_U7016;
  assign n2463 = ~new_P3_U7015 | ~new_P3_U7014 | ~new_P3_U7013;
  assign n2458 = ~new_P3_U7012 | ~new_P3_U7011 | ~new_P3_U7010;
  assign n2453 = ~new_P3_U7009 | ~new_P3_U7008 | ~new_P3_U7007;
  assign n2448 = ~new_P3_U7006 | ~new_P3_U7005 | ~new_P3_U7004;
  assign n2443 = ~new_P3_U7003 | ~new_P3_U7002 | ~new_P3_U7001;
  assign n2438 = ~new_P3_U7000 | ~new_P3_U6999 | ~new_P3_U6998;
  assign n2433 = ~new_P3_U6994 | ~new_P3_U6995 | ~new_P3_U6993;
  assign n2428 = ~new_P3_U6991 | ~new_P3_U6990 | ~new_P3_U6992 | ~new_P3_U6989 | ~new_P3_U6988;
  assign n2423 = ~new_P3_U6986 | ~new_P3_U6985 | ~new_P3_U6987 | ~new_P3_U6984 | ~new_P3_U6983;
  assign n2418 = ~new_P3_U6981 | ~new_P3_U6980 | ~new_P3_U6982 | ~new_P3_U6979 | ~new_P3_U6978;
  assign n2413 = ~new_P3_U6976 | ~new_P3_U4029 | ~new_P3_U6974 | ~new_P3_U6973;
  assign n2408 = ~new_P3_U6971 | ~new_P3_U4028 | ~new_P3_U6969 | ~new_P3_U6968;
  assign n2403 = ~new_P3_U6966 | ~new_P3_U4027 | ~new_P3_U6964 | ~new_P3_U6963;
  assign n2398 = ~new_P3_U6961 | ~new_P3_U4026 | ~new_P3_U6959 | ~new_P3_U6958;
  assign n2393 = ~new_P3_U6956 | ~new_P3_U4025 | ~new_P3_U6954 | ~new_P3_U6953;
  assign n2388 = ~new_P3_U6951 | ~new_P3_U4024 | ~new_P3_U6949 | ~new_P3_U6948;
  assign n2383 = ~new_P3_U6946 | ~new_P3_U4023 | ~new_P3_U6944 | ~new_P3_U6943;
  assign n2378 = ~new_P3_U6941 | ~new_P3_U4022 | ~new_P3_U6939 | ~new_P3_U6938;
  assign n2373 = ~new_P3_U6936 | ~new_P3_U4021 | ~new_P3_U6934 | ~new_P3_U6933;
  assign n2368 = ~new_P3_U6931 | ~new_P3_U4020 | ~new_P3_U6929 | ~new_P3_U6928;
  assign n2363 = ~new_P3_U6926 | ~new_P3_U4019 | ~new_P3_U6924 | ~new_P3_U6923;
  assign n2358 = ~new_P3_U6921 | ~new_P3_U4018 | ~new_P3_U6919 | ~new_P3_U6918;
  assign n2353 = ~new_P3_U6916 | ~new_P3_U6914 | ~new_P3_U4017;
  assign n2348 = ~new_P3_U6912 | ~new_P3_U6910 | ~new_P3_U4016;
  assign n2343 = ~new_P3_U6908 | ~new_P3_U6906 | ~new_P3_U4015;
  assign n2338 = ~new_P3_U4014 | ~new_P3_U6903 | ~new_P3_U6902;
  assign n2333 = ~new_P3_U4013 | ~new_P3_U6899 | ~new_P3_U6898;
  assign n2328 = ~new_P3_U4012 | ~new_P3_U6895 | ~new_P3_U6894;
  assign n2323 = ~new_P3_U4011 | ~new_P3_U6891 | ~new_P3_U6890;
  assign n2318 = ~new_P3_U4010 | ~new_P3_U6887 | ~new_P3_U6886;
  assign n2313 = ~new_P3_U4009 | ~new_P3_U6883 | ~new_P3_U6882;
  assign n2308 = ~new_P3_U4008 | ~new_P3_U6879 | ~new_P3_U6878;
  assign n2303 = ~new_P3_U4007 | ~new_P3_U6875 | ~new_P3_U6874;
  assign n2298 = ~new_P3_U4006 | ~new_P3_U6871 | ~new_P3_U6870;
  assign n2293 = ~new_P3_U4005 | ~new_P3_U6867 | ~new_P3_U6866;
  assign n2288 = ~new_P3_U4004 | ~new_P3_U6863 | ~new_P3_U6862;
  assign n2283 = ~new_P3_U4003 | ~new_P3_U6859 | ~new_P3_U6858;
  assign n2278 = ~new_P3_U4002 | ~new_P3_U6855 | ~new_P3_U6854;
  assign n2274 = P3_DATAO_REG_31_ & new_P3_U6759;
  assign n2270 = ~new_P3_U4001 | ~new_P3_U6850;
  assign n2266 = ~new_P3_U4000 | ~new_P3_U6847;
  assign n2262 = ~new_P3_U3999 | ~new_P3_U6844;
  assign n2258 = ~new_P3_U3998 | ~new_P3_U6841;
  assign n2254 = ~new_P3_U3997 | ~new_P3_U6838;
  assign n2250 = ~new_P3_U3996 | ~new_P3_U6835;
  assign n2246 = ~new_P3_U3995 | ~new_P3_U6832;
  assign n2242 = ~new_P3_U3994 | ~new_P3_U6829;
  assign n2238 = ~new_P3_U3993 | ~new_P3_U6826;
  assign n2234 = ~new_P3_U3992 | ~new_P3_U6823;
  assign n2230 = ~new_P3_U3991 | ~new_P3_U6820;
  assign n2226 = ~new_P3_U3990 | ~new_P3_U6817;
  assign n2222 = ~new_P3_U3989 | ~new_P3_U6814;
  assign n2218 = ~new_P3_U3988 | ~new_P3_U6811;
  assign n2214 = ~new_P3_U3987 | ~new_P3_U6808;
  assign n2210 = ~new_P3_U6807 | ~new_P3_U6806 | ~new_P3_U6805;
  assign n2206 = ~new_P3_U6804 | ~new_P3_U6803 | ~new_P3_U6802;
  assign n2202 = ~new_P3_U6801 | ~new_P3_U6800 | ~new_P3_U6799;
  assign n2198 = ~new_P3_U6798 | ~new_P3_U6797 | ~new_P3_U6796;
  assign n2194 = ~new_P3_U6795 | ~new_P3_U6794 | ~new_P3_U6793;
  assign n2190 = ~new_P3_U6792 | ~new_P3_U6791 | ~new_P3_U6790;
  assign n2186 = ~new_P3_U6789 | ~new_P3_U6788 | ~new_P3_U6787;
  assign n2182 = ~new_P3_U6786 | ~new_P3_U6785 | ~new_P3_U6784;
  assign n2178 = ~new_P3_U6783 | ~new_P3_U6782 | ~new_P3_U6781;
  assign n2174 = ~new_P3_U6780 | ~new_P3_U6779 | ~new_P3_U6778;
  assign n2170 = ~new_P3_U6777 | ~new_P3_U6776 | ~new_P3_U6775;
  assign n2166 = ~new_P3_U6774 | ~new_P3_U6773 | ~new_P3_U6772;
  assign n2162 = ~new_P3_U6771 | ~new_P3_U6770 | ~new_P3_U6769;
  assign n2158 = ~new_P3_U6768 | ~new_P3_U6767 | ~new_P3_U6766;
  assign n2154 = ~new_P3_U6765 | ~new_P3_U6764 | ~new_P3_U6763;
  assign n2150 = ~new_P3_U6762 | ~new_P3_U6761 | ~new_P3_U6760;
  assign n2145 = ~new_P3_U6756 | ~new_P3_U6755 | ~new_P3_U6754;
  assign n2140 = ~new_P3_U6753 | ~new_P3_U6752 | ~new_P3_U6751;
  assign n2135 = ~new_P3_U6750 | ~new_P3_U6749 | ~new_P3_U6748;
  assign n2130 = ~new_P3_U6747 | ~new_P3_U6746 | ~new_P3_U6745;
  assign n2125 = ~new_P3_U6744 | ~new_P3_U6743 | ~new_P3_U6742;
  assign n2120 = ~new_P3_U6741 | ~new_P3_U6740 | ~new_P3_U6739;
  assign n2115 = ~new_P3_U6738 | ~new_P3_U6737 | ~new_P3_U6736;
  assign n2110 = ~new_P3_U6735 | ~new_P3_U6734 | ~new_P3_U6733;
  assign n2105 = ~new_P3_U6732 | ~new_P3_U6731 | ~new_P3_U6730;
  assign n2100 = ~new_P3_U6729 | ~new_P3_U6728 | ~new_P3_U6727;
  assign n2095 = ~new_P3_U6726 | ~new_P3_U6725 | ~new_P3_U6724;
  assign n2090 = ~new_P3_U6723 | ~new_P3_U6722 | ~new_P3_U6721;
  assign n2085 = ~new_P3_U6720 | ~new_P3_U6719 | ~new_P3_U6718;
  assign n2080 = ~new_P3_U6717 | ~new_P3_U6716 | ~new_P3_U6715;
  assign n2075 = ~new_P3_U6714 | ~new_P3_U6713 | ~new_P3_U6712;
  assign n2070 = ~new_P3_U6711 | ~new_P3_U6710 | ~new_P3_U6709;
  assign n2065 = ~new_P3_U6708 | ~new_P3_U6707 | ~new_P3_U6706;
  assign n2060 = ~new_P3_U6705 | ~new_P3_U6704 | ~new_P3_U6703;
  assign n2055 = ~new_P3_U6702 | ~new_P3_U6701 | ~new_P3_U6700;
  assign n2050 = ~new_P3_U6699 | ~new_P3_U6698 | ~new_P3_U6697;
  assign n2045 = ~new_P3_U6696 | ~new_P3_U6695 | ~new_P3_U6694;
  assign n2040 = ~new_P3_U6693 | ~new_P3_U6692 | ~new_P3_U6691;
  assign n2035 = ~new_P3_U6690 | ~new_P3_U6689 | ~new_P3_U6688;
  assign n2030 = ~new_P3_U6687 | ~new_P3_U6686 | ~new_P3_U6685;
  assign n2025 = ~new_P3_U6684 | ~new_P3_U6683 | ~new_P3_U6682;
  assign n2020 = ~new_P3_U6681 | ~new_P3_U6680 | ~new_P3_U6679;
  assign n2015 = ~new_P3_U6678 | ~new_P3_U6677 | ~new_P3_U6676;
  assign n2010 = ~new_P3_U6675 | ~new_P3_U6674 | ~new_P3_U6673;
  assign n2005 = ~new_P3_U6672 | ~new_P3_U6671 | ~new_P3_U6670;
  assign n2000 = ~new_P3_U6669 | ~new_P3_U6668 | ~new_P3_U6667;
  assign n1995 = ~new_P3_U6666 | ~new_P3_U6665 | ~new_P3_U6664;
  assign n1990 = ~new_P3_U3985 | ~new_P3_U6653 | ~new_P3_U6655 | ~new_P3_U6656 | ~new_P3_U6654;
  assign n1985 = ~new_P3_U3984 | ~new_P3_U6645 | ~new_P3_U6646 | ~new_P3_U6648 | ~new_P3_U6647;
  assign n1980 = ~new_P3_U3983 | ~new_P3_U6637 | ~new_P3_U6638 | ~new_P3_U6640 | ~new_P3_U6639;
  assign n1975 = ~new_P3_U3982 | ~new_P3_U6629 | ~new_P3_U6630 | ~new_P3_U6632 | ~new_P3_U6631;
  assign n1970 = ~new_P3_U3981 | ~new_P3_U6623 | ~new_P3_U6621 | ~new_P3_U6622 | ~new_P3_U6624;
  assign n1965 = ~new_P3_U3980 | ~new_P3_U6615 | ~new_P3_U6613 | ~new_P3_U6614 | ~new_P3_U6616;
  assign n1960 = ~new_P3_U3979 | ~new_P3_U6607 | ~new_P3_U6605 | ~new_P3_U6606 | ~new_P3_U6608;
  assign n1955 = ~new_P3_U3978 | ~new_P3_U6599 | ~new_P3_U6597 | ~new_P3_U6598 | ~new_P3_U6600;
  assign n1950 = ~new_P3_U3977 | ~new_P3_U6591 | ~new_P3_U6592 | ~new_P3_U6590 | ~new_P3_U6589;
  assign n1945 = ~new_P3_U3976 | ~new_P3_U6583 | ~new_P3_U6584 | ~new_P3_U6582 | ~new_P3_U6581;
  assign n1940 = ~new_P3_U6576 | ~new_P3_U3975 | ~new_P3_U6575 | ~new_P3_U6574 | ~new_P3_U6573;
  assign n1935 = ~new_P3_U6568 | ~new_P3_U3974 | ~new_P3_U6567 | ~new_P3_U6566 | ~new_P3_U6565;
  assign n1930 = ~new_P3_U3973 | ~new_P3_U6560 | ~new_P3_U6559 | ~new_P3_U6558 | ~new_P3_U6557;
  assign n1925 = ~new_P3_U3972 | ~new_P3_U6552 | ~new_P3_U6551 | ~new_P3_U6550 | ~new_P3_U6549;
  assign n1920 = ~new_P3_U3971 | ~new_P3_U6544 | ~new_P3_U6543 | ~new_P3_U6542 | ~new_P3_U6541;
  assign n1915 = ~new_P3_U3970 | ~new_P3_U6536 | ~new_P3_U6535 | ~new_P3_U6534 | ~new_P3_U6533;
  assign n1910 = ~new_P3_U3969 | ~new_P3_U6527 | ~new_P3_U6528 | ~new_P3_U6526 | ~new_P3_U6525;
  assign n1905 = ~new_P3_U3968 | ~new_P3_U6519 | ~new_P3_U6520 | ~new_P3_U6518 | ~new_P3_U6517;
  assign n1900 = ~new_P3_U3967 | ~new_P3_U6511 | ~new_P3_U6512 | ~new_P3_U6510 | ~new_P3_U6509;
  assign n1895 = ~new_P3_U3966 | ~new_P3_U6503 | ~new_P3_U6504 | ~new_P3_U6502 | ~new_P3_U6501;
  assign n1890 = ~new_P3_U3965 | ~new_P3_U6496 | ~new_P3_U6495 | ~new_P3_U6494 | ~new_P3_U6493;
  assign n1885 = ~new_P3_U3964 | ~new_P3_U6488 | ~new_P3_U6487 | ~new_P3_U6486 | ~new_P3_U6485;
  assign n1880 = ~new_P3_U3963 | ~new_P3_U6479 | ~new_P3_U6480 | ~new_P3_U6478 | ~new_P3_U6477;
  assign n1875 = ~new_P3_U3962 | ~new_P3_U6471 | ~new_P3_U6472 | ~new_P3_U6470 | ~new_P3_U6469;
  assign n1870 = ~new_P3_U3961 | ~new_P3_U6463 | ~new_P3_U6464 | ~new_P3_U6462 | ~new_P3_U6461;
  assign n1865 = ~new_P3_U3960 | ~new_P3_U6455 | ~new_P3_U6456 | ~new_P3_U6454 | ~new_P3_U6453;
  assign n1860 = ~new_P3_U3959 | ~new_P3_U6447 | ~new_P3_U6448 | ~new_P3_U6446 | ~new_P3_U6445;
  assign n1855 = ~new_P3_U3958 | ~new_P3_U6440 | ~new_P3_U6439 | ~new_P3_U6438 | ~new_P3_U6437;
  assign n1850 = ~new_P3_U3957 | ~new_P3_U6429 | ~new_P3_U6430 | ~new_P3_U6432 | ~new_P3_U6431;
  assign n1845 = ~new_P3_U3956 | ~new_P3_U6421 | ~new_P3_U6422 | ~new_P3_U6424 | ~new_P3_U6423;
  assign n1840 = ~new_P3_U3955 | ~new_P3_U6413 | ~new_P3_U6414 | ~new_P3_U6416 | ~new_P3_U6415;
  assign n1835 = ~new_P3_U3954 | ~new_P3_U6405 | ~new_P3_U6406 | ~new_P3_U6408 | ~new_P3_U6407;
  assign n1830 = new_P3_U6396 & new_P3_U7906;
  assign n1825 = ~new_P3_U6374 | ~new_P3_U6375 | ~new_P3_U6373;
  assign n1820 = ~new_P3_U6350 | ~new_P3_U6351 | ~new_P3_U6349;
  assign n1815 = ~new_P3_U6326 | ~new_P3_U6327 | ~new_P3_U6325;
  assign n1810 = ~new_P3_U6302 | ~new_P3_U6303 | ~new_P3_U6301;
  assign n1805 = ~new_P3_U6278 | ~new_P3_U6279 | ~new_P3_U6277;
  assign n1800 = ~new_P3_U3893 | ~new_P3_U6254;
  assign n1795 = ~new_P3_U3883 | ~new_P3_U6230;
  assign n1790 = ~new_P3_U3873 | ~new_P3_U6206;
  assign n1785 = ~new_P3_U3863 | ~new_P3_U6182;
  assign n1780 = ~new_P3_U3853 | ~new_P3_U6158;
  assign n1775 = ~new_P3_U3845 | ~new_P3_U6134;
  assign n1770 = ~new_P3_U6110 | ~new_P3_U6111 | ~new_P3_U6109;
  assign n1765 = ~new_P3_U6086 | ~new_P3_U6087 | ~new_P3_U6085;
  assign n1760 = ~new_P3_U6062 | ~new_P3_U6063 | ~new_P3_U6061;
  assign n1755 = ~new_P3_U6038 | ~new_P3_U6039 | ~new_P3_U6037;
  assign n1750 = ~new_P3_U3811 | ~new_P3_U6014;
  assign n1745 = ~new_P3_U3803 | ~new_P3_U5990;
  assign n1740 = ~new_P3_U5966 | ~new_P3_U5967 | ~new_P3_U5965;
  assign n1735 = ~new_P3_U5942 | ~new_P3_U5943 | ~new_P3_U5941;
  assign n1730 = ~new_P3_U5918 | ~new_P3_U5919 | ~new_P3_U5917;
  assign n1725 = ~new_P3_U5894 | ~new_P3_U5895 | ~new_P3_U5893;
  assign n1720 = ~new_P3_U5870 | ~new_P3_U5871 | ~new_P3_U5869;
  assign n1715 = ~new_P3_U5846 | ~new_P3_U5847 | ~new_P3_U5845;
  assign n1710 = ~new_P3_U5822 | ~new_P3_U5823 | ~new_P3_U5821;
  assign n1705 = ~new_P3_U5798 | ~new_P3_U5799 | ~new_P3_U5797;
  assign n1700 = ~new_P3_U5774 | ~new_P3_U5775 | ~new_P3_U5773;
  assign n1695 = ~new_P3_U5750 | ~new_P3_U5751 | ~new_P3_U5749;
  assign n1690 = ~new_P3_U5726 | ~new_P3_U5727 | ~new_P3_U5725;
  assign n1685 = ~new_P3_U5702 | ~new_P3_U5703 | ~new_P3_U5701;
  assign n1680 = ~new_P3_U5678 | ~new_P3_U5679 | ~new_P3_U5677;
  assign n1675 = ~new_P3_U5655 | ~new_P3_U5654 | ~new_P3_U5653;
  assign n1670 = ~new_P3_U5616 | ~new_P3_U5615;
  assign n1665 = ~new_P3_U5610 | ~new_P3_U5609;
  assign n1660 = ~new_P3_U5599 | ~new_P3_U5598;
  assign n1655 = ~new_P3_U5591 | ~new_P3_U5590;
  assign n1650 = P3_INSTQUEUEWR_ADDR_REG_4_ & new_P3_U5579;
  assign n1620 = ~new_P3_U3651 | ~new_P3_U5482;
  assign n1615 = ~new_P3_U3649 | ~new_P3_U5477;
  assign n1610 = ~new_P3_U3647 | ~new_P3_U5472;
  assign n1605 = ~new_P3_U3645 | ~new_P3_U5467;
  assign n1600 = ~new_P3_U3643 | ~new_P3_U5462;
  assign n1595 = ~new_P3_U3641 | ~new_P3_U5457;
  assign n1590 = ~new_P3_U3639 | ~new_P3_U5452;
  assign n1585 = ~new_P3_U3637 | ~new_P3_U5447;
  assign n1580 = ~new_P3_U3633 | ~new_P3_U5432;
  assign n1575 = ~new_P3_U3631 | ~new_P3_U5427;
  assign n1570 = ~new_P3_U3629 | ~new_P3_U5422;
  assign n1565 = ~new_P3_U3627 | ~new_P3_U5417;
  assign n1560 = ~new_P3_U3625 | ~new_P3_U5412;
  assign n1555 = ~new_P3_U3623 | ~new_P3_U5407;
  assign n1550 = ~new_P3_U3621 | ~new_P3_U5402;
  assign n1545 = ~new_P3_U3619 | ~new_P3_U5397;
  assign n1540 = ~new_P3_U3615 | ~new_P3_U5381;
  assign n1535 = ~new_P3_U3613 | ~new_P3_U5376;
  assign n1530 = ~new_P3_U3611 | ~new_P3_U5371;
  assign n1525 = ~new_P3_U3609 | ~new_P3_U5366;
  assign n1520 = ~new_P3_U3607 | ~new_P3_U5361;
  assign n1515 = ~new_P3_U3605 | ~new_P3_U5356;
  assign n1510 = ~new_P3_U3603 | ~new_P3_U5351;
  assign n1505 = ~new_P3_U3601 | ~new_P3_U5346;
  assign n1500 = ~new_P3_U3598 | ~new_P3_U5330;
  assign n1495 = ~new_P3_U3596 | ~new_P3_U5325;
  assign n1490 = ~new_P3_U3594 | ~new_P3_U5320;
  assign n1485 = ~new_P3_U3592 | ~new_P3_U5315;
  assign n1480 = ~new_P3_U3590 | ~new_P3_U5310;
  assign n1475 = ~new_P3_U3588 | ~new_P3_U5305;
  assign n1470 = ~new_P3_U3586 | ~new_P3_U5300;
  assign n1465 = ~new_P3_U3584 | ~new_P3_U5295;
  assign n1460 = ~new_P3_U3580 | ~new_P3_U5279;
  assign n1455 = ~new_P3_U3578 | ~new_P3_U5274;
  assign n1450 = ~new_P3_U3576 | ~new_P3_U5269;
  assign n1445 = ~new_P3_U3574 | ~new_P3_U5264;
  assign n1440 = ~new_P3_U3572 | ~new_P3_U5259;
  assign n1435 = ~new_P3_U3570 | ~new_P3_U5254;
  assign n1430 = ~new_P3_U3568 | ~new_P3_U5249;
  assign n1425 = ~new_P3_U3566 | ~new_P3_U5244;
  assign n1420 = ~new_P3_U5228 | ~new_P3_U5229 | ~new_P3_U3562;
  assign n1415 = ~new_P3_U5223 | ~new_P3_U5224 | ~new_P3_U3560;
  assign n1410 = ~new_P3_U5218 | ~new_P3_U5219 | ~new_P3_U3558;
  assign n1405 = ~new_P3_U5213 | ~new_P3_U5214 | ~new_P3_U3556;
  assign n1400 = ~new_P3_U5208 | ~new_P3_U5209 | ~new_P3_U3554;
  assign n1395 = ~new_P3_U5203 | ~new_P3_U5204 | ~new_P3_U3552;
  assign n1390 = ~new_P3_U5198 | ~new_P3_U5199 | ~new_P3_U3550;
  assign n1385 = ~new_P3_U5193 | ~new_P3_U5194 | ~new_P3_U3548;
  assign n1380 = ~new_P3_U5176 | ~new_P3_U5177 | ~new_P3_U3544;
  assign n1375 = ~new_P3_U5171 | ~new_P3_U5172 | ~new_P3_U3542;
  assign n1370 = ~new_P3_U5166 | ~new_P3_U5167 | ~new_P3_U3540;
  assign n1365 = ~new_P3_U5161 | ~new_P3_U5162 | ~new_P3_U3538;
  assign n1360 = ~new_P3_U5156 | ~new_P3_U5157 | ~new_P3_U3536;
  assign n1355 = ~new_P3_U5151 | ~new_P3_U5152 | ~new_P3_U3534;
  assign n1350 = ~new_P3_U5146 | ~new_P3_U5147 | ~new_P3_U3532;
  assign n1345 = ~new_P3_U5141 | ~new_P3_U5142 | ~new_P3_U3530;
  assign n1340 = ~new_P3_U5124 | ~new_P3_U5125 | ~new_P3_U3526;
  assign n1335 = ~new_P3_U5119 | ~new_P3_U5120 | ~new_P3_U3524;
  assign n1330 = ~new_P3_U5114 | ~new_P3_U5115 | ~new_P3_U3522;
  assign n1325 = ~new_P3_U5109 | ~new_P3_U5110 | ~new_P3_U3520;
  assign n1320 = ~new_P3_U5104 | ~new_P3_U5105 | ~new_P3_U3518;
  assign n1315 = ~new_P3_U5099 | ~new_P3_U5100 | ~new_P3_U3516;
  assign n1310 = ~new_P3_U5094 | ~new_P3_U5095 | ~new_P3_U3514;
  assign n1305 = ~new_P3_U5089 | ~new_P3_U5090 | ~new_P3_U3512;
  assign n1300 = ~new_P3_U5075 | ~new_P3_U5076 | ~new_P3_U3509;
  assign n1295 = ~new_P3_U5070 | ~new_P3_U5071 | ~new_P3_U3507;
  assign n1290 = ~new_P3_U5065 | ~new_P3_U5066 | ~new_P3_U3505;
  assign n1285 = ~new_P3_U5060 | ~new_P3_U5061 | ~new_P3_U3503;
  assign n1280 = ~new_P3_U5055 | ~new_P3_U5056 | ~new_P3_U3501;
  assign n1275 = ~new_P3_U5050 | ~new_P3_U5051 | ~new_P3_U3499;
  assign n1270 = ~new_P3_U5045 | ~new_P3_U5046 | ~new_P3_U3497;
  assign n1265 = ~new_P3_U5040 | ~new_P3_U5041 | ~new_P3_U3495;
  assign n1260 = ~new_P3_U5024 | ~new_P3_U5025 | ~new_P3_U3492;
  assign n1255 = ~new_P3_U5019 | ~new_P3_U5020 | ~new_P3_U3490;
  assign n1250 = ~new_P3_U5014 | ~new_P3_U5015 | ~new_P3_U3488;
  assign n1245 = ~new_P3_U5009 | ~new_P3_U5010 | ~new_P3_U3486;
  assign n1240 = ~new_P3_U5004 | ~new_P3_U5005 | ~new_P3_U3484;
  assign n1235 = ~new_P3_U4999 | ~new_P3_U5000 | ~new_P3_U3482;
  assign n1230 = ~new_P3_U4994 | ~new_P3_U4995 | ~new_P3_U3480;
  assign n1225 = ~new_P3_U4989 | ~new_P3_U4990 | ~new_P3_U3478;
  assign n1220 = ~new_P3_U4972 | ~new_P3_U4973 | ~new_P3_U3474;
  assign n1215 = ~new_P3_U4967 | ~new_P3_U4968 | ~new_P3_U3472;
  assign n1210 = ~new_P3_U4962 | ~new_P3_U4963 | ~new_P3_U3470;
  assign n1205 = ~new_P3_U4957 | ~new_P3_U4958 | ~new_P3_U3468;
  assign n1200 = ~new_P3_U4952 | ~new_P3_U4953 | ~new_P3_U3466;
  assign n1195 = ~new_P3_U4947 | ~new_P3_U4948 | ~new_P3_U3464;
  assign n1190 = ~new_P3_U4942 | ~new_P3_U4943 | ~new_P3_U3462;
  assign n1185 = ~new_P3_U4937 | ~new_P3_U4938 | ~new_P3_U3460;
  assign n1180 = ~new_P3_U4920 | ~new_P3_U4921 | ~new_P3_U3456;
  assign n1175 = ~new_P3_U4915 | ~new_P3_U4916 | ~new_P3_U3454;
  assign n1170 = ~new_P3_U4910 | ~new_P3_U4911 | ~new_P3_U3452;
  assign n1165 = ~new_P3_U4905 | ~new_P3_U4906 | ~new_P3_U3450;
  assign n1160 = ~new_P3_U4900 | ~new_P3_U4901 | ~new_P3_U3448;
  assign n1155 = ~new_P3_U4895 | ~new_P3_U4896 | ~new_P3_U3446;
  assign n1150 = ~new_P3_U4890 | ~new_P3_U4891 | ~new_P3_U3444;
  assign n1145 = ~new_P3_U4885 | ~new_P3_U4886 | ~new_P3_U3442;
  assign n1140 = ~new_P3_U4868 | ~new_P3_U4869 | ~new_P3_U3439;
  assign n1135 = ~new_P3_U4863 | ~new_P3_U4864 | ~new_P3_U3437;
  assign n1130 = ~new_P3_U4858 | ~new_P3_U4859 | ~new_P3_U3435;
  assign n1125 = ~new_P3_U4853 | ~new_P3_U4854 | ~new_P3_U3433;
  assign n1120 = ~new_P3_U4848 | ~new_P3_U4849 | ~new_P3_U3431;
  assign n1115 = ~new_P3_U4843 | ~new_P3_U4844 | ~new_P3_U3429;
  assign n1110 = ~new_P3_U4838 | ~new_P3_U4839 | ~new_P3_U3427;
  assign n1105 = ~new_P3_U4833 | ~new_P3_U4834 | ~new_P3_U3425;
  assign n1100 = ~new_P3_U4817 | ~new_P3_U4818 | ~new_P3_U3421;
  assign n1095 = ~new_P3_U4812 | ~new_P3_U4813 | ~new_P3_U3419;
  assign n1090 = ~new_P3_U4807 | ~new_P3_U4808 | ~new_P3_U3417;
  assign n1085 = ~new_P3_U4802 | ~new_P3_U4803 | ~new_P3_U3415;
  assign n1080 = ~new_P3_U4797 | ~new_P3_U4798 | ~new_P3_U3413;
  assign n1075 = ~new_P3_U4792 | ~new_P3_U4793 | ~new_P3_U3411;
  assign n1070 = ~new_P3_U4787 | ~new_P3_U4788 | ~new_P3_U3409;
  assign n1065 = ~new_P3_U4782 | ~new_P3_U4783 | ~new_P3_U3407;
  assign n1060 = ~new_P3_U4765 | ~new_P3_U4766 | ~new_P3_U3403;
  assign n1055 = ~new_P3_U4760 | ~new_P3_U4761 | ~new_P3_U3401;
  assign n1050 = ~new_P3_U4755 | ~new_P3_U4756 | ~new_P3_U3399;
  assign n1045 = ~new_P3_U4750 | ~new_P3_U4751 | ~new_P3_U3397;
  assign n1040 = ~new_P3_U4745 | ~new_P3_U4746 | ~new_P3_U3395;
  assign n1035 = ~new_P3_U4740 | ~new_P3_U4741 | ~new_P3_U3393;
  assign n1030 = ~new_P3_U4735 | ~new_P3_U4736 | ~new_P3_U3391;
  assign n1025 = ~new_P3_U4730 | ~new_P3_U4731 | ~new_P3_U3389;
  assign n1020 = ~new_P3_U4713 | ~new_P3_U4714 | ~new_P3_U3385;
  assign n1015 = ~new_P3_U4708 | ~new_P3_U4709 | ~new_P3_U3383;
  assign n1010 = ~new_P3_U4703 | ~new_P3_U4704 | ~new_P3_U3381;
  assign n1005 = ~new_P3_U4698 | ~new_P3_U4699 | ~new_P3_U3379;
  assign n1000 = ~new_P3_U4693 | ~new_P3_U4694 | ~new_P3_U3377;
  assign n995 = ~new_P3_U4688 | ~new_P3_U4689 | ~new_P3_U3375;
  assign n990 = ~new_P3_U4683 | ~new_P3_U4684 | ~new_P3_U3373;
  assign n985 = ~new_P3_U4678 | ~new_P3_U4679 | ~new_P3_U3371;
  assign n980 = ~new_P3_U3367 | ~new_P3_U7959 | ~new_P3_U7958;
  assign n975 = ~new_P3_U4329 | ~new_P3_U4634 | ~new_P3_U4636 | ~new_P3_U4635;
  assign n970 = ~new_P3_U3363 | ~new_P3_U4632;
  assign n960 = P3_DATAWIDTH_REG_31_ & new_P3_U7937;
  assign n955 = P3_DATAWIDTH_REG_30_ & new_P3_U7937;
  assign n950 = P3_DATAWIDTH_REG_29_ & new_P3_U7937;
  assign n945 = P3_DATAWIDTH_REG_28_ & new_P3_U7937;
  assign n940 = P3_DATAWIDTH_REG_27_ & new_P3_U7937;
  assign n935 = P3_DATAWIDTH_REG_26_ & new_P3_U7937;
  assign n930 = P3_DATAWIDTH_REG_25_ & new_P3_U7937;
  assign n925 = P3_DATAWIDTH_REG_24_ & new_P3_U7937;
  assign n920 = P3_DATAWIDTH_REG_23_ & new_P3_U7937;
  assign n915 = P3_DATAWIDTH_REG_22_ & new_P3_U7937;
  assign n910 = P3_DATAWIDTH_REG_21_ & new_P3_U7937;
  assign n905 = P3_DATAWIDTH_REG_20_ & new_P3_U7937;
  assign n900 = P3_DATAWIDTH_REG_19_ & new_P3_U7937;
  assign n895 = P3_DATAWIDTH_REG_18_ & new_P3_U7937;
  assign n890 = P3_DATAWIDTH_REG_17_ & new_P3_U7937;
  assign n885 = P3_DATAWIDTH_REG_16_ & new_P3_U7937;
  assign n880 = P3_DATAWIDTH_REG_15_ & new_P3_U7937;
  assign n875 = P3_DATAWIDTH_REG_14_ & new_P3_U7937;
  assign n870 = P3_DATAWIDTH_REG_13_ & new_P3_U7937;
  assign n865 = P3_DATAWIDTH_REG_12_ & new_P3_U7937;
  assign n860 = P3_DATAWIDTH_REG_11_ & new_P3_U7937;
  assign n855 = P3_DATAWIDTH_REG_10_ & new_P3_U7937;
  assign n850 = P3_DATAWIDTH_REG_9_ & new_P3_U7937;
  assign n845 = P3_DATAWIDTH_REG_8_ & new_P3_U7937;
  assign n840 = P3_DATAWIDTH_REG_7_ & new_P3_U7937;
  assign n835 = P3_DATAWIDTH_REG_6_ & new_P3_U7937;
  assign n830 = P3_DATAWIDTH_REG_5_ & new_P3_U7937;
  assign n825 = P3_DATAWIDTH_REG_4_ & new_P3_U7937;
  assign n820 = P3_DATAWIDTH_REG_3_ & new_P3_U7937;
  assign n815 = P3_DATAWIDTH_REG_2_ & new_P3_U7937;
  assign n800 = ~new_P3_U4463 | ~new_P3_U7934 | ~new_P3_U7933;
  assign n795 = ~new_P3_U3311 | ~new_P3_U7932 | ~new_P3_U7931;
  assign n790 = ~new_P3_U3310 | ~new_P3_U4457;
  assign n785 = ~new_P3_U4444 | ~new_P3_U4443 | ~new_P3_U4442;
  assign n780 = ~new_P3_U4441 | ~new_P3_U4440 | ~new_P3_U4439;
  assign n775 = ~new_P3_U4438 | ~new_P3_U4437 | ~new_P3_U4436;
  assign n770 = ~new_P3_U4435 | ~new_P3_U4434 | ~new_P3_U4433;
  assign n765 = ~new_P3_U4432 | ~new_P3_U4431 | ~new_P3_U4430;
  assign n760 = ~new_P3_U4429 | ~new_P3_U4428 | ~new_P3_U4427;
  assign n755 = ~new_P3_U4426 | ~new_P3_U4425 | ~new_P3_U4424;
  assign n750 = ~new_P3_U4423 | ~new_P3_U4422 | ~new_P3_U4421;
  assign n745 = ~new_P3_U4420 | ~new_P3_U4419 | ~new_P3_U4418;
  assign n740 = ~new_P3_U4417 | ~new_P3_U4416 | ~new_P3_U4415;
  assign n735 = ~new_P3_U4414 | ~new_P3_U4413 | ~new_P3_U4412;
  assign n730 = ~new_P3_U4411 | ~new_P3_U4410 | ~new_P3_U4409;
  assign n725 = ~new_P3_U4408 | ~new_P3_U4407 | ~new_P3_U4406;
  assign n720 = ~new_P3_U4405 | ~new_P3_U4404 | ~new_P3_U4403;
  assign n715 = ~new_P3_U4402 | ~new_P3_U4401 | ~new_P3_U4400;
  assign n710 = ~new_P3_U4399 | ~new_P3_U4398 | ~new_P3_U4397;
  assign n705 = ~new_P3_U4396 | ~new_P3_U4395 | ~new_P3_U4394;
  assign n700 = ~new_P3_U4393 | ~new_P3_U4392 | ~new_P3_U4391;
  assign n695 = ~new_P3_U4390 | ~new_P3_U4389 | ~new_P3_U4388;
  assign n690 = ~new_P3_U4387 | ~new_P3_U4386 | ~new_P3_U4385;
  assign n685 = ~new_P3_U4384 | ~new_P3_U4383 | ~new_P3_U4382;
  assign n680 = ~new_P3_U4381 | ~new_P3_U4380 | ~new_P3_U4379;
  assign n675 = ~new_P3_U4378 | ~new_P3_U4377 | ~new_P3_U4376;
  assign n670 = ~new_P3_U4375 | ~new_P3_U4374 | ~new_P3_U4373;
  assign n665 = ~new_P3_U4372 | ~new_P3_U4371 | ~new_P3_U4370;
  assign n660 = ~new_P3_U4369 | ~new_P3_U4368 | ~new_P3_U4367;
  assign n655 = ~new_P3_U4366 | ~new_P3_U4365 | ~new_P3_U4364;
  assign n650 = ~new_P3_U4363 | ~new_P3_U4362 | ~new_P3_U4361;
  assign n645 = ~new_P3_U4360 | ~new_P3_U4359 | ~new_P3_U4358;
  assign n640 = ~new_P3_U4357 | ~new_P3_U4356 | ~new_P3_U4355;
  assign new_P3_U3062 = ~new_P3_U4244 | ~new_P3_U4245 | ~new_P3_U4247 | ~new_P3_U4246;
  assign new_P3_U3063 = ~new_P3_U4240 | ~new_P3_U4241 | ~new_P3_U4243 | ~new_P3_U4242;
  assign new_P3_U3064 = ~new_P3_U4236 | ~new_P3_U4237 | ~new_P3_U4239 | ~new_P3_U4238;
  assign new_P3_U3065 = ~new_P3_U4232 | ~new_P3_U4233 | ~new_P3_U4235 | ~new_P3_U4234;
  assign new_P3_U3066 = ~new_P3_U4228 | ~new_P3_U4229 | ~new_P3_U4231 | ~new_P3_U4230;
  assign new_P3_U3067 = ~new_P3_U4224 | ~new_P3_U4225 | ~new_P3_U4227 | ~new_P3_U4226;
  assign new_P3_U3068 = ~new_P3_U4220 | ~new_P3_U4221 | ~new_P3_U4223 | ~new_P3_U4222;
  assign new_P3_U3069 = ~new_P3_U4216 | ~new_P3_U4217 | ~new_P3_U4219 | ~new_P3_U4218;
  assign new_P3_U3070 = ~new_P3_U2457 | ~new_P3_U4642;
  assign new_P3_U3071 = ~new_P3_U2459 | ~new_P3_U4642;
  assign new_P3_U3072 = ~new_P3_U2458 | ~new_P3_U4642;
  assign new_P3_U3073 = ~new_P3_U2460 | ~new_P3_U4642;
  assign new_P3_U3074 = ~new_P3_U3343 | ~new_P3_U3344 | ~new_P3_U3347 | ~new_P3_U3346 | ~new_P3_U3345;
  assign new_P3_U3075 = ~P3_REQUESTPENDING_REG;
  assign new_P3_U3076 = ~P3_STATE_REG_1_;
  assign new_P3_U3077 = ~P3_STATE_REG_1_ | ~new_P3_U3085;
  assign new_P3_U3078 = ~new_P3_U4308 | ~new_P3_U3079;
  assign new_P3_U3079 = ~P3_STATE_REG_2_;
  assign new_P3_U3080 = ~P3_STATE_REG_2_ | ~new_P3_U4308;
  assign new_P3_U3081 = ~P3_REIP_REG_1_;
  assign new_P3_U3082 = ~P3_STATE_REG_1_ | ~new_P3_U3079;
  assign new_P3_U3083 = P3_STATE_REG_1_ | P3_STATE_REG_2_;
  assign new_P3_U3084 = ~HOLD;
  assign new_P3_U3085 = ~P3_STATE_REG_0_;
  assign new_P3_U3086 = ~P3_STATE_REG_0_ | ~new_P3_U3087;
  assign new_P3_U3087 = ~P3_REQUESTPENDING_REG | ~new_P3_U3084;
  assign new_P3_U3088 = HOLD | P3_REQUESTPENDING_REG;
  assign new_P3_U3089 = ~P3_STATE2_REG_1_;
  assign new_P3_U3090 = ~P3_STATE2_REG_2_;
  assign new_P3_U3091 = P3_INSTQUEUERD_ADDR_REG_1_ | P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_U3092 = ~new_P3_U4467 | ~new_P3_U3097;
  assign new_P3_U3093 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_U3094 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_U3095 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_U3096 = ~new_P3_U4332 | ~new_P3_U3097;
  assign new_P3_U3097 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_U3098 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U3100;
  assign new_P3_U3099 = ~new_P3_U4470 | ~new_P3_U4332;
  assign new_P3_U3100 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_U3101 = ~new_P3_U3338 | ~new_P3_U3339 | ~new_P3_U3342 | ~new_P3_U3341 | ~new_P3_U3340;
  assign new_P3_U3102 = ~new_P3_U3323 | ~new_P3_U3324 | ~new_P3_U3327 | ~new_P3_U3326 | ~new_P3_U3325;
  assign new_P3_U3103 = ~new_P3_U3074 | ~new_P3_U3110;
  assign new_P3_U3104 = ~new_P3_U3318 | ~new_P3_U3319 | ~new_P3_U3322 | ~new_P3_U3321 | ~new_P3_U3320;
  assign new_P3_U3105 = ~new_P3_U4466 | ~new_P3_U3085;
  assign new_P3_U3106 = ~new_P3_U4293 | ~new_P3_U2630;
  assign new_P3_U3107 = ~new_P3_U3328 | ~new_P3_U3329 | ~new_P3_U3332 | ~new_P3_U3331 | ~new_P3_U3330;
  assign new_P3_U3108 = ~new_P3_U3313 | ~new_P3_U3314 | ~new_P3_U3317 | ~new_P3_U3316 | ~new_P3_U3315;
  assign new_P3_U3109 = ~new_P3_U2353 | ~new_P3_U4488;
  assign new_P3_U3110 = ~new_P3_U3348 | ~new_P3_U3349 | ~new_P3_U3352 | ~new_P3_U3351 | ~new_P3_U3350;
  assign new_P3_U3111 = ~new_P3_U3104 | ~new_P3_U3108;
  assign new_P3_U3112 = ~new_P3_U4505 | ~new_P3_U3108;
  assign new_P3_U3113 = ~new_P3_U4607 | ~new_P3_U3110;
  assign new_P3_U3114 = ~new_P3_U4488 | ~new_P3_U4505;
  assign new_P3_U3115 = ~new_P3_U2451 | ~new_P3_U4297;
  assign new_P3_U3116 = ~new_P3_U2452 | ~new_P3_U4297;
  assign new_P3_U3117 = ~new_P3_U2452 | ~new_P3_U4296;
  assign new_P3_U3118 = ~new_P3_U4488 | ~new_P3_U3104;
  assign new_P3_U3119 = ~new_P3_U3356 | ~new_P3_U2353;
  assign new_P3_U3120 = ~new_P3_LT_563_U6 | ~new_P3_U4313 | ~new_P3_U3262 | ~new_P3_U7949 | ~new_P3_U7948;
  assign new_P3_U3121 = ~P3_STATE2_REG_0_;
  assign new_P3_U3122 = ~P3_STATE2_REG_0_ | ~new_P3_U4629;
  assign new_P3_U3123 = P3_STATE2_REG_3_ | P3_STATE2_REG_1_;
  assign new_P3_U3124 = ~P3_STATE2_REG_2_ | ~new_P3_U3089;
  assign new_P3_U3125 = P3_STATE2_REG_2_ | P3_STATE2_REG_1_;
  assign new_P3_U3126 = ~new_P3_LTE_597_U6 | ~P3_STATE2_REG_3_;
  assign new_P3_U3127 = ~new_P3_U4666 | ~new_P3_U3121;
  assign new_P3_U3128 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_U3129 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_U3130 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_U3131 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_U3132 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_U4648;
  assign new_P3_U3133 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_U3134 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_U4649;
  assign new_P3_U3135 = P3_STATE2_REG_3_ | P3_STATE2_REG_2_;
  assign new_P3_U3136 = ~new_P3_U4295 | ~P3_STATEBS16_REG;
  assign new_P3_U3137 = ~new_P3_U3153 | ~new_P3_U4641;
  assign new_P3_U3138 = ~new_P3_U3137 | ~new_P3_U3128;
  assign new_P3_U3139 = ~new_P3_U3180 | ~new_P3_U4651;
  assign new_P3_U3140 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_U3141;
  assign new_P3_U3141 = ~new_P3_U3150 | ~new_P3_U3158;
  assign new_P3_U3142 = ~new_P3_U4331 | ~new_P3_U4655;
  assign new_P3_U3143 = ~new_P3_U3156 | ~new_P3_U3128;
  assign new_P3_U3144 = ~new_P3_U4647 | ~new_P3_U2486;
  assign new_P3_U3145 = ~new_P3_U3144 | ~new_P3_U4667;
  assign new_P3_U3146 = ~new_P3_U3134 | ~new_P3_U4663;
  assign new_P3_U3147 = ~new_P3_U3386 | ~new_P3_U2492;
  assign new_P3_U3148 = ~new_P3_U3141 | ~new_P3_U3128;
  assign new_P3_U3149 = ~new_P3_U2490 | ~new_P3_U2486;
  assign new_P3_U3150 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_U3137;
  assign new_P3_U3151 = ~new_P3_U3149 | ~new_P3_U4719;
  assign new_P3_U3152 = ~new_P3_U3147 | ~new_P3_U4717;
  assign new_P3_U3153 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_U3129;
  assign new_P3_U3154 = ~new_P3_U3404 | ~new_P3_U4640;
  assign new_P3_U3155 = ~new_P3_U4643 | ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_U3156 = ~new_P3_U3148 | ~new_P3_U3155;
  assign new_P3_U3157 = ~new_P3_U2493 | ~new_P3_U2486;
  assign new_P3_U3158 = ~new_P3_U4642 | ~new_P3_U3128;
  assign new_P3_U3159 = ~new_P3_U3157 | ~new_P3_U4771;
  assign new_P3_U3160 = ~new_P3_U3154 | ~new_P3_U4769;
  assign new_P3_U3161 = ~new_P3_U3422 | ~new_P3_U2492;
  assign new_P3_U3162 = ~new_P3_U2495 | ~new_P3_U2486;
  assign new_P3_U3163 = ~new_P3_U3162 | ~new_P3_U4822;
  assign new_P3_U3164 = ~new_P3_U4648 | ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_U3131;
  assign new_P3_U3165 = ~new_P3_U7965 | ~new_P3_U3142;
  assign new_P3_U3166 = ~new_P3_U2498 | ~new_P3_U4647;
  assign new_P3_U3167 = ~new_P3_U3166 | ~new_P3_U4874;
  assign new_P3_U3168 = ~new_P3_U3164 | ~new_P3_U4872;
  assign new_P3_U3169 = ~new_P3_U3457 | ~new_P3_U2501;
  assign new_P3_U3170 = ~new_P3_U2498 | ~new_P3_U2490;
  assign new_P3_U3171 = ~new_P3_U3170 | ~new_P3_U4926;
  assign new_P3_U3172 = ~new_P3_U3169 | ~new_P3_U4924;
  assign new_P3_U3173 = ~new_P3_U3475 | ~new_P3_U4640;
  assign new_P3_U3174 = ~new_P3_U2498 | ~new_P3_U2493;
  assign new_P3_U3175 = ~new_P3_U3174 | ~new_P3_U4978;
  assign new_P3_U3176 = ~new_P3_U3173 | ~new_P3_U4976;
  assign new_P3_U3177 = ~new_P3_U2501 | ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_U3129;
  assign new_P3_U3178 = ~new_P3_U2498 | ~new_P3_U2495;
  assign new_P3_U3179 = ~new_P3_U3178 | ~new_P3_U5029;
  assign new_P3_U3180 = ~new_P3_U4649 | ~new_P3_U3133;
  assign new_P3_U3181 = ~new_P3_U2485 | ~new_P3_U4657;
  assign new_P3_U3182 = ~new_P3_U3368 | ~new_P3_U3181;
  assign new_P3_U3183 = ~new_P3_U2504 | ~new_P3_U4647;
  assign new_P3_U3184 = ~new_P3_U3183 | ~new_P3_U3181;
  assign new_P3_U3185 = ~new_P3_U3180 | ~new_P3_U4331;
  assign new_P3_U3186 = ~new_P3_U3527 | ~new_P3_U2492;
  assign new_P3_U3187 = ~new_P3_U2504 | ~new_P3_U2490;
  assign new_P3_U3188 = ~new_P3_U3187 | ~new_P3_U5130;
  assign new_P3_U3189 = ~new_P3_U3186 | ~new_P3_U5128;
  assign new_P3_U3190 = ~new_P3_U3545 | ~new_P3_U4640;
  assign new_P3_U3191 = ~new_P3_U2504 | ~new_P3_U2493;
  assign new_P3_U3192 = ~new_P3_U3191 | ~new_P3_U5182;
  assign new_P3_U3193 = ~new_P3_U3190 | ~new_P3_U5180;
  assign new_P3_U3194 = ~new_P3_U3563 | ~new_P3_U2492;
  assign new_P3_U3195 = ~new_P3_U2504 | ~new_P3_U2495;
  assign new_P3_U3196 = ~new_P3_U3581 | ~new_P3_U4648;
  assign new_P3_U3197 = ~new_P3_U2508 | ~new_P3_U4647;
  assign new_P3_U3198 = ~new_P3_U3196 | ~new_P3_U5282;
  assign new_P3_U3199 = ~new_P3_U2501 | ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_U3133;
  assign new_P3_U3200 = ~new_P3_U2508 | ~new_P3_U2490;
  assign new_P3_U3201 = ~new_P3_U3199 | ~new_P3_U5333;
  assign new_P3_U3202 = ~new_P3_U3616 | ~new_P3_U4640;
  assign new_P3_U3203 = ~new_P3_U2508 | ~new_P3_U2493;
  assign new_P3_U3204 = ~new_P3_U3202 | ~new_P3_U5384;
  assign new_P3_U3205 = ~new_P3_U3634 | ~new_P3_U2501;
  assign new_P3_U3206 = ~new_P3_U2508 | ~new_P3_U2495;
  assign new_P3_U3207 = ~P3_FLUSH_REG;
  assign new_P3_U3208 = ~new_P3_U4539 | ~new_P3_U3102;
  assign new_P3_U3209 = ~new_P3_U2514 | ~new_P3_U3113;
  assign new_P3_U3210 = ~new_P3_GTE_412_U6;
  assign new_P3_U3211 = ~new_P3_GTE_485_U6;
  assign new_P3_U3212 = ~new_P3_GTE_390_U6;
  assign new_P3_U3213 = ~new_P3_GTE_450_U6;
  assign new_P3_U3214 = ~new_P3_GTE_504_U6;
  assign new_P3_U3215 = ~new_P3_GTE_401_U6;
  assign new_P3_U3216 = ~new_P3_U4590 | ~new_P3_U3074;
  assign new_P3_U3217 = ~new_P3_U2450 | ~new_P3_U4323;
  assign new_P3_U3218 = ~new_P3_U3333 | ~new_P3_U3334 | ~new_P3_U3337 | ~new_P3_U3336 | ~new_P3_U3335;
  assign new_P3_U3219 = ~new_P3_U3662 | ~new_P3_U2461;
  assign new_P3_U3220 = ~new_P3_U3667 | ~new_P3_U7976 | ~new_P3_U7975;
  assign new_P3_U3221 = ~new_P3_U5524 | ~new_P3_U3222 | ~new_P3_U3119;
  assign new_P3_U3222 = ~new_P3_U4314 | ~new_P3_U3218;
  assign new_P3_U3223 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_U5503;
  assign new_P3_U3224 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_U5505;
  assign new_P3_U3225 = ~new_P3_U3096 | ~new_P3_U3227;
  assign new_P3_U3226 = ~new_P3_U3674 | ~new_P3_U2517;
  assign new_P3_U3227 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U3095;
  assign new_P3_U3228 = ~new_P3_U3091 | ~new_P3_U3095;
  assign new_P3_U3229 = ~new_P3_U4350 | ~new_P3_U4323 | ~new_P3_U3218;
  assign new_P3_U3230 = ~new_P3_U2518 | ~new_P3_U3243;
  assign new_P3_U3231 = ~new_P3_U3115 | ~new_P3_U5559;
  assign new_P3_U3232 = ~new_P3_LT_589_U6;
  assign new_P3_U3233 = ~new_P3_U5578 | ~new_P3_U4330 | ~new_P3_U3127;
  assign new_P3_U3234 = ~new_P3_U3135 | ~new_P3_U3123;
  assign new_P3_U3235 = ~new_P3_U4294 | ~new_P3_U3101 | ~new_P3_U3104;
  assign new_P3_U3236 = ~new_P3_U4505 | ~new_P3_U3101 | ~new_P3_U2630;
  assign new_P3_U3237 = ~new_P3_GTE_370_U6;
  assign new_P3_U3238 = ~new_P3_GTE_355_U6;
  assign new_P3_U3239 = ~new_P3_U4295 | ~new_P3_U3089;
  assign new_P3_U3240 = ~P3_REIP_REG_0_;
  assign new_P3_U3241 = ~new_P3_U2628;
  assign new_P3_U3242 = ~new_P3_U3661 | ~new_P3_U2450;
  assign new_P3_U3243 = ~new_P3_U2461 | ~new_P3_U4314;
  assign new_P3_U3244 = ~new_P3_U4352 | ~new_P3_U4522;
  assign new_P3_U3245 = ~new_P3_U4352 | ~new_P3_U3102;
  assign new_P3_U3246 = ~new_P3_U3664 | ~new_P3_U3663 | ~new_P3_U2449;
  assign new_P3_U3247 = ~P3_STATE2_REG_2_ | ~new_P3_U3248;
  assign new_P3_U3248 = ~new_P3_U4336 | ~new_P3_U5630;
  assign new_P3_U3249 = ~new_P3_U6403 | ~new_P3_U6402;
  assign new_P3_U3250 = ~new_P3_U2390 | ~new_P3_U6663;
  assign new_P3_U3251 = ~new_P3_U6758 | ~new_P3_U6757;
  assign new_P3_U3252 = ~new_P3_U2390 | ~new_P3_U6853;
  assign new_P3_U3253 = ~new_P3_U2390 | ~new_P3_U6997;
  assign new_P3_U3254 = ~new_P3_U5490 | ~new_P3_U5489;
  assign new_P3_U3255 = ~new_P3_U5487 | ~new_P3_U5486;
  assign new_P3_U3256 = ~P3_EBX_REG_31_;
  assign new_P3_U3257 = P3_STATEBS16_REG | new_U209;
  assign new_P3_U3258 = ~new_P3_ADD_318_U69;
  assign new_P3_U3259 = ~new_P3_ADD_318_U69 | ~new_P3_U2385;
  assign new_P3_U3260 = ~new_P3_U4030 | ~new_P3_U4334;
  assign new_P3_U3261 = ~new_P3_U4138 | ~new_P3_U4141 | ~new_P3_U4148 | ~new_P3_U4144;
  assign new_P3_U3262 = ~new_P3_U4282 | ~new_P3_U2462 | ~new_P3_U3108;
  assign new_P3_U3263 = ~P3_CODEFETCH_REG;
  assign new_P3_U3264 = ~P3_READREQUEST_REG;
  assign new_P3_U3265 = ~new_P3_U3099 | ~new_P3_U3224;
  assign new_P3_U3266 = ~new_P3_U3223 | ~new_P3_U7515;
  assign new_P3_U3267 = ~new_P3_U4289 | ~new_P3_U3092;
  assign new_P3_U3268 = ~new_P3_U3098 | ~new_P3_U7774;
  assign new_P3_U3269 = ~new_P3_U7961 | ~new_P3_U7960;
  assign new_P3_U3270 = ~new_P3_U7964 | ~new_P3_U7963;
  assign new_P3_U3271 = ~new_P3_U7967 | ~new_P3_U7966;
  assign new_P3_U3272 = ~new_P3_U8033 | ~new_P3_U8032;
  assign new_P3_U3273 = ~new_P3_U8036 | ~new_P3_U8035;
  assign n620 = ~new_P3_U7921 | ~new_P3_U7920;
  assign n625 = ~new_P3_U7923 | ~new_P3_U7922;
  assign n630 = ~new_P3_U7925 | ~new_P3_U7924;
  assign n635 = ~new_P3_U7927 | ~new_P3_U7926;
  assign new_P3_U3278 = ~new_P3_U7936 | ~new_P3_U7935;
  assign new_P3_U3279 = new_P3_U3083 & new_P3_U4286;
  assign n805 = ~new_P3_U7939 | ~new_P3_U7938;
  assign n810 = ~new_P3_U7941 | ~new_P3_U7940;
  assign n965 = ~new_P3_U7955 | ~new_P3_U7954;
  assign new_P3_U3283 = new_P3_U3652 & new_P3_U2356;
  assign n1625 = ~new_P3_U7972 | ~new_P3_U7971;
  assign n1630 = ~new_P3_U7980 | ~new_P3_U7979;
  assign new_P3_U3286 = ~new_P3_U7987 | ~new_P3_U7986;
  assign new_P3_U3287 = ~new_P3_U7984 | ~new_P3_U7983;
  assign n1635 = ~new_P3_U7990 | ~new_P3_U7989;
  assign n1640 = ~new_P3_U7992 | ~new_P3_U7991;
  assign n1645 = ~new_P3_U7996 | ~new_P3_U7995;
  assign new_P3_U3291 = ~P3_DATAWIDTH_REG_1_ & ~P3_REIP_REG_1_;
  assign n2763 = ~new_P3_U8011 | ~new_P3_U8010;
  assign n2773 = ~new_P3_U8015 | ~new_P3_U8014;
  assign n2778 = ~new_P3_U8017 | ~new_P3_U8016;
  assign n2787 = ~new_P3_U8019 | ~new_P3_U8018;
  assign n2797 = ~new_P3_U8023 | ~new_P3_U8022;
  assign n2806 = ~new_P3_U8027 | ~new_P3_U8026;
  assign n2819 = ~new_P3_U8029 | ~new_P3_U8028;
  assign n2824 = ~new_P3_U8031 | ~new_P3_U8030;
  assign new_P3_U3300 = ~new_P3_U8039 | ~new_P3_U8038;
  assign new_P3_U3301 = ~new_P3_U8041 | ~new_P3_U8040;
  assign new_P3_U3302 = ~new_P3_U8043 | ~new_P3_U8042;
  assign new_P3_U3303 = new_P3_ADD_495_U8 & new_P3_U2356;
  assign new_P3_U3304 = ~new_P3_U8045 | ~new_P3_U8044;
  assign new_P3_U3305 = ~new_P3_U8047 | ~new_P3_U8046;
  assign new_P3_U3306 = ~new_P3_U8049 | ~new_P3_U8048;
  assign new_P3_U3307 = ~new_P3_U8051 | ~new_P3_U8050;
  assign new_P3_U3308 = ~new_P3_U8053 | ~new_P3_U8052;
  assign new_P3_U3309 = P3_STATE_REG_0_ & new_P3_U4447;
  assign new_P3_U3310 = new_P3_U4456 & new_P3_U3080;
  assign new_P3_U3311 = new_P3_U4458 & new_P3_U3078;
  assign new_P3_U3312 = P3_REQUESTPENDING_REG & P3_STATE_REG_0_;
  assign new_P3_U3313 = new_P3_U4472 & new_P3_U4473 & new_P3_U4475 & new_P3_U4474;
  assign new_P3_U3314 = new_P3_U4476 & new_P3_U4477 & new_P3_U4479 & new_P3_U4478;
  assign new_P3_U3315 = new_P3_U4481 & new_P3_U4480;
  assign new_P3_U3316 = new_P3_U4483 & new_P3_U4482;
  assign new_P3_U3317 = new_P3_U4484 & new_P3_U4485 & new_P3_U4487 & new_P3_U4486;
  assign new_P3_U3318 = new_P3_U4489 & new_P3_U4490 & new_P3_U4492 & new_P3_U4491;
  assign new_P3_U3319 = new_P3_U4493 & new_P3_U4494 & new_P3_U4496 & new_P3_U4495;
  assign new_P3_U3320 = new_P3_U4498 & new_P3_U4497;
  assign new_P3_U3321 = new_P3_U4500 & new_P3_U4499;
  assign new_P3_U3322 = new_P3_U4501 & new_P3_U4502 & new_P3_U4504 & new_P3_U4503;
  assign new_P3_U3323 = new_P3_U4506 & new_P3_U4507 & new_P3_U4509 & new_P3_U4508;
  assign new_P3_U3324 = new_P3_U4510 & new_P3_U4511 & new_P3_U4513 & new_P3_U4512;
  assign new_P3_U3325 = new_P3_U4515 & new_P3_U4514;
  assign new_P3_U3326 = new_P3_U4517 & new_P3_U4516;
  assign new_P3_U3327 = new_P3_U4518 & new_P3_U4519 & new_P3_U4521 & new_P3_U4520;
  assign new_P3_U3328 = new_P3_U4540 & new_P3_U4541 & new_P3_U4543 & new_P3_U4542;
  assign new_P3_U3329 = new_P3_U4544 & new_P3_U4545 & new_P3_U4547 & new_P3_U4546;
  assign new_P3_U3330 = new_P3_U4549 & new_P3_U4548;
  assign new_P3_U3331 = new_P3_U4551 & new_P3_U4550;
  assign new_P3_U3332 = new_P3_U4552 & new_P3_U4553 & new_P3_U4555 & new_P3_U4554;
  assign new_P3_U3333 = new_P3_U4557 & new_P3_U4558 & new_P3_U4560 & new_P3_U4559;
  assign new_P3_U3334 = new_P3_U4561 & new_P3_U4562 & new_P3_U4564 & new_P3_U4563;
  assign new_P3_U3335 = new_P3_U4566 & new_P3_U4565;
  assign new_P3_U3336 = new_P3_U4568 & new_P3_U4567;
  assign new_P3_U3337 = new_P3_U4569 & new_P3_U4570 & new_P3_U4572 & new_P3_U4571;
  assign new_P3_U3338 = new_P3_U4523 & new_P3_U4524 & new_P3_U4526 & new_P3_U4525;
  assign new_P3_U3339 = new_P3_U4527 & new_P3_U4528 & new_P3_U4530 & new_P3_U4529;
  assign new_P3_U3340 = new_P3_U4532 & new_P3_U4531;
  assign new_P3_U3341 = new_P3_U4534 & new_P3_U4533;
  assign new_P3_U3342 = new_P3_U4535 & new_P3_U4536 & new_P3_U4538 & new_P3_U4537;
  assign new_P3_U3343 = new_P3_U4591 & new_P3_U4592 & new_P3_U4594 & new_P3_U4593;
  assign new_P3_U3344 = new_P3_U4595 & new_P3_U4596 & new_P3_U4598 & new_P3_U4597;
  assign new_P3_U3345 = new_P3_U4600 & new_P3_U4599;
  assign new_P3_U3346 = new_P3_U4602 & new_P3_U4601;
  assign new_P3_U3347 = new_P3_U4603 & new_P3_U4604 & new_P3_U4606 & new_P3_U4605;
  assign new_P3_U3348 = new_P3_U4574 & new_P3_U4575 & new_P3_U4577 & new_P3_U4576;
  assign new_P3_U3349 = new_P3_U4578 & new_P3_U4579 & new_P3_U4581 & new_P3_U4580;
  assign new_P3_U3350 = new_P3_U4583 & new_P3_U4582;
  assign new_P3_U3351 = new_P3_U4585 & new_P3_U4584;
  assign new_P3_U3352 = new_P3_U4586 & new_P3_U4587 & new_P3_U4589 & new_P3_U4588;
  assign new_P3_U3353 = new_P3_U2352 & new_P3_U4293;
  assign new_P3_U3354 = new_P3_U4556 & new_P3_U3218;
  assign new_P3_U3355 = new_P3_U4323 & new_P3_U3101;
  assign new_P3_U3356 = new_P3_U4324 & new_P3_U3101;
  assign new_P3_U3357 = new_P3_U4609 & new_P3_U4610 & new_P3_U4612 & new_P3_U4611;
  assign new_P3_U3358 = new_P3_U4613 & new_P3_U4614 & new_P3_U4616 & new_P3_U4615;
  assign new_P3_U3359 = new_P3_U4539 & new_P3_U2630;
  assign new_P3_U3360 = new_P3_U3218 & new_P3_U3107 & new_P3_U3108;
  assign new_P3_U3361 = new_P3_U4621 & new_P3_U3235 & new_P3_U3236;
  assign new_P3_U3362 = new_P3_U4626 & new_P3_U3089;
  assign new_P3_U3363 = new_P3_U4631 & new_P3_U3124;
  assign new_P3_U3364 = new_P3_U4340 & new_P3_U2630;
  assign new_P3_U3365 = P3_STATE2_REG_3_ & P3_STATE2_REG_0_;
  assign new_P3_U3366 = new_P3_U4338 & new_P3_U4328;
  assign new_P3_U3367 = new_P3_U3366 & new_P3_U4639;
  assign new_P3_U3368 = new_P3_U3165 & new_P3_U4659;
  assign new_P3_U3369 = new_P3_U4671 & new_P3_U4312;
  assign new_P3_U3370 = new_P3_U4676 & new_P3_U4675;
  assign new_P3_U3371 = new_P3_U3370 & new_P3_U4677;
  assign new_P3_U3372 = new_P3_U4681 & new_P3_U4680;
  assign new_P3_U3373 = new_P3_U3372 & new_P3_U4682;
  assign new_P3_U3374 = new_P3_U4686 & new_P3_U4685;
  assign new_P3_U3375 = new_P3_U3374 & new_P3_U4687;
  assign new_P3_U3376 = new_P3_U4691 & new_P3_U4690;
  assign new_P3_U3377 = new_P3_U3376 & new_P3_U4692;
  assign new_P3_U3378 = new_P3_U4696 & new_P3_U4695;
  assign new_P3_U3379 = new_P3_U3378 & new_P3_U4697;
  assign new_P3_U3380 = new_P3_U4701 & new_P3_U4700;
  assign new_P3_U3381 = new_P3_U3380 & new_P3_U4702;
  assign new_P3_U3382 = new_P3_U4706 & new_P3_U4705;
  assign new_P3_U3383 = new_P3_U3382 & new_P3_U4707;
  assign new_P3_U3384 = new_P3_U4711 & new_P3_U4710;
  assign new_P3_U3385 = new_P3_U3384 & new_P3_U4712;
  assign new_P3_U3386 = P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_U3387 = new_P3_U4723 & new_P3_U4312;
  assign new_P3_U3388 = new_P3_U4728 & new_P3_U4727;
  assign new_P3_U3389 = new_P3_U3388 & new_P3_U4729;
  assign new_P3_U3390 = new_P3_U4733 & new_P3_U4732;
  assign new_P3_U3391 = new_P3_U3390 & new_P3_U4734;
  assign new_P3_U3392 = new_P3_U4738 & new_P3_U4737;
  assign new_P3_U3393 = new_P3_U3392 & new_P3_U4739;
  assign new_P3_U3394 = new_P3_U4743 & new_P3_U4742;
  assign new_P3_U3395 = new_P3_U3394 & new_P3_U4744;
  assign new_P3_U3396 = new_P3_U4748 & new_P3_U4747;
  assign new_P3_U3397 = new_P3_U3396 & new_P3_U4749;
  assign new_P3_U3398 = new_P3_U4753 & new_P3_U4752;
  assign new_P3_U3399 = new_P3_U3398 & new_P3_U4754;
  assign new_P3_U3400 = new_P3_U4758 & new_P3_U4757;
  assign new_P3_U3401 = new_P3_U3400 & new_P3_U4759;
  assign new_P3_U3402 = new_P3_U4763 & new_P3_U4762;
  assign new_P3_U3403 = new_P3_U3402 & new_P3_U4764;
  assign new_P3_U3404 = P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_U3405 = new_P3_U4775 & new_P3_U4312;
  assign new_P3_U3406 = new_P3_U4780 & new_P3_U4779;
  assign new_P3_U3407 = new_P3_U3406 & new_P3_U4781;
  assign new_P3_U3408 = new_P3_U4785 & new_P3_U4784;
  assign new_P3_U3409 = new_P3_U3408 & new_P3_U4786;
  assign new_P3_U3410 = new_P3_U4790 & new_P3_U4789;
  assign new_P3_U3411 = new_P3_U3410 & new_P3_U4791;
  assign new_P3_U3412 = new_P3_U4795 & new_P3_U4794;
  assign new_P3_U3413 = new_P3_U3412 & new_P3_U4796;
  assign new_P3_U3414 = new_P3_U4800 & new_P3_U4799;
  assign new_P3_U3415 = new_P3_U3414 & new_P3_U4801;
  assign new_P3_U3416 = new_P3_U4805 & new_P3_U4804;
  assign new_P3_U3417 = new_P3_U3416 & new_P3_U4806;
  assign new_P3_U3418 = new_P3_U4810 & new_P3_U4809;
  assign new_P3_U3419 = new_P3_U3418 & new_P3_U4811;
  assign new_P3_U3420 = new_P3_U4815 & new_P3_U4814;
  assign new_P3_U3421 = new_P3_U3420 & new_P3_U4816;
  assign new_P3_U3422 = P3_INSTQUEUEWR_ADDR_REG_3_ & new_P3_U3129;
  assign new_P3_U3423 = new_P3_U4826 & new_P3_U4312;
  assign new_P3_U3424 = new_P3_U4831 & new_P3_U4830;
  assign new_P3_U3425 = new_P3_U3424 & new_P3_U4832;
  assign new_P3_U3426 = new_P3_U4836 & new_P3_U4835;
  assign new_P3_U3427 = new_P3_U3426 & new_P3_U4837;
  assign new_P3_U3428 = new_P3_U4841 & new_P3_U4840;
  assign new_P3_U3429 = new_P3_U3428 & new_P3_U4842;
  assign new_P3_U3430 = new_P3_U4846 & new_P3_U4845;
  assign new_P3_U3431 = new_P3_U3430 & new_P3_U4847;
  assign new_P3_U3432 = new_P3_U4851 & new_P3_U4850;
  assign new_P3_U3433 = new_P3_U3432 & new_P3_U4852;
  assign new_P3_U3434 = new_P3_U4856 & new_P3_U4855;
  assign new_P3_U3435 = new_P3_U3434 & new_P3_U4857;
  assign new_P3_U3436 = new_P3_U4861 & new_P3_U4860;
  assign new_P3_U3437 = new_P3_U3436 & new_P3_U4862;
  assign new_P3_U3438 = new_P3_U4866 & new_P3_U4865;
  assign new_P3_U3439 = new_P3_U3438 & new_P3_U4867;
  assign new_P3_U3440 = new_P3_U4878 & new_P3_U4312;
  assign new_P3_U3441 = new_P3_U4883 & new_P3_U4882;
  assign new_P3_U3442 = new_P3_U3441 & new_P3_U4884;
  assign new_P3_U3443 = new_P3_U4888 & new_P3_U4887;
  assign new_P3_U3444 = new_P3_U3443 & new_P3_U4889;
  assign new_P3_U3445 = new_P3_U4893 & new_P3_U4892;
  assign new_P3_U3446 = new_P3_U3445 & new_P3_U4894;
  assign new_P3_U3447 = new_P3_U4898 & new_P3_U4897;
  assign new_P3_U3448 = new_P3_U3447 & new_P3_U4899;
  assign new_P3_U3449 = new_P3_U4903 & new_P3_U4902;
  assign new_P3_U3450 = new_P3_U3449 & new_P3_U4904;
  assign new_P3_U3451 = new_P3_U4908 & new_P3_U4907;
  assign new_P3_U3452 = new_P3_U3451 & new_P3_U4909;
  assign new_P3_U3453 = new_P3_U4913 & new_P3_U4912;
  assign new_P3_U3454 = new_P3_U3453 & new_P3_U4914;
  assign new_P3_U3455 = new_P3_U4918 & new_P3_U4917;
  assign new_P3_U3456 = new_P3_U3455 & new_P3_U4919;
  assign new_P3_U3457 = P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_U3458 = new_P3_U4930 & new_P3_U4312;
  assign new_P3_U3459 = new_P3_U4935 & new_P3_U4934;
  assign new_P3_U3460 = new_P3_U3459 & new_P3_U4936;
  assign new_P3_U3461 = new_P3_U4940 & new_P3_U4939;
  assign new_P3_U3462 = new_P3_U3461 & new_P3_U4941;
  assign new_P3_U3463 = new_P3_U4945 & new_P3_U4944;
  assign new_P3_U3464 = new_P3_U3463 & new_P3_U4946;
  assign new_P3_U3465 = new_P3_U4950 & new_P3_U4949;
  assign new_P3_U3466 = new_P3_U3465 & new_P3_U4951;
  assign new_P3_U3467 = new_P3_U4955 & new_P3_U4954;
  assign new_P3_U3468 = new_P3_U3467 & new_P3_U4956;
  assign new_P3_U3469 = new_P3_U4960 & new_P3_U4959;
  assign new_P3_U3470 = new_P3_U3469 & new_P3_U4961;
  assign new_P3_U3471 = new_P3_U4965 & new_P3_U4964;
  assign new_P3_U3472 = new_P3_U3471 & new_P3_U4966;
  assign new_P3_U3473 = new_P3_U4970 & new_P3_U4969;
  assign new_P3_U3474 = new_P3_U3473 & new_P3_U4971;
  assign new_P3_U3475 = P3_INSTQUEUEWR_ADDR_REG_3_ & new_P3_U3131;
  assign new_P3_U3476 = new_P3_U4982 & new_P3_U4312;
  assign new_P3_U3477 = new_P3_U4987 & new_P3_U4986;
  assign new_P3_U3478 = new_P3_U3477 & new_P3_U4988;
  assign new_P3_U3479 = new_P3_U4992 & new_P3_U4991;
  assign new_P3_U3480 = new_P3_U3479 & new_P3_U4993;
  assign new_P3_U3481 = new_P3_U4997 & new_P3_U4996;
  assign new_P3_U3482 = new_P3_U3481 & new_P3_U4998;
  assign new_P3_U3483 = new_P3_U5002 & new_P3_U5001;
  assign new_P3_U3484 = new_P3_U3483 & new_P3_U5003;
  assign new_P3_U3485 = new_P3_U5007 & new_P3_U5006;
  assign new_P3_U3486 = new_P3_U3485 & new_P3_U5008;
  assign new_P3_U3487 = new_P3_U5012 & new_P3_U5011;
  assign new_P3_U3488 = new_P3_U3487 & new_P3_U5013;
  assign new_P3_U3489 = new_P3_U5017 & new_P3_U5016;
  assign new_P3_U3490 = new_P3_U3489 & new_P3_U5018;
  assign new_P3_U3491 = new_P3_U5022 & new_P3_U5021;
  assign new_P3_U3492 = new_P3_U3491 & new_P3_U5023;
  assign new_P3_U3493 = new_P3_U5033 & new_P3_U4312;
  assign new_P3_U3494 = new_P3_U5038 & new_P3_U5037;
  assign new_P3_U3495 = new_P3_U3494 & new_P3_U5039;
  assign new_P3_U3496 = new_P3_U5043 & new_P3_U5042;
  assign new_P3_U3497 = new_P3_U3496 & new_P3_U5044;
  assign new_P3_U3498 = new_P3_U5048 & new_P3_U5047;
  assign new_P3_U3499 = new_P3_U3498 & new_P3_U5049;
  assign new_P3_U3500 = new_P3_U5053 & new_P3_U5052;
  assign new_P3_U3501 = new_P3_U3500 & new_P3_U5054;
  assign new_P3_U3502 = new_P3_U5058 & new_P3_U5057;
  assign new_P3_U3503 = new_P3_U3502 & new_P3_U5059;
  assign new_P3_U3504 = new_P3_U5063 & new_P3_U5062;
  assign new_P3_U3505 = new_P3_U3504 & new_P3_U5064;
  assign new_P3_U3506 = new_P3_U5068 & new_P3_U5067;
  assign new_P3_U3507 = new_P3_U3506 & new_P3_U5069;
  assign new_P3_U3508 = new_P3_U5073 & new_P3_U5072;
  assign new_P3_U3509 = new_P3_U3508 & new_P3_U5074;
  assign new_P3_U3510 = new_P3_U5082 & new_P3_U4312;
  assign new_P3_U3511 = new_P3_U5087 & new_P3_U5086;
  assign new_P3_U3512 = new_P3_U3511 & new_P3_U5088;
  assign new_P3_U3513 = new_P3_U5092 & new_P3_U5091;
  assign new_P3_U3514 = new_P3_U3513 & new_P3_U5093;
  assign new_P3_U3515 = new_P3_U5097 & new_P3_U5096;
  assign new_P3_U3516 = new_P3_U3515 & new_P3_U5098;
  assign new_P3_U3517 = new_P3_U5102 & new_P3_U5101;
  assign new_P3_U3518 = new_P3_U3517 & new_P3_U5103;
  assign new_P3_U3519 = new_P3_U5107 & new_P3_U5106;
  assign new_P3_U3520 = new_P3_U3519 & new_P3_U5108;
  assign new_P3_U3521 = new_P3_U5112 & new_P3_U5111;
  assign new_P3_U3522 = new_P3_U3521 & new_P3_U5113;
  assign new_P3_U3523 = new_P3_U5117 & new_P3_U5116;
  assign new_P3_U3524 = new_P3_U3523 & new_P3_U5118;
  assign new_P3_U3525 = new_P3_U5122 & new_P3_U5121;
  assign new_P3_U3526 = new_P3_U3525 & new_P3_U5123;
  assign new_P3_U3527 = P3_INSTQUEUEWR_ADDR_REG_1_ & new_P3_U3133;
  assign new_P3_U3528 = new_P3_U5134 & new_P3_U4312;
  assign new_P3_U3529 = new_P3_U5139 & new_P3_U5138;
  assign new_P3_U3530 = new_P3_U3529 & new_P3_U5140;
  assign new_P3_U3531 = new_P3_U5144 & new_P3_U5143;
  assign new_P3_U3532 = new_P3_U3531 & new_P3_U5145;
  assign new_P3_U3533 = new_P3_U5149 & new_P3_U5148;
  assign new_P3_U3534 = new_P3_U3533 & new_P3_U5150;
  assign new_P3_U3535 = new_P3_U5154 & new_P3_U5153;
  assign new_P3_U3536 = new_P3_U3535 & new_P3_U5155;
  assign new_P3_U3537 = new_P3_U5159 & new_P3_U5158;
  assign new_P3_U3538 = new_P3_U3537 & new_P3_U5160;
  assign new_P3_U3539 = new_P3_U5164 & new_P3_U5163;
  assign new_P3_U3540 = new_P3_U3539 & new_P3_U5165;
  assign new_P3_U3541 = new_P3_U5169 & new_P3_U5168;
  assign new_P3_U3542 = new_P3_U3541 & new_P3_U5170;
  assign new_P3_U3543 = new_P3_U5174 & new_P3_U5173;
  assign new_P3_U3544 = new_P3_U3543 & new_P3_U5175;
  assign new_P3_U3545 = P3_INSTQUEUEWR_ADDR_REG_2_ & new_P3_U3133;
  assign new_P3_U3546 = new_P3_U5186 & new_P3_U4312;
  assign new_P3_U3547 = new_P3_U5191 & new_P3_U5190;
  assign new_P3_U3548 = new_P3_U3547 & new_P3_U5192;
  assign new_P3_U3549 = new_P3_U5196 & new_P3_U5195;
  assign new_P3_U3550 = new_P3_U3549 & new_P3_U5197;
  assign new_P3_U3551 = new_P3_U5201 & new_P3_U5200;
  assign new_P3_U3552 = new_P3_U3551 & new_P3_U5202;
  assign new_P3_U3553 = new_P3_U5206 & new_P3_U5205;
  assign new_P3_U3554 = new_P3_U3553 & new_P3_U5207;
  assign new_P3_U3555 = new_P3_U5211 & new_P3_U5210;
  assign new_P3_U3556 = new_P3_U3555 & new_P3_U5212;
  assign new_P3_U3557 = new_P3_U5216 & new_P3_U5215;
  assign new_P3_U3558 = new_P3_U3557 & new_P3_U5217;
  assign new_P3_U3559 = new_P3_U5221 & new_P3_U5220;
  assign new_P3_U3560 = new_P3_U3559 & new_P3_U5222;
  assign new_P3_U3561 = new_P3_U5226 & new_P3_U5225;
  assign new_P3_U3562 = new_P3_U3561 & new_P3_U5227;
  assign new_P3_U3563 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_U3564 = new_P3_U5237 & new_P3_U4312;
  assign new_P3_U3565 = new_P3_U5243 & new_P3_U5241 & new_P3_U5240;
  assign new_P3_U3566 = new_P3_U3565 & new_P3_U5242;
  assign new_P3_U3567 = new_P3_U5248 & new_P3_U5246 & new_P3_U5245;
  assign new_P3_U3568 = new_P3_U3567 & new_P3_U5247;
  assign new_P3_U3569 = new_P3_U5253 & new_P3_U5251 & new_P3_U5250;
  assign new_P3_U3570 = new_P3_U3569 & new_P3_U5252;
  assign new_P3_U3571 = new_P3_U5258 & new_P3_U5256 & new_P3_U5255;
  assign new_P3_U3572 = new_P3_U3571 & new_P3_U5257;
  assign new_P3_U3573 = new_P3_U5263 & new_P3_U5261 & new_P3_U5260;
  assign new_P3_U3574 = new_P3_U3573 & new_P3_U5262;
  assign new_P3_U3575 = new_P3_U5268 & new_P3_U5266 & new_P3_U5265;
  assign new_P3_U3576 = new_P3_U3575 & new_P3_U5267;
  assign new_P3_U3577 = new_P3_U5273 & new_P3_U5271 & new_P3_U5270;
  assign new_P3_U3578 = new_P3_U3577 & new_P3_U5272;
  assign new_P3_U3579 = new_P3_U5278 & new_P3_U5276 & new_P3_U5275;
  assign new_P3_U3580 = new_P3_U3579 & new_P3_U5277;
  assign new_P3_U3581 = ~P3_INSTQUEUEWR_ADDR_REG_2_ & ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_U3582 = new_P3_U5288 & new_P3_U4312;
  assign new_P3_U3583 = new_P3_U5294 & new_P3_U5292 & new_P3_U5291;
  assign new_P3_U3584 = new_P3_U3583 & new_P3_U5293;
  assign new_P3_U3585 = new_P3_U5299 & new_P3_U5297 & new_P3_U5296;
  assign new_P3_U3586 = new_P3_U3585 & new_P3_U5298;
  assign new_P3_U3587 = new_P3_U5304 & new_P3_U5302 & new_P3_U5301;
  assign new_P3_U3588 = new_P3_U3587 & new_P3_U5303;
  assign new_P3_U3589 = new_P3_U5309 & new_P3_U5307 & new_P3_U5306;
  assign new_P3_U3590 = new_P3_U3589 & new_P3_U5308;
  assign new_P3_U3591 = new_P3_U5314 & new_P3_U5312 & new_P3_U5311;
  assign new_P3_U3592 = new_P3_U3591 & new_P3_U5313;
  assign new_P3_U3593 = new_P3_U5319 & new_P3_U5317 & new_P3_U5316;
  assign new_P3_U3594 = new_P3_U3593 & new_P3_U5318;
  assign new_P3_U3595 = new_P3_U5324 & new_P3_U5322 & new_P3_U5321;
  assign new_P3_U3596 = new_P3_U3595 & new_P3_U5323;
  assign new_P3_U3597 = new_P3_U5329 & new_P3_U5327 & new_P3_U5326;
  assign new_P3_U3598 = new_P3_U3597 & new_P3_U5328;
  assign new_P3_U3599 = new_P3_U5339 & new_P3_U4312;
  assign new_P3_U3600 = new_P3_U5345 & new_P3_U5343 & new_P3_U5342;
  assign new_P3_U3601 = new_P3_U3600 & new_P3_U5344;
  assign new_P3_U3602 = new_P3_U5350 & new_P3_U5348 & new_P3_U5347;
  assign new_P3_U3603 = new_P3_U3602 & new_P3_U5349;
  assign new_P3_U3604 = new_P3_U5355 & new_P3_U5353 & new_P3_U5352;
  assign new_P3_U3605 = new_P3_U3604 & new_P3_U5354;
  assign new_P3_U3606 = new_P3_U5360 & new_P3_U5358 & new_P3_U5357;
  assign new_P3_U3607 = new_P3_U3606 & new_P3_U5359;
  assign new_P3_U3608 = new_P3_U5365 & new_P3_U5363 & new_P3_U5362;
  assign new_P3_U3609 = new_P3_U3608 & new_P3_U5364;
  assign new_P3_U3610 = new_P3_U5370 & new_P3_U5368 & new_P3_U5367;
  assign new_P3_U3611 = new_P3_U3610 & new_P3_U5369;
  assign new_P3_U3612 = new_P3_U5375 & new_P3_U5373 & new_P3_U5372;
  assign new_P3_U3613 = new_P3_U3612 & new_P3_U5374;
  assign new_P3_U3614 = new_P3_U5380 & new_P3_U5378 & new_P3_U5377;
  assign new_P3_U3615 = new_P3_U3614 & new_P3_U5379;
  assign new_P3_U3616 = ~P3_INSTQUEUEWR_ADDR_REG_2_ & ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_U3617 = new_P3_U5390 & new_P3_U4312;
  assign new_P3_U3618 = new_P3_U5396 & new_P3_U5394 & new_P3_U5393;
  assign new_P3_U3619 = new_P3_U3618 & new_P3_U5395;
  assign new_P3_U3620 = new_P3_U5401 & new_P3_U5399 & new_P3_U5398;
  assign new_P3_U3621 = new_P3_U3620 & new_P3_U5400;
  assign new_P3_U3622 = new_P3_U5406 & new_P3_U5404 & new_P3_U5403;
  assign new_P3_U3623 = new_P3_U3622 & new_P3_U5405;
  assign new_P3_U3624 = new_P3_U5411 & new_P3_U5409 & new_P3_U5408;
  assign new_P3_U3625 = new_P3_U3624 & new_P3_U5410;
  assign new_P3_U3626 = new_P3_U5416 & new_P3_U5414 & new_P3_U5413;
  assign new_P3_U3627 = new_P3_U3626 & new_P3_U5415;
  assign new_P3_U3628 = new_P3_U5421 & new_P3_U5419 & new_P3_U5418;
  assign new_P3_U3629 = new_P3_U3628 & new_P3_U5420;
  assign new_P3_U3630 = new_P3_U5426 & new_P3_U5424 & new_P3_U5423;
  assign new_P3_U3631 = new_P3_U3630 & new_P3_U5425;
  assign new_P3_U3632 = new_P3_U5431 & new_P3_U5429 & new_P3_U5428;
  assign new_P3_U3633 = new_P3_U3632 & new_P3_U5430;
  assign new_P3_U3634 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_U3635 = new_P3_U5440 & new_P3_U4312;
  assign new_P3_U3636 = new_P3_U5446 & new_P3_U5444 & new_P3_U5443;
  assign new_P3_U3637 = new_P3_U3636 & new_P3_U5445;
  assign new_P3_U3638 = new_P3_U5451 & new_P3_U5449 & new_P3_U5448;
  assign new_P3_U3639 = new_P3_U3638 & new_P3_U5450;
  assign new_P3_U3640 = new_P3_U5456 & new_P3_U5454 & new_P3_U5453;
  assign new_P3_U3641 = new_P3_U3640 & new_P3_U5455;
  assign new_P3_U3642 = new_P3_U5461 & new_P3_U5459 & new_P3_U5458;
  assign new_P3_U3643 = new_P3_U3642 & new_P3_U5460;
  assign new_P3_U3644 = new_P3_U5466 & new_P3_U5464 & new_P3_U5463;
  assign new_P3_U3645 = new_P3_U3644 & new_P3_U5465;
  assign new_P3_U3646 = new_P3_U5471 & new_P3_U5469 & new_P3_U5468;
  assign new_P3_U3647 = new_P3_U3646 & new_P3_U5470;
  assign new_P3_U3648 = new_P3_U5476 & new_P3_U5474 & new_P3_U5473;
  assign new_P3_U3649 = new_P3_U3648 & new_P3_U5475;
  assign new_P3_U3650 = new_P3_U5481 & new_P3_U5479 & new_P3_U5478;
  assign new_P3_U3651 = new_P3_U3650 & new_P3_U5480;
  assign new_P3_U3652 = new_P3_U4340 & new_P3_ADD_495_U8;
  assign new_P3_U3653 = P3_FLUSH_REG & P3_STATE2_REG_0_;
  assign new_P3_U3654 = new_P3_U4522 & new_P3_U3104;
  assign new_P3_U3655 = new_P3_U3107 & new_P3_U3118;
  assign new_P3_U3656 = new_P3_U5495 & new_P3_U4333;
  assign new_P3_U3657 = new_P3_U3656 & new_P3_U5494;
  assign new_P3_U3658 = new_P3_U5498 & new_P3_U4330;
  assign new_P3_U3659 = new_P3_U5502 & new_P3_U5501;
  assign new_P3_U3660 = new_P3_U4556 & new_P3_U4539;
  assign new_P3_U3661 = new_P3_U2461 & new_P3_U4297;
  assign new_P3_U3662 = new_P3_U4590 & new_P3_U3101;
  assign new_P3_U3663 = new_P3_U4556 & new_P3_U3101;
  assign new_P3_U3664 = new_P3_U4573 & new_P3_U4324;
  assign new_P3_U3665 = new_P3_U5508 & new_P3_U5511 & new_P3_U5510;
  assign new_P3_U3666 = new_P3_U5520 & new_P3_U5519 & new_P3_U4339;
  assign new_P3_U3667 = new_P3_U3666 & new_P3_U5521 & new_P3_U7978 & new_P3_U7977;
  assign new_P3_U3668 = new_P3_U2517 & new_P3_U5528 & new_P3_U3242;
  assign new_P3_U3669 = P3_INSTQUEUERD_ADDR_REG_1_ & new_P3_U4470;
  assign new_P3_U3670 = P3_INSTQUEUERD_ADDR_REG_3_ & new_P3_U3093;
  assign new_P3_U3671 = new_P3_U3119 & new_P3_U3116 & new_P3_U3117;
  assign new_P3_U3672 = new_P3_U3671 & new_P3_U3245 & new_P3_U3244;
  assign new_P3_U3673 = new_P3_U4505 & new_P3_U2456;
  assign new_P3_U3674 = new_P3_U5533 & new_P3_U5532;
  assign new_P3_U3675 = new_P3_U5538 & new_P3_U5536;
  assign new_P3_U3676 = new_P3_U3675 & new_P3_U3677 & new_P3_U5539;
  assign new_P3_U3677 = new_P3_U5540 & new_P3_U5541;
  assign new_P3_U3678 = new_P3_U5552 & new_P3_U5550;
  assign new_P3_U3679 = new_P3_U3678 & new_P3_U5551;
  assign new_P3_U3680 = new_P3_U5555 & new_P3_U5554;
  assign new_P3_U3681 = new_P3_U3682 & new_P3_U5562;
  assign new_P3_U3682 = new_P3_U5565 & new_P3_U5564;
  assign new_P3_U3683 = new_P3_U5568 & new_P3_U5567;
  assign new_P3_U3684 = new_P3_U5576 & new_P3_U5574;
  assign new_P3_U3685 = new_P3_U5587 & new_P3_U5588;
  assign new_P3_U3686 = new_P3_U5594 & new_P3_U5592;
  assign new_P3_U3687 = new_P3_U5626 & new_P3_U5625 & new_P3_U4333;
  assign new_P3_U3688 = new_P3_U2456 & new_P3_U4296;
  assign new_P3_U3689 = new_P3_U2456 & new_P3_U4323;
  assign new_P3_U3690 = new_P3_U4608 & new_P3_U4556;
  assign new_P3_U3691 = new_P3_U2456 & new_P3_U4590;
  assign new_P3_U3692 = new_P3_U5636 & new_P3_U5635;
  assign new_P3_U3693 = new_P3_U5632 & new_P3_U5633 & new_P3_U3694 & new_P3_U5638 & new_P3_U5637;
  assign new_P3_U3694 = new_P3_U3695 & new_P3_U5641;
  assign new_P3_U3695 = new_P3_U5639 & new_P3_U5640;
  assign new_P3_U3696 = new_P3_U5645 & new_P3_U5646 & new_P3_U5644 & new_P3_U5643 & new_P3_U5642;
  assign new_P3_U3697 = new_P3_U5650 & new_P3_U5651 & new_P3_U5647 & new_P3_U5648 & new_P3_U5649;
  assign new_P3_U3698 = new_P3_U3697 & new_P3_U3696;
  assign new_P3_U3699 = new_P3_U5660 & new_P3_U5659;
  assign new_P3_U3700 = new_P3_U5657 & new_P3_U3701 & new_P3_U5662 & new_P3_U5661;
  assign new_P3_U3701 = new_P3_U3702 & new_P3_U5665;
  assign new_P3_U3702 = new_P3_U5663 & new_P3_U5664;
  assign new_P3_U3703 = new_P3_U5669 & new_P3_U5670 & new_P3_U5668 & new_P3_U5667 & new_P3_U5666;
  assign new_P3_U3704 = new_P3_U5673 & new_P3_U5672 & new_P3_U5674 & new_P3_U5671;
  assign new_P3_U3705 = new_P3_U5675 & new_P3_U3704 & new_P3_U3703;
  assign new_P3_U3706 = new_P3_U3707 & new_P3_U5681;
  assign new_P3_U3707 = new_P3_U5684 & new_P3_U5683;
  assign new_P3_U3708 = new_P3_U3709 & new_P3_U5689;
  assign new_P3_U3709 = new_P3_U5687 & new_P3_U5688;
  assign new_P3_U3710 = new_P3_U3708 & new_P3_U5686 & new_P3_U5685;
  assign new_P3_U3711 = new_P3_U5693 & new_P3_U5694 & new_P3_U5692 & new_P3_U5691 & new_P3_U5690;
  assign new_P3_U3712 = new_P3_U5697 & new_P3_U5696 & new_P3_U5698 & new_P3_U5695;
  assign new_P3_U3713 = new_P3_U5699 & new_P3_U3712 & new_P3_U3711;
  assign new_P3_U3714 = new_P3_U5705 & new_P3_U5704;
  assign new_P3_U3715 = new_P3_U5708 & new_P3_U5707;
  assign new_P3_U3716 = new_P3_U3717 & new_P3_U5713;
  assign new_P3_U3717 = new_P3_U5711 & new_P3_U5712;
  assign new_P3_U3718 = new_P3_U3716 & new_P3_U5710 & new_P3_U5709;
  assign new_P3_U3719 = new_P3_U5717 & new_P3_U5718 & new_P3_U5716 & new_P3_U5715 & new_P3_U5714;
  assign new_P3_U3720 = new_P3_U5721 & new_P3_U5720 & new_P3_U5722 & new_P3_U5719;
  assign new_P3_U3721 = new_P3_U5723 & new_P3_U3720 & new_P3_U3719;
  assign new_P3_U3722 = new_P3_U3723 & new_P3_U5729;
  assign new_P3_U3723 = new_P3_U5732 & new_P3_U5731;
  assign new_P3_U3724 = new_P3_U3725 & new_P3_U5737;
  assign new_P3_U3725 = new_P3_U5735 & new_P3_U5736;
  assign new_P3_U3726 = new_P3_U3724 & new_P3_U5734 & new_P3_U5733;
  assign new_P3_U3727 = new_P3_U5741 & new_P3_U5742 & new_P3_U5740 & new_P3_U5739 & new_P3_U5738;
  assign new_P3_U3728 = new_P3_U5745 & new_P3_U5744 & new_P3_U5746 & new_P3_U5743;
  assign new_P3_U3729 = new_P3_U5747 & new_P3_U3728 & new_P3_U3727;
  assign new_P3_U3730 = new_P3_U3731 & new_P3_U5752;
  assign new_P3_U3731 = new_P3_U5756 & new_P3_U5755;
  assign new_P3_U3732 = new_P3_U3733 & new_P3_U5761;
  assign new_P3_U3733 = new_P3_U5759 & new_P3_U5760;
  assign new_P3_U3734 = new_P3_U3732 & new_P3_U5758 & new_P3_U5757;
  assign new_P3_U3735 = new_P3_U5765 & new_P3_U5766 & new_P3_U5764 & new_P3_U5763 & new_P3_U5762;
  assign new_P3_U3736 = new_P3_U5769 & new_P3_U5768 & new_P3_U5770 & new_P3_U5767;
  assign new_P3_U3737 = new_P3_U5771 & new_P3_U3736 & new_P3_U3735;
  assign new_P3_U3738 = new_P3_U3739 & new_P3_U5776;
  assign new_P3_U3739 = new_P3_U5780 & new_P3_U5779;
  assign new_P3_U3740 = new_P3_U3741 & new_P3_U5785;
  assign new_P3_U3741 = new_P3_U5783 & new_P3_U5784;
  assign new_P3_U3742 = new_P3_U3740 & new_P3_U5782 & new_P3_U5781;
  assign new_P3_U3743 = new_P3_U5789 & new_P3_U5790 & new_P3_U5788 & new_P3_U5787 & new_P3_U5786;
  assign new_P3_U3744 = new_P3_U5793 & new_P3_U5792 & new_P3_U5794 & new_P3_U5791;
  assign new_P3_U3745 = new_P3_U5795 & new_P3_U3744 & new_P3_U3743;
  assign new_P3_U3746 = new_P3_U3747 & new_P3_U5800;
  assign new_P3_U3747 = new_P3_U5804 & new_P3_U5803;
  assign new_P3_U3748 = new_P3_U3749 & new_P3_U5809;
  assign new_P3_U3749 = new_P3_U5807 & new_P3_U5808;
  assign new_P3_U3750 = new_P3_U3748 & new_P3_U5806 & new_P3_U5805;
  assign new_P3_U3751 = new_P3_U5813 & new_P3_U5814 & new_P3_U5812 & new_P3_U5811 & new_P3_U5810;
  assign new_P3_U3752 = new_P3_U5817 & new_P3_U5816 & new_P3_U5818 & new_P3_U5815;
  assign new_P3_U3753 = new_P3_U5819 & new_P3_U3752 & new_P3_U3751;
  assign new_P3_U3754 = new_P3_U3755 & new_P3_U5824;
  assign new_P3_U3755 = new_P3_U5828 & new_P3_U5827;
  assign new_P3_U3756 = new_P3_U5831 & new_P3_U5833 & new_P3_U5832;
  assign new_P3_U3757 = new_P3_U3756 & new_P3_U5830 & new_P3_U5829;
  assign new_P3_U3758 = new_P3_U5837 & new_P3_U5838 & new_P3_U5836 & new_P3_U5835 & new_P3_U5834;
  assign new_P3_U3759 = new_P3_U5839 & new_P3_U5840 & new_P3_U5842 & new_P3_U5841;
  assign new_P3_U3760 = new_P3_U5843 & new_P3_U3759 & new_P3_U3758;
  assign new_P3_U3761 = new_P3_U3762 & new_P3_U5848;
  assign new_P3_U3762 = new_P3_U5852 & new_P3_U5851;
  assign new_P3_U3763 = new_P3_U5857 & new_P3_U5856;
  assign new_P3_U3764 = new_P3_U3763 & new_P3_U5855 & new_P3_U5854 & new_P3_U5853;
  assign new_P3_U3765 = new_P3_U5861 & new_P3_U5862 & new_P3_U5860 & new_P3_U5859 & new_P3_U5858;
  assign new_P3_U3766 = new_P3_U5863 & new_P3_U5864 & new_P3_U5866 & new_P3_U5865;
  assign new_P3_U3767 = new_P3_U5867 & new_P3_U3766 & new_P3_U3765;
  assign new_P3_U3768 = new_P3_U3769 & new_P3_U5873;
  assign new_P3_U3769 = new_P3_U5876 & new_P3_U5875;
  assign new_P3_U3770 = new_P3_U5881 & new_P3_U5880;
  assign new_P3_U3771 = new_P3_U3770 & new_P3_U5879 & new_P3_U5878 & new_P3_U5877;
  assign new_P3_U3772 = new_P3_U5885 & new_P3_U5886 & new_P3_U5884 & new_P3_U5883 & new_P3_U5882;
  assign new_P3_U3773 = new_P3_U5887 & new_P3_U5888 & new_P3_U5890 & new_P3_U5889;
  assign new_P3_U3774 = new_P3_U5891 & new_P3_U3773 & new_P3_U3772;
  assign new_P3_U3775 = new_P3_U3776 & new_P3_U5897;
  assign new_P3_U3776 = new_P3_U5900 & new_P3_U5899;
  assign new_P3_U3777 = new_P3_U5905 & new_P3_U5904;
  assign new_P3_U3778 = new_P3_U3777 & new_P3_U5903 & new_P3_U5902 & new_P3_U5901;
  assign new_P3_U3779 = new_P3_U5909 & new_P3_U5910 & new_P3_U5908 & new_P3_U5907 & new_P3_U5906;
  assign new_P3_U3780 = new_P3_U5911 & new_P3_U5912 & new_P3_U5914 & new_P3_U5913;
  assign new_P3_U3781 = new_P3_U5915 & new_P3_U3780 & new_P3_U3779;
  assign new_P3_U3782 = new_P3_U3783 & new_P3_U5920;
  assign new_P3_U3783 = new_P3_U5924 & new_P3_U5923;
  assign new_P3_U3784 = new_P3_U5929 & new_P3_U5928;
  assign new_P3_U3785 = new_P3_U3784 & new_P3_U5927 & new_P3_U5926 & new_P3_U5925;
  assign new_P3_U3786 = new_P3_U5933 & new_P3_U5934 & new_P3_U5932 & new_P3_U5931 & new_P3_U5930;
  assign new_P3_U3787 = new_P3_U5935 & new_P3_U5936 & new_P3_U5938 & new_P3_U5937;
  assign new_P3_U3788 = new_P3_U5939 & new_P3_U3787 & new_P3_U3786;
  assign new_P3_U3789 = new_P3_U3790 & new_P3_U5944;
  assign new_P3_U3790 = new_P3_U5948 & new_P3_U5947;
  assign new_P3_U3791 = new_P3_U5953 & new_P3_U5952;
  assign new_P3_U3792 = new_P3_U3791 & new_P3_U5951 & new_P3_U5950 & new_P3_U5949;
  assign new_P3_U3793 = new_P3_U5957 & new_P3_U5958 & new_P3_U5956 & new_P3_U5955 & new_P3_U5954;
  assign new_P3_U3794 = new_P3_U5959 & new_P3_U5960 & new_P3_U5962 & new_P3_U5961;
  assign new_P3_U3795 = new_P3_U5963 & new_P3_U3794 & new_P3_U3793;
  assign new_P3_U3796 = new_P3_U5972 & new_P3_U5971;
  assign new_P3_U3797 = new_P3_U5977 & new_P3_U5976;
  assign new_P3_U3798 = new_P3_U3797 & new_P3_U5975 & new_P3_U5974 & new_P3_U5973;
  assign new_P3_U3799 = new_P3_U5968 & new_P3_U5969 & new_P3_U3798 & new_P3_U3796 & new_P3_U5970;
  assign new_P3_U3800 = new_P3_U5981 & new_P3_U5982 & new_P3_U5980 & new_P3_U5979 & new_P3_U5978;
  assign new_P3_U3801 = new_P3_U5983 & new_P3_U5984 & new_P3_U5986 & new_P3_U5985;
  assign new_P3_U3802 = new_P3_U5987 & new_P3_U3801 & new_P3_U3800;
  assign new_P3_U3803 = new_P3_U5991 & new_P3_U5989;
  assign new_P3_U3804 = new_P3_U5996 & new_P3_U5995;
  assign new_P3_U3805 = new_P3_U6001 & new_P3_U6000;
  assign new_P3_U3806 = new_P3_U3805 & new_P3_U5999 & new_P3_U5998 & new_P3_U5997;
  assign new_P3_U3807 = new_P3_U5992 & new_P3_U5993 & new_P3_U3806 & new_P3_U3804 & new_P3_U5994;
  assign new_P3_U3808 = new_P3_U6005 & new_P3_U6006 & new_P3_U6004 & new_P3_U6003 & new_P3_U6002;
  assign new_P3_U3809 = new_P3_U6007 & new_P3_U6008 & new_P3_U6010 & new_P3_U6009;
  assign new_P3_U3810 = new_P3_U6011 & new_P3_U3809 & new_P3_U3808;
  assign new_P3_U3811 = new_P3_U6015 & new_P3_U6013;
  assign new_P3_U3812 = new_P3_U3813 & new_P3_U6017;
  assign new_P3_U3813 = new_P3_U6020 & new_P3_U6019;
  assign new_P3_U3814 = new_P3_U6025 & new_P3_U6024;
  assign new_P3_U3815 = new_P3_U3814 & new_P3_U6023 & new_P3_U6022 & new_P3_U6021;
  assign new_P3_U3816 = new_P3_U6029 & new_P3_U6030 & new_P3_U6028 & new_P3_U6027 & new_P3_U6026;
  assign new_P3_U3817 = new_P3_U6031 & new_P3_U6032 & new_P3_U6034 & new_P3_U6033;
  assign new_P3_U3818 = new_P3_U6035 & new_P3_U3817 & new_P3_U3816;
  assign new_P3_U3819 = new_P3_U6044 & new_P3_U6043;
  assign new_P3_U3820 = new_P3_U6041 & new_P3_U3821 & new_P3_U6047 & new_P3_U6046 & new_P3_U6045;
  assign new_P3_U3821 = new_P3_U6049 & new_P3_U6048;
  assign new_P3_U3822 = new_P3_U6053 & new_P3_U6054 & new_P3_U6052 & new_P3_U6051 & new_P3_U6050;
  assign new_P3_U3823 = new_P3_U6055 & new_P3_U6056 & new_P3_U6058 & new_P3_U6057;
  assign new_P3_U3824 = new_P3_U6059 & new_P3_U3823 & new_P3_U3822;
  assign new_P3_U3825 = new_P3_U3826 & new_P3_U6065;
  assign new_P3_U3826 = new_P3_U6068 & new_P3_U6067;
  assign new_P3_U3827 = new_P3_U6073 & new_P3_U6072;
  assign new_P3_U3828 = new_P3_U3827 & new_P3_U6071 & new_P3_U6070 & new_P3_U6069;
  assign new_P3_U3829 = new_P3_U6077 & new_P3_U6078 & new_P3_U6076 & new_P3_U6075 & new_P3_U6074;
  assign new_P3_U3830 = new_P3_U6079 & new_P3_U6080 & new_P3_U6082 & new_P3_U6081;
  assign new_P3_U3831 = new_P3_U6083 & new_P3_U3830 & new_P3_U3829;
  assign new_P3_U3832 = new_P3_U6092 & new_P3_U6091;
  assign new_P3_U3833 = new_P3_U6089 & new_P3_U3834 & new_P3_U6095 & new_P3_U6094 & new_P3_U6093;
  assign new_P3_U3834 = new_P3_U6097 & new_P3_U6096;
  assign new_P3_U3835 = new_P3_U6101 & new_P3_U6102 & new_P3_U6100 & new_P3_U6099 & new_P3_U6098;
  assign new_P3_U3836 = new_P3_U6103 & new_P3_U6104 & new_P3_U6106 & new_P3_U6105;
  assign new_P3_U3837 = new_P3_U6107 & new_P3_U3836 & new_P3_U3835;
  assign new_P3_U3838 = new_P3_U6116 & new_P3_U6115;
  assign new_P3_U3839 = new_P3_U6121 & new_P3_U6120;
  assign new_P3_U3840 = new_P3_U3839 & new_P3_U6119 & new_P3_U6118 & new_P3_U6117;
  assign new_P3_U3841 = new_P3_U3844 & new_P3_U6112 & new_P3_U3840 & new_P3_U6114 & new_P3_U3838;
  assign new_P3_U3842 = new_P3_U6125 & new_P3_U6126 & new_P3_U6124 & new_P3_U6123 & new_P3_U6122;
  assign new_P3_U3843 = new_P3_U6127 & new_P3_U6128 & new_P3_U6130 & new_P3_U6129;
  assign new_P3_U3844 = new_P3_U6131 & new_P3_U3843 & new_P3_U3842;
  assign new_P3_U3845 = new_P3_U6135 & new_P3_U6133;
  assign new_P3_U3846 = new_P3_U6140 & new_P3_U6139;
  assign new_P3_U3847 = new_P3_U6145 & new_P3_U6144;
  assign new_P3_U3848 = new_P3_U3847 & new_P3_U6143 & new_P3_U6142 & new_P3_U6141;
  assign new_P3_U3849 = new_P3_U3852 & new_P3_U6136 & new_P3_U3848 & new_P3_U6138 & new_P3_U3846;
  assign new_P3_U3850 = new_P3_U6149 & new_P3_U6150 & new_P3_U6148 & new_P3_U6147 & new_P3_U6146;
  assign new_P3_U3851 = new_P3_U6151 & new_P3_U6152 & new_P3_U6154 & new_P3_U6153;
  assign new_P3_U3852 = new_P3_U6155 & new_P3_U3850 & new_P3_U3851;
  assign new_P3_U3853 = new_P3_U6159 & new_P3_U6157;
  assign new_P3_U3854 = new_P3_U6164 & new_P3_U6163;
  assign new_P3_U3855 = new_P3_U6169 & new_P3_U6168;
  assign new_P3_U3856 = new_P3_U3855 & new_P3_U6167 & new_P3_U6166 & new_P3_U6165;
  assign new_P3_U3857 = new_P3_U6160 & new_P3_U3856 & new_P3_U3854 & new_P3_U6161 & new_P3_U6162;
  assign new_P3_U3858 = new_P3_U6172 & new_P3_U6171 & new_P3_U6170;
  assign new_P3_U3859 = new_P3_U6174 & new_P3_U6173;
  assign new_P3_U3860 = new_P3_U6177 & new_P3_U6176 & new_P3_U6175;
  assign new_P3_U3861 = new_P3_U6179 & new_P3_U6178;
  assign new_P3_U3862 = new_P3_U3861 & new_P3_U3860 & new_P3_U3859 & new_P3_U3858;
  assign new_P3_U3863 = new_P3_U6183 & new_P3_U6181;
  assign new_P3_U3864 = new_P3_U6188 & new_P3_U6187;
  assign new_P3_U3865 = new_P3_U6193 & new_P3_U6192;
  assign new_P3_U3866 = new_P3_U3865 & new_P3_U6191 & new_P3_U6190 & new_P3_U6189;
  assign new_P3_U3867 = new_P3_U6184 & new_P3_U3866 & new_P3_U3864 & new_P3_U6185 & new_P3_U6186;
  assign new_P3_U3868 = new_P3_U6196 & new_P3_U6195 & new_P3_U6194;
  assign new_P3_U3869 = new_P3_U6198 & new_P3_U6197;
  assign new_P3_U3870 = new_P3_U6201 & new_P3_U6200 & new_P3_U6199;
  assign new_P3_U3871 = new_P3_U6203 & new_P3_U6202;
  assign new_P3_U3872 = new_P3_U3871 & new_P3_U3870 & new_P3_U3869 & new_P3_U3868;
  assign new_P3_U3873 = new_P3_U6207 & new_P3_U6205;
  assign new_P3_U3874 = new_P3_U6212 & new_P3_U6211;
  assign new_P3_U3875 = new_P3_U6217 & new_P3_U6216;
  assign new_P3_U3876 = new_P3_U3875 & new_P3_U6215 & new_P3_U6214 & new_P3_U6213;
  assign new_P3_U3877 = new_P3_U3876 & new_P3_U6208 & new_P3_U3874 & new_P3_U6209 & new_P3_U6210;
  assign new_P3_U3878 = new_P3_U6220 & new_P3_U6219 & new_P3_U6218;
  assign new_P3_U3879 = new_P3_U6222 & new_P3_U6221;
  assign new_P3_U3880 = new_P3_U6225 & new_P3_U6224 & new_P3_U6223;
  assign new_P3_U3881 = new_P3_U6227 & new_P3_U6226;
  assign new_P3_U3882 = new_P3_U3880 & new_P3_U3881 & new_P3_U3879 & new_P3_U3878;
  assign new_P3_U3883 = new_P3_U6231 & new_P3_U6229;
  assign new_P3_U3884 = new_P3_U6236 & new_P3_U6235;
  assign new_P3_U3885 = new_P3_U6241 & new_P3_U6240;
  assign new_P3_U3886 = new_P3_U3885 & new_P3_U6239 & new_P3_U6238 & new_P3_U6237;
  assign new_P3_U3887 = new_P3_U3886 & new_P3_U3884 & new_P3_U6232 & new_P3_U6233 & new_P3_U6234;
  assign new_P3_U3888 = new_P3_U6244 & new_P3_U6243 & new_P3_U6242;
  assign new_P3_U3889 = new_P3_U6246 & new_P3_U6245;
  assign new_P3_U3890 = new_P3_U6249 & new_P3_U6248 & new_P3_U6247;
  assign new_P3_U3891 = new_P3_U6251 & new_P3_U6250;
  assign new_P3_U3892 = new_P3_U3890 & new_P3_U3891 & new_P3_U3889 & new_P3_U3888;
  assign new_P3_U3893 = new_P3_U6255 & new_P3_U6253;
  assign new_P3_U3894 = new_P3_U6257 & new_P3_U6256;
  assign new_P3_U3895 = new_P3_U6260 & new_P3_U6259;
  assign new_P3_U3896 = new_P3_U6265 & new_P3_U6264;
  assign new_P3_U3897 = new_P3_U3896 & new_P3_U6263 & new_P3_U6262 & new_P3_U6261;
  assign new_P3_U3898 = new_P3_U6268 & new_P3_U6267 & new_P3_U6266;
  assign new_P3_U3899 = new_P3_U6270 & new_P3_U6269;
  assign new_P3_U3900 = new_P3_U6273 & new_P3_U6272 & new_P3_U6271;
  assign new_P3_U3901 = new_P3_U6275 & new_P3_U6274;
  assign new_P3_U3902 = new_P3_U3900 & new_P3_U3901 & new_P3_U3899 & new_P3_U3898;
  assign new_P3_U3903 = new_P3_U6281 & new_P3_U6280;
  assign new_P3_U3904 = new_P3_U6284 & new_P3_U6283;
  assign new_P3_U3905 = new_P3_U6289 & new_P3_U6288;
  assign new_P3_U3906 = new_P3_U3905 & new_P3_U6287 & new_P3_U6286 & new_P3_U6285;
  assign new_P3_U3907 = new_P3_U6292 & new_P3_U6291 & new_P3_U6290;
  assign new_P3_U3908 = new_P3_U6294 & new_P3_U6293;
  assign new_P3_U3909 = new_P3_U6297 & new_P3_U6296 & new_P3_U6295;
  assign new_P3_U3910 = new_P3_U6299 & new_P3_U6298;
  assign new_P3_U3911 = new_P3_U3909 & new_P3_U3910 & new_P3_U3908 & new_P3_U3907;
  assign new_P3_U3912 = new_P3_U6305 & new_P3_U6304;
  assign new_P3_U3913 = new_P3_U6308 & new_P3_U6307;
  assign new_P3_U3914 = new_P3_U6313 & new_P3_U6312;
  assign new_P3_U3915 = new_P3_U3914 & new_P3_U6311 & new_P3_U6310 & new_P3_U6309;
  assign new_P3_U3916 = new_P3_U6316 & new_P3_U6315 & new_P3_U6314;
  assign new_P3_U3917 = new_P3_U6318 & new_P3_U6317;
  assign new_P3_U3918 = new_P3_U6321 & new_P3_U6320 & new_P3_U6319;
  assign new_P3_U3919 = new_P3_U6323 & new_P3_U6322;
  assign new_P3_U3920 = new_P3_U3918 & new_P3_U3919 & new_P3_U3917 & new_P3_U3916;
  assign new_P3_U3921 = new_P3_U6329 & new_P3_U6328;
  assign new_P3_U3922 = new_P3_U6332 & new_P3_U6331;
  assign new_P3_U3923 = new_P3_U6337 & new_P3_U6336;
  assign new_P3_U3924 = new_P3_U3923 & new_P3_U6335 & new_P3_U6334 & new_P3_U6333;
  assign new_P3_U3925 = new_P3_U6340 & new_P3_U6339 & new_P3_U6338;
  assign new_P3_U3926 = new_P3_U6342 & new_P3_U6341;
  assign new_P3_U3927 = new_P3_U6345 & new_P3_U6344 & new_P3_U6343;
  assign new_P3_U3928 = new_P3_U6347 & new_P3_U6346;
  assign new_P3_U3929 = new_P3_U3927 & new_P3_U3928 & new_P3_U3926 & new_P3_U3925;
  assign new_P3_U3930 = new_P3_U6353 & new_P3_U6352;
  assign new_P3_U3931 = new_P3_U6356 & new_P3_U6355;
  assign new_P3_U3932 = new_P3_U6361 & new_P3_U6360;
  assign new_P3_U3933 = new_P3_U3932 & new_P3_U6359 & new_P3_U6358 & new_P3_U6357;
  assign new_P3_U3934 = new_P3_U6364 & new_P3_U6363 & new_P3_U6362;
  assign new_P3_U3935 = new_P3_U6366 & new_P3_U6365;
  assign new_P3_U3936 = new_P3_U6369 & new_P3_U6368 & new_P3_U6367;
  assign new_P3_U3937 = new_P3_U6371 & new_P3_U6370;
  assign new_P3_U3938 = new_P3_U3936 & new_P3_U3937 & new_P3_U3935 & new_P3_U3934;
  assign new_P3_U3939 = new_P3_U6398 & new_P3_U3247;
  assign new_P3_U3940 = new_P3_U6377 & new_P3_U6376;
  assign new_P3_U3941 = new_P3_U6380 & new_P3_U6379;
  assign new_P3_U3942 = new_P3_U3941 & new_P3_U6381;
  assign new_P3_U3943 = new_P3_U6384 & new_P3_U6386 & new_P3_U6385;
  assign new_P3_U3944 = new_P3_U3943 & new_P3_U6383 & new_P3_U6382;
  assign new_P3_U3945 = new_P3_U3944 & new_P3_U3942 & new_P3_U3940 & new_P3_U6378;
  assign new_P3_U3946 = new_P3_U6389 & new_P3_U6388 & new_P3_U6387;
  assign new_P3_U3947 = new_P3_U6391 & new_P3_U6390;
  assign new_P3_U3948 = new_P3_U3947 & new_P3_U3946 & new_P3_U6392;
  assign new_P3_U3949 = new_P3_U6394 & new_P3_U6393;
  assign new_P3_U3950 = new_P3_U3948 & new_P3_U3949 & new_P3_U6395 & new_P3_U6398 & new_P3_U6397;
  assign new_P3_U3951 = P3_STATE2_REG_0_ & new_P3_U3104;
  assign new_P3_U3952 = P3_STATE2_REG_2_ & new_P3_U3121;
  assign new_P3_U3953 = new_P3_U4505 & P3_STATE2_REG_0_;
  assign new_P3_U3954 = new_P3_U6409 & new_P3_U6410 & new_P3_U6412 & new_P3_U6411;
  assign new_P3_U3955 = new_P3_U6417 & new_P3_U6418 & new_P3_U6420 & new_P3_U6419;
  assign new_P3_U3956 = new_P3_U6427 & new_P3_U6428 & new_P3_U6426 & new_P3_U6425;
  assign new_P3_U3957 = new_P3_U6435 & new_P3_U6436 & new_P3_U6434 & new_P3_U6433;
  assign new_P3_U3958 = new_P3_U6443 & new_P3_U6444 & new_P3_U6442 & new_P3_U6441;
  assign new_P3_U3959 = new_P3_U6451 & new_P3_U6452 & new_P3_U6450 & new_P3_U6449;
  assign new_P3_U3960 = new_P3_U6459 & new_P3_U6460 & new_P3_U6458 & new_P3_U6457;
  assign new_P3_U3961 = new_P3_U6467 & new_P3_U6468 & new_P3_U6466 & new_P3_U6465;
  assign new_P3_U3962 = new_P3_U6475 & new_P3_U6476 & new_P3_U6474 & new_P3_U6473;
  assign new_P3_U3963 = new_P3_U6483 & new_P3_U6484 & new_P3_U6482 & new_P3_U6481;
  assign new_P3_U3964 = new_P3_U6491 & new_P3_U6492 & new_P3_U6490 & new_P3_U6489;
  assign new_P3_U3965 = new_P3_U6499 & new_P3_U6500 & new_P3_U6498 & new_P3_U6497;
  assign new_P3_U3966 = new_P3_U6507 & new_P3_U6506 & new_P3_U6508 & new_P3_U6505;
  assign new_P3_U3967 = new_P3_U6515 & new_P3_U6514 & new_P3_U6516 & new_P3_U6513;
  assign new_P3_U3968 = new_P3_U6523 & new_P3_U6522 & new_P3_U6524 & new_P3_U6521;
  assign new_P3_U3969 = new_P3_U6531 & new_P3_U6530 & new_P3_U6532 & new_P3_U6529;
  assign new_P3_U3970 = new_P3_U6539 & new_P3_U6538 & new_P3_U6540 & new_P3_U6537;
  assign new_P3_U3971 = new_P3_U6547 & new_P3_U6546 & new_P3_U6548 & new_P3_U6545;
  assign new_P3_U3972 = new_P3_U6555 & new_P3_U6554 & new_P3_U6556 & new_P3_U6553;
  assign new_P3_U3973 = new_P3_U6563 & new_P3_U6562 & new_P3_U6564 & new_P3_U6561;
  assign new_P3_U3974 = new_P3_U6571 & new_P3_U6570 & new_P3_U6572 & new_P3_U6569;
  assign new_P3_U3975 = new_P3_U6579 & new_P3_U6578 & new_P3_U6580 & new_P3_U6577;
  assign new_P3_U3976 = new_P3_U6587 & new_P3_U6586 & new_P3_U6588 & new_P3_U6585;
  assign new_P3_U3977 = new_P3_U6595 & new_P3_U6594 & new_P3_U6596 & new_P3_U6593;
  assign new_P3_U3978 = new_P3_U6603 & new_P3_U6602 & new_P3_U6604 & new_P3_U6601;
  assign new_P3_U3979 = new_P3_U6611 & new_P3_U6610 & new_P3_U6612 & new_P3_U6609;
  assign new_P3_U3980 = new_P3_U6617 & new_P3_U6618 & new_P3_U6620 & new_P3_U6619;
  assign new_P3_U3981 = new_P3_U6625 & new_P3_U6626 & new_P3_U6628 & new_P3_U6627;
  assign new_P3_U3982 = new_P3_U6633 & new_P3_U6634 & new_P3_U6636 & new_P3_U6635;
  assign new_P3_U3983 = new_P3_U6642 & new_P3_U6643 & new_P3_U6644 & new_P3_U6641;
  assign new_P3_U3984 = new_P3_U6650 & new_P3_U6651 & new_P3_U6652 & new_P3_U6649;
  assign new_P3_U3985 = new_P3_U6658 & new_P3_U6659 & new_P3_U6660 & new_P3_U6657;
  assign new_P3_U3986 = new_P3_U4293 & new_P3_U2390;
  assign new_P3_U3987 = new_P3_U6809 & new_P3_U6810;
  assign new_P3_U3988 = new_P3_U6812 & new_P3_U6813;
  assign new_P3_U3989 = new_P3_U6815 & new_P3_U6816;
  assign new_P3_U3990 = new_P3_U6818 & new_P3_U6819;
  assign new_P3_U3991 = new_P3_U6821 & new_P3_U6822;
  assign new_P3_U3992 = new_P3_U6824 & new_P3_U6825;
  assign new_P3_U3993 = new_P3_U6827 & new_P3_U6828;
  assign new_P3_U3994 = new_P3_U6830 & new_P3_U6831;
  assign new_P3_U3995 = new_P3_U6833 & new_P3_U6834;
  assign new_P3_U3996 = new_P3_U6836 & new_P3_U6837;
  assign new_P3_U3997 = new_P3_U6839 & new_P3_U6840;
  assign new_P3_U3998 = new_P3_U6842 & new_P3_U6843;
  assign new_P3_U3999 = new_P3_U6845 & new_P3_U6846;
  assign new_P3_U4000 = new_P3_U6848 & new_P3_U6849;
  assign new_P3_U4001 = new_P3_U6851 & new_P3_U6852;
  assign new_P3_U4002 = new_P3_U6857 & new_P3_U6856;
  assign new_P3_U4003 = new_P3_U6861 & new_P3_U6860;
  assign new_P3_U4004 = new_P3_U6865 & new_P3_U6864;
  assign new_P3_U4005 = new_P3_U6869 & new_P3_U6868;
  assign new_P3_U4006 = new_P3_U6873 & new_P3_U6872;
  assign new_P3_U4007 = new_P3_U6877 & new_P3_U6876;
  assign new_P3_U4008 = new_P3_U6881 & new_P3_U6880;
  assign new_P3_U4009 = new_P3_U6885 & new_P3_U6884;
  assign new_P3_U4010 = new_P3_U6889 & new_P3_U6888;
  assign new_P3_U4011 = new_P3_U6893 & new_P3_U6892;
  assign new_P3_U4012 = new_P3_U6897 & new_P3_U6896;
  assign new_P3_U4013 = new_P3_U6901 & new_P3_U6900;
  assign new_P3_U4014 = new_P3_U6905 & new_P3_U6904;
  assign new_P3_U4015 = new_P3_U6907 & new_P3_U6909;
  assign new_P3_U4016 = new_P3_U6911 & new_P3_U6913;
  assign new_P3_U4017 = new_P3_U6915 & new_P3_U6917;
  assign new_P3_U4018 = new_P3_U6922 & new_P3_U6920;
  assign new_P3_U4019 = new_P3_U6927 & new_P3_U6925;
  assign new_P3_U4020 = new_P3_U6932 & new_P3_U6930;
  assign new_P3_U4021 = new_P3_U6937 & new_P3_U6935;
  assign new_P3_U4022 = new_P3_U6942 & new_P3_U6940;
  assign new_P3_U4023 = new_P3_U6947 & new_P3_U6945;
  assign new_P3_U4024 = new_P3_U6952 & new_P3_U6950;
  assign new_P3_U4025 = new_P3_U6957 & new_P3_U6955;
  assign new_P3_U4026 = new_P3_U6962 & new_P3_U6960;
  assign new_P3_U4027 = new_P3_U6967 & new_P3_U6965;
  assign new_P3_U4028 = new_P3_U6972 & new_P3_U6970;
  assign new_P3_U4029 = new_P3_U6977 & new_P3_U6975;
  assign new_P3_U4030 = new_P3_U4336 & new_P3_U4329 & new_P3_U4328;
  assign new_P3_U4031 = new_P3_U4032 & new_P3_U7098 & new_P3_U7097;
  assign new_P3_U4032 = new_P3_U7101 & new_P3_U7100;
  assign new_P3_U4033 = new_P3_U4034 & new_P3_U7104;
  assign new_P3_U4034 = new_P3_U7106 & new_P3_U7105;
  assign new_P3_U4035 = new_P3_U4036 & new_P3_U7108 & new_P3_U7107;
  assign new_P3_U4036 = new_P3_U7111 & new_P3_U7110;
  assign new_P3_U4037 = new_P3_U4038 & new_P3_U7114;
  assign new_P3_U4038 = new_P3_U7116 & new_P3_U7115;
  assign new_P3_U4039 = new_P3_U4040 & new_P3_U7118 & new_P3_U7117;
  assign new_P3_U4040 = new_P3_U7121 & new_P3_U7120;
  assign new_P3_U4041 = new_P3_U4042 & new_P3_U7124;
  assign new_P3_U4042 = new_P3_U7126 & new_P3_U7125;
  assign new_P3_U4043 = new_P3_U4044 & new_P3_U7128 & new_P3_U7127;
  assign new_P3_U4044 = new_P3_U7131 & new_P3_U7130;
  assign new_P3_U4045 = new_P3_U4046 & new_P3_U7134;
  assign new_P3_U4046 = new_P3_U7136 & new_P3_U7135;
  assign new_P3_U4047 = new_P3_U7138 & new_P3_U7137 & new_P3_U4316;
  assign new_P3_U4048 = new_P3_U7140 & new_P3_U7141;
  assign new_P3_U4049 = new_P3_U4050 & new_P3_U7144;
  assign new_P3_U4050 = new_P3_U7146 & new_P3_U7145;
  assign new_P3_U4051 = new_P3_U7143 & new_P3_U7142 & new_P3_U4047 & new_P3_U4048 & new_P3_U7139;
  assign new_P3_U4052 = new_P3_U7148 & new_P3_U7147 & new_P3_U4316;
  assign new_P3_U4053 = new_P3_U7150 & new_P3_U7151;
  assign new_P3_U4054 = new_P3_U4055 & new_P3_U7154;
  assign new_P3_U4055 = new_P3_U7156 & new_P3_U7155;
  assign new_P3_U4056 = new_P3_U7153 & new_P3_U7152 & new_P3_U4052 & new_P3_U4053 & new_P3_U7149;
  assign new_P3_U4057 = new_P3_U7158 & new_P3_U7157 & new_P3_U4316;
  assign new_P3_U4058 = new_P3_U4059 & new_P3_U7161;
  assign new_P3_U4059 = new_P3_U7164 & new_P3_U7163;
  assign new_P3_U4060 = new_P3_U7166 & new_P3_U7165 & new_P3_U4316;
  assign new_P3_U4061 = new_P3_U4062 & new_P3_U7169;
  assign new_P3_U4062 = new_P3_U7172 & new_P3_U7171;
  assign new_P3_U4063 = new_P3_U7174 & new_P3_U7173 & new_P3_U4316;
  assign new_P3_U4064 = new_P3_U4065 & new_P3_U7177;
  assign new_P3_U4065 = new_P3_U7180 & new_P3_U7179;
  assign new_P3_U4066 = new_P3_U7182 & new_P3_U7181 & new_P3_U4316;
  assign new_P3_U4067 = new_P3_U4068 & new_P3_U7185;
  assign new_P3_U4068 = new_P3_U7188 & new_P3_U7187;
  assign new_P3_U4069 = new_P3_U7190 & new_P3_U7189 & new_P3_U4316;
  assign new_P3_U4070 = new_P3_U4071 & new_P3_U7193;
  assign new_P3_U4071 = new_P3_U7196 & new_P3_U7195;
  assign new_P3_U4072 = new_P3_U7198 & new_P3_U7197 & new_P3_U4316;
  assign new_P3_U4073 = new_P3_U4074 & new_P3_U7201;
  assign new_P3_U4074 = new_P3_U7204 & new_P3_U7203;
  assign new_P3_U4075 = new_P3_U7206 & new_P3_U7205 & new_P3_U4316;
  assign new_P3_U4076 = new_P3_U4077 & new_P3_U7209;
  assign new_P3_U4077 = new_P3_U7212 & new_P3_U7211;
  assign new_P3_U4078 = new_P3_U7214 & new_P3_U7213 & new_P3_U4316;
  assign new_P3_U4079 = new_P3_U4080 & new_P3_U7217;
  assign new_P3_U4080 = new_P3_U7220 & new_P3_U7219;
  assign new_P3_U4081 = new_P3_U7222 & new_P3_U7221 & new_P3_U4316;
  assign new_P3_U4082 = new_P3_U4083 & new_P3_U7225;
  assign new_P3_U4083 = new_P3_U7228 & new_P3_U7227;
  assign new_P3_U4084 = new_P3_U7230 & new_P3_U7229 & new_P3_U4316;
  assign new_P3_U4085 = new_P3_U4086 & new_P3_U7233;
  assign new_P3_U4086 = new_P3_U7236 & new_P3_U7235;
  assign new_P3_U4087 = new_P3_U7238 & new_P3_U7237 & new_P3_U4316;
  assign new_P3_U4088 = new_P3_U4089 & new_P3_U7241;
  assign new_P3_U4089 = new_P3_U7244 & new_P3_U7243;
  assign new_P3_U4090 = new_P3_U7246 & new_P3_U7245 & new_P3_U4316;
  assign new_P3_U4091 = new_P3_U4092 & new_P3_U7249;
  assign new_P3_U4092 = new_P3_U7252 & new_P3_U7251;
  assign new_P3_U4093 = new_P3_U7254 & new_P3_U7253 & new_P3_U4316;
  assign new_P3_U4094 = new_P3_U4095 & new_P3_U7257;
  assign new_P3_U4095 = new_P3_U7260 & new_P3_U7259;
  assign new_P3_U4096 = new_P3_U7262 & new_P3_U7261 & new_P3_U4316;
  assign new_P3_U4097 = new_P3_U4098 & new_P3_U7265;
  assign new_P3_U4098 = new_P3_U7268 & new_P3_U7267;
  assign new_P3_U4099 = new_P3_U7270 & new_P3_U7269;
  assign new_P3_U4100 = new_P3_U4101 & new_P3_U7273;
  assign new_P3_U4101 = new_P3_U7276 & new_P3_U7275;
  assign new_P3_U4102 = new_P3_U7278 & new_P3_U7277;
  assign new_P3_U4103 = new_P3_U4104 & new_P3_U7281;
  assign new_P3_U4104 = new_P3_U7284 & new_P3_U7283;
  assign new_P3_U4105 = new_P3_U7286 & new_P3_U7285;
  assign new_P3_U4106 = new_P3_U4107 & new_P3_U7289;
  assign new_P3_U4107 = new_P3_U7292 & new_P3_U7291;
  assign new_P3_U4108 = new_P3_U7294 & new_P3_U7293;
  assign new_P3_U4109 = new_P3_U4110 & new_P3_U7297;
  assign new_P3_U4110 = new_P3_U7300 & new_P3_U7299;
  assign new_P3_U4111 = new_P3_U7302 & new_P3_U7301;
  assign new_P3_U4112 = new_P3_U4113 & new_P3_U7305;
  assign new_P3_U4113 = new_P3_U7308 & new_P3_U7307;
  assign new_P3_U4114 = new_P3_U7310 & new_P3_U7309;
  assign new_P3_U4115 = new_P3_U4116 & new_P3_U7313;
  assign new_P3_U4116 = new_P3_U7316 & new_P3_U7315;
  assign new_P3_U4117 = new_P3_U7318 & new_P3_U7317;
  assign new_P3_U4118 = new_P3_U4119 & new_P3_U7321;
  assign new_P3_U4119 = new_P3_U7324 & new_P3_U7323;
  assign new_P3_U4120 = new_P3_U7326 & new_P3_U7325;
  assign new_P3_U4121 = new_P3_U4122 & new_P3_U7329;
  assign new_P3_U4122 = new_P3_U7332 & new_P3_U7331;
  assign new_P3_U4123 = new_P3_U7334 & new_P3_U7333;
  assign new_P3_U4124 = new_P3_U4125 & new_P3_U7337;
  assign new_P3_U4125 = new_P3_U7340 & new_P3_U7339;
  assign new_P3_U4126 = new_P3_U7342 & new_P3_U7341;
  assign new_P3_U4127 = new_P3_U4128 & new_P3_U7345;
  assign new_P3_U4128 = new_P3_U7348 & new_P3_U7347;
  assign new_P3_U4129 = new_P3_U7350 & new_P3_U7349;
  assign new_P3_U4130 = new_P3_U4131 & new_P3_U7353;
  assign new_P3_U4131 = new_P3_U7356 & new_P3_U7355;
  assign new_P3_U4132 = new_P3_U7364 & new_P3_U7365;
  assign new_P3_U4133 = new_P3_U4132 & new_P3_U7361;
  assign new_P3_U4134 = new_P3_U7362 & new_P3_U3259;
  assign new_P3_U4135 = ~new_P3_SUB_320_U51 & ~new_P3_U7363;
  assign new_P3_U4136 = ~P3_DATAWIDTH_REG_5_ & ~P3_DATAWIDTH_REG_4_ & ~P3_DATAWIDTH_REG_2_ & ~P3_DATAWIDTH_REG_3_;
  assign new_P3_U4137 = ~P3_DATAWIDTH_REG_9_ & ~P3_DATAWIDTH_REG_8_ & ~P3_DATAWIDTH_REG_6_ & ~P3_DATAWIDTH_REG_7_;
  assign new_P3_U4138 = new_P3_U4137 & new_P3_U4136;
  assign new_P3_U4139 = ~P3_DATAWIDTH_REG_13_ & ~P3_DATAWIDTH_REG_12_ & ~P3_DATAWIDTH_REG_10_ & ~P3_DATAWIDTH_REG_11_;
  assign new_P3_U4140 = ~P3_DATAWIDTH_REG_17_ & ~P3_DATAWIDTH_REG_16_ & ~P3_DATAWIDTH_REG_14_ & ~P3_DATAWIDTH_REG_15_;
  assign new_P3_U4141 = new_P3_U4140 & new_P3_U4139;
  assign new_P3_U4142 = ~P3_DATAWIDTH_REG_21_ & ~P3_DATAWIDTH_REG_20_ & ~P3_DATAWIDTH_REG_18_ & ~P3_DATAWIDTH_REG_19_;
  assign new_P3_U4143 = ~P3_DATAWIDTH_REG_25_ & ~P3_DATAWIDTH_REG_24_ & ~P3_DATAWIDTH_REG_22_ & ~P3_DATAWIDTH_REG_23_;
  assign new_P3_U4144 = new_P3_U4143 & new_P3_U4142;
  assign new_P3_U4145 = ~P3_DATAWIDTH_REG_26_ & ~P3_DATAWIDTH_REG_27_;
  assign new_P3_U4146 = ~P3_DATAWIDTH_REG_28_ & ~P3_DATAWIDTH_REG_29_;
  assign new_P3_U4147 = ~P3_DATAWIDTH_REG_30_ & ~P3_DATAWIDTH_REG_31_;
  assign new_P3_U4148 = new_P3_U4145 & new_P3_U4146 & new_P3_U4147 & new_P3_U7366;
  assign new_P3_U4149 = ~P3_DATAWIDTH_REG_1_ & ~P3_REIP_REG_0_ & ~P3_DATAWIDTH_REG_0_;
  assign new_P3_U4150 = new_P3_U7375 & new_P3_U2630;
  assign new_P3_U4151 = new_P3_U7373 & new_P3_U3135;
  assign new_P3_U4152 = new_P3_U7387 & new_P3_U7388 & new_P3_U7390 & new_P3_U7389;
  assign new_P3_U4153 = new_P3_U7391 & new_P3_U7392 & new_P3_U7394 & new_P3_U7393;
  assign new_P3_U4154 = new_P3_U7395 & new_P3_U7396 & new_P3_U7398 & new_P3_U7397;
  assign new_P3_U4155 = new_P3_U7399 & new_P3_U7400 & new_P3_U7402 & new_P3_U7401;
  assign new_P3_U4156 = new_P3_U7403 & new_P3_U7404 & new_P3_U7406 & new_P3_U7405;
  assign new_P3_U4157 = new_P3_U7407 & new_P3_U7408 & new_P3_U7410 & new_P3_U7409;
  assign new_P3_U4158 = new_P3_U7411 & new_P3_U7412 & new_P3_U7414 & new_P3_U7413;
  assign new_P3_U4159 = new_P3_U7415 & new_P3_U7416 & new_P3_U7418 & new_P3_U7417;
  assign new_P3_U4160 = new_P3_U7419 & new_P3_U7420 & new_P3_U7422 & new_P3_U7421;
  assign new_P3_U4161 = new_P3_U7423 & new_P3_U7424 & new_P3_U7426 & new_P3_U7425;
  assign new_P3_U4162 = new_P3_U7427 & new_P3_U7428 & new_P3_U7430 & new_P3_U7429;
  assign new_P3_U4163 = new_P3_U7431 & new_P3_U7432 & new_P3_U7434 & new_P3_U7433;
  assign new_P3_U4164 = new_P3_U7435 & new_P3_U7436 & new_P3_U7438 & new_P3_U7437;
  assign new_P3_U4165 = new_P3_U7439 & new_P3_U7440 & new_P3_U7442 & new_P3_U7441;
  assign new_P3_U4166 = new_P3_U7443 & new_P3_U7444 & new_P3_U7446 & new_P3_U7445;
  assign new_P3_U4167 = new_P3_U7447 & new_P3_U7448 & new_P3_U7450 & new_P3_U7449;
  assign new_P3_U4168 = new_P3_U7451 & new_P3_U7452 & new_P3_U7454 & new_P3_U7453;
  assign new_P3_U4169 = new_P3_U7455 & new_P3_U7456 & new_P3_U7458 & new_P3_U7457;
  assign new_P3_U4170 = new_P3_U7459 & new_P3_U7460 & new_P3_U7462 & new_P3_U7461;
  assign new_P3_U4171 = new_P3_U7463 & new_P3_U7464 & new_P3_U7466 & new_P3_U7465;
  assign new_P3_U4172 = new_P3_U7467 & new_P3_U7468 & new_P3_U7470 & new_P3_U7469;
  assign new_P3_U4173 = new_P3_U7471 & new_P3_U7472 & new_P3_U7474 & new_P3_U7473;
  assign new_P3_U4174 = new_P3_U7475 & new_P3_U7476 & new_P3_U7478 & new_P3_U7477;
  assign new_P3_U4175 = new_P3_U7479 & new_P3_U7480 & new_P3_U7482 & new_P3_U7481;
  assign new_P3_U4176 = new_P3_U7483 & new_P3_U7484 & new_P3_U7486 & new_P3_U7485;
  assign new_P3_U4177 = new_P3_U7487 & new_P3_U7488 & new_P3_U7490 & new_P3_U7489;
  assign new_P3_U4178 = new_P3_U7491 & new_P3_U7492 & new_P3_U7494 & new_P3_U7493;
  assign new_P3_U4179 = new_P3_U7495 & new_P3_U7496 & new_P3_U7498 & new_P3_U7497;
  assign new_P3_U4180 = new_P3_U7499 & new_P3_U7500 & new_P3_U7502 & new_P3_U7501;
  assign new_P3_U4181 = new_P3_U7503 & new_P3_U7504 & new_P3_U7506 & new_P3_U7505;
  assign new_P3_U4182 = new_P3_U7507 & new_P3_U7508 & new_P3_U7510 & new_P3_U7509;
  assign new_P3_U4183 = new_P3_U7511 & new_P3_U7512 & new_P3_U7514 & new_P3_U7513;
  assign new_P3_U4184 = new_P3_U7517 & new_P3_U7518 & new_P3_U7520 & new_P3_U7519;
  assign new_P3_U4185 = new_P3_U7521 & new_P3_U7522 & new_P3_U7524 & new_P3_U7523;
  assign new_P3_U4186 = new_P3_U7525 & new_P3_U7526 & new_P3_U7528 & new_P3_U7527;
  assign new_P3_U4187 = new_P3_U7529 & new_P3_U7530 & new_P3_U7532 & new_P3_U7531;
  assign new_P3_U4188 = new_P3_U7533 & new_P3_U7534 & new_P3_U7536 & new_P3_U7535;
  assign new_P3_U4189 = new_P3_U7537 & new_P3_U7538 & new_P3_U7540 & new_P3_U7539;
  assign new_P3_U4190 = new_P3_U7541 & new_P3_U7542 & new_P3_U7544 & new_P3_U7543;
  assign new_P3_U4191 = new_P3_U7545 & new_P3_U7546 & new_P3_U7548 & new_P3_U7547;
  assign new_P3_U4192 = new_P3_U7549 & new_P3_U7550 & new_P3_U7552 & new_P3_U7551;
  assign new_P3_U4193 = new_P3_U7553 & new_P3_U7554 & new_P3_U7556 & new_P3_U7555;
  assign new_P3_U4194 = new_P3_U7557 & new_P3_U7558 & new_P3_U7560 & new_P3_U7559;
  assign new_P3_U4195 = new_P3_U7561 & new_P3_U7562 & new_P3_U7564 & new_P3_U7563;
  assign new_P3_U4196 = new_P3_U7565 & new_P3_U7566 & new_P3_U7568 & new_P3_U7567;
  assign new_P3_U4197 = new_P3_U7569 & new_P3_U7570 & new_P3_U7572 & new_P3_U7571;
  assign new_P3_U4198 = new_P3_U7573 & new_P3_U7574 & new_P3_U7576 & new_P3_U7575;
  assign new_P3_U4199 = new_P3_U7577 & new_P3_U7578 & new_P3_U7580 & new_P3_U7579;
  assign new_P3_U4200 = new_P3_U7581 & new_P3_U7582 & new_P3_U7584 & new_P3_U7583;
  assign new_P3_U4201 = new_P3_U7585 & new_P3_U7586 & new_P3_U7588 & new_P3_U7587;
  assign new_P3_U4202 = new_P3_U7589 & new_P3_U7590 & new_P3_U7592 & new_P3_U7591;
  assign new_P3_U4203 = new_P3_U7593 & new_P3_U7594 & new_P3_U7596 & new_P3_U7595;
  assign new_P3_U4204 = new_P3_U7597 & new_P3_U7598 & new_P3_U7600 & new_P3_U7599;
  assign new_P3_U4205 = new_P3_U7601 & new_P3_U7602 & new_P3_U7604 & new_P3_U7603;
  assign new_P3_U4206 = new_P3_U7605 & new_P3_U7606 & new_P3_U7608 & new_P3_U7607;
  assign new_P3_U4207 = new_P3_U7609 & new_P3_U7610 & new_P3_U7612 & new_P3_U7611;
  assign new_P3_U4208 = new_P3_U7613 & new_P3_U7614 & new_P3_U7616 & new_P3_U7615;
  assign new_P3_U4209 = new_P3_U7617 & new_P3_U7618 & new_P3_U7620 & new_P3_U7619;
  assign new_P3_U4210 = new_P3_U7621 & new_P3_U7622 & new_P3_U7624 & new_P3_U7623;
  assign new_P3_U4211 = new_P3_U7625 & new_P3_U7626 & new_P3_U7628 & new_P3_U7627;
  assign new_P3_U4212 = new_P3_U7629 & new_P3_U7630 & new_P3_U7632 & new_P3_U7631;
  assign new_P3_U4213 = new_P3_U7633 & new_P3_U7634 & new_P3_U7636 & new_P3_U7635;
  assign new_P3_U4214 = new_P3_U7637 & new_P3_U7638 & new_P3_U7640 & new_P3_U7639;
  assign new_P3_U4215 = new_P3_U7641 & new_P3_U7642 & new_P3_U7644 & new_P3_U7643;
  assign new_P3_U4216 = new_P3_U7646 & new_P3_U7647 & new_P3_U7649 & new_P3_U7648;
  assign new_P3_U4217 = new_P3_U7650 & new_P3_U7651 & new_P3_U7653 & new_P3_U7652;
  assign new_P3_U4218 = new_P3_U7654 & new_P3_U7655 & new_P3_U7657 & new_P3_U7656;
  assign new_P3_U4219 = new_P3_U7658 & new_P3_U7659 & new_P3_U7661 & new_P3_U7660;
  assign new_P3_U4220 = new_P3_U7662 & new_P3_U7663 & new_P3_U7665 & new_P3_U7664;
  assign new_P3_U4221 = new_P3_U7666 & new_P3_U7667 & new_P3_U7669 & new_P3_U7668;
  assign new_P3_U4222 = new_P3_U7670 & new_P3_U7671 & new_P3_U7673 & new_P3_U7672;
  assign new_P3_U4223 = new_P3_U7674 & new_P3_U7675 & new_P3_U7677 & new_P3_U7676;
  assign new_P3_U4224 = new_P3_U7678 & new_P3_U7679 & new_P3_U7681 & new_P3_U7680;
  assign new_P3_U4225 = new_P3_U7682 & new_P3_U7683 & new_P3_U7685 & new_P3_U7684;
  assign new_P3_U4226 = new_P3_U7686 & new_P3_U7687 & new_P3_U7689 & new_P3_U7688;
  assign new_P3_U4227 = new_P3_U7690 & new_P3_U7691 & new_P3_U7693 & new_P3_U7692;
  assign new_P3_U4228 = new_P3_U7694 & new_P3_U7695 & new_P3_U7697 & new_P3_U7696;
  assign new_P3_U4229 = new_P3_U7698 & new_P3_U7699 & new_P3_U7701 & new_P3_U7700;
  assign new_P3_U4230 = new_P3_U7702 & new_P3_U7703 & new_P3_U7705 & new_P3_U7704;
  assign new_P3_U4231 = new_P3_U7706 & new_P3_U7707 & new_P3_U7709 & new_P3_U7708;
  assign new_P3_U4232 = new_P3_U7710 & new_P3_U7711 & new_P3_U7713 & new_P3_U7712;
  assign new_P3_U4233 = new_P3_U7714 & new_P3_U7715 & new_P3_U7717 & new_P3_U7716;
  assign new_P3_U4234 = new_P3_U7718 & new_P3_U7719 & new_P3_U7721 & new_P3_U7720;
  assign new_P3_U4235 = new_P3_U7722 & new_P3_U7723 & new_P3_U7725 & new_P3_U7724;
  assign new_P3_U4236 = new_P3_U7726 & new_P3_U7727 & new_P3_U7729 & new_P3_U7728;
  assign new_P3_U4237 = new_P3_U7730 & new_P3_U7731 & new_P3_U7733 & new_P3_U7732;
  assign new_P3_U4238 = new_P3_U7734 & new_P3_U7735 & new_P3_U7737 & new_P3_U7736;
  assign new_P3_U4239 = new_P3_U7738 & new_P3_U7739 & new_P3_U7741 & new_P3_U7740;
  assign new_P3_U4240 = new_P3_U7742 & new_P3_U7743 & new_P3_U7745 & new_P3_U7744;
  assign new_P3_U4241 = new_P3_U7746 & new_P3_U7747 & new_P3_U7749 & new_P3_U7748;
  assign new_P3_U4242 = new_P3_U7750 & new_P3_U7751 & new_P3_U7753 & new_P3_U7752;
  assign new_P3_U4243 = new_P3_U7754 & new_P3_U7755 & new_P3_U7757 & new_P3_U7756;
  assign new_P3_U4244 = new_P3_U7758 & new_P3_U7759 & new_P3_U7761 & new_P3_U7760;
  assign new_P3_U4245 = new_P3_U7762 & new_P3_U7763 & new_P3_U7765 & new_P3_U7764;
  assign new_P3_U4246 = new_P3_U7766 & new_P3_U7767 & new_P3_U7769 & new_P3_U7768;
  assign new_P3_U4247 = new_P3_U7770 & new_P3_U7771 & new_P3_U7773 & new_P3_U7772;
  assign new_P3_U4248 = new_P3_U7776 & new_P3_U7777 & new_P3_U7779 & new_P3_U7778;
  assign new_P3_U4249 = new_P3_U7780 & new_P3_U7781 & new_P3_U7783 & new_P3_U7782;
  assign new_P3_U4250 = new_P3_U7784 & new_P3_U7785 & new_P3_U7787 & new_P3_U7786;
  assign new_P3_U4251 = new_P3_U7788 & new_P3_U7789 & new_P3_U7791 & new_P3_U7790;
  assign new_P3_U4252 = new_P3_U7792 & new_P3_U7793 & new_P3_U7795 & new_P3_U7794;
  assign new_P3_U4253 = new_P3_U7796 & new_P3_U7797 & new_P3_U7799 & new_P3_U7798;
  assign new_P3_U4254 = new_P3_U7800 & new_P3_U7801 & new_P3_U7803 & new_P3_U7802;
  assign new_P3_U4255 = new_P3_U7804 & new_P3_U7805 & new_P3_U7807 & new_P3_U7806;
  assign new_P3_U4256 = new_P3_U7808 & new_P3_U7809 & new_P3_U7811 & new_P3_U7810;
  assign new_P3_U4257 = new_P3_U7812 & new_P3_U7813 & new_P3_U7815 & new_P3_U7814;
  assign new_P3_U4258 = new_P3_U7816 & new_P3_U7817 & new_P3_U7819 & new_P3_U7818;
  assign new_P3_U4259 = new_P3_U7820 & new_P3_U7821 & new_P3_U7823 & new_P3_U7822;
  assign new_P3_U4260 = new_P3_U7824 & new_P3_U7825 & new_P3_U7827 & new_P3_U7826;
  assign new_P3_U4261 = new_P3_U7828 & new_P3_U7829 & new_P3_U7831 & new_P3_U7830;
  assign new_P3_U4262 = new_P3_U7832 & new_P3_U7833 & new_P3_U7835 & new_P3_U7834;
  assign new_P3_U4263 = new_P3_U7836 & new_P3_U7837 & new_P3_U7839 & new_P3_U7838;
  assign new_P3_U4264 = new_P3_U7840 & new_P3_U7841 & new_P3_U7843 & new_P3_U7842;
  assign new_P3_U4265 = new_P3_U7844 & new_P3_U7845 & new_P3_U7847 & new_P3_U7846;
  assign new_P3_U4266 = new_P3_U7848 & new_P3_U7849 & new_P3_U7851 & new_P3_U7850;
  assign new_P3_U4267 = new_P3_U7852 & new_P3_U7853 & new_P3_U7855 & new_P3_U7854;
  assign new_P3_U4268 = new_P3_U7856 & new_P3_U7857 & new_P3_U7859 & new_P3_U7858;
  assign new_P3_U4269 = new_P3_U7860 & new_P3_U7861 & new_P3_U7863 & new_P3_U7862;
  assign new_P3_U4270 = new_P3_U7864 & new_P3_U7865 & new_P3_U7867 & new_P3_U7866;
  assign new_P3_U4271 = new_P3_U7868 & new_P3_U7869 & new_P3_U7871 & new_P3_U7870;
  assign new_P3_U4272 = new_P3_U7872 & new_P3_U7873 & new_P3_U7875 & new_P3_U7874;
  assign new_P3_U4273 = new_P3_U7876 & new_P3_U7877 & new_P3_U7879 & new_P3_U7878;
  assign new_P3_U4274 = new_P3_U7880 & new_P3_U7881 & new_P3_U7883 & new_P3_U7882;
  assign new_P3_U4275 = new_P3_U7884 & new_P3_U7885 & new_P3_U7887 & new_P3_U7886;
  assign new_P3_U4276 = new_P3_U7888 & new_P3_U7889 & new_P3_U7891 & new_P3_U7890;
  assign new_P3_U4277 = new_P3_U7892 & new_P3_U7893 & new_P3_U7895 & new_P3_U7894;
  assign new_P3_U4278 = new_P3_U7896 & new_P3_U7897 & new_P3_U7899 & new_P3_U7898;
  assign new_P3_U4279 = new_P3_U7900 & new_P3_U7901 & new_P3_U7903 & new_P3_U7902;
  assign new_P3_U4280 = new_P3_U7943 & new_P3_U7942;
  assign new_P3_U4281 = ~new_P3_U3361 | ~new_P3_U2604;
  assign new_P3_U4282 = new_P3_U7951 & new_P3_U7950;
  assign new_P3_U4283 = ~new_P3_U3658 | ~new_P3_U5497;
  assign new_P3_U4284 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_U4285 = ~new_P3_U2390 | ~new_P3_U4281;
  assign new_P3_U4286 = ~BS16;
  assign new_P3_U4287 = ~new_P3_U4151 | ~new_P3_U4334;
  assign new_P3_U4288 = ~new_P3_U4334 | ~new_P3_U3239;
  assign new_P3_U4289 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U3091;
  assign new_P3_U4290 = ~new_P3_U3657 | ~new_P3_U2515 | ~new_P3_U2516;
  assign new_P3_U4291 = ~new_P3_U3267;
  assign new_P3_U4292 = ~HOLD | ~new_P3_U2630;
  assign new_P3_U4293 = ~new_P3_U3105;
  assign new_P3_U4294 = ~new_P3_U3106;
  assign new_P3_U4295 = ~new_P3_U3135;
  assign new_P3_U4296 = ~new_P3_U3112;
  assign new_P3_U4297 = ~new_P3_U3111;
  assign new_P3_U4298 = ~new_P3_U3242;
  assign new_P3_U4299 = ~new_P3_U3243;
  assign new_P3_U4300 = ~new_P3_U3244;
  assign new_P3_U4301 = ~new_P3_U3245;
  assign new_P3_U4302 = ~new_P3_U3119;
  assign new_P3_U4303 = ~new_P3_U3117;
  assign new_P3_U4304 = ~new_P3_U3116;
  assign new_P3_U4305 = ~new_P3_U3115;
  assign new_P3_U4306 = ~new_P3_U3246;
  assign new_P3_U4307 = ~new_P3_U3261;
  assign new_P3_U4308 = ~new_P3_U3077;
  assign new_P3_U4309 = ~new_P3_U3253;
  assign new_P3_U4310 = ~new_P3_U3252;
  assign new_P3_U4311 = ~new_P3_U3250;
  assign new_P3_U4312 = ~new_P3_U3127;
  assign new_P3_U4313 = ~new_P3_LT_563_1260_U6;
  assign new_P3_U4314 = ~new_P3_U3217;
  assign new_P3_U4315 = ~new_P3_U4295 | ~new_P3_U2631;
  assign new_P3_U4316 = ~new_P3_U4347 | ~new_P3_U3260;
  assign new_P3_U4317 = ~new_P3_U2383 | ~new_P3_U3105;
  assign new_P3_U4318 = ~new_P3_U3247;
  assign new_P3_U4319 = ~new_P3_U3259;
  assign new_P3_U4320 = ~new_P3_U3080;
  assign new_P3_U4321 = ~new_P3_U3078;
  assign new_P3_U4322 = ~new_P3_U3136;
  assign new_P3_U4323 = ~new_P3_U3114;
  assign new_P3_U4324 = ~new_P3_U3118;
  assign new_P3_U4325 = ~new_P3_U3219;
  assign new_P3_U4326 = ~new_P3_U3181;
  assign new_P3_U4327 = ~new_P3_U4149 | ~new_P3_U4307;
  assign new_P3_U4328 = ~new_P3_U3365 | ~new_P3_U4354;
  assign new_P3_U4329 = ~new_P3_U2631 | ~new_P3_U3090 | ~P3_STATE2_REG_1_ | ~new_P3_U3121;
  assign new_P3_U4330 = ~new_P3_U3653 | ~new_P3_U2453;
  assign new_P3_U4331 = ~new_P3_U2458 | ~new_P3_U4653;
  assign new_P3_U4332 = ~new_P3_U3095;
  assign new_P3_U4333 = ~new_P3_U4350 | ~new_P3_U3113;
  assign new_P3_U4334 = ~new_P3_U2390 | ~new_P3_U7093;
  assign new_P3_U4335 = ~new_P3_U4452 | ~new_P3_U3085;
  assign new_P3_U4336 = ~new_P3_U4347 | ~new_P3_U3121;
  assign new_P3_U4337 = ~new_P3_U2453 | ~new_P3_U3232;
  assign new_P3_U4338 = ~new_U209 | ~new_P3_U3090 | ~P3_STATE2_REG_0_;
  assign new_P3_U4339 = ~new_P3_U3654 | ~new_P3_U4608;
  assign new_P3_U4340 = ~new_P3_U3123;
  assign new_P3_U4341 = ~new_P3_U3229;
  assign new_P3_U4342 = ~new_P3_U3150;
  assign new_P3_U4343 = ~new_P3_U3158;
  assign new_P3_U4344 = ~new_P3_U3103;
  assign new_P3_U4345 = ~new_P3_U3126;
  assign new_P3_U4346 = ~new_P3_U3082;
  assign new_P3_U4347 = ~new_P3_U3239;
  assign new_P3_U4348 = ~new_P3_U3236;
  assign new_P3_U4349 = ~new_P3_U3235;
  assign new_P3_U4350 = ~new_P3_U3208;
  assign new_P3_U4351 = ~new_P3_U3216;
  assign new_P3_U4352 = ~new_P3_U3222;
  assign new_P3_U4353 = ~new_P3_U3124;
  assign new_P3_U4354 = ~new_P3_U3125;
  assign new_P3_U4355 = ~P3_REIP_REG_31_ | ~new_P3_U4321;
  assign new_P3_U4356 = ~P3_REIP_REG_30_ | ~new_P3_U4320;
  assign new_P3_U4357 = ~P3_ADDRESS_REG_29_ | ~new_P3_U3077;
  assign new_P3_U4358 = ~P3_REIP_REG_30_ | ~new_P3_U4321;
  assign new_P3_U4359 = ~P3_REIP_REG_29_ | ~new_P3_U4320;
  assign new_P3_U4360 = ~P3_ADDRESS_REG_28_ | ~new_P3_U3077;
  assign new_P3_U4361 = ~P3_REIP_REG_29_ | ~new_P3_U4321;
  assign new_P3_U4362 = ~P3_REIP_REG_28_ | ~new_P3_U4320;
  assign new_P3_U4363 = ~P3_ADDRESS_REG_27_ | ~new_P3_U3077;
  assign new_P3_U4364 = ~P3_REIP_REG_28_ | ~new_P3_U4321;
  assign new_P3_U4365 = ~P3_REIP_REG_27_ | ~new_P3_U4320;
  assign new_P3_U4366 = ~P3_ADDRESS_REG_26_ | ~new_P3_U3077;
  assign new_P3_U4367 = ~P3_REIP_REG_27_ | ~new_P3_U4321;
  assign new_P3_U4368 = ~P3_REIP_REG_26_ | ~new_P3_U4320;
  assign new_P3_U4369 = ~P3_ADDRESS_REG_25_ | ~new_P3_U3077;
  assign new_P3_U4370 = ~P3_REIP_REG_26_ | ~new_P3_U4321;
  assign new_P3_U4371 = ~P3_REIP_REG_25_ | ~new_P3_U4320;
  assign new_P3_U4372 = ~P3_ADDRESS_REG_24_ | ~new_P3_U3077;
  assign new_P3_U4373 = ~P3_REIP_REG_25_ | ~new_P3_U4321;
  assign new_P3_U4374 = ~P3_REIP_REG_24_ | ~new_P3_U4320;
  assign new_P3_U4375 = ~P3_ADDRESS_REG_23_ | ~new_P3_U3077;
  assign new_P3_U4376 = ~P3_REIP_REG_24_ | ~new_P3_U4321;
  assign new_P3_U4377 = ~P3_REIP_REG_23_ | ~new_P3_U4320;
  assign new_P3_U4378 = ~P3_ADDRESS_REG_22_ | ~new_P3_U3077;
  assign new_P3_U4379 = ~P3_REIP_REG_23_ | ~new_P3_U4321;
  assign new_P3_U4380 = ~P3_REIP_REG_22_ | ~new_P3_U4320;
  assign new_P3_U4381 = ~P3_ADDRESS_REG_21_ | ~new_P3_U3077;
  assign new_P3_U4382 = ~P3_REIP_REG_22_ | ~new_P3_U4321;
  assign new_P3_U4383 = ~P3_REIP_REG_21_ | ~new_P3_U4320;
  assign new_P3_U4384 = ~P3_ADDRESS_REG_20_ | ~new_P3_U3077;
  assign new_P3_U4385 = ~P3_REIP_REG_21_ | ~new_P3_U4321;
  assign new_P3_U4386 = ~P3_REIP_REG_20_ | ~new_P3_U4320;
  assign new_P3_U4387 = ~P3_ADDRESS_REG_19_ | ~new_P3_U3077;
  assign new_P3_U4388 = ~P3_REIP_REG_20_ | ~new_P3_U4321;
  assign new_P3_U4389 = ~P3_REIP_REG_19_ | ~new_P3_U4320;
  assign new_P3_U4390 = ~P3_ADDRESS_REG_18_ | ~new_P3_U3077;
  assign new_P3_U4391 = ~P3_REIP_REG_19_ | ~new_P3_U4321;
  assign new_P3_U4392 = ~P3_REIP_REG_18_ | ~new_P3_U4320;
  assign new_P3_U4393 = ~P3_ADDRESS_REG_17_ | ~new_P3_U3077;
  assign new_P3_U4394 = ~P3_REIP_REG_18_ | ~new_P3_U4321;
  assign new_P3_U4395 = ~P3_REIP_REG_17_ | ~new_P3_U4320;
  assign new_P3_U4396 = ~P3_ADDRESS_REG_16_ | ~new_P3_U3077;
  assign new_P3_U4397 = ~P3_REIP_REG_17_ | ~new_P3_U4321;
  assign new_P3_U4398 = ~P3_REIP_REG_16_ | ~new_P3_U4320;
  assign new_P3_U4399 = ~P3_ADDRESS_REG_15_ | ~new_P3_U3077;
  assign new_P3_U4400 = ~P3_REIP_REG_16_ | ~new_P3_U4321;
  assign new_P3_U4401 = ~P3_REIP_REG_15_ | ~new_P3_U4320;
  assign new_P3_U4402 = ~P3_ADDRESS_REG_14_ | ~new_P3_U3077;
  assign new_P3_U4403 = ~P3_REIP_REG_15_ | ~new_P3_U4321;
  assign new_P3_U4404 = ~P3_REIP_REG_14_ | ~new_P3_U4320;
  assign new_P3_U4405 = ~P3_ADDRESS_REG_13_ | ~new_P3_U3077;
  assign new_P3_U4406 = ~P3_REIP_REG_14_ | ~new_P3_U4321;
  assign new_P3_U4407 = ~P3_REIP_REG_13_ | ~new_P3_U4320;
  assign new_P3_U4408 = ~P3_ADDRESS_REG_12_ | ~new_P3_U3077;
  assign new_P3_U4409 = ~P3_REIP_REG_13_ | ~new_P3_U4321;
  assign new_P3_U4410 = ~P3_REIP_REG_12_ | ~new_P3_U4320;
  assign new_P3_U4411 = ~P3_ADDRESS_REG_11_ | ~new_P3_U3077;
  assign new_P3_U4412 = ~P3_REIP_REG_12_ | ~new_P3_U4321;
  assign new_P3_U4413 = ~P3_REIP_REG_11_ | ~new_P3_U4320;
  assign new_P3_U4414 = ~P3_ADDRESS_REG_10_ | ~new_P3_U3077;
  assign new_P3_U4415 = ~P3_REIP_REG_11_ | ~new_P3_U4321;
  assign new_P3_U4416 = ~P3_REIP_REG_10_ | ~new_P3_U4320;
  assign new_P3_U4417 = ~P3_ADDRESS_REG_9_ | ~new_P3_U3077;
  assign new_P3_U4418 = ~P3_REIP_REG_10_ | ~new_P3_U4321;
  assign new_P3_U4419 = ~P3_REIP_REG_9_ | ~new_P3_U4320;
  assign new_P3_U4420 = ~P3_ADDRESS_REG_8_ | ~new_P3_U3077;
  assign new_P3_U4421 = ~P3_REIP_REG_9_ | ~new_P3_U4321;
  assign new_P3_U4422 = ~P3_REIP_REG_8_ | ~new_P3_U4320;
  assign new_P3_U4423 = ~P3_ADDRESS_REG_7_ | ~new_P3_U3077;
  assign new_P3_U4424 = ~P3_REIP_REG_8_ | ~new_P3_U4321;
  assign new_P3_U4425 = ~P3_REIP_REG_7_ | ~new_P3_U4320;
  assign new_P3_U4426 = ~P3_ADDRESS_REG_6_ | ~new_P3_U3077;
  assign new_P3_U4427 = ~P3_REIP_REG_7_ | ~new_P3_U4321;
  assign new_P3_U4428 = ~P3_REIP_REG_6_ | ~new_P3_U4320;
  assign new_P3_U4429 = ~P3_ADDRESS_REG_5_ | ~new_P3_U3077;
  assign new_P3_U4430 = ~P3_REIP_REG_6_ | ~new_P3_U4321;
  assign new_P3_U4431 = ~P3_REIP_REG_5_ | ~new_P3_U4320;
  assign new_P3_U4432 = ~P3_ADDRESS_REG_4_ | ~new_P3_U3077;
  assign new_P3_U4433 = ~P3_REIP_REG_5_ | ~new_P3_U4321;
  assign new_P3_U4434 = ~P3_REIP_REG_4_ | ~new_P3_U4320;
  assign new_P3_U4435 = ~P3_ADDRESS_REG_3_ | ~new_P3_U3077;
  assign new_P3_U4436 = ~P3_REIP_REG_4_ | ~new_P3_U4321;
  assign new_P3_U4437 = ~P3_REIP_REG_3_ | ~new_P3_U4320;
  assign new_P3_U4438 = ~P3_ADDRESS_REG_2_ | ~new_P3_U3077;
  assign new_P3_U4439 = ~P3_REIP_REG_3_ | ~new_P3_U4321;
  assign new_P3_U4440 = ~P3_REIP_REG_2_ | ~new_P3_U4320;
  assign new_P3_U4441 = ~P3_ADDRESS_REG_1_ | ~new_P3_U3077;
  assign new_P3_U4442 = ~P3_REIP_REG_2_ | ~new_P3_U4321;
  assign new_P3_U4443 = ~P3_REIP_REG_1_ | ~new_P3_U4320;
  assign new_P3_U4444 = ~P3_ADDRESS_REG_0_ | ~new_P3_U3077;
  assign new_P3_U4445 = ~new_P3_U3087;
  assign new_P3_U4446 = ~new_P3_U4445 | ~new_P3_U2630;
  assign new_P3_U4447 = ~NA | ~new_P3_U4346;
  assign new_P3_U4448 = ~new_P3_U3088;
  assign new_P3_U4449 = ~new_P3_U4448 | ~new_P3_U2630;
  assign new_P3_U4450 = P3_STATE_REG_0_ | NA;
  assign new_P3_U4451 = ~new_P3_U7913 | ~new_P3_U7912 | ~new_P3_U4450;
  assign new_P3_U4452 = ~new_P3_U3083;
  assign new_P3_U4453 = ~new_P3_U4346 | ~new_P3_U3088 | ~new_U209;
  assign new_P3_U4454 = ~new_P3_U4452 | ~HOLD | ~new_P3_U3075;
  assign new_P3_U4455 = ~new_P3_U4453 | ~new_P3_U4454;
  assign new_P3_U4456 = ~new_P3_U3309 | ~new_P3_U4455;
  assign new_P3_U4457 = ~P3_STATE_REG_2_ | ~new_P3_U4451;
  assign new_P3_U4458 = ~new_P3_U4308 | ~new_U209;
  assign new_P3_U4459 = ~new_P3_U3312 | ~new_P3_U7915;
  assign new_P3_U4460 = ~P3_STATE_REG_2_ | ~new_P3_U3087;
  assign new_P3_U4461 = ~NA | ~new_P3_U3085;
  assign new_P3_U4462 = ~new_P3_U4461 | ~new_P3_U4460;
  assign new_P3_U4463 = ~new_P3_U4462 | ~new_P3_U3076;
  assign new_P3_U4464 = ~new_P3_U4286 | ~new_P3_U3083;
  assign new_P3_U4465 = ~P3_STATE_REG_2_ | ~new_P3_U3076;
  assign new_P3_U4466 = ~new_P3_U3082 | ~new_P3_U4465;
  assign new_P3_U4467 = ~new_P3_U3091;
  assign new_P3_U4468 = ~new_P3_U3096;
  assign new_P3_U4469 = ~new_P3_U3092;
  assign new_P3_U4470 = ~new_P3_U3098;
  assign new_P3_U4471 = ~new_P3_U3099;
  assign new_P3_U4472 = ~P3_INSTQUEUE_REG_0__0_ | ~new_P3_U2484;
  assign new_P3_U4473 = ~P3_INSTQUEUE_REG_1__0_ | ~new_P3_U2483;
  assign new_P3_U4474 = ~P3_INSTQUEUE_REG_2__0_ | ~new_P3_U2482;
  assign new_P3_U4475 = ~P3_INSTQUEUE_REG_3__0_ | ~new_P3_U2480;
  assign new_P3_U4476 = ~P3_INSTQUEUE_REG_4__0_ | ~new_P3_U2479;
  assign new_P3_U4477 = ~P3_INSTQUEUE_REG_5__0_ | ~new_P3_U2478;
  assign new_P3_U4478 = ~P3_INSTQUEUE_REG_6__0_ | ~new_P3_U2477;
  assign new_P3_U4479 = ~P3_INSTQUEUE_REG_7__0_ | ~new_P3_U4471;
  assign new_P3_U4480 = ~P3_INSTQUEUE_REG_8__0_ | ~new_P3_U2476;
  assign new_P3_U4481 = ~P3_INSTQUEUE_REG_9__0_ | ~new_P3_U2475;
  assign new_P3_U4482 = ~P3_INSTQUEUE_REG_10__0_ | ~new_P3_U2473;
  assign new_P3_U4483 = ~P3_INSTQUEUE_REG_11__0_ | ~new_P3_U2471;
  assign new_P3_U4484 = ~P3_INSTQUEUE_REG_12__0_ | ~new_P3_U2470;
  assign new_P3_U4485 = ~P3_INSTQUEUE_REG_13__0_ | ~new_P3_U2469;
  assign new_P3_U4486 = ~P3_INSTQUEUE_REG_14__0_ | ~new_P3_U2467;
  assign new_P3_U4487 = ~P3_INSTQUEUE_REG_15__0_ | ~new_P3_U2465;
  assign new_P3_U4488 = ~new_P3_U3108;
  assign new_P3_U4489 = ~P3_INSTQUEUE_REG_0__1_ | ~new_P3_U2484;
  assign new_P3_U4490 = ~P3_INSTQUEUE_REG_1__1_ | ~new_P3_U2483;
  assign new_P3_U4491 = ~P3_INSTQUEUE_REG_2__1_ | ~new_P3_U2482;
  assign new_P3_U4492 = ~P3_INSTQUEUE_REG_3__1_ | ~new_P3_U2480;
  assign new_P3_U4493 = ~P3_INSTQUEUE_REG_4__1_ | ~new_P3_U2479;
  assign new_P3_U4494 = ~P3_INSTQUEUE_REG_5__1_ | ~new_P3_U2478;
  assign new_P3_U4495 = ~P3_INSTQUEUE_REG_6__1_ | ~new_P3_U2477;
  assign new_P3_U4496 = ~P3_INSTQUEUE_REG_7__1_ | ~new_P3_U4471;
  assign new_P3_U4497 = ~P3_INSTQUEUE_REG_8__1_ | ~new_P3_U2476;
  assign new_P3_U4498 = ~P3_INSTQUEUE_REG_9__1_ | ~new_P3_U2475;
  assign new_P3_U4499 = ~P3_INSTQUEUE_REG_10__1_ | ~new_P3_U2473;
  assign new_P3_U4500 = ~P3_INSTQUEUE_REG_11__1_ | ~new_P3_U2471;
  assign new_P3_U4501 = ~P3_INSTQUEUE_REG_12__1_ | ~new_P3_U2470;
  assign new_P3_U4502 = ~P3_INSTQUEUE_REG_13__1_ | ~new_P3_U2469;
  assign new_P3_U4503 = ~P3_INSTQUEUE_REG_14__1_ | ~new_P3_U2467;
  assign new_P3_U4504 = ~P3_INSTQUEUE_REG_15__1_ | ~new_P3_U2465;
  assign new_P3_U4505 = ~new_P3_U3104;
  assign new_P3_U4506 = ~P3_INSTQUEUE_REG_0__4_ | ~new_P3_U2484;
  assign new_P3_U4507 = ~P3_INSTQUEUE_REG_1__4_ | ~new_P3_U2483;
  assign new_P3_U4508 = ~P3_INSTQUEUE_REG_2__4_ | ~new_P3_U2482;
  assign new_P3_U4509 = ~P3_INSTQUEUE_REG_3__4_ | ~new_P3_U2480;
  assign new_P3_U4510 = ~P3_INSTQUEUE_REG_4__4_ | ~new_P3_U2479;
  assign new_P3_U4511 = ~P3_INSTQUEUE_REG_5__4_ | ~new_P3_U2478;
  assign new_P3_U4512 = ~P3_INSTQUEUE_REG_6__4_ | ~new_P3_U2477;
  assign new_P3_U4513 = ~P3_INSTQUEUE_REG_7__4_ | ~new_P3_U4471;
  assign new_P3_U4514 = ~P3_INSTQUEUE_REG_8__4_ | ~new_P3_U2476;
  assign new_P3_U4515 = ~P3_INSTQUEUE_REG_9__4_ | ~new_P3_U2475;
  assign new_P3_U4516 = ~P3_INSTQUEUE_REG_10__4_ | ~new_P3_U2473;
  assign new_P3_U4517 = ~P3_INSTQUEUE_REG_11__4_ | ~new_P3_U2471;
  assign new_P3_U4518 = ~P3_INSTQUEUE_REG_12__4_ | ~new_P3_U2470;
  assign new_P3_U4519 = ~P3_INSTQUEUE_REG_13__4_ | ~new_P3_U2469;
  assign new_P3_U4520 = ~P3_INSTQUEUE_REG_14__4_ | ~new_P3_U2467;
  assign new_P3_U4521 = ~P3_INSTQUEUE_REG_15__4_ | ~new_P3_U2465;
  assign new_P3_U4522 = ~new_P3_U3102;
  assign new_P3_U4523 = ~P3_INSTQUEUE_REG_0__2_ | ~new_P3_U2484;
  assign new_P3_U4524 = ~P3_INSTQUEUE_REG_1__2_ | ~new_P3_U2483;
  assign new_P3_U4525 = ~P3_INSTQUEUE_REG_2__2_ | ~new_P3_U2482;
  assign new_P3_U4526 = ~P3_INSTQUEUE_REG_3__2_ | ~new_P3_U2480;
  assign new_P3_U4527 = ~P3_INSTQUEUE_REG_4__2_ | ~new_P3_U2479;
  assign new_P3_U4528 = ~P3_INSTQUEUE_REG_5__2_ | ~new_P3_U2478;
  assign new_P3_U4529 = ~P3_INSTQUEUE_REG_6__2_ | ~new_P3_U2477;
  assign new_P3_U4530 = ~P3_INSTQUEUE_REG_7__2_ | ~new_P3_U4471;
  assign new_P3_U4531 = ~P3_INSTQUEUE_REG_8__2_ | ~new_P3_U2476;
  assign new_P3_U4532 = ~P3_INSTQUEUE_REG_9__2_ | ~new_P3_U2475;
  assign new_P3_U4533 = ~P3_INSTQUEUE_REG_10__2_ | ~new_P3_U2473;
  assign new_P3_U4534 = ~P3_INSTQUEUE_REG_11__2_ | ~new_P3_U2471;
  assign new_P3_U4535 = ~P3_INSTQUEUE_REG_12__2_ | ~new_P3_U2470;
  assign new_P3_U4536 = ~P3_INSTQUEUE_REG_13__2_ | ~new_P3_U2469;
  assign new_P3_U4537 = ~P3_INSTQUEUE_REG_14__2_ | ~new_P3_U2467;
  assign new_P3_U4538 = ~P3_INSTQUEUE_REG_15__2_ | ~new_P3_U2465;
  assign new_P3_U4539 = ~new_P3_U3101;
  assign new_P3_U4540 = ~P3_INSTQUEUE_REG_0__3_ | ~new_P3_U2484;
  assign new_P3_U4541 = ~P3_INSTQUEUE_REG_1__3_ | ~new_P3_U2483;
  assign new_P3_U4542 = ~P3_INSTQUEUE_REG_2__3_ | ~new_P3_U2482;
  assign new_P3_U4543 = ~P3_INSTQUEUE_REG_3__3_ | ~new_P3_U2480;
  assign new_P3_U4544 = ~P3_INSTQUEUE_REG_4__3_ | ~new_P3_U2479;
  assign new_P3_U4545 = ~P3_INSTQUEUE_REG_5__3_ | ~new_P3_U2478;
  assign new_P3_U4546 = ~P3_INSTQUEUE_REG_6__3_ | ~new_P3_U2477;
  assign new_P3_U4547 = ~P3_INSTQUEUE_REG_7__3_ | ~new_P3_U4471;
  assign new_P3_U4548 = ~P3_INSTQUEUE_REG_8__3_ | ~new_P3_U2476;
  assign new_P3_U4549 = ~P3_INSTQUEUE_REG_9__3_ | ~new_P3_U2475;
  assign new_P3_U4550 = ~P3_INSTQUEUE_REG_10__3_ | ~new_P3_U2473;
  assign new_P3_U4551 = ~P3_INSTQUEUE_REG_11__3_ | ~new_P3_U2471;
  assign new_P3_U4552 = ~P3_INSTQUEUE_REG_12__3_ | ~new_P3_U2470;
  assign new_P3_U4553 = ~P3_INSTQUEUE_REG_13__3_ | ~new_P3_U2469;
  assign new_P3_U4554 = ~P3_INSTQUEUE_REG_14__3_ | ~new_P3_U2467;
  assign new_P3_U4555 = ~P3_INSTQUEUE_REG_15__3_ | ~new_P3_U2465;
  assign new_P3_U4556 = ~new_P3_U3107;
  assign new_P3_U4557 = ~P3_INSTQUEUE_REG_0__7_ | ~new_P3_U2484;
  assign new_P3_U4558 = ~P3_INSTQUEUE_REG_1__7_ | ~new_P3_U2483;
  assign new_P3_U4559 = ~P3_INSTQUEUE_REG_2__7_ | ~new_P3_U2482;
  assign new_P3_U4560 = ~P3_INSTQUEUE_REG_3__7_ | ~new_P3_U2480;
  assign new_P3_U4561 = ~P3_INSTQUEUE_REG_4__7_ | ~new_P3_U2479;
  assign new_P3_U4562 = ~P3_INSTQUEUE_REG_5__7_ | ~new_P3_U2478;
  assign new_P3_U4563 = ~P3_INSTQUEUE_REG_6__7_ | ~new_P3_U2477;
  assign new_P3_U4564 = ~P3_INSTQUEUE_REG_7__7_ | ~new_P3_U4471;
  assign new_P3_U4565 = ~P3_INSTQUEUE_REG_8__7_ | ~new_P3_U2476;
  assign new_P3_U4566 = ~P3_INSTQUEUE_REG_9__7_ | ~new_P3_U2475;
  assign new_P3_U4567 = ~P3_INSTQUEUE_REG_10__7_ | ~new_P3_U2473;
  assign new_P3_U4568 = ~P3_INSTQUEUE_REG_11__7_ | ~new_P3_U2471;
  assign new_P3_U4569 = ~P3_INSTQUEUE_REG_12__7_ | ~new_P3_U2470;
  assign new_P3_U4570 = ~P3_INSTQUEUE_REG_13__7_ | ~new_P3_U2469;
  assign new_P3_U4571 = ~P3_INSTQUEUE_REG_14__7_ | ~new_P3_U2467;
  assign new_P3_U4572 = ~P3_INSTQUEUE_REG_15__7_ | ~new_P3_U2465;
  assign new_P3_U4573 = ~new_P3_U3218;
  assign new_P3_U4574 = ~P3_INSTQUEUE_REG_0__5_ | ~new_P3_U2484;
  assign new_P3_U4575 = ~P3_INSTQUEUE_REG_1__5_ | ~new_P3_U2483;
  assign new_P3_U4576 = ~P3_INSTQUEUE_REG_2__5_ | ~new_P3_U2482;
  assign new_P3_U4577 = ~P3_INSTQUEUE_REG_3__5_ | ~new_P3_U2480;
  assign new_P3_U4578 = ~P3_INSTQUEUE_REG_4__5_ | ~new_P3_U2479;
  assign new_P3_U4579 = ~P3_INSTQUEUE_REG_5__5_ | ~new_P3_U2478;
  assign new_P3_U4580 = ~P3_INSTQUEUE_REG_6__5_ | ~new_P3_U2477;
  assign new_P3_U4581 = ~P3_INSTQUEUE_REG_7__5_ | ~new_P3_U4471;
  assign new_P3_U4582 = ~P3_INSTQUEUE_REG_8__5_ | ~new_P3_U2476;
  assign new_P3_U4583 = ~P3_INSTQUEUE_REG_9__5_ | ~new_P3_U2475;
  assign new_P3_U4584 = ~P3_INSTQUEUE_REG_10__5_ | ~new_P3_U2473;
  assign new_P3_U4585 = ~P3_INSTQUEUE_REG_11__5_ | ~new_P3_U2471;
  assign new_P3_U4586 = ~P3_INSTQUEUE_REG_12__5_ | ~new_P3_U2470;
  assign new_P3_U4587 = ~P3_INSTQUEUE_REG_13__5_ | ~new_P3_U2469;
  assign new_P3_U4588 = ~P3_INSTQUEUE_REG_14__5_ | ~new_P3_U2467;
  assign new_P3_U4589 = ~P3_INSTQUEUE_REG_15__5_ | ~new_P3_U2465;
  assign new_P3_U4590 = ~new_P3_U3110;
  assign new_P3_U4591 = ~P3_INSTQUEUE_REG_0__6_ | ~new_P3_U2484;
  assign new_P3_U4592 = ~P3_INSTQUEUE_REG_1__6_ | ~new_P3_U2483;
  assign new_P3_U4593 = ~P3_INSTQUEUE_REG_2__6_ | ~new_P3_U2482;
  assign new_P3_U4594 = ~P3_INSTQUEUE_REG_3__6_ | ~new_P3_U2480;
  assign new_P3_U4595 = ~P3_INSTQUEUE_REG_4__6_ | ~new_P3_U2479;
  assign new_P3_U4596 = ~P3_INSTQUEUE_REG_5__6_ | ~new_P3_U2478;
  assign new_P3_U4597 = ~P3_INSTQUEUE_REG_6__6_ | ~new_P3_U2477;
  assign new_P3_U4598 = ~P3_INSTQUEUE_REG_7__6_ | ~new_P3_U4471;
  assign new_P3_U4599 = ~P3_INSTQUEUE_REG_8__6_ | ~new_P3_U2476;
  assign new_P3_U4600 = ~P3_INSTQUEUE_REG_9__6_ | ~new_P3_U2475;
  assign new_P3_U4601 = ~P3_INSTQUEUE_REG_10__6_ | ~new_P3_U2473;
  assign new_P3_U4602 = ~P3_INSTQUEUE_REG_11__6_ | ~new_P3_U2471;
  assign new_P3_U4603 = ~P3_INSTQUEUE_REG_12__6_ | ~new_P3_U2470;
  assign new_P3_U4604 = ~P3_INSTQUEUE_REG_13__6_ | ~new_P3_U2469;
  assign new_P3_U4605 = ~P3_INSTQUEUE_REG_14__6_ | ~new_P3_U2467;
  assign new_P3_U4606 = ~P3_INSTQUEUE_REG_15__6_ | ~new_P3_U2465;
  assign new_P3_U4607 = ~new_P3_U3074;
  assign new_P3_U4608 = ~new_P3_U3113;
  assign new_P3_U4609 = ~new_P3_U2361 | ~new_P3_U3238;
  assign new_P3_U4610 = ~new_P3_U2360 | ~new_P3_U3237;
  assign new_P3_U4611 = ~new_P3_U2357 | ~new_P3_U3212;
  assign new_P3_U4612 = ~new_P3_U4305 | ~new_P3_U3215;
  assign new_P3_U4613 = ~new_P3_U4304 | ~new_P3_U3210;
  assign new_P3_U4614 = ~new_P3_U4303 | ~new_P3_U3213;
  assign new_P3_U4615 = ~new_P3_U2356 | ~new_P3_U3211;
  assign new_P3_U4616 = ~new_P3_U4302 | ~new_P3_U3214;
  assign new_P3_U4617 = ~new_P3_U3358 | ~new_P3_U3357;
  assign new_P3_U4618 = ~new_P3_U7944 | ~new_P3_U7945 | ~new_P3_U3360 | ~new_P3_U2463 | ~new_P3_U4522;
  assign new_P3_U4619 = ~new_P3_U3109;
  assign new_P3_U4620 = ~new_P3_U4280 | ~new_P3_U4619;
  assign new_P3_U4621 = ~new_P3_U3359 | ~new_P3_U7916;
  assign new_P3_U4622 = ~new_P3_U4281;
  assign new_P3_U4623 = ~new_P3_U3262;
  assign new_P3_U4624 = P3_MORE_REG | P3_FLUSH_REG;
  assign new_P3_U4625 = ~new_P3_U3120;
  assign new_P3_U4626 = ~new_P3_U3353 | ~new_P3_U4303;
  assign new_P3_U4627 = ~new_P3_U3362 | ~new_P3_U4625;
  assign new_P3_U4628 = ~P3_STATE2_REG_1_ | ~new_U209;
  assign new_P3_U4629 = ~P3_STATE2_REG_2_ | ~new_P3_U7953 | ~new_P3_U7952;
  assign new_P3_U4630 = ~new_P3_U3122;
  assign new_P3_U4631 = ~P3_STATE2_REG_1_ | ~new_P3_U7957 | ~new_P3_U7956;
  assign new_P3_U4632 = ~P3_STATE2_REG_2_ | ~new_P3_U3122;
  assign new_P3_U4633 = ~new_P3_U4629 | ~new_P3_U4338;
  assign new_P3_U4634 = ~new_P3_U3364 | ~new_P3_U4630;
  assign new_P3_U4635 = ~P3_STATE2_REG_1_ | ~new_P3_U4633;
  assign new_P3_U4636 = ~new_P3_U2390 | ~new_P3_U4629;
  assign new_P3_U4637 = ~new_P3_U4345 | ~new_P3_U4354;
  assign new_P3_U4638 = ~new_P3_U4629 | ~new_P3_U4337;
  assign new_P3_U4639 = ~new_P3_U2390 | ~new_P3_U3120;
  assign new_P3_U4640 = ~new_P3_U3153;
  assign new_P3_U4641 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_U3128;
  assign new_P3_U4642 = ~new_P3_U3137;
  assign new_P3_U4643 = ~new_P3_U3141;
  assign new_P3_U4644 = ~new_P3_U3148;
  assign new_P3_U4645 = ~new_P3_U3155;
  assign new_P3_U4646 = ~new_P3_U3156;
  assign new_P3_U4647 = ~new_P3_U3143;
  assign new_P3_U4648 = ~new_P3_U3130;
  assign new_P3_U4649 = ~new_P3_U3132;
  assign new_P3_U4650 = ~new_P3_U3180;
  assign new_P3_U4651 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_U3132;
  assign new_P3_U4652 = ~new_P3_U3139;
  assign new_P3_U4653 = ~new_P3_U3138;
  assign new_P3_U4654 = ~new_P3_U4653 | ~new_P3_U3269;
  assign new_P3_U4655 = ~new_P3_U4654 | ~new_P3_U3139;
  assign new_P3_U4656 = ~new_P3_U3142;
  assign new_P3_U4657 = ~new_P3_U3140;
  assign new_P3_U4658 = ~new_P3_U3165;
  assign new_P3_U4659 = ~new_P3_U3140 | ~new_P3_U3142;
  assign new_P3_U4660 = ~new_P3_U3182;
  assign new_P3_U4661 = ~new_P3_U3144;
  assign new_P3_U4662 = ~new_P3_U3134;
  assign new_P3_U4663 = ~new_P3_U2457 | ~new_P3_U4653;
  assign new_P3_U4664 = ~new_P3_U3146;
  assign new_P3_U4665 = ~P3_STATE2_REG_1_ | ~new_P3_U3090;
  assign new_P3_U4666 = ~new_P3_U3126 | ~new_P3_U3124 | ~new_P3_U4665;
  assign new_P3_U4667 = ~new_P3_U4657 | ~new_P3_U2487;
  assign new_P3_U4668 = ~new_P3_U3145;
  assign new_P3_U4669 = ~new_P3_U2489 | ~new_P3_U3145;
  assign new_P3_U4670 = ~new_P3_U4664 | ~new_P3_U4669;
  assign new_P3_U4671 = ~P3_STATE2_REG_3_ | ~new_P3_U3134;
  assign new_P3_U4672 = ~new_P3_U3369 | ~new_P3_U4670;
  assign new_P3_U4673 = ~new_P3_U4668 | ~new_P3_U4322;
  assign new_P3_U4674 = ~new_P3_U2489 | ~new_P3_U4673;
  assign new_P3_U4675 = ~new_P3_U2445 | ~new_P3_U4662;
  assign new_P3_U4676 = ~new_P3_U2436 | ~new_P3_U2488;
  assign new_P3_U4677 = ~new_P3_U2435 | ~new_P3_U4661;
  assign new_P3_U4678 = ~new_P3_U2378 | ~new_P3_U2420;
  assign new_P3_U4679 = ~P3_INSTQUEUE_REG_15__7_ | ~new_P3_U4672;
  assign new_P3_U4680 = ~new_P3_U2443 | ~new_P3_U4662;
  assign new_P3_U4681 = ~new_P3_U2434 | ~new_P3_U2488;
  assign new_P3_U4682 = ~new_P3_U2433 | ~new_P3_U4661;
  assign new_P3_U4683 = ~new_P3_U2419 | ~new_P3_U2378;
  assign new_P3_U4684 = ~P3_INSTQUEUE_REG_15__6_ | ~new_P3_U4672;
  assign new_P3_U4685 = ~new_P3_U2442 | ~new_P3_U4662;
  assign new_P3_U4686 = ~new_P3_U2432 | ~new_P3_U2488;
  assign new_P3_U4687 = ~new_P3_U2431 | ~new_P3_U4661;
  assign new_P3_U4688 = ~new_P3_U2418 | ~new_P3_U2378;
  assign new_P3_U4689 = ~P3_INSTQUEUE_REG_15__5_ | ~new_P3_U4672;
  assign new_P3_U4690 = ~new_P3_U2441 | ~new_P3_U4662;
  assign new_P3_U4691 = ~new_P3_U2430 | ~new_P3_U2488;
  assign new_P3_U4692 = ~new_P3_U2429 | ~new_P3_U4661;
  assign new_P3_U4693 = ~new_P3_U2417 | ~new_P3_U2378;
  assign new_P3_U4694 = ~P3_INSTQUEUE_REG_15__4_ | ~new_P3_U4672;
  assign new_P3_U4695 = ~new_P3_U2440 | ~new_P3_U4662;
  assign new_P3_U4696 = ~new_P3_U2428 | ~new_P3_U2488;
  assign new_P3_U4697 = ~new_P3_U2427 | ~new_P3_U4661;
  assign new_P3_U4698 = ~new_P3_U2416 | ~new_P3_U2378;
  assign new_P3_U4699 = ~P3_INSTQUEUE_REG_15__3_ | ~new_P3_U4672;
  assign new_P3_U4700 = ~new_P3_U2439 | ~new_P3_U4662;
  assign new_P3_U4701 = ~new_P3_U2426 | ~new_P3_U2488;
  assign new_P3_U4702 = ~new_P3_U2425 | ~new_P3_U4661;
  assign new_P3_U4703 = ~new_P3_U2415 | ~new_P3_U2378;
  assign new_P3_U4704 = ~P3_INSTQUEUE_REG_15__2_ | ~new_P3_U4672;
  assign new_P3_U4705 = ~new_P3_U2438 | ~new_P3_U4662;
  assign new_P3_U4706 = ~new_P3_U2424 | ~new_P3_U2488;
  assign new_P3_U4707 = ~new_P3_U2423 | ~new_P3_U4661;
  assign new_P3_U4708 = ~new_P3_U2414 | ~new_P3_U2378;
  assign new_P3_U4709 = ~P3_INSTQUEUE_REG_15__1_ | ~new_P3_U4672;
  assign new_P3_U4710 = ~new_P3_U2437 | ~new_P3_U4662;
  assign new_P3_U4711 = ~new_P3_U2422 | ~new_P3_U2488;
  assign new_P3_U4712 = ~new_P3_U2421 | ~new_P3_U4661;
  assign new_P3_U4713 = ~new_P3_U2413 | ~new_P3_U2378;
  assign new_P3_U4714 = ~P3_INSTQUEUE_REG_15__0_ | ~new_P3_U4672;
  assign new_P3_U4715 = ~new_P3_U3149;
  assign new_P3_U4716 = ~new_P3_U3147;
  assign new_P3_U4717 = ~new_P3_U4342 | ~new_P3_U2457;
  assign new_P3_U4718 = ~new_P3_U3152;
  assign new_P3_U4719 = ~new_P3_U4644 | ~new_P3_U2487;
  assign new_P3_U4720 = ~new_P3_U3151;
  assign new_P3_U4721 = ~new_P3_U2489 | ~new_P3_U3151;
  assign new_P3_U4722 = ~new_P3_U4718 | ~new_P3_U4721;
  assign new_P3_U4723 = ~P3_STATE2_REG_3_ | ~new_P3_U3147;
  assign new_P3_U4724 = ~new_P3_U3387 | ~new_P3_U4722;
  assign new_P3_U4725 = ~new_P3_U4720 | ~new_P3_U4322;
  assign new_P3_U4726 = ~new_P3_U2489 | ~new_P3_U4725;
  assign new_P3_U4727 = ~new_P3_U4716 | ~new_P3_U2445;
  assign new_P3_U4728 = ~new_P3_U2491 | ~new_P3_U2436;
  assign new_P3_U4729 = ~new_P3_U4715 | ~new_P3_U2435;
  assign new_P3_U4730 = ~new_P3_U2377 | ~new_P3_U2420;
  assign new_P3_U4731 = ~P3_INSTQUEUE_REG_14__7_ | ~new_P3_U4724;
  assign new_P3_U4732 = ~new_P3_U4716 | ~new_P3_U2443;
  assign new_P3_U4733 = ~new_P3_U2491 | ~new_P3_U2434;
  assign new_P3_U4734 = ~new_P3_U4715 | ~new_P3_U2433;
  assign new_P3_U4735 = ~new_P3_U2377 | ~new_P3_U2419;
  assign new_P3_U4736 = ~P3_INSTQUEUE_REG_14__6_ | ~new_P3_U4724;
  assign new_P3_U4737 = ~new_P3_U4716 | ~new_P3_U2442;
  assign new_P3_U4738 = ~new_P3_U2491 | ~new_P3_U2432;
  assign new_P3_U4739 = ~new_P3_U4715 | ~new_P3_U2431;
  assign new_P3_U4740 = ~new_P3_U2377 | ~new_P3_U2418;
  assign new_P3_U4741 = ~P3_INSTQUEUE_REG_14__5_ | ~new_P3_U4724;
  assign new_P3_U4742 = ~new_P3_U4716 | ~new_P3_U2441;
  assign new_P3_U4743 = ~new_P3_U2491 | ~new_P3_U2430;
  assign new_P3_U4744 = ~new_P3_U4715 | ~new_P3_U2429;
  assign new_P3_U4745 = ~new_P3_U2377 | ~new_P3_U2417;
  assign new_P3_U4746 = ~P3_INSTQUEUE_REG_14__4_ | ~new_P3_U4724;
  assign new_P3_U4747 = ~new_P3_U4716 | ~new_P3_U2440;
  assign new_P3_U4748 = ~new_P3_U2491 | ~new_P3_U2428;
  assign new_P3_U4749 = ~new_P3_U4715 | ~new_P3_U2427;
  assign new_P3_U4750 = ~new_P3_U2377 | ~new_P3_U2416;
  assign new_P3_U4751 = ~P3_INSTQUEUE_REG_14__3_ | ~new_P3_U4724;
  assign new_P3_U4752 = ~new_P3_U4716 | ~new_P3_U2439;
  assign new_P3_U4753 = ~new_P3_U2491 | ~new_P3_U2426;
  assign new_P3_U4754 = ~new_P3_U4715 | ~new_P3_U2425;
  assign new_P3_U4755 = ~new_P3_U2377 | ~new_P3_U2415;
  assign new_P3_U4756 = ~P3_INSTQUEUE_REG_14__2_ | ~new_P3_U4724;
  assign new_P3_U4757 = ~new_P3_U4716 | ~new_P3_U2438;
  assign new_P3_U4758 = ~new_P3_U2491 | ~new_P3_U2424;
  assign new_P3_U4759 = ~new_P3_U4715 | ~new_P3_U2423;
  assign new_P3_U4760 = ~new_P3_U2377 | ~new_P3_U2414;
  assign new_P3_U4761 = ~P3_INSTQUEUE_REG_14__1_ | ~new_P3_U4724;
  assign new_P3_U4762 = ~new_P3_U4716 | ~new_P3_U2437;
  assign new_P3_U4763 = ~new_P3_U2491 | ~new_P3_U2422;
  assign new_P3_U4764 = ~new_P3_U4715 | ~new_P3_U2421;
  assign new_P3_U4765 = ~new_P3_U2377 | ~new_P3_U2413;
  assign new_P3_U4766 = ~P3_INSTQUEUE_REG_14__0_ | ~new_P3_U4724;
  assign new_P3_U4767 = ~new_P3_U3157;
  assign new_P3_U4768 = ~new_P3_U3154;
  assign new_P3_U4769 = ~new_P3_U4343 | ~new_P3_U2457;
  assign new_P3_U4770 = ~new_P3_U3160;
  assign new_P3_U4771 = ~new_P3_U4645 | ~new_P3_U2487;
  assign new_P3_U4772 = ~new_P3_U3159;
  assign new_P3_U4773 = ~new_P3_U2489 | ~new_P3_U3159;
  assign new_P3_U4774 = ~new_P3_U4770 | ~new_P3_U4773;
  assign new_P3_U4775 = ~P3_STATE2_REG_3_ | ~new_P3_U3154;
  assign new_P3_U4776 = ~new_P3_U3405 | ~new_P3_U4774;
  assign new_P3_U4777 = ~new_P3_U4772 | ~new_P3_U4322;
  assign new_P3_U4778 = ~new_P3_U2489 | ~new_P3_U4777;
  assign new_P3_U4779 = ~new_P3_U4768 | ~new_P3_U2445;
  assign new_P3_U4780 = ~new_P3_U2494 | ~new_P3_U2436;
  assign new_P3_U4781 = ~new_P3_U4767 | ~new_P3_U2435;
  assign new_P3_U4782 = ~new_P3_U2376 | ~new_P3_U2420;
  assign new_P3_U4783 = ~P3_INSTQUEUE_REG_13__7_ | ~new_P3_U4776;
  assign new_P3_U4784 = ~new_P3_U4768 | ~new_P3_U2443;
  assign new_P3_U4785 = ~new_P3_U2494 | ~new_P3_U2434;
  assign new_P3_U4786 = ~new_P3_U4767 | ~new_P3_U2433;
  assign new_P3_U4787 = ~new_P3_U2376 | ~new_P3_U2419;
  assign new_P3_U4788 = ~P3_INSTQUEUE_REG_13__6_ | ~new_P3_U4776;
  assign new_P3_U4789 = ~new_P3_U4768 | ~new_P3_U2442;
  assign new_P3_U4790 = ~new_P3_U2494 | ~new_P3_U2432;
  assign new_P3_U4791 = ~new_P3_U4767 | ~new_P3_U2431;
  assign new_P3_U4792 = ~new_P3_U2376 | ~new_P3_U2418;
  assign new_P3_U4793 = ~P3_INSTQUEUE_REG_13__5_ | ~new_P3_U4776;
  assign new_P3_U4794 = ~new_P3_U4768 | ~new_P3_U2441;
  assign new_P3_U4795 = ~new_P3_U2494 | ~new_P3_U2430;
  assign new_P3_U4796 = ~new_P3_U4767 | ~new_P3_U2429;
  assign new_P3_U4797 = ~new_P3_U2376 | ~new_P3_U2417;
  assign new_P3_U4798 = ~P3_INSTQUEUE_REG_13__4_ | ~new_P3_U4776;
  assign new_P3_U4799 = ~new_P3_U4768 | ~new_P3_U2440;
  assign new_P3_U4800 = ~new_P3_U2494 | ~new_P3_U2428;
  assign new_P3_U4801 = ~new_P3_U4767 | ~new_P3_U2427;
  assign new_P3_U4802 = ~new_P3_U2376 | ~new_P3_U2416;
  assign new_P3_U4803 = ~P3_INSTQUEUE_REG_13__3_ | ~new_P3_U4776;
  assign new_P3_U4804 = ~new_P3_U4768 | ~new_P3_U2439;
  assign new_P3_U4805 = ~new_P3_U2494 | ~new_P3_U2426;
  assign new_P3_U4806 = ~new_P3_U4767 | ~new_P3_U2425;
  assign new_P3_U4807 = ~new_P3_U2376 | ~new_P3_U2415;
  assign new_P3_U4808 = ~P3_INSTQUEUE_REG_13__2_ | ~new_P3_U4776;
  assign new_P3_U4809 = ~new_P3_U4768 | ~new_P3_U2438;
  assign new_P3_U4810 = ~new_P3_U2494 | ~new_P3_U2424;
  assign new_P3_U4811 = ~new_P3_U4767 | ~new_P3_U2423;
  assign new_P3_U4812 = ~new_P3_U2376 | ~new_P3_U2414;
  assign new_P3_U4813 = ~P3_INSTQUEUE_REG_13__1_ | ~new_P3_U4776;
  assign new_P3_U4814 = ~new_P3_U4768 | ~new_P3_U2437;
  assign new_P3_U4815 = ~new_P3_U2494 | ~new_P3_U2422;
  assign new_P3_U4816 = ~new_P3_U4767 | ~new_P3_U2421;
  assign new_P3_U4817 = ~new_P3_U2376 | ~new_P3_U2413;
  assign new_P3_U4818 = ~P3_INSTQUEUE_REG_13__0_ | ~new_P3_U4776;
  assign new_P3_U4819 = ~new_P3_U3162;
  assign new_P3_U4820 = ~new_P3_U3161;
  assign new_P3_U4821 = ~new_P3_U3070;
  assign new_P3_U4822 = ~new_P3_U2496 | ~new_P3_U2487;
  assign new_P3_U4823 = ~new_P3_U3163;
  assign new_P3_U4824 = ~new_P3_U2489 | ~new_P3_U3163;
  assign new_P3_U4825 = ~new_P3_U4824 | ~new_P3_U3070;
  assign new_P3_U4826 = ~P3_STATE2_REG_3_ | ~new_P3_U3161;
  assign new_P3_U4827 = ~new_P3_U3423 | ~new_P3_U4825;
  assign new_P3_U4828 = ~new_P3_U4823 | ~new_P3_U4322;
  assign new_P3_U4829 = ~new_P3_U2489 | ~new_P3_U4828;
  assign new_P3_U4830 = ~new_P3_U4820 | ~new_P3_U2445;
  assign new_P3_U4831 = ~new_P3_U2497 | ~new_P3_U2436;
  assign new_P3_U4832 = ~new_P3_U4819 | ~new_P3_U2435;
  assign new_P3_U4833 = ~new_P3_U2375 | ~new_P3_U2420;
  assign new_P3_U4834 = ~P3_INSTQUEUE_REG_12__7_ | ~new_P3_U4827;
  assign new_P3_U4835 = ~new_P3_U4820 | ~new_P3_U2443;
  assign new_P3_U4836 = ~new_P3_U2497 | ~new_P3_U2434;
  assign new_P3_U4837 = ~new_P3_U4819 | ~new_P3_U2433;
  assign new_P3_U4838 = ~new_P3_U2375 | ~new_P3_U2419;
  assign new_P3_U4839 = ~P3_INSTQUEUE_REG_12__6_ | ~new_P3_U4827;
  assign new_P3_U4840 = ~new_P3_U4820 | ~new_P3_U2442;
  assign new_P3_U4841 = ~new_P3_U2497 | ~new_P3_U2432;
  assign new_P3_U4842 = ~new_P3_U4819 | ~new_P3_U2431;
  assign new_P3_U4843 = ~new_P3_U2375 | ~new_P3_U2418;
  assign new_P3_U4844 = ~P3_INSTQUEUE_REG_12__5_ | ~new_P3_U4827;
  assign new_P3_U4845 = ~new_P3_U4820 | ~new_P3_U2441;
  assign new_P3_U4846 = ~new_P3_U2497 | ~new_P3_U2430;
  assign new_P3_U4847 = ~new_P3_U4819 | ~new_P3_U2429;
  assign new_P3_U4848 = ~new_P3_U2375 | ~new_P3_U2417;
  assign new_P3_U4849 = ~P3_INSTQUEUE_REG_12__4_ | ~new_P3_U4827;
  assign new_P3_U4850 = ~new_P3_U4820 | ~new_P3_U2440;
  assign new_P3_U4851 = ~new_P3_U2497 | ~new_P3_U2428;
  assign new_P3_U4852 = ~new_P3_U4819 | ~new_P3_U2427;
  assign new_P3_U4853 = ~new_P3_U2375 | ~new_P3_U2416;
  assign new_P3_U4854 = ~P3_INSTQUEUE_REG_12__3_ | ~new_P3_U4827;
  assign new_P3_U4855 = ~new_P3_U4820 | ~new_P3_U2439;
  assign new_P3_U4856 = ~new_P3_U2497 | ~new_P3_U2426;
  assign new_P3_U4857 = ~new_P3_U4819 | ~new_P3_U2425;
  assign new_P3_U4858 = ~new_P3_U2375 | ~new_P3_U2415;
  assign new_P3_U4859 = ~P3_INSTQUEUE_REG_12__2_ | ~new_P3_U4827;
  assign new_P3_U4860 = ~new_P3_U4820 | ~new_P3_U2438;
  assign new_P3_U4861 = ~new_P3_U2497 | ~new_P3_U2424;
  assign new_P3_U4862 = ~new_P3_U4819 | ~new_P3_U2423;
  assign new_P3_U4863 = ~new_P3_U2375 | ~new_P3_U2414;
  assign new_P3_U4864 = ~P3_INSTQUEUE_REG_12__1_ | ~new_P3_U4827;
  assign new_P3_U4865 = ~new_P3_U4820 | ~new_P3_U2437;
  assign new_P3_U4866 = ~new_P3_U2497 | ~new_P3_U2422;
  assign new_P3_U4867 = ~new_P3_U4819 | ~new_P3_U2421;
  assign new_P3_U4868 = ~new_P3_U2375 | ~new_P3_U2413;
  assign new_P3_U4869 = ~P3_INSTQUEUE_REG_12__0_ | ~new_P3_U4827;
  assign new_P3_U4870 = ~new_P3_U3166;
  assign new_P3_U4871 = ~new_P3_U3164;
  assign new_P3_U4872 = ~new_P3_U2459 | ~new_P3_U4653;
  assign new_P3_U4873 = ~new_P3_U3168;
  assign new_P3_U4874 = ~new_P3_U4658 | ~new_P3_U4657;
  assign new_P3_U4875 = ~new_P3_U3167;
  assign new_P3_U4876 = ~new_P3_U2489 | ~new_P3_U3167;
  assign new_P3_U4877 = ~new_P3_U4873 | ~new_P3_U4876;
  assign new_P3_U4878 = ~P3_STATE2_REG_3_ | ~new_P3_U3164;
  assign new_P3_U4879 = ~new_P3_U3440 | ~new_P3_U4877;
  assign new_P3_U4880 = ~new_P3_U4875 | ~new_P3_U4322;
  assign new_P3_U4881 = ~new_P3_U2489 | ~new_P3_U4880;
  assign new_P3_U4882 = ~new_P3_U4871 | ~new_P3_U2445;
  assign new_P3_U4883 = ~new_P3_U2499 | ~new_P3_U2436;
  assign new_P3_U4884 = ~new_P3_U4870 | ~new_P3_U2435;
  assign new_P3_U4885 = ~new_P3_U2374 | ~new_P3_U2420;
  assign new_P3_U4886 = ~P3_INSTQUEUE_REG_11__7_ | ~new_P3_U4879;
  assign new_P3_U4887 = ~new_P3_U4871 | ~new_P3_U2443;
  assign new_P3_U4888 = ~new_P3_U2499 | ~new_P3_U2434;
  assign new_P3_U4889 = ~new_P3_U4870 | ~new_P3_U2433;
  assign new_P3_U4890 = ~new_P3_U2374 | ~new_P3_U2419;
  assign new_P3_U4891 = ~P3_INSTQUEUE_REG_11__6_ | ~new_P3_U4879;
  assign new_P3_U4892 = ~new_P3_U4871 | ~new_P3_U2442;
  assign new_P3_U4893 = ~new_P3_U2499 | ~new_P3_U2432;
  assign new_P3_U4894 = ~new_P3_U4870 | ~new_P3_U2431;
  assign new_P3_U4895 = ~new_P3_U2374 | ~new_P3_U2418;
  assign new_P3_U4896 = ~P3_INSTQUEUE_REG_11__5_ | ~new_P3_U4879;
  assign new_P3_U4897 = ~new_P3_U4871 | ~new_P3_U2441;
  assign new_P3_U4898 = ~new_P3_U2499 | ~new_P3_U2430;
  assign new_P3_U4899 = ~new_P3_U4870 | ~new_P3_U2429;
  assign new_P3_U4900 = ~new_P3_U2374 | ~new_P3_U2417;
  assign new_P3_U4901 = ~P3_INSTQUEUE_REG_11__4_ | ~new_P3_U4879;
  assign new_P3_U4902 = ~new_P3_U4871 | ~new_P3_U2440;
  assign new_P3_U4903 = ~new_P3_U2499 | ~new_P3_U2428;
  assign new_P3_U4904 = ~new_P3_U4870 | ~new_P3_U2427;
  assign new_P3_U4905 = ~new_P3_U2374 | ~new_P3_U2416;
  assign new_P3_U4906 = ~P3_INSTQUEUE_REG_11__3_ | ~new_P3_U4879;
  assign new_P3_U4907 = ~new_P3_U4871 | ~new_P3_U2439;
  assign new_P3_U4908 = ~new_P3_U2499 | ~new_P3_U2426;
  assign new_P3_U4909 = ~new_P3_U4870 | ~new_P3_U2425;
  assign new_P3_U4910 = ~new_P3_U2374 | ~new_P3_U2415;
  assign new_P3_U4911 = ~P3_INSTQUEUE_REG_11__2_ | ~new_P3_U4879;
  assign new_P3_U4912 = ~new_P3_U4871 | ~new_P3_U2438;
  assign new_P3_U4913 = ~new_P3_U2499 | ~new_P3_U2424;
  assign new_P3_U4914 = ~new_P3_U4870 | ~new_P3_U2423;
  assign new_P3_U4915 = ~new_P3_U2374 | ~new_P3_U2414;
  assign new_P3_U4916 = ~P3_INSTQUEUE_REG_11__1_ | ~new_P3_U4879;
  assign new_P3_U4917 = ~new_P3_U4871 | ~new_P3_U2437;
  assign new_P3_U4918 = ~new_P3_U2499 | ~new_P3_U2422;
  assign new_P3_U4919 = ~new_P3_U4870 | ~new_P3_U2421;
  assign new_P3_U4920 = ~new_P3_U2374 | ~new_P3_U2413;
  assign new_P3_U4921 = ~P3_INSTQUEUE_REG_11__0_ | ~new_P3_U4879;
  assign new_P3_U4922 = ~new_P3_U3170;
  assign new_P3_U4923 = ~new_P3_U3169;
  assign new_P3_U4924 = ~new_P3_U2459 | ~new_P3_U4342;
  assign new_P3_U4925 = ~new_P3_U3172;
  assign new_P3_U4926 = ~new_P3_U4658 | ~new_P3_U4644;
  assign new_P3_U4927 = ~new_P3_U3171;
  assign new_P3_U4928 = ~new_P3_U2489 | ~new_P3_U3171;
  assign new_P3_U4929 = ~new_P3_U4925 | ~new_P3_U4928;
  assign new_P3_U4930 = ~P3_STATE2_REG_3_ | ~new_P3_U3169;
  assign new_P3_U4931 = ~new_P3_U3458 | ~new_P3_U4929;
  assign new_P3_U4932 = ~new_P3_U4927 | ~new_P3_U4322;
  assign new_P3_U4933 = ~new_P3_U2489 | ~new_P3_U4932;
  assign new_P3_U4934 = ~new_P3_U4923 | ~new_P3_U2445;
  assign new_P3_U4935 = ~new_P3_U2500 | ~new_P3_U2436;
  assign new_P3_U4936 = ~new_P3_U4922 | ~new_P3_U2435;
  assign new_P3_U4937 = ~new_P3_U2373 | ~new_P3_U2420;
  assign new_P3_U4938 = ~P3_INSTQUEUE_REG_10__7_ | ~new_P3_U4931;
  assign new_P3_U4939 = ~new_P3_U4923 | ~new_P3_U2443;
  assign new_P3_U4940 = ~new_P3_U2500 | ~new_P3_U2434;
  assign new_P3_U4941 = ~new_P3_U4922 | ~new_P3_U2433;
  assign new_P3_U4942 = ~new_P3_U2373 | ~new_P3_U2419;
  assign new_P3_U4943 = ~P3_INSTQUEUE_REG_10__6_ | ~new_P3_U4931;
  assign new_P3_U4944 = ~new_P3_U4923 | ~new_P3_U2442;
  assign new_P3_U4945 = ~new_P3_U2500 | ~new_P3_U2432;
  assign new_P3_U4946 = ~new_P3_U4922 | ~new_P3_U2431;
  assign new_P3_U4947 = ~new_P3_U2373 | ~new_P3_U2418;
  assign new_P3_U4948 = ~P3_INSTQUEUE_REG_10__5_ | ~new_P3_U4931;
  assign new_P3_U4949 = ~new_P3_U4923 | ~new_P3_U2441;
  assign new_P3_U4950 = ~new_P3_U2500 | ~new_P3_U2430;
  assign new_P3_U4951 = ~new_P3_U4922 | ~new_P3_U2429;
  assign new_P3_U4952 = ~new_P3_U2373 | ~new_P3_U2417;
  assign new_P3_U4953 = ~P3_INSTQUEUE_REG_10__4_ | ~new_P3_U4931;
  assign new_P3_U4954 = ~new_P3_U4923 | ~new_P3_U2440;
  assign new_P3_U4955 = ~new_P3_U2500 | ~new_P3_U2428;
  assign new_P3_U4956 = ~new_P3_U4922 | ~new_P3_U2427;
  assign new_P3_U4957 = ~new_P3_U2373 | ~new_P3_U2416;
  assign new_P3_U4958 = ~P3_INSTQUEUE_REG_10__3_ | ~new_P3_U4931;
  assign new_P3_U4959 = ~new_P3_U4923 | ~new_P3_U2439;
  assign new_P3_U4960 = ~new_P3_U2500 | ~new_P3_U2426;
  assign new_P3_U4961 = ~new_P3_U4922 | ~new_P3_U2425;
  assign new_P3_U4962 = ~new_P3_U2373 | ~new_P3_U2415;
  assign new_P3_U4963 = ~P3_INSTQUEUE_REG_10__2_ | ~new_P3_U4931;
  assign new_P3_U4964 = ~new_P3_U4923 | ~new_P3_U2438;
  assign new_P3_U4965 = ~new_P3_U2500 | ~new_P3_U2424;
  assign new_P3_U4966 = ~new_P3_U4922 | ~new_P3_U2423;
  assign new_P3_U4967 = ~new_P3_U2373 | ~new_P3_U2414;
  assign new_P3_U4968 = ~P3_INSTQUEUE_REG_10__1_ | ~new_P3_U4931;
  assign new_P3_U4969 = ~new_P3_U4923 | ~new_P3_U2437;
  assign new_P3_U4970 = ~new_P3_U2500 | ~new_P3_U2422;
  assign new_P3_U4971 = ~new_P3_U4922 | ~new_P3_U2421;
  assign new_P3_U4972 = ~new_P3_U2373 | ~new_P3_U2413;
  assign new_P3_U4973 = ~P3_INSTQUEUE_REG_10__0_ | ~new_P3_U4931;
  assign new_P3_U4974 = ~new_P3_U3174;
  assign new_P3_U4975 = ~new_P3_U3173;
  assign new_P3_U4976 = ~new_P3_U2459 | ~new_P3_U4343;
  assign new_P3_U4977 = ~new_P3_U3176;
  assign new_P3_U4978 = ~new_P3_U4658 | ~new_P3_U4645;
  assign new_P3_U4979 = ~new_P3_U3175;
  assign new_P3_U4980 = ~new_P3_U2489 | ~new_P3_U3175;
  assign new_P3_U4981 = ~new_P3_U4977 | ~new_P3_U4980;
  assign new_P3_U4982 = ~P3_STATE2_REG_3_ | ~new_P3_U3173;
  assign new_P3_U4983 = ~new_P3_U3476 | ~new_P3_U4981;
  assign new_P3_U4984 = ~new_P3_U4979 | ~new_P3_U4322;
  assign new_P3_U4985 = ~new_P3_U2489 | ~new_P3_U4984;
  assign new_P3_U4986 = ~new_P3_U4975 | ~new_P3_U2445;
  assign new_P3_U4987 = ~new_P3_U2502 | ~new_P3_U2436;
  assign new_P3_U4988 = ~new_P3_U4974 | ~new_P3_U2435;
  assign new_P3_U4989 = ~new_P3_U2372 | ~new_P3_U2420;
  assign new_P3_U4990 = ~P3_INSTQUEUE_REG_9__7_ | ~new_P3_U4983;
  assign new_P3_U4991 = ~new_P3_U4975 | ~new_P3_U2443;
  assign new_P3_U4992 = ~new_P3_U2502 | ~new_P3_U2434;
  assign new_P3_U4993 = ~new_P3_U4974 | ~new_P3_U2433;
  assign new_P3_U4994 = ~new_P3_U2372 | ~new_P3_U2419;
  assign new_P3_U4995 = ~P3_INSTQUEUE_REG_9__6_ | ~new_P3_U4983;
  assign new_P3_U4996 = ~new_P3_U4975 | ~new_P3_U2442;
  assign new_P3_U4997 = ~new_P3_U2502 | ~new_P3_U2432;
  assign new_P3_U4998 = ~new_P3_U4974 | ~new_P3_U2431;
  assign new_P3_U4999 = ~new_P3_U2372 | ~new_P3_U2418;
  assign new_P3_U5000 = ~P3_INSTQUEUE_REG_9__5_ | ~new_P3_U4983;
  assign new_P3_U5001 = ~new_P3_U4975 | ~new_P3_U2441;
  assign new_P3_U5002 = ~new_P3_U2502 | ~new_P3_U2430;
  assign new_P3_U5003 = ~new_P3_U4974 | ~new_P3_U2429;
  assign new_P3_U5004 = ~new_P3_U2372 | ~new_P3_U2417;
  assign new_P3_U5005 = ~P3_INSTQUEUE_REG_9__4_ | ~new_P3_U4983;
  assign new_P3_U5006 = ~new_P3_U4975 | ~new_P3_U2440;
  assign new_P3_U5007 = ~new_P3_U2502 | ~new_P3_U2428;
  assign new_P3_U5008 = ~new_P3_U4974 | ~new_P3_U2427;
  assign new_P3_U5009 = ~new_P3_U2372 | ~new_P3_U2416;
  assign new_P3_U5010 = ~P3_INSTQUEUE_REG_9__3_ | ~new_P3_U4983;
  assign new_P3_U5011 = ~new_P3_U4975 | ~new_P3_U2439;
  assign new_P3_U5012 = ~new_P3_U2502 | ~new_P3_U2426;
  assign new_P3_U5013 = ~new_P3_U4974 | ~new_P3_U2425;
  assign new_P3_U5014 = ~new_P3_U2372 | ~new_P3_U2415;
  assign new_P3_U5015 = ~P3_INSTQUEUE_REG_9__2_ | ~new_P3_U4983;
  assign new_P3_U5016 = ~new_P3_U4975 | ~new_P3_U2438;
  assign new_P3_U5017 = ~new_P3_U2502 | ~new_P3_U2424;
  assign new_P3_U5018 = ~new_P3_U4974 | ~new_P3_U2423;
  assign new_P3_U5019 = ~new_P3_U2372 | ~new_P3_U2414;
  assign new_P3_U5020 = ~P3_INSTQUEUE_REG_9__1_ | ~new_P3_U4983;
  assign new_P3_U5021 = ~new_P3_U4975 | ~new_P3_U2437;
  assign new_P3_U5022 = ~new_P3_U2502 | ~new_P3_U2422;
  assign new_P3_U5023 = ~new_P3_U4974 | ~new_P3_U2421;
  assign new_P3_U5024 = ~new_P3_U2372 | ~new_P3_U2413;
  assign new_P3_U5025 = ~P3_INSTQUEUE_REG_9__0_ | ~new_P3_U4983;
  assign new_P3_U5026 = ~new_P3_U3178;
  assign new_P3_U5027 = ~new_P3_U3177;
  assign new_P3_U5028 = ~new_P3_U3071;
  assign new_P3_U5029 = ~new_P3_U4658 | ~new_P3_U2496;
  assign new_P3_U5030 = ~new_P3_U3179;
  assign new_P3_U5031 = ~new_P3_U2489 | ~new_P3_U3179;
  assign new_P3_U5032 = ~new_P3_U5031 | ~new_P3_U3071;
  assign new_P3_U5033 = ~P3_STATE2_REG_3_ | ~new_P3_U3177;
  assign new_P3_U5034 = ~new_P3_U3493 | ~new_P3_U5032;
  assign new_P3_U5035 = ~new_P3_U5030 | ~new_P3_U4322;
  assign new_P3_U5036 = ~new_P3_U2489 | ~new_P3_U5035;
  assign new_P3_U5037 = ~new_P3_U5027 | ~new_P3_U2445;
  assign new_P3_U5038 = ~new_P3_U2503 | ~new_P3_U2436;
  assign new_P3_U5039 = ~new_P3_U5026 | ~new_P3_U2435;
  assign new_P3_U5040 = ~new_P3_U2371 | ~new_P3_U2420;
  assign new_P3_U5041 = ~P3_INSTQUEUE_REG_8__7_ | ~new_P3_U5034;
  assign new_P3_U5042 = ~new_P3_U5027 | ~new_P3_U2443;
  assign new_P3_U5043 = ~new_P3_U2503 | ~new_P3_U2434;
  assign new_P3_U5044 = ~new_P3_U5026 | ~new_P3_U2433;
  assign new_P3_U5045 = ~new_P3_U2371 | ~new_P3_U2419;
  assign new_P3_U5046 = ~P3_INSTQUEUE_REG_8__6_ | ~new_P3_U5034;
  assign new_P3_U5047 = ~new_P3_U5027 | ~new_P3_U2442;
  assign new_P3_U5048 = ~new_P3_U2503 | ~new_P3_U2432;
  assign new_P3_U5049 = ~new_P3_U5026 | ~new_P3_U2431;
  assign new_P3_U5050 = ~new_P3_U2371 | ~new_P3_U2418;
  assign new_P3_U5051 = ~P3_INSTQUEUE_REG_8__5_ | ~new_P3_U5034;
  assign new_P3_U5052 = ~new_P3_U5027 | ~new_P3_U2441;
  assign new_P3_U5053 = ~new_P3_U2503 | ~new_P3_U2430;
  assign new_P3_U5054 = ~new_P3_U5026 | ~new_P3_U2429;
  assign new_P3_U5055 = ~new_P3_U2371 | ~new_P3_U2417;
  assign new_P3_U5056 = ~P3_INSTQUEUE_REG_8__4_ | ~new_P3_U5034;
  assign new_P3_U5057 = ~new_P3_U5027 | ~new_P3_U2440;
  assign new_P3_U5058 = ~new_P3_U2503 | ~new_P3_U2428;
  assign new_P3_U5059 = ~new_P3_U5026 | ~new_P3_U2427;
  assign new_P3_U5060 = ~new_P3_U2371 | ~new_P3_U2416;
  assign new_P3_U5061 = ~P3_INSTQUEUE_REG_8__3_ | ~new_P3_U5034;
  assign new_P3_U5062 = ~new_P3_U5027 | ~new_P3_U2439;
  assign new_P3_U5063 = ~new_P3_U2503 | ~new_P3_U2426;
  assign new_P3_U5064 = ~new_P3_U5026 | ~new_P3_U2425;
  assign new_P3_U5065 = ~new_P3_U2371 | ~new_P3_U2415;
  assign new_P3_U5066 = ~P3_INSTQUEUE_REG_8__2_ | ~new_P3_U5034;
  assign new_P3_U5067 = ~new_P3_U5027 | ~new_P3_U2438;
  assign new_P3_U5068 = ~new_P3_U2503 | ~new_P3_U2424;
  assign new_P3_U5069 = ~new_P3_U5026 | ~new_P3_U2423;
  assign new_P3_U5070 = ~new_P3_U2371 | ~new_P3_U2414;
  assign new_P3_U5071 = ~P3_INSTQUEUE_REG_8__1_ | ~new_P3_U5034;
  assign new_P3_U5072 = ~new_P3_U5027 | ~new_P3_U2437;
  assign new_P3_U5073 = ~new_P3_U2503 | ~new_P3_U2422;
  assign new_P3_U5074 = ~new_P3_U5026 | ~new_P3_U2421;
  assign new_P3_U5075 = ~new_P3_U2371 | ~new_P3_U2413;
  assign new_P3_U5076 = ~P3_INSTQUEUE_REG_8__0_ | ~new_P3_U5034;
  assign new_P3_U5077 = ~new_P3_U3183;
  assign new_P3_U5078 = ~new_P3_U3185;
  assign new_P3_U5079 = ~new_P3_U3184;
  assign new_P3_U5080 = ~new_P3_U2489 | ~new_P3_U3184;
  assign new_P3_U5081 = ~new_P3_U5078 | ~new_P3_U5080;
  assign new_P3_U5082 = ~P3_STATE2_REG_3_ | ~new_P3_U3180;
  assign new_P3_U5083 = ~new_P3_U3510 | ~new_P3_U5081;
  assign new_P3_U5084 = ~new_P3_U5079 | ~new_P3_U4322;
  assign new_P3_U5085 = ~new_P3_U2489 | ~new_P3_U5084;
  assign new_P3_U5086 = ~new_P3_U4650 | ~new_P3_U2445;
  assign new_P3_U5087 = ~new_P3_U4326 | ~new_P3_U2436;
  assign new_P3_U5088 = ~new_P3_U5077 | ~new_P3_U2435;
  assign new_P3_U5089 = ~new_P3_U2370 | ~new_P3_U2420;
  assign new_P3_U5090 = ~P3_INSTQUEUE_REG_7__7_ | ~new_P3_U5083;
  assign new_P3_U5091 = ~new_P3_U4650 | ~new_P3_U2443;
  assign new_P3_U5092 = ~new_P3_U4326 | ~new_P3_U2434;
  assign new_P3_U5093 = ~new_P3_U5077 | ~new_P3_U2433;
  assign new_P3_U5094 = ~new_P3_U2370 | ~new_P3_U2419;
  assign new_P3_U5095 = ~P3_INSTQUEUE_REG_7__6_ | ~new_P3_U5083;
  assign new_P3_U5096 = ~new_P3_U4650 | ~new_P3_U2442;
  assign new_P3_U5097 = ~new_P3_U4326 | ~new_P3_U2432;
  assign new_P3_U5098 = ~new_P3_U5077 | ~new_P3_U2431;
  assign new_P3_U5099 = ~new_P3_U2370 | ~new_P3_U2418;
  assign new_P3_U5100 = ~P3_INSTQUEUE_REG_7__5_ | ~new_P3_U5083;
  assign new_P3_U5101 = ~new_P3_U4650 | ~new_P3_U2441;
  assign new_P3_U5102 = ~new_P3_U4326 | ~new_P3_U2430;
  assign new_P3_U5103 = ~new_P3_U5077 | ~new_P3_U2429;
  assign new_P3_U5104 = ~new_P3_U2370 | ~new_P3_U2417;
  assign new_P3_U5105 = ~P3_INSTQUEUE_REG_7__4_ | ~new_P3_U5083;
  assign new_P3_U5106 = ~new_P3_U4650 | ~new_P3_U2440;
  assign new_P3_U5107 = ~new_P3_U4326 | ~new_P3_U2428;
  assign new_P3_U5108 = ~new_P3_U5077 | ~new_P3_U2427;
  assign new_P3_U5109 = ~new_P3_U2370 | ~new_P3_U2416;
  assign new_P3_U5110 = ~P3_INSTQUEUE_REG_7__3_ | ~new_P3_U5083;
  assign new_P3_U5111 = ~new_P3_U4650 | ~new_P3_U2439;
  assign new_P3_U5112 = ~new_P3_U4326 | ~new_P3_U2426;
  assign new_P3_U5113 = ~new_P3_U5077 | ~new_P3_U2425;
  assign new_P3_U5114 = ~new_P3_U2370 | ~new_P3_U2415;
  assign new_P3_U5115 = ~P3_INSTQUEUE_REG_7__2_ | ~new_P3_U5083;
  assign new_P3_U5116 = ~new_P3_U4650 | ~new_P3_U2438;
  assign new_P3_U5117 = ~new_P3_U4326 | ~new_P3_U2424;
  assign new_P3_U5118 = ~new_P3_U5077 | ~new_P3_U2423;
  assign new_P3_U5119 = ~new_P3_U2370 | ~new_P3_U2414;
  assign new_P3_U5120 = ~P3_INSTQUEUE_REG_7__1_ | ~new_P3_U5083;
  assign new_P3_U5121 = ~new_P3_U4650 | ~new_P3_U2437;
  assign new_P3_U5122 = ~new_P3_U4326 | ~new_P3_U2422;
  assign new_P3_U5123 = ~new_P3_U5077 | ~new_P3_U2421;
  assign new_P3_U5124 = ~new_P3_U2370 | ~new_P3_U2413;
  assign new_P3_U5125 = ~P3_INSTQUEUE_REG_7__0_ | ~new_P3_U5083;
  assign new_P3_U5126 = ~new_P3_U3187;
  assign new_P3_U5127 = ~new_P3_U3186;
  assign new_P3_U5128 = ~new_P3_U4342 | ~new_P3_U2458;
  assign new_P3_U5129 = ~new_P3_U3189;
  assign new_P3_U5130 = ~new_P3_U4644 | ~new_P3_U2485;
  assign new_P3_U5131 = ~new_P3_U3188;
  assign new_P3_U5132 = ~new_P3_U2489 | ~new_P3_U3188;
  assign new_P3_U5133 = ~new_P3_U5129 | ~new_P3_U5132;
  assign new_P3_U5134 = ~P3_STATE2_REG_3_ | ~new_P3_U3186;
  assign new_P3_U5135 = ~new_P3_U3528 | ~new_P3_U5133;
  assign new_P3_U5136 = ~new_P3_U5131 | ~new_P3_U4322;
  assign new_P3_U5137 = ~new_P3_U2489 | ~new_P3_U5136;
  assign new_P3_U5138 = ~new_P3_U5127 | ~new_P3_U2445;
  assign new_P3_U5139 = ~new_P3_U2505 | ~new_P3_U2436;
  assign new_P3_U5140 = ~new_P3_U5126 | ~new_P3_U2435;
  assign new_P3_U5141 = ~new_P3_U2369 | ~new_P3_U2420;
  assign new_P3_U5142 = ~P3_INSTQUEUE_REG_6__7_ | ~new_P3_U5135;
  assign new_P3_U5143 = ~new_P3_U5127 | ~new_P3_U2443;
  assign new_P3_U5144 = ~new_P3_U2505 | ~new_P3_U2434;
  assign new_P3_U5145 = ~new_P3_U5126 | ~new_P3_U2433;
  assign new_P3_U5146 = ~new_P3_U2369 | ~new_P3_U2419;
  assign new_P3_U5147 = ~P3_INSTQUEUE_REG_6__6_ | ~new_P3_U5135;
  assign new_P3_U5148 = ~new_P3_U5127 | ~new_P3_U2442;
  assign new_P3_U5149 = ~new_P3_U2505 | ~new_P3_U2432;
  assign new_P3_U5150 = ~new_P3_U5126 | ~new_P3_U2431;
  assign new_P3_U5151 = ~new_P3_U2369 | ~new_P3_U2418;
  assign new_P3_U5152 = ~P3_INSTQUEUE_REG_6__5_ | ~new_P3_U5135;
  assign new_P3_U5153 = ~new_P3_U5127 | ~new_P3_U2441;
  assign new_P3_U5154 = ~new_P3_U2505 | ~new_P3_U2430;
  assign new_P3_U5155 = ~new_P3_U5126 | ~new_P3_U2429;
  assign new_P3_U5156 = ~new_P3_U2369 | ~new_P3_U2417;
  assign new_P3_U5157 = ~P3_INSTQUEUE_REG_6__4_ | ~new_P3_U5135;
  assign new_P3_U5158 = ~new_P3_U5127 | ~new_P3_U2440;
  assign new_P3_U5159 = ~new_P3_U2505 | ~new_P3_U2428;
  assign new_P3_U5160 = ~new_P3_U5126 | ~new_P3_U2427;
  assign new_P3_U5161 = ~new_P3_U2369 | ~new_P3_U2416;
  assign new_P3_U5162 = ~P3_INSTQUEUE_REG_6__3_ | ~new_P3_U5135;
  assign new_P3_U5163 = ~new_P3_U5127 | ~new_P3_U2439;
  assign new_P3_U5164 = ~new_P3_U2505 | ~new_P3_U2426;
  assign new_P3_U5165 = ~new_P3_U5126 | ~new_P3_U2425;
  assign new_P3_U5166 = ~new_P3_U2369 | ~new_P3_U2415;
  assign new_P3_U5167 = ~P3_INSTQUEUE_REG_6__2_ | ~new_P3_U5135;
  assign new_P3_U5168 = ~new_P3_U5127 | ~new_P3_U2438;
  assign new_P3_U5169 = ~new_P3_U2505 | ~new_P3_U2424;
  assign new_P3_U5170 = ~new_P3_U5126 | ~new_P3_U2423;
  assign new_P3_U5171 = ~new_P3_U2369 | ~new_P3_U2414;
  assign new_P3_U5172 = ~P3_INSTQUEUE_REG_6__1_ | ~new_P3_U5135;
  assign new_P3_U5173 = ~new_P3_U5127 | ~new_P3_U2437;
  assign new_P3_U5174 = ~new_P3_U2505 | ~new_P3_U2422;
  assign new_P3_U5175 = ~new_P3_U5126 | ~new_P3_U2421;
  assign new_P3_U5176 = ~new_P3_U2369 | ~new_P3_U2413;
  assign new_P3_U5177 = ~P3_INSTQUEUE_REG_6__0_ | ~new_P3_U5135;
  assign new_P3_U5178 = ~new_P3_U3191;
  assign new_P3_U5179 = ~new_P3_U3190;
  assign new_P3_U5180 = ~new_P3_U4343 | ~new_P3_U2458;
  assign new_P3_U5181 = ~new_P3_U3193;
  assign new_P3_U5182 = ~new_P3_U4645 | ~new_P3_U2485;
  assign new_P3_U5183 = ~new_P3_U3192;
  assign new_P3_U5184 = ~new_P3_U2489 | ~new_P3_U3192;
  assign new_P3_U5185 = ~new_P3_U5181 | ~new_P3_U5184;
  assign new_P3_U5186 = ~P3_STATE2_REG_3_ | ~new_P3_U3190;
  assign new_P3_U5187 = ~new_P3_U3546 | ~new_P3_U5185;
  assign new_P3_U5188 = ~new_P3_U5183 | ~new_P3_U4322;
  assign new_P3_U5189 = ~new_P3_U2489 | ~new_P3_U5188;
  assign new_P3_U5190 = ~new_P3_U5179 | ~new_P3_U2445;
  assign new_P3_U5191 = ~new_P3_U2506 | ~new_P3_U2436;
  assign new_P3_U5192 = ~new_P3_U5178 | ~new_P3_U2435;
  assign new_P3_U5193 = ~new_P3_U2368 | ~new_P3_U2420;
  assign new_P3_U5194 = ~P3_INSTQUEUE_REG_5__7_ | ~new_P3_U5187;
  assign new_P3_U5195 = ~new_P3_U5179 | ~new_P3_U2443;
  assign new_P3_U5196 = ~new_P3_U2506 | ~new_P3_U2434;
  assign new_P3_U5197 = ~new_P3_U5178 | ~new_P3_U2433;
  assign new_P3_U5198 = ~new_P3_U2368 | ~new_P3_U2419;
  assign new_P3_U5199 = ~P3_INSTQUEUE_REG_5__6_ | ~new_P3_U5187;
  assign new_P3_U5200 = ~new_P3_U5179 | ~new_P3_U2442;
  assign new_P3_U5201 = ~new_P3_U2506 | ~new_P3_U2432;
  assign new_P3_U5202 = ~new_P3_U5178 | ~new_P3_U2431;
  assign new_P3_U5203 = ~new_P3_U2368 | ~new_P3_U2418;
  assign new_P3_U5204 = ~P3_INSTQUEUE_REG_5__5_ | ~new_P3_U5187;
  assign new_P3_U5205 = ~new_P3_U5179 | ~new_P3_U2441;
  assign new_P3_U5206 = ~new_P3_U2506 | ~new_P3_U2430;
  assign new_P3_U5207 = ~new_P3_U5178 | ~new_P3_U2429;
  assign new_P3_U5208 = ~new_P3_U2368 | ~new_P3_U2417;
  assign new_P3_U5209 = ~P3_INSTQUEUE_REG_5__4_ | ~new_P3_U5187;
  assign new_P3_U5210 = ~new_P3_U5179 | ~new_P3_U2440;
  assign new_P3_U5211 = ~new_P3_U2506 | ~new_P3_U2428;
  assign new_P3_U5212 = ~new_P3_U5178 | ~new_P3_U2427;
  assign new_P3_U5213 = ~new_P3_U2368 | ~new_P3_U2416;
  assign new_P3_U5214 = ~P3_INSTQUEUE_REG_5__3_ | ~new_P3_U5187;
  assign new_P3_U5215 = ~new_P3_U5179 | ~new_P3_U2439;
  assign new_P3_U5216 = ~new_P3_U2506 | ~new_P3_U2426;
  assign new_P3_U5217 = ~new_P3_U5178 | ~new_P3_U2425;
  assign new_P3_U5218 = ~new_P3_U2368 | ~new_P3_U2415;
  assign new_P3_U5219 = ~P3_INSTQUEUE_REG_5__2_ | ~new_P3_U5187;
  assign new_P3_U5220 = ~new_P3_U5179 | ~new_P3_U2438;
  assign new_P3_U5221 = ~new_P3_U2506 | ~new_P3_U2424;
  assign new_P3_U5222 = ~new_P3_U5178 | ~new_P3_U2423;
  assign new_P3_U5223 = ~new_P3_U2368 | ~new_P3_U2414;
  assign new_P3_U5224 = ~P3_INSTQUEUE_REG_5__1_ | ~new_P3_U5187;
  assign new_P3_U5225 = ~new_P3_U5179 | ~new_P3_U2437;
  assign new_P3_U5226 = ~new_P3_U2506 | ~new_P3_U2422;
  assign new_P3_U5227 = ~new_P3_U5178 | ~new_P3_U2421;
  assign new_P3_U5228 = ~new_P3_U2368 | ~new_P3_U2413;
  assign new_P3_U5229 = ~P3_INSTQUEUE_REG_5__0_ | ~new_P3_U5187;
  assign new_P3_U5230 = ~new_P3_U3195;
  assign new_P3_U5231 = ~new_P3_U3194;
  assign new_P3_U5232 = ~new_P3_U3072;
  assign new_P3_U5233 = ~new_P3_U2496 | ~new_P3_U2485;
  assign new_P3_U5234 = ~new_P3_U3195 | ~new_P3_U5233;
  assign new_P3_U5235 = ~new_P3_U2489 | ~new_P3_U5234;
  assign new_P3_U5236 = ~new_P3_U5235 | ~new_P3_U3072;
  assign new_P3_U5237 = ~P3_STATE2_REG_3_ | ~new_P3_U3194;
  assign new_P3_U5238 = ~new_P3_U3564 | ~new_P3_U5236;
  assign new_P3_U5239 = ~new_P3_U2489 | ~new_P3_U3136;
  assign new_P3_U5240 = ~new_P3_U5231 | ~new_P3_U2445;
  assign new_P3_U5241 = ~new_P3_U2507 | ~new_P3_U2436;
  assign new_P3_U5242 = ~new_P3_U5230 | ~new_P3_U2435;
  assign new_P3_U5243 = ~new_P3_U2367 | ~new_P3_U2420;
  assign new_P3_U5244 = ~P3_INSTQUEUE_REG_4__7_ | ~new_P3_U5238;
  assign new_P3_U5245 = ~new_P3_U5231 | ~new_P3_U2443;
  assign new_P3_U5246 = ~new_P3_U2507 | ~new_P3_U2434;
  assign new_P3_U5247 = ~new_P3_U5230 | ~new_P3_U2433;
  assign new_P3_U5248 = ~new_P3_U2367 | ~new_P3_U2419;
  assign new_P3_U5249 = ~P3_INSTQUEUE_REG_4__6_ | ~new_P3_U5238;
  assign new_P3_U5250 = ~new_P3_U5231 | ~new_P3_U2442;
  assign new_P3_U5251 = ~new_P3_U2507 | ~new_P3_U2432;
  assign new_P3_U5252 = ~new_P3_U5230 | ~new_P3_U2431;
  assign new_P3_U5253 = ~new_P3_U2367 | ~new_P3_U2418;
  assign new_P3_U5254 = ~P3_INSTQUEUE_REG_4__5_ | ~new_P3_U5238;
  assign new_P3_U5255 = ~new_P3_U5231 | ~new_P3_U2441;
  assign new_P3_U5256 = ~new_P3_U2507 | ~new_P3_U2430;
  assign new_P3_U5257 = ~new_P3_U5230 | ~new_P3_U2429;
  assign new_P3_U5258 = ~new_P3_U2367 | ~new_P3_U2417;
  assign new_P3_U5259 = ~P3_INSTQUEUE_REG_4__4_ | ~new_P3_U5238;
  assign new_P3_U5260 = ~new_P3_U5231 | ~new_P3_U2440;
  assign new_P3_U5261 = ~new_P3_U2507 | ~new_P3_U2428;
  assign new_P3_U5262 = ~new_P3_U5230 | ~new_P3_U2427;
  assign new_P3_U5263 = ~new_P3_U2367 | ~new_P3_U2416;
  assign new_P3_U5264 = ~P3_INSTQUEUE_REG_4__3_ | ~new_P3_U5238;
  assign new_P3_U5265 = ~new_P3_U5231 | ~new_P3_U2439;
  assign new_P3_U5266 = ~new_P3_U2507 | ~new_P3_U2426;
  assign new_P3_U5267 = ~new_P3_U5230 | ~new_P3_U2425;
  assign new_P3_U5268 = ~new_P3_U2367 | ~new_P3_U2415;
  assign new_P3_U5269 = ~P3_INSTQUEUE_REG_4__2_ | ~new_P3_U5238;
  assign new_P3_U5270 = ~new_P3_U5231 | ~new_P3_U2438;
  assign new_P3_U5271 = ~new_P3_U2507 | ~new_P3_U2424;
  assign new_P3_U5272 = ~new_P3_U5230 | ~new_P3_U2423;
  assign new_P3_U5273 = ~new_P3_U2367 | ~new_P3_U2414;
  assign new_P3_U5274 = ~P3_INSTQUEUE_REG_4__1_ | ~new_P3_U5238;
  assign new_P3_U5275 = ~new_P3_U5231 | ~new_P3_U2437;
  assign new_P3_U5276 = ~new_P3_U2507 | ~new_P3_U2422;
  assign new_P3_U5277 = ~new_P3_U5230 | ~new_P3_U2421;
  assign new_P3_U5278 = ~new_P3_U2367 | ~new_P3_U2413;
  assign new_P3_U5279 = ~P3_INSTQUEUE_REG_4__0_ | ~new_P3_U5238;
  assign new_P3_U5280 = ~new_P3_U3197;
  assign new_P3_U5281 = ~new_P3_U3196;
  assign new_P3_U5282 = ~new_P3_U2460 | ~new_P3_U4653;
  assign new_P3_U5283 = ~new_P3_U3198;
  assign new_P3_U5284 = ~new_P3_U2509 | ~new_P3_U4657;
  assign new_P3_U5285 = ~new_P3_U3197 | ~new_P3_U5284;
  assign new_P3_U5286 = ~new_P3_U2489 | ~new_P3_U5285;
  assign new_P3_U5287 = ~new_P3_U5283 | ~new_P3_U5286;
  assign new_P3_U5288 = ~P3_STATE2_REG_3_ | ~new_P3_U3196;
  assign new_P3_U5289 = ~new_P3_U3582 | ~new_P3_U5287;
  assign new_P3_U5290 = ~new_P3_U2489 | ~new_P3_U3136;
  assign new_P3_U5291 = ~new_P3_U5281 | ~new_P3_U2445;
  assign new_P3_U5292 = ~new_P3_U2510 | ~new_P3_U2436;
  assign new_P3_U5293 = ~new_P3_U5280 | ~new_P3_U2435;
  assign new_P3_U5294 = ~new_P3_U2366 | ~new_P3_U2420;
  assign new_P3_U5295 = ~P3_INSTQUEUE_REG_3__7_ | ~new_P3_U5289;
  assign new_P3_U5296 = ~new_P3_U5281 | ~new_P3_U2443;
  assign new_P3_U5297 = ~new_P3_U2510 | ~new_P3_U2434;
  assign new_P3_U5298 = ~new_P3_U5280 | ~new_P3_U2433;
  assign new_P3_U5299 = ~new_P3_U2366 | ~new_P3_U2419;
  assign new_P3_U5300 = ~P3_INSTQUEUE_REG_3__6_ | ~new_P3_U5289;
  assign new_P3_U5301 = ~new_P3_U5281 | ~new_P3_U2442;
  assign new_P3_U5302 = ~new_P3_U2510 | ~new_P3_U2432;
  assign new_P3_U5303 = ~new_P3_U5280 | ~new_P3_U2431;
  assign new_P3_U5304 = ~new_P3_U2366 | ~new_P3_U2418;
  assign new_P3_U5305 = ~P3_INSTQUEUE_REG_3__5_ | ~new_P3_U5289;
  assign new_P3_U5306 = ~new_P3_U5281 | ~new_P3_U2441;
  assign new_P3_U5307 = ~new_P3_U2510 | ~new_P3_U2430;
  assign new_P3_U5308 = ~new_P3_U5280 | ~new_P3_U2429;
  assign new_P3_U5309 = ~new_P3_U2366 | ~new_P3_U2417;
  assign new_P3_U5310 = ~P3_INSTQUEUE_REG_3__4_ | ~new_P3_U5289;
  assign new_P3_U5311 = ~new_P3_U5281 | ~new_P3_U2440;
  assign new_P3_U5312 = ~new_P3_U2510 | ~new_P3_U2428;
  assign new_P3_U5313 = ~new_P3_U5280 | ~new_P3_U2427;
  assign new_P3_U5314 = ~new_P3_U2366 | ~new_P3_U2416;
  assign new_P3_U5315 = ~P3_INSTQUEUE_REG_3__3_ | ~new_P3_U5289;
  assign new_P3_U5316 = ~new_P3_U5281 | ~new_P3_U2439;
  assign new_P3_U5317 = ~new_P3_U2510 | ~new_P3_U2426;
  assign new_P3_U5318 = ~new_P3_U5280 | ~new_P3_U2425;
  assign new_P3_U5319 = ~new_P3_U2366 | ~new_P3_U2415;
  assign new_P3_U5320 = ~P3_INSTQUEUE_REG_3__2_ | ~new_P3_U5289;
  assign new_P3_U5321 = ~new_P3_U5281 | ~new_P3_U2438;
  assign new_P3_U5322 = ~new_P3_U2510 | ~new_P3_U2424;
  assign new_P3_U5323 = ~new_P3_U5280 | ~new_P3_U2423;
  assign new_P3_U5324 = ~new_P3_U2366 | ~new_P3_U2414;
  assign new_P3_U5325 = ~P3_INSTQUEUE_REG_3__1_ | ~new_P3_U5289;
  assign new_P3_U5326 = ~new_P3_U5281 | ~new_P3_U2437;
  assign new_P3_U5327 = ~new_P3_U2510 | ~new_P3_U2422;
  assign new_P3_U5328 = ~new_P3_U5280 | ~new_P3_U2421;
  assign new_P3_U5329 = ~new_P3_U2366 | ~new_P3_U2413;
  assign new_P3_U5330 = ~P3_INSTQUEUE_REG_3__0_ | ~new_P3_U5289;
  assign new_P3_U5331 = ~new_P3_U3200;
  assign new_P3_U5332 = ~new_P3_U3199;
  assign new_P3_U5333 = ~new_P3_U2460 | ~new_P3_U4342;
  assign new_P3_U5334 = ~new_P3_U3201;
  assign new_P3_U5335 = ~new_P3_U2509 | ~new_P3_U4644;
  assign new_P3_U5336 = ~new_P3_U3200 | ~new_P3_U5335;
  assign new_P3_U5337 = ~new_P3_U2489 | ~new_P3_U5336;
  assign new_P3_U5338 = ~new_P3_U5334 | ~new_P3_U5337;
  assign new_P3_U5339 = ~P3_STATE2_REG_3_ | ~new_P3_U3199;
  assign new_P3_U5340 = ~new_P3_U3599 | ~new_P3_U5338;
  assign new_P3_U5341 = ~new_P3_U2489 | ~new_P3_U3136;
  assign new_P3_U5342 = ~new_P3_U5332 | ~new_P3_U2445;
  assign new_P3_U5343 = ~new_P3_U2511 | ~new_P3_U2436;
  assign new_P3_U5344 = ~new_P3_U5331 | ~new_P3_U2435;
  assign new_P3_U5345 = ~new_P3_U2365 | ~new_P3_U2420;
  assign new_P3_U5346 = ~P3_INSTQUEUE_REG_2__7_ | ~new_P3_U5340;
  assign new_P3_U5347 = ~new_P3_U5332 | ~new_P3_U2443;
  assign new_P3_U5348 = ~new_P3_U2511 | ~new_P3_U2434;
  assign new_P3_U5349 = ~new_P3_U5331 | ~new_P3_U2433;
  assign new_P3_U5350 = ~new_P3_U2365 | ~new_P3_U2419;
  assign new_P3_U5351 = ~P3_INSTQUEUE_REG_2__6_ | ~new_P3_U5340;
  assign new_P3_U5352 = ~new_P3_U5332 | ~new_P3_U2442;
  assign new_P3_U5353 = ~new_P3_U2511 | ~new_P3_U2432;
  assign new_P3_U5354 = ~new_P3_U5331 | ~new_P3_U2431;
  assign new_P3_U5355 = ~new_P3_U2365 | ~new_P3_U2418;
  assign new_P3_U5356 = ~P3_INSTQUEUE_REG_2__5_ | ~new_P3_U5340;
  assign new_P3_U5357 = ~new_P3_U5332 | ~new_P3_U2441;
  assign new_P3_U5358 = ~new_P3_U2511 | ~new_P3_U2430;
  assign new_P3_U5359 = ~new_P3_U5331 | ~new_P3_U2429;
  assign new_P3_U5360 = ~new_P3_U2365 | ~new_P3_U2417;
  assign new_P3_U5361 = ~P3_INSTQUEUE_REG_2__4_ | ~new_P3_U5340;
  assign new_P3_U5362 = ~new_P3_U5332 | ~new_P3_U2440;
  assign new_P3_U5363 = ~new_P3_U2511 | ~new_P3_U2428;
  assign new_P3_U5364 = ~new_P3_U5331 | ~new_P3_U2427;
  assign new_P3_U5365 = ~new_P3_U2365 | ~new_P3_U2416;
  assign new_P3_U5366 = ~P3_INSTQUEUE_REG_2__3_ | ~new_P3_U5340;
  assign new_P3_U5367 = ~new_P3_U5332 | ~new_P3_U2439;
  assign new_P3_U5368 = ~new_P3_U2511 | ~new_P3_U2426;
  assign new_P3_U5369 = ~new_P3_U5331 | ~new_P3_U2425;
  assign new_P3_U5370 = ~new_P3_U2365 | ~new_P3_U2415;
  assign new_P3_U5371 = ~P3_INSTQUEUE_REG_2__2_ | ~new_P3_U5340;
  assign new_P3_U5372 = ~new_P3_U5332 | ~new_P3_U2438;
  assign new_P3_U5373 = ~new_P3_U2511 | ~new_P3_U2424;
  assign new_P3_U5374 = ~new_P3_U5331 | ~new_P3_U2423;
  assign new_P3_U5375 = ~new_P3_U2365 | ~new_P3_U2414;
  assign new_P3_U5376 = ~P3_INSTQUEUE_REG_2__1_ | ~new_P3_U5340;
  assign new_P3_U5377 = ~new_P3_U5332 | ~new_P3_U2437;
  assign new_P3_U5378 = ~new_P3_U2511 | ~new_P3_U2422;
  assign new_P3_U5379 = ~new_P3_U5331 | ~new_P3_U2421;
  assign new_P3_U5380 = ~new_P3_U2365 | ~new_P3_U2413;
  assign new_P3_U5381 = ~P3_INSTQUEUE_REG_2__0_ | ~new_P3_U5340;
  assign new_P3_U5382 = ~new_P3_U3203;
  assign new_P3_U5383 = ~new_P3_U3202;
  assign new_P3_U5384 = ~new_P3_U2460 | ~new_P3_U4343;
  assign new_P3_U5385 = ~new_P3_U3204;
  assign new_P3_U5386 = ~new_P3_U2509 | ~new_P3_U4645;
  assign new_P3_U5387 = ~new_P3_U3203 | ~new_P3_U5386;
  assign new_P3_U5388 = ~new_P3_U2489 | ~new_P3_U5387;
  assign new_P3_U5389 = ~new_P3_U5385 | ~new_P3_U5388;
  assign new_P3_U5390 = ~P3_STATE2_REG_3_ | ~new_P3_U3202;
  assign new_P3_U5391 = ~new_P3_U3617 | ~new_P3_U5389;
  assign new_P3_U5392 = ~new_P3_U2489 | ~new_P3_U3136;
  assign new_P3_U5393 = ~new_P3_U5383 | ~new_P3_U2445;
  assign new_P3_U5394 = ~new_P3_U2512 | ~new_P3_U2436;
  assign new_P3_U5395 = ~new_P3_U5382 | ~new_P3_U2435;
  assign new_P3_U5396 = ~new_P3_U2364 | ~new_P3_U2420;
  assign new_P3_U5397 = ~P3_INSTQUEUE_REG_1__7_ | ~new_P3_U5391;
  assign new_P3_U5398 = ~new_P3_U5383 | ~new_P3_U2443;
  assign new_P3_U5399 = ~new_P3_U2512 | ~new_P3_U2434;
  assign new_P3_U5400 = ~new_P3_U5382 | ~new_P3_U2433;
  assign new_P3_U5401 = ~new_P3_U2364 | ~new_P3_U2419;
  assign new_P3_U5402 = ~P3_INSTQUEUE_REG_1__6_ | ~new_P3_U5391;
  assign new_P3_U5403 = ~new_P3_U5383 | ~new_P3_U2442;
  assign new_P3_U5404 = ~new_P3_U2512 | ~new_P3_U2432;
  assign new_P3_U5405 = ~new_P3_U5382 | ~new_P3_U2431;
  assign new_P3_U5406 = ~new_P3_U2364 | ~new_P3_U2418;
  assign new_P3_U5407 = ~P3_INSTQUEUE_REG_1__5_ | ~new_P3_U5391;
  assign new_P3_U5408 = ~new_P3_U5383 | ~new_P3_U2441;
  assign new_P3_U5409 = ~new_P3_U2512 | ~new_P3_U2430;
  assign new_P3_U5410 = ~new_P3_U5382 | ~new_P3_U2429;
  assign new_P3_U5411 = ~new_P3_U2364 | ~new_P3_U2417;
  assign new_P3_U5412 = ~P3_INSTQUEUE_REG_1__4_ | ~new_P3_U5391;
  assign new_P3_U5413 = ~new_P3_U5383 | ~new_P3_U2440;
  assign new_P3_U5414 = ~new_P3_U2512 | ~new_P3_U2428;
  assign new_P3_U5415 = ~new_P3_U5382 | ~new_P3_U2427;
  assign new_P3_U5416 = ~new_P3_U2364 | ~new_P3_U2416;
  assign new_P3_U5417 = ~P3_INSTQUEUE_REG_1__3_ | ~new_P3_U5391;
  assign new_P3_U5418 = ~new_P3_U5383 | ~new_P3_U2439;
  assign new_P3_U5419 = ~new_P3_U2512 | ~new_P3_U2426;
  assign new_P3_U5420 = ~new_P3_U5382 | ~new_P3_U2425;
  assign new_P3_U5421 = ~new_P3_U2364 | ~new_P3_U2415;
  assign new_P3_U5422 = ~P3_INSTQUEUE_REG_1__2_ | ~new_P3_U5391;
  assign new_P3_U5423 = ~new_P3_U5383 | ~new_P3_U2438;
  assign new_P3_U5424 = ~new_P3_U2512 | ~new_P3_U2424;
  assign new_P3_U5425 = ~new_P3_U5382 | ~new_P3_U2423;
  assign new_P3_U5426 = ~new_P3_U2364 | ~new_P3_U2414;
  assign new_P3_U5427 = ~P3_INSTQUEUE_REG_1__1_ | ~new_P3_U5391;
  assign new_P3_U5428 = ~new_P3_U5383 | ~new_P3_U2437;
  assign new_P3_U5429 = ~new_P3_U2512 | ~new_P3_U2422;
  assign new_P3_U5430 = ~new_P3_U5382 | ~new_P3_U2421;
  assign new_P3_U5431 = ~new_P3_U2364 | ~new_P3_U2413;
  assign new_P3_U5432 = ~P3_INSTQUEUE_REG_1__0_ | ~new_P3_U5391;
  assign new_P3_U5433 = ~new_P3_U3206;
  assign new_P3_U5434 = ~new_P3_U3205;
  assign new_P3_U5435 = ~new_P3_U3073;
  assign new_P3_U5436 = ~new_P3_U2509 | ~new_P3_U2496;
  assign new_P3_U5437 = ~new_P3_U3206 | ~new_P3_U5436;
  assign new_P3_U5438 = ~new_P3_U2489 | ~new_P3_U5437;
  assign new_P3_U5439 = ~new_P3_U5438 | ~new_P3_U3073;
  assign new_P3_U5440 = ~P3_STATE2_REG_3_ | ~new_P3_U3205;
  assign new_P3_U5441 = ~new_P3_U3635 | ~new_P3_U5439;
  assign new_P3_U5442 = ~new_P3_U2489 | ~new_P3_U3136;
  assign new_P3_U5443 = ~new_P3_U5434 | ~new_P3_U2445;
  assign new_P3_U5444 = ~new_P3_U2513 | ~new_P3_U2436;
  assign new_P3_U5445 = ~new_P3_U5433 | ~new_P3_U2435;
  assign new_P3_U5446 = ~new_P3_U2363 | ~new_P3_U2420;
  assign new_P3_U5447 = ~P3_INSTQUEUE_REG_0__7_ | ~new_P3_U5441;
  assign new_P3_U5448 = ~new_P3_U5434 | ~new_P3_U2443;
  assign new_P3_U5449 = ~new_P3_U2513 | ~new_P3_U2434;
  assign new_P3_U5450 = ~new_P3_U5433 | ~new_P3_U2433;
  assign new_P3_U5451 = ~new_P3_U2363 | ~new_P3_U2419;
  assign new_P3_U5452 = ~P3_INSTQUEUE_REG_0__6_ | ~new_P3_U5441;
  assign new_P3_U5453 = ~new_P3_U5434 | ~new_P3_U2442;
  assign new_P3_U5454 = ~new_P3_U2513 | ~new_P3_U2432;
  assign new_P3_U5455 = ~new_P3_U5433 | ~new_P3_U2431;
  assign new_P3_U5456 = ~new_P3_U2363 | ~new_P3_U2418;
  assign new_P3_U5457 = ~P3_INSTQUEUE_REG_0__5_ | ~new_P3_U5441;
  assign new_P3_U5458 = ~new_P3_U5434 | ~new_P3_U2441;
  assign new_P3_U5459 = ~new_P3_U2513 | ~new_P3_U2430;
  assign new_P3_U5460 = ~new_P3_U5433 | ~new_P3_U2429;
  assign new_P3_U5461 = ~new_P3_U2363 | ~new_P3_U2417;
  assign new_P3_U5462 = ~P3_INSTQUEUE_REG_0__4_ | ~new_P3_U5441;
  assign new_P3_U5463 = ~new_P3_U5434 | ~new_P3_U2440;
  assign new_P3_U5464 = ~new_P3_U2513 | ~new_P3_U2428;
  assign new_P3_U5465 = ~new_P3_U5433 | ~new_P3_U2427;
  assign new_P3_U5466 = ~new_P3_U2363 | ~new_P3_U2416;
  assign new_P3_U5467 = ~P3_INSTQUEUE_REG_0__3_ | ~new_P3_U5441;
  assign new_P3_U5468 = ~new_P3_U5434 | ~new_P3_U2439;
  assign new_P3_U5469 = ~new_P3_U2513 | ~new_P3_U2426;
  assign new_P3_U5470 = ~new_P3_U5433 | ~new_P3_U2425;
  assign new_P3_U5471 = ~new_P3_U2363 | ~new_P3_U2415;
  assign new_P3_U5472 = ~P3_INSTQUEUE_REG_0__2_ | ~new_P3_U5441;
  assign new_P3_U5473 = ~new_P3_U5434 | ~new_P3_U2438;
  assign new_P3_U5474 = ~new_P3_U2513 | ~new_P3_U2424;
  assign new_P3_U5475 = ~new_P3_U5433 | ~new_P3_U2423;
  assign new_P3_U5476 = ~new_P3_U2363 | ~new_P3_U2414;
  assign new_P3_U5477 = ~P3_INSTQUEUE_REG_0__1_ | ~new_P3_U5441;
  assign new_P3_U5478 = ~new_P3_U5434 | ~new_P3_U2437;
  assign new_P3_U5479 = ~new_P3_U2513 | ~new_P3_U2422;
  assign new_P3_U5480 = ~new_P3_U5433 | ~new_P3_U2421;
  assign new_P3_U5481 = ~new_P3_U2363 | ~new_P3_U2413;
  assign new_P3_U5482 = ~P3_INSTQUEUE_REG_0__0_ | ~new_P3_U5441;
  assign new_P3_U5483 = ~new_P3_U4339 | ~new_P3_U3655 | ~new_P3_U7917 | ~new_P3_U2514;
  assign new_P3_U5484 = ~new_P3_U3209;
  assign new_P3_U5485 = ~new_P3_U4296 | ~new_P3_U3209;
  assign new_P3_U5486 = ~new_P3_GTE_450_U6 | ~new_P3_U4303;
  assign new_P3_U5487 = ~new_P3_GTE_504_U6 | ~new_P3_U4302;
  assign new_P3_U5488 = ~new_P3_U3255;
  assign new_P3_U5489 = ~new_P3_GTE_412_U6 | ~new_P3_U4304;
  assign new_P3_U5490 = ~new_P3_GTE_485_U6 | ~new_P3_U2356;
  assign new_P3_U5491 = ~new_P3_U3254;
  assign new_P3_U5492 = ~new_P3_U3254 | ~new_P3_U2630;
  assign new_P3_U5493 = ~new_P3_GTE_390_U6 | ~new_P3_U2357;
  assign new_P3_U5494 = ~new_P3_U4294 | ~new_P3_U3255;
  assign new_P3_U5495 = ~new_P3_GTE_401_U6 | ~new_P3_U4305;
  assign new_P3_U5496 = ~new_P3_U4290;
  assign new_P3_U5497 = ~new_P3_U2390 | ~new_P3_U4290;
  assign new_P3_U5498 = ~P3_STATE2_REG_3_ | ~new_P3_U3121;
  assign new_P3_U5499 = ~new_P3_U4283;
  assign new_P3_U5500 = ~new_P3_U3095 | ~new_P3_U3097;
  assign new_P3_U5501 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_U5500;
  assign new_P3_U5502 = ~new_P3_U2481 | ~new_P3_U3095;
  assign new_P3_U5503 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_U5504 = ~new_P3_U3223;
  assign new_P3_U5505 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U4332;
  assign new_P3_U5506 = ~new_P3_U3224;
  assign new_P3_U5507 = ~new_P3_U5484 | ~new_P3_U3107;
  assign new_P3_U5508 = ~new_P3_U4488 | ~new_P3_U4522 | ~new_P3_U4607;
  assign new_P3_U5509 = ~new_P3_U4296 | ~new_P3_U5507;
  assign new_P3_U5510 = ~new_P3_U3104 | ~new_P3_U7974 | ~new_P3_U7973;
  assign new_P3_U5511 = ~new_P3_U4323 | ~new_P3_U4344;
  assign new_P3_U5512 = ~new_P3_U5509 | ~new_P3_U3665;
  assign new_P3_U5513 = ~new_P3_U4522 | ~new_P3_U4607;
  assign new_P3_U5514 = ~new_P3_U4607 | ~new_P3_U3218;
  assign new_P3_U5515 = ~new_P3_U4556 | ~new_P3_U5514 | ~new_P3_U3216;
  assign new_P3_U5516 = ~new_P3_U4573 | ~new_P3_U4505;
  assign new_P3_U5517 = ~new_P3_U4488 | ~new_P3_U5516;
  assign new_P3_U5518 = ~new_P3_U3112 | ~new_P3_U3103 | ~new_P3_U3218;
  assign new_P3_U5519 = ~new_P3_U4573 | ~new_P3_U4607 | ~new_P3_U3104;
  assign new_P3_U5520 = ~new_P3_U4324 | ~new_P3_U3103;
  assign new_P3_U5521 = ~new_P3_U5518 | ~new_P3_U3102;
  assign new_P3_U5522 = ~new_P3_U3220;
  assign new_P3_U5523 = ~new_P3_U3111 | ~new_P3_U3114;
  assign new_P3_U5524 = ~new_P3_U2452 | ~new_P3_U3108;
  assign new_P3_U5525 = ~new_P3_U3221;
  assign new_P3_U5526 = ~new_P3_U2462 | ~new_P3_U3104;
  assign new_P3_U5527 = ~new_P3_U3229 | ~new_P3_U3219;
  assign new_P3_U5528 = ~new_P3_U2456 | ~new_P3_U5527;
  assign new_P3_U5529 = ~new_P3_U2518 | ~new_P3_U3217;
  assign new_P3_U5530 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_U5529;
  assign new_P3_U5531 = ~new_P3_U5525 | ~new_P3_U5530;
  assign new_P3_U5532 = ~new_P3_U2450 | ~new_P3_U2461 | ~new_P3_U5523;
  assign new_P3_U5533 = ~new_P3_U3673 | ~new_P3_U7918;
  assign new_P3_U5534 = ~new_P3_U3226;
  assign new_P3_U5535 = ~new_P3_U3672 | ~new_P3_U5522;
  assign new_P3_U5536 = ~new_P3_U2451 | ~new_P3_U3659 | ~new_P3_U5523;
  assign new_P3_U5537 = ~new_P3_U3669 | ~new_P3_U5531;
  assign new_P3_U5538 = ~new_P3_U3670 | ~new_P3_U3220;
  assign new_P3_U5539 = ~new_P3_U5504 | ~new_P3_U5535;
  assign new_P3_U5540 = ~new_P3_U5506 | ~new_P3_U3226;
  assign new_P3_U5541 = ~new_P3_ADD_495_U9 | ~new_P3_U2356;
  assign new_P3_U5542 = ~new_P3_U5537 | ~new_P3_U3676;
  assign new_P3_U5543 = ~new_P3_U3265;
  assign new_P3_U5544 = ~new_P3_U4345 | ~new_P3_U3265;
  assign new_P3_U5545 = ~new_P3_U4340 | ~new_P3_U5542;
  assign new_P3_U5546 = ~new_P3_U5545 | ~new_P3_U5544;
  assign new_P3_U5547 = ~new_P3_U3227;
  assign new_P3_U5548 = ~new_P3_U3225;
  assign new_P3_U5549 = ~new_P3_U5534 | ~new_P3_U5522;
  assign new_P3_U5550 = ~new_P3_U2451 | ~new_P3_U5548 | ~new_P3_U5523;
  assign new_P3_U5551 = ~new_P3_U5547 | ~new_P3_U5549;
  assign new_P3_U5552 = ~new_P3_ADD_495_U10 | ~new_P3_U2356;
  assign new_P3_U5553 = ~new_P3_U3679 | ~new_P3_U7982 | ~new_P3_U7981;
  assign new_P3_U5554 = ~new_P3_U3287 | ~P3_STATE2_REG_1_ | ~new_P3_U3286;
  assign new_P3_U5555 = ~new_P3_U4345 | ~new_P3_U3225;
  assign new_P3_U5556 = ~new_P3_U4340 | ~new_P3_U5553;
  assign new_P3_U5557 = ~new_P3_U3680 | ~new_P3_U5556;
  assign new_P3_U5558 = ~new_P3_U3228;
  assign new_P3_U5559 = ~new_P3_U4341 | ~new_P3_U4608;
  assign new_P3_U5560 = ~new_P3_U3231;
  assign new_P3_U5561 = ~new_P3_U3230;
  assign new_P3_U5562 = ~new_P3_U2466 | ~new_P3_U3230;
  assign new_P3_U5563 = ~new_P3_U5531 | ~new_P3_U3094;
  assign new_P3_U5564 = ~new_P3_U5558 | ~new_P3_U3231;
  assign new_P3_U5565 = ~new_P3_ADD_495_U4 | ~new_P3_U2356;
  assign new_P3_U5566 = ~new_P3_U5563 | ~new_P3_U3681;
  assign new_P3_U5567 = ~new_P3_U7985 | ~P3_STATE2_REG_1_ | ~new_P3_U3286;
  assign new_P3_U5568 = ~new_P3_U5558 | ~new_P3_U4345;
  assign new_P3_U5569 = ~new_P3_U4340 | ~new_P3_U5566;
  assign new_P3_U5570 = ~new_P3_U3683 | ~new_P3_U5569;
  assign new_P3_U5571 = ~new_P3_U5560 | ~new_P3_U5561;
  assign new_P3_U5572 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_U2356;
  assign new_P3_U5573 = ~new_P3_U5572 | ~new_P3_U7994 | ~new_P3_U7993;
  assign new_P3_U5574 = ~new_P3_U4345 | ~new_P3_U3093;
  assign new_P3_U5575 = ~new_P3_U4340 | ~new_P3_U5573;
  assign new_P3_U5576 = ~new_P3_U7988 | ~P3_STATE2_REG_1_;
  assign new_P3_U5577 = ~new_P3_U3684 | ~new_P3_U5575;
  assign new_P3_U5578 = ~new_P3_LT_589_U6 | ~new_P3_U2453 | ~P3_STATE2_REG_0_;
  assign new_P3_U5579 = ~new_P3_U3233;
  assign new_P3_U5580 = ~P3_STATE2_REG_3_ | ~new_P3_U3132;
  assign new_P3_U5581 = ~new_P3_U3233 | ~new_P3_U5580;
  assign new_P3_U5582 = ~new_P3_U4315 | ~new_P3_U3123;
  assign new_P3_U5583 = ~new_P3_U4647 | ~new_P3_U3271;
  assign new_P3_U5584 = ~new_P3_U3182 | ~new_P3_U5583;
  assign new_P3_U5585 = ~new_P3_U3183 | ~new_P3_U5584;
  assign new_P3_U5586 = ~new_P3_U4322 | ~new_P3_U5585;
  assign new_P3_U5587 = ~new_P3_U5582 | ~new_P3_U3142;
  assign new_P3_U5588 = ~new_P3_U4650 | ~P3_STATE2_REG_3_;
  assign new_P3_U5589 = ~new_P3_U3685 | ~new_P3_U5586;
  assign new_P3_U5590 = ~new_P3_U5589 | ~new_P3_U3233;
  assign new_P3_U5591 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_U5581;
  assign new_P3_U5592 = ~new_P3_U4648 | ~P3_STATE2_REG_3_ | ~new_P3_U3131;
  assign new_P3_U5593 = ~new_P3_U4322 | ~new_P3_U7999;
  assign new_P3_U5594 = ~new_P3_U3270 | ~new_P3_U5582;
  assign new_P3_U5595 = ~new_P3_U3686 | ~new_P3_U5593;
  assign new_P3_U5596 = ~P3_STATE2_REG_3_ | ~new_P3_U3130;
  assign new_P3_U5597 = ~new_P3_U3233 | ~new_P3_U5596;
  assign new_P3_U5598 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_U5597;
  assign new_P3_U5599 = ~new_P3_U5595 | ~new_P3_U3233;
  assign new_P3_U5600 = ~new_P3_U4322 | ~new_P3_U3156;
  assign new_P3_U5601 = ~P3_STATE2_REG_3_ | ~new_P3_U3129;
  assign new_P3_U5602 = ~new_P3_U5601 | ~new_P3_U5600;
  assign new_P3_U5603 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_U5602;
  assign new_P3_U5604 = ~new_P3_U2493 | ~new_P3_U4322;
  assign new_P3_U5605 = ~new_P3_U5582 | ~new_P3_U3141;
  assign new_P3_U5606 = ~new_P3_U5604 | ~new_P3_U5605 | ~new_P3_U5603;
  assign new_P3_U5607 = ~P3_STATE2_REG_3_ | ~new_P3_U3128;
  assign new_P3_U5608 = ~new_P3_U3233 | ~new_P3_U5607;
  assign new_P3_U5609 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_U5608;
  assign new_P3_U5610 = ~new_P3_U5606 | ~new_P3_U3233;
  assign new_P3_U5611 = ~new_P3_U3234;
  assign new_P3_U5612 = ~new_P3_U5611 | ~new_P3_U3233;
  assign new_P3_U5613 = ~P3_STATE2_REG_3_ | ~new_P3_U3128;
  assign new_P3_U5614 = ~new_P3_U4337 | ~new_P3_U5613;
  assign new_P3_U5615 = ~new_P3_U5614 | ~new_P3_U3233;
  assign new_P3_U5616 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_U5612;
  assign new_P3_U5617 = ~new_P3_GTE_450_U6 | ~new_P3_U2463 | ~new_P3_U4294;
  assign new_P3_U5618 = ~new_P3_GTE_370_U6 | ~new_P3_U4344;
  assign new_P3_U5619 = ~new_P3_U5618 | ~new_P3_U5617;
  assign new_P3_U5620 = ~new_P3_GTE_412_U6 | ~new_P3_U4590 | ~new_P3_U2630;
  assign new_P3_U5621 = ~new_P3_GTE_355_U6 | ~new_P3_U3074;
  assign new_P3_U5622 = ~new_P3_U5621 | ~new_P3_U5620;
  assign new_P3_U5623 = ~new_P3_GTE_390_U6 | ~new_P3_U4488;
  assign new_P3_U5624 = ~new_P3_U5623 | ~new_P3_U8001 | ~new_P3_U8000;
  assign new_P3_U5625 = ~new_P3_GTE_401_U6 | ~new_P3_U3102 | ~new_P3_U3108;
  assign new_P3_U5626 = ~new_P3_U4349 | ~new_P3_GTE_504_U6;
  assign new_P3_U5627 = ~new_P3_U4348 | ~new_P3_GTE_485_U6;
  assign new_P3_U5628 = ~new_P3_U4539 | ~new_P3_U5624;
  assign new_P3_U5629 = ~new_P3_U5628 | ~new_P3_U3687 | ~new_P3_U2515 | ~new_P3_U5627;
  assign new_P3_U5630 = ~new_P3_U2390 | ~new_P3_U5629;
  assign new_P3_U5631 = ~new_P3_U3248;
  assign new_P3_U5632 = ~new_P3_ADD_360_1242_U85 | ~new_P3_U2395;
  assign new_P3_U5633 = ~new_P3_SUB_357_1258_U69 | ~new_P3_U2393;
  assign new_P3_U5634 = ~new_P3_ADD_558_U5 | ~new_P3_U3220;
  assign new_P3_U5635 = ~new_P3_U4298 | ~new_P3_ADD_553_U5;
  assign new_P3_U5636 = ~new_P3_U4299 | ~new_P3_ADD_547_U5;
  assign new_P3_U5637 = ~new_P3_U4300 | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_U5638 = ~new_P3_U4301 | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_U5639 = ~new_P3_U2354 | ~new_P3_ADD_531_U5;
  assign new_P3_U5640 = ~new_P3_U2355 | ~new_P3_ADD_526_U5;
  assign new_P3_U5641 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_U4302;
  assign new_P3_U5642 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_U2356;
  assign new_P3_U5643 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_U4303;
  assign new_P3_U5644 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_U4304;
  assign new_P3_U5645 = ~new_P3_ADD_405_U4 | ~new_P3_U4305;
  assign new_P3_U5646 = ~new_P3_ADD_394_U4 | ~new_P3_U2357;
  assign new_P3_U5647 = ~new_P3_U2358 | ~new_P3_ADD_385_U5;
  assign new_P3_U5648 = ~new_P3_U2359 | ~new_P3_ADD_380_U5;
  assign new_P3_U5649 = ~new_P3_U4306 | ~new_P3_ADD_349_U5;
  assign new_P3_U5650 = ~new_P3_U2362 | ~new_P3_ADD_344_U5;
  assign new_P3_U5651 = ~new_P3_ADD_371_1212_U87 | ~new_P3_U2360;
  assign new_P3_U5652 = ~new_P3_U3698 | ~new_P3_U3693 | ~new_P3_U3692 | ~new_P3_U5634;
  assign new_P3_U5653 = ~P3_REIP_REG_0_ | ~new_P3_U2402;
  assign new_P3_U5654 = ~new_P3_U4318 | ~new_P3_U5652;
  assign new_P3_U5655 = ~new_P3_U5631 | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_U5656 = ~new_P3_ADD_360_1242_U19 | ~new_P3_U2395;
  assign new_P3_U5657 = ~new_P3_SUB_357_1258_U21 | ~new_P3_U2393;
  assign new_P3_U5658 = ~new_P3_ADD_558_U85 | ~new_P3_U3220;
  assign new_P3_U5659 = ~new_P3_ADD_553_U85 | ~new_P3_U4298;
  assign new_P3_U5660 = ~new_P3_ADD_547_U85 | ~new_P3_U4299;
  assign new_P3_U5661 = ~new_P3_ADD_541_U4 | ~new_P3_U4300;
  assign new_P3_U5662 = ~new_P3_ADD_536_U4 | ~new_P3_U4301;
  assign new_P3_U5663 = ~new_P3_ADD_531_U85 | ~new_P3_U2354;
  assign new_P3_U5664 = ~new_P3_ADD_526_U71 | ~new_P3_U2355;
  assign new_P3_U5665 = ~new_P3_ADD_515_U4 | ~new_P3_U4302;
  assign new_P3_U5666 = ~new_P3_ADD_494_U4 | ~new_P3_U2356;
  assign new_P3_U5667 = ~new_P3_ADD_476_U4 | ~new_P3_U4303;
  assign new_P3_U5668 = ~new_P3_ADD_441_U4 | ~new_P3_U4304;
  assign new_P3_U5669 = ~new_P3_ADD_405_U81 | ~new_P3_U4305;
  assign new_P3_U5670 = ~new_P3_ADD_394_U81 | ~new_P3_U2357;
  assign new_P3_U5671 = ~new_P3_ADD_385_U85 | ~new_P3_U2358;
  assign new_P3_U5672 = ~new_P3_ADD_380_U85 | ~new_P3_U2359;
  assign new_P3_U5673 = ~new_P3_ADD_349_U85 | ~new_P3_U4306;
  assign new_P3_U5674 = ~new_P3_ADD_344_U85 | ~new_P3_U2362;
  assign new_P3_U5675 = ~new_P3_ADD_371_1212_U20 | ~new_P3_U2360;
  assign new_P3_U5676 = ~new_P3_U3700 | ~new_P3_U3705 | ~new_P3_U5656 | ~new_P3_U5658 | ~new_P3_U3699;
  assign new_P3_U5677 = ~new_P3_U2402 | ~P3_REIP_REG_1_;
  assign new_P3_U5678 = ~new_P3_U4318 | ~new_P3_U5676;
  assign new_P3_U5679 = ~new_P3_U5631 | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_U5680 = ~new_P3_ADD_360_1242_U91 | ~new_P3_U2395;
  assign new_P3_U5681 = ~new_P3_SUB_357_1258_U78 | ~new_P3_U2393;
  assign new_P3_U5682 = ~new_P3_ADD_558_U74 | ~new_P3_U3220;
  assign new_P3_U5683 = ~new_P3_ADD_553_U74 | ~new_P3_U4298;
  assign new_P3_U5684 = ~new_P3_ADD_547_U74 | ~new_P3_U4299;
  assign new_P3_U5685 = ~new_P3_ADD_541_U71 | ~new_P3_U4300;
  assign new_P3_U5686 = ~new_P3_ADD_536_U71 | ~new_P3_U4301;
  assign new_P3_U5687 = ~new_P3_ADD_531_U74 | ~new_P3_U2354;
  assign new_P3_U5688 = ~new_P3_ADD_526_U60 | ~new_P3_U2355;
  assign new_P3_U5689 = ~new_P3_ADD_515_U71 | ~new_P3_U4302;
  assign new_P3_U5690 = ~new_P3_ADD_494_U71 | ~new_P3_U2356;
  assign new_P3_U5691 = ~new_P3_ADD_476_U71 | ~new_P3_U4303;
  assign new_P3_U5692 = ~new_P3_ADD_441_U71 | ~new_P3_U4304;
  assign new_P3_U5693 = ~new_P3_ADD_405_U5 | ~new_P3_U4305;
  assign new_P3_U5694 = ~new_P3_ADD_394_U5 | ~new_P3_U2357;
  assign new_P3_U5695 = ~new_P3_ADD_385_U74 | ~new_P3_U2358;
  assign new_P3_U5696 = ~new_P3_ADD_380_U74 | ~new_P3_U2359;
  assign new_P3_U5697 = ~new_P3_ADD_349_U74 | ~new_P3_U4306;
  assign new_P3_U5698 = ~new_P3_ADD_344_U74 | ~new_P3_U2362;
  assign new_P3_U5699 = ~new_P3_ADD_371_1212_U93 | ~new_P3_U2360;
  assign new_P3_U5700 = ~new_P3_U3713 | ~new_P3_U3706 | ~new_P3_U5680 | ~new_P3_U5682 | ~new_P3_U3710;
  assign new_P3_U5701 = ~new_P3_U2402 | ~P3_REIP_REG_2_;
  assign new_P3_U5702 = ~new_P3_U4318 | ~new_P3_U5700;
  assign new_P3_U5703 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_U5631;
  assign new_P3_U5704 = ~new_P3_ADD_360_1242_U17 | ~new_P3_U2395;
  assign new_P3_U5705 = ~new_P3_SUB_357_1258_U76 | ~new_P3_U2393;
  assign new_P3_U5706 = ~new_P3_ADD_558_U71 | ~new_P3_U3220;
  assign new_P3_U5707 = ~new_P3_ADD_553_U71 | ~new_P3_U4298;
  assign new_P3_U5708 = ~new_P3_ADD_547_U71 | ~new_P3_U4299;
  assign new_P3_U5709 = ~new_P3_ADD_541_U68 | ~new_P3_U4300;
  assign new_P3_U5710 = ~new_P3_ADD_536_U68 | ~new_P3_U4301;
  assign new_P3_U5711 = ~new_P3_ADD_531_U71 | ~new_P3_U2354;
  assign new_P3_U5712 = ~new_P3_ADD_526_U57 | ~new_P3_U2355;
  assign new_P3_U5713 = ~new_P3_ADD_515_U68 | ~new_P3_U4302;
  assign new_P3_U5714 = ~new_P3_ADD_494_U68 | ~new_P3_U2356;
  assign new_P3_U5715 = ~new_P3_ADD_476_U68 | ~new_P3_U4303;
  assign new_P3_U5716 = ~new_P3_ADD_441_U68 | ~new_P3_U4304;
  assign new_P3_U5717 = ~new_P3_ADD_405_U93 | ~new_P3_U4305;
  assign new_P3_U5718 = ~new_P3_ADD_394_U93 | ~new_P3_U2357;
  assign new_P3_U5719 = ~new_P3_ADD_385_U71 | ~new_P3_U2358;
  assign new_P3_U5720 = ~new_P3_ADD_380_U71 | ~new_P3_U2359;
  assign new_P3_U5721 = ~new_P3_ADD_349_U71 | ~new_P3_U4306;
  assign new_P3_U5722 = ~new_P3_ADD_344_U71 | ~new_P3_U2362;
  assign new_P3_U5723 = ~new_P3_ADD_371_1212_U18 | ~new_P3_U2360;
  assign new_P3_U5724 = ~new_P3_U3721 | ~new_P3_U3714 | ~new_P3_U3718 | ~new_P3_U3715 | ~new_P3_U5706;
  assign new_P3_U5725 = ~new_P3_U2402 | ~P3_REIP_REG_3_;
  assign new_P3_U5726 = ~new_P3_U4318 | ~new_P3_U5724;
  assign new_P3_U5727 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_U5631;
  assign new_P3_U5728 = ~new_P3_ADD_360_1242_U18 | ~new_P3_U2395;
  assign new_P3_U5729 = ~new_P3_SUB_357_1258_U75 | ~new_P3_U2393;
  assign new_P3_U5730 = ~new_P3_ADD_558_U70 | ~new_P3_U3220;
  assign new_P3_U5731 = ~new_P3_ADD_553_U70 | ~new_P3_U4298;
  assign new_P3_U5732 = ~new_P3_ADD_547_U70 | ~new_P3_U4299;
  assign new_P3_U5733 = ~new_P3_ADD_541_U67 | ~new_P3_U4300;
  assign new_P3_U5734 = ~new_P3_ADD_536_U67 | ~new_P3_U4301;
  assign new_P3_U5735 = ~new_P3_ADD_531_U70 | ~new_P3_U2354;
  assign new_P3_U5736 = ~new_P3_ADD_526_U56 | ~new_P3_U2355;
  assign new_P3_U5737 = ~new_P3_ADD_515_U67 | ~new_P3_U4302;
  assign new_P3_U5738 = ~new_P3_ADD_494_U67 | ~new_P3_U2356;
  assign new_P3_U5739 = ~new_P3_ADD_476_U67 | ~new_P3_U4303;
  assign new_P3_U5740 = ~new_P3_ADD_441_U67 | ~new_P3_U4304;
  assign new_P3_U5741 = ~new_P3_ADD_405_U68 | ~new_P3_U4305;
  assign new_P3_U5742 = ~new_P3_ADD_394_U68 | ~new_P3_U2357;
  assign new_P3_U5743 = ~new_P3_ADD_385_U70 | ~new_P3_U2358;
  assign new_P3_U5744 = ~new_P3_ADD_380_U70 | ~new_P3_U2359;
  assign new_P3_U5745 = ~new_P3_ADD_349_U70 | ~new_P3_U4306;
  assign new_P3_U5746 = ~new_P3_ADD_344_U70 | ~new_P3_U2362;
  assign new_P3_U5747 = ~new_P3_ADD_371_1212_U91 | ~new_P3_U2360;
  assign new_P3_U5748 = ~new_P3_U3729 | ~new_P3_U3722 | ~new_P3_U5728 | ~new_P3_U5730 | ~new_P3_U3726;
  assign new_P3_U5749 = ~new_P3_U2402 | ~P3_REIP_REG_4_;
  assign new_P3_U5750 = ~new_P3_U4318 | ~new_P3_U5748;
  assign new_P3_U5751 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_U5631;
  assign new_P3_U5752 = ~new_P3_ADD_360_1242_U89 | ~new_P3_U2395;
  assign new_P3_U5753 = ~new_P3_SUB_357_1258_U74 | ~new_P3_U2393;
  assign new_P3_U5754 = ~new_P3_ADD_558_U69 | ~new_P3_U3220;
  assign new_P3_U5755 = ~new_P3_ADD_553_U69 | ~new_P3_U4298;
  assign new_P3_U5756 = ~new_P3_ADD_547_U69 | ~new_P3_U4299;
  assign new_P3_U5757 = ~new_P3_ADD_541_U66 | ~new_P3_U4300;
  assign new_P3_U5758 = ~new_P3_ADD_536_U66 | ~new_P3_U4301;
  assign new_P3_U5759 = ~new_P3_ADD_531_U69 | ~new_P3_U2354;
  assign new_P3_U5760 = ~new_P3_ADD_526_U55 | ~new_P3_U2355;
  assign new_P3_U5761 = ~new_P3_ADD_515_U66 | ~new_P3_U4302;
  assign new_P3_U5762 = ~new_P3_ADD_494_U66 | ~new_P3_U2356;
  assign new_P3_U5763 = ~new_P3_ADD_476_U66 | ~new_P3_U4303;
  assign new_P3_U5764 = ~new_P3_ADD_441_U66 | ~new_P3_U4304;
  assign new_P3_U5765 = ~new_P3_ADD_405_U67 | ~new_P3_U4305;
  assign new_P3_U5766 = ~new_P3_ADD_394_U67 | ~new_P3_U2357;
  assign new_P3_U5767 = ~new_P3_ADD_385_U69 | ~new_P3_U2358;
  assign new_P3_U5768 = ~new_P3_ADD_380_U69 | ~new_P3_U2359;
  assign new_P3_U5769 = ~new_P3_ADD_349_U69 | ~new_P3_U4306;
  assign new_P3_U5770 = ~new_P3_ADD_344_U69 | ~new_P3_U2362;
  assign new_P3_U5771 = ~new_P3_ADD_371_1212_U19 | ~new_P3_U2360;
  assign new_P3_U5772 = ~new_P3_U3737 | ~new_P3_U3730 | ~new_P3_U5753 | ~new_P3_U3734 | ~new_P3_U5754;
  assign new_P3_U5773 = ~new_P3_U2402 | ~P3_REIP_REG_5_;
  assign new_P3_U5774 = ~new_P3_U4318 | ~new_P3_U5772;
  assign new_P3_U5775 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_U5631;
  assign new_P3_U5776 = ~new_P3_ADD_360_1242_U88 | ~new_P3_U2395;
  assign new_P3_U5777 = ~new_P3_SUB_357_1258_U73 | ~new_P3_U2393;
  assign new_P3_U5778 = ~new_P3_ADD_558_U68 | ~new_P3_U3220;
  assign new_P3_U5779 = ~new_P3_ADD_553_U68 | ~new_P3_U4298;
  assign new_P3_U5780 = ~new_P3_ADD_547_U68 | ~new_P3_U4299;
  assign new_P3_U5781 = ~new_P3_ADD_541_U65 | ~new_P3_U4300;
  assign new_P3_U5782 = ~new_P3_ADD_536_U65 | ~new_P3_U4301;
  assign new_P3_U5783 = ~new_P3_ADD_531_U68 | ~new_P3_U2354;
  assign new_P3_U5784 = ~new_P3_ADD_526_U54 | ~new_P3_U2355;
  assign new_P3_U5785 = ~new_P3_ADD_515_U65 | ~new_P3_U4302;
  assign new_P3_U5786 = ~new_P3_ADD_494_U65 | ~new_P3_U2356;
  assign new_P3_U5787 = ~new_P3_ADD_476_U65 | ~new_P3_U4303;
  assign new_P3_U5788 = ~new_P3_ADD_441_U65 | ~new_P3_U4304;
  assign new_P3_U5789 = ~new_P3_ADD_405_U66 | ~new_P3_U4305;
  assign new_P3_U5790 = ~new_P3_ADD_394_U66 | ~new_P3_U2357;
  assign new_P3_U5791 = ~new_P3_ADD_385_U68 | ~new_P3_U2358;
  assign new_P3_U5792 = ~new_P3_ADD_380_U68 | ~new_P3_U2359;
  assign new_P3_U5793 = ~new_P3_ADD_349_U68 | ~new_P3_U4306;
  assign new_P3_U5794 = ~new_P3_ADD_344_U68 | ~new_P3_U2362;
  assign new_P3_U5795 = ~new_P3_ADD_371_1212_U90 | ~new_P3_U2360;
  assign new_P3_U5796 = ~new_P3_U3745 | ~new_P3_U3738 | ~new_P3_U5777 | ~new_P3_U3742 | ~new_P3_U5778;
  assign new_P3_U5797 = ~new_P3_U2402 | ~P3_REIP_REG_6_;
  assign new_P3_U5798 = ~new_P3_U4318 | ~new_P3_U5796;
  assign new_P3_U5799 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_U5631;
  assign new_P3_U5800 = ~new_P3_ADD_360_1242_U87 | ~new_P3_U2395;
  assign new_P3_U5801 = ~new_P3_SUB_357_1258_U72 | ~new_P3_U2393;
  assign new_P3_U5802 = ~new_P3_ADD_558_U67 | ~new_P3_U3220;
  assign new_P3_U5803 = ~new_P3_ADD_553_U67 | ~new_P3_U4298;
  assign new_P3_U5804 = ~new_P3_ADD_547_U67 | ~new_P3_U4299;
  assign new_P3_U5805 = ~new_P3_ADD_541_U64 | ~new_P3_U4300;
  assign new_P3_U5806 = ~new_P3_ADD_536_U64 | ~new_P3_U4301;
  assign new_P3_U5807 = ~new_P3_ADD_531_U67 | ~new_P3_U2354;
  assign new_P3_U5808 = ~new_P3_ADD_526_U53 | ~new_P3_U2355;
  assign new_P3_U5809 = ~new_P3_ADD_515_U64 | ~new_P3_U4302;
  assign new_P3_U5810 = ~new_P3_ADD_494_U64 | ~new_P3_U2356;
  assign new_P3_U5811 = ~new_P3_ADD_476_U64 | ~new_P3_U4303;
  assign new_P3_U5812 = ~new_P3_ADD_441_U64 | ~new_P3_U4304;
  assign new_P3_U5813 = ~new_P3_ADD_405_U65 | ~new_P3_U4305;
  assign new_P3_U5814 = ~new_P3_ADD_394_U65 | ~new_P3_U2357;
  assign new_P3_U5815 = ~new_P3_ADD_385_U67 | ~new_P3_U2358;
  assign new_P3_U5816 = ~new_P3_ADD_380_U67 | ~new_P3_U2359;
  assign new_P3_U5817 = ~new_P3_ADD_349_U67 | ~new_P3_U4306;
  assign new_P3_U5818 = ~new_P3_ADD_344_U67 | ~new_P3_U2362;
  assign new_P3_U5819 = ~new_P3_ADD_371_1212_U89 | ~new_P3_U2360;
  assign new_P3_U5820 = ~new_P3_U3753 | ~new_P3_U3746 | ~new_P3_U5801 | ~new_P3_U3750 | ~new_P3_U5802;
  assign new_P3_U5821 = ~new_P3_U2402 | ~P3_REIP_REG_7_;
  assign new_P3_U5822 = ~new_P3_U4318 | ~new_P3_U5820;
  assign new_P3_U5823 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_U5631;
  assign new_P3_U5824 = ~new_P3_ADD_360_1242_U86 | ~new_P3_U2395;
  assign new_P3_U5825 = ~new_P3_SUB_357_1258_U71 | ~new_P3_U2393;
  assign new_P3_U5826 = ~new_P3_ADD_558_U66 | ~new_P3_U3220;
  assign new_P3_U5827 = ~new_P3_ADD_553_U66 | ~new_P3_U4298;
  assign new_P3_U5828 = ~new_P3_ADD_547_U66 | ~new_P3_U4299;
  assign new_P3_U5829 = ~new_P3_ADD_541_U63 | ~new_P3_U4300;
  assign new_P3_U5830 = ~new_P3_ADD_536_U63 | ~new_P3_U4301;
  assign new_P3_U5831 = ~new_P3_ADD_531_U66 | ~new_P3_U2354;
  assign new_P3_U5832 = ~new_P3_ADD_526_U52 | ~new_P3_U2355;
  assign new_P3_U5833 = ~new_P3_ADD_515_U63 | ~new_P3_U4302;
  assign new_P3_U5834 = ~new_P3_ADD_494_U63 | ~new_P3_U2356;
  assign new_P3_U5835 = ~new_P3_ADD_476_U63 | ~new_P3_U4303;
  assign new_P3_U5836 = ~new_P3_ADD_441_U63 | ~new_P3_U4304;
  assign new_P3_U5837 = ~new_P3_ADD_405_U64 | ~new_P3_U4305;
  assign new_P3_U5838 = ~new_P3_ADD_394_U64 | ~new_P3_U2357;
  assign new_P3_U5839 = ~new_P3_ADD_385_U66 | ~new_P3_U2358;
  assign new_P3_U5840 = ~new_P3_ADD_380_U66 | ~new_P3_U2359;
  assign new_P3_U5841 = ~new_P3_ADD_349_U66 | ~new_P3_U4306;
  assign new_P3_U5842 = ~new_P3_ADD_344_U66 | ~new_P3_U2362;
  assign new_P3_U5843 = ~new_P3_ADD_371_1212_U88 | ~new_P3_U2360;
  assign new_P3_U5844 = ~new_P3_U3760 | ~new_P3_U3754 | ~new_P3_U5825 | ~new_P3_U3757 | ~new_P3_U5826;
  assign new_P3_U5845 = ~new_P3_U2402 | ~P3_REIP_REG_8_;
  assign new_P3_U5846 = ~new_P3_U4318 | ~new_P3_U5844;
  assign new_P3_U5847 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_U5631;
  assign new_P3_U5848 = ~new_P3_ADD_360_1242_U106 | ~new_P3_U2395;
  assign new_P3_U5849 = ~new_P3_SUB_357_1258_U70 | ~new_P3_U2393;
  assign new_P3_U5850 = ~new_P3_ADD_558_U65 | ~new_P3_U3220;
  assign new_P3_U5851 = ~new_P3_ADD_553_U65 | ~new_P3_U4298;
  assign new_P3_U5852 = ~new_P3_ADD_547_U65 | ~new_P3_U4299;
  assign new_P3_U5853 = ~new_P3_ADD_541_U62 | ~new_P3_U4300;
  assign new_P3_U5854 = ~new_P3_ADD_536_U62 | ~new_P3_U4301;
  assign new_P3_U5855 = ~new_P3_ADD_531_U65 | ~new_P3_U2354;
  assign new_P3_U5856 = ~new_P3_ADD_526_U51 | ~new_P3_U2355;
  assign new_P3_U5857 = ~new_P3_ADD_515_U62 | ~new_P3_U4302;
  assign new_P3_U5858 = ~new_P3_ADD_494_U62 | ~new_P3_U2356;
  assign new_P3_U5859 = ~new_P3_ADD_476_U62 | ~new_P3_U4303;
  assign new_P3_U5860 = ~new_P3_ADD_441_U62 | ~new_P3_U4304;
  assign new_P3_U5861 = ~new_P3_ADD_405_U63 | ~new_P3_U4305;
  assign new_P3_U5862 = ~new_P3_ADD_394_U63 | ~new_P3_U2357;
  assign new_P3_U5863 = ~new_P3_ADD_385_U65 | ~new_P3_U2358;
  assign new_P3_U5864 = ~new_P3_ADD_380_U65 | ~new_P3_U2359;
  assign new_P3_U5865 = ~new_P3_ADD_349_U65 | ~new_P3_U4306;
  assign new_P3_U5866 = ~new_P3_ADD_344_U65 | ~new_P3_U2362;
  assign new_P3_U5867 = ~new_P3_ADD_371_1212_U109 | ~new_P3_U2360;
  assign new_P3_U5868 = ~new_P3_U3767 | ~new_P3_U3761 | ~new_P3_U5849 | ~new_P3_U3764 | ~new_P3_U5850;
  assign new_P3_U5869 = ~new_P3_U2402 | ~P3_REIP_REG_9_;
  assign new_P3_U5870 = ~new_P3_U4318 | ~new_P3_U5868;
  assign new_P3_U5871 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_U5631;
  assign new_P3_U5872 = ~new_P3_ADD_360_1242_U4 | ~new_P3_U2395;
  assign new_P3_U5873 = ~new_P3_SUB_357_1258_U93 | ~new_P3_U2393;
  assign new_P3_U5874 = ~new_P3_ADD_558_U95 | ~new_P3_U3220;
  assign new_P3_U5875 = ~new_P3_ADD_553_U95 | ~new_P3_U4298;
  assign new_P3_U5876 = ~new_P3_ADD_547_U95 | ~new_P3_U4299;
  assign new_P3_U5877 = ~new_P3_ADD_541_U91 | ~new_P3_U4300;
  assign new_P3_U5878 = ~new_P3_ADD_536_U91 | ~new_P3_U4301;
  assign new_P3_U5879 = ~new_P3_ADD_531_U95 | ~new_P3_U2354;
  assign new_P3_U5880 = ~new_P3_ADD_526_U81 | ~new_P3_U2355;
  assign new_P3_U5881 = ~new_P3_ADD_515_U91 | ~new_P3_U4302;
  assign new_P3_U5882 = ~new_P3_ADD_494_U91 | ~new_P3_U2356;
  assign new_P3_U5883 = ~new_P3_ADD_476_U91 | ~new_P3_U4303;
  assign new_P3_U5884 = ~new_P3_ADD_441_U91 | ~new_P3_U4304;
  assign new_P3_U5885 = ~new_P3_ADD_405_U91 | ~new_P3_U4305;
  assign new_P3_U5886 = ~new_P3_ADD_394_U91 | ~new_P3_U2357;
  assign new_P3_U5887 = ~new_P3_ADD_385_U95 | ~new_P3_U2358;
  assign new_P3_U5888 = ~new_P3_ADD_380_U95 | ~new_P3_U2359;
  assign new_P3_U5889 = ~new_P3_ADD_349_U95 | ~new_P3_U4306;
  assign new_P3_U5890 = ~new_P3_ADD_344_U95 | ~new_P3_U2362;
  assign new_P3_U5891 = ~new_P3_ADD_371_1212_U5 | ~new_P3_U2360;
  assign new_P3_U5892 = ~new_P3_U3768 | ~new_P3_U3774 | ~new_P3_U5872 | ~new_P3_U5874 | ~new_P3_U3771;
  assign new_P3_U5893 = ~new_P3_U2402 | ~P3_REIP_REG_10_;
  assign new_P3_U5894 = ~new_P3_U4318 | ~new_P3_U5892;
  assign new_P3_U5895 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_U5631;
  assign new_P3_U5896 = ~new_P3_ADD_360_1242_U84 | ~new_P3_U2395;
  assign new_P3_U5897 = ~new_P3_SUB_357_1258_U92 | ~new_P3_U2393;
  assign new_P3_U5898 = ~new_P3_ADD_558_U94 | ~new_P3_U3220;
  assign new_P3_U5899 = ~new_P3_ADD_553_U94 | ~new_P3_U4298;
  assign new_P3_U5900 = ~new_P3_ADD_547_U94 | ~new_P3_U4299;
  assign new_P3_U5901 = ~new_P3_ADD_541_U90 | ~new_P3_U4300;
  assign new_P3_U5902 = ~new_P3_ADD_536_U90 | ~new_P3_U4301;
  assign new_P3_U5903 = ~new_P3_ADD_531_U94 | ~new_P3_U2354;
  assign new_P3_U5904 = ~new_P3_ADD_526_U80 | ~new_P3_U2355;
  assign new_P3_U5905 = ~new_P3_ADD_515_U90 | ~new_P3_U4302;
  assign new_P3_U5906 = ~new_P3_ADD_494_U90 | ~new_P3_U2356;
  assign new_P3_U5907 = ~new_P3_ADD_476_U90 | ~new_P3_U4303;
  assign new_P3_U5908 = ~new_P3_ADD_441_U90 | ~new_P3_U4304;
  assign new_P3_U5909 = ~new_P3_ADD_405_U90 | ~new_P3_U4305;
  assign new_P3_U5910 = ~new_P3_ADD_394_U90 | ~new_P3_U2357;
  assign new_P3_U5911 = ~new_P3_ADD_385_U94 | ~new_P3_U2358;
  assign new_P3_U5912 = ~new_P3_ADD_380_U94 | ~new_P3_U2359;
  assign new_P3_U5913 = ~new_P3_ADD_349_U94 | ~new_P3_U4306;
  assign new_P3_U5914 = ~new_P3_ADD_344_U94 | ~new_P3_U2362;
  assign new_P3_U5915 = ~new_P3_ADD_371_1212_U86 | ~new_P3_U2360;
  assign new_P3_U5916 = ~new_P3_U3781 | ~new_P3_U3775 | ~new_P3_U5896 | ~new_P3_U5898 | ~new_P3_U3778;
  assign new_P3_U5917 = ~new_P3_U2402 | ~P3_REIP_REG_11_;
  assign new_P3_U5918 = ~new_P3_U4318 | ~new_P3_U5916;
  assign new_P3_U5919 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_U5631;
  assign new_P3_U5920 = ~new_P3_ADD_360_1242_U5 | ~new_P3_U2395;
  assign new_P3_U5921 = ~new_P3_SUB_357_1258_U91 | ~new_P3_U2393;
  assign new_P3_U5922 = ~new_P3_ADD_558_U93 | ~new_P3_U3220;
  assign new_P3_U5923 = ~new_P3_ADD_553_U93 | ~new_P3_U4298;
  assign new_P3_U5924 = ~new_P3_ADD_547_U93 | ~new_P3_U4299;
  assign new_P3_U5925 = ~new_P3_ADD_541_U89 | ~new_P3_U4300;
  assign new_P3_U5926 = ~new_P3_ADD_536_U89 | ~new_P3_U4301;
  assign new_P3_U5927 = ~new_P3_ADD_531_U93 | ~new_P3_U2354;
  assign new_P3_U5928 = ~new_P3_ADD_526_U79 | ~new_P3_U2355;
  assign new_P3_U5929 = ~new_P3_ADD_515_U89 | ~new_P3_U4302;
  assign new_P3_U5930 = ~new_P3_ADD_494_U89 | ~new_P3_U2356;
  assign new_P3_U5931 = ~new_P3_ADD_476_U89 | ~new_P3_U4303;
  assign new_P3_U5932 = ~new_P3_ADD_441_U89 | ~new_P3_U4304;
  assign new_P3_U5933 = ~new_P3_ADD_405_U89 | ~new_P3_U4305;
  assign new_P3_U5934 = ~new_P3_ADD_394_U89 | ~new_P3_U2357;
  assign new_P3_U5935 = ~new_P3_ADD_385_U93 | ~new_P3_U2358;
  assign new_P3_U5936 = ~new_P3_ADD_380_U93 | ~new_P3_U2359;
  assign new_P3_U5937 = ~new_P3_ADD_349_U93 | ~new_P3_U4306;
  assign new_P3_U5938 = ~new_P3_ADD_344_U93 | ~new_P3_U2362;
  assign new_P3_U5939 = ~new_P3_ADD_371_1212_U6 | ~new_P3_U2360;
  assign new_P3_U5940 = ~new_P3_U3788 | ~new_P3_U3782 | ~new_P3_U5921 | ~new_P3_U3785 | ~new_P3_U5922;
  assign new_P3_U5941 = ~new_P3_U2402 | ~P3_REIP_REG_12_;
  assign new_P3_U5942 = ~new_P3_U4318 | ~new_P3_U5940;
  assign new_P3_U5943 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_U5631;
  assign new_P3_U5944 = ~new_P3_ADD_360_1242_U6 | ~new_P3_U2395;
  assign new_P3_U5945 = ~new_P3_SUB_357_1258_U15 | ~new_P3_U2393;
  assign new_P3_U5946 = ~new_P3_ADD_558_U92 | ~new_P3_U3220;
  assign new_P3_U5947 = ~new_P3_ADD_553_U92 | ~new_P3_U4298;
  assign new_P3_U5948 = ~new_P3_ADD_547_U92 | ~new_P3_U4299;
  assign new_P3_U5949 = ~new_P3_ADD_541_U88 | ~new_P3_U4300;
  assign new_P3_U5950 = ~new_P3_ADD_536_U88 | ~new_P3_U4301;
  assign new_P3_U5951 = ~new_P3_ADD_531_U92 | ~new_P3_U2354;
  assign new_P3_U5952 = ~new_P3_ADD_526_U78 | ~new_P3_U2355;
  assign new_P3_U5953 = ~new_P3_ADD_515_U88 | ~new_P3_U4302;
  assign new_P3_U5954 = ~new_P3_ADD_494_U88 | ~new_P3_U2356;
  assign new_P3_U5955 = ~new_P3_ADD_476_U88 | ~new_P3_U4303;
  assign new_P3_U5956 = ~new_P3_ADD_441_U88 | ~new_P3_U4304;
  assign new_P3_U5957 = ~new_P3_ADD_405_U88 | ~new_P3_U4305;
  assign new_P3_U5958 = ~new_P3_ADD_394_U88 | ~new_P3_U2357;
  assign new_P3_U5959 = ~new_P3_ADD_385_U92 | ~new_P3_U2358;
  assign new_P3_U5960 = ~new_P3_ADD_380_U92 | ~new_P3_U2359;
  assign new_P3_U5961 = ~new_P3_ADD_349_U92 | ~new_P3_U4306;
  assign new_P3_U5962 = ~new_P3_ADD_344_U92 | ~new_P3_U2362;
  assign new_P3_U5963 = ~new_P3_ADD_371_1212_U7 | ~new_P3_U2360;
  assign new_P3_U5964 = ~new_P3_U3795 | ~new_P3_U3789 | ~new_P3_U5945 | ~new_P3_U3792 | ~new_P3_U5946;
  assign new_P3_U5965 = ~new_P3_U2402 | ~P3_REIP_REG_13_;
  assign new_P3_U5966 = ~new_P3_U4318 | ~new_P3_U5964;
  assign new_P3_U5967 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_U5631;
  assign new_P3_U5968 = ~new_P3_ADD_360_1242_U83 | ~new_P3_U2395;
  assign new_P3_U5969 = ~new_P3_SUB_357_1258_U90 | ~new_P3_U2393;
  assign new_P3_U5970 = ~new_P3_ADD_558_U91 | ~new_P3_U3220;
  assign new_P3_U5971 = ~new_P3_ADD_553_U91 | ~new_P3_U4298;
  assign new_P3_U5972 = ~new_P3_ADD_547_U91 | ~new_P3_U4299;
  assign new_P3_U5973 = ~new_P3_ADD_541_U87 | ~new_P3_U4300;
  assign new_P3_U5974 = ~new_P3_ADD_536_U87 | ~new_P3_U4301;
  assign new_P3_U5975 = ~new_P3_ADD_531_U91 | ~new_P3_U2354;
  assign new_P3_U5976 = ~new_P3_ADD_526_U77 | ~new_P3_U2355;
  assign new_P3_U5977 = ~new_P3_ADD_515_U87 | ~new_P3_U4302;
  assign new_P3_U5978 = ~new_P3_ADD_494_U87 | ~new_P3_U2356;
  assign new_P3_U5979 = ~new_P3_ADD_476_U87 | ~new_P3_U4303;
  assign new_P3_U5980 = ~new_P3_ADD_441_U87 | ~new_P3_U4304;
  assign new_P3_U5981 = ~new_P3_ADD_405_U87 | ~new_P3_U4305;
  assign new_P3_U5982 = ~new_P3_ADD_394_U87 | ~new_P3_U2357;
  assign new_P3_U5983 = ~new_P3_ADD_385_U91 | ~new_P3_U2358;
  assign new_P3_U5984 = ~new_P3_ADD_380_U91 | ~new_P3_U2359;
  assign new_P3_U5985 = ~new_P3_ADD_349_U91 | ~new_P3_U4306;
  assign new_P3_U5986 = ~new_P3_ADD_344_U91 | ~new_P3_U2362;
  assign new_P3_U5987 = ~new_P3_ADD_371_1212_U85 | ~new_P3_U2360;
  assign new_P3_U5988 = ~new_P3_U3802 | ~new_P3_U3799;
  assign new_P3_U5989 = ~new_P3_U2402 | ~P3_REIP_REG_14_;
  assign new_P3_U5990 = ~new_P3_U4318 | ~new_P3_U5988;
  assign new_P3_U5991 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_U5631;
  assign new_P3_U5992 = ~new_P3_ADD_360_1242_U7 | ~new_P3_U2395;
  assign new_P3_U5993 = ~new_P3_SUB_357_1258_U89 | ~new_P3_U2393;
  assign new_P3_U5994 = ~new_P3_ADD_558_U90 | ~new_P3_U3220;
  assign new_P3_U5995 = ~new_P3_ADD_553_U90 | ~new_P3_U4298;
  assign new_P3_U5996 = ~new_P3_ADD_547_U90 | ~new_P3_U4299;
  assign new_P3_U5997 = ~new_P3_ADD_541_U86 | ~new_P3_U4300;
  assign new_P3_U5998 = ~new_P3_ADD_536_U86 | ~new_P3_U4301;
  assign new_P3_U5999 = ~new_P3_ADD_531_U90 | ~new_P3_U2354;
  assign new_P3_U6000 = ~new_P3_ADD_526_U76 | ~new_P3_U2355;
  assign new_P3_U6001 = ~new_P3_ADD_515_U86 | ~new_P3_U4302;
  assign new_P3_U6002 = ~new_P3_ADD_494_U86 | ~new_P3_U2356;
  assign new_P3_U6003 = ~new_P3_ADD_476_U86 | ~new_P3_U4303;
  assign new_P3_U6004 = ~new_P3_ADD_441_U86 | ~new_P3_U4304;
  assign new_P3_U6005 = ~new_P3_ADD_405_U86 | ~new_P3_U4305;
  assign new_P3_U6006 = ~new_P3_ADD_394_U86 | ~new_P3_U2357;
  assign new_P3_U6007 = ~new_P3_ADD_385_U90 | ~new_P3_U2358;
  assign new_P3_U6008 = ~new_P3_ADD_380_U90 | ~new_P3_U2359;
  assign new_P3_U6009 = ~new_P3_ADD_349_U90 | ~new_P3_U4306;
  assign new_P3_U6010 = ~new_P3_ADD_344_U90 | ~new_P3_U2362;
  assign new_P3_U6011 = ~new_P3_ADD_371_1212_U8 | ~new_P3_U2360;
  assign new_P3_U6012 = ~new_P3_U3810 | ~new_P3_U3807;
  assign new_P3_U6013 = ~new_P3_U2402 | ~P3_REIP_REG_15_;
  assign new_P3_U6014 = ~new_P3_U4318 | ~new_P3_U6012;
  assign new_P3_U6015 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_U5631;
  assign new_P3_U6016 = ~new_P3_ADD_360_1242_U82 | ~new_P3_U2395;
  assign new_P3_U6017 = ~new_P3_SUB_357_1258_U88 | ~new_P3_U2393;
  assign new_P3_U6018 = ~new_P3_ADD_558_U89 | ~new_P3_U3220;
  assign new_P3_U6019 = ~new_P3_ADD_553_U89 | ~new_P3_U4298;
  assign new_P3_U6020 = ~new_P3_ADD_547_U89 | ~new_P3_U4299;
  assign new_P3_U6021 = ~new_P3_ADD_541_U85 | ~new_P3_U4300;
  assign new_P3_U6022 = ~new_P3_ADD_536_U85 | ~new_P3_U4301;
  assign new_P3_U6023 = ~new_P3_ADD_531_U89 | ~new_P3_U2354;
  assign new_P3_U6024 = ~new_P3_ADD_526_U75 | ~new_P3_U2355;
  assign new_P3_U6025 = ~new_P3_ADD_515_U85 | ~new_P3_U4302;
  assign new_P3_U6026 = ~new_P3_ADD_494_U85 | ~new_P3_U2356;
  assign new_P3_U6027 = ~new_P3_ADD_476_U85 | ~new_P3_U4303;
  assign new_P3_U6028 = ~new_P3_ADD_441_U85 | ~new_P3_U4304;
  assign new_P3_U6029 = ~new_P3_ADD_405_U85 | ~new_P3_U4305;
  assign new_P3_U6030 = ~new_P3_ADD_394_U85 | ~new_P3_U2357;
  assign new_P3_U6031 = ~new_P3_ADD_385_U89 | ~new_P3_U2358;
  assign new_P3_U6032 = ~new_P3_ADD_380_U89 | ~new_P3_U2359;
  assign new_P3_U6033 = ~new_P3_ADD_349_U89 | ~new_P3_U4306;
  assign new_P3_U6034 = ~new_P3_ADD_344_U89 | ~new_P3_U2362;
  assign new_P3_U6035 = ~new_P3_ADD_371_1212_U84 | ~new_P3_U2360;
  assign new_P3_U6036 = ~new_P3_U3818 | ~new_P3_U3812 | ~new_P3_U6016 | ~new_P3_U6018 | ~new_P3_U3815;
  assign new_P3_U6037 = ~new_P3_U2402 | ~P3_REIP_REG_16_;
  assign new_P3_U6038 = ~new_P3_U4318 | ~new_P3_U6036;
  assign new_P3_U6039 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_U5631;
  assign new_P3_U6040 = ~new_P3_ADD_360_1242_U8 | ~new_P3_U2395;
  assign new_P3_U6041 = ~new_P3_SUB_357_1258_U16 | ~new_P3_U2393;
  assign new_P3_U6042 = ~new_P3_ADD_558_U88 | ~new_P3_U3220;
  assign new_P3_U6043 = ~new_P3_ADD_553_U88 | ~new_P3_U4298;
  assign new_P3_U6044 = ~new_P3_ADD_547_U88 | ~new_P3_U4299;
  assign new_P3_U6045 = ~new_P3_ADD_541_U84 | ~new_P3_U4300;
  assign new_P3_U6046 = ~new_P3_ADD_536_U84 | ~new_P3_U4301;
  assign new_P3_U6047 = ~new_P3_ADD_531_U88 | ~new_P3_U2354;
  assign new_P3_U6048 = ~new_P3_ADD_526_U74 | ~new_P3_U2355;
  assign new_P3_U6049 = ~new_P3_ADD_515_U84 | ~new_P3_U4302;
  assign new_P3_U6050 = ~new_P3_ADD_494_U84 | ~new_P3_U2356;
  assign new_P3_U6051 = ~new_P3_ADD_476_U84 | ~new_P3_U4303;
  assign new_P3_U6052 = ~new_P3_ADD_441_U84 | ~new_P3_U4304;
  assign new_P3_U6053 = ~new_P3_ADD_405_U84 | ~new_P3_U4305;
  assign new_P3_U6054 = ~new_P3_ADD_394_U84 | ~new_P3_U2357;
  assign new_P3_U6055 = ~new_P3_ADD_385_U88 | ~new_P3_U2358;
  assign new_P3_U6056 = ~new_P3_ADD_380_U88 | ~new_P3_U2359;
  assign new_P3_U6057 = ~new_P3_ADD_349_U88 | ~new_P3_U4306;
  assign new_P3_U6058 = ~new_P3_ADD_344_U88 | ~new_P3_U2362;
  assign new_P3_U6059 = ~new_P3_ADD_371_1212_U9 | ~new_P3_U2360;
  assign new_P3_U6060 = ~new_P3_U3820 | ~new_P3_U3824 | ~new_P3_U6040 | ~new_P3_U6042 | ~new_P3_U3819;
  assign new_P3_U6061 = ~new_P3_U2402 | ~P3_REIP_REG_17_;
  assign new_P3_U6062 = ~new_P3_U4318 | ~new_P3_U6060;
  assign new_P3_U6063 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_U5631;
  assign new_P3_U6064 = ~new_P3_ADD_360_1242_U81 | ~new_P3_U2395;
  assign new_P3_U6065 = ~new_P3_SUB_357_1258_U87 | ~new_P3_U2393;
  assign new_P3_U6066 = ~new_P3_ADD_558_U87 | ~new_P3_U3220;
  assign new_P3_U6067 = ~new_P3_ADD_553_U87 | ~new_P3_U4298;
  assign new_P3_U6068 = ~new_P3_ADD_547_U87 | ~new_P3_U4299;
  assign new_P3_U6069 = ~new_P3_ADD_541_U83 | ~new_P3_U4300;
  assign new_P3_U6070 = ~new_P3_ADD_536_U83 | ~new_P3_U4301;
  assign new_P3_U6071 = ~new_P3_ADD_531_U87 | ~new_P3_U2354;
  assign new_P3_U6072 = ~new_P3_ADD_526_U73 | ~new_P3_U2355;
  assign new_P3_U6073 = ~new_P3_ADD_515_U83 | ~new_P3_U4302;
  assign new_P3_U6074 = ~new_P3_ADD_494_U83 | ~new_P3_U2356;
  assign new_P3_U6075 = ~new_P3_ADD_476_U83 | ~new_P3_U4303;
  assign new_P3_U6076 = ~new_P3_ADD_441_U83 | ~new_P3_U4304;
  assign new_P3_U6077 = ~new_P3_ADD_405_U83 | ~new_P3_U4305;
  assign new_P3_U6078 = ~new_P3_ADD_394_U83 | ~new_P3_U2357;
  assign new_P3_U6079 = ~new_P3_ADD_385_U87 | ~new_P3_U2358;
  assign new_P3_U6080 = ~new_P3_ADD_380_U87 | ~new_P3_U2359;
  assign new_P3_U6081 = ~new_P3_ADD_349_U87 | ~new_P3_U4306;
  assign new_P3_U6082 = ~new_P3_ADD_344_U87 | ~new_P3_U2362;
  assign new_P3_U6083 = ~new_P3_ADD_371_1212_U83 | ~new_P3_U2360;
  assign new_P3_U6084 = ~new_P3_U3831 | ~new_P3_U3825 | ~new_P3_U6064 | ~new_P3_U6066 | ~new_P3_U3828;
  assign new_P3_U6085 = ~new_P3_U2402 | ~P3_REIP_REG_18_;
  assign new_P3_U6086 = ~new_P3_U4318 | ~new_P3_U6084;
  assign new_P3_U6087 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_U5631;
  assign new_P3_U6088 = ~new_P3_ADD_360_1242_U9 | ~new_P3_U2395;
  assign new_P3_U6089 = ~new_P3_SUB_357_1258_U86 | ~new_P3_U2393;
  assign new_P3_U6090 = ~new_P3_ADD_558_U86 | ~new_P3_U3220;
  assign new_P3_U6091 = ~new_P3_ADD_553_U86 | ~new_P3_U4298;
  assign new_P3_U6092 = ~new_P3_ADD_547_U86 | ~new_P3_U4299;
  assign new_P3_U6093 = ~new_P3_ADD_541_U82 | ~new_P3_U4300;
  assign new_P3_U6094 = ~new_P3_ADD_536_U82 | ~new_P3_U4301;
  assign new_P3_U6095 = ~new_P3_ADD_531_U86 | ~new_P3_U2354;
  assign new_P3_U6096 = ~new_P3_ADD_526_U72 | ~new_P3_U2355;
  assign new_P3_U6097 = ~new_P3_ADD_515_U82 | ~new_P3_U4302;
  assign new_P3_U6098 = ~new_P3_ADD_494_U82 | ~new_P3_U2356;
  assign new_P3_U6099 = ~new_P3_ADD_476_U82 | ~new_P3_U4303;
  assign new_P3_U6100 = ~new_P3_ADD_441_U82 | ~new_P3_U4304;
  assign new_P3_U6101 = ~new_P3_ADD_405_U82 | ~new_P3_U4305;
  assign new_P3_U6102 = ~new_P3_ADD_394_U82 | ~new_P3_U2357;
  assign new_P3_U6103 = ~new_P3_ADD_385_U86 | ~new_P3_U2358;
  assign new_P3_U6104 = ~new_P3_ADD_380_U86 | ~new_P3_U2359;
  assign new_P3_U6105 = ~new_P3_ADD_349_U86 | ~new_P3_U4306;
  assign new_P3_U6106 = ~new_P3_ADD_344_U86 | ~new_P3_U2362;
  assign new_P3_U6107 = ~new_P3_ADD_371_1212_U10 | ~new_P3_U2360;
  assign new_P3_U6108 = ~new_P3_U3833 | ~new_P3_U3837 | ~new_P3_U6088 | ~new_P3_U6090 | ~new_P3_U3832;
  assign new_P3_U6109 = ~new_P3_U2402 | ~P3_REIP_REG_19_;
  assign new_P3_U6110 = ~new_P3_U4318 | ~new_P3_U6108;
  assign new_P3_U6111 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_U5631;
  assign new_P3_U6112 = ~new_P3_ADD_360_1242_U10 | ~new_P3_U2395;
  assign new_P3_U6113 = ~new_P3_SUB_357_1258_U17 | ~new_P3_U2393;
  assign new_P3_U6114 = ~new_P3_ADD_558_U84 | ~new_P3_U3220;
  assign new_P3_U6115 = ~new_P3_ADD_553_U84 | ~new_P3_U4298;
  assign new_P3_U6116 = ~new_P3_ADD_547_U84 | ~new_P3_U4299;
  assign new_P3_U6117 = ~new_P3_ADD_541_U81 | ~new_P3_U4300;
  assign new_P3_U6118 = ~new_P3_ADD_536_U81 | ~new_P3_U4301;
  assign new_P3_U6119 = ~new_P3_ADD_531_U84 | ~new_P3_U2354;
  assign new_P3_U6120 = ~new_P3_ADD_526_U70 | ~new_P3_U2355;
  assign new_P3_U6121 = ~new_P3_ADD_515_U81 | ~new_P3_U4302;
  assign new_P3_U6122 = ~new_P3_ADD_494_U81 | ~new_P3_U2356;
  assign new_P3_U6123 = ~new_P3_ADD_476_U81 | ~new_P3_U4303;
  assign new_P3_U6124 = ~new_P3_ADD_441_U81 | ~new_P3_U4304;
  assign new_P3_U6125 = ~new_P3_ADD_405_U80 | ~new_P3_U4305;
  assign new_P3_U6126 = ~new_P3_ADD_394_U80 | ~new_P3_U2357;
  assign new_P3_U6127 = ~new_P3_ADD_385_U84 | ~new_P3_U2358;
  assign new_P3_U6128 = ~new_P3_ADD_380_U84 | ~new_P3_U2359;
  assign new_P3_U6129 = ~new_P3_ADD_349_U84 | ~new_P3_U4306;
  assign new_P3_U6130 = ~new_P3_ADD_344_U84 | ~new_P3_U2362;
  assign new_P3_U6131 = ~new_P3_ADD_371_1212_U11 | ~new_P3_U2360;
  assign new_P3_U6132 = ~new_P3_U6113 | ~new_P3_U3841;
  assign new_P3_U6133 = ~new_P3_U2402 | ~P3_REIP_REG_20_;
  assign new_P3_U6134 = ~new_P3_U4318 | ~new_P3_U6132;
  assign new_P3_U6135 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_U5631;
  assign new_P3_U6136 = ~new_P3_ADD_360_1242_U11 | ~new_P3_U2395;
  assign new_P3_U6137 = ~new_P3_SUB_357_1258_U85 | ~new_P3_U2393;
  assign new_P3_U6138 = ~new_P3_ADD_558_U83 | ~new_P3_U3220;
  assign new_P3_U6139 = ~new_P3_ADD_553_U83 | ~new_P3_U4298;
  assign new_P3_U6140 = ~new_P3_ADD_547_U83 | ~new_P3_U4299;
  assign new_P3_U6141 = ~new_P3_ADD_541_U80 | ~new_P3_U4300;
  assign new_P3_U6142 = ~new_P3_ADD_536_U80 | ~new_P3_U4301;
  assign new_P3_U6143 = ~new_P3_ADD_531_U83 | ~new_P3_U2354;
  assign new_P3_U6144 = ~new_P3_ADD_526_U69 | ~new_P3_U2355;
  assign new_P3_U6145 = ~new_P3_ADD_515_U80 | ~new_P3_U4302;
  assign new_P3_U6146 = ~new_P3_ADD_494_U80 | ~new_P3_U2356;
  assign new_P3_U6147 = ~new_P3_ADD_476_U80 | ~new_P3_U4303;
  assign new_P3_U6148 = ~new_P3_ADD_441_U80 | ~new_P3_U4304;
  assign new_P3_U6149 = ~new_P3_ADD_405_U79 | ~new_P3_U4305;
  assign new_P3_U6150 = ~new_P3_ADD_394_U79 | ~new_P3_U2357;
  assign new_P3_U6151 = ~new_P3_ADD_385_U83 | ~new_P3_U2358;
  assign new_P3_U6152 = ~new_P3_ADD_380_U83 | ~new_P3_U2359;
  assign new_P3_U6153 = ~new_P3_ADD_349_U83 | ~new_P3_U4306;
  assign new_P3_U6154 = ~new_P3_ADD_344_U83 | ~new_P3_U2362;
  assign new_P3_U6155 = ~new_P3_ADD_371_1212_U12 | ~new_P3_U2360;
  assign new_P3_U6156 = ~new_P3_U6137 | ~new_P3_U3849;
  assign new_P3_U6157 = ~new_P3_U2402 | ~P3_REIP_REG_21_;
  assign new_P3_U6158 = ~new_P3_U4318 | ~new_P3_U6156;
  assign new_P3_U6159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_U5631;
  assign new_P3_U6160 = ~new_P3_ADD_360_1242_U80 | ~new_P3_U2395;
  assign new_P3_U6161 = ~new_P3_SUB_357_1258_U84 | ~new_P3_U2393;
  assign new_P3_U6162 = ~new_P3_ADD_558_U82 | ~new_P3_U3220;
  assign new_P3_U6163 = ~new_P3_ADD_553_U82 | ~new_P3_U4298;
  assign new_P3_U6164 = ~new_P3_ADD_547_U82 | ~new_P3_U4299;
  assign new_P3_U6165 = ~new_P3_ADD_541_U79 | ~new_P3_U4300;
  assign new_P3_U6166 = ~new_P3_ADD_536_U79 | ~new_P3_U4301;
  assign new_P3_U6167 = ~new_P3_ADD_531_U82 | ~new_P3_U2354;
  assign new_P3_U6168 = ~new_P3_ADD_526_U68 | ~new_P3_U2355;
  assign new_P3_U6169 = ~new_P3_ADD_515_U79 | ~new_P3_U4302;
  assign new_P3_U6170 = ~new_P3_ADD_494_U79 | ~new_P3_U2356;
  assign new_P3_U6171 = ~new_P3_ADD_476_U79 | ~new_P3_U4303;
  assign new_P3_U6172 = ~new_P3_ADD_441_U79 | ~new_P3_U4304;
  assign new_P3_U6173 = ~new_P3_ADD_405_U78 | ~new_P3_U4305;
  assign new_P3_U6174 = ~new_P3_ADD_394_U78 | ~new_P3_U2357;
  assign new_P3_U6175 = ~new_P3_ADD_385_U82 | ~new_P3_U2358;
  assign new_P3_U6176 = ~new_P3_ADD_380_U82 | ~new_P3_U2359;
  assign new_P3_U6177 = ~new_P3_ADD_349_U82 | ~new_P3_U4306;
  assign new_P3_U6178 = ~new_P3_ADD_344_U82 | ~new_P3_U2362;
  assign new_P3_U6179 = ~new_P3_ADD_371_1212_U82 | ~new_P3_U2360;
  assign new_P3_U6180 = ~new_P3_U3862 | ~new_P3_U3857;
  assign new_P3_U6181 = ~new_P3_U2402 | ~P3_REIP_REG_22_;
  assign new_P3_U6182 = ~new_P3_U4318 | ~new_P3_U6180;
  assign new_P3_U6183 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_U5631;
  assign new_P3_U6184 = ~new_P3_ADD_360_1242_U12 | ~new_P3_U2395;
  assign new_P3_U6185 = ~new_P3_SUB_357_1258_U83 | ~new_P3_U2393;
  assign new_P3_U6186 = ~new_P3_ADD_558_U81 | ~new_P3_U3220;
  assign new_P3_U6187 = ~new_P3_ADD_553_U81 | ~new_P3_U4298;
  assign new_P3_U6188 = ~new_P3_ADD_547_U81 | ~new_P3_U4299;
  assign new_P3_U6189 = ~new_P3_ADD_541_U78 | ~new_P3_U4300;
  assign new_P3_U6190 = ~new_P3_ADD_536_U78 | ~new_P3_U4301;
  assign new_P3_U6191 = ~new_P3_ADD_531_U81 | ~new_P3_U2354;
  assign new_P3_U6192 = ~new_P3_ADD_526_U67 | ~new_P3_U2355;
  assign new_P3_U6193 = ~new_P3_ADD_515_U78 | ~new_P3_U4302;
  assign new_P3_U6194 = ~new_P3_ADD_494_U78 | ~new_P3_U2356;
  assign new_P3_U6195 = ~new_P3_ADD_476_U78 | ~new_P3_U4303;
  assign new_P3_U6196 = ~new_P3_ADD_441_U78 | ~new_P3_U4304;
  assign new_P3_U6197 = ~new_P3_ADD_405_U77 | ~new_P3_U4305;
  assign new_P3_U6198 = ~new_P3_ADD_394_U77 | ~new_P3_U2357;
  assign new_P3_U6199 = ~new_P3_ADD_385_U81 | ~new_P3_U2358;
  assign new_P3_U6200 = ~new_P3_ADD_380_U81 | ~new_P3_U2359;
  assign new_P3_U6201 = ~new_P3_ADD_349_U81 | ~new_P3_U4306;
  assign new_P3_U6202 = ~new_P3_ADD_344_U81 | ~new_P3_U2362;
  assign new_P3_U6203 = ~new_P3_ADD_371_1212_U13 | ~new_P3_U2360;
  assign new_P3_U6204 = ~new_P3_U3872 | ~new_P3_U3867;
  assign new_P3_U6205 = ~new_P3_U2402 | ~P3_REIP_REG_23_;
  assign new_P3_U6206 = ~new_P3_U4318 | ~new_P3_U6204;
  assign new_P3_U6207 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_U5631;
  assign new_P3_U6208 = ~new_P3_ADD_360_1242_U79 | ~new_P3_U2395;
  assign new_P3_U6209 = ~new_P3_SUB_357_1258_U82 | ~new_P3_U2393;
  assign new_P3_U6210 = ~new_P3_ADD_558_U80 | ~new_P3_U3220;
  assign new_P3_U6211 = ~new_P3_ADD_553_U80 | ~new_P3_U4298;
  assign new_P3_U6212 = ~new_P3_ADD_547_U80 | ~new_P3_U4299;
  assign new_P3_U6213 = ~new_P3_ADD_541_U77 | ~new_P3_U4300;
  assign new_P3_U6214 = ~new_P3_ADD_536_U77 | ~new_P3_U4301;
  assign new_P3_U6215 = ~new_P3_ADD_531_U80 | ~new_P3_U2354;
  assign new_P3_U6216 = ~new_P3_ADD_526_U66 | ~new_P3_U2355;
  assign new_P3_U6217 = ~new_P3_ADD_515_U77 | ~new_P3_U4302;
  assign new_P3_U6218 = ~new_P3_ADD_494_U77 | ~new_P3_U2356;
  assign new_P3_U6219 = ~new_P3_ADD_476_U77 | ~new_P3_U4303;
  assign new_P3_U6220 = ~new_P3_ADD_441_U77 | ~new_P3_U4304;
  assign new_P3_U6221 = ~new_P3_ADD_405_U76 | ~new_P3_U4305;
  assign new_P3_U6222 = ~new_P3_ADD_394_U76 | ~new_P3_U2357;
  assign new_P3_U6223 = ~new_P3_ADD_385_U80 | ~new_P3_U2358;
  assign new_P3_U6224 = ~new_P3_ADD_380_U80 | ~new_P3_U2359;
  assign new_P3_U6225 = ~new_P3_ADD_349_U80 | ~new_P3_U4306;
  assign new_P3_U6226 = ~new_P3_ADD_344_U80 | ~new_P3_U2362;
  assign new_P3_U6227 = ~new_P3_ADD_371_1212_U81 | ~new_P3_U2360;
  assign new_P3_U6228 = ~new_P3_U3882 | ~new_P3_U3877;
  assign new_P3_U6229 = ~new_P3_U2402 | ~P3_REIP_REG_24_;
  assign new_P3_U6230 = ~new_P3_U4318 | ~new_P3_U6228;
  assign new_P3_U6231 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_U5631;
  assign new_P3_U6232 = ~new_P3_ADD_360_1242_U13 | ~new_P3_U2395;
  assign new_P3_U6233 = ~new_P3_SUB_357_1258_U81 | ~new_P3_U2393;
  assign new_P3_U6234 = ~new_P3_ADD_558_U79 | ~new_P3_U3220;
  assign new_P3_U6235 = ~new_P3_ADD_553_U79 | ~new_P3_U4298;
  assign new_P3_U6236 = ~new_P3_ADD_547_U79 | ~new_P3_U4299;
  assign new_P3_U6237 = ~new_P3_ADD_541_U76 | ~new_P3_U4300;
  assign new_P3_U6238 = ~new_P3_ADD_536_U76 | ~new_P3_U4301;
  assign new_P3_U6239 = ~new_P3_ADD_531_U79 | ~new_P3_U2354;
  assign new_P3_U6240 = ~new_P3_ADD_526_U65 | ~new_P3_U2355;
  assign new_P3_U6241 = ~new_P3_ADD_515_U76 | ~new_P3_U4302;
  assign new_P3_U6242 = ~new_P3_ADD_494_U76 | ~new_P3_U2356;
  assign new_P3_U6243 = ~new_P3_ADD_476_U76 | ~new_P3_U4303;
  assign new_P3_U6244 = ~new_P3_ADD_441_U76 | ~new_P3_U4304;
  assign new_P3_U6245 = ~new_P3_ADD_405_U75 | ~new_P3_U4305;
  assign new_P3_U6246 = ~new_P3_ADD_394_U75 | ~new_P3_U2357;
  assign new_P3_U6247 = ~new_P3_ADD_385_U79 | ~new_P3_U2358;
  assign new_P3_U6248 = ~new_P3_ADD_380_U79 | ~new_P3_U2359;
  assign new_P3_U6249 = ~new_P3_ADD_349_U79 | ~new_P3_U4306;
  assign new_P3_U6250 = ~new_P3_ADD_344_U79 | ~new_P3_U2362;
  assign new_P3_U6251 = ~new_P3_ADD_371_1212_U14 | ~new_P3_U2360;
  assign new_P3_U6252 = ~new_P3_U3892 | ~new_P3_U3887;
  assign new_P3_U6253 = ~new_P3_U2402 | ~P3_REIP_REG_25_;
  assign new_P3_U6254 = ~new_P3_U4318 | ~new_P3_U6252;
  assign new_P3_U6255 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_U5631;
  assign new_P3_U6256 = ~new_P3_ADD_360_1242_U14 | ~new_P3_U2395;
  assign new_P3_U6257 = ~new_P3_SUB_357_1258_U18 | ~new_P3_U2393;
  assign new_P3_U6258 = ~new_P3_ADD_558_U78 | ~new_P3_U3220;
  assign new_P3_U6259 = ~new_P3_ADD_553_U78 | ~new_P3_U4298;
  assign new_P3_U6260 = ~new_P3_ADD_547_U78 | ~new_P3_U4299;
  assign new_P3_U6261 = ~new_P3_ADD_541_U75 | ~new_P3_U4300;
  assign new_P3_U6262 = ~new_P3_ADD_536_U75 | ~new_P3_U4301;
  assign new_P3_U6263 = ~new_P3_ADD_531_U78 | ~new_P3_U2354;
  assign new_P3_U6264 = ~new_P3_ADD_526_U64 | ~new_P3_U2355;
  assign new_P3_U6265 = ~new_P3_ADD_515_U75 | ~new_P3_U4302;
  assign new_P3_U6266 = ~new_P3_ADD_494_U75 | ~new_P3_U2356;
  assign new_P3_U6267 = ~new_P3_ADD_476_U75 | ~new_P3_U4303;
  assign new_P3_U6268 = ~new_P3_ADD_441_U75 | ~new_P3_U4304;
  assign new_P3_U6269 = ~new_P3_ADD_405_U74 | ~new_P3_U4305;
  assign new_P3_U6270 = ~new_P3_ADD_394_U74 | ~new_P3_U2357;
  assign new_P3_U6271 = ~new_P3_ADD_385_U78 | ~new_P3_U2358;
  assign new_P3_U6272 = ~new_P3_ADD_380_U78 | ~new_P3_U2359;
  assign new_P3_U6273 = ~new_P3_ADD_349_U78 | ~new_P3_U4306;
  assign new_P3_U6274 = ~new_P3_ADD_344_U78 | ~new_P3_U2362;
  assign new_P3_U6275 = ~new_P3_ADD_371_1212_U15 | ~new_P3_U2360;
  assign new_P3_U6276 = ~new_P3_U3902 | ~new_P3_U3897 | ~new_P3_U3895 | ~new_P3_U3894 | ~new_P3_U6258;
  assign new_P3_U6277 = ~new_P3_U2402 | ~P3_REIP_REG_26_;
  assign new_P3_U6278 = ~new_P3_U4318 | ~new_P3_U6276;
  assign new_P3_U6279 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_U5631;
  assign new_P3_U6280 = ~new_P3_ADD_360_1242_U78 | ~new_P3_U2395;
  assign new_P3_U6281 = ~new_P3_SUB_357_1258_U80 | ~new_P3_U2393;
  assign new_P3_U6282 = ~new_P3_ADD_558_U77 | ~new_P3_U3220;
  assign new_P3_U6283 = ~new_P3_ADD_553_U77 | ~new_P3_U4298;
  assign new_P3_U6284 = ~new_P3_ADD_547_U77 | ~new_P3_U4299;
  assign new_P3_U6285 = ~new_P3_ADD_541_U74 | ~new_P3_U4300;
  assign new_P3_U6286 = ~new_P3_ADD_536_U74 | ~new_P3_U4301;
  assign new_P3_U6287 = ~new_P3_ADD_531_U77 | ~new_P3_U2354;
  assign new_P3_U6288 = ~new_P3_ADD_526_U63 | ~new_P3_U2355;
  assign new_P3_U6289 = ~new_P3_ADD_515_U74 | ~new_P3_U4302;
  assign new_P3_U6290 = ~new_P3_ADD_494_U74 | ~new_P3_U2356;
  assign new_P3_U6291 = ~new_P3_ADD_476_U74 | ~new_P3_U4303;
  assign new_P3_U6292 = ~new_P3_ADD_441_U74 | ~new_P3_U4304;
  assign new_P3_U6293 = ~new_P3_ADD_405_U73 | ~new_P3_U4305;
  assign new_P3_U6294 = ~new_P3_ADD_394_U73 | ~new_P3_U2357;
  assign new_P3_U6295 = ~new_P3_ADD_385_U77 | ~new_P3_U2358;
  assign new_P3_U6296 = ~new_P3_ADD_380_U77 | ~new_P3_U2359;
  assign new_P3_U6297 = ~new_P3_ADD_349_U77 | ~new_P3_U4306;
  assign new_P3_U6298 = ~new_P3_ADD_344_U77 | ~new_P3_U2362;
  assign new_P3_U6299 = ~new_P3_ADD_371_1212_U80 | ~new_P3_U2360;
  assign new_P3_U6300 = ~new_P3_U3911 | ~new_P3_U3906 | ~new_P3_U3904 | ~new_P3_U3903 | ~new_P3_U6282;
  assign new_P3_U6301 = ~new_P3_U2402 | ~P3_REIP_REG_27_;
  assign new_P3_U6302 = ~new_P3_U4318 | ~new_P3_U6300;
  assign new_P3_U6303 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_U5631;
  assign new_P3_U6304 = ~new_P3_ADD_360_1242_U15 | ~new_P3_U2395;
  assign new_P3_U6305 = ~new_P3_SUB_357_1258_U19 | ~new_P3_U2393;
  assign new_P3_U6306 = ~new_P3_ADD_558_U76 | ~new_P3_U3220;
  assign new_P3_U6307 = ~new_P3_ADD_553_U76 | ~new_P3_U4298;
  assign new_P3_U6308 = ~new_P3_ADD_547_U76 | ~new_P3_U4299;
  assign new_P3_U6309 = ~new_P3_ADD_541_U73 | ~new_P3_U4300;
  assign new_P3_U6310 = ~new_P3_ADD_536_U73 | ~new_P3_U4301;
  assign new_P3_U6311 = ~new_P3_ADD_531_U76 | ~new_P3_U2354;
  assign new_P3_U6312 = ~new_P3_ADD_526_U62 | ~new_P3_U2355;
  assign new_P3_U6313 = ~new_P3_ADD_515_U73 | ~new_P3_U4302;
  assign new_P3_U6314 = ~new_P3_ADD_494_U73 | ~new_P3_U2356;
  assign new_P3_U6315 = ~new_P3_ADD_476_U73 | ~new_P3_U4303;
  assign new_P3_U6316 = ~new_P3_ADD_441_U73 | ~new_P3_U4304;
  assign new_P3_U6317 = ~new_P3_ADD_405_U72 | ~new_P3_U4305;
  assign new_P3_U6318 = ~new_P3_ADD_394_U72 | ~new_P3_U2357;
  assign new_P3_U6319 = ~new_P3_ADD_385_U76 | ~new_P3_U2358;
  assign new_P3_U6320 = ~new_P3_ADD_380_U76 | ~new_P3_U2359;
  assign new_P3_U6321 = ~new_P3_ADD_349_U76 | ~new_P3_U4306;
  assign new_P3_U6322 = ~new_P3_ADD_344_U76 | ~new_P3_U2362;
  assign new_P3_U6323 = ~new_P3_ADD_371_1212_U16 | ~new_P3_U2360;
  assign new_P3_U6324 = ~new_P3_U3920 | ~new_P3_U3915 | ~new_P3_U3913 | ~new_P3_U3912 | ~new_P3_U6306;
  assign new_P3_U6325 = ~new_P3_U2402 | ~P3_REIP_REG_28_;
  assign new_P3_U6326 = ~new_P3_U4318 | ~new_P3_U6324;
  assign new_P3_U6327 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_U5631;
  assign new_P3_U6328 = ~new_P3_ADD_360_1242_U16 | ~new_P3_U2395;
  assign new_P3_U6329 = ~new_P3_SUB_357_1258_U79 | ~new_P3_U2393;
  assign new_P3_U6330 = ~new_P3_ADD_558_U75 | ~new_P3_U3220;
  assign new_P3_U6331 = ~new_P3_ADD_553_U75 | ~new_P3_U4298;
  assign new_P3_U6332 = ~new_P3_ADD_547_U75 | ~new_P3_U4299;
  assign new_P3_U6333 = ~new_P3_ADD_541_U72 | ~new_P3_U4300;
  assign new_P3_U6334 = ~new_P3_ADD_536_U72 | ~new_P3_U4301;
  assign new_P3_U6335 = ~new_P3_ADD_531_U75 | ~new_P3_U2354;
  assign new_P3_U6336 = ~new_P3_ADD_526_U61 | ~new_P3_U2355;
  assign new_P3_U6337 = ~new_P3_ADD_515_U72 | ~new_P3_U4302;
  assign new_P3_U6338 = ~new_P3_ADD_494_U72 | ~new_P3_U2356;
  assign new_P3_U6339 = ~new_P3_ADD_476_U72 | ~new_P3_U4303;
  assign new_P3_U6340 = ~new_P3_ADD_441_U72 | ~new_P3_U4304;
  assign new_P3_U6341 = ~new_P3_ADD_405_U71 | ~new_P3_U4305;
  assign new_P3_U6342 = ~new_P3_ADD_394_U71 | ~new_P3_U2357;
  assign new_P3_U6343 = ~new_P3_ADD_385_U75 | ~new_P3_U2358;
  assign new_P3_U6344 = ~new_P3_ADD_380_U75 | ~new_P3_U2359;
  assign new_P3_U6345 = ~new_P3_ADD_349_U75 | ~new_P3_U4306;
  assign new_P3_U6346 = ~new_P3_ADD_344_U75 | ~new_P3_U2362;
  assign new_P3_U6347 = ~new_P3_ADD_371_1212_U17 | ~new_P3_U2360;
  assign new_P3_U6348 = ~new_P3_U3929 | ~new_P3_U3924 | ~new_P3_U3922 | ~new_P3_U3921 | ~new_P3_U6330;
  assign new_P3_U6349 = ~new_P3_U2402 | ~P3_REIP_REG_29_;
  assign new_P3_U6350 = ~new_P3_U4318 | ~new_P3_U6348;
  assign new_P3_U6351 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_U5631;
  assign new_P3_U6352 = ~new_P3_ADD_360_1242_U77 | ~new_P3_U2395;
  assign new_P3_U6353 = ~new_P3_SUB_357_1258_U77 | ~new_P3_U2393;
  assign new_P3_U6354 = ~new_P3_ADD_558_U73 | ~new_P3_U3220;
  assign new_P3_U6355 = ~new_P3_ADD_553_U73 | ~new_P3_U4298;
  assign new_P3_U6356 = ~new_P3_ADD_547_U73 | ~new_P3_U4299;
  assign new_P3_U6357 = ~new_P3_ADD_541_U70 | ~new_P3_U4300;
  assign new_P3_U6358 = ~new_P3_ADD_536_U70 | ~new_P3_U4301;
  assign new_P3_U6359 = ~new_P3_ADD_531_U73 | ~new_P3_U2354;
  assign new_P3_U6360 = ~new_P3_ADD_526_U59 | ~new_P3_U2355;
  assign new_P3_U6361 = ~new_P3_ADD_515_U70 | ~new_P3_U4302;
  assign new_P3_U6362 = ~new_P3_ADD_494_U70 | ~new_P3_U2356;
  assign new_P3_U6363 = ~new_P3_ADD_476_U70 | ~new_P3_U4303;
  assign new_P3_U6364 = ~new_P3_ADD_441_U70 | ~new_P3_U4304;
  assign new_P3_U6365 = ~new_P3_ADD_405_U70 | ~new_P3_U4305;
  assign new_P3_U6366 = ~new_P3_ADD_394_U70 | ~new_P3_U2357;
  assign new_P3_U6367 = ~new_P3_ADD_385_U73 | ~new_P3_U2358;
  assign new_P3_U6368 = ~new_P3_ADD_380_U73 | ~new_P3_U2359;
  assign new_P3_U6369 = ~new_P3_ADD_349_U73 | ~new_P3_U4306;
  assign new_P3_U6370 = ~new_P3_ADD_344_U73 | ~new_P3_U2362;
  assign new_P3_U6371 = ~new_P3_ADD_371_1212_U79 | ~new_P3_U2360;
  assign new_P3_U6372 = ~new_P3_U3938 | ~new_P3_U3933 | ~new_P3_U3931 | ~new_P3_U3930 | ~new_P3_U6354;
  assign new_P3_U6373 = ~new_P3_U2402 | ~P3_REIP_REG_30_;
  assign new_P3_U6374 = ~new_P3_U4318 | ~new_P3_U6372;
  assign new_P3_U6375 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_U5631;
  assign new_P3_U6376 = ~new_P3_ADD_360_1242_U90 | ~new_P3_U2395;
  assign new_P3_U6377 = ~new_P3_SUB_357_1258_U20 | ~new_P3_U2393;
  assign new_P3_U6378 = ~new_P3_ADD_558_U72 | ~new_P3_U3220;
  assign new_P3_U6379 = ~new_P3_ADD_553_U72 | ~new_P3_U4298;
  assign new_P3_U6380 = ~new_P3_ADD_547_U72 | ~new_P3_U4299;
  assign new_P3_U6381 = ~new_P3_ADD_541_U69 | ~new_P3_U4300;
  assign new_P3_U6382 = ~new_P3_ADD_536_U69 | ~new_P3_U4301;
  assign new_P3_U6383 = ~new_P3_ADD_531_U72 | ~new_P3_U2354;
  assign new_P3_U6384 = ~new_P3_ADD_526_U58 | ~new_P3_U2355;
  assign new_P3_U6385 = ~new_P3_ADD_515_U69 | ~new_P3_U4302;
  assign new_P3_U6386 = ~new_P3_ADD_494_U69 | ~new_P3_U2356;
  assign new_P3_U6387 = ~new_P3_ADD_476_U69 | ~new_P3_U4303;
  assign new_P3_U6388 = ~new_P3_ADD_441_U69 | ~new_P3_U4304;
  assign new_P3_U6389 = ~new_P3_ADD_405_U69 | ~new_P3_U4305;
  assign new_P3_U6390 = ~new_P3_ADD_394_U69 | ~new_P3_U2357;
  assign new_P3_U6391 = ~new_P3_ADD_385_U72 | ~new_P3_U2358;
  assign new_P3_U6392 = ~new_P3_ADD_380_U72 | ~new_P3_U2359;
  assign new_P3_U6393 = ~new_P3_ADD_349_U72 | ~new_P3_U4306;
  assign new_P3_U6394 = ~new_P3_ADD_344_U72 | ~new_P3_U2362;
  assign new_P3_U6395 = ~new_P3_ADD_371_1212_U92 | ~new_P3_U2360;
  assign new_P3_U6396 = ~new_P3_U3950 | ~new_P3_U3945;
  assign new_P3_U6397 = ~new_P3_U2402 | ~P3_REIP_REG_31_;
  assign new_P3_U6398 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_U5631;
  assign new_P3_U6399 = ~new_P3_GTE_355_U6 | ~new_P3_U2361;
  assign new_P3_U6400 = ~new_P3_GTE_370_U6 | ~new_P3_U2360;
  assign new_P3_U6401 = ~new_P3_U6400 | ~new_P3_U6399;
  assign new_P3_U6402 = ~new_P3_U2390 | ~new_P3_U6401;
  assign new_P3_U6403 = ~new_P3_U3234 | ~new_P3_U3121;
  assign new_P3_U6404 = ~new_P3_U3249;
  assign new_P3_U6405 = ~P3_PHYADDRPOINTER_REG_0_ | ~new_P3_U2398;
  assign new_P3_U6406 = ~P3_PHYADDRPOINTER_REG_0_ | ~new_P3_U2397;
  assign new_P3_U6407 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U85;
  assign new_P3_U6408 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U69;
  assign new_P3_U6409 = ~new_P3_U2389 | ~P3_REIP_REG_0_;
  assign new_P3_U6410 = ~P3_PHYADDRPOINTER_REG_0_ | ~new_P3_U2388;
  assign new_P3_U6411 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U87;
  assign new_P3_U6412 = ~P3_PHYADDRPOINTER_REG_0_ | ~new_P3_U6404;
  assign new_P3_U6413 = ~new_P3_ADD_318_U4 | ~new_P3_U2398;
  assign new_P3_U6414 = ~P3_PHYADDRPOINTER_REG_1_ | ~new_P3_U2397;
  assign new_P3_U6415 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U19;
  assign new_P3_U6416 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U21;
  assign new_P3_U6417 = ~new_P3_U2389 | ~P3_REIP_REG_1_;
  assign new_P3_U6418 = ~new_P3_ADD_339_U4 | ~new_P3_U2388;
  assign new_P3_U6419 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U20;
  assign new_P3_U6420 = ~P3_PHYADDRPOINTER_REG_1_ | ~new_P3_U6404;
  assign new_P3_U6421 = ~new_P3_ADD_318_U71 | ~new_P3_U2398;
  assign new_P3_U6422 = ~new_P3_ADD_315_U4 | ~new_P3_U2397;
  assign new_P3_U6423 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U91;
  assign new_P3_U6424 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U78;
  assign new_P3_U6425 = ~new_P3_U2389 | ~P3_REIP_REG_2_;
  assign new_P3_U6426 = ~new_P3_ADD_339_U71 | ~new_P3_U2388;
  assign new_P3_U6427 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U93;
  assign new_P3_U6428 = ~P3_PHYADDRPOINTER_REG_2_ | ~new_P3_U6404;
  assign new_P3_U6429 = ~new_P3_ADD_318_U68 | ~new_P3_U2398;
  assign new_P3_U6430 = ~new_P3_ADD_315_U66 | ~new_P3_U2397;
  assign new_P3_U6431 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U17;
  assign new_P3_U6432 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U76;
  assign new_P3_U6433 = ~new_P3_U2389 | ~P3_REIP_REG_3_;
  assign new_P3_U6434 = ~new_P3_ADD_339_U68 | ~new_P3_U2388;
  assign new_P3_U6435 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U18;
  assign new_P3_U6436 = ~P3_PHYADDRPOINTER_REG_3_ | ~new_P3_U6404;
  assign new_P3_U6437 = ~new_P3_ADD_318_U67 | ~new_P3_U2398;
  assign new_P3_U6438 = ~new_P3_ADD_315_U65 | ~new_P3_U2397;
  assign new_P3_U6439 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U18;
  assign new_P3_U6440 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U75;
  assign new_P3_U6441 = ~new_P3_U2389 | ~P3_REIP_REG_4_;
  assign new_P3_U6442 = ~new_P3_ADD_339_U67 | ~new_P3_U2388;
  assign new_P3_U6443 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U91;
  assign new_P3_U6444 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_U6404;
  assign new_P3_U6445 = ~new_P3_ADD_318_U66 | ~new_P3_U2398;
  assign new_P3_U6446 = ~new_P3_ADD_315_U64 | ~new_P3_U2397;
  assign new_P3_U6447 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U89;
  assign new_P3_U6448 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U74;
  assign new_P3_U6449 = ~new_P3_U2389 | ~P3_REIP_REG_5_;
  assign new_P3_U6450 = ~new_P3_ADD_339_U66 | ~new_P3_U2388;
  assign new_P3_U6451 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U19;
  assign new_P3_U6452 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_U6404;
  assign new_P3_U6453 = ~new_P3_ADD_318_U65 | ~new_P3_U2398;
  assign new_P3_U6454 = ~new_P3_ADD_315_U63 | ~new_P3_U2397;
  assign new_P3_U6455 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U88;
  assign new_P3_U6456 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U73;
  assign new_P3_U6457 = ~new_P3_U2389 | ~P3_REIP_REG_6_;
  assign new_P3_U6458 = ~new_P3_ADD_339_U65 | ~new_P3_U2388;
  assign new_P3_U6459 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U90;
  assign new_P3_U6460 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_U6404;
  assign new_P3_U6461 = ~new_P3_ADD_318_U64 | ~new_P3_U2398;
  assign new_P3_U6462 = ~new_P3_ADD_315_U62 | ~new_P3_U2397;
  assign new_P3_U6463 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U87;
  assign new_P3_U6464 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U72;
  assign new_P3_U6465 = ~new_P3_U2389 | ~P3_REIP_REG_7_;
  assign new_P3_U6466 = ~new_P3_ADD_339_U64 | ~new_P3_U2388;
  assign new_P3_U6467 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U89;
  assign new_P3_U6468 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_U6404;
  assign new_P3_U6469 = ~new_P3_ADD_318_U63 | ~new_P3_U2398;
  assign new_P3_U6470 = ~new_P3_ADD_315_U61 | ~new_P3_U2397;
  assign new_P3_U6471 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U86;
  assign new_P3_U6472 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U71;
  assign new_P3_U6473 = ~new_P3_U2389 | ~P3_REIP_REG_8_;
  assign new_P3_U6474 = ~new_P3_ADD_339_U63 | ~new_P3_U2388;
  assign new_P3_U6475 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U88;
  assign new_P3_U6476 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_U6404;
  assign new_P3_U6477 = ~new_P3_ADD_318_U62 | ~new_P3_U2398;
  assign new_P3_U6478 = ~new_P3_ADD_315_U60 | ~new_P3_U2397;
  assign new_P3_U6479 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U106;
  assign new_P3_U6480 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U70;
  assign new_P3_U6481 = ~new_P3_U2389 | ~P3_REIP_REG_9_;
  assign new_P3_U6482 = ~new_P3_ADD_339_U62 | ~new_P3_U2388;
  assign new_P3_U6483 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U109;
  assign new_P3_U6484 = ~P3_PHYADDRPOINTER_REG_9_ | ~new_P3_U6404;
  assign new_P3_U6485 = ~new_P3_ADD_318_U91 | ~new_P3_U2398;
  assign new_P3_U6486 = ~new_P3_ADD_315_U88 | ~new_P3_U2397;
  assign new_P3_U6487 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U4;
  assign new_P3_U6488 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U93;
  assign new_P3_U6489 = ~new_P3_U2389 | ~P3_REIP_REG_10_;
  assign new_P3_U6490 = ~new_P3_ADD_339_U91 | ~new_P3_U2388;
  assign new_P3_U6491 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U5;
  assign new_P3_U6492 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_U6404;
  assign new_P3_U6493 = ~new_P3_ADD_318_U90 | ~new_P3_U2398;
  assign new_P3_U6494 = ~new_P3_ADD_315_U87 | ~new_P3_U2397;
  assign new_P3_U6495 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U84;
  assign new_P3_U6496 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U92;
  assign new_P3_U6497 = ~new_P3_U2389 | ~P3_REIP_REG_11_;
  assign new_P3_U6498 = ~new_P3_ADD_339_U90 | ~new_P3_U2388;
  assign new_P3_U6499 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U86;
  assign new_P3_U6500 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_U6404;
  assign new_P3_U6501 = ~new_P3_ADD_318_U89 | ~new_P3_U2398;
  assign new_P3_U6502 = ~new_P3_ADD_315_U86 | ~new_P3_U2397;
  assign new_P3_U6503 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U5;
  assign new_P3_U6504 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U91;
  assign new_P3_U6505 = ~new_P3_U2389 | ~P3_REIP_REG_12_;
  assign new_P3_U6506 = ~new_P3_ADD_339_U89 | ~new_P3_U2388;
  assign new_P3_U6507 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U6;
  assign new_P3_U6508 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_U6404;
  assign new_P3_U6509 = ~new_P3_ADD_318_U88 | ~new_P3_U2398;
  assign new_P3_U6510 = ~new_P3_ADD_315_U85 | ~new_P3_U2397;
  assign new_P3_U6511 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U6;
  assign new_P3_U6512 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U15;
  assign new_P3_U6513 = ~new_P3_U2389 | ~P3_REIP_REG_13_;
  assign new_P3_U6514 = ~new_P3_ADD_339_U88 | ~new_P3_U2388;
  assign new_P3_U6515 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U7;
  assign new_P3_U6516 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_U6404;
  assign new_P3_U6517 = ~new_P3_ADD_318_U87 | ~new_P3_U2398;
  assign new_P3_U6518 = ~new_P3_ADD_315_U84 | ~new_P3_U2397;
  assign new_P3_U6519 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U83;
  assign new_P3_U6520 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U90;
  assign new_P3_U6521 = ~new_P3_U2389 | ~P3_REIP_REG_14_;
  assign new_P3_U6522 = ~new_P3_ADD_339_U87 | ~new_P3_U2388;
  assign new_P3_U6523 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U85;
  assign new_P3_U6524 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_U6404;
  assign new_P3_U6525 = ~new_P3_ADD_318_U86 | ~new_P3_U2398;
  assign new_P3_U6526 = ~new_P3_ADD_315_U83 | ~new_P3_U2397;
  assign new_P3_U6527 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U7;
  assign new_P3_U6528 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U89;
  assign new_P3_U6529 = ~new_P3_U2389 | ~P3_REIP_REG_15_;
  assign new_P3_U6530 = ~new_P3_ADD_339_U86 | ~new_P3_U2388;
  assign new_P3_U6531 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U8;
  assign new_P3_U6532 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_U6404;
  assign new_P3_U6533 = ~new_P3_ADD_318_U85 | ~new_P3_U2398;
  assign new_P3_U6534 = ~new_P3_ADD_315_U82 | ~new_P3_U2397;
  assign new_P3_U6535 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U82;
  assign new_P3_U6536 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U88;
  assign new_P3_U6537 = ~new_P3_U2389 | ~P3_REIP_REG_16_;
  assign new_P3_U6538 = ~new_P3_ADD_339_U85 | ~new_P3_U2388;
  assign new_P3_U6539 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U84;
  assign new_P3_U6540 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_U6404;
  assign new_P3_U6541 = ~new_P3_ADD_318_U84 | ~new_P3_U2398;
  assign new_P3_U6542 = ~new_P3_ADD_315_U81 | ~new_P3_U2397;
  assign new_P3_U6543 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U8;
  assign new_P3_U6544 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U16;
  assign new_P3_U6545 = ~new_P3_U2389 | ~P3_REIP_REG_17_;
  assign new_P3_U6546 = ~new_P3_ADD_339_U84 | ~new_P3_U2388;
  assign new_P3_U6547 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U9;
  assign new_P3_U6548 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_U6404;
  assign new_P3_U6549 = ~new_P3_ADD_318_U83 | ~new_P3_U2398;
  assign new_P3_U6550 = ~new_P3_ADD_315_U80 | ~new_P3_U2397;
  assign new_P3_U6551 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U81;
  assign new_P3_U6552 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U87;
  assign new_P3_U6553 = ~new_P3_U2389 | ~P3_REIP_REG_18_;
  assign new_P3_U6554 = ~new_P3_ADD_339_U83 | ~new_P3_U2388;
  assign new_P3_U6555 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U83;
  assign new_P3_U6556 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_U6404;
  assign new_P3_U6557 = ~new_P3_ADD_318_U82 | ~new_P3_U2398;
  assign new_P3_U6558 = ~new_P3_ADD_315_U79 | ~new_P3_U2397;
  assign new_P3_U6559 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U9;
  assign new_P3_U6560 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U86;
  assign new_P3_U6561 = ~new_P3_U2389 | ~P3_REIP_REG_19_;
  assign new_P3_U6562 = ~new_P3_ADD_339_U82 | ~new_P3_U2388;
  assign new_P3_U6563 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U10;
  assign new_P3_U6564 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_U6404;
  assign new_P3_U6565 = ~new_P3_ADD_318_U81 | ~new_P3_U2398;
  assign new_P3_U6566 = ~new_P3_ADD_315_U78 | ~new_P3_U2397;
  assign new_P3_U6567 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U10;
  assign new_P3_U6568 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U17;
  assign new_P3_U6569 = ~new_P3_U2389 | ~P3_REIP_REG_20_;
  assign new_P3_U6570 = ~new_P3_ADD_339_U81 | ~new_P3_U2388;
  assign new_P3_U6571 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U11;
  assign new_P3_U6572 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_U6404;
  assign new_P3_U6573 = ~new_P3_ADD_318_U80 | ~new_P3_U2398;
  assign new_P3_U6574 = ~new_P3_ADD_315_U77 | ~new_P3_U2397;
  assign new_P3_U6575 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U11;
  assign new_P3_U6576 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U85;
  assign new_P3_U6577 = ~new_P3_U2389 | ~P3_REIP_REG_21_;
  assign new_P3_U6578 = ~new_P3_ADD_339_U80 | ~new_P3_U2388;
  assign new_P3_U6579 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U12;
  assign new_P3_U6580 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_U6404;
  assign new_P3_U6581 = ~new_P3_ADD_318_U79 | ~new_P3_U2398;
  assign new_P3_U6582 = ~new_P3_ADD_315_U76 | ~new_P3_U2397;
  assign new_P3_U6583 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U80;
  assign new_P3_U6584 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U84;
  assign new_P3_U6585 = ~new_P3_U2389 | ~P3_REIP_REG_22_;
  assign new_P3_U6586 = ~new_P3_ADD_339_U79 | ~new_P3_U2388;
  assign new_P3_U6587 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U82;
  assign new_P3_U6588 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_U6404;
  assign new_P3_U6589 = ~new_P3_ADD_318_U78 | ~new_P3_U2398;
  assign new_P3_U6590 = ~new_P3_ADD_315_U75 | ~new_P3_U2397;
  assign new_P3_U6591 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U12;
  assign new_P3_U6592 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U83;
  assign new_P3_U6593 = ~new_P3_U2389 | ~P3_REIP_REG_23_;
  assign new_P3_U6594 = ~new_P3_ADD_339_U78 | ~new_P3_U2388;
  assign new_P3_U6595 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U13;
  assign new_P3_U6596 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_U6404;
  assign new_P3_U6597 = ~new_P3_ADD_318_U77 | ~new_P3_U2398;
  assign new_P3_U6598 = ~new_P3_ADD_315_U74 | ~new_P3_U2397;
  assign new_P3_U6599 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U79;
  assign new_P3_U6600 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U82;
  assign new_P3_U6601 = ~new_P3_U2389 | ~P3_REIP_REG_24_;
  assign new_P3_U6602 = ~new_P3_ADD_339_U77 | ~new_P3_U2388;
  assign new_P3_U6603 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U81;
  assign new_P3_U6604 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_U6404;
  assign new_P3_U6605 = ~new_P3_ADD_318_U76 | ~new_P3_U2398;
  assign new_P3_U6606 = ~new_P3_ADD_315_U73 | ~new_P3_U2397;
  assign new_P3_U6607 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U13;
  assign new_P3_U6608 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U81;
  assign new_P3_U6609 = ~new_P3_U2389 | ~P3_REIP_REG_25_;
  assign new_P3_U6610 = ~new_P3_ADD_339_U76 | ~new_P3_U2388;
  assign new_P3_U6611 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U14;
  assign new_P3_U6612 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_U6404;
  assign new_P3_U6613 = ~new_P3_ADD_318_U75 | ~new_P3_U2398;
  assign new_P3_U6614 = ~new_P3_ADD_315_U72 | ~new_P3_U2397;
  assign new_P3_U6615 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U14;
  assign new_P3_U6616 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U18;
  assign new_P3_U6617 = ~new_P3_U2389 | ~P3_REIP_REG_26_;
  assign new_P3_U6618 = ~new_P3_ADD_339_U75 | ~new_P3_U2388;
  assign new_P3_U6619 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U15;
  assign new_P3_U6620 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_U6404;
  assign new_P3_U6621 = ~new_P3_ADD_318_U74 | ~new_P3_U2398;
  assign new_P3_U6622 = ~new_P3_ADD_315_U71 | ~new_P3_U2397;
  assign new_P3_U6623 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U78;
  assign new_P3_U6624 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U80;
  assign new_P3_U6625 = ~new_P3_U2389 | ~P3_REIP_REG_27_;
  assign new_P3_U6626 = ~new_P3_ADD_339_U74 | ~new_P3_U2388;
  assign new_P3_U6627 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U80;
  assign new_P3_U6628 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_U6404;
  assign new_P3_U6629 = ~new_P3_ADD_318_U73 | ~new_P3_U2398;
  assign new_P3_U6630 = ~new_P3_ADD_315_U70 | ~new_P3_U2397;
  assign new_P3_U6631 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U15;
  assign new_P3_U6632 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U19;
  assign new_P3_U6633 = ~new_P3_U2389 | ~P3_REIP_REG_28_;
  assign new_P3_U6634 = ~new_P3_ADD_339_U73 | ~new_P3_U2388;
  assign new_P3_U6635 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U16;
  assign new_P3_U6636 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_U6404;
  assign new_P3_U6637 = ~new_P3_ADD_318_U72 | ~new_P3_U2398;
  assign new_P3_U6638 = ~new_P3_ADD_315_U69 | ~new_P3_U2397;
  assign new_P3_U6639 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U16;
  assign new_P3_U6640 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U79;
  assign new_P3_U6641 = ~new_P3_U2389 | ~P3_REIP_REG_29_;
  assign new_P3_U6642 = ~new_P3_ADD_339_U72 | ~new_P3_U2388;
  assign new_P3_U6643 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U17;
  assign new_P3_U6644 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_U6404;
  assign new_P3_U6645 = ~new_P3_ADD_318_U70 | ~new_P3_U2398;
  assign new_P3_U6646 = ~new_P3_ADD_315_U68 | ~new_P3_U2397;
  assign new_P3_U6647 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U77;
  assign new_P3_U6648 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U77;
  assign new_P3_U6649 = ~new_P3_U2389 | ~P3_REIP_REG_30_;
  assign new_P3_U6650 = ~new_P3_ADD_339_U70 | ~new_P3_U2388;
  assign new_P3_U6651 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U79;
  assign new_P3_U6652 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_U6404;
  assign new_P3_U6653 = ~new_P3_ADD_318_U69 | ~new_P3_U2398;
  assign new_P3_U6654 = ~new_P3_ADD_315_U67 | ~new_P3_U2397;
  assign new_P3_U6655 = ~new_P3_U2396 | ~new_P3_ADD_360_1242_U90;
  assign new_P3_U6656 = ~new_P3_U2394 | ~new_P3_SUB_357_1258_U20;
  assign new_P3_U6657 = ~new_P3_U2389 | ~P3_REIP_REG_31_;
  assign new_P3_U6658 = ~new_P3_ADD_339_U69 | ~new_P3_U2388;
  assign new_P3_U6659 = ~new_P3_U2387 | ~new_P3_ADD_371_1212_U92;
  assign new_P3_U6660 = ~P3_PHYADDRPOINTER_REG_31_ | ~new_P3_U6404;
  assign new_P3_U6661 = ~new_P3_GTE_412_U6 | ~new_P3_U4304 | ~new_P3_U2630;
  assign new_P3_U6662 = ~new_P3_GTE_450_U6 | ~new_P3_U4303;
  assign new_P3_U6663 = ~new_P3_U6662 | ~new_P3_U6661;
  assign new_P3_U6664 = ~P3_EAX_REG_15_ | ~new_P3_U2407;
  assign new_P3_U6665 = ~BUF2_REG_15_ | ~new_P3_U2406;
  assign new_P3_U6666 = ~P3_LWORD_REG_15_ | ~new_P3_U3250;
  assign new_P3_U6667 = ~P3_EAX_REG_14_ | ~new_P3_U2407;
  assign new_P3_U6668 = ~BUF2_REG_14_ | ~new_P3_U2406;
  assign new_P3_U6669 = ~P3_LWORD_REG_14_ | ~new_P3_U3250;
  assign new_P3_U6670 = ~P3_EAX_REG_13_ | ~new_P3_U2407;
  assign new_P3_U6671 = ~BUF2_REG_13_ | ~new_P3_U2406;
  assign new_P3_U6672 = ~P3_LWORD_REG_13_ | ~new_P3_U3250;
  assign new_P3_U6673 = ~P3_EAX_REG_12_ | ~new_P3_U2407;
  assign new_P3_U6674 = ~BUF2_REG_12_ | ~new_P3_U2406;
  assign new_P3_U6675 = ~P3_LWORD_REG_12_ | ~new_P3_U3250;
  assign new_P3_U6676 = ~P3_EAX_REG_11_ | ~new_P3_U2407;
  assign new_P3_U6677 = ~BUF2_REG_11_ | ~new_P3_U2406;
  assign new_P3_U6678 = ~P3_LWORD_REG_11_ | ~new_P3_U3250;
  assign new_P3_U6679 = ~P3_EAX_REG_10_ | ~new_P3_U2407;
  assign new_P3_U6680 = ~BUF2_REG_10_ | ~new_P3_U2406;
  assign new_P3_U6681 = ~P3_LWORD_REG_10_ | ~new_P3_U3250;
  assign new_P3_U6682 = ~P3_EAX_REG_9_ | ~new_P3_U2407;
  assign new_P3_U6683 = ~BUF2_REG_9_ | ~new_P3_U2406;
  assign new_P3_U6684 = ~P3_LWORD_REG_9_ | ~new_P3_U3250;
  assign new_P3_U6685 = ~P3_EAX_REG_8_ | ~new_P3_U2407;
  assign new_P3_U6686 = ~BUF2_REG_8_ | ~new_P3_U2406;
  assign new_P3_U6687 = ~P3_LWORD_REG_8_ | ~new_P3_U3250;
  assign new_P3_U6688 = ~P3_EAX_REG_7_ | ~new_P3_U2407;
  assign new_P3_U6689 = ~new_P3_U2406 | ~BUF2_REG_7_;
  assign new_P3_U6690 = ~P3_LWORD_REG_7_ | ~new_P3_U3250;
  assign new_P3_U6691 = ~P3_EAX_REG_6_ | ~new_P3_U2407;
  assign new_P3_U6692 = ~new_P3_U2406 | ~BUF2_REG_6_;
  assign new_P3_U6693 = ~P3_LWORD_REG_6_ | ~new_P3_U3250;
  assign new_P3_U6694 = ~P3_EAX_REG_5_ | ~new_P3_U2407;
  assign new_P3_U6695 = ~new_P3_U2406 | ~BUF2_REG_5_;
  assign new_P3_U6696 = ~P3_LWORD_REG_5_ | ~new_P3_U3250;
  assign new_P3_U6697 = ~P3_EAX_REG_4_ | ~new_P3_U2407;
  assign new_P3_U6698 = ~new_P3_U2406 | ~BUF2_REG_4_;
  assign new_P3_U6699 = ~P3_LWORD_REG_4_ | ~new_P3_U3250;
  assign new_P3_U6700 = ~P3_EAX_REG_3_ | ~new_P3_U2407;
  assign new_P3_U6701 = ~new_P3_U2406 | ~BUF2_REG_3_;
  assign new_P3_U6702 = ~P3_LWORD_REG_3_ | ~new_P3_U3250;
  assign new_P3_U6703 = ~P3_EAX_REG_2_ | ~new_P3_U2407;
  assign new_P3_U6704 = ~new_P3_U2406 | ~BUF2_REG_2_;
  assign new_P3_U6705 = ~P3_LWORD_REG_2_ | ~new_P3_U3250;
  assign new_P3_U6706 = ~P3_EAX_REG_1_ | ~new_P3_U2407;
  assign new_P3_U6707 = ~new_P3_U2406 | ~BUF2_REG_1_;
  assign new_P3_U6708 = ~P3_LWORD_REG_1_ | ~new_P3_U3250;
  assign new_P3_U6709 = ~P3_EAX_REG_0_ | ~new_P3_U2407;
  assign new_P3_U6710 = ~new_P3_U2406 | ~BUF2_REG_0_;
  assign new_P3_U6711 = ~P3_LWORD_REG_0_ | ~new_P3_U3250;
  assign new_P3_U6712 = ~P3_EAX_REG_30_ | ~new_P3_U2407;
  assign new_P3_U6713 = ~BUF2_REG_14_ | ~new_P3_U2406;
  assign new_P3_U6714 = ~P3_UWORD_REG_14_ | ~new_P3_U3250;
  assign new_P3_U6715 = ~P3_EAX_REG_29_ | ~new_P3_U2407;
  assign new_P3_U6716 = ~BUF2_REG_13_ | ~new_P3_U2406;
  assign new_P3_U6717 = ~P3_UWORD_REG_13_ | ~new_P3_U3250;
  assign new_P3_U6718 = ~P3_EAX_REG_28_ | ~new_P3_U2407;
  assign new_P3_U6719 = ~BUF2_REG_12_ | ~new_P3_U2406;
  assign new_P3_U6720 = ~P3_UWORD_REG_12_ | ~new_P3_U3250;
  assign new_P3_U6721 = ~P3_EAX_REG_27_ | ~new_P3_U2407;
  assign new_P3_U6722 = ~BUF2_REG_11_ | ~new_P3_U2406;
  assign new_P3_U6723 = ~P3_UWORD_REG_11_ | ~new_P3_U3250;
  assign new_P3_U6724 = ~P3_EAX_REG_26_ | ~new_P3_U2407;
  assign new_P3_U6725 = ~BUF2_REG_10_ | ~new_P3_U2406;
  assign new_P3_U6726 = ~P3_UWORD_REG_10_ | ~new_P3_U3250;
  assign new_P3_U6727 = ~P3_EAX_REG_25_ | ~new_P3_U2407;
  assign new_P3_U6728 = ~BUF2_REG_9_ | ~new_P3_U2406;
  assign new_P3_U6729 = ~P3_UWORD_REG_9_ | ~new_P3_U3250;
  assign new_P3_U6730 = ~P3_EAX_REG_24_ | ~new_P3_U2407;
  assign new_P3_U6731 = ~BUF2_REG_8_ | ~new_P3_U2406;
  assign new_P3_U6732 = ~P3_UWORD_REG_8_ | ~new_P3_U3250;
  assign new_P3_U6733 = ~P3_EAX_REG_23_ | ~new_P3_U2407;
  assign new_P3_U6734 = ~new_P3_U2406 | ~BUF2_REG_7_;
  assign new_P3_U6735 = ~P3_UWORD_REG_7_ | ~new_P3_U3250;
  assign new_P3_U6736 = ~P3_EAX_REG_22_ | ~new_P3_U2407;
  assign new_P3_U6737 = ~new_P3_U2406 | ~BUF2_REG_6_;
  assign new_P3_U6738 = ~P3_UWORD_REG_6_ | ~new_P3_U3250;
  assign new_P3_U6739 = ~P3_EAX_REG_21_ | ~new_P3_U2407;
  assign new_P3_U6740 = ~new_P3_U2406 | ~BUF2_REG_5_;
  assign new_P3_U6741 = ~P3_UWORD_REG_5_ | ~new_P3_U3250;
  assign new_P3_U6742 = ~P3_EAX_REG_20_ | ~new_P3_U2407;
  assign new_P3_U6743 = ~new_P3_U2406 | ~BUF2_REG_4_;
  assign new_P3_U6744 = ~P3_UWORD_REG_4_ | ~new_P3_U3250;
  assign new_P3_U6745 = ~P3_EAX_REG_19_ | ~new_P3_U2407;
  assign new_P3_U6746 = ~new_P3_U2406 | ~BUF2_REG_3_;
  assign new_P3_U6747 = ~P3_UWORD_REG_3_ | ~new_P3_U3250;
  assign new_P3_U6748 = ~P3_EAX_REG_18_ | ~new_P3_U2407;
  assign new_P3_U6749 = ~new_P3_U2406 | ~BUF2_REG_2_;
  assign new_P3_U6750 = ~P3_UWORD_REG_2_ | ~new_P3_U3250;
  assign new_P3_U6751 = ~P3_EAX_REG_17_ | ~new_P3_U2407;
  assign new_P3_U6752 = ~new_P3_U2406 | ~BUF2_REG_1_;
  assign new_P3_U6753 = ~P3_UWORD_REG_1_ | ~new_P3_U3250;
  assign new_P3_U6754 = ~P3_EAX_REG_16_ | ~new_P3_U2407;
  assign new_P3_U6755 = ~new_P3_U2406 | ~BUF2_REG_0_;
  assign new_P3_U6756 = ~P3_UWORD_REG_0_ | ~new_P3_U3250;
  assign new_P3_U6757 = ~new_P3_U3986 | ~new_P3_U3255;
  assign new_P3_U6758 = ~new_P3_U2453 | ~new_P3_U3121;
  assign new_P3_U6759 = ~new_P3_U3251;
  assign new_P3_U6760 = ~new_P3_U2410 | ~P3_LWORD_REG_0_;
  assign new_P3_U6761 = ~new_P3_U2409 | ~P3_EAX_REG_0_;
  assign new_P3_U6762 = ~P3_DATAO_REG_0_ | ~new_P3_U6759;
  assign new_P3_U6763 = ~new_P3_U2410 | ~P3_LWORD_REG_1_;
  assign new_P3_U6764 = ~new_P3_U2409 | ~P3_EAX_REG_1_;
  assign new_P3_U6765 = ~P3_DATAO_REG_1_ | ~new_P3_U6759;
  assign new_P3_U6766 = ~new_P3_U2410 | ~P3_LWORD_REG_2_;
  assign new_P3_U6767 = ~new_P3_U2409 | ~P3_EAX_REG_2_;
  assign new_P3_U6768 = ~P3_DATAO_REG_2_ | ~new_P3_U6759;
  assign new_P3_U6769 = ~new_P3_U2410 | ~P3_LWORD_REG_3_;
  assign new_P3_U6770 = ~new_P3_U2409 | ~P3_EAX_REG_3_;
  assign new_P3_U6771 = ~P3_DATAO_REG_3_ | ~new_P3_U6759;
  assign new_P3_U6772 = ~new_P3_U2410 | ~P3_LWORD_REG_4_;
  assign new_P3_U6773 = ~new_P3_U2409 | ~P3_EAX_REG_4_;
  assign new_P3_U6774 = ~P3_DATAO_REG_4_ | ~new_P3_U6759;
  assign new_P3_U6775 = ~new_P3_U2410 | ~P3_LWORD_REG_5_;
  assign new_P3_U6776 = ~new_P3_U2409 | ~P3_EAX_REG_5_;
  assign new_P3_U6777 = ~P3_DATAO_REG_5_ | ~new_P3_U6759;
  assign new_P3_U6778 = ~new_P3_U2410 | ~P3_LWORD_REG_6_;
  assign new_P3_U6779 = ~new_P3_U2409 | ~P3_EAX_REG_6_;
  assign new_P3_U6780 = ~P3_DATAO_REG_6_ | ~new_P3_U6759;
  assign new_P3_U6781 = ~new_P3_U2410 | ~P3_LWORD_REG_7_;
  assign new_P3_U6782 = ~new_P3_U2409 | ~P3_EAX_REG_7_;
  assign new_P3_U6783 = ~P3_DATAO_REG_7_ | ~new_P3_U6759;
  assign new_P3_U6784 = ~new_P3_U2410 | ~P3_LWORD_REG_8_;
  assign new_P3_U6785 = ~new_P3_U2409 | ~P3_EAX_REG_8_;
  assign new_P3_U6786 = ~P3_DATAO_REG_8_ | ~new_P3_U6759;
  assign new_P3_U6787 = ~new_P3_U2410 | ~P3_LWORD_REG_9_;
  assign new_P3_U6788 = ~new_P3_U2409 | ~P3_EAX_REG_9_;
  assign new_P3_U6789 = ~P3_DATAO_REG_9_ | ~new_P3_U6759;
  assign new_P3_U6790 = ~new_P3_U2410 | ~P3_LWORD_REG_10_;
  assign new_P3_U6791 = ~new_P3_U2409 | ~P3_EAX_REG_10_;
  assign new_P3_U6792 = ~P3_DATAO_REG_10_ | ~new_P3_U6759;
  assign new_P3_U6793 = ~new_P3_U2410 | ~P3_LWORD_REG_11_;
  assign new_P3_U6794 = ~new_P3_U2409 | ~P3_EAX_REG_11_;
  assign new_P3_U6795 = ~P3_DATAO_REG_11_ | ~new_P3_U6759;
  assign new_P3_U6796 = ~new_P3_U2410 | ~P3_LWORD_REG_12_;
  assign new_P3_U6797 = ~new_P3_U2409 | ~P3_EAX_REG_12_;
  assign new_P3_U6798 = ~P3_DATAO_REG_12_ | ~new_P3_U6759;
  assign new_P3_U6799 = ~new_P3_U2410 | ~P3_LWORD_REG_13_;
  assign new_P3_U6800 = ~new_P3_U2409 | ~P3_EAX_REG_13_;
  assign new_P3_U6801 = ~P3_DATAO_REG_13_ | ~new_P3_U6759;
  assign new_P3_U6802 = ~new_P3_U2410 | ~P3_LWORD_REG_14_;
  assign new_P3_U6803 = ~new_P3_U2409 | ~P3_EAX_REG_14_;
  assign new_P3_U6804 = ~P3_DATAO_REG_14_ | ~new_P3_U6759;
  assign new_P3_U6805 = ~new_P3_U2410 | ~P3_LWORD_REG_15_;
  assign new_P3_U6806 = ~new_P3_U2409 | ~P3_EAX_REG_15_;
  assign new_P3_U6807 = ~P3_DATAO_REG_15_ | ~new_P3_U6759;
  assign new_P3_U6808 = ~new_P3_U2447 | ~P3_EAX_REG_16_;
  assign new_P3_U6809 = ~new_P3_U2410 | ~P3_UWORD_REG_0_;
  assign new_P3_U6810 = ~P3_DATAO_REG_16_ | ~new_P3_U6759;
  assign new_P3_U6811 = ~new_P3_U2447 | ~P3_EAX_REG_17_;
  assign new_P3_U6812 = ~new_P3_U2410 | ~P3_UWORD_REG_1_;
  assign new_P3_U6813 = ~P3_DATAO_REG_17_ | ~new_P3_U6759;
  assign new_P3_U6814 = ~new_P3_U2447 | ~P3_EAX_REG_18_;
  assign new_P3_U6815 = ~new_P3_U2410 | ~P3_UWORD_REG_2_;
  assign new_P3_U6816 = ~P3_DATAO_REG_18_ | ~new_P3_U6759;
  assign new_P3_U6817 = ~new_P3_U2447 | ~P3_EAX_REG_19_;
  assign new_P3_U6818 = ~new_P3_U2410 | ~P3_UWORD_REG_3_;
  assign new_P3_U6819 = ~P3_DATAO_REG_19_ | ~new_P3_U6759;
  assign new_P3_U6820 = ~new_P3_U2447 | ~P3_EAX_REG_20_;
  assign new_P3_U6821 = ~new_P3_U2410 | ~P3_UWORD_REG_4_;
  assign new_P3_U6822 = ~P3_DATAO_REG_20_ | ~new_P3_U6759;
  assign new_P3_U6823 = ~new_P3_U2447 | ~P3_EAX_REG_21_;
  assign new_P3_U6824 = ~new_P3_U2410 | ~P3_UWORD_REG_5_;
  assign new_P3_U6825 = ~P3_DATAO_REG_21_ | ~new_P3_U6759;
  assign new_P3_U6826 = ~new_P3_U2447 | ~P3_EAX_REG_22_;
  assign new_P3_U6827 = ~new_P3_U2410 | ~P3_UWORD_REG_6_;
  assign new_P3_U6828 = ~P3_DATAO_REG_22_ | ~new_P3_U6759;
  assign new_P3_U6829 = ~new_P3_U2447 | ~P3_EAX_REG_23_;
  assign new_P3_U6830 = ~new_P3_U2410 | ~P3_UWORD_REG_7_;
  assign new_P3_U6831 = ~P3_DATAO_REG_23_ | ~new_P3_U6759;
  assign new_P3_U6832 = ~new_P3_U2447 | ~P3_EAX_REG_24_;
  assign new_P3_U6833 = ~new_P3_U2410 | ~P3_UWORD_REG_8_;
  assign new_P3_U6834 = ~P3_DATAO_REG_24_ | ~new_P3_U6759;
  assign new_P3_U6835 = ~new_P3_U2447 | ~P3_EAX_REG_25_;
  assign new_P3_U6836 = ~new_P3_U2410 | ~P3_UWORD_REG_9_;
  assign new_P3_U6837 = ~P3_DATAO_REG_25_ | ~new_P3_U6759;
  assign new_P3_U6838 = ~new_P3_U2447 | ~P3_EAX_REG_26_;
  assign new_P3_U6839 = ~new_P3_U2410 | ~P3_UWORD_REG_10_;
  assign new_P3_U6840 = ~P3_DATAO_REG_26_ | ~new_P3_U6759;
  assign new_P3_U6841 = ~new_P3_U2447 | ~P3_EAX_REG_27_;
  assign new_P3_U6842 = ~new_P3_U2410 | ~P3_UWORD_REG_11_;
  assign new_P3_U6843 = ~P3_DATAO_REG_27_ | ~new_P3_U6759;
  assign new_P3_U6844 = ~new_P3_U2447 | ~P3_EAX_REG_28_;
  assign new_P3_U6845 = ~new_P3_U2410 | ~P3_UWORD_REG_12_;
  assign new_P3_U6846 = ~P3_DATAO_REG_28_ | ~new_P3_U6759;
  assign new_P3_U6847 = ~new_P3_U2447 | ~P3_EAX_REG_29_;
  assign new_P3_U6848 = ~new_P3_U2410 | ~P3_UWORD_REG_13_;
  assign new_P3_U6849 = ~P3_DATAO_REG_29_ | ~new_P3_U6759;
  assign new_P3_U6850 = ~new_P3_U2447 | ~P3_EAX_REG_30_;
  assign new_P3_U6851 = ~new_P3_U2410 | ~P3_UWORD_REG_14_;
  assign new_P3_U6852 = ~P3_DATAO_REG_30_ | ~new_P3_U6759;
  assign new_P3_U6853 = ~new_P3_U2516 | ~new_P3_U3243;
  assign new_P3_U6854 = ~new_P3_U2446 | ~BUF2_REG_0_;
  assign new_P3_U6855 = ~new_P3_U2621 | ~new_P3_U2411;
  assign new_P3_U6856 = ~new_P3_ADD_546_U5 | ~new_P3_U2400;
  assign new_P3_U6857 = ~P3_EAX_REG_0_ | ~new_P3_U3252;
  assign new_P3_U6858 = ~new_P3_U2446 | ~BUF2_REG_1_;
  assign new_P3_U6859 = ~new_P3_U2622 | ~new_P3_U2411;
  assign new_P3_U6860 = ~new_P3_ADD_546_U71 | ~new_P3_U2400;
  assign new_P3_U6861 = ~P3_EAX_REG_1_ | ~new_P3_U3252;
  assign new_P3_U6862 = ~new_P3_U2446 | ~BUF2_REG_2_;
  assign new_P3_U6863 = ~new_P3_U2623 | ~new_P3_U2411;
  assign new_P3_U6864 = ~new_P3_ADD_546_U60 | ~new_P3_U2400;
  assign new_P3_U6865 = ~P3_EAX_REG_2_ | ~new_P3_U3252;
  assign new_P3_U6866 = ~new_P3_U2446 | ~BUF2_REG_3_;
  assign new_P3_U6867 = ~new_P3_U2624 | ~new_P3_U2411;
  assign new_P3_U6868 = ~new_P3_ADD_546_U57 | ~new_P3_U2400;
  assign new_P3_U6869 = ~P3_EAX_REG_3_ | ~new_P3_U3252;
  assign new_P3_U6870 = ~new_P3_U2446 | ~BUF2_REG_4_;
  assign new_P3_U6871 = ~new_P3_U2625 | ~new_P3_U2411;
  assign new_P3_U6872 = ~new_P3_ADD_546_U56 | ~new_P3_U2400;
  assign new_P3_U6873 = ~P3_EAX_REG_4_ | ~new_P3_U3252;
  assign new_P3_U6874 = ~new_P3_U2446 | ~BUF2_REG_5_;
  assign new_P3_U6875 = ~new_P3_U2626 | ~new_P3_U2411;
  assign new_P3_U6876 = ~new_P3_ADD_546_U55 | ~new_P3_U2400;
  assign new_P3_U6877 = ~P3_EAX_REG_5_ | ~new_P3_U3252;
  assign new_P3_U6878 = ~new_P3_U2446 | ~BUF2_REG_6_;
  assign new_P3_U6879 = ~new_P3_U2627 | ~new_P3_U2411;
  assign new_P3_U6880 = ~new_P3_ADD_546_U54 | ~new_P3_U2400;
  assign new_P3_U6881 = ~P3_EAX_REG_6_ | ~new_P3_U3252;
  assign new_P3_U6882 = ~new_P3_U2446 | ~BUF2_REG_7_;
  assign new_P3_U6883 = ~new_P3_U2628 | ~new_P3_U2411;
  assign new_P3_U6884 = ~new_P3_ADD_546_U53 | ~new_P3_U2400;
  assign new_P3_U6885 = ~P3_EAX_REG_7_ | ~new_P3_U3252;
  assign new_P3_U6886 = ~new_P3_U2446 | ~BUF2_REG_8_;
  assign new_P3_U6887 = ~new_P3_U2605 | ~new_P3_U2411;
  assign new_P3_U6888 = ~new_P3_ADD_546_U52 | ~new_P3_U2400;
  assign new_P3_U6889 = ~P3_EAX_REG_8_ | ~new_P3_U3252;
  assign new_P3_U6890 = ~new_P3_U2446 | ~BUF2_REG_9_;
  assign new_P3_U6891 = ~new_P3_U2606 | ~new_P3_U2411;
  assign new_P3_U6892 = ~new_P3_ADD_546_U51 | ~new_P3_U2400;
  assign new_P3_U6893 = ~P3_EAX_REG_9_ | ~new_P3_U3252;
  assign new_P3_U6894 = ~new_P3_U2446 | ~BUF2_REG_10_;
  assign new_P3_U6895 = ~new_P3_U2607 | ~new_P3_U2411;
  assign new_P3_U6896 = ~new_P3_ADD_546_U81 | ~new_P3_U2400;
  assign new_P3_U6897 = ~P3_EAX_REG_10_ | ~new_P3_U3252;
  assign new_P3_U6898 = ~new_P3_U2446 | ~BUF2_REG_11_;
  assign new_P3_U6899 = ~new_P3_U2608 | ~new_P3_U2411;
  assign new_P3_U6900 = ~new_P3_ADD_546_U80 | ~new_P3_U2400;
  assign new_P3_U6901 = ~P3_EAX_REG_11_ | ~new_P3_U3252;
  assign new_P3_U6902 = ~new_P3_U2446 | ~BUF2_REG_12_;
  assign new_P3_U6903 = ~new_P3_U2609 | ~new_P3_U2411;
  assign new_P3_U6904 = ~new_P3_ADD_546_U79 | ~new_P3_U2400;
  assign new_P3_U6905 = ~P3_EAX_REG_12_ | ~new_P3_U3252;
  assign new_P3_U6906 = ~new_P3_U2446 | ~BUF2_REG_13_;
  assign new_P3_U6907 = ~new_P3_U2610 | ~new_P3_U2411;
  assign new_P3_U6908 = ~new_P3_ADD_546_U78 | ~new_P3_U2400;
  assign new_P3_U6909 = ~P3_EAX_REG_13_ | ~new_P3_U3252;
  assign new_P3_U6910 = ~new_P3_U2446 | ~BUF2_REG_14_;
  assign new_P3_U6911 = ~new_P3_U2611 | ~new_P3_U2411;
  assign new_P3_U6912 = ~new_P3_ADD_546_U77 | ~new_P3_U2400;
  assign new_P3_U6913 = ~P3_EAX_REG_14_ | ~new_P3_U3252;
  assign new_P3_U6914 = ~new_P3_U2446 | ~BUF2_REG_15_;
  assign new_P3_U6915 = ~new_P3_U2612 | ~new_P3_U2411;
  assign new_P3_U6916 = ~new_P3_ADD_546_U76 | ~new_P3_U2400;
  assign new_P3_U6917 = ~P3_EAX_REG_15_ | ~new_P3_U3252;
  assign new_P3_U6918 = ~new_P3_U2448 | ~BUF2_REG_0_;
  assign new_P3_U6919 = ~new_P3_U2444 | ~BUF2_REG_16_;
  assign new_P3_U6920 = ~new_P3_U3062 | ~new_P3_U2411;
  assign new_P3_U6921 = ~new_P3_ADD_546_U75 | ~new_P3_U2400;
  assign new_P3_U6922 = ~P3_EAX_REG_16_ | ~new_P3_U3252;
  assign new_P3_U6923 = ~new_P3_U2448 | ~BUF2_REG_1_;
  assign new_P3_U6924 = ~new_P3_U2444 | ~BUF2_REG_17_;
  assign new_P3_U6925 = ~new_P3_U3063 | ~new_P3_U2411;
  assign new_P3_U6926 = ~new_P3_ADD_546_U74 | ~new_P3_U2400;
  assign new_P3_U6927 = ~P3_EAX_REG_17_ | ~new_P3_U3252;
  assign new_P3_U6928 = ~new_P3_U2448 | ~BUF2_REG_2_;
  assign new_P3_U6929 = ~new_P3_U2444 | ~BUF2_REG_18_;
  assign new_P3_U6930 = ~new_P3_U3064 | ~new_P3_U2411;
  assign new_P3_U6931 = ~new_P3_ADD_546_U73 | ~new_P3_U2400;
  assign new_P3_U6932 = ~P3_EAX_REG_18_ | ~new_P3_U3252;
  assign new_P3_U6933 = ~new_P3_U2448 | ~BUF2_REG_3_;
  assign new_P3_U6934 = ~new_P3_U2444 | ~BUF2_REG_19_;
  assign new_P3_U6935 = ~new_P3_U3065 | ~new_P3_U2411;
  assign new_P3_U6936 = ~new_P3_ADD_546_U72 | ~new_P3_U2400;
  assign new_P3_U6937 = ~P3_EAX_REG_19_ | ~new_P3_U3252;
  assign new_P3_U6938 = ~new_P3_U2448 | ~BUF2_REG_4_;
  assign new_P3_U6939 = ~new_P3_U2444 | ~BUF2_REG_20_;
  assign new_P3_U6940 = ~new_P3_U3066 | ~new_P3_U2411;
  assign new_P3_U6941 = ~new_P3_ADD_546_U70 | ~new_P3_U2400;
  assign new_P3_U6942 = ~P3_EAX_REG_20_ | ~new_P3_U3252;
  assign new_P3_U6943 = ~new_P3_U2448 | ~BUF2_REG_5_;
  assign new_P3_U6944 = ~new_P3_U2444 | ~BUF2_REG_21_;
  assign new_P3_U6945 = ~new_P3_U3067 | ~new_P3_U2411;
  assign new_P3_U6946 = ~new_P3_ADD_546_U69 | ~new_P3_U2400;
  assign new_P3_U6947 = ~P3_EAX_REG_21_ | ~new_P3_U3252;
  assign new_P3_U6948 = ~new_P3_U2448 | ~BUF2_REG_6_;
  assign new_P3_U6949 = ~new_P3_U2444 | ~BUF2_REG_22_;
  assign new_P3_U6950 = ~new_P3_U3068 | ~new_P3_U2411;
  assign new_P3_U6951 = ~new_P3_ADD_546_U68 | ~new_P3_U2400;
  assign new_P3_U6952 = ~P3_EAX_REG_22_ | ~new_P3_U3252;
  assign new_P3_U6953 = ~new_P3_U2448 | ~BUF2_REG_7_;
  assign new_P3_U6954 = ~new_P3_U2444 | ~BUF2_REG_23_;
  assign new_P3_U6955 = ~new_P3_ADD_391_1180_U25 | ~new_P3_U2411;
  assign new_P3_U6956 = ~new_P3_ADD_546_U67 | ~new_P3_U2400;
  assign new_P3_U6957 = ~P3_EAX_REG_23_ | ~new_P3_U3252;
  assign new_P3_U6958 = ~new_P3_U2448 | ~BUF2_REG_8_;
  assign new_P3_U6959 = ~new_P3_U2444 | ~BUF2_REG_24_;
  assign new_P3_U6960 = ~new_P3_ADD_391_1180_U24 | ~new_P3_U2411;
  assign new_P3_U6961 = ~new_P3_ADD_546_U66 | ~new_P3_U2400;
  assign new_P3_U6962 = ~P3_EAX_REG_24_ | ~new_P3_U3252;
  assign new_P3_U6963 = ~new_P3_U2448 | ~BUF2_REG_9_;
  assign new_P3_U6964 = ~new_P3_U2444 | ~BUF2_REG_25_;
  assign new_P3_U6965 = ~new_P3_ADD_391_1180_U23 | ~new_P3_U2411;
  assign new_P3_U6966 = ~new_P3_ADD_546_U65 | ~new_P3_U2400;
  assign new_P3_U6967 = ~P3_EAX_REG_25_ | ~new_P3_U3252;
  assign new_P3_U6968 = ~new_P3_U2448 | ~BUF2_REG_10_;
  assign new_P3_U6969 = ~new_P3_U2444 | ~BUF2_REG_26_;
  assign new_P3_U6970 = ~new_P3_ADD_391_1180_U22 | ~new_P3_U2411;
  assign new_P3_U6971 = ~new_P3_ADD_546_U64 | ~new_P3_U2400;
  assign new_P3_U6972 = ~P3_EAX_REG_26_ | ~new_P3_U3252;
  assign new_P3_U6973 = ~new_P3_U2448 | ~BUF2_REG_11_;
  assign new_P3_U6974 = ~new_P3_U2444 | ~BUF2_REG_27_;
  assign new_P3_U6975 = ~new_P3_ADD_391_1180_U21 | ~new_P3_U2411;
  assign new_P3_U6976 = ~new_P3_ADD_546_U63 | ~new_P3_U2400;
  assign new_P3_U6977 = ~P3_EAX_REG_27_ | ~new_P3_U3252;
  assign new_P3_U6978 = ~new_P3_U2448 | ~BUF2_REG_12_;
  assign new_P3_U6979 = ~new_P3_U2444 | ~BUF2_REG_28_;
  assign new_P3_U6980 = ~new_P3_ADD_391_1180_U20 | ~new_P3_U2411;
  assign new_P3_U6981 = ~new_P3_ADD_546_U62 | ~new_P3_U2400;
  assign new_P3_U6982 = ~P3_EAX_REG_28_ | ~new_P3_U3252;
  assign new_P3_U6983 = ~new_P3_U2448 | ~BUF2_REG_13_;
  assign new_P3_U6984 = ~new_P3_U2444 | ~BUF2_REG_29_;
  assign new_P3_U6985 = ~new_P3_ADD_391_1180_U19 | ~new_P3_U2411;
  assign new_P3_U6986 = ~new_P3_ADD_546_U61 | ~new_P3_U2400;
  assign new_P3_U6987 = ~P3_EAX_REG_29_ | ~new_P3_U3252;
  assign new_P3_U6988 = ~new_P3_U2448 | ~BUF2_REG_14_;
  assign new_P3_U6989 = ~new_P3_U2444 | ~BUF2_REG_30_;
  assign new_P3_U6990 = ~new_P3_ADD_391_1180_U18 | ~new_P3_U2411;
  assign new_P3_U6991 = ~new_P3_ADD_546_U59 | ~new_P3_U2400;
  assign new_P3_U6992 = ~P3_EAX_REG_30_ | ~new_P3_U3252;
  assign new_P3_U6993 = ~new_P3_U2444 | ~BUF2_REG_31_;
  assign new_P3_U6994 = ~new_P3_ADD_546_U58 | ~new_P3_U2400;
  assign new_P3_U6995 = ~P3_EAX_REG_31_ | ~new_P3_U3252;
  assign new_P3_U6996 = ~new_P3_GTE_401_U6 | ~new_P3_U4305;
  assign new_P3_U6997 = ~new_P3_U3242 | ~new_P3_U6996;
  assign new_P3_U6998 = ~P3_INSTQUEUE_REG_0__0_ | ~new_P3_U2408;
  assign new_P3_U6999 = ~new_P3_ADD_552_U5 | ~new_P3_U2399;
  assign new_P3_U7000 = ~P3_EBX_REG_0_ | ~new_P3_U3253;
  assign new_P3_U7001 = ~P3_INSTQUEUE_REG_0__1_ | ~new_P3_U2408;
  assign new_P3_U7002 = ~new_P3_ADD_552_U71 | ~new_P3_U2399;
  assign new_P3_U7003 = ~P3_EBX_REG_1_ | ~new_P3_U3253;
  assign new_P3_U7004 = ~P3_INSTQUEUE_REG_0__2_ | ~new_P3_U2408;
  assign new_P3_U7005 = ~new_P3_ADD_552_U60 | ~new_P3_U2399;
  assign new_P3_U7006 = ~P3_EBX_REG_2_ | ~new_P3_U3253;
  assign new_P3_U7007 = ~P3_INSTQUEUE_REG_0__3_ | ~new_P3_U2408;
  assign new_P3_U7008 = ~new_P3_ADD_552_U57 | ~new_P3_U2399;
  assign new_P3_U7009 = ~P3_EBX_REG_3_ | ~new_P3_U3253;
  assign new_P3_U7010 = ~P3_INSTQUEUE_REG_0__4_ | ~new_P3_U2408;
  assign new_P3_U7011 = ~new_P3_ADD_552_U56 | ~new_P3_U2399;
  assign new_P3_U7012 = ~P3_EBX_REG_4_ | ~new_P3_U3253;
  assign new_P3_U7013 = ~P3_INSTQUEUE_REG_0__5_ | ~new_P3_U2408;
  assign new_P3_U7014 = ~new_P3_ADD_552_U55 | ~new_P3_U2399;
  assign new_P3_U7015 = ~P3_EBX_REG_5_ | ~new_P3_U3253;
  assign new_P3_U7016 = ~P3_INSTQUEUE_REG_0__6_ | ~new_P3_U2408;
  assign new_P3_U7017 = ~new_P3_ADD_552_U54 | ~new_P3_U2399;
  assign new_P3_U7018 = ~P3_EBX_REG_6_ | ~new_P3_U3253;
  assign new_P3_U7019 = ~P3_INSTQUEUE_REG_0__7_ | ~new_P3_U2408;
  assign new_P3_U7020 = ~new_P3_ADD_552_U53 | ~new_P3_U2399;
  assign new_P3_U7021 = ~P3_EBX_REG_7_ | ~new_P3_U3253;
  assign new_P3_U7022 = ~new_P3_U2605 | ~new_P3_U2408;
  assign new_P3_U7023 = ~new_P3_ADD_552_U52 | ~new_P3_U2399;
  assign new_P3_U7024 = ~P3_EBX_REG_8_ | ~new_P3_U3253;
  assign new_P3_U7025 = ~new_P3_U2606 | ~new_P3_U2408;
  assign new_P3_U7026 = ~new_P3_ADD_552_U51 | ~new_P3_U2399;
  assign new_P3_U7027 = ~P3_EBX_REG_9_ | ~new_P3_U3253;
  assign new_P3_U7028 = ~new_P3_U2607 | ~new_P3_U2408;
  assign new_P3_U7029 = ~new_P3_ADD_552_U81 | ~new_P3_U2399;
  assign new_P3_U7030 = ~P3_EBX_REG_10_ | ~new_P3_U3253;
  assign new_P3_U7031 = ~new_P3_U2608 | ~new_P3_U2408;
  assign new_P3_U7032 = ~new_P3_ADD_552_U80 | ~new_P3_U2399;
  assign new_P3_U7033 = ~P3_EBX_REG_11_ | ~new_P3_U3253;
  assign new_P3_U7034 = ~new_P3_U2609 | ~new_P3_U2408;
  assign new_P3_U7035 = ~new_P3_ADD_552_U79 | ~new_P3_U2399;
  assign new_P3_U7036 = ~P3_EBX_REG_12_ | ~new_P3_U3253;
  assign new_P3_U7037 = ~new_P3_U2610 | ~new_P3_U2408;
  assign new_P3_U7038 = ~new_P3_ADD_552_U78 | ~new_P3_U2399;
  assign new_P3_U7039 = ~P3_EBX_REG_13_ | ~new_P3_U3253;
  assign new_P3_U7040 = ~new_P3_U2611 | ~new_P3_U2408;
  assign new_P3_U7041 = ~new_P3_ADD_552_U77 | ~new_P3_U2399;
  assign new_P3_U7042 = ~P3_EBX_REG_14_ | ~new_P3_U3253;
  assign new_P3_U7043 = ~new_P3_U2612 | ~new_P3_U2408;
  assign new_P3_U7044 = ~new_P3_ADD_552_U76 | ~new_P3_U2399;
  assign new_P3_U7045 = ~P3_EBX_REG_15_ | ~new_P3_U3253;
  assign new_P3_U7046 = ~new_P3_U3062 | ~new_P3_U2408;
  assign new_P3_U7047 = ~new_P3_ADD_552_U75 | ~new_P3_U2399;
  assign new_P3_U7048 = ~P3_EBX_REG_16_ | ~new_P3_U3253;
  assign new_P3_U7049 = ~new_P3_U3063 | ~new_P3_U2408;
  assign new_P3_U7050 = ~new_P3_ADD_552_U74 | ~new_P3_U2399;
  assign new_P3_U7051 = ~P3_EBX_REG_17_ | ~new_P3_U3253;
  assign new_P3_U7052 = ~new_P3_U3064 | ~new_P3_U2408;
  assign new_P3_U7053 = ~new_P3_ADD_552_U73 | ~new_P3_U2399;
  assign new_P3_U7054 = ~P3_EBX_REG_18_ | ~new_P3_U3253;
  assign new_P3_U7055 = ~new_P3_U3065 | ~new_P3_U2408;
  assign new_P3_U7056 = ~new_P3_ADD_552_U72 | ~new_P3_U2399;
  assign new_P3_U7057 = ~P3_EBX_REG_19_ | ~new_P3_U3253;
  assign new_P3_U7058 = ~new_P3_U3066 | ~new_P3_U2408;
  assign new_P3_U7059 = ~new_P3_ADD_552_U70 | ~new_P3_U2399;
  assign new_P3_U7060 = ~P3_EBX_REG_20_ | ~new_P3_U3253;
  assign new_P3_U7061 = ~new_P3_U3067 | ~new_P3_U2408;
  assign new_P3_U7062 = ~new_P3_ADD_552_U69 | ~new_P3_U2399;
  assign new_P3_U7063 = ~P3_EBX_REG_21_ | ~new_P3_U3253;
  assign new_P3_U7064 = ~new_P3_U3068 | ~new_P3_U2408;
  assign new_P3_U7065 = ~new_P3_ADD_552_U68 | ~new_P3_U2399;
  assign new_P3_U7066 = ~P3_EBX_REG_22_ | ~new_P3_U3253;
  assign new_P3_U7067 = ~new_P3_ADD_402_1132_U25 | ~new_P3_U2408;
  assign new_P3_U7068 = ~new_P3_ADD_552_U67 | ~new_P3_U2399;
  assign new_P3_U7069 = ~P3_EBX_REG_23_ | ~new_P3_U3253;
  assign new_P3_U7070 = ~new_P3_ADD_402_1132_U24 | ~new_P3_U2408;
  assign new_P3_U7071 = ~new_P3_ADD_552_U66 | ~new_P3_U2399;
  assign new_P3_U7072 = ~P3_EBX_REG_24_ | ~new_P3_U3253;
  assign new_P3_U7073 = ~new_P3_ADD_402_1132_U23 | ~new_P3_U2408;
  assign new_P3_U7074 = ~new_P3_ADD_552_U65 | ~new_P3_U2399;
  assign new_P3_U7075 = ~P3_EBX_REG_25_ | ~new_P3_U3253;
  assign new_P3_U7076 = ~new_P3_ADD_402_1132_U22 | ~new_P3_U2408;
  assign new_P3_U7077 = ~new_P3_ADD_552_U64 | ~new_P3_U2399;
  assign new_P3_U7078 = ~P3_EBX_REG_26_ | ~new_P3_U3253;
  assign new_P3_U7079 = ~new_P3_ADD_402_1132_U21 | ~new_P3_U2408;
  assign new_P3_U7080 = ~new_P3_ADD_552_U63 | ~new_P3_U2399;
  assign new_P3_U7081 = ~P3_EBX_REG_27_ | ~new_P3_U3253;
  assign new_P3_U7082 = ~new_P3_ADD_402_1132_U20 | ~new_P3_U2408;
  assign new_P3_U7083 = ~new_P3_ADD_552_U62 | ~new_P3_U2399;
  assign new_P3_U7084 = ~P3_EBX_REG_28_ | ~new_P3_U3253;
  assign new_P3_U7085 = ~new_P3_ADD_402_1132_U19 | ~new_P3_U2408;
  assign new_P3_U7086 = ~new_P3_ADD_552_U61 | ~new_P3_U2399;
  assign new_P3_U7087 = ~P3_EBX_REG_29_ | ~new_P3_U3253;
  assign new_P3_U7088 = ~new_P3_ADD_402_1132_U18 | ~new_P3_U2408;
  assign new_P3_U7089 = ~new_P3_ADD_552_U59 | ~new_P3_U2399;
  assign new_P3_U7090 = ~P3_EBX_REG_30_ | ~new_P3_U3253;
  assign new_P3_U7091 = ~new_P3_ADD_552_U58 | ~new_P3_U2399;
  assign new_P3_U7092 = ~P3_EBX_REG_31_ | ~new_P3_U3253;
  assign new_P3_U7093 = ~new_P3_U5488 | ~new_P3_U5491;
  assign new_P3_U7094 = ~new_P3_U3260;
  assign new_P3_U7095 = ~new_P3_U3257;
  assign new_P3_U7096 = P3_STATEBS16_REG | new_U209;
  assign new_P3_U7097 = ~P3_EBX_REG_0_ | ~new_P3_U2602;
  assign new_P3_U7098 = ~P3_REIP_REG_0_ | ~new_P3_U2601;
  assign new_P3_U7099 = ~P3_EBX_REG_0_ | ~new_P3_U7910;
  assign new_P3_U7100 = ~new_P3_ADD_505_U5 | ~new_P3_U2455;
  assign new_P3_U7101 = ~new_P3_ADD_486_U5 | ~new_P3_U2454;
  assign new_P3_U7102 = ~P3_REIP_REG_0_ | ~new_P3_U2405;
  assign new_P3_U7103 = ~new_P3_U2403 | ~P3_PHYADDRPOINTER_REG_0_;
  assign new_P3_U7104 = ~P3_PHYADDRPOINTER_REG_0_ | ~new_P3_U4319;
  assign new_P3_U7105 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_0_;
  assign new_P3_U7106 = ~new_P3_U7094 | ~P3_REIP_REG_0_;
  assign new_P3_U7107 = ~new_P3_SUB_414_U50 | ~new_P3_U2602;
  assign new_P3_U7108 = ~new_P3_ADD_467_U4 | ~new_P3_U2601;
  assign new_P3_U7109 = ~P3_EBX_REG_1_ | ~new_P3_U7910;
  assign new_P3_U7110 = ~new_P3_ADD_505_U17 | ~new_P3_U2455;
  assign new_P3_U7111 = ~new_P3_ADD_486_U17 | ~new_P3_U2454;
  assign new_P3_U7112 = ~new_P3_ADD_430_U4 | ~new_P3_U2405;
  assign new_P3_U7113 = ~new_P3_U2403 | ~new_P3_ADD_318_U4;
  assign new_P3_U7114 = ~new_P3_SUB_320_U50 | ~new_P3_U4319;
  assign new_P3_U7115 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_1_;
  assign new_P3_U7116 = ~new_P3_U7094 | ~P3_REIP_REG_1_;
  assign new_P3_U7117 = ~new_P3_SUB_414_U17 | ~new_P3_U2602;
  assign new_P3_U7118 = ~new_P3_ADD_467_U71 | ~new_P3_U2601;
  assign new_P3_U7119 = ~P3_EBX_REG_2_ | ~new_P3_U7910;
  assign new_P3_U7120 = ~new_P3_ADD_505_U16 | ~new_P3_U2455;
  assign new_P3_U7121 = ~new_P3_ADD_486_U16 | ~new_P3_U2454;
  assign new_P3_U7122 = ~new_P3_ADD_430_U71 | ~new_P3_U2405;
  assign new_P3_U7123 = ~new_P3_U2403 | ~new_P3_ADD_318_U71;
  assign new_P3_U7124 = ~new_P3_SUB_320_U17 | ~new_P3_U4319;
  assign new_P3_U7125 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_2_;
  assign new_P3_U7126 = ~new_P3_U7094 | ~P3_REIP_REG_2_;
  assign new_P3_U7127 = ~new_P3_SUB_414_U59 | ~new_P3_U2602;
  assign new_P3_U7128 = ~new_P3_ADD_467_U68 | ~new_P3_U2601;
  assign new_P3_U7129 = ~P3_EBX_REG_3_ | ~new_P3_U7910;
  assign new_P3_U7130 = ~new_P3_ADD_505_U15 | ~new_P3_U2455;
  assign new_P3_U7131 = ~new_P3_ADD_486_U15 | ~new_P3_U2454;
  assign new_P3_U7132 = ~new_P3_ADD_430_U68 | ~new_P3_U2405;
  assign new_P3_U7133 = ~new_P3_U2403 | ~new_P3_ADD_318_U68;
  assign new_P3_U7134 = ~new_P3_SUB_320_U59 | ~new_P3_U4319;
  assign new_P3_U7135 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_3_;
  assign new_P3_U7136 = ~new_P3_U7094 | ~P3_REIP_REG_3_;
  assign new_P3_U7137 = ~new_P3_SUB_414_U18 | ~new_P3_U2602;
  assign new_P3_U7138 = ~new_P3_ADD_467_U67 | ~new_P3_U2601;
  assign new_P3_U7139 = ~P3_EBX_REG_4_ | ~new_P3_U7910;
  assign new_P3_U7140 = ~new_P3_ADD_505_U14 | ~new_P3_U2455;
  assign new_P3_U7141 = ~new_P3_ADD_486_U14 | ~new_P3_U2454;
  assign new_P3_U7142 = ~new_P3_ADD_430_U67 | ~new_P3_U2405;
  assign new_P3_U7143 = ~new_P3_U2403 | ~new_P3_ADD_318_U67;
  assign new_P3_U7144 = ~new_P3_SUB_320_U18 | ~new_P3_U4319;
  assign new_P3_U7145 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_4_;
  assign new_P3_U7146 = ~new_P3_U7094 | ~P3_REIP_REG_4_;
  assign new_P3_U7147 = ~new_P3_SUB_414_U57 | ~new_P3_U2602;
  assign new_P3_U7148 = ~new_P3_ADD_467_U66 | ~new_P3_U2601;
  assign new_P3_U7149 = ~P3_EBX_REG_5_ | ~new_P3_U7910;
  assign new_P3_U7150 = ~new_P3_ADD_505_U6 | ~new_P3_U2455;
  assign new_P3_U7151 = ~new_P3_ADD_486_U6 | ~new_P3_U2454;
  assign new_P3_U7152 = ~new_P3_ADD_430_U66 | ~new_P3_U2405;
  assign new_P3_U7153 = ~new_P3_U2403 | ~new_P3_ADD_318_U66;
  assign new_P3_U7154 = ~new_P3_SUB_320_U57 | ~new_P3_U4319;
  assign new_P3_U7155 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_5_;
  assign new_P3_U7156 = ~new_P3_U7094 | ~P3_REIP_REG_5_;
  assign new_P3_U7157 = ~new_P3_SUB_414_U19 | ~new_P3_U2602;
  assign new_P3_U7158 = ~new_P3_ADD_467_U65 | ~new_P3_U2601;
  assign new_P3_U7159 = ~P3_EBX_REG_6_ | ~new_P3_U7910;
  assign new_P3_U7160 = ~new_P3_ADD_430_U65 | ~new_P3_U2405;
  assign new_P3_U7161 = ~new_P3_U2403 | ~new_P3_ADD_318_U65;
  assign new_P3_U7162 = ~new_P3_SUB_320_U19 | ~new_P3_U4319;
  assign new_P3_U7163 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_6_;
  assign new_P3_U7164 = ~new_P3_U7094 | ~P3_REIP_REG_6_;
  assign new_P3_U7165 = ~new_P3_SUB_414_U55 | ~new_P3_U2602;
  assign new_P3_U7166 = ~new_P3_ADD_467_U64 | ~new_P3_U2601;
  assign new_P3_U7167 = ~P3_EBX_REG_7_ | ~new_P3_U7910;
  assign new_P3_U7168 = ~new_P3_ADD_430_U64 | ~new_P3_U2405;
  assign new_P3_U7169 = ~new_P3_U2403 | ~new_P3_ADD_318_U64;
  assign new_P3_U7170 = ~new_P3_SUB_320_U55 | ~new_P3_U4319;
  assign new_P3_U7171 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_7_;
  assign new_P3_U7172 = ~new_P3_U7094 | ~P3_REIP_REG_7_;
  assign new_P3_U7173 = ~new_P3_SUB_414_U20 | ~new_P3_U2602;
  assign new_P3_U7174 = ~new_P3_ADD_467_U63 | ~new_P3_U2601;
  assign new_P3_U7175 = ~P3_EBX_REG_8_ | ~new_P3_U7910;
  assign new_P3_U7176 = ~new_P3_ADD_430_U63 | ~new_P3_U2405;
  assign new_P3_U7177 = ~new_P3_U2403 | ~new_P3_ADD_318_U63;
  assign new_P3_U7178 = ~new_P3_SUB_320_U20 | ~new_P3_U4319;
  assign new_P3_U7179 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_8_;
  assign new_P3_U7180 = ~new_P3_U7094 | ~P3_REIP_REG_8_;
  assign new_P3_U7181 = ~new_P3_SUB_414_U53 | ~new_P3_U2602;
  assign new_P3_U7182 = ~new_P3_ADD_467_U62 | ~new_P3_U2601;
  assign new_P3_U7183 = ~P3_EBX_REG_9_ | ~new_P3_U7910;
  assign new_P3_U7184 = ~new_P3_ADD_430_U62 | ~new_P3_U2405;
  assign new_P3_U7185 = ~new_P3_U2403 | ~new_P3_ADD_318_U62;
  assign new_P3_U7186 = ~new_P3_SUB_320_U53 | ~new_P3_U4319;
  assign new_P3_U7187 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_U7188 = ~new_P3_U7094 | ~P3_REIP_REG_9_;
  assign new_P3_U7189 = ~new_P3_SUB_414_U6 | ~new_P3_U2602;
  assign new_P3_U7190 = ~new_P3_ADD_467_U91 | ~new_P3_U2601;
  assign new_P3_U7191 = ~P3_EBX_REG_10_ | ~new_P3_U7910;
  assign new_P3_U7192 = ~new_P3_ADD_430_U91 | ~new_P3_U2405;
  assign new_P3_U7193 = ~new_P3_U2403 | ~new_P3_ADD_318_U91;
  assign new_P3_U7194 = ~new_P3_SUB_320_U6 | ~new_P3_U4319;
  assign new_P3_U7195 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_10_;
  assign new_P3_U7196 = ~new_P3_U7094 | ~P3_REIP_REG_10_;
  assign new_P3_U7197 = ~new_P3_SUB_414_U82 | ~new_P3_U2602;
  assign new_P3_U7198 = ~new_P3_ADD_467_U90 | ~new_P3_U2601;
  assign new_P3_U7199 = ~P3_EBX_REG_11_ | ~new_P3_U7910;
  assign new_P3_U7200 = ~new_P3_ADD_430_U90 | ~new_P3_U2405;
  assign new_P3_U7201 = ~new_P3_U2403 | ~new_P3_ADD_318_U90;
  assign new_P3_U7202 = ~new_P3_SUB_320_U82 | ~new_P3_U4319;
  assign new_P3_U7203 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_11_;
  assign new_P3_U7204 = ~new_P3_U7094 | ~P3_REIP_REG_11_;
  assign new_P3_U7205 = ~new_P3_SUB_414_U7 | ~new_P3_U2602;
  assign new_P3_U7206 = ~new_P3_ADD_467_U89 | ~new_P3_U2601;
  assign new_P3_U7207 = ~P3_EBX_REG_12_ | ~new_P3_U7910;
  assign new_P3_U7208 = ~new_P3_ADD_430_U89 | ~new_P3_U2405;
  assign new_P3_U7209 = ~new_P3_U2403 | ~new_P3_ADD_318_U89;
  assign new_P3_U7210 = ~new_P3_SUB_320_U7 | ~new_P3_U4319;
  assign new_P3_U7211 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_12_;
  assign new_P3_U7212 = ~new_P3_U7094 | ~P3_REIP_REG_12_;
  assign new_P3_U7213 = ~new_P3_SUB_414_U80 | ~new_P3_U2602;
  assign new_P3_U7214 = ~new_P3_ADD_467_U88 | ~new_P3_U2601;
  assign new_P3_U7215 = ~P3_EBX_REG_13_ | ~new_P3_U7910;
  assign new_P3_U7216 = ~new_P3_ADD_430_U88 | ~new_P3_U2405;
  assign new_P3_U7217 = ~new_P3_U2403 | ~new_P3_ADD_318_U88;
  assign new_P3_U7218 = ~new_P3_SUB_320_U80 | ~new_P3_U4319;
  assign new_P3_U7219 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_13_;
  assign new_P3_U7220 = ~new_P3_U7094 | ~P3_REIP_REG_13_;
  assign new_P3_U7221 = ~new_P3_SUB_414_U8 | ~new_P3_U2602;
  assign new_P3_U7222 = ~new_P3_ADD_467_U87 | ~new_P3_U2601;
  assign new_P3_U7223 = ~P3_EBX_REG_14_ | ~new_P3_U7910;
  assign new_P3_U7224 = ~new_P3_ADD_430_U87 | ~new_P3_U2405;
  assign new_P3_U7225 = ~new_P3_U2403 | ~new_P3_ADD_318_U87;
  assign new_P3_U7226 = ~new_P3_SUB_320_U8 | ~new_P3_U4319;
  assign new_P3_U7227 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_14_;
  assign new_P3_U7228 = ~new_P3_U7094 | ~P3_REIP_REG_14_;
  assign new_P3_U7229 = ~new_P3_SUB_414_U78 | ~new_P3_U2602;
  assign new_P3_U7230 = ~new_P3_ADD_467_U86 | ~new_P3_U2601;
  assign new_P3_U7231 = ~P3_EBX_REG_15_ | ~new_P3_U7910;
  assign new_P3_U7232 = ~new_P3_ADD_430_U86 | ~new_P3_U2405;
  assign new_P3_U7233 = ~new_P3_U2403 | ~new_P3_ADD_318_U86;
  assign new_P3_U7234 = ~new_P3_SUB_320_U78 | ~new_P3_U4319;
  assign new_P3_U7235 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_15_;
  assign new_P3_U7236 = ~new_P3_U7094 | ~P3_REIP_REG_15_;
  assign new_P3_U7237 = ~new_P3_SUB_414_U9 | ~new_P3_U2602;
  assign new_P3_U7238 = ~new_P3_ADD_467_U85 | ~new_P3_U2601;
  assign new_P3_U7239 = ~P3_EBX_REG_16_ | ~new_P3_U7910;
  assign new_P3_U7240 = ~new_P3_ADD_430_U85 | ~new_P3_U2405;
  assign new_P3_U7241 = ~new_P3_U2403 | ~new_P3_ADD_318_U85;
  assign new_P3_U7242 = ~new_P3_SUB_320_U9 | ~new_P3_U4319;
  assign new_P3_U7243 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_16_;
  assign new_P3_U7244 = ~new_P3_U7094 | ~P3_REIP_REG_16_;
  assign new_P3_U7245 = ~new_P3_SUB_414_U76 | ~new_P3_U2602;
  assign new_P3_U7246 = ~new_P3_ADD_467_U84 | ~new_P3_U2601;
  assign new_P3_U7247 = ~P3_EBX_REG_17_ | ~new_P3_U7910;
  assign new_P3_U7248 = ~new_P3_ADD_430_U84 | ~new_P3_U2405;
  assign new_P3_U7249 = ~new_P3_U2403 | ~new_P3_ADD_318_U84;
  assign new_P3_U7250 = ~new_P3_SUB_320_U76 | ~new_P3_U4319;
  assign new_P3_U7251 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_17_;
  assign new_P3_U7252 = ~new_P3_U7094 | ~P3_REIP_REG_17_;
  assign new_P3_U7253 = ~new_P3_SUB_414_U10 | ~new_P3_U2602;
  assign new_P3_U7254 = ~new_P3_ADD_467_U83 | ~new_P3_U2601;
  assign new_P3_U7255 = ~P3_EBX_REG_18_ | ~new_P3_U7910;
  assign new_P3_U7256 = ~new_P3_ADD_430_U83 | ~new_P3_U2405;
  assign new_P3_U7257 = ~new_P3_U2403 | ~new_P3_ADD_318_U83;
  assign new_P3_U7258 = ~new_P3_SUB_320_U10 | ~new_P3_U4319;
  assign new_P3_U7259 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_18_;
  assign new_P3_U7260 = ~new_P3_U7094 | ~P3_REIP_REG_18_;
  assign new_P3_U7261 = ~new_P3_SUB_414_U74 | ~new_P3_U2602;
  assign new_P3_U7262 = ~new_P3_ADD_467_U82 | ~new_P3_U2601;
  assign new_P3_U7263 = ~P3_EBX_REG_19_ | ~new_P3_U7910;
  assign new_P3_U7264 = ~new_P3_ADD_430_U82 | ~new_P3_U2405;
  assign new_P3_U7265 = ~new_P3_U2403 | ~new_P3_ADD_318_U82;
  assign new_P3_U7266 = ~new_P3_SUB_320_U74 | ~new_P3_U4319;
  assign new_P3_U7267 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_19_;
  assign new_P3_U7268 = ~new_P3_U7094 | ~P3_REIP_REG_19_;
  assign new_P3_U7269 = ~new_P3_SUB_414_U11 | ~new_P3_U2602;
  assign new_P3_U7270 = ~new_P3_ADD_467_U81 | ~new_P3_U2601;
  assign new_P3_U7271 = ~P3_EBX_REG_20_ | ~new_P3_U7910;
  assign new_P3_U7272 = ~new_P3_ADD_430_U81 | ~new_P3_U2405;
  assign new_P3_U7273 = ~new_P3_U2403 | ~new_P3_ADD_318_U81;
  assign new_P3_U7274 = ~new_P3_SUB_320_U11 | ~new_P3_U4319;
  assign new_P3_U7275 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_20_;
  assign new_P3_U7276 = ~new_P3_U7094 | ~P3_REIP_REG_20_;
  assign new_P3_U7277 = ~new_P3_SUB_414_U70 | ~new_P3_U2602;
  assign new_P3_U7278 = ~new_P3_ADD_467_U80 | ~new_P3_U2601;
  assign new_P3_U7279 = ~P3_EBX_REG_21_ | ~new_P3_U7910;
  assign new_P3_U7280 = ~new_P3_ADD_430_U80 | ~new_P3_U2405;
  assign new_P3_U7281 = ~new_P3_U2403 | ~new_P3_ADD_318_U80;
  assign new_P3_U7282 = ~new_P3_SUB_320_U70 | ~new_P3_U4319;
  assign new_P3_U7283 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_21_;
  assign new_P3_U7284 = ~new_P3_U7094 | ~P3_REIP_REG_21_;
  assign new_P3_U7285 = ~new_P3_SUB_414_U12 | ~new_P3_U2602;
  assign new_P3_U7286 = ~new_P3_ADD_467_U79 | ~new_P3_U2601;
  assign new_P3_U7287 = ~P3_EBX_REG_22_ | ~new_P3_U7910;
  assign new_P3_U7288 = ~new_P3_ADD_430_U79 | ~new_P3_U2405;
  assign new_P3_U7289 = ~new_P3_U2403 | ~new_P3_ADD_318_U79;
  assign new_P3_U7290 = ~new_P3_SUB_320_U12 | ~new_P3_U4319;
  assign new_P3_U7291 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_22_;
  assign new_P3_U7292 = ~new_P3_U7094 | ~P3_REIP_REG_22_;
  assign new_P3_U7293 = ~new_P3_SUB_414_U68 | ~new_P3_U2602;
  assign new_P3_U7294 = ~new_P3_ADD_467_U78 | ~new_P3_U2601;
  assign new_P3_U7295 = ~P3_EBX_REG_23_ | ~new_P3_U7910;
  assign new_P3_U7296 = ~new_P3_ADD_430_U78 | ~new_P3_U2405;
  assign new_P3_U7297 = ~new_P3_U2403 | ~new_P3_ADD_318_U78;
  assign new_P3_U7298 = ~new_P3_SUB_320_U68 | ~new_P3_U4319;
  assign new_P3_U7299 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_23_;
  assign new_P3_U7300 = ~new_P3_U7094 | ~P3_REIP_REG_23_;
  assign new_P3_U7301 = ~new_P3_SUB_414_U13 | ~new_P3_U2602;
  assign new_P3_U7302 = ~new_P3_ADD_467_U77 | ~new_P3_U2601;
  assign new_P3_U7303 = ~P3_EBX_REG_24_ | ~new_P3_U7910;
  assign new_P3_U7304 = ~new_P3_ADD_430_U77 | ~new_P3_U2405;
  assign new_P3_U7305 = ~new_P3_U2403 | ~new_P3_ADD_318_U77;
  assign new_P3_U7306 = ~new_P3_SUB_320_U13 | ~new_P3_U4319;
  assign new_P3_U7307 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_24_;
  assign new_P3_U7308 = ~new_P3_U7094 | ~P3_REIP_REG_24_;
  assign new_P3_U7309 = ~new_P3_SUB_414_U66 | ~new_P3_U2602;
  assign new_P3_U7310 = ~new_P3_ADD_467_U76 | ~new_P3_U2601;
  assign new_P3_U7311 = ~P3_EBX_REG_25_ | ~new_P3_U7910;
  assign new_P3_U7312 = ~new_P3_ADD_430_U76 | ~new_P3_U2405;
  assign new_P3_U7313 = ~new_P3_U2403 | ~new_P3_ADD_318_U76;
  assign new_P3_U7314 = ~new_P3_SUB_320_U66 | ~new_P3_U4319;
  assign new_P3_U7315 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_25_;
  assign new_P3_U7316 = ~new_P3_U7094 | ~P3_REIP_REG_25_;
  assign new_P3_U7317 = ~new_P3_SUB_414_U14 | ~new_P3_U2602;
  assign new_P3_U7318 = ~new_P3_ADD_467_U75 | ~new_P3_U2601;
  assign new_P3_U7319 = ~P3_EBX_REG_26_ | ~new_P3_U7910;
  assign new_P3_U7320 = ~new_P3_ADD_430_U75 | ~new_P3_U2405;
  assign new_P3_U7321 = ~new_P3_U2403 | ~new_P3_ADD_318_U75;
  assign new_P3_U7322 = ~new_P3_SUB_320_U14 | ~new_P3_U4319;
  assign new_P3_U7323 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_26_;
  assign new_P3_U7324 = ~new_P3_U7094 | ~P3_REIP_REG_26_;
  assign new_P3_U7325 = ~new_P3_SUB_414_U64 | ~new_P3_U2602;
  assign new_P3_U7326 = ~new_P3_ADD_467_U74 | ~new_P3_U2601;
  assign new_P3_U7327 = ~P3_EBX_REG_27_ | ~new_P3_U7910;
  assign new_P3_U7328 = ~new_P3_ADD_430_U74 | ~new_P3_U2405;
  assign new_P3_U7329 = ~new_P3_U2403 | ~new_P3_ADD_318_U74;
  assign new_P3_U7330 = ~new_P3_SUB_320_U64 | ~new_P3_U4319;
  assign new_P3_U7331 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_27_;
  assign new_P3_U7332 = ~new_P3_U7094 | ~P3_REIP_REG_27_;
  assign new_P3_U7333 = ~new_P3_SUB_414_U15 | ~new_P3_U2602;
  assign new_P3_U7334 = ~new_P3_ADD_467_U73 | ~new_P3_U2601;
  assign new_P3_U7335 = ~P3_EBX_REG_28_ | ~new_P3_U7910;
  assign new_P3_U7336 = ~new_P3_ADD_430_U73 | ~new_P3_U2405;
  assign new_P3_U7337 = ~new_P3_U2403 | ~new_P3_ADD_318_U73;
  assign new_P3_U7338 = ~new_P3_SUB_320_U15 | ~new_P3_U4319;
  assign new_P3_U7339 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_28_;
  assign new_P3_U7340 = ~new_P3_U7094 | ~P3_REIP_REG_28_;
  assign new_P3_U7341 = ~new_P3_SUB_414_U16 | ~new_P3_U2602;
  assign new_P3_U7342 = ~new_P3_ADD_467_U72 | ~new_P3_U2601;
  assign new_P3_U7343 = ~P3_EBX_REG_29_ | ~new_P3_U7910;
  assign new_P3_U7344 = ~new_P3_ADD_430_U72 | ~new_P3_U2405;
  assign new_P3_U7345 = ~new_P3_U2403 | ~new_P3_ADD_318_U72;
  assign new_P3_U7346 = ~new_P3_SUB_320_U16 | ~new_P3_U4319;
  assign new_P3_U7347 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_29_;
  assign new_P3_U7348 = ~new_P3_U7094 | ~P3_REIP_REG_29_;
  assign new_P3_U7349 = ~new_P3_SUB_414_U62 | ~new_P3_U2602;
  assign new_P3_U7350 = ~new_P3_ADD_467_U70 | ~new_P3_U2601;
  assign new_P3_U7351 = ~P3_EBX_REG_30_ | ~new_P3_U7910;
  assign new_P3_U7352 = ~new_P3_ADD_430_U70 | ~new_P3_U2405;
  assign new_P3_U7353 = ~new_P3_U2403 | ~new_P3_ADD_318_U70;
  assign new_P3_U7354 = ~new_P3_SUB_320_U62 | ~new_P3_U4319;
  assign new_P3_U7355 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_30_;
  assign new_P3_U7356 = ~new_P3_U7094 | ~P3_REIP_REG_30_;
  assign new_P3_U7357 = ~new_P3_U4135 | ~new_P3_U2603;
  assign new_P3_U7358 = ~new_P3_SUB_414_U51 | ~new_P3_U2602;
  assign new_P3_U7359 = ~new_P3_ADD_467_U69 | ~new_P3_U2601;
  assign new_P3_U7360 = ~P3_EBX_REG_31_ | ~new_P3_U7910;
  assign new_P3_U7361 = ~new_P3_ADD_430_U69 | ~new_P3_U2405;
  assign new_P3_U7362 = ~new_P3_U2403 | ~new_P3_ADD_318_U69;
  assign new_P3_U7363 = ~new_P3_U7362;
  assign new_P3_U7364 = ~new_P3_U2401 | ~P3_PHYADDRPOINTER_REG_31_;
  assign new_P3_U7365 = ~new_P3_U7094 | ~P3_REIP_REG_31_;
  assign new_P3_U7366 = ~P3_DATAWIDTH_REG_1_ | ~P3_DATAWIDTH_REG_0_;
  assign new_P3_U7367 = P3_REIP_REG_1_ | P3_REIP_REG_0_;
  assign new_P3_U7368 = ~new_P3_U4285;
  assign new_P3_U7369 = ~P3_FLUSH_REG | ~new_P3_U4285;
  assign new_P3_U7370 = ~new_P3_U4623 | ~new_P3_U2390;
  assign new_P3_U7371 = ~new_P3_U2453 | ~new_P3_U2630;
  assign new_P3_U7372 = ~new_P3_U3123 | ~new_P3_U7371;
  assign new_P3_U7373 = ~new_P3_U7372 | ~new_P3_U3121;
  assign new_P3_U7374 = ~new_P3_U4287;
  assign new_P3_U7375 = ~new_P3_U4296 | ~new_P3_U2631;
  assign new_P3_U7376 = ~new_P3_U3112 | ~new_P3_U3118;
  assign new_P3_U7377 = ~new_P3_U4150 | ~P3_STATE2_REG_2_ | ~new_P3_U7919;
  assign new_P3_U7378 = ~P3_STATE2_REG_0_ | ~new_P3_U7377;
  assign new_P3_U7379 = ~new_P3_U3125 | ~new_P3_U7378;
  assign new_P3_U7380 = ~new_P3_U2390 | ~new_P3_U2604;
  assign new_P3_U7381 = ~P3_CODEFETCH_REG | ~new_P3_U7380;
  assign new_P3_U7382 = ~new_P3_U4347 | ~P3_STATE2_REG_0_;
  assign new_P3_U7383 = ~P3_ADS_N_REG | ~P3_STATE_REG_0_;
  assign new_P3_U7384 = ~new_P3_U4288;
  assign new_P3_U7385 = ~new_P3_U3114 | ~P3_STATE2_REG_2_ | ~new_P3_U3111;
  assign new_P3_U7386 = ~new_P3_U4488 | ~P3_STATE2_REG_2_;
  assign new_P3_U7387 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__7_;
  assign new_P3_U7388 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__7_;
  assign new_P3_U7389 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__7_;
  assign new_P3_U7390 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__7_;
  assign new_P3_U7391 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__7_;
  assign new_P3_U7392 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__7_;
  assign new_P3_U7393 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__7_;
  assign new_P3_U7394 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__7_;
  assign new_P3_U7395 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__7_;
  assign new_P3_U7396 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__7_;
  assign new_P3_U7397 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__7_;
  assign new_P3_U7398 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__7_;
  assign new_P3_U7399 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__7_;
  assign new_P3_U7400 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__7_;
  assign new_P3_U7401 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__7_;
  assign new_P3_U7402 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__7_;
  assign new_P3_U7403 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__6_;
  assign new_P3_U7404 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__6_;
  assign new_P3_U7405 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__6_;
  assign new_P3_U7406 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__6_;
  assign new_P3_U7407 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__6_;
  assign new_P3_U7408 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__6_;
  assign new_P3_U7409 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__6_;
  assign new_P3_U7410 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__6_;
  assign new_P3_U7411 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__6_;
  assign new_P3_U7412 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__6_;
  assign new_P3_U7413 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__6_;
  assign new_P3_U7414 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__6_;
  assign new_P3_U7415 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__6_;
  assign new_P3_U7416 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__6_;
  assign new_P3_U7417 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__6_;
  assign new_P3_U7418 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__6_;
  assign new_P3_U7419 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__5_;
  assign new_P3_U7420 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__5_;
  assign new_P3_U7421 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__5_;
  assign new_P3_U7422 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__5_;
  assign new_P3_U7423 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__5_;
  assign new_P3_U7424 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__5_;
  assign new_P3_U7425 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__5_;
  assign new_P3_U7426 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__5_;
  assign new_P3_U7427 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__5_;
  assign new_P3_U7428 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__5_;
  assign new_P3_U7429 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__5_;
  assign new_P3_U7430 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__5_;
  assign new_P3_U7431 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__5_;
  assign new_P3_U7432 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__5_;
  assign new_P3_U7433 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__5_;
  assign new_P3_U7434 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__5_;
  assign new_P3_U7435 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__4_;
  assign new_P3_U7436 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__4_;
  assign new_P3_U7437 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__4_;
  assign new_P3_U7438 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__4_;
  assign new_P3_U7439 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__4_;
  assign new_P3_U7440 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__4_;
  assign new_P3_U7441 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__4_;
  assign new_P3_U7442 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__4_;
  assign new_P3_U7443 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__4_;
  assign new_P3_U7444 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__4_;
  assign new_P3_U7445 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__4_;
  assign new_P3_U7446 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__4_;
  assign new_P3_U7447 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__4_;
  assign new_P3_U7448 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__4_;
  assign new_P3_U7449 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__4_;
  assign new_P3_U7450 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__4_;
  assign new_P3_U7451 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__3_;
  assign new_P3_U7452 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__3_;
  assign new_P3_U7453 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__3_;
  assign new_P3_U7454 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__3_;
  assign new_P3_U7455 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__3_;
  assign new_P3_U7456 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__3_;
  assign new_P3_U7457 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__3_;
  assign new_P3_U7458 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__3_;
  assign new_P3_U7459 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__3_;
  assign new_P3_U7460 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__3_;
  assign new_P3_U7461 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__3_;
  assign new_P3_U7462 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__3_;
  assign new_P3_U7463 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__3_;
  assign new_P3_U7464 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__3_;
  assign new_P3_U7465 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__3_;
  assign new_P3_U7466 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__3_;
  assign new_P3_U7467 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__2_;
  assign new_P3_U7468 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__2_;
  assign new_P3_U7469 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__2_;
  assign new_P3_U7470 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__2_;
  assign new_P3_U7471 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__2_;
  assign new_P3_U7472 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__2_;
  assign new_P3_U7473 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__2_;
  assign new_P3_U7474 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__2_;
  assign new_P3_U7475 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__2_;
  assign new_P3_U7476 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__2_;
  assign new_P3_U7477 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__2_;
  assign new_P3_U7478 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__2_;
  assign new_P3_U7479 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__2_;
  assign new_P3_U7480 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__2_;
  assign new_P3_U7481 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__2_;
  assign new_P3_U7482 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__2_;
  assign new_P3_U7483 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__1_;
  assign new_P3_U7484 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__1_;
  assign new_P3_U7485 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__1_;
  assign new_P3_U7486 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__1_;
  assign new_P3_U7487 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__1_;
  assign new_P3_U7488 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__1_;
  assign new_P3_U7489 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__1_;
  assign new_P3_U7490 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__1_;
  assign new_P3_U7491 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__1_;
  assign new_P3_U7492 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__1_;
  assign new_P3_U7493 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__1_;
  assign new_P3_U7494 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__1_;
  assign new_P3_U7495 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__1_;
  assign new_P3_U7496 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__1_;
  assign new_P3_U7497 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__1_;
  assign new_P3_U7498 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__1_;
  assign new_P3_U7499 = ~new_P3_U2542 | ~P3_INSTQUEUE_REG_15__0_;
  assign new_P3_U7500 = ~new_P3_U2541 | ~P3_INSTQUEUE_REG_14__0_;
  assign new_P3_U7501 = ~new_P3_U2540 | ~P3_INSTQUEUE_REG_13__0_;
  assign new_P3_U7502 = ~new_P3_U2539 | ~P3_INSTQUEUE_REG_12__0_;
  assign new_P3_U7503 = ~new_P3_U2537 | ~P3_INSTQUEUE_REG_11__0_;
  assign new_P3_U7504 = ~new_P3_U2536 | ~P3_INSTQUEUE_REG_10__0_;
  assign new_P3_U7505 = ~new_P3_U2535 | ~P3_INSTQUEUE_REG_9__0_;
  assign new_P3_U7506 = ~new_P3_U2534 | ~P3_INSTQUEUE_REG_8__0_;
  assign new_P3_U7507 = ~new_P3_U2532 | ~P3_INSTQUEUE_REG_7__0_;
  assign new_P3_U7508 = ~new_P3_U2531 | ~P3_INSTQUEUE_REG_6__0_;
  assign new_P3_U7509 = ~new_P3_U2530 | ~P3_INSTQUEUE_REG_5__0_;
  assign new_P3_U7510 = ~new_P3_U2529 | ~P3_INSTQUEUE_REG_4__0_;
  assign new_P3_U7511 = ~new_P3_U2527 | ~P3_INSTQUEUE_REG_3__0_;
  assign new_P3_U7512 = ~new_P3_U2525 | ~P3_INSTQUEUE_REG_2__0_;
  assign new_P3_U7513 = ~new_P3_U2523 | ~P3_INSTQUEUE_REG_1__0_;
  assign new_P3_U7514 = ~new_P3_U2521 | ~P3_INSTQUEUE_REG_0__0_;
  assign new_P3_U7515 = ~new_P3_U4470 | ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_U7516 = ~new_P3_U3266;
  assign new_P3_U7517 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__7_;
  assign new_P3_U7518 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__7_;
  assign new_P3_U7519 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__7_;
  assign new_P3_U7520 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__7_;
  assign new_P3_U7521 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__7_;
  assign new_P3_U7522 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__7_;
  assign new_P3_U7523 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__7_;
  assign new_P3_U7524 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__7_;
  assign new_P3_U7525 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__7_;
  assign new_P3_U7526 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__7_;
  assign new_P3_U7527 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__7_;
  assign new_P3_U7528 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__7_;
  assign new_P3_U7529 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__7_;
  assign new_P3_U7530 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__7_;
  assign new_P3_U7531 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__7_;
  assign new_P3_U7532 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__7_;
  assign new_P3_U7533 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__6_;
  assign new_P3_U7534 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__6_;
  assign new_P3_U7535 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__6_;
  assign new_P3_U7536 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__6_;
  assign new_P3_U7537 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__6_;
  assign new_P3_U7538 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__6_;
  assign new_P3_U7539 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__6_;
  assign new_P3_U7540 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__6_;
  assign new_P3_U7541 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__6_;
  assign new_P3_U7542 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__6_;
  assign new_P3_U7543 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__6_;
  assign new_P3_U7544 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__6_;
  assign new_P3_U7545 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__6_;
  assign new_P3_U7546 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__6_;
  assign new_P3_U7547 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__6_;
  assign new_P3_U7548 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__6_;
  assign new_P3_U7549 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__5_;
  assign new_P3_U7550 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__5_;
  assign new_P3_U7551 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__5_;
  assign new_P3_U7552 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__5_;
  assign new_P3_U7553 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__5_;
  assign new_P3_U7554 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__5_;
  assign new_P3_U7555 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__5_;
  assign new_P3_U7556 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__5_;
  assign new_P3_U7557 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__5_;
  assign new_P3_U7558 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__5_;
  assign new_P3_U7559 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__5_;
  assign new_P3_U7560 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__5_;
  assign new_P3_U7561 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__5_;
  assign new_P3_U7562 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__5_;
  assign new_P3_U7563 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__5_;
  assign new_P3_U7564 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__5_;
  assign new_P3_U7565 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__4_;
  assign new_P3_U7566 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__4_;
  assign new_P3_U7567 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__4_;
  assign new_P3_U7568 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__4_;
  assign new_P3_U7569 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__4_;
  assign new_P3_U7570 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__4_;
  assign new_P3_U7571 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__4_;
  assign new_P3_U7572 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__4_;
  assign new_P3_U7573 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__4_;
  assign new_P3_U7574 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__4_;
  assign new_P3_U7575 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__4_;
  assign new_P3_U7576 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__4_;
  assign new_P3_U7577 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__4_;
  assign new_P3_U7578 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__4_;
  assign new_P3_U7579 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__4_;
  assign new_P3_U7580 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__4_;
  assign new_P3_U7581 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__3_;
  assign new_P3_U7582 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__3_;
  assign new_P3_U7583 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__3_;
  assign new_P3_U7584 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__3_;
  assign new_P3_U7585 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__3_;
  assign new_P3_U7586 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__3_;
  assign new_P3_U7587 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__3_;
  assign new_P3_U7588 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__3_;
  assign new_P3_U7589 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__3_;
  assign new_P3_U7590 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__3_;
  assign new_P3_U7591 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__3_;
  assign new_P3_U7592 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__3_;
  assign new_P3_U7593 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__3_;
  assign new_P3_U7594 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__3_;
  assign new_P3_U7595 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__3_;
  assign new_P3_U7596 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__3_;
  assign new_P3_U7597 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__2_;
  assign new_P3_U7598 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__2_;
  assign new_P3_U7599 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__2_;
  assign new_P3_U7600 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__2_;
  assign new_P3_U7601 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__2_;
  assign new_P3_U7602 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__2_;
  assign new_P3_U7603 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__2_;
  assign new_P3_U7604 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__2_;
  assign new_P3_U7605 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__2_;
  assign new_P3_U7606 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__2_;
  assign new_P3_U7607 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__2_;
  assign new_P3_U7608 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__2_;
  assign new_P3_U7609 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__2_;
  assign new_P3_U7610 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__2_;
  assign new_P3_U7611 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__2_;
  assign new_P3_U7612 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__2_;
  assign new_P3_U7613 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__1_;
  assign new_P3_U7614 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__1_;
  assign new_P3_U7615 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__1_;
  assign new_P3_U7616 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__1_;
  assign new_P3_U7617 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__1_;
  assign new_P3_U7618 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__1_;
  assign new_P3_U7619 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__1_;
  assign new_P3_U7620 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__1_;
  assign new_P3_U7621 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__1_;
  assign new_P3_U7622 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__1_;
  assign new_P3_U7623 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__1_;
  assign new_P3_U7624 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__1_;
  assign new_P3_U7625 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__1_;
  assign new_P3_U7626 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__1_;
  assign new_P3_U7627 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__1_;
  assign new_P3_U7628 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__1_;
  assign new_P3_U7629 = ~new_P3_U2562 | ~P3_INSTQUEUE_REG_0__0_;
  assign new_P3_U7630 = ~new_P3_U2561 | ~P3_INSTQUEUE_REG_1__0_;
  assign new_P3_U7631 = ~new_P3_U2560 | ~P3_INSTQUEUE_REG_2__0_;
  assign new_P3_U7632 = ~new_P3_U2559 | ~P3_INSTQUEUE_REG_3__0_;
  assign new_P3_U7633 = ~new_P3_U2557 | ~P3_INSTQUEUE_REG_4__0_;
  assign new_P3_U7634 = ~new_P3_U2556 | ~P3_INSTQUEUE_REG_5__0_;
  assign new_P3_U7635 = ~new_P3_U2555 | ~P3_INSTQUEUE_REG_6__0_;
  assign new_P3_U7636 = ~new_P3_U2554 | ~P3_INSTQUEUE_REG_7__0_;
  assign new_P3_U7637 = ~new_P3_U2552 | ~P3_INSTQUEUE_REG_8__0_;
  assign new_P3_U7638 = ~new_P3_U2551 | ~P3_INSTQUEUE_REG_9__0_;
  assign new_P3_U7639 = ~new_P3_U2550 | ~P3_INSTQUEUE_REG_10__0_;
  assign new_P3_U7640 = ~new_P3_U2549 | ~P3_INSTQUEUE_REG_11__0_;
  assign new_P3_U7641 = ~new_P3_U2547 | ~P3_INSTQUEUE_REG_12__0_;
  assign new_P3_U7642 = ~new_P3_U2546 | ~P3_INSTQUEUE_REG_13__0_;
  assign new_P3_U7643 = ~new_P3_U2545 | ~P3_INSTQUEUE_REG_14__0_;
  assign new_P3_U7644 = ~new_P3_U2544 | ~P3_INSTQUEUE_REG_15__0_;
  assign new_P3_U7645 = ~new_P3_U4289;
  assign new_P3_U7646 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__7_;
  assign new_P3_U7647 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__7_;
  assign new_P3_U7648 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__7_;
  assign new_P3_U7649 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__7_;
  assign new_P3_U7650 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__7_;
  assign new_P3_U7651 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__7_;
  assign new_P3_U7652 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__7_;
  assign new_P3_U7653 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__7_;
  assign new_P3_U7654 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__7_;
  assign new_P3_U7655 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__7_;
  assign new_P3_U7656 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__7_;
  assign new_P3_U7657 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__7_;
  assign new_P3_U7658 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__7_;
  assign new_P3_U7659 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__7_;
  assign new_P3_U7660 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__7_;
  assign new_P3_U7661 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__7_;
  assign new_P3_U7662 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__6_;
  assign new_P3_U7663 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__6_;
  assign new_P3_U7664 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__6_;
  assign new_P3_U7665 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__6_;
  assign new_P3_U7666 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__6_;
  assign new_P3_U7667 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__6_;
  assign new_P3_U7668 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__6_;
  assign new_P3_U7669 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__6_;
  assign new_P3_U7670 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__6_;
  assign new_P3_U7671 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__6_;
  assign new_P3_U7672 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__6_;
  assign new_P3_U7673 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__6_;
  assign new_P3_U7674 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__6_;
  assign new_P3_U7675 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__6_;
  assign new_P3_U7676 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__6_;
  assign new_P3_U7677 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__6_;
  assign new_P3_U7678 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__5_;
  assign new_P3_U7679 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__5_;
  assign new_P3_U7680 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__5_;
  assign new_P3_U7681 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__5_;
  assign new_P3_U7682 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__5_;
  assign new_P3_U7683 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__5_;
  assign new_P3_U7684 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__5_;
  assign new_P3_U7685 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__5_;
  assign new_P3_U7686 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__5_;
  assign new_P3_U7687 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__5_;
  assign new_P3_U7688 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__5_;
  assign new_P3_U7689 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__5_;
  assign new_P3_U7690 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__5_;
  assign new_P3_U7691 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__5_;
  assign new_P3_U7692 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__5_;
  assign new_P3_U7693 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__5_;
  assign new_P3_U7694 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__4_;
  assign new_P3_U7695 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__4_;
  assign new_P3_U7696 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__4_;
  assign new_P3_U7697 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__4_;
  assign new_P3_U7698 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__4_;
  assign new_P3_U7699 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__4_;
  assign new_P3_U7700 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__4_;
  assign new_P3_U7701 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__4_;
  assign new_P3_U7702 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__4_;
  assign new_P3_U7703 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__4_;
  assign new_P3_U7704 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__4_;
  assign new_P3_U7705 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__4_;
  assign new_P3_U7706 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__4_;
  assign new_P3_U7707 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__4_;
  assign new_P3_U7708 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__4_;
  assign new_P3_U7709 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__4_;
  assign new_P3_U7710 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__3_;
  assign new_P3_U7711 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__3_;
  assign new_P3_U7712 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__3_;
  assign new_P3_U7713 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__3_;
  assign new_P3_U7714 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__3_;
  assign new_P3_U7715 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__3_;
  assign new_P3_U7716 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__3_;
  assign new_P3_U7717 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__3_;
  assign new_P3_U7718 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__3_;
  assign new_P3_U7719 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__3_;
  assign new_P3_U7720 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__3_;
  assign new_P3_U7721 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__3_;
  assign new_P3_U7722 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__3_;
  assign new_P3_U7723 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__3_;
  assign new_P3_U7724 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__3_;
  assign new_P3_U7725 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__3_;
  assign new_P3_U7726 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__2_;
  assign new_P3_U7727 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__2_;
  assign new_P3_U7728 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__2_;
  assign new_P3_U7729 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__2_;
  assign new_P3_U7730 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__2_;
  assign new_P3_U7731 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__2_;
  assign new_P3_U7732 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__2_;
  assign new_P3_U7733 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__2_;
  assign new_P3_U7734 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__2_;
  assign new_P3_U7735 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__2_;
  assign new_P3_U7736 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__2_;
  assign new_P3_U7737 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__2_;
  assign new_P3_U7738 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__2_;
  assign new_P3_U7739 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__2_;
  assign new_P3_U7740 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__2_;
  assign new_P3_U7741 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__2_;
  assign new_P3_U7742 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__1_;
  assign new_P3_U7743 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__1_;
  assign new_P3_U7744 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__1_;
  assign new_P3_U7745 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__1_;
  assign new_P3_U7746 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__1_;
  assign new_P3_U7747 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__1_;
  assign new_P3_U7748 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__1_;
  assign new_P3_U7749 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__1_;
  assign new_P3_U7750 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__1_;
  assign new_P3_U7751 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__1_;
  assign new_P3_U7752 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__1_;
  assign new_P3_U7753 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__1_;
  assign new_P3_U7754 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__1_;
  assign new_P3_U7755 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__1_;
  assign new_P3_U7756 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__1_;
  assign new_P3_U7757 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__1_;
  assign new_P3_U7758 = ~new_P3_U2582 | ~P3_INSTQUEUE_REG_8__0_;
  assign new_P3_U7759 = ~new_P3_U2581 | ~P3_INSTQUEUE_REG_9__0_;
  assign new_P3_U7760 = ~new_P3_U2580 | ~P3_INSTQUEUE_REG_10__0_;
  assign new_P3_U7761 = ~new_P3_U2579 | ~P3_INSTQUEUE_REG_11__0_;
  assign new_P3_U7762 = ~new_P3_U2577 | ~P3_INSTQUEUE_REG_12__0_;
  assign new_P3_U7763 = ~new_P3_U2576 | ~P3_INSTQUEUE_REG_13__0_;
  assign new_P3_U7764 = ~new_P3_U2575 | ~P3_INSTQUEUE_REG_14__0_;
  assign new_P3_U7765 = ~new_P3_U2574 | ~P3_INSTQUEUE_REG_15__0_;
  assign new_P3_U7766 = ~new_P3_U2572 | ~P3_INSTQUEUE_REG_0__0_;
  assign new_P3_U7767 = ~new_P3_U2571 | ~P3_INSTQUEUE_REG_1__0_;
  assign new_P3_U7768 = ~new_P3_U2570 | ~P3_INSTQUEUE_REG_2__0_;
  assign new_P3_U7769 = ~new_P3_U2569 | ~P3_INSTQUEUE_REG_3__0_;
  assign new_P3_U7770 = ~new_P3_U2567 | ~P3_INSTQUEUE_REG_4__0_;
  assign new_P3_U7771 = ~new_P3_U2566 | ~P3_INSTQUEUE_REG_5__0_;
  assign new_P3_U7772 = ~new_P3_U2565 | ~P3_INSTQUEUE_REG_6__0_;
  assign new_P3_U7773 = ~new_P3_U2564 | ~P3_INSTQUEUE_REG_7__0_;
  assign new_P3_U7774 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_U3097;
  assign new_P3_U7775 = ~new_P3_U3268;
  assign new_P3_U7776 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__7_;
  assign new_P3_U7777 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__7_;
  assign new_P3_U7778 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__7_;
  assign new_P3_U7779 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__7_;
  assign new_P3_U7780 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__7_;
  assign new_P3_U7781 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__7_;
  assign new_P3_U7782 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__7_;
  assign new_P3_U7783 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__7_;
  assign new_P3_U7784 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__7_;
  assign new_P3_U7785 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__7_;
  assign new_P3_U7786 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__7_;
  assign new_P3_U7787 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__7_;
  assign new_P3_U7788 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__7_;
  assign new_P3_U7789 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__7_;
  assign new_P3_U7790 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__7_;
  assign new_P3_U7791 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__7_;
  assign new_P3_U7792 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__6_;
  assign new_P3_U7793 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__6_;
  assign new_P3_U7794 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__6_;
  assign new_P3_U7795 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__6_;
  assign new_P3_U7796 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__6_;
  assign new_P3_U7797 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__6_;
  assign new_P3_U7798 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__6_;
  assign new_P3_U7799 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__6_;
  assign new_P3_U7800 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__6_;
  assign new_P3_U7801 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__6_;
  assign new_P3_U7802 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__6_;
  assign new_P3_U7803 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__6_;
  assign new_P3_U7804 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__6_;
  assign new_P3_U7805 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__6_;
  assign new_P3_U7806 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__6_;
  assign new_P3_U7807 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__6_;
  assign new_P3_U7808 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__5_;
  assign new_P3_U7809 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__5_;
  assign new_P3_U7810 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__5_;
  assign new_P3_U7811 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__5_;
  assign new_P3_U7812 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__5_;
  assign new_P3_U7813 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__5_;
  assign new_P3_U7814 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__5_;
  assign new_P3_U7815 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__5_;
  assign new_P3_U7816 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__5_;
  assign new_P3_U7817 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__5_;
  assign new_P3_U7818 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__5_;
  assign new_P3_U7819 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__5_;
  assign new_P3_U7820 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__5_;
  assign new_P3_U7821 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__5_;
  assign new_P3_U7822 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__5_;
  assign new_P3_U7823 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__5_;
  assign new_P3_U7824 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__4_;
  assign new_P3_U7825 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__4_;
  assign new_P3_U7826 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__4_;
  assign new_P3_U7827 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__4_;
  assign new_P3_U7828 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__4_;
  assign new_P3_U7829 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__4_;
  assign new_P3_U7830 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__4_;
  assign new_P3_U7831 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__4_;
  assign new_P3_U7832 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__4_;
  assign new_P3_U7833 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__4_;
  assign new_P3_U7834 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__4_;
  assign new_P3_U7835 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__4_;
  assign new_P3_U7836 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__4_;
  assign new_P3_U7837 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__4_;
  assign new_P3_U7838 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__4_;
  assign new_P3_U7839 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__4_;
  assign new_P3_U7840 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__3_;
  assign new_P3_U7841 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__3_;
  assign new_P3_U7842 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__3_;
  assign new_P3_U7843 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__3_;
  assign new_P3_U7844 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__3_;
  assign new_P3_U7845 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__3_;
  assign new_P3_U7846 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__3_;
  assign new_P3_U7847 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__3_;
  assign new_P3_U7848 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__3_;
  assign new_P3_U7849 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__3_;
  assign new_P3_U7850 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__3_;
  assign new_P3_U7851 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__3_;
  assign new_P3_U7852 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__3_;
  assign new_P3_U7853 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__3_;
  assign new_P3_U7854 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__3_;
  assign new_P3_U7855 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__3_;
  assign new_P3_U7856 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__2_;
  assign new_P3_U7857 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__2_;
  assign new_P3_U7858 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__2_;
  assign new_P3_U7859 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__2_;
  assign new_P3_U7860 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__2_;
  assign new_P3_U7861 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__2_;
  assign new_P3_U7862 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__2_;
  assign new_P3_U7863 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__2_;
  assign new_P3_U7864 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__2_;
  assign new_P3_U7865 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__2_;
  assign new_P3_U7866 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__2_;
  assign new_P3_U7867 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__2_;
  assign new_P3_U7868 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__2_;
  assign new_P3_U7869 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__2_;
  assign new_P3_U7870 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__2_;
  assign new_P3_U7871 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__2_;
  assign new_P3_U7872 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__1_;
  assign new_P3_U7873 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__1_;
  assign new_P3_U7874 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__1_;
  assign new_P3_U7875 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__1_;
  assign new_P3_U7876 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__1_;
  assign new_P3_U7877 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__1_;
  assign new_P3_U7878 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__1_;
  assign new_P3_U7879 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__1_;
  assign new_P3_U7880 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__1_;
  assign new_P3_U7881 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__1_;
  assign new_P3_U7882 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__1_;
  assign new_P3_U7883 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__1_;
  assign new_P3_U7884 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__1_;
  assign new_P3_U7885 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__1_;
  assign new_P3_U7886 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__1_;
  assign new_P3_U7887 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__1_;
  assign new_P3_U7888 = ~new_P3_U2600 | ~P3_INSTQUEUE_REG_8__0_;
  assign new_P3_U7889 = ~new_P3_U2599 | ~P3_INSTQUEUE_REG_9__0_;
  assign new_P3_U7890 = ~new_P3_U2598 | ~P3_INSTQUEUE_REG_10__0_;
  assign new_P3_U7891 = ~new_P3_U2597 | ~P3_INSTQUEUE_REG_11__0_;
  assign new_P3_U7892 = ~new_P3_U2595 | ~P3_INSTQUEUE_REG_12__0_;
  assign new_P3_U7893 = ~new_P3_U2594 | ~P3_INSTQUEUE_REG_13__0_;
  assign new_P3_U7894 = ~new_P3_U2593 | ~P3_INSTQUEUE_REG_14__0_;
  assign new_P3_U7895 = ~new_P3_U2592 | ~P3_INSTQUEUE_REG_15__0_;
  assign new_P3_U7896 = ~new_P3_U2591 | ~P3_INSTQUEUE_REG_0__0_;
  assign new_P3_U7897 = ~new_P3_U2590 | ~P3_INSTQUEUE_REG_1__0_;
  assign new_P3_U7898 = ~new_P3_U2589 | ~P3_INSTQUEUE_REG_2__0_;
  assign new_P3_U7899 = ~new_P3_U2588 | ~P3_INSTQUEUE_REG_3__0_;
  assign new_P3_U7900 = ~new_P3_U2586 | ~P3_INSTQUEUE_REG_4__0_;
  assign new_P3_U7901 = ~new_P3_U2585 | ~P3_INSTQUEUE_REG_5__0_;
  assign new_P3_U7902 = ~new_P3_U2584 | ~P3_INSTQUEUE_REG_6__0_;
  assign new_P3_U7903 = ~new_P3_U2583 | ~P3_INSTQUEUE_REG_7__0_;
  assign new_P3_U7904 = ~P3_STATE_REG_0_ | ~new_P3_U4292;
  assign new_P3_U7905 = new_U209 | P3_STATE2_REG_2_;
  assign new_P3_U7906 = ~new_P3_U3939 | ~new_P3_U6397;
  assign new_P3_U7907 = ~new_P3_U4134 | ~new_P3_U2603;
  assign new_P3_U7908 = ~new_P3_U2404 | ~new_P3_U3256;
  assign new_P3_U7909 = ~new_P3_U2392 | ~new_P3_U7096;
  assign new_P3_U7910 = ~new_P3_U7909 | ~new_P3_U7908 | ~new_P3_U4317;
  assign new_P3_U7911 = ~new_P3_U3086;
  assign new_P3_U7912 = ~new_P3_U7911 | ~new_P3_U3088;
  assign new_P3_U7913 = ~new_P3_U4446 | ~new_P3_U4449 | ~P3_STATE_REG_1_;
  assign new_P3_U7914 = ~P3_STATE_REG_2_ | ~new_P3_U7904;
  assign new_P3_U7915 = ~P3_STATE_REG_1_ | ~new_P3_U4446;
  assign new_P3_U7916 = ~new_P3_U4505 | ~new_P3_U3106;
  assign new_P3_U7917 = ~new_P3_U4488 | ~new_P3_U4522;
  assign new_P3_U7918 = ~new_P3_U3208 | ~new_P3_U3219;
  assign new_P3_U7919 = ~new_P3_U7376 | ~new_P3_U3105;
  assign new_P3_U7920 = ~P3_BE_N_REG_3_ | ~new_P3_U3077;
  assign new_P3_U7921 = ~P3_BYTEENABLE_REG_3_ | ~new_P3_U4308;
  assign new_P3_U7922 = ~P3_BE_N_REG_2_ | ~new_P3_U3077;
  assign new_P3_U7923 = ~P3_BYTEENABLE_REG_2_ | ~new_P3_U4308;
  assign new_P3_U7924 = ~P3_BE_N_REG_1_ | ~new_P3_U3077;
  assign new_P3_U7925 = ~P3_BYTEENABLE_REG_1_ | ~new_P3_U4308;
  assign new_P3_U7926 = ~P3_BE_N_REG_0_ | ~new_P3_U3077;
  assign new_P3_U7927 = ~P3_BYTEENABLE_REG_0_ | ~new_P3_U4308;
  assign new_P3_U7928 = ~new_P3_U3079 | ~P3_STATE_REG_0_ | ~P3_REQUESTPENDING_REG;
  assign new_P3_U7929 = ~P3_STATE_REG_2_ | ~new_P3_U3086;
  assign new_P3_U7930 = ~new_P3_U7929 | ~new_P3_U7928;
  assign new_P3_U7931 = ~P3_STATE_REG_1_ | ~new_P3_U7914 | ~new_P3_U4449;
  assign new_P3_U7932 = ~new_P3_U7930 | ~new_P3_U3076;
  assign new_P3_U7933 = ~P3_STATE_REG_2_ | ~P3_STATE_REG_0_ | ~new_P3_U3087;
  assign new_P3_U7934 = ~new_P3_U4459 | ~new_P3_U3079;
  assign new_P3_U7935 = P3_STATE_REG_0_ | P3_STATE_REG_1_;
  assign new_P3_U7936 = ~P3_STATE_REG_0_ | ~new_P3_U4346;
  assign new_P3_U7937 = ~new_P3_U3278;
  assign new_P3_U7938 = ~new_P3_U7937 | ~P3_DATAWIDTH_REG_0_;
  assign new_P3_U7939 = ~new_P3_U3279 | ~new_P3_U3278;
  assign new_P3_U7940 = ~new_P3_U3278 | ~new_P3_U4464;
  assign new_P3_U7941 = ~new_P3_U7937 | ~P3_DATAWIDTH_REG_1_;
  assign new_P3_U7942 = ~new_P3_U4505 | ~new_P3_U3211;
  assign new_P3_U7943 = ~new_P3_U3104 | ~new_P3_U3214;
  assign new_P3_U7944 = ~new_P3_U4505 | ~new_P3_U3213;
  assign new_P3_U7945 = ~new_P3_U3104 | ~new_P3_U3210;
  assign new_P3_U7946 = ~new_P3_U4539 | ~new_P3_U4618;
  assign new_P3_U7947 = ~new_P3_U4620 | ~new_P3_U3101;
  assign new_P3_U7948 = ~new_P3_U4281 | ~new_P3_U4617;
  assign new_P3_U7949 = ~new_P3_U4622 | ~new_P3_U4624;
  assign new_P3_U7950 = ~new_P3_U4505 | ~new_P3_U3237;
  assign new_P3_U7951 = ~new_P3_U3104 | ~new_P3_U3238;
  assign new_P3_U7952 = ~P3_STATE2_REG_0_ | ~new_P3_U4627;
  assign new_P3_U7953 = ~new_P3_U4628 | ~new_P3_U3121;
  assign new_P3_U7954 = ~P3_STATE2_REG_3_ | ~new_P3_U3122;
  assign new_P3_U7955 = ~new_P3_U2453 | ~new_P3_U4630;
  assign new_P3_U7956 = P3_STATEBS16_REG | P3_STATE2_REG_0_;
  assign new_P3_U7957 = ~P3_STATE2_REG_0_ | ~new_P3_U7905;
  assign new_P3_U7958 = ~P3_STATE2_REG_0_ | ~new_P3_U4638;
  assign new_P3_U7959 = ~new_P3_U3121 | ~new_P3_U4637 | ~new_P3_U4629;
  assign new_P3_U7960 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_U3130;
  assign new_P3_U7961 = ~new_P3_U4648 | ~new_P3_U3131;
  assign new_P3_U7962 = ~new_P3_U3269;
  assign new_P3_U7963 = ~new_P3_U7962 | ~new_P3_U4653;
  assign new_P3_U7964 = ~new_P3_U3269 | ~new_P3_U3138;
  assign new_P3_U7965 = ~new_P3_U3270;
  assign new_P3_U7966 = ~new_P3_U7965 | ~new_P3_U4657;
  assign new_P3_U7967 = ~new_P3_U3270 | ~new_P3_U3140;
  assign new_P3_U7968 = ~new_P3_U3271;
  assign new_P3_U7969 = ~new_P3_U3109 | ~new_P3_U3101;
  assign new_P3_U7970 = ~new_P3_U4539 | ~new_P3_U5483;
  assign new_P3_U7971 = ~new_P3_U3283 | ~new_P3_U4283;
  assign new_P3_U7972 = ~new_P3_U5499 | ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_U7973 = ~new_P3_U3218 | ~new_P3_U3107;
  assign new_P3_U7974 = ~new_P3_U4573 | ~new_P3_U4590;
  assign new_P3_U7975 = ~new_P3_U4539 | ~new_P3_U5512;
  assign new_P3_U7976 = ~new_P3_U5515 | ~new_P3_U3101;
  assign new_P3_U7977 = ~new_P3_U3110 | ~new_P3_U4556 | ~new_P3_U5517;
  assign new_P3_U7978 = ~new_P3_U4590 | ~new_P3_U5513 | ~new_P3_U3107;
  assign new_P3_U7979 = ~new_P3_U5499 | ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_U7980 = ~new_P3_U5546 | ~new_P3_U4283;
  assign new_P3_U7981 = ~new_P3_U3094 | ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U3221;
  assign new_P3_U7982 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_U5531 | ~new_P3_U3097;
  assign new_P3_U7983 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_U4284;
  assign new_P3_U7984 = ~new_P3_SUB_580_U6 | ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_U7985 = ~new_P3_U3287;
  assign new_P3_U7986 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_U4284;
  assign new_P3_U7987 = ~P3_INSTADDRPOINTER_REG_0_ | ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_U7988 = ~new_P3_U3286;
  assign new_P3_U7989 = ~new_P3_U5499 | ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_U7990 = ~new_P3_U5557 | ~new_P3_U4283;
  assign new_P3_U7991 = ~new_P3_U5499 | ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_U7992 = ~new_P3_U5570 | ~new_P3_U4283;
  assign new_P3_U7993 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_U3221;
  assign new_P3_U7994 = ~new_P3_U5571 | ~new_P3_U3093;
  assign new_P3_U7995 = ~new_P3_U5499 | ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_U7996 = ~new_P3_U5577 | ~new_P3_U4283;
  assign new_P3_U7997 = ~new_P3_U7968 | ~new_P3_U4647;
  assign new_P3_U7998 = ~new_P3_U3271 | ~new_P3_U3143;
  assign new_P3_U7999 = ~new_P3_U7998 | ~new_P3_U7997;
  assign new_P3_U8000 = ~new_P3_U5622 | ~new_P3_U3104;
  assign new_P3_U8001 = ~new_P3_U4505 | ~new_P3_U5619;
  assign new_P3_U8002 = ~P3_BYTEENABLE_REG_3_ | ~new_P3_U3261;
  assign new_P3_U8003 = ~new_P3_U3291 | ~new_P3_U4307;
  assign new_P3_U8004 = P3_DATAWIDTH_REG_0_ | P3_DATAWIDTH_REG_1_;
  assign new_P3_U8005 = ~P3_DATAWIDTH_REG_0_ | ~new_P3_U3240;
  assign new_P3_U8006 = ~new_P3_U8005 | ~new_P3_U8004;
  assign new_P3_U8007 = ~new_P3_U8006 | ~new_P3_U3081;
  assign new_P3_U8008 = ~P3_REIP_REG_0_ | ~P3_REIP_REG_1_;
  assign new_P3_U8009 = ~new_P3_U8008 | ~new_P3_U8007;
  assign new_P3_U8010 = ~P3_BYTEENABLE_REG_2_ | ~new_P3_U3261;
  assign new_P3_U8011 = ~new_P3_U8009 | ~new_P3_U4307;
  assign new_P3_U8012 = ~P3_BYTEENABLE_REG_1_ | ~new_P3_U3261;
  assign new_P3_U8013 = ~new_P3_U4307 | ~P3_REIP_REG_1_;
  assign new_P3_U8014 = ~P3_BYTEENABLE_REG_0_ | ~new_P3_U3261;
  assign new_P3_U8015 = ~new_P3_U4307 | ~new_P3_U7367;
  assign new_P3_U8016 = ~new_P3_U4308 | ~new_P3_U3264;
  assign new_P3_U8017 = ~P3_W_R_N_REG | ~new_P3_U3077;
  assign new_P3_U8018 = ~new_P3_U7368 | ~new_P3_U4617;
  assign new_P3_U8019 = ~P3_MORE_REG | ~new_P3_U4285;
  assign new_P3_U8020 = ~new_P3_U7937 | ~P3_STATEBS16_REG;
  assign new_P3_U8021 = ~BS16 | ~new_P3_U3278;
  assign new_P3_U8022 = ~new_P3_U7374 | ~P3_REQUESTPENDING_REG;
  assign new_P3_U8023 = ~new_P3_U7379 | ~new_P3_U4287;
  assign new_P3_U8024 = ~new_P3_U4308 | ~new_P3_U3263;
  assign new_P3_U8025 = ~P3_D_C_N_REG | ~new_P3_U3077;
  assign new_P3_U8026 = ~P3_M_IO_N_REG | ~new_P3_U3077;
  assign new_P3_U8027 = ~P3_MEMORYFETCH_REG | ~new_P3_U4308;
  assign new_P3_U8028 = ~new_P3_U7384 | ~P3_READREQUEST_REG;
  assign new_P3_U8029 = ~new_P3_U7385 | ~new_P3_U4288;
  assign new_P3_U8030 = ~new_P3_U7384 | ~P3_MEMORYFETCH_REG;
  assign new_P3_U8031 = ~new_P3_U7386 | ~new_P3_U4288;
  assign new_P3_U8032 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_U3097;
  assign new_P3_U8033 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U3094;
  assign new_P3_U8034 = ~new_P3_U3272;
  assign new_P3_U8035 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_U4289;
  assign new_P3_U8036 = ~new_P3_U7645 | ~new_P3_U3100;
  assign new_P3_U8037 = ~new_P3_U3273;
  assign new_P3_U8038 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_U3207;
  assign new_P3_U8039 = ~P3_FLUSH_REG | ~new_P3_U3287 | ~new_P3_U3286;
  assign new_P3_U8040 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_U3207;
  assign new_P3_U8041 = ~P3_FLUSH_REG | ~new_P3_U3286 | ~new_P3_U7985;
  assign new_P3_U8042 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_U3207;
  assign new_P3_U8043 = ~new_P3_U7988 | ~P3_FLUSH_REG;
  assign new_P3_U8044 = ~new_P3_U3303 | ~new_P3_U4290;
  assign new_P3_U8045 = ~new_P3_U5496 | ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_U8046 = ~new_P3_U5496 | ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_U8047 = ~new_P3_U5542 | ~new_P3_U4290;
  assign new_P3_U8048 = ~new_P3_U5496 | ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_U8049 = ~new_P3_U5553 | ~new_P3_U4290;
  assign new_P3_U8050 = ~new_P3_U5496 | ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_U8051 = ~new_P3_U5566 | ~new_P3_U4290;
  assign new_P3_U8052 = ~new_P3_U5496 | ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_U8053 = ~new_P3_U5573 | ~new_P3_U4290;
  assign new_P1_ADD_515_U170 = ~new_P1_ADD_515_U94 | ~new_P1_ADD_515_U7;
  assign new_P1_ADD_515_U169 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_ADD_515_U6;
  assign new_P1_ADD_515_U168 = ~new_P1_ADD_515_U122 | ~new_P1_ADD_515_U92;
  assign new_P1_ADD_515_U167 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_ADD_515_U93;
  assign new_P1_ADD_515_U166 = ~new_P1_ADD_515_U101 | ~new_P1_ADD_515_U21;
  assign new_P1_ADD_515_U165 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_ADD_515_U20;
  assign new_P1_ADD_515_U164 = ~new_P1_ADD_515_U110 | ~new_P1_ADD_515_U39;
  assign new_P1_ADD_515_U163 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_ADD_515_U38;
  assign new_P1_ADD_515_U162 = ~new_P1_ADD_515_U114 | ~new_P1_ADD_515_U47;
  assign new_P1_ADD_515_U161 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_ADD_515_U46;
  assign new_P1_ADD_515_U160 = ~new_P1_ADD_515_U99 | ~new_P1_ADD_515_U17;
  assign new_P1_ADD_515_U159 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_ADD_515_U16;
  assign new_P1_ADD_515_U158 = ~new_P1_ADD_515_U96 | ~new_P1_ADD_515_U11;
  assign new_P1_ADD_515_U157 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_ADD_515_U10;
  assign new_P1_ADD_515_U156 = ~new_P1_ADD_515_U105 | ~new_P1_ADD_515_U29;
  assign new_P1_ADD_515_U155 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_ADD_515_U28;
  assign new_P1_ADD_515_U154 = ~new_P1_ADD_515_U118 | ~new_P1_ADD_515_U55;
  assign new_P1_ADD_515_U153 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_ADD_515_U54;
  assign new_P1_ADD_515_U152 = ~new_P1_ADD_515_U95 | ~new_P1_ADD_515_U9;
  assign new_P1_ADD_515_U151 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_ADD_515_U8;
  assign new_P1_ADD_515_U150 = ~new_P1_ADD_515_U106 | ~new_P1_ADD_515_U31;
  assign new_P1_ADD_515_U149 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_ADD_515_U30;
  assign new_P1_ADD_515_U148 = ~new_P1_ADD_515_U117 | ~new_P1_ADD_515_U53;
  assign new_P1_ADD_515_U147 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_ADD_515_U52;
  assign new_P1_ADD_515_U146 = ~new_P1_ADD_515_U102 | ~new_P1_ADD_515_U23;
  assign new_P1_ADD_515_U145 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_ADD_515_U22;
  assign new_P1_ADD_515_U144 = ~new_P1_ADD_515_U109 | ~new_P1_ADD_515_U37;
  assign new_P1_ADD_515_U143 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_ADD_515_U36;
  assign new_P1_ADD_515_U142 = ~new_P1_ADD_515_U113 | ~new_P1_ADD_515_U45;
  assign new_P1_ADD_515_U141 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_ADD_515_U44;
  assign new_P1_ADD_515_U140 = ~new_P1_ADD_515_U100 | ~new_P1_ADD_515_U19;
  assign new_P1_ADD_515_U139 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_ADD_515_U18;
  assign new_P1_ADD_515_U138 = ~new_P1_ADD_515_U104 | ~new_P1_ADD_515_U27;
  assign new_P1_ADD_515_U137 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_ADD_515_U26;
  assign new_P1_ADD_515_U136 = ~new_P1_ADD_515_U111 | ~new_P1_ADD_515_U41;
  assign new_P1_ADD_515_U135 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_ADD_515_U40;
  assign new_P1_ADD_515_U134 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_ADD_515_U5;
  assign new_P1_ADD_515_U133 = ~P1_INSTADDRPOINTER_REG_2_ | ~new_P1_ADD_515_U4;
  assign new_P1_ADD_515_U132 = ~new_P1_ADD_515_U108 | ~new_P1_ADD_515_U35;
  assign new_P1_ADD_515_U131 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_ADD_515_U34;
  assign new_P1_ADD_515_U130 = ~new_P1_ADD_515_U115 | ~new_P1_ADD_515_U49;
  assign new_P1_ADD_515_U129 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_ADD_515_U48;
  assign new_P1_ADD_515_U128 = ~new_P1_ADD_515_U120 | ~new_P1_ADD_515_U59;
  assign new_P1_ADD_515_U127 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_ADD_515_U58;
  assign new_P1_ADD_515_U126 = ~new_P1_ADD_515_U121 | ~new_P1_ADD_515_U60;
  assign new_P1_ADD_515_U125 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_ADD_515_U61;
  assign new_P1_ADD_515_U124 = ~new_P1_ADD_515_U97 | ~new_P1_ADD_515_U12;
  assign new_P1_ADD_515_U123 = ~P1_INSTADDRPOINTER_REG_6_ | ~new_P1_ADD_515_U13;
  assign new_P1_ADD_515_U122 = ~new_P1_ADD_515_U93;
  assign new_P1_ADD_515_U121 = ~new_P1_ADD_515_U61;
  assign new_P1_ADD_515_U120 = ~new_P1_ADD_515_U58;
  assign new_P1_ADD_515_U119 = ~new_P1_ADD_515_U56;
  assign new_P1_ADD_515_U118 = ~new_P1_ADD_515_U54;
  assign new_P1_ADD_515_U117 = ~new_P1_ADD_515_U52;
  assign new_P1_ADD_515_U116 = ~new_P1_ADD_515_U50;
  assign new_P1_ADD_515_U115 = ~new_P1_ADD_515_U48;
  assign new_P1_ADD_515_U114 = ~new_P1_ADD_515_U46;
  assign new_P1_ADD_515_U113 = ~new_P1_ADD_515_U44;
  assign new_P1_ADD_515_U112 = ~new_P1_ADD_515_U42;
  assign new_P1_ADD_515_U111 = ~new_P1_ADD_515_U40;
  assign new_P1_ADD_515_U110 = ~new_P1_ADD_515_U38;
  assign new_P1_ADD_515_U109 = ~new_P1_ADD_515_U36;
  assign new_P1_ADD_515_U108 = ~new_P1_ADD_515_U34;
  assign new_P1_ADD_515_U107 = ~new_P1_ADD_515_U32;
  assign new_P1_ADD_515_U106 = ~new_P1_ADD_515_U30;
  assign new_P1_ADD_515_U105 = ~new_P1_ADD_515_U28;
  assign new_P1_ADD_515_U104 = ~new_P1_ADD_515_U26;
  assign new_P1_ADD_515_U103 = ~new_P1_ADD_515_U24;
  assign new_P1_ADD_515_U102 = ~new_P1_ADD_515_U22;
  assign new_P1_ADD_515_U101 = ~new_P1_ADD_515_U20;
  assign new_P1_ADD_515_U100 = ~new_P1_ADD_515_U18;
  assign new_P1_ADD_515_U99 = ~new_P1_ADD_515_U16;
  assign new_P1_ADD_515_U98 = ~new_P1_ADD_515_U14;
  assign new_P1_ADD_515_U97 = ~new_P1_ADD_515_U13;
  assign new_P1_ADD_515_U96 = ~new_P1_ADD_515_U10;
  assign new_P1_ADD_515_U95 = ~new_P1_ADD_515_U8;
  assign new_P1_ADD_515_U94 = ~new_P1_ADD_515_U6;
  assign new_P1_ADD_515_U93 = ~new_P1_ADD_515_U121 | ~P1_INSTADDRPOINTER_REG_30_;
  assign new_P1_ADD_515_U92 = ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_ADD_515_U91 = ~new_P1_ADD_515_U182 | ~new_P1_ADD_515_U181;
  assign new_P1_ADD_515_U90 = ~new_P1_ADD_515_U180 | ~new_P1_ADD_515_U179;
  assign new_P1_ADD_515_U89 = ~new_P1_ADD_515_U178 | ~new_P1_ADD_515_U177;
  assign new_P1_ADD_515_U88 = ~new_P1_ADD_515_U176 | ~new_P1_ADD_515_U175;
  assign new_P1_ADD_515_U87 = ~new_P1_ADD_515_U174 | ~new_P1_ADD_515_U173;
  assign new_P1_ADD_515_U86 = ~new_P1_ADD_515_U172 | ~new_P1_ADD_515_U171;
  assign new_P1_ADD_515_U85 = ~new_P1_ADD_515_U170 | ~new_P1_ADD_515_U169;
  assign new_P1_ADD_515_U84 = ~new_P1_ADD_515_U168 | ~new_P1_ADD_515_U167;
  assign new_P1_ADD_515_U83 = ~new_P1_ADD_515_U166 | ~new_P1_ADD_515_U165;
  assign new_P1_ADD_515_U82 = ~new_P1_ADD_515_U164 | ~new_P1_ADD_515_U163;
  assign new_P1_ADD_515_U81 = ~new_P1_ADD_515_U162 | ~new_P1_ADD_515_U161;
  assign new_P1_ADD_515_U80 = ~new_P1_ADD_515_U160 | ~new_P1_ADD_515_U159;
  assign new_P1_ADD_515_U79 = ~new_P1_ADD_515_U158 | ~new_P1_ADD_515_U157;
  assign new_P1_ADD_515_U78 = ~new_P1_ADD_515_U156 | ~new_P1_ADD_515_U155;
  assign new_P1_ADD_515_U77 = ~new_P1_ADD_515_U154 | ~new_P1_ADD_515_U153;
  assign new_P1_ADD_515_U76 = ~new_P1_ADD_515_U152 | ~new_P1_ADD_515_U151;
  assign new_P1_ADD_515_U75 = ~new_P1_ADD_515_U150 | ~new_P1_ADD_515_U149;
  assign new_P1_ADD_515_U74 = ~new_P1_ADD_515_U148 | ~new_P1_ADD_515_U147;
  assign new_P1_ADD_515_U73 = ~new_P1_ADD_515_U146 | ~new_P1_ADD_515_U145;
  assign new_P1_ADD_515_U72 = ~new_P1_ADD_515_U144 | ~new_P1_ADD_515_U143;
  assign new_P1_ADD_515_U71 = ~new_P1_ADD_515_U142 | ~new_P1_ADD_515_U141;
  assign new_P1_ADD_515_U70 = ~new_P1_ADD_515_U140 | ~new_P1_ADD_515_U139;
  assign new_P1_ADD_515_U69 = ~new_P1_ADD_515_U138 | ~new_P1_ADD_515_U137;
  assign new_P1_ADD_515_U68 = ~new_P1_ADD_515_U136 | ~new_P1_ADD_515_U135;
  assign new_P1_ADD_515_U67 = ~new_P1_ADD_515_U134 | ~new_P1_ADD_515_U133;
  assign new_P1_ADD_515_U66 = ~new_P1_ADD_515_U132 | ~new_P1_ADD_515_U131;
  assign new_P1_ADD_515_U65 = ~new_P1_ADD_515_U130 | ~new_P1_ADD_515_U129;
  assign new_P1_ADD_515_U64 = ~new_P1_ADD_515_U128 | ~new_P1_ADD_515_U127;
  assign new_P1_ADD_515_U63 = ~new_P1_ADD_515_U126 | ~new_P1_ADD_515_U125;
  assign new_P1_ADD_515_U62 = ~new_P1_ADD_515_U124 | ~new_P1_ADD_515_U123;
  assign new_P1_ADD_515_U61 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_ADD_515_U120;
  assign new_P1_ADD_515_U60 = ~P1_INSTADDRPOINTER_REG_30_;
  assign new_P1_ADD_515_U59 = ~P1_INSTADDRPOINTER_REG_29_;
  assign new_P1_ADD_515_U58 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_ADD_515_U119;
  assign new_P1_ADD_515_U57 = ~P1_INSTADDRPOINTER_REG_28_;
  assign new_P1_ADD_515_U56 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_ADD_515_U118;
  assign new_P1_ADD_515_U55 = ~P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_ADD_515_U54 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_ADD_515_U117;
  assign new_P1_ADD_515_U53 = ~P1_INSTADDRPOINTER_REG_26_;
  assign new_P1_ADD_515_U52 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_ADD_515_U116;
  assign new_P1_ADD_515_U51 = ~P1_INSTADDRPOINTER_REG_25_;
  assign new_P1_ADD_515_U50 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_ADD_515_U115;
  assign new_P1_ADD_515_U49 = ~P1_INSTADDRPOINTER_REG_24_;
  assign new_P1_ADD_515_U48 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_ADD_515_U114;
  assign new_P1_ADD_515_U47 = ~P1_INSTADDRPOINTER_REG_23_;
  assign new_P1_ADD_515_U46 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_ADD_515_U113;
  assign new_P1_ADD_515_U45 = ~P1_INSTADDRPOINTER_REG_22_;
  assign new_P1_ADD_515_U44 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_ADD_515_U112;
  assign new_P1_ADD_515_U43 = ~P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_ADD_515_U42 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_ADD_515_U111;
  assign new_P1_ADD_515_U41 = ~P1_INSTADDRPOINTER_REG_20_;
  assign new_P1_ADD_515_U40 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_ADD_515_U110;
  assign new_P1_ADD_515_U39 = ~P1_INSTADDRPOINTER_REG_19_;
  assign new_P1_ADD_515_U38 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_ADD_515_U109;
  assign new_P1_ADD_515_U37 = ~P1_INSTADDRPOINTER_REG_18_;
  assign new_P1_ADD_515_U36 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_ADD_515_U108;
  assign new_P1_ADD_515_U35 = ~P1_INSTADDRPOINTER_REG_17_;
  assign new_P1_ADD_515_U34 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_ADD_515_U107;
  assign new_P1_ADD_515_U33 = ~P1_INSTADDRPOINTER_REG_16_;
  assign new_P1_ADD_515_U32 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_ADD_515_U106;
  assign new_P1_ADD_515_U31 = ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_ADD_515_U30 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_ADD_515_U105;
  assign new_P1_ADD_515_U29 = ~P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_ADD_515_U28 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_ADD_515_U104;
  assign new_P1_ADD_515_U27 = ~P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_ADD_515_U26 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_ADD_515_U103;
  assign new_P1_ADD_515_U25 = ~P1_INSTADDRPOINTER_REG_12_;
  assign new_P1_ADD_515_U24 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_ADD_515_U102;
  assign new_P1_ADD_515_U23 = ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_ADD_515_U22 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_ADD_515_U101;
  assign new_P1_ADD_515_U21 = ~P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_ADD_515_U20 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_ADD_515_U100;
  assign new_P1_ADD_515_U19 = ~P1_INSTADDRPOINTER_REG_9_;
  assign new_P1_ADD_515_U18 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_ADD_515_U99;
  assign new_P1_ADD_515_U17 = ~P1_INSTADDRPOINTER_REG_8_;
  assign new_P1_ADD_515_U16 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_ADD_515_U98;
  assign new_P1_ADD_515_U15 = ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_ADD_515_U14 = ~new_P1_ADD_515_U97 | ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_ADD_515_U13 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_ADD_515_U96;
  assign new_P1_ADD_515_U12 = ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_ADD_515_U11 = ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_ADD_515_U10 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_ADD_515_U95;
  assign new_P1_ADD_515_U9 = ~P1_INSTADDRPOINTER_REG_4_;
  assign new_P1_ADD_515_U8 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_ADD_515_U94;
  assign new_P1_ADD_515_U7 = ~P1_INSTADDRPOINTER_REG_3_;
  assign new_P1_ADD_515_U6 = ~P1_INSTADDRPOINTER_REG_2_ | ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_ADD_515_U5 = ~P1_INSTADDRPOINTER_REG_2_;
  assign new_P1_ADD_515_U4 = ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_GTE_485_U7 = ~new_P1_R2238_U21 & ~new_P1_R2238_U22 & ~new_P1_R2238_U19 & ~new_P1_R2238_U20;
  assign new_P1_GTE_485_U6 = ~new_P1_R2238_U6 & ~new_P1_GTE_485_U7;
  assign new_P1_ADD_405_U186 = ~new_P1_ADD_405_U110 | ~new_P1_ADD_405_U33;
  assign new_P1_ADD_405_U185 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_ADD_405_U32;
  assign new_P1_ADD_405_U184 = ~new_P1_ADD_405_U119 | ~new_P1_ADD_405_U51;
  assign new_P1_ADD_405_U183 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_ADD_405_U50;
  assign new_P1_ADD_405_U182 = ~new_P1_ADD_405_U101 | ~new_P1_ADD_405_U15;
  assign new_P1_ADD_405_U181 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_ADD_405_U14;
  assign new_P1_ADD_405_U180 = ~new_P1_ADD_405_U106 | ~new_P1_ADD_405_U25;
  assign new_P1_ADD_405_U179 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_ADD_405_U24;
  assign new_P1_ADD_405_U178 = ~new_P1_ADD_405_U115 | ~new_P1_ADD_405_U43;
  assign new_P1_ADD_405_U177 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_ADD_405_U42;
  assign new_P1_ADD_405_U176 = ~new_P1_ADD_405_U122 | ~new_P1_ADD_405_U57;
  assign new_P1_ADD_405_U175 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_ADD_405_U56;
  assign new_P1_ADD_405_U174 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_ADD_405_U6;
  assign new_P1_ADD_405_U173 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_ADD_405_U4;
  assign new_P2_U2352 = new_P2_U7873 & new_P2_U2617 & new_P2_U3300;
  assign new_P2_U2353 = new_P2_U4343 & new_P2_U2439;
  assign new_P2_U2354 = P2_STATE2_REG_0_ & new_P2_U7861 & new_P2_U7873;
  assign new_P2_U2355 = new_P2_U2447 & new_P2_U7861;
  assign new_P2_U2356 = P2_STATE2_REG_0_ & new_P2_U3253;
  assign new_P2_U2357 = new_P2_U3712 & new_P2_U2458;
  assign new_P2_U2358 = new_P2_U4431 & P2_STATE2_REG_0_;
  assign new_P2_U2359 = new_P2_U4411 & new_P2_U3265;
  assign new_P2_U2360 = ~new_U211 & ~P2_STATEBS16_REG;
  assign new_P2_U2361 = new_P2_R2238_U6 & new_P2_U2356;
  assign new_P2_U2362 = new_P2_U2398 & new_P2_U4443;
  assign new_P2_U2363 = P2_STATE2_REG_2_ & new_P2_U3535;
  assign new_P2_U2364 = P2_STATE2_REG_2_ & new_P2_U3546;
  assign new_P2_U2365 = new_P2_U4443 & P2_STATE2_REG_3_;
  assign new_P2_U2366 = P2_STATE2_REG_1_ & new_P2_U3546;
  assign new_P2_U2367 = new_P2_U2364 & new_P2_U4417;
  assign new_P2_U2368 = new_P2_U2363 & new_P2_U4420;
  assign new_P2_U2369 = new_P2_U2364 & new_P2_U4428;
  assign new_P2_U2370 = new_P2_U2447 & new_P2_U3537;
  assign new_P2_U2371 = new_P2_U3990 & new_P2_U3537;
  assign new_P2_U2372 = new_P2_U3989 & new_P2_U3537;
  assign new_P2_U2373 = new_P2_U4419 & new_P2_U3537;
  assign new_P2_U2374 = new_P2_U4468 & P2_STATE2_REG_0_;
  assign new_P2_U2375 = new_P2_U4441 & new_P2_U3521;
  assign new_P2_U2376 = new_P2_U3873 & new_P2_U2436;
  assign new_P2_U2377 = new_P2_U2367 & new_P2_U4411;
  assign new_P2_U2378 = P2_STATE2_REG_3_ & new_P2_U3546;
  assign new_P2_U2379 = new_P2_U4440 & new_P2_U7865;
  assign new_P2_U2380 = new_P2_U4441 & new_P2_U7865;
  assign new_P2_U2381 = new_P2_U3535 & new_P2_U3270;
  assign new_P2_U2382 = new_P2_U2366 & new_P2_U3647;
  assign new_P2_U2383 = new_P2_U2366 & new_P2_U3528;
  assign new_P2_U2384 = new_P2_U2368 & new_P2_U4417;
  assign new_P2_U2385 = new_P2_U2368 & new_P2_U4428;
  assign new_P2_U2386 = new_P2_U2363 & new_P2_U4436;
  assign new_P2_U2387 = new_P2_U5940 & new_P2_U3537;
  assign new_P2_U2388 = new_P2_U2363 & new_P2_U5675;
  assign new_P2_U2389 = new_P2_U2363 & new_P2_U5677;
  assign new_P2_U2390 = new_P2_U2363 & new_P2_U5679;
  assign new_P2_U2391 = new_P2_U2369 & new_P2_U3545;
  assign new_P2_U2392 = new_P2_U6571 & new_P2_U2369;
  assign new_P2_U2393 = new_P2_U4440 & new_P2_U3521;
  assign new_P2_U2394 = new_P2_U4442 & new_P2_U2616;
  assign new_P2_U2395 = new_P2_U4442 & new_P2_U7873;
  assign new_P2_U2396 = new_P2_U3541 & new_P2_U3284;
  assign new_P2_U2397 = new_P2_U4441 & new_P2_U4601;
  assign new_P2_U2398 = new_P2_U4430 & P2_STATEBS16_REG;
  assign new_P2_U2399 = new_U314 & new_P2_U4443;
  assign new_P2_U2400 = new_U303 & new_P2_U4443;
  assign new_P2_U2401 = new_U292 & new_P2_U4443;
  assign new_P2_U2402 = new_U289 & new_P2_U4443;
  assign new_P2_U2403 = new_U288 & new_P2_U4443;
  assign new_P2_U2404 = new_U287 & new_P2_U4443;
  assign new_P2_U2405 = new_U286 & new_P2_U4443;
  assign new_P2_U2406 = new_U285 & new_P2_U4443;
  assign new_P2_U2407 = new_U298 & new_P2_U2362;
  assign new_P2_U2408 = new_U307 & new_P2_U2362;
  assign new_P2_U2409 = new_U297 & new_P2_U2362;
  assign new_P2_U2410 = new_U306 & new_P2_U2362;
  assign new_P2_U2411 = new_U296 & new_P2_U2362;
  assign new_P2_U2412 = new_U305 & new_P2_U2362;
  assign new_P2_U2413 = new_U295 & new_P2_U2362;
  assign new_P2_U2414 = new_U304 & new_P2_U2362;
  assign new_P2_U2415 = new_U294 & new_P2_U2362;
  assign new_P2_U2416 = new_U302 & new_P2_U2362;
  assign new_P2_U2417 = new_U293 & new_P2_U2362;
  assign new_P2_U2418 = new_U301 & new_P2_U2362;
  assign new_P2_U2419 = new_U291 & new_P2_U2362;
  assign new_P2_U2420 = new_U300 & new_P2_U2362;
  assign new_P2_U2421 = new_U290 & new_P2_U2362;
  assign new_P2_U2422 = new_U299 & new_P2_U2362;
  assign new_P2_U2423 = new_P2_U2365 & new_P2_U3255;
  assign new_P2_U2424 = new_P2_U2365 & new_P2_U3278;
  assign new_P2_U2425 = new_P2_U2365 & new_P2_U3521;
  assign new_P2_U2426 = new_P2_U2365 & new_P2_U3279;
  assign new_P2_U2427 = new_P2_U2375 & new_P2_U3279;
  assign new_P2_U2428 = new_P2_U2365 & new_P2_U2616;
  assign new_P2_U2429 = new_P2_U2365 & new_P2_U2617;
  assign new_P2_U2430 = P2_STATE2_REG_0_ & new_P2_U3541;
  assign new_P2_U2431 = new_P2_U2365 & new_P2_U3253;
  assign new_P2_U2432 = new_P2_U2365 & new_P2_U3280;
  assign new_P2_U2433 = new_P2_U2375 & new_P2_U3295;
  assign new_P2_U2434 = new_P2_U2375 & new_P2_U7869;
  assign new_P2_U2435 = new_P2_U2356 & new_P2_U3541;
  assign new_P2_U2436 = new_P2_U7859 & new_P2_U7867;
  assign new_P2_U2437 = new_P2_U2364 & new_P2_U7871;
  assign new_P2_U2438 = new_P2_U7859 & new_P2_U3278;
  assign new_P2_U2439 = new_P2_U4339 & new_P2_U3521;
  assign new_P2_U2440 = new_P2_U3580 & new_P2_U3428;
  assign new_P2_U2441 = new_P2_U4647 & new_P2_U3580;
  assign new_P2_U2442 = new_P2_U8067 & new_P2_U3428;
  assign new_P2_U2443 = new_P2_U4647 & new_P2_U8067;
  assign new_P2_U2444 = new_P2_U3243 & new_P2_U3307;
  assign new_P2_U2445 = new_P2_U4650 & new_P2_U3307;
  assign new_P2_U2446 = new_P2_R2088_U6 & new_P2_U4424;
  assign new_P2_U2447 = P2_STATE2_REG_0_ & new_P2_U2616;
  assign new_P2_U2448 = P2_STATE2_REG_2_ & P2_STATE2_REG_1_;
  assign new_P2_U2449 = new_P2_U3278 & new_P2_U3521;
  assign new_P2_U2450 = new_P2_U2354 & new_P2_U7871;
  assign new_P2_U2451 = new_P2_U2438 & new_P2_U4601 & new_P2_U2457;
  assign new_P2_U2452 = P2_INSTQUEUERD_ADDR_REG_2_ & P2_INSTQUEUERD_ADDR_REG_1_ & new_P2_U3272;
  assign new_P2_U2453 = P2_INSTQUEUERD_ADDR_REG_2_ & P2_INSTQUEUERD_ADDR_REG_0_ & new_P2_U3271;
  assign new_P2_U2454 = P2_INSTQUEUERD_ADDR_REG_2_ & new_P2_U3271 & new_P2_U3272;
  assign new_P2_U2455 = P2_INSTQUEUERD_ADDR_REG_1_ & new_P2_U3276 & new_P2_U3272;
  assign new_P2_U2456 = P2_INSTQUEUERD_ADDR_REG_0_ & new_P2_U3276 & new_P2_U3271;
  assign new_P2_U2457 = new_P2_U3521 & new_P2_U3255;
  assign new_P2_U2458 = new_P2_U7863 & new_P2_U2617 & new_P2_U3279;
  assign new_P2_U2459 = new_P2_U4393 & new_P2_U8053 & new_P2_U8052;
  assign new_P2_U2460 = new_P2_R2182_U40 & new_P2_U3317;
  assign new_P2_U2461 = new_P2_U3579 & new_P2_U3426;
  assign new_P2_U2462 = new_P2_R2182_U76 & new_P2_R2182_U40;
  assign new_P2_U2463 = new_P2_U4637 & new_P2_U2462;
  assign new_P2_U2464 = P2_INSTQUEUEWR_ADDR_REG_2_ & P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_U2465 = P2_INSTQUEUEWR_ADDR_REG_2_ & new_P2_U3309;
  assign new_P2_U2466 = new_P2_R2099_U96 & new_P2_R2099_U95;
  assign new_P2_U2467 = new_P2_R2099_U5 & new_P2_R2099_U94;
  assign new_P2_U2468 = new_P2_U3320 & new_P2_U4657;
  assign new_P2_U2469 = new_P2_U4633 & new_P2_U2462;
  assign new_P2_U2470 = new_P2_R2099_U5 & new_P2_U3323;
  assign new_P2_U2471 = new_P2_U3339 & new_P2_U4715;
  assign new_P2_U2472 = new_P2_U4634 & new_P2_U2462;
  assign new_P2_U2473 = new_P2_R2099_U94 & new_P2_U3324;
  assign new_P2_U2474 = new_P2_U3354 & new_P2_U4774;
  assign new_P2_U2475 = new_P2_U4635 & new_P2_R2182_U69;
  assign new_P2_U2476 = ~new_P2_R2182_U69 & ~new_P2_R2182_U68;
  assign new_P2_U2477 = new_P2_U2476 & new_P2_U2462;
  assign new_P2_U2478 = ~P2_INSTQUEUEWR_ADDR_REG_0_ & ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_U2479 = ~new_P2_R2099_U94 & ~new_P2_R2099_U5;
  assign new_P2_U2480 = new_P2_U3366 & new_P2_U4831;
  assign new_P2_U2481 = new_P2_U8064 & new_P2_U3426;
  assign new_P2_U2482 = new_P2_U4638 & new_P2_U4637;
  assign new_P2_U2483 = new_P2_R2099_U95 & new_P2_U3322;
  assign new_P2_U2484 = new_P2_U3379 & new_P2_U4889;
  assign new_P2_U2485 = new_P2_U4638 & new_P2_U4633;
  assign new_P2_U2486 = new_P2_U3391 & new_P2_U4946;
  assign new_P2_U2487 = new_P2_U4638 & new_P2_U4634;
  assign new_P2_U2488 = new_P2_U3402 & new_P2_U5004;
  assign new_P2_U2489 = new_P2_U4638 & new_P2_U2476;
  assign new_P2_U2490 = new_P2_U3414 & new_P2_U5061;
  assign new_P2_U2491 = new_P2_U4640 & new_P2_U3579;
  assign new_P2_U2492 = new_P2_R2099_U96 & new_P2_U3321;
  assign new_P2_U2493 = new_P2_U3427 & new_P2_U3425;
  assign new_P2_U2494 = new_P2_U4633 & new_P2_U2460;
  assign new_P2_U2495 = new_P2_U3440 & new_P2_U5174;
  assign new_P2_U2496 = new_P2_U4634 & new_P2_U2460;
  assign new_P2_U2497 = new_P2_U3451 & new_P2_U5232;
  assign new_P2_U2498 = new_P2_U2476 & new_P2_U2460;
  assign new_P2_U2499 = new_P2_U3463 & new_P2_U5289;
  assign new_P2_U2500 = new_P2_U4640 & new_P2_U8064;
  assign new_P2_U2501 = ~new_P2_R2182_U40 & ~new_P2_R2182_U76;
  assign new_P2_U2502 = new_P2_U2501 & new_P2_U4637;
  assign new_P2_U2503 = ~P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P2_U2504 = ~new_P2_R2099_U95 & ~new_P2_R2099_U96;
  assign new_P2_U2505 = new_P2_U3474 & new_P2_U5347;
  assign new_P2_U2506 = new_P2_U2501 & new_P2_U4633;
  assign new_P2_U2507 = new_P2_U3486 & new_P2_U5404;
  assign new_P2_U2508 = new_P2_U2501 & new_P2_U4634;
  assign new_P2_U2509 = new_P2_U3497 & new_P2_U5462;
  assign new_P2_U2510 = new_P2_U2501 & new_P2_U2476;
  assign new_P2_U2511 = new_P2_U3509 & new_P2_U5519;
  assign new_P2_U2512 = new_P2_U3869 & new_P2_U8069 & new_P2_U8068;
  assign new_P2_U2513 = new_P2_U5580 & new_P2_U5579;
  assign new_P2_U2514 = new_P2_U3882 & new_P2_U3881 & new_P2_U7896;
  assign new_P2_U2515 = new_P2_U8082 & new_P2_U8100;
  assign new_P2_U2516 = new_P2_U5616 & P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_U2517 = new_P2_U2515 & new_P2_U2516;
  assign new_P2_U2518 = new_P2_U5616 & new_P2_U3272;
  assign new_P2_U2519 = new_P2_U2515 & new_P2_U2518;
  assign new_P2_U2520 = new_P2_U8082 & new_P2_U3582;
  assign new_P2_U2521 = new_P2_U2520 & new_P2_U2516;
  assign new_P2_U2522 = new_P2_U2520 & new_P2_U2518;
  assign new_P2_U2523 = P2_INSTQUEUERD_ADDR_REG_0_ & new_P2_U3530;
  assign new_P2_U2524 = new_P2_U2515 & new_P2_U2523;
  assign new_P2_U2525 = new_P2_U3272 & new_P2_U3530;
  assign new_P2_U2526 = new_P2_U2515 & new_P2_U2525;
  assign new_P2_U2527 = new_P2_U2520 & new_P2_U2523;
  assign new_P2_U2528 = new_P2_U2520 & new_P2_U2525;
  assign new_P2_U2529 = new_P2_U3582 & new_P2_U3581;
  assign new_P2_U2530 = new_P2_U2525 & new_P2_U2529;
  assign new_P2_U2531 = new_P2_U2523 & new_P2_U2529;
  assign new_P2_U2532 = new_P2_U8100 & new_P2_U3581;
  assign new_P2_U2533 = new_P2_U2525 & new_P2_U2532;
  assign new_P2_U2534 = new_P2_U2523 & new_P2_U2532;
  assign new_P2_U2535 = new_P2_U2529 & new_P2_U2518;
  assign new_P2_U2536 = new_P2_U2529 & new_P2_U2516;
  assign new_P2_U2537 = new_P2_U2518 & new_P2_U2532;
  assign new_P2_U2538 = new_P2_U2516 & new_P2_U2532;
  assign new_P2_U2539 = ~new_P2_R2147_U8 & ~new_P2_R2147_U4;
  assign new_P2_U2540 = ~P2_INSTQUEUERD_ADDR_REG_0_ & ~new_P2_R2147_U9;
  assign new_P2_U2541 = new_P2_U2539 & new_P2_U2540;
  assign new_P2_U2542 = P2_INSTQUEUERD_ADDR_REG_0_ & new_P2_U3529;
  assign new_P2_U2543 = new_P2_U2539 & new_P2_U2542;
  assign new_P2_U2544 = new_P2_R2147_U4 & new_P2_U3526;
  assign new_P2_U2545 = new_P2_U2544 & new_P2_U2540;
  assign new_P2_U2546 = new_P2_U2544 & new_P2_U2542;
  assign new_P2_U2547 = new_P2_R2147_U9 & new_P2_U3532;
  assign new_P2_U2548 = new_P2_U2539 & new_P2_U2547;
  assign new_P2_U2549 = P2_INSTQUEUERD_ADDR_REG_0_ & new_P2_R2147_U9;
  assign new_P2_U2550 = new_P2_U2539 & new_P2_U2549;
  assign new_P2_U2551 = new_P2_U2544 & new_P2_U2547;
  assign new_P2_U2552 = new_P2_U2544 & new_P2_U2549;
  assign new_P2_U2553 = new_P2_R2147_U8 & new_P2_U3531;
  assign new_P2_U2554 = new_P2_U2540 & new_P2_U2553;
  assign new_P2_U2555 = new_P2_U2542 & new_P2_U2553;
  assign new_P2_U2556 = new_P2_R2147_U4 & new_P2_R2147_U8;
  assign new_P2_U2557 = new_P2_U2540 & new_P2_U2556;
  assign new_P2_U2558 = new_P2_U2542 & new_P2_U2556;
  assign new_P2_U2559 = new_P2_U2553 & new_P2_U2547;
  assign new_P2_U2560 = new_P2_U2553 & new_P2_U2549;
  assign new_P2_U2561 = new_P2_U2547 & new_P2_U2556;
  assign new_P2_U2562 = new_P2_U2549 & new_P2_U2556;
  assign new_P2_U2563 = new_P2_U8100 & new_P2_U3272;
  assign new_P2_U2564 = new_P2_U4409 & new_P2_U3583;
  assign new_P2_U2565 = new_P2_U2564 & new_P2_U2563;
  assign new_P2_U2566 = new_P2_U8100 & P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_U2567 = new_P2_U2564 & new_P2_U2566;
  assign new_P2_U2568 = new_P2_U3582 & new_P2_U3272;
  assign new_P2_U2569 = new_P2_U2564 & new_P2_U2568;
  assign new_P2_U2570 = P2_INSTQUEUERD_ADDR_REG_0_ & new_P2_U3582;
  assign new_P2_U2571 = new_P2_U2564 & new_P2_U2570;
  assign new_P2_U2572 = new_P2_U3583 & new_P2_U3553;
  assign new_P2_U2573 = new_P2_U2572 & new_P2_U2563;
  assign new_P2_U2574 = new_P2_U2572 & new_P2_U2566;
  assign new_P2_U2575 = new_P2_U2572 & new_P2_U2568;
  assign new_P2_U2576 = new_P2_U2572 & new_P2_U2570;
  assign new_P2_U2577 = new_P2_U4409 & new_P2_U8149;
  assign new_P2_U2578 = new_P2_U2577 & new_P2_U2563;
  assign new_P2_U2579 = new_P2_U2577 & new_P2_U2566;
  assign new_P2_U2580 = new_P2_U2577 & new_P2_U2568;
  assign new_P2_U2581 = new_P2_U2577 & new_P2_U2570;
  assign new_P2_U2582 = new_P2_U8149 & new_P2_U3553;
  assign new_P2_U2583 = new_P2_U2563 & new_P2_U2582;
  assign new_P2_U2584 = new_P2_U2566 & new_P2_U2582;
  assign new_P2_U2585 = new_P2_U2568 & new_P2_U2582;
  assign new_P2_U2586 = new_P2_U2570 & new_P2_U2582;
  assign new_P2_U2587 = P2_EBX_REG_31_ & new_P2_U2391;
  assign new_P2_U2588 = new_P2_U2377 & new_P2_U2360;
  assign new_P2_U2589 = new_P2_U3549 & new_P2_U4457 & new_P2_U7581 & new_P2_U3550;
  assign new_P2_U2590 = new_P2_U5590 & new_P2_U2436;
  assign new_P2_U2591 = ~new_P2_U4274 | ~new_P2_U4273;
  assign new_P2_U2592 = ~new_P2_U4272 | ~new_P2_U4271;
  assign new_P2_U2593 = ~new_P2_U4270 | ~new_P2_U4269;
  assign new_P2_U2594 = ~new_P2_U4268 | ~new_P2_U4267;
  assign new_P2_U2595 = ~new_P2_U4266 | ~new_P2_U4265;
  assign new_P2_U2596 = ~new_P2_U4264 | ~new_P2_U4263;
  assign new_P2_U2597 = ~new_P2_U4262 | ~new_P2_U4261;
  assign new_P2_U2598 = ~new_P2_U4260 | ~new_P2_U4259;
  assign new_P2_U2599 = ~new_P2_U4255 | ~new_P2_U4256 | ~new_P2_U4258 | ~new_P2_U4257;
  assign new_P2_U2600 = ~new_P2_U4251 | ~new_P2_U4252 | ~new_P2_U4254 | ~new_P2_U4253;
  assign new_P2_U2601 = ~new_P2_U4247 | ~new_P2_U4248 | ~new_P2_U4250 | ~new_P2_U4249;
  assign new_P2_U2602 = ~new_P2_U4243 | ~new_P2_U4244 | ~new_P2_U4246 | ~new_P2_U4245;
  assign new_P2_U2603 = ~new_P2_U4239 | ~new_P2_U4240 | ~new_P2_U4242 | ~new_P2_U4241;
  assign new_P2_U2604 = ~new_P2_U4235 | ~new_P2_U4236 | ~new_P2_U4238 | ~new_P2_U4237;
  assign new_P2_U2605 = ~new_P2_U4231 | ~new_P2_U4232 | ~new_P2_U4234 | ~new_P2_U4233;
  assign new_P2_U2606 = ~new_P2_U4227 | ~new_P2_U4228 | ~new_P2_U4230 | ~new_P2_U4229;
  assign new_P2_U2607 = ~new_P2_U4223 | ~new_P2_U4224 | ~new_P2_U4226 | ~new_P2_U4225;
  assign new_P2_U2608 = ~new_P2_U4219 | ~new_P2_U4220 | ~new_P2_U4222 | ~new_P2_U4221;
  assign new_P2_U2609 = ~new_P2_U4215 | ~new_P2_U4216 | ~new_P2_U4218 | ~new_P2_U4217;
  assign new_P2_U2610 = ~new_P2_U4211 | ~new_P2_U4212 | ~new_P2_U4214 | ~new_P2_U4213;
  assign new_P2_U2611 = ~new_P2_U4207 | ~new_P2_U4208 | ~new_P2_U4210 | ~new_P2_U4209;
  assign new_P2_U2612 = ~new_P2_U4203 | ~new_P2_U4204 | ~new_P2_U4206 | ~new_P2_U4205;
  assign new_P2_U2613 = ~new_P2_U4199 | ~new_P2_U4200 | ~new_P2_U4202 | ~new_P2_U4201;
  assign new_P2_U2614 = ~new_P2_U4195 | ~new_P2_U4196 | ~new_P2_U4198 | ~new_P2_U4197;
  assign new_P2_U2615 = P2_INSTQUEUERD_ADDR_REG_4_ & new_P2_U3519;
  assign new_P2_U2616 = ~new_P2_U3706 | ~new_P2_U3705;
  assign new_P2_U2617 = ~new_P2_U3694 | ~new_P2_U3693;
  assign new_P2_U2618 = ~new_P2_U4350 | ~new_P2_U7453;
  assign new_P2_U2619 = ~new_P2_U4351 | ~new_P2_U7456;
  assign new_P2_U2620 = ~new_P2_U4353 | ~new_P2_U7462;
  assign new_P2_U2621 = ~new_P2_U4354 | ~new_P2_U7465;
  assign new_P2_U2622 = ~new_P2_U4355 | ~new_P2_U7468;
  assign new_P2_U2623 = ~new_P2_U4356 | ~new_P2_U7471;
  assign new_P2_U2624 = ~new_P2_U4357 | ~new_P2_U7474;
  assign new_P2_U2625 = ~new_P2_U4358 | ~new_P2_U7477;
  assign new_P2_U2626 = ~new_P2_U4359 | ~new_P2_U7480;
  assign new_P2_U2627 = ~new_P2_U4360 | ~new_P2_U7483;
  assign new_P2_U2628 = ~new_P2_U4361 | ~new_P2_U7486;
  assign new_P2_U2629 = ~new_P2_U4362 | ~new_P2_U7489;
  assign new_P2_U2630 = ~new_P2_U4364 | ~new_P2_U7495;
  assign new_P2_U2631 = ~new_P2_U4365 | ~new_P2_U7498;
  assign new_P2_U2632 = ~new_P2_U4366 | ~new_P2_U7501;
  assign new_P2_U2633 = ~new_P2_U4367 | ~new_P2_U7504;
  assign new_P2_U2634 = ~new_P2_U4368 | ~new_P2_U7508 | ~new_P2_U7507;
  assign new_P2_U2635 = ~new_P2_U4369 | ~new_P2_U7512 | ~new_P2_U7511;
  assign new_P2_U2636 = ~new_P2_U4370 | ~new_P2_U7516 | ~new_P2_U7515;
  assign new_P2_U2637 = ~new_P2_U4371 | ~new_P2_U7520 | ~new_P2_U7519;
  assign new_P2_U2638 = ~new_P2_U4372 | ~new_P2_U7524 | ~new_P2_U7523;
  assign new_P2_U2639 = ~new_P2_U4373 | ~new_P2_U7528 | ~new_P2_U7527;
  assign new_P2_U2640 = ~new_P2_U4344 | ~new_P2_U7434 | ~new_P2_U7433;
  assign new_P2_U2641 = ~new_P2_U4345 | ~new_P2_U7438 | ~new_P2_U7437;
  assign new_P2_U2642 = ~new_P2_U4346 | ~new_P2_U7441;
  assign new_P2_U2643 = ~new_P2_U4347 | ~new_P2_U7444;
  assign new_P2_U2644 = ~new_P2_U4348 | ~new_P2_U7447;
  assign new_P2_U2645 = ~new_P2_U4349 | ~new_P2_U7450;
  assign new_P2_U2646 = ~new_P2_U4352 | ~new_P2_U7459;
  assign new_P2_U2647 = ~new_P2_U4363 | ~new_P2_U7492;
  assign new_P2_U2648 = ~new_P2_U4374 | ~new_P2_U7531;
  assign new_P2_U2649 = ~new_P2_U4375 | ~new_P2_U7534 | ~new_P2_U3300;
  assign new_P2_U2650 = new_P2_U2352 & new_P2_U3242;
  assign new_P2_U2651 = new_P2_U2352 & new_P2_U7217;
  assign new_P2_U2652 = new_P2_U2352 & new_P2_U7251;
  assign new_P2_U2653 = new_P2_U2352 & new_P2_U7285;
  assign new_P2_U2654 = ~new_P2_U7423 | ~new_P2_U7422;
  assign new_P2_U2655 = ~new_P2_U4338 | ~new_P2_U7424;
  assign new_P2_U2656 = ~new_P2_U4340 | ~new_P2_U7427;
  assign new_P2_U2657 = ~new_P2_U4342 | ~new_P2_U7429;
  assign new_P2_U2658 = new_P2_U2354 & new_P2_U2598;
  assign new_P2_U2659 = new_P2_U2354 & new_P2_U2597;
  assign new_P2_U2660 = new_P2_U2354 & new_P2_U2596;
  assign new_P2_U2661 = new_P2_U2354 & new_P2_U2595;
  assign new_P2_U2662 = new_P2_U2354 & new_P2_U2594;
  assign new_P2_U2663 = new_P2_U2354 & new_P2_U2593;
  assign new_P2_U2664 = new_P2_U2354 & new_P2_U2592;
  assign new_P2_U2665 = new_P2_U2354 & new_P2_U2591;
  assign new_P2_U2666 = new_P2_U2614 & new_P2_U2355;
  assign new_P2_U2667 = new_P2_U2613 & new_P2_U2355;
  assign new_P2_U2668 = new_P2_U2612 & new_P2_U2355;
  assign new_P2_U2669 = new_P2_U2611 & new_P2_U2355;
  assign new_P2_U2670 = new_P2_U2610 & new_P2_U2355;
  assign new_P2_U2671 = new_P2_U2609 & new_P2_U2355;
  assign new_P2_U2672 = new_P2_U2608 & new_P2_U2355;
  assign new_P2_U2673 = new_P2_U2607 & new_P2_U2355;
  assign new_P2_U2674 = P2_INSTQUEUE_REG_0__7_ & new_P2_U2355;
  assign new_P2_U2675 = P2_INSTQUEUE_REG_0__6_ & new_P2_U2355;
  assign new_P2_U2676 = P2_INSTQUEUE_REG_0__5_ & new_P2_U2355;
  assign new_P2_U2677 = P2_INSTQUEUE_REG_0__4_ & new_P2_U2355;
  assign new_P2_U2678 = P2_INSTQUEUE_REG_0__3_ & new_P2_U2355;
  assign new_P2_U2679 = P2_INSTQUEUE_REG_0__2_ & new_P2_U2355;
  assign new_P2_U2680 = P2_INSTQUEUE_REG_0__1_ & new_P2_U2355;
  assign new_P2_U2681 = ~new_P2_U7166 | ~new_P2_U4275;
  assign new_P2_U2682 = new_P2_U2355 & new_P2_ADD_402_1132_U18;
  assign new_P2_U2683 = new_P2_ADD_402_1132_U19 & new_P2_U2355;
  assign new_P2_U2684 = new_P2_ADD_402_1132_U24 & new_P2_U2355;
  assign new_P2_U2685 = new_P2_ADD_402_1132_U22 & new_P2_U2355;
  assign new_P2_U2686 = new_P2_ADD_402_1132_U21 & new_P2_U2355;
  assign new_P2_U2687 = new_P2_ADD_402_1132_U25 & new_P2_U2355;
  assign new_P2_U2688 = new_P2_ADD_402_1132_U20 & new_P2_U2355;
  assign new_P2_U2689 = ~new_P2_U7142 | ~new_P2_U7141;
  assign new_P2_U2690 = ~new_P2_U7144 | ~new_P2_U7143;
  assign new_P2_U2691 = ~new_P2_U7146 | ~new_P2_U7145;
  assign new_P2_U2692 = ~new_P2_U7148 | ~new_P2_U7147;
  assign new_P2_U2693 = ~new_P2_U7153 | ~new_P2_U7152;
  assign new_P2_U2694 = ~new_P2_U7155 | ~new_P2_U7154;
  assign new_P2_U2695 = ~new_P2_U7157 | ~new_P2_U7156;
  assign new_P2_U2696 = ~new_P2_U7159 | ~new_P2_U7158;
  assign new_P1_ADD_405_U172 = ~new_P1_ADD_405_U97 | ~new_P1_ADD_405_U7;
  assign new_P2_U2698 = P2_INSTQUEUERD_ADDR_REG_4_ & new_P2_U3554;
  assign new_P2_U2699 = ~new_P2_U7138 | ~new_P2_U7139 | ~new_P2_U7140;
  assign new_P2_U2700 = ~new_P2_U7149 | ~new_P2_U7150 | ~new_P2_U7151;
  assign new_P2_U2701 = ~new_P2_U7160 | ~new_P2_U7161 | ~new_P2_U7162;
  assign new_P2_U2702 = ~new_P2_U7163 | ~new_P2_U7164 | ~new_P2_U7165;
  assign new_P2_U2703 = ~new_P2_U7727 | ~new_P2_U7726;
  assign new_P2_U2704 = ~new_P2_U7729 | ~new_P2_U7728;
  assign new_P2_U2705 = ~new_P2_U4390 | ~new_P2_U7730;
  assign new_P2_U2706 = ~new_P2_U3550 | ~new_P2_U7732 | ~new_P2_U7733;
  assign new_P2_U2707 = ~new_P2_U4391 | ~new_P2_U7734;
  assign new_P2_U2708 = new_P2_R2219_U25 & new_P2_U7723;
  assign new_P2_U2709 = new_P2_R2219_U26 & new_P2_U7723;
  assign new_P2_U2710 = new_P2_R2219_U27 & new_P2_U7723;
  assign new_P2_U2711 = ~P2_STATE2_REG_0_ | ~new_P2_U7724;
  assign new_P2_U2712 = ~new_P2_U4407 | ~new_P2_U7871 | ~P2_STATE2_REG_0_;
  assign new_P2_U2713 = ~P2_STATE2_REG_0_ | ~new_P2_U7725;
  assign new_P2_U2714 = ~new_P2_U4408 | ~new_P2_U7871 | ~P2_STATE2_REG_0_;
  assign new_P2_U2715 = ~new_P2_U2356 | ~new_P2_U2616;
  assign new_P2_U2716 = ~new_P2_U7617 | ~new_P2_U7618 | ~new_P2_U7620 | ~new_P2_U7619;
  assign new_P2_U2717 = ~new_P2_U7621 | ~new_P2_U7622 | ~new_P2_U7624 | ~new_P2_U7623;
  assign new_P2_U2718 = ~new_P2_U7629 | ~new_P2_U7630 | ~new_P2_U7632 | ~new_P2_U7631;
  assign new_P2_U2719 = ~new_P2_U7633 | ~new_P2_U7634 | ~new_P2_U7636 | ~new_P2_U7635;
  assign new_P2_U2720 = ~new_P2_U7637 | ~new_P2_U7638 | ~new_P2_U7640 | ~new_P2_U7639;
  assign new_P2_U2721 = ~new_P2_U7641 | ~new_P2_U7642 | ~new_P2_U7644 | ~new_P2_U7643;
  assign new_P2_U2722 = ~new_P2_U7645 | ~new_P2_U7646 | ~new_P2_U7648 | ~new_P2_U7647;
  assign new_P2_U2723 = ~new_P2_U7649 | ~new_P2_U7650 | ~new_P2_U7652 | ~new_P2_U7651;
  assign new_P2_U2724 = ~new_P2_U7653 | ~new_P2_U7654 | ~new_P2_U7656 | ~new_P2_U7655;
  assign new_P2_U2725 = ~new_P2_U7657 | ~new_P2_U7658 | ~new_P2_U7660 | ~new_P2_U7659;
  assign new_P2_U2726 = ~new_P2_U7661 | ~new_P2_U7662 | ~new_P2_U7664 | ~new_P2_U7663;
  assign new_P2_U2727 = ~new_P2_U7665 | ~new_P2_U7666 | ~new_P2_U7668 | ~new_P2_U7667;
  assign new_P2_U2728 = ~new_P2_U7673 | ~new_P2_U7674 | ~new_P2_U7676 | ~new_P2_U7675;
  assign new_P2_U2729 = ~new_P2_U7677 | ~new_P2_U7678 | ~new_P2_U7680 | ~new_P2_U7679;
  assign new_P2_U2730 = ~new_P2_U7681 | ~new_P2_U7682 | ~new_P2_U7684 | ~new_P2_U7683;
  assign new_P2_U2731 = ~new_P2_U7685 | ~new_P2_U7686 | ~new_P2_U7688 | ~new_P2_U7687;
  assign new_P2_U2732 = ~new_P2_U7689 | ~new_P2_U7690 | ~new_P2_U7692 | ~new_P2_U7691;
  assign new_P2_U2733 = ~new_P2_U7693 | ~new_P2_U7694 | ~new_P2_U7696 | ~new_P2_U7695;
  assign new_P2_U2734 = ~new_P2_U7697 | ~new_P2_U7698 | ~new_P2_U7700 | ~new_P2_U7699;
  assign new_P2_U2735 = ~new_P2_U7701 | ~new_P2_U7702 | ~new_P2_U7704 | ~new_P2_U7703;
  assign new_P2_U2736 = ~new_P2_U7705 | ~new_P2_U7706 | ~new_P2_U7708 | ~new_P2_U7707;
  assign new_P2_U2737 = ~new_P2_U7709 | ~new_P2_U7710 | ~new_P2_U7712 | ~new_P2_U7711;
  assign new_P2_U2738 = ~new_P2_U7593 | ~new_P2_U7594 | ~new_P2_U7596 | ~new_P2_U7595;
  assign new_P2_U2739 = ~new_P2_U7597 | ~new_P2_U7598 | ~new_P2_U7600 | ~new_P2_U7599;
  assign new_P2_U2740 = ~new_P2_U7601 | ~new_P2_U7602 | ~new_P2_U7604 | ~new_P2_U7603;
  assign new_P2_U2741 = ~new_P2_U7605 | ~new_P2_U7606 | ~new_P2_U7608 | ~new_P2_U7607;
  assign new_P2_U2742 = ~new_P2_U7609 | ~new_P2_U7610 | ~new_P2_U7612 | ~new_P2_U7611;
  assign new_P2_U2743 = ~new_P2_U7613 | ~new_P2_U7614 | ~new_P2_U7616 | ~new_P2_U7615;
  assign new_P2_U2744 = ~new_P2_U7625 | ~new_P2_U7626 | ~new_P2_U7628 | ~new_P2_U7627;
  assign new_P2_U2745 = ~new_P2_U7669 | ~new_P2_U7670 | ~new_P2_U7672 | ~new_P2_U7671;
  assign new_P2_U2746 = ~new_P2_U7713 | ~new_P2_U7714 | ~new_P2_U7716 | ~new_P2_U7715;
  assign new_P2_U2747 = ~new_P2_U7717 | ~new_P2_U4388 | ~new_P2_U4389 | ~new_P2_U7886 | ~new_P2_U7721;
  assign new_P2_U2748 = ~new_P2_U7583 | ~new_P2_U7582;
  assign new_P2_U2749 = ~new_P2_U4380 | ~new_P2_U7584;
  assign new_P2_U2750 = ~new_P2_U4382 | ~new_P2_U7588;
  assign new_P2_U2751 = new_P2_U7888 & new_P2_U7737;
  assign new_P2_U2752 = new_P2_U7873 & new_P2_U3280 & P2_INSTQUEUERD_ADDR_REG_4_;
  assign new_P2_U2753 = ~new_P2_U3286 | ~new_P2_U7572;
  assign new_P2_U2754 = ~new_P2_U3286 | ~new_P2_U7573;
  assign new_P2_U2755 = ~new_P2_U3286 | ~new_P2_U7574;
  assign new_P2_U2756 = ~new_P2_U3286 | ~new_P2_U7575;
  assign new_P2_U2757 = ~new_P2_U3286 | ~new_P2_U7576;
  assign new_P2_U2758 = new_P2_U4428 & new_P2_U3242;
  assign new_P2_U2759 = new_P2_U4428 & new_P2_U7217;
  assign new_P2_U2760 = new_P2_U4428 & new_P2_U7251;
  assign new_P2_U2761 = ~new_P2_U7563 | ~new_P2_U7562;
  assign new_P2_U2762 = ~new_P2_U7565 | ~new_P2_U7564;
  assign new_P2_U2763 = ~new_P2_U7567 | ~new_P2_U7566;
  assign new_P2_U2764 = ~new_P2_U7569 | ~new_P2_U7568;
  assign new_P2_U2765 = ~new_P2_U7571 | ~new_P2_U7570;
  assign new_P2_U2766 = ~new_P2_U4447 | ~new_P2_U7539;
  assign new_P2_U2767 = ~new_P2_U4447 | ~new_P2_U7540;
  assign new_P2_U2768 = ~new_P2_U4447 | ~new_P2_U7541;
  assign new_P2_U2769 = ~new_P2_U4447 | ~new_P2_U7542;
  assign new_P2_U2770 = ~new_P2_U4447 | ~new_P2_U7543;
  assign new_P2_U2771 = ~new_P2_U4447 | ~new_P2_U7544;
  assign new_P2_U2772 = ~new_P2_U4447 | ~new_P2_U7545;
  assign new_P2_U2773 = ~new_P2_U4447 | ~new_P2_U7546;
  assign new_P2_U2774 = ~new_P2_U4447 | ~new_P2_U7547;
  assign new_P2_U2775 = ~new_P2_U4447 | ~new_P2_U7548;
  assign new_P2_U2776 = ~new_P2_U4447 | ~new_P2_U7549;
  assign new_P2_U2777 = ~new_P2_U4447 | ~new_P2_U7550;
  assign new_P2_U2778 = ~new_P2_U4447 | ~new_P2_U7551;
  assign new_P2_U2779 = ~new_P2_U4447 | ~new_P2_U7552;
  assign new_P2_U2780 = ~new_P2_U4447 | ~new_P2_U7553;
  assign new_P2_U2781 = ~new_P2_U4447 | ~new_P2_U7554;
  assign new_P2_U2782 = ~new_P2_U4447 | ~new_P2_U7555;
  assign new_P2_U2783 = ~new_P2_U4447 | ~new_P2_U7556;
  assign new_P2_U2784 = ~new_P2_U4447 | ~new_P2_U7557;
  assign new_P2_U2785 = ~new_P2_U4447 | ~new_P2_U7558;
  assign new_P2_U2786 = ~new_P2_U4447 | ~new_P2_U7559;
  assign new_P2_U2787 = ~new_P2_U4447 | ~new_P2_U7560;
  assign new_P2_U2788 = ~new_P2_U4447 | ~new_P2_U7537;
  assign new_P2_U2789 = ~new_P2_U4447 | ~new_P2_U7538;
  assign new_P2_U2790 = new_P2_U3242 & new_P2_R2267_U63;
  assign new_P2_U2791 = new_P2_U3242 & new_P2_R2267_U16;
  assign new_P2_U2792 = new_P2_U3242 & new_P2_R2267_U15;
  assign new_P2_U2793 = new_P2_U3242 & new_P2_R2267_U67;
  assign new_P2_U2794 = new_P2_U3242 & new_P2_R2267_U14;
  assign new_P2_U2795 = new_P2_U3242 & new_P2_R2267_U69;
  assign new_P2_U2796 = new_P2_U3242 & new_P2_R2267_U13;
  assign new_P2_U2797 = new_P2_U3242 & new_P2_R2267_U71;
  assign new_P2_U2798 = new_P2_U3242 & new_P2_R2267_U12;
  assign new_P2_U2799 = new_P2_U3242 & new_P2_R2267_U73;
  assign new_P2_U2800 = new_P2_U3242 & new_P2_R2267_U11;
  assign new_P2_U2801 = new_P2_U3242 & new_P2_R2267_U75;
  assign new_P2_U2802 = new_P2_U3242 & new_P2_R2267_U10;
  assign new_P2_U2803 = new_P2_U3242 & new_P2_R2267_U79;
  assign new_P2_U2804 = new_P2_U3242 & new_P2_R2267_U9;
  assign new_P2_U2805 = new_P2_U3242 & new_P2_R2267_U81;
  assign new_P2_U2806 = new_P2_U3242 & new_P2_R2267_U8;
  assign new_P2_U2807 = new_P2_U3242 & new_P2_R2267_U83;
  assign new_P2_U2808 = new_P2_U3242 & new_P2_R2267_U7;
  assign new_P2_U2809 = new_P2_U3242 & new_P2_R2267_U85;
  assign new_P2_U2810 = new_P2_U3242 & new_P2_R2267_U6;
  assign new_P2_U2811 = new_P2_U3242 & new_P2_R2267_U87;
  assign new_P2_U2812 = new_P2_U3242 & new_P2_R2267_U20;
  assign new_P2_U2813 = P2_INSTQUEUERD_ADDR_REG_3_ & new_P2_U3519;
  assign n5069 = ~new_P2_U4190 | ~new_P2_U6861;
  assign n5059 = ~new_P2_U7917 | ~new_P2_U6856;
  assign n5054 = ~new_P2_U6855 | ~new_P2_U6854;
  assign n5044 = ~new_P2_U4463 | ~new_P2_U8140 | ~new_P2_U8139;
  assign n5034 = ~new_P2_U4463 | ~new_P2_U8136 | ~new_P2_U8135;
  assign n5024 = ~new_P2_U6840 | ~new_P2_U6839;
  assign n5014 = ~new_P2_U3548 | ~new_P2_U8128 | ~new_P2_U8127;
  assign n5009 = ~new_P2_U6837 | ~new_P2_U3548 | ~new_P2_U4452;
  assign n5004 = ~new_P2_U4398 | ~new_P2_U6836;
  assign n4999 = ~new_P2_U4452 | ~new_P2_U8124 | ~new_P2_U8123;
  assign n4994 = ~new_P2_U6828 | ~new_P2_U6830 | ~new_P2_U4168 | ~new_P2_U6827 | ~new_P2_U6829;
  assign n4989 = ~new_P2_U6820 | ~new_P2_U6822 | ~new_P2_U4166 | ~new_P2_U6819 | ~new_P2_U6821;
  assign n4984 = ~new_P2_U6812 | ~new_P2_U6814 | ~new_P2_U4164 | ~new_P2_U6811 | ~new_P2_U6813;
  assign n4979 = ~new_P2_U6804 | ~new_P2_U6806 | ~new_P2_U4162 | ~new_P2_U6803 | ~new_P2_U6805;
  assign n4974 = ~new_P2_U6796 | ~new_P2_U6798 | ~new_P2_U4160 | ~new_P2_U6795 | ~new_P2_U6797;
  assign n4969 = ~new_P2_U6788 | ~new_P2_U6790 | ~new_P2_U4158 | ~new_P2_U6787 | ~new_P2_U6789;
  assign n4964 = ~new_P2_U6780 | ~new_P2_U4156 | ~new_P2_U6782 | ~new_P2_U6779 | ~new_P2_U6781;
  assign n4959 = ~new_P2_U6772 | ~new_P2_U4152;
  assign n4954 = ~new_P2_U6764 | ~new_P2_U4149;
  assign n4949 = ~new_P2_U4148 | ~new_P2_U6756 | ~new_P2_U6758 | ~new_P2_U6755 | ~new_P2_U6757;
  assign n4944 = ~new_P2_U4146 | ~new_P2_U4144;
  assign n4939 = ~new_P2_U4143 | ~new_P2_U4141;
  assign n4934 = ~new_P2_U4140 | ~new_P2_U4138;
  assign n4929 = ~new_P2_U4136 | ~new_P2_U4134;
  assign n4924 = ~new_P2_U4132 | ~new_P2_U4130;
  assign n4919 = ~new_P2_U4128 | ~new_P2_U4126;
  assign n4914 = ~new_P2_U4124 | ~new_P2_U4122;
  assign n4909 = ~new_P2_U4119 | ~new_P2_U6696 | ~new_P2_U6692 | ~new_P2_U6693 | ~new_P2_U4118;
  assign n4904 = ~new_P2_U4116 | ~new_P2_U6688 | ~new_P2_U6684 | ~new_P2_U6685 | ~new_P2_U4115;
  assign n4899 = ~new_P2_U4113 | ~new_P2_U6680 | ~new_P2_U6676 | ~new_P2_U6677 | ~new_P2_U4112;
  assign n4894 = ~new_P2_U4110 | ~new_P2_U6672 | ~new_P2_U4109 | ~new_P2_U6670 | ~new_P2_U6669;
  assign n4889 = ~new_P2_U4107 | ~new_P2_U6664 | ~new_P2_U4106 | ~new_P2_U6662 | ~new_P2_U6661;
  assign n4884 = ~new_P2_U4104 | ~new_P2_U6656 | ~new_P2_U4103 | ~new_P2_U6654 | ~new_P2_U6653;
  assign n4879 = ~new_P2_U4101 | ~new_P2_U6648 | ~new_P2_U4100 | ~new_P2_U6646 | ~new_P2_U6645;
  assign n4874 = ~new_P2_U4098 | ~new_P2_U6640 | ~new_P2_U4097 | ~new_P2_U6638 | ~new_P2_U6637;
  assign n4869 = ~new_P2_U4095 | ~new_P2_U6632 | ~new_P2_U4094 | ~new_P2_U6630 | ~new_P2_U6629;
  assign n4864 = ~new_P2_U4093 | ~new_P2_U4091;
  assign n4859 = ~new_P2_U4089 | ~new_P2_U4087;
  assign n4854 = ~new_P2_U4084 | ~new_P2_U6606 | ~new_P2_U6602 | ~new_P2_U4082;
  assign n4849 = ~new_P2_U4080 | ~new_P2_U6597 | ~new_P2_U6593 | ~new_P2_U4078;
  assign n4844 = ~new_P2_U4076 | ~new_P2_U6588 | ~new_P2_U6584 | ~new_P2_U4074;
  assign n4839 = ~new_P2_U4072 | ~new_P2_U6579 | ~new_P2_U6575 | ~new_P2_U4070;
  assign n4834 = ~new_P2_U6565 | ~new_P2_U6564;
  assign n4829 = ~new_P2_U6561 | ~new_P2_U6562 | ~new_P2_U6563;
  assign n4824 = ~new_P2_U6558 | ~new_P2_U6559 | ~new_P2_U6560;
  assign n4819 = ~new_P2_U6555 | ~new_P2_U6556 | ~new_P2_U6557;
  assign n4814 = ~new_P2_U6552 | ~new_P2_U6553 | ~new_P2_U6554;
  assign n4809 = ~new_P2_U6549 | ~new_P2_U6550 | ~new_P2_U6551;
  assign n4804 = ~new_P2_U6546 | ~new_P2_U6547 | ~new_P2_U6548;
  assign n4799 = ~new_P2_U6543 | ~new_P2_U6544 | ~new_P2_U6545;
  assign n4794 = ~new_P2_U6540 | ~new_P2_U6541 | ~new_P2_U6542;
  assign n4789 = ~new_P2_U6537 | ~new_P2_U6538 | ~new_P2_U6539;
  assign n4784 = ~new_P2_U6534 | ~new_P2_U6535 | ~new_P2_U6536;
  assign n4779 = ~new_P2_U6531 | ~new_P2_U6532 | ~new_P2_U6533;
  assign n4774 = ~new_P2_U6528 | ~new_P2_U6529 | ~new_P2_U6530;
  assign n4769 = ~new_P2_U6525 | ~new_P2_U6526 | ~new_P2_U6527;
  assign n4764 = ~new_P2_U6522 | ~new_P2_U6523 | ~new_P2_U6524;
  assign n4759 = ~new_P2_U6519 | ~new_P2_U6520 | ~new_P2_U6521;
  assign n4754 = ~new_P2_U6516 | ~new_P2_U6517 | ~new_P2_U6518;
  assign n4749 = ~new_P2_U6513 | ~new_P2_U6514 | ~new_P2_U6515;
  assign n4744 = ~new_P2_U6510 | ~new_P2_U6511 | ~new_P2_U6512;
  assign n4739 = ~new_P2_U6507 | ~new_P2_U6508 | ~new_P2_U6509;
  assign n4734 = ~new_P2_U6504 | ~new_P2_U6505 | ~new_P2_U6506;
  assign n4729 = ~new_P2_U6501 | ~new_P2_U6502 | ~new_P2_U6503;
  assign n4724 = ~new_P2_U6498 | ~new_P2_U6499 | ~new_P2_U6500;
  assign n4719 = ~new_P2_U6495 | ~new_P2_U6496 | ~new_P2_U6497;
  assign n4714 = ~new_P2_U6494 | ~new_P2_U6493 | ~new_P2_U6492;
  assign n4709 = ~new_P2_U6491 | ~new_P2_U6490 | ~new_P2_U6489;
  assign n4704 = ~new_P2_U6488 | ~new_P2_U6487 | ~new_P2_U6486;
  assign n4699 = ~new_P2_U6485 | ~new_P2_U6484 | ~new_P2_U6483;
  assign n4694 = ~new_P2_U6482 | ~new_P2_U6481 | ~new_P2_U6480;
  assign n4689 = ~new_P2_U6479 | ~new_P2_U6478 | ~new_P2_U6477;
  assign n4684 = ~new_P2_U6476 | ~new_P2_U6475 | ~new_P2_U6474;
  assign n4679 = ~new_P2_U6473 | ~new_P2_U6472 | ~new_P2_U6471;
  assign n4674 = ~new_P2_U6467 | ~new_P2_U6468 | ~new_P2_U6466;
  assign n4669 = ~new_P2_U6463 | ~new_P2_U6464 | ~new_P2_U6465 | ~new_P2_U6462 | ~new_P2_U6461;
  assign n4664 = ~new_P2_U6458 | ~new_P2_U6459 | ~new_P2_U6460 | ~new_P2_U6457 | ~new_P2_U6456;
  assign n4659 = ~new_P2_U6453 | ~new_P2_U6454 | ~new_P2_U6455 | ~new_P2_U6452 | ~new_P2_U6451;
  assign n4654 = ~new_P2_U6448 | ~new_P2_U6449 | ~new_P2_U6450 | ~new_P2_U6447 | ~new_P2_U6446;
  assign n4649 = ~new_P2_U6443 | ~new_P2_U6444 | ~new_P2_U6445 | ~new_P2_U6442 | ~new_P2_U6441;
  assign n4644 = ~new_P2_U6438 | ~new_P2_U6439 | ~new_P2_U6440 | ~new_P2_U6437 | ~new_P2_U6436;
  assign n4639 = ~new_P2_U6433 | ~new_P2_U6434 | ~new_P2_U6435 | ~new_P2_U6432 | ~new_P2_U6431;
  assign n4634 = ~new_P2_U6428 | ~new_P2_U6429 | ~new_P2_U6430 | ~new_P2_U6427 | ~new_P2_U6426;
  assign n4629 = ~new_P2_U6423 | ~new_P2_U6424 | ~new_P2_U6425 | ~new_P2_U6422 | ~new_P2_U6421;
  assign n4624 = ~new_P2_U6418 | ~new_P2_U6419 | ~new_P2_U6420 | ~new_P2_U6417 | ~new_P2_U6416;
  assign n4619 = ~new_P2_U6413 | ~new_P2_U6414 | ~new_P2_U6415 | ~new_P2_U6412 | ~new_P2_U6411;
  assign n4614 = ~new_P2_U6408 | ~new_P2_U6409 | ~new_P2_U6410 | ~new_P2_U6407 | ~new_P2_U6406;
  assign n4609 = ~new_P2_U6403 | ~new_P2_U6404 | ~new_P2_U6405 | ~new_P2_U6402 | ~new_P2_U6401;
  assign n4604 = ~new_P2_U6398 | ~new_P2_U6399 | ~new_P2_U6400 | ~new_P2_U6397 | ~new_P2_U6396;
  assign n4599 = ~new_P2_U6393 | ~new_P2_U6394 | ~new_P2_U6395 | ~new_P2_U6392 | ~new_P2_U6391;
  assign n4594 = ~new_P2_U6388 | ~new_P2_U6389 | ~new_P2_U6390 | ~new_P2_U6387;
  assign n4589 = ~new_P2_U6384 | ~new_P2_U6385 | ~new_P2_U6386 | ~new_P2_U6383;
  assign n4584 = ~new_P2_U6380 | ~new_P2_U6381 | ~new_P2_U6382 | ~new_P2_U6379;
  assign n4579 = ~new_P2_U6376 | ~new_P2_U6377 | ~new_P2_U6378 | ~new_P2_U6375;
  assign n4574 = ~new_P2_U6372 | ~new_P2_U6373 | ~new_P2_U6374 | ~new_P2_U6371;
  assign n4569 = ~new_P2_U6368 | ~new_P2_U6369 | ~new_P2_U6370 | ~new_P2_U6367;
  assign n4564 = ~new_P2_U6364 | ~new_P2_U4068 | ~new_P2_U6363;
  assign n4559 = ~new_P2_U6360 | ~new_P2_U4067 | ~new_P2_U6359;
  assign n4554 = ~new_P2_U6356 | ~new_P2_U4066 | ~new_P2_U6355;
  assign n4549 = ~new_P2_U4065 | ~new_P2_U6352 | ~new_P2_U6351;
  assign n4544 = ~new_P2_U4064 | ~new_P2_U6348 | ~new_P2_U6347;
  assign n4539 = ~new_P2_U4063 | ~new_P2_U6344 | ~new_P2_U6343;
  assign n4534 = ~new_P2_U4062 | ~new_P2_U6340 | ~new_P2_U6339;
  assign n4529 = ~new_P2_U4061 | ~new_P2_U6336 | ~new_P2_U6335;
  assign n4524 = ~new_P2_U4060 | ~new_P2_U6332 | ~new_P2_U6331;
  assign n4519 = ~new_P2_U4059 | ~new_P2_U6328 | ~new_P2_U6327;
  assign n4514 = P2_DATAO_REG_31_ & new_P2_U6232;
  assign n4509 = ~new_P2_U6325 | ~new_P2_U6324 | ~new_P2_U6323;
  assign n4504 = ~new_P2_U6322 | ~new_P2_U6321 | ~new_P2_U6320;
  assign n4499 = ~new_P2_U6319 | ~new_P2_U6318 | ~new_P2_U6317;
  assign n4494 = ~new_P2_U6316 | ~new_P2_U6315 | ~new_P2_U6314;
  assign n4489 = ~new_P2_U6313 | ~new_P2_U6312 | ~new_P2_U6311;
  assign n4484 = ~new_P2_U6310 | ~new_P2_U6309 | ~new_P2_U6308;
  assign n4479 = ~new_P2_U6307 | ~new_P2_U6306 | ~new_P2_U6305;
  assign n4474 = ~new_P2_U6304 | ~new_P2_U6303 | ~new_P2_U6302;
  assign n4469 = ~new_P2_U6301 | ~new_P2_U6300 | ~new_P2_U6299;
  assign n4464 = ~new_P2_U6298 | ~new_P2_U6297 | ~new_P2_U6296;
  assign n4459 = ~new_P2_U6295 | ~new_P2_U6294 | ~new_P2_U6293;
  assign n4454 = ~new_P2_U6292 | ~new_P2_U6291 | ~new_P2_U6290;
  assign n4449 = ~new_P2_U6289 | ~new_P2_U6288 | ~new_P2_U6287;
  assign n4444 = ~new_P2_U6286 | ~new_P2_U6285 | ~new_P2_U6284;
  assign n4439 = ~new_P2_U6283 | ~new_P2_U6282 | ~new_P2_U6281;
  assign n4434 = ~new_P2_U6280 | ~new_P2_U6279 | ~new_P2_U6278;
  assign n4429 = ~new_P2_U6277 | ~new_P2_U6276 | ~new_P2_U6275;
  assign n4424 = ~new_P2_U6274 | ~new_P2_U6273 | ~new_P2_U6272;
  assign n4419 = ~new_P2_U6271 | ~new_P2_U6270 | ~new_P2_U6269;
  assign n4414 = ~new_P2_U6268 | ~new_P2_U6267 | ~new_P2_U6266;
  assign n4409 = ~new_P2_U6265 | ~new_P2_U6264 | ~new_P2_U6263;
  assign n4404 = ~new_P2_U6262 | ~new_P2_U6261 | ~new_P2_U6260;
  assign n4399 = ~new_P2_U6259 | ~new_P2_U6258 | ~new_P2_U6257;
  assign n4394 = ~new_P2_U6256 | ~new_P2_U6255 | ~new_P2_U6254;
  assign n4389 = ~new_P2_U6253 | ~new_P2_U6252 | ~new_P2_U6251;
  assign n4384 = ~new_P2_U6250 | ~new_P2_U6249 | ~new_P2_U6248;
  assign n4379 = ~new_P2_U6247 | ~new_P2_U6246 | ~new_P2_U6245;
  assign n4374 = ~new_P2_U6244 | ~new_P2_U6243 | ~new_P2_U6242;
  assign n4369 = ~new_P2_U6241 | ~new_P2_U6240 | ~new_P2_U6239;
  assign n4364 = ~new_P2_U6238 | ~new_P2_U6237 | ~new_P2_U6236;
  assign n4359 = ~new_P2_U6235 | ~new_P2_U6234 | ~new_P2_U6233;
  assign n4354 = ~new_P2_U6226 | ~new_P2_U6225 | ~new_P2_U6224;
  assign n4349 = ~new_P2_U6223 | ~new_P2_U6222 | ~new_P2_U6221;
  assign n4344 = ~new_P2_U6220 | ~new_P2_U6219 | ~new_P2_U6218;
  assign n4339 = ~new_P2_U6217 | ~new_P2_U6216 | ~new_P2_U6215;
  assign n4334 = ~new_P2_U6214 | ~new_P2_U6213 | ~new_P2_U6212;
  assign n4329 = ~new_P2_U6211 | ~new_P2_U6210 | ~new_P2_U6209;
  assign n4324 = ~new_P2_U6208 | ~new_P2_U6207 | ~new_P2_U6206;
  assign n4319 = ~new_P2_U6205 | ~new_P2_U6204 | ~new_P2_U6203;
  assign n4314 = ~new_P2_U6202 | ~new_P2_U6201 | ~new_P2_U6200;
  assign n4309 = ~new_P2_U6199 | ~new_P2_U6198 | ~new_P2_U6197;
  assign n4304 = ~new_P2_U6196 | ~new_P2_U6195 | ~new_P2_U6194;
  assign n4299 = ~new_P2_U6193 | ~new_P2_U6192 | ~new_P2_U6191;
  assign n4294 = ~new_P2_U6190 | ~new_P2_U6189 | ~new_P2_U6188;
  assign n4289 = ~new_P2_U6187 | ~new_P2_U6186 | ~new_P2_U6185;
  assign n4284 = ~new_P2_U6184 | ~new_P2_U6183 | ~new_P2_U6182;
  assign n4279 = ~new_P2_U6181 | ~new_P2_U6180 | ~new_P2_U6179;
  assign n4274 = ~new_P2_U6178 | ~new_P2_U6177 | ~new_P2_U6176;
  assign n4269 = ~new_P2_U6175 | ~new_P2_U6174 | ~new_P2_U6173;
  assign n4264 = ~new_P2_U6172 | ~new_P2_U6171 | ~new_P2_U6170;
  assign n4259 = ~new_P2_U6169 | ~new_P2_U6168 | ~new_P2_U6167;
  assign n4254 = ~new_P2_U6166 | ~new_P2_U6165 | ~new_P2_U6164;
  assign n4249 = ~new_P2_U6163 | ~new_P2_U6162 | ~new_P2_U6161;
  assign n4244 = ~new_P2_U6160 | ~new_P2_U6159 | ~new_P2_U6158;
  assign n4239 = ~new_P2_U6157 | ~new_P2_U6156 | ~new_P2_U6155;
  assign n4234 = ~new_P2_U6154 | ~new_P2_U6153 | ~new_P2_U6152;
  assign n4229 = ~new_P2_U6151 | ~new_P2_U6150 | ~new_P2_U6149;
  assign n4224 = ~new_P2_U6148 | ~new_P2_U6147 | ~new_P2_U6146;
  assign n4219 = ~new_P2_U6145 | ~new_P2_U6144 | ~new_P2_U6143;
  assign n4214 = ~new_P2_U6142 | ~new_P2_U6141 | ~new_P2_U6140;
  assign n4209 = ~new_P2_U6139 | ~new_P2_U6138 | ~new_P2_U6137;
  assign n4204 = ~new_P2_U6136 | ~new_P2_U6135 | ~new_P2_U6134;
  assign n4199 = ~new_P2_U4054 | ~new_P2_U4053;
  assign n4194 = ~new_P2_U4052 | ~new_P2_U4051;
  assign n4189 = ~new_P2_U4050 | ~new_P2_U4049;
  assign n4184 = ~new_P2_U4048 | ~new_P2_U4047;
  assign n4179 = ~new_P2_U4046 | ~new_P2_U4045;
  assign n4174 = ~new_P2_U4044 | ~new_P2_U4043;
  assign n4169 = ~new_P2_U4042 | ~new_P2_U4041;
  assign n4164 = ~new_P2_U4040 | ~new_P2_U4039;
  assign n4159 = ~new_P2_U4038 | ~new_P2_U4037;
  assign n4154 = ~new_P2_U4036 | ~new_P2_U4035;
  assign n4149 = ~new_P2_U4034 | ~new_P2_U4033;
  assign n4144 = ~new_P2_U4032 | ~new_P2_U4031;
  assign n4139 = ~new_P2_U4030 | ~new_P2_U4029;
  assign n4134 = ~new_P2_U4028 | ~new_P2_U4027;
  assign n4129 = ~new_P2_U4026 | ~new_P2_U4025;
  assign n4124 = ~new_P2_U4024 | ~new_P2_U4023;
  assign n4119 = ~new_P2_U4022 | ~new_P2_U4021;
  assign n4114 = ~new_P2_U4020 | ~new_P2_U4019;
  assign n4109 = ~new_P2_U4018 | ~new_P2_U4017;
  assign n4104 = ~new_P2_U4016 | ~new_P2_U4015;
  assign n4099 = ~new_P2_U4014 | ~new_P2_U4013;
  assign n4094 = ~new_P2_U4012 | ~new_P2_U4011;
  assign n4089 = ~new_P2_U4010 | ~new_P2_U4009;
  assign n4084 = ~new_P2_U4008 | ~new_P2_U4007;
  assign n4079 = ~new_P2_U4006 | ~new_P2_U4005;
  assign n4074 = ~new_P2_U4004 | ~new_P2_U4003;
  assign n4069 = ~new_P2_U4002 | ~new_P2_U4001;
  assign n4064 = ~new_P2_U4000 | ~new_P2_U3999;
  assign n4059 = ~new_P2_U3998 | ~new_P2_U3997;
  assign n4054 = ~new_P2_U3996 | ~new_P2_U3995;
  assign n4049 = ~new_P2_U3994 | ~new_P2_U3993;
  assign n4044 = ~new_P2_U3992 | ~new_P2_U3991;
  assign n4039 = ~new_P2_U5928 | ~new_P2_U3987 | ~new_P2_U3988 | ~new_P2_U5933 | ~new_P2_U5932;
  assign n4034 = ~new_P2_U5920 | ~new_P2_U3985 | ~new_P2_U3986 | ~new_P2_U5925 | ~new_P2_U5924;
  assign n4029 = ~new_P2_U3983 | ~new_P2_U3984 | ~new_P2_U5917 | ~new_P2_U5916;
  assign n4024 = ~new_P2_U3980 | ~new_P2_U3981 | ~new_P2_U3982 | ~new_P2_U5909 | ~new_P2_U5908;
  assign n4019 = ~new_P2_U3977 | ~new_P2_U3978 | ~new_P2_U3979 | ~new_P2_U5901 | ~new_P2_U5900;
  assign n4014 = ~new_P2_U3974 | ~new_P2_U3975 | ~new_P2_U3976 | ~new_P2_U5893 | ~new_P2_U5892;
  assign n4009 = ~new_P2_U3971 | ~new_P2_U3972 | ~new_P2_U3973 | ~new_P2_U5885 | ~new_P2_U5884;
  assign n4004 = ~new_P2_U3968 | ~new_P2_U3969 | ~new_P2_U3970 | ~new_P2_U5877 | ~new_P2_U5876;
  assign n3999 = ~new_P2_U3965 | ~new_P2_U3966 | ~new_P2_U3967 | ~new_P2_U5869 | ~new_P2_U5868;
  assign n3994 = ~new_P2_U3962 | ~new_P2_U3963 | ~new_P2_U3964 | ~new_P2_U5861 | ~new_P2_U5860;
  assign n3989 = ~new_P2_U3959 | ~new_P2_U3960 | ~new_P2_U3961 | ~new_P2_U5853 | ~new_P2_U5852;
  assign n3984 = ~new_P2_U3956 | ~new_P2_U3957 | ~new_P2_U3958 | ~new_P2_U5845 | ~new_P2_U5844;
  assign n3979 = ~new_P2_U3953 | ~new_P2_U3954 | ~new_P2_U3955 | ~new_P2_U5837 | ~new_P2_U5836;
  assign n3974 = ~new_P2_U3950 | ~new_P2_U3951 | ~new_P2_U3952 | ~new_P2_U5829 | ~new_P2_U5828;
  assign n3969 = ~new_P2_U3947 | ~new_P2_U3948 | ~new_P2_U3949 | ~new_P2_U5821 | ~new_P2_U5820;
  assign n3964 = ~new_P2_U3944 | ~new_P2_U3945 | ~new_P2_U3946 | ~new_P2_U5813 | ~new_P2_U5812;
  assign n3959 = ~new_P2_U3941 | ~new_P2_U3942 | ~new_P2_U3943 | ~new_P2_U5805 | ~new_P2_U5804;
  assign n3954 = ~new_P2_U3938 | ~new_P2_U3939 | ~new_P2_U3940 | ~new_P2_U5797 | ~new_P2_U5796;
  assign n3949 = ~new_P2_U3935 | ~new_P2_U3936 | ~new_P2_U3937 | ~new_P2_U5789 | ~new_P2_U5788;
  assign n3944 = ~new_P2_U3932 | ~new_P2_U3933 | ~new_P2_U3934 | ~new_P2_U5781 | ~new_P2_U5780;
  assign n3939 = ~new_P2_U3929 | ~new_P2_U3930 | ~new_P2_U3931 | ~new_P2_U5773 | ~new_P2_U5772;
  assign n3934 = ~new_P2_U3926 | ~new_P2_U3927 | ~new_P2_U3928 | ~new_P2_U5765 | ~new_P2_U5764;
  assign n3929 = ~new_P2_U3923 | ~new_P2_U3924 | ~new_P2_U3925 | ~new_P2_U5757 | ~new_P2_U5756;
  assign n3924 = ~new_P2_U3920 | ~new_P2_U3921 | ~new_P2_U3922 | ~new_P2_U5749 | ~new_P2_U5748;
  assign n3919 = ~new_P2_U3917 | ~new_P2_U3918 | ~new_P2_U3919 | ~new_P2_U5741 | ~new_P2_U5740;
  assign n3914 = ~new_P2_U3914 | ~new_P2_U3915 | ~new_P2_U3916 | ~new_P2_U5733 | ~new_P2_U5732;
  assign n3909 = ~new_P2_U3911 | ~new_P2_U3912 | ~new_P2_U3913 | ~new_P2_U5725 | ~new_P2_U5724;
  assign n3904 = ~new_P2_U3908 | ~new_P2_U3909 | ~new_P2_U3910 | ~new_P2_U5717 | ~new_P2_U5716;
  assign n3899 = ~new_P2_U3905 | ~new_P2_U3906 | ~new_P2_U3907 | ~new_P2_U5709 | ~new_P2_U5708;
  assign n3894 = ~new_P2_U3902 | ~new_P2_U3903 | ~new_P2_U3904 | ~new_P2_U5701 | ~new_P2_U5700;
  assign n3889 = ~new_P2_U3899 | ~new_P2_U3900 | ~new_P2_U3901 | ~new_P2_U5693 | ~new_P2_U5692;
  assign n3884 = ~new_P2_U3896 | ~new_P2_U3897 | ~new_P2_U3898 | ~new_P2_U5685 | ~new_P2_U5684;
  assign n3859 = P2_INSTQUEUEWR_ADDR_REG_4_ & new_P2_U5643;
  assign n3829 = ~new_P2_U3865 | ~new_P2_U5570 | ~new_P2_U5569;
  assign n3824 = ~new_P2_U3864 | ~new_P2_U5565 | ~new_P2_U5564;
  assign n3819 = ~new_P2_U3863 | ~new_P2_U5560 | ~new_P2_U5559;
  assign n3814 = ~new_P2_U3862 | ~new_P2_U5555 | ~new_P2_U5554;
  assign n3809 = ~new_P2_U3861 | ~new_P2_U5550 | ~new_P2_U5549;
  assign n3804 = ~new_P2_U3860 | ~new_P2_U5545 | ~new_P2_U5544;
  assign n3799 = ~new_P2_U3859 | ~new_P2_U5540 | ~new_P2_U5539;
  assign n3794 = ~new_P2_U3858 | ~new_P2_U5535 | ~new_P2_U5534;
  assign n3789 = ~new_P2_U3856 | ~new_P2_U5513 | ~new_P2_U5512;
  assign n3784 = ~new_P2_U3855 | ~new_P2_U5508 | ~new_P2_U5507;
  assign n3779 = ~new_P2_U3854 | ~new_P2_U5503 | ~new_P2_U5502;
  assign n3774 = ~new_P2_U3853 | ~new_P2_U5498 | ~new_P2_U5497;
  assign n3769 = ~new_P2_U3852 | ~new_P2_U5493 | ~new_P2_U5492;
  assign n3764 = ~new_P2_U3851 | ~new_P2_U5488 | ~new_P2_U5487;
  assign n3759 = ~new_P2_U3850 | ~new_P2_U5483 | ~new_P2_U5482;
  assign n3754 = ~new_P2_U3849 | ~new_P2_U5478 | ~new_P2_U5477;
  assign n3749 = ~new_P2_U3847 | ~new_P2_U5455 | ~new_P2_U5454;
  assign n3744 = ~new_P2_U3846 | ~new_P2_U5450 | ~new_P2_U5449;
  assign n3739 = ~new_P2_U3845 | ~new_P2_U5445 | ~new_P2_U5444;
  assign n3734 = ~new_P2_U3844 | ~new_P2_U5440 | ~new_P2_U5439;
  assign n3729 = ~new_P2_U3843 | ~new_P2_U5435 | ~new_P2_U5434;
  assign n3724 = ~new_P2_U3842 | ~new_P2_U5430 | ~new_P2_U5429;
  assign n3719 = ~new_P2_U3841 | ~new_P2_U5425 | ~new_P2_U5424;
  assign n3714 = ~new_P2_U3840 | ~new_P2_U5420 | ~new_P2_U5419;
  assign n3709 = ~new_P2_U3838 | ~new_P2_U5398 | ~new_P2_U5397;
  assign n3704 = ~new_P2_U3837 | ~new_P2_U5393 | ~new_P2_U5392;
  assign n3699 = ~new_P2_U3836 | ~new_P2_U5388 | ~new_P2_U5387;
  assign n3694 = ~new_P2_U3835 | ~new_P2_U5383 | ~new_P2_U5382;
  assign n3689 = ~new_P2_U3834 | ~new_P2_U5378 | ~new_P2_U5377;
  assign n3684 = ~new_P2_U3833 | ~new_P2_U5373 | ~new_P2_U5372;
  assign n3679 = ~new_P2_U3832 | ~new_P2_U5368 | ~new_P2_U5367;
  assign n3674 = ~new_P2_U3831 | ~new_P2_U5363 | ~new_P2_U5362;
  assign n3669 = ~new_P2_U3829 | ~new_P2_U5340 | ~new_P2_U5339;
  assign n3664 = ~new_P2_U3828 | ~new_P2_U5335 | ~new_P2_U5334;
  assign n3659 = ~new_P2_U3827 | ~new_P2_U5330 | ~new_P2_U5329;
  assign n3654 = ~new_P2_U3826 | ~new_P2_U5325 | ~new_P2_U5324;
  assign n3649 = ~new_P2_U3825 | ~new_P2_U5320 | ~new_P2_U5319;
  assign n3644 = ~new_P2_U3824 | ~new_P2_U5315 | ~new_P2_U5314;
  assign n3639 = ~new_P2_U3823 | ~new_P2_U5310 | ~new_P2_U5309;
  assign n3634 = ~new_P2_U3822 | ~new_P2_U5305 | ~new_P2_U5304;
  assign n3629 = ~new_P2_U3820 | ~new_P2_U5283 | ~new_P2_U5282;
  assign n3624 = ~new_P2_U3819 | ~new_P2_U5278 | ~new_P2_U5277;
  assign n3619 = ~new_P2_U3818 | ~new_P2_U5273 | ~new_P2_U5272;
  assign n3614 = ~new_P2_U3817 | ~new_P2_U5268 | ~new_P2_U5267;
  assign n3609 = ~new_P2_U3816 | ~new_P2_U5263 | ~new_P2_U5262;
  assign n3604 = ~new_P2_U3815 | ~new_P2_U5258 | ~new_P2_U5257;
  assign n3599 = ~new_P2_U3814 | ~new_P2_U5253 | ~new_P2_U5252;
  assign n3594 = ~new_P2_U3813 | ~new_P2_U5248 | ~new_P2_U5247;
  assign n3589 = ~new_P2_U3811 | ~new_P2_U5225 | ~new_P2_U5224;
  assign n3584 = ~new_P2_U3810 | ~new_P2_U5220 | ~new_P2_U5219;
  assign n3579 = ~new_P2_U3809 | ~new_P2_U5215 | ~new_P2_U5214;
  assign n3574 = ~new_P2_U3808 | ~new_P2_U5210 | ~new_P2_U5209;
  assign n3569 = ~new_P2_U3807 | ~new_P2_U5205 | ~new_P2_U5204;
  assign n3564 = ~new_P2_U3806 | ~new_P2_U5200 | ~new_P2_U5199;
  assign n3559 = ~new_P2_U3805 | ~new_P2_U5195 | ~new_P2_U5194;
  assign n3554 = ~new_P2_U3804 | ~new_P2_U5190 | ~new_P2_U5189;
  assign n3549 = ~new_P2_U3802 | ~new_P2_U5168 | ~new_P2_U5167;
  assign n3544 = ~new_P2_U3801 | ~new_P2_U5163 | ~new_P2_U5162;
  assign n3539 = ~new_P2_U3800 | ~new_P2_U5158 | ~new_P2_U5157;
  assign n3534 = ~new_P2_U3799 | ~new_P2_U5153 | ~new_P2_U5152;
  assign n3529 = ~new_P2_U3798 | ~new_P2_U5148 | ~new_P2_U5147;
  assign n3524 = ~new_P2_U3797 | ~new_P2_U5143 | ~new_P2_U5142;
  assign n3519 = ~new_P2_U3796 | ~new_P2_U5138 | ~new_P2_U5137;
  assign n3514 = ~new_P2_U3795 | ~new_P2_U5133 | ~new_P2_U5132;
  assign n3509 = ~new_P2_U3793 | ~new_P2_U5112 | ~new_P2_U5111;
  assign n3504 = ~new_P2_U3792 | ~new_P2_U5107 | ~new_P2_U5106;
  assign n3499 = ~new_P2_U3791 | ~new_P2_U5102 | ~new_P2_U5101;
  assign n3494 = ~new_P2_U3790 | ~new_P2_U5097 | ~new_P2_U5096;
  assign n3489 = ~new_P2_U3789 | ~new_P2_U5092 | ~new_P2_U5091;
  assign n3484 = ~new_P2_U3788 | ~new_P2_U5087 | ~new_P2_U5086;
  assign n3479 = ~new_P2_U3787 | ~new_P2_U5082 | ~new_P2_U5081;
  assign n3474 = ~new_P2_U3786 | ~new_P2_U5077 | ~new_P2_U5076;
  assign n3469 = ~new_P2_U3784 | ~new_P2_U5055 | ~new_P2_U5054;
  assign n3464 = ~new_P2_U3783 | ~new_P2_U5050 | ~new_P2_U5049;
  assign n3459 = ~new_P2_U3782 | ~new_P2_U5045 | ~new_P2_U5044;
  assign n3454 = ~new_P2_U3781 | ~new_P2_U5040 | ~new_P2_U5039;
  assign n3449 = ~new_P2_U3780 | ~new_P2_U5035 | ~new_P2_U5034;
  assign n3444 = ~new_P2_U3779 | ~new_P2_U5030 | ~new_P2_U5029;
  assign n3439 = ~new_P2_U3778 | ~new_P2_U5025 | ~new_P2_U5024;
  assign n3434 = ~new_P2_U3777 | ~new_P2_U5020 | ~new_P2_U5019;
  assign n3429 = ~new_P2_U3775 | ~new_P2_U4997 | ~new_P2_U4996;
  assign n3424 = ~new_P2_U3774 | ~new_P2_U4992 | ~new_P2_U4991;
  assign n3419 = ~new_P2_U3773 | ~new_P2_U4987 | ~new_P2_U4986;
  assign n3414 = ~new_P2_U3772 | ~new_P2_U4982 | ~new_P2_U4981;
  assign n3409 = ~new_P2_U3771 | ~new_P2_U4977 | ~new_P2_U4976;
  assign n3404 = ~new_P2_U3770 | ~new_P2_U4972 | ~new_P2_U4971;
  assign n3399 = ~new_P2_U3769 | ~new_P2_U4967 | ~new_P2_U4966;
  assign n3394 = ~new_P2_U3768 | ~new_P2_U4962 | ~new_P2_U4961;
  assign n3389 = ~new_P2_U3766 | ~new_P2_U4940 | ~new_P2_U4939;
  assign n3384 = ~new_P2_U3765 | ~new_P2_U4935 | ~new_P2_U4934;
  assign n3379 = ~new_P2_U3764 | ~new_P2_U4930 | ~new_P2_U4929;
  assign n3374 = ~new_P2_U3763 | ~new_P2_U4925 | ~new_P2_U4924;
  assign n3369 = ~new_P2_U3762 | ~new_P2_U4920 | ~new_P2_U4919;
  assign n3364 = ~new_P2_U3761 | ~new_P2_U4915 | ~new_P2_U4914;
  assign n3359 = ~new_P2_U3760 | ~new_P2_U4910 | ~new_P2_U4909;
  assign n3354 = ~new_P2_U3759 | ~new_P2_U4905 | ~new_P2_U4904;
  assign n3349 = ~new_P2_U3757 | ~new_P2_U4882 | ~new_P2_U4881;
  assign n3344 = ~new_P2_U3756 | ~new_P2_U4877 | ~new_P2_U4876;
  assign n3339 = ~new_P2_U3755 | ~new_P2_U4872 | ~new_P2_U4871;
  assign n3334 = ~new_P2_U3754 | ~new_P2_U4867 | ~new_P2_U4866;
  assign n3329 = ~new_P2_U3753 | ~new_P2_U4862 | ~new_P2_U4861;
  assign n3324 = ~new_P2_U3752 | ~new_P2_U4857 | ~new_P2_U4856;
  assign n3319 = ~new_P2_U3751 | ~new_P2_U4852 | ~new_P2_U4851;
  assign n3314 = ~new_P2_U3750 | ~new_P2_U4847 | ~new_P2_U4846;
  assign n3309 = ~new_P2_U3748 | ~new_P2_U4825 | ~new_P2_U4824;
  assign n3304 = ~new_P2_U3747 | ~new_P2_U4820 | ~new_P2_U4819;
  assign n3299 = ~new_P2_U3746 | ~new_P2_U4815 | ~new_P2_U4814;
  assign n3294 = ~new_P2_U3745 | ~new_P2_U4810 | ~new_P2_U4809;
  assign n3289 = ~new_P2_U3744 | ~new_P2_U4805 | ~new_P2_U4804;
  assign n3284 = ~new_P2_U3743 | ~new_P2_U4800 | ~new_P2_U4799;
  assign n3279 = ~new_P2_U3742 | ~new_P2_U4795 | ~new_P2_U4794;
  assign n3274 = ~new_P2_U3741 | ~new_P2_U4790 | ~new_P2_U4789;
  assign n3269 = ~new_P2_U3739 | ~new_P2_U4766 | ~new_P2_U4765;
  assign n3264 = ~new_P2_U3738 | ~new_P2_U4761 | ~new_P2_U4760;
  assign n3259 = ~new_P2_U3737 | ~new_P2_U4756 | ~new_P2_U4755;
  assign n3254 = ~new_P2_U3736 | ~new_P2_U4751 | ~new_P2_U4750;
  assign n3249 = ~new_P2_U3735 | ~new_P2_U4746 | ~new_P2_U4745;
  assign n3244 = ~new_P2_U3734 | ~new_P2_U4741 | ~new_P2_U4740;
  assign n3239 = ~new_P2_U3733 | ~new_P2_U4736 | ~new_P2_U4735;
  assign n3234 = ~new_P2_U3732 | ~new_P2_U4731 | ~new_P2_U4730;
  assign n3229 = ~new_P2_U3730 | ~new_P2_U4708 | ~new_P2_U4707;
  assign n3224 = ~new_P2_U3729 | ~new_P2_U4703 | ~new_P2_U4702;
  assign n3219 = ~new_P2_U3728 | ~new_P2_U4698 | ~new_P2_U4697;
  assign n3214 = ~new_P2_U3727 | ~new_P2_U4693 | ~new_P2_U4692;
  assign n3209 = ~new_P2_U3726 | ~new_P2_U4688 | ~new_P2_U4687;
  assign n3204 = ~new_P2_U3725 | ~new_P2_U4683 | ~new_P2_U4682;
  assign n3199 = ~new_P2_U3724 | ~new_P2_U4678 | ~new_P2_U4677;
  assign n3194 = ~new_P2_U3723 | ~new_P2_U4673 | ~new_P2_U4672;
  assign n3189 = ~new_P2_U3721 | ~new_P2_U8061 | ~new_P2_U8060;
  assign n3184 = ~new_P2_U4454 | ~new_P2_U4627 | ~new_P2_U4629 | ~new_P2_U4628;
  assign n3179 = ~new_P2_U3716 | ~new_P2_U4625;
  assign n3169 = P2_DATAWIDTH_REG_31_ & new_P2_U7917;
  assign n3164 = P2_DATAWIDTH_REG_30_ & new_P2_U7917;
  assign n3159 = P2_DATAWIDTH_REG_29_ & new_P2_U7917;
  assign n3154 = P2_DATAWIDTH_REG_28_ & new_P2_U7917;
  assign n3149 = P2_DATAWIDTH_REG_27_ & new_P2_U7917;
  assign n3144 = P2_DATAWIDTH_REG_26_ & new_P2_U7917;
  assign n3139 = P2_DATAWIDTH_REG_25_ & new_P2_U7917;
  assign n3134 = P2_DATAWIDTH_REG_24_ & new_P2_U7917;
  assign n3129 = P2_DATAWIDTH_REG_23_ & new_P2_U7917;
  assign n3124 = P2_DATAWIDTH_REG_22_ & new_P2_U7917;
  assign n3119 = P2_DATAWIDTH_REG_21_ & new_P2_U7917;
  assign n3114 = P2_DATAWIDTH_REG_20_ & new_P2_U7917;
  assign n3109 = P2_DATAWIDTH_REG_19_ & new_P2_U7917;
  assign n3104 = P2_DATAWIDTH_REG_18_ & new_P2_U7917;
  assign n3099 = P2_DATAWIDTH_REG_17_ & new_P2_U7917;
  assign n3094 = P2_DATAWIDTH_REG_16_ & new_P2_U7917;
  assign n3089 = P2_DATAWIDTH_REG_15_ & new_P2_U7917;
  assign n3084 = P2_DATAWIDTH_REG_14_ & new_P2_U7917;
  assign n3079 = P2_DATAWIDTH_REG_13_ & new_P2_U7917;
  assign n3074 = P2_DATAWIDTH_REG_12_ & new_P2_U7917;
  assign n3069 = P2_DATAWIDTH_REG_11_ & new_P2_U7917;
  assign n3064 = P2_DATAWIDTH_REG_10_ & new_P2_U7917;
  assign n3059 = P2_DATAWIDTH_REG_9_ & new_P2_U7917;
  assign n3054 = P2_DATAWIDTH_REG_8_ & new_P2_U7917;
  assign n3049 = P2_DATAWIDTH_REG_7_ & new_P2_U7917;
  assign n3044 = P2_DATAWIDTH_REG_6_ & new_P2_U7917;
  assign n3039 = P2_DATAWIDTH_REG_5_ & new_P2_U7917;
  assign n3034 = P2_DATAWIDTH_REG_4_ & new_P2_U7917;
  assign n3029 = P2_DATAWIDTH_REG_3_ & new_P2_U7917;
  assign n3024 = P2_DATAWIDTH_REG_2_ & new_P2_U7917;
  assign n3009 = ~new_P2_U4588 | ~new_P2_U7914 | ~new_P2_U7913;
  assign n3004 = ~new_P2_U3691 | ~new_P2_U7912 | ~new_P2_U7911;
  assign n2999 = ~new_P2_U3690 | ~new_P2_U4579;
  assign n2994 = ~new_P2_U4567 | ~new_P2_U4566 | ~new_P2_U4565;
  assign n2989 = ~new_P2_U4564 | ~new_P2_U4563 | ~new_P2_U4562;
  assign n2984 = ~new_P2_U4561 | ~new_P2_U4560 | ~new_P2_U4559;
  assign n2979 = ~new_P2_U4558 | ~new_P2_U4557 | ~new_P2_U4556;
  assign n2974 = ~new_P2_U4555 | ~new_P2_U4554 | ~new_P2_U4553;
  assign n2969 = ~new_P2_U4552 | ~new_P2_U4551 | ~new_P2_U4550;
  assign n2964 = ~new_P2_U4549 | ~new_P2_U4548 | ~new_P2_U4547;
  assign n2959 = ~new_P2_U4546 | ~new_P2_U4545 | ~new_P2_U4544;
  assign n2954 = ~new_P2_U4543 | ~new_P2_U4542 | ~new_P2_U4541;
  assign n2949 = ~new_P2_U4540 | ~new_P2_U4539 | ~new_P2_U4538;
  assign n2944 = ~new_P2_U4537 | ~new_P2_U4536 | ~new_P2_U4535;
  assign n2939 = ~new_P2_U4534 | ~new_P2_U4533 | ~new_P2_U4532;
  assign n2934 = ~new_P2_U4531 | ~new_P2_U4530 | ~new_P2_U4529;
  assign n2929 = ~new_P2_U4528 | ~new_P2_U4527 | ~new_P2_U4526;
  assign n2924 = ~new_P2_U4525 | ~new_P2_U4524 | ~new_P2_U4523;
  assign n2919 = ~new_P2_U4522 | ~new_P2_U4521 | ~new_P2_U4520;
  assign n2914 = ~new_P2_U4519 | ~new_P2_U4518 | ~new_P2_U4517;
  assign n2909 = ~new_P2_U4516 | ~new_P2_U4515 | ~new_P2_U4514;
  assign n2904 = ~new_P2_U4513 | ~new_P2_U4512 | ~new_P2_U4511;
  assign n2899 = ~new_P2_U4510 | ~new_P2_U4509 | ~new_P2_U4508;
  assign n2894 = ~new_P2_U4507 | ~new_P2_U4506 | ~new_P2_U4505;
  assign n2889 = ~new_P2_U4504 | ~new_P2_U4503 | ~new_P2_U4502;
  assign n2884 = ~new_P2_U4501 | ~new_P2_U4500 | ~new_P2_U4499;
  assign n2879 = ~new_P2_U4498 | ~new_P2_U4497 | ~new_P2_U4496;
  assign n2874 = ~new_P2_U4495 | ~new_P2_U4494 | ~new_P2_U4493;
  assign n2869 = ~new_P2_U4492 | ~new_P2_U4491 | ~new_P2_U4490;
  assign n2864 = ~new_P2_U4489 | ~new_P2_U4488 | ~new_P2_U4487;
  assign n2859 = ~new_P2_U4486 | ~new_P2_U4485 | ~new_P2_U4484;
  assign n2854 = ~new_P2_U4483 | ~new_P2_U4482 | ~new_P2_U4481;
  assign n2849 = ~new_P2_U4480 | ~new_P2_U4479 | ~new_P2_U4478;
  assign new_P2_U3242 = ~new_P2_U4191 | ~new_P2_U4192 | ~new_P2_U4194 | ~new_P2_U4193;
  assign new_P2_U3243 = ~new_P2_U3349 | ~new_P2_U3335;
  assign new_P2_U3244 = ~P2_STATE_REG_2_;
  assign new_P2_U3245 = ~new_P2_U2440 | ~new_P2_U3243;
  assign new_P2_U3246 = ~new_P2_U2440 | ~new_P2_U4650;
  assign new_P2_U3247 = ~new_P2_U2442 | ~new_P2_U3243;
  assign new_P2_U3248 = ~new_P2_U2442 | ~new_P2_U4650;
  assign new_P2_U3249 = ~new_P2_U2441 | ~new_P2_U3243;
  assign new_P2_U3250 = ~new_P2_U2441 | ~new_P2_U4650;
  assign new_P2_U3251 = ~new_P2_U2443 | ~new_P2_U3243;
  assign new_P2_U3252 = ~new_P2_U2443 | ~new_P2_U4650;
  assign new_P2_U3253 = ~new_P2_U3708 | ~new_P2_U3707;
  assign new_P2_U3254 = ~new_P2_U2590 | ~new_P2_U4429;
  assign new_P2_U3255 = ~new_P2_U3696 | ~new_P2_U3695;
  assign new_P2_U3256 = ~P2_REQUESTPENDING_REG;
  assign new_P2_U3257 = ~new_P2_U4608 | ~new_P2_U4609 | ~new_P2_U8051 | ~new_P2_U8050;
  assign new_P2_U3258 = ~P2_STATE_REG_1_;
  assign new_P2_U3259 = ~P2_STATE_REG_1_ | ~new_P2_U3266;
  assign new_P2_U3260 = ~new_P2_U4439 | ~new_P2_U3244;
  assign new_P2_U3261 = ~new_P2_U4439 | ~P2_STATE_REG_2_;
  assign new_P2_U3262 = ~P2_STATE_REG_1_ | ~new_P2_U3244;
  assign new_P2_U3263 = P2_STATE_REG_2_ | P2_STATE_REG_1_;
  assign new_P2_U3264 = ~HOLD;
  assign new_P2_U3265 = ~new_U211;
  assign new_P2_U3266 = ~P2_STATE_REG_0_;
  assign new_P2_U3267 = ~P2_REQUESTPENDING_REG | ~new_P2_U3264;
  assign new_P2_U3268 = HOLD | P2_REQUESTPENDING_REG;
  assign new_P2_U3269 = ~P2_STATE2_REG_1_;
  assign new_P2_U3270 = ~P2_STATE2_REG_2_;
  assign new_P2_U3271 = ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U3272 = ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_U3273 = ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign new_P2_U3274 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U3276;
  assign new_P2_U3275 = P2_INSTQUEUERD_ADDR_REG_2_ | P2_INSTQUEUERD_ADDR_REG_0_ | P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U3276 = ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign new_P2_U3277 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~P2_INSTQUEUERD_ADDR_REG_0_ | ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U3278 = ~new_P2_U3700 | ~new_P2_U3699;
  assign new_P2_U3279 = ~new_P2_U3702 | ~new_P2_U3701;
  assign new_P2_U3280 = ~new_P2_U3704 | ~new_P2_U3703;
  assign new_P2_U3281 = ~new_P2_U7859 | ~new_P2_U7861 | ~new_P2_U7863;
  assign new_P2_U3282 = ~new_P2_U4476 | ~new_P2_U2457 | ~new_P2_U7869;
  assign new_P2_U3283 = ~new_P2_U3253 | ~new_P2_U7873;
  assign new_P2_U3284 = ~P2_STATE2_REG_0_;
  assign new_P2_U3285 = ~new_P2_U4424 | ~new_P2_U3709;
  assign new_P2_U3286 = ~new_P2_U3253 | ~new_P2_U2616;
  assign new_P2_U3287 = ~new_P2_GTE_370_U6;
  assign new_P2_U3288 = ~new_P2_U2458 | ~new_P2_U2457 | ~new_P2_U7859;
  assign new_P2_U3289 = ~new_P2_U2616 | ~new_P2_U7871;
  assign new_P2_U3290 = ~new_P2_U4595 | ~new_P2_U3266;
  assign new_P2_U3291 = ~new_P2_U3713 | ~new_P2_U2459;
  assign new_P2_U3292 = ~new_P2_R2243_U8;
  assign new_P2_U3293 = ~new_P2_U2357 | ~new_P2_U3280;
  assign new_P2_U3294 = ~new_P2_U7871 | ~new_P2_U7873;
  assign new_P2_U3295 = ~new_P2_U7861 | ~new_P2_U2617;
  assign new_P2_U3296 = ~new_P2_U2451 | ~new_P2_U4428;
  assign new_P2_U3297 = ~new_P2_R2167_U6;
  assign new_P2_U3298 = ~new_P2_U4610 | ~new_P2_U4614 | ~new_P2_LT_563_U6 | ~new_P2_U7894 | ~new_P2_U4444;
  assign new_P2_U3299 = ~P2_STATE2_REG_0_ | ~new_P2_U4619;
  assign new_P2_U3300 = ~P2_STATE2_REG_3_;
  assign new_P2_U3301 = ~P2_STATE2_REG_0_ | ~new_P2_U3270;
  assign new_P2_U3302 = ~P2_STATEBS16_REG;
  assign new_P2_U3303 = P2_STATE2_REG_3_ | P2_STATE2_REG_1_;
  assign new_P2_U3304 = ~P2_STATE2_REG_2_ | ~new_P2_U3269;
  assign new_P2_U3305 = ~P2_STATE2_REG_3_ | ~new_P2_R2167_U6;
  assign new_P2_U3306 = ~new_P2_U4656 | ~new_P2_U3284;
  assign new_P2_U3307 = ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P2_U3308 = ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_U3309 = ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_U3310 = ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P2_U3311 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P2_U3312 = ~new_P2_U4642 | ~new_P2_U2464;
  assign new_P2_U3313 = P2_STATE2_REG_3_ | P2_STATE2_REG_2_;
  assign new_P2_U3314 = ~new_P2_R2182_U69;
  assign new_P2_U3315 = ~new_P2_R2182_U68;
  assign new_P2_U3316 = ~new_P2_R2182_U40;
  assign new_P2_U3317 = ~new_P2_R2182_U76;
  assign new_P2_U3318 = ~new_P2_R2182_U68 | ~new_P2_R2182_U69;
  assign new_P2_U3319 = ~new_P2_U3352 | ~new_P2_U3314;
  assign new_P2_U3320 = ~new_P2_U4636 | ~new_P2_U2461;
  assign new_P2_U3321 = ~new_P2_R2099_U95;
  assign new_P2_U3322 = ~new_P2_R2099_U96;
  assign new_P2_U3323 = ~new_P2_R2099_U94;
  assign new_P2_U3324 = ~new_P2_R2099_U5;
  assign new_P2_U3325 = ~new_P2_U3312 | ~new_P2_U4651;
  assign new_P2_U3326 = ~new_P2_U3570 | ~new_P2_U3312;
  assign new_P2_U3327 = ~P2_INSTQUEUE_REG_15__7_;
  assign new_P2_U3328 = ~P2_INSTQUEUE_REG_15__6_;
  assign new_P2_U3329 = ~P2_INSTQUEUE_REG_15__5_;
  assign new_P2_U3330 = ~P2_INSTQUEUE_REG_15__4_;
  assign new_P2_U3331 = ~P2_INSTQUEUE_REG_15__3_;
  assign new_P2_U3332 = ~P2_INSTQUEUE_REG_15__2_;
  assign new_P2_U3333 = ~P2_INSTQUEUE_REG_15__1_;
  assign new_P2_U3334 = ~P2_INSTQUEUE_REG_15__0_;
  assign new_P2_U3335 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_U3307;
  assign new_P2_U3336 = ~new_P2_U4649 | ~new_P2_U2464;
  assign new_P2_U3337 = ~new_P2_R2182_U68 | ~new_P2_U3314;
  assign new_P2_U3338 = ~new_P2_R2182_U69 | ~new_P2_U3352;
  assign new_P2_U3339 = ~new_P2_U4709 | ~new_P2_U2461;
  assign new_P2_U3340 = ~new_P2_U3569 | ~new_P2_U3336;
  assign new_P2_U3341 = ~P2_INSTQUEUE_REG_14__7_;
  assign new_P2_U3342 = ~P2_INSTQUEUE_REG_14__6_;
  assign new_P2_U3343 = ~P2_INSTQUEUE_REG_14__5_;
  assign new_P2_U3344 = ~P2_INSTQUEUE_REG_14__4_;
  assign new_P2_U3345 = ~P2_INSTQUEUE_REG_14__3_;
  assign new_P2_U3346 = ~P2_INSTQUEUE_REG_14__2_;
  assign new_P2_U3347 = ~P2_INSTQUEUE_REG_14__1_;
  assign new_P2_U3348 = ~P2_INSTQUEUE_REG_14__0_;
  assign new_P2_U3349 = ~P2_INSTQUEUEWR_ADDR_REG_0_ | ~new_P2_U3308;
  assign new_P2_U3350 = ~new_P2_U4648 | ~new_P2_U2464;
  assign new_P2_U3351 = ~new_P2_R2182_U69 | ~new_P2_U3315;
  assign new_P2_U3352 = ~new_P2_U3337 | ~new_P2_U3351;
  assign new_P2_U3353 = ~new_P2_U4635 | ~new_P2_U3314;
  assign new_P2_U3354 = ~new_P2_U4767 | ~new_P2_U2461;
  assign new_P2_U3355 = ~new_P2_U3350 | ~new_P2_U4770;
  assign new_P2_U3356 = ~new_P2_U3568 | ~new_P2_U3350;
  assign new_P2_U3357 = ~P2_INSTQUEUE_REG_13__7_;
  assign new_P2_U3358 = ~P2_INSTQUEUE_REG_13__6_;
  assign new_P2_U3359 = ~P2_INSTQUEUE_REG_13__5_;
  assign new_P2_U3360 = ~P2_INSTQUEUE_REG_13__4_;
  assign new_P2_U3361 = ~P2_INSTQUEUE_REG_13__3_;
  assign new_P2_U3362 = ~P2_INSTQUEUE_REG_13__2_;
  assign new_P2_U3363 = ~P2_INSTQUEUE_REG_13__1_;
  assign new_P2_U3364 = ~P2_INSTQUEUE_REG_13__0_;
  assign new_P2_U3365 = ~new_P2_U2478 | ~new_P2_U2464;
  assign new_P2_U3366 = ~new_P2_U2475 | ~new_P2_U2461;
  assign new_P2_U3367 = ~new_P2_U3567 | ~new_P2_U3365;
  assign new_P2_U3368 = ~P2_INSTQUEUE_REG_12__7_;
  assign new_P2_U3369 = ~P2_INSTQUEUE_REG_12__6_;
  assign new_P2_U3370 = ~P2_INSTQUEUE_REG_12__5_;
  assign new_P2_U3371 = ~P2_INSTQUEUE_REG_12__4_;
  assign new_P2_U3372 = ~P2_INSTQUEUE_REG_12__3_;
  assign new_P2_U3373 = ~P2_INSTQUEUE_REG_12__2_;
  assign new_P2_U3374 = ~P2_INSTQUEUE_REG_12__1_;
  assign new_P2_U3375 = ~P2_INSTQUEUE_REG_12__0_;
  assign new_P2_U3376 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_U3310;
  assign new_P2_U3377 = ~new_P2_U4645 | ~new_P2_U4642;
  assign new_P2_U3378 = ~new_P2_R2182_U76 | ~new_P2_U3316;
  assign new_P2_U3379 = ~new_P2_U2481 | ~new_P2_U4636;
  assign new_P2_U3380 = ~new_P2_U3377 | ~new_P2_U4885;
  assign new_P2_U3381 = ~new_P2_U3566 | ~new_P2_U3377;
  assign new_P2_U3382 = ~P2_INSTQUEUE_REG_11__7_;
  assign new_P2_U3383 = ~P2_INSTQUEUE_REG_11__6_;
  assign new_P2_U3384 = ~P2_INSTQUEUE_REG_11__5_;
  assign new_P2_U3385 = ~P2_INSTQUEUE_REG_11__4_;
  assign new_P2_U3386 = ~P2_INSTQUEUE_REG_11__3_;
  assign new_P2_U3387 = ~P2_INSTQUEUE_REG_11__2_;
  assign new_P2_U3388 = ~P2_INSTQUEUE_REG_11__1_;
  assign new_P2_U3389 = ~P2_INSTQUEUE_REG_11__0_;
  assign new_P2_U3390 = ~new_P2_U4645 | ~new_P2_U4649;
  assign new_P2_U3391 = ~new_P2_U2481 | ~new_P2_U4709;
  assign new_P2_U3392 = ~new_P2_U3565 | ~new_P2_U3390;
  assign new_P2_U3393 = ~P2_INSTQUEUE_REG_10__7_;
  assign new_P2_U3394 = ~P2_INSTQUEUE_REG_10__6_;
  assign new_P2_U3395 = ~P2_INSTQUEUE_REG_10__5_;
  assign new_P2_U3396 = ~P2_INSTQUEUE_REG_10__4_;
  assign new_P2_U3397 = ~P2_INSTQUEUE_REG_10__3_;
  assign new_P2_U3398 = ~P2_INSTQUEUE_REG_10__2_;
  assign new_P2_U3399 = ~P2_INSTQUEUE_REG_10__1_;
  assign new_P2_U3400 = ~P2_INSTQUEUE_REG_10__0_;
  assign new_P2_U3401 = ~new_P2_U4645 | ~new_P2_U4648;
  assign new_P2_U3402 = ~new_P2_U2481 | ~new_P2_U4767;
  assign new_P2_U3403 = ~new_P2_U3401 | ~new_P2_U5000;
  assign new_P2_U3404 = ~new_P2_U3564 | ~new_P2_U3401;
  assign new_P2_U3405 = ~P2_INSTQUEUE_REG_9__7_;
  assign new_P2_U3406 = ~P2_INSTQUEUE_REG_9__6_;
  assign new_P2_U3407 = ~P2_INSTQUEUE_REG_9__5_;
  assign new_P2_U3408 = ~P2_INSTQUEUE_REG_9__4_;
  assign new_P2_U3409 = ~P2_INSTQUEUE_REG_9__3_;
  assign new_P2_U3410 = ~P2_INSTQUEUE_REG_9__2_;
  assign new_P2_U3411 = ~P2_INSTQUEUE_REG_9__1_;
  assign new_P2_U3412 = ~P2_INSTQUEUE_REG_9__0_;
  assign new_P2_U3413 = ~new_P2_U4645 | ~new_P2_U2478;
  assign new_P2_U3414 = ~new_P2_U2481 | ~new_P2_U2475;
  assign new_P2_U3415 = ~new_P2_U3563 | ~new_P2_U3413;
  assign new_P2_U3416 = ~P2_INSTQUEUE_REG_8__7_;
  assign new_P2_U3417 = ~P2_INSTQUEUE_REG_8__6_;
  assign new_P2_U3418 = ~P2_INSTQUEUE_REG_8__5_;
  assign new_P2_U3419 = ~P2_INSTQUEUE_REG_8__4_;
  assign new_P2_U3420 = ~P2_INSTQUEUE_REG_8__3_;
  assign new_P2_U3421 = ~P2_INSTQUEUE_REG_8__2_;
  assign new_P2_U3422 = ~P2_INSTQUEUE_REG_8__1_;
  assign new_P2_U3423 = ~P2_INSTQUEUE_REG_8__0_;
  assign new_P2_U3424 = ~new_P2_U2465 | ~new_P2_U4642;
  assign new_P2_U3425 = ~new_P2_U2460 | ~new_P2_U4637;
  assign new_P2_U3426 = ~new_P2_U3425 | ~new_P2_U3378 | ~new_P2_U4639;
  assign new_P2_U3427 = ~new_P2_U2491 | ~new_P2_U4636;
  assign new_P2_U3428 = ~new_P2_U3424 | ~new_P2_U3376 | ~new_P2_U4646;
  assign new_P2_U3429 = ~new_P2_U3424 | ~new_P2_U5114;
  assign new_P2_U3430 = ~new_P2_U3562 | ~new_P2_U3424;
  assign new_P2_U3431 = ~P2_INSTQUEUE_REG_7__7_;
  assign new_P2_U3432 = ~P2_INSTQUEUE_REG_7__6_;
  assign new_P2_U3433 = ~P2_INSTQUEUE_REG_7__5_;
  assign new_P2_U3434 = ~P2_INSTQUEUE_REG_7__4_;
  assign new_P2_U3435 = ~P2_INSTQUEUE_REG_7__3_;
  assign new_P2_U3436 = ~P2_INSTQUEUE_REG_7__2_;
  assign new_P2_U3437 = ~P2_INSTQUEUE_REG_7__1_;
  assign new_P2_U3438 = ~P2_INSTQUEUE_REG_7__0_;
  assign new_P2_U3439 = ~new_P2_U4649 | ~new_P2_U2465;
  assign new_P2_U3440 = ~new_P2_U2491 | ~new_P2_U4709;
  assign new_P2_U3441 = ~new_P2_U3561 | ~new_P2_U3439;
  assign new_P2_U3442 = ~P2_INSTQUEUE_REG_6__7_;
  assign new_P2_U3443 = ~P2_INSTQUEUE_REG_6__6_;
  assign new_P2_U3444 = ~P2_INSTQUEUE_REG_6__5_;
  assign new_P2_U3445 = ~P2_INSTQUEUE_REG_6__4_;
  assign new_P2_U3446 = ~P2_INSTQUEUE_REG_6__3_;
  assign new_P2_U3447 = ~P2_INSTQUEUE_REG_6__2_;
  assign new_P2_U3448 = ~P2_INSTQUEUE_REG_6__1_;
  assign new_P2_U3449 = ~P2_INSTQUEUE_REG_6__0_;
  assign new_P2_U3450 = ~new_P2_U4648 | ~new_P2_U2465;
  assign new_P2_U3451 = ~new_P2_U2491 | ~new_P2_U4767;
  assign new_P2_U3452 = ~new_P2_U3450 | ~new_P2_U5228;
  assign new_P2_U3453 = ~new_P2_U3560 | ~new_P2_U3450;
  assign new_P2_U3454 = ~P2_INSTQUEUE_REG_5__7_;
  assign new_P2_U3455 = ~P2_INSTQUEUE_REG_5__6_;
  assign new_P2_U3456 = ~P2_INSTQUEUE_REG_5__5_;
  assign new_P2_U3457 = ~P2_INSTQUEUE_REG_5__4_;
  assign new_P2_U3458 = ~P2_INSTQUEUE_REG_5__3_;
  assign new_P2_U3459 = ~P2_INSTQUEUE_REG_5__2_;
  assign new_P2_U3460 = ~P2_INSTQUEUE_REG_5__1_;
  assign new_P2_U3461 = ~P2_INSTQUEUE_REG_5__0_;
  assign new_P2_U3462 = ~new_P2_U2478 | ~new_P2_U2465;
  assign new_P2_U3463 = ~new_P2_U2491 | ~new_P2_U2475;
  assign new_P2_U3464 = ~new_P2_U3559 | ~new_P2_U3462;
  assign new_P2_U3465 = ~P2_INSTQUEUE_REG_4__7_;
  assign new_P2_U3466 = ~P2_INSTQUEUE_REG_4__6_;
  assign new_P2_U3467 = ~P2_INSTQUEUE_REG_4__5_;
  assign new_P2_U3468 = ~P2_INSTQUEUE_REG_4__4_;
  assign new_P2_U3469 = ~P2_INSTQUEUE_REG_4__3_;
  assign new_P2_U3470 = ~P2_INSTQUEUE_REG_4__2_;
  assign new_P2_U3471 = ~P2_INSTQUEUE_REG_4__1_;
  assign new_P2_U3472 = ~P2_INSTQUEUE_REG_4__0_;
  assign new_P2_U3473 = ~new_P2_U2503 | ~new_P2_U4642;
  assign new_P2_U3474 = ~new_P2_U2500 | ~new_P2_U4636;
  assign new_P2_U3475 = ~new_P2_U3473 | ~new_P2_U5343;
  assign new_P2_U3476 = ~new_P2_U3558 | ~new_P2_U3473;
  assign new_P2_U3477 = ~P2_INSTQUEUE_REG_3__7_;
  assign new_P2_U3478 = ~P2_INSTQUEUE_REG_3__6_;
  assign new_P2_U3479 = ~P2_INSTQUEUE_REG_3__5_;
  assign new_P2_U3480 = ~P2_INSTQUEUE_REG_3__4_;
  assign new_P2_U3481 = ~P2_INSTQUEUE_REG_3__3_;
  assign new_P2_U3482 = ~P2_INSTQUEUE_REG_3__2_;
  assign new_P2_U3483 = ~P2_INSTQUEUE_REG_3__1_;
  assign new_P2_U3484 = ~P2_INSTQUEUE_REG_3__0_;
  assign new_P2_U3485 = ~new_P2_U2503 | ~new_P2_U4649;
  assign new_P2_U3486 = ~new_P2_U2500 | ~new_P2_U4709;
  assign new_P2_U3487 = ~new_P2_U3557 | ~new_P2_U3485;
  assign new_P2_U3488 = ~P2_INSTQUEUE_REG_2__7_;
  assign new_P2_U3489 = ~P2_INSTQUEUE_REG_2__6_;
  assign new_P2_U3490 = ~P2_INSTQUEUE_REG_2__5_;
  assign new_P2_U3491 = ~P2_INSTQUEUE_REG_2__4_;
  assign new_P2_U3492 = ~P2_INSTQUEUE_REG_2__3_;
  assign new_P2_U3493 = ~P2_INSTQUEUE_REG_2__2_;
  assign new_P2_U3494 = ~P2_INSTQUEUE_REG_2__1_;
  assign new_P2_U3495 = ~P2_INSTQUEUE_REG_2__0_;
  assign new_P2_U3496 = ~new_P2_U2503 | ~new_P2_U4648;
  assign new_P2_U3497 = ~new_P2_U2500 | ~new_P2_U4767;
  assign new_P2_U3498 = ~new_P2_U3496 | ~new_P2_U5458;
  assign new_P2_U3499 = ~new_P2_U3556 | ~new_P2_U3496;
  assign new_P2_U3500 = ~P2_INSTQUEUE_REG_1__7_;
  assign new_P2_U3501 = ~P2_INSTQUEUE_REG_1__6_;
  assign new_P2_U3502 = ~P2_INSTQUEUE_REG_1__5_;
  assign new_P2_U3503 = ~P2_INSTQUEUE_REG_1__4_;
  assign new_P2_U3504 = ~P2_INSTQUEUE_REG_1__3_;
  assign new_P2_U3505 = ~P2_INSTQUEUE_REG_1__2_;
  assign new_P2_U3506 = ~P2_INSTQUEUE_REG_1__1_;
  assign new_P2_U3507 = ~P2_INSTQUEUE_REG_1__0_;
  assign new_P2_U3508 = ~new_P2_U2503 | ~new_P2_U2478;
  assign new_P2_U3509 = ~new_P2_U2500 | ~new_P2_U2475;
  assign new_P2_U3510 = ~new_P2_U3555 | ~new_P2_U3508;
  assign new_P2_U3511 = ~P2_INSTQUEUE_REG_0__7_;
  assign new_P2_U3512 = ~P2_INSTQUEUE_REG_0__6_;
  assign new_P2_U3513 = ~P2_INSTQUEUE_REG_0__5_;
  assign new_P2_U3514 = ~P2_INSTQUEUE_REG_0__4_;
  assign new_P2_U3515 = ~P2_INSTQUEUE_REG_0__3_;
  assign new_P2_U3516 = ~P2_INSTQUEUE_REG_0__2_;
  assign new_P2_U3517 = ~P2_INSTQUEUE_REG_0__1_;
  assign new_P2_U3518 = ~P2_INSTQUEUE_REG_0__0_;
  assign new_P2_U3519 = ~P2_FLUSH_REG;
  assign new_P2_U3520 = ~new_P2_R2088_U6;
  assign new_P2_U3521 = ~new_P2_U3698 | ~new_P2_U3697;
  assign new_P2_U3522 = ~new_P2_U2451 | ~new_P2_U4429;
  assign new_P2_U3523 = ~new_P2_U4475 | ~new_P2_U4427;
  assign new_P2_U3524 = ~new_P2_U4429 | ~new_P2_U4475;
  assign new_P2_U3525 = ~new_P2_U7869 | ~new_P2_U3279 | ~new_P2_U7865 | ~new_P2_U7863;
  assign new_P2_U3526 = ~new_P2_R2147_U8;
  assign new_P2_U3527 = ~new_P2_U3283 | ~new_P2_U3289;
  assign new_P2_U3528 = ~new_P2_U3647;
  assign new_P2_U3529 = ~new_P2_R2147_U9;
  assign new_P2_U3530 = ~new_P2_U3274 | ~new_P2_U5615;
  assign new_P2_U3531 = ~new_P2_R2147_U4;
  assign new_P2_U3532 = ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_U3533 = ~new_P2_U5642 | ~new_P2_U4455 | ~new_P2_U3306;
  assign new_P2_U3534 = ~new_P2_U4430 | ~new_P2_U3269;
  assign new_P2_U3535 = ~new_P2_U5672 | ~new_P2_U5671;
  assign new_P2_U3536 = ~P2_STATE2_REG_0_ | ~new_P2_U7873;
  assign new_P2_U3537 = ~new_P2_U5937 | ~new_P2_U5936;
  assign new_P2_U3538 = ~new_P2_U4055 | ~new_P2_U2446;
  assign new_P2_U3539 = ~new_P2_U4056 | ~new_P2_U2357;
  assign new_P2_U3540 = ~P2_STATE2_REG_2_ | ~new_P2_U3284;
  assign new_P2_U3541 = ~new_P2_U6231 | ~new_P2_U6230;
  assign new_P2_U3542 = ~new_P2_U2374 | ~new_P2_U6326;
  assign new_P2_U3543 = ~new_P2_U2374 | ~new_P2_U6470;
  assign new_P2_U3544 = ~P2_EBX_REG_31_;
  assign new_P2_U3545 = P2_STATEBS16_REG | new_U211;
  assign new_P2_U3546 = ~new_P2_U4069 | ~new_P2_U4462;
  assign new_P2_U3547 = ~new_P2_U4171 | ~new_P2_U4174 | ~new_P2_U4181 | ~new_P2_U4177;
  assign new_P2_U3548 = ~new_P2_U4438 | ~P2_REIP_REG_1_;
  assign new_P2_U3549 = ~new_P2_U2356 | ~new_P2_U4420;
  assign new_P2_U3550 = ~new_P2_U4427 | ~P2_STATE2_REG_0_;
  assign new_P2_U3551 = ~P2_CODEFETCH_REG;
  assign new_P2_U3552 = ~P2_READREQUEST_REG;
  assign new_P2_U3553 = ~new_P2_U4405 | ~new_P2_U3275;
  assign new_P2_U3554 = ~new_P2_U4415 | ~new_P2_U3576;
  assign new_P2_U3555 = ~new_P2_U2504 | ~new_P2_U2479;
  assign new_P2_U3556 = ~new_P2_U2504 | ~new_P2_U2473;
  assign new_P2_U3557 = ~new_P2_U2504 | ~new_P2_U2470;
  assign new_P2_U3558 = ~new_P2_U2504 | ~new_P2_U2467;
  assign new_P2_U3559 = ~new_P2_U2492 | ~new_P2_U2479;
  assign new_P2_U3560 = ~new_P2_U2492 | ~new_P2_U2473;
  assign new_P2_U3561 = ~new_P2_U2492 | ~new_P2_U2470;
  assign new_P2_U3562 = ~new_P2_U2492 | ~new_P2_U2467;
  assign new_P2_U3563 = ~new_P2_U2483 | ~new_P2_U2479;
  assign new_P2_U3564 = ~new_P2_U2483 | ~new_P2_U2473;
  assign new_P2_U3565 = ~new_P2_U2483 | ~new_P2_U2470;
  assign new_P2_U3566 = ~new_P2_U2483 | ~new_P2_U2467;
  assign new_P2_U3567 = ~new_P2_U2479 | ~new_P2_U2466;
  assign new_P2_U3568 = ~new_P2_U2473 | ~new_P2_U2466;
  assign new_P2_U3569 = ~new_P2_U2470 | ~new_P2_U2466;
  assign new_P2_U3570 = ~new_P2_U2466 | ~new_P2_U2467;
  assign new_P2_U3571 = ~new_P2_U7865 | ~new_P2_U3300;
  assign new_P2_U3572 = ~new_P2_U3242;
  assign new_P2_U3573 = P2_STATE2_REG_0_ | P2_STATE2_REG_1_;
  assign new_P2_U3574 = ~new_P2_U3521 | ~new_P2_U5571 | ~new_P2_U3295;
  assign new_P2_U3575 = ~new_P2_U4419 | ~new_P2_U7871;
  assign new_P2_U3576 = ~new_P2_U4419 | ~new_P2_U3279;
  assign new_P2_U3577 = ~new_P2_U4424 | ~new_P2_U6845;
  assign new_P2_U3578 = ~new_P2_U2590 | ~new_P2_U4428;
  assign new_P2_U3579 = ~new_P2_U8063 | ~new_P2_U8062;
  assign new_P2_U3580 = ~new_P2_U8066 | ~new_P2_U8065;
  assign new_P2_U3581 = ~new_P2_U8081 | ~new_P2_U8080;
  assign new_P2_U3582 = ~new_P2_U8099 | ~new_P2_U8098;
  assign new_P2_U3583 = ~new_P2_U8148 | ~new_P2_U8147;
  assign new_P2_U3584 = ~new_P2_U8151 | ~new_P2_U8150;
  assign n2829 = ~new_P2_U7900 | ~new_P2_U7899;
  assign n2834 = ~new_P2_U7902 | ~new_P2_U7901;
  assign n2839 = ~new_P2_U7904 | ~new_P2_U7903;
  assign n2844 = ~new_P2_U7906 | ~new_P2_U7905;
  assign new_P2_U3589 = ~new_P2_U7916 | ~new_P2_U7915;
  assign new_P2_U3590 = new_P2_U3263 & new_P2_U4401;
  assign n3014 = ~new_P2_U7919 | ~new_P2_U7918;
  assign n3019 = ~new_P2_U7921 | ~new_P2_U7920;
  assign n3174 = ~new_P2_U8059 | ~new_P2_U8058;
  assign new_P2_U3594 = new_P2_U3866 & new_P2_U4434;
  assign n3834 = ~new_P2_U8073 | ~new_P2_U8072;
  assign n3839 = ~new_P2_U8084 | ~new_P2_U8083;
  assign new_P2_U3597 = ~new_P2_U8086 | ~new_P2_U8085;
  assign new_P2_U3598 = ~new_P2_U8089 | ~new_P2_U8088;
  assign n3844 = ~new_P2_U8094 | ~new_P2_U8093;
  assign n3849 = ~new_P2_U8102 | ~new_P2_U8101;
  assign n3854 = ~new_P2_U8104 | ~new_P2_U8103;
  assign n3864 = ~new_P2_U8106 | ~new_P2_U8105;
  assign n3869 = ~new_P2_U8111 | ~new_P2_U8110;
  assign n3874 = ~new_P2_U8113 | ~new_P2_U8112;
  assign n3879 = ~new_P2_U8115 | ~new_P2_U8114;
  assign new_P2_U3606 = ~P2_REIP_REG_1_ & ~P2_DATAWIDTH_REG_1_;
  assign new_P2_U3607 = new_P2_U4183 & new_P2_U7898;
  assign n5019 = ~new_P2_U8130 | ~new_P2_U8129;
  assign n5029 = ~new_P2_U8134 | ~new_P2_U8133;
  assign n5039 = ~new_P2_U8138 | ~new_P2_U8137;
  assign n5049 = ~new_P2_U8142 | ~new_P2_U8141;
  assign n5064 = ~new_P2_U8144 | ~new_P2_U8143;
  assign new_P2_U3613 = ~new_P2_U8282 | ~new_P2_U8281;
  assign new_P2_U3614 = ~new_P2_U8284 | ~new_P2_U8283;
  assign new_P2_U3615 = ~new_P2_U8286 | ~new_P2_U8285;
  assign new_P2_U3616 = new_P2_U4434 & new_P2_R2147_U7;
  assign new_P2_U3617 = ~new_P2_U8288 | ~new_P2_U8287;
  assign new_P2_U3618 = ~new_P2_U8290 | ~new_P2_U8289;
  assign new_P2_U3619 = ~new_P2_U8292 | ~new_P2_U8291;
  assign new_P2_U3620 = ~new_P2_U8294 | ~new_P2_U8293;
  assign new_P2_U3621 = ~new_P2_U8296 | ~new_P2_U8295;
  assign new_P2_U3622 = ~new_P2_U8298 | ~new_P2_U8297;
  assign new_P2_U3623 = ~new_P2_U8300 | ~new_P2_U8299;
  assign new_P2_U3624 = ~new_P2_U8302 | ~new_P2_U8301;
  assign new_P2_U3625 = ~new_P2_U8304 | ~new_P2_U8303;
  assign new_P2_U3626 = ~new_P2_U8306 | ~new_P2_U8305;
  assign new_P2_U3627 = ~new_P2_U8308 | ~new_P2_U8307;
  assign new_P2_U3628 = ~new_P2_U8310 | ~new_P2_U8309;
  assign new_P2_U3629 = ~new_P2_U8312 | ~new_P2_U8311;
  assign new_P2_U3630 = ~new_P2_U8314 | ~new_P2_U8313;
  assign new_P2_U3631 = ~new_P2_U8316 | ~new_P2_U8315;
  assign new_P2_U3632 = ~new_P2_U8318 | ~new_P2_U8317;
  assign new_P2_U3633 = ~new_P2_U8320 | ~new_P2_U8319;
  assign new_P2_U3634 = ~new_P2_U8322 | ~new_P2_U8321;
  assign new_P2_U3635 = ~new_P2_U8324 | ~new_P2_U8323;
  assign new_P2_U3636 = ~new_P2_U8326 | ~new_P2_U8325;
  assign new_P2_U3637 = ~new_P2_U8328 | ~new_P2_U8327;
  assign new_P2_U3638 = ~new_P2_U8330 | ~new_P2_U8329;
  assign new_P2_U3639 = ~new_P2_U8332 | ~new_P2_U8331;
  assign new_P2_U3640 = ~new_P2_U8334 | ~new_P2_U8333;
  assign new_P2_U3641 = ~new_P2_U8336 | ~new_P2_U8335;
  assign new_P2_U3642 = ~new_P2_U8338 | ~new_P2_U8337;
  assign new_P2_U3643 = ~new_P2_U8340 | ~new_P2_U8339;
  assign new_P2_U3644 = ~new_P2_U8342 | ~new_P2_U8341;
  assign new_P2_U3645 = ~new_P2_U8344 | ~new_P2_U8343;
  assign new_P2_U3646 = ~new_P2_U8346 | ~new_P2_U8345;
  assign new_P2_U3647 = ~new_P2_U8350 | ~new_P2_U8349;
  assign new_P2_U3648 = ~new_P2_U8352 | ~new_P2_U8351;
  assign new_P2_U3649 = ~new_P2_U8354 | ~new_P2_U8353;
  assign new_P2_U3650 = ~new_P2_U8356 | ~new_P2_U8355;
  assign new_P2_U3651 = ~new_P2_U8358 | ~new_P2_U8357;
  assign new_P2_U3652 = ~new_P2_U8360 | ~new_P2_U8359;
  assign new_P2_U3653 = ~new_P2_U8362 | ~new_P2_U8361;
  assign new_P2_U3654 = ~new_P2_U8364 | ~new_P2_U8363;
  assign new_P2_U3655 = ~new_P2_U8366 | ~new_P2_U8365;
  assign new_P2_U3656 = ~new_P2_U8368 | ~new_P2_U8367;
  assign new_P2_U3657 = ~new_P2_U8370 | ~new_P2_U8369;
  assign new_P2_U3658 = ~new_P2_U8372 | ~new_P2_U8371;
  assign new_P2_U3659 = ~new_P2_U8374 | ~new_P2_U8373;
  assign new_P2_U3660 = ~new_P2_U8376 | ~new_P2_U8375;
  assign new_P2_U3661 = ~new_P2_U8378 | ~new_P2_U8377;
  assign new_P2_U3662 = ~new_P2_U8380 | ~new_P2_U8379;
  assign new_P2_U3663 = ~new_P2_U8382 | ~new_P2_U8381;
  assign new_P2_U3664 = ~new_P2_U8384 | ~new_P2_U8383;
  assign new_P2_U3665 = ~new_P2_U8386 | ~new_P2_U8385;
  assign new_P2_U3666 = ~new_P2_U8388 | ~new_P2_U8387;
  assign new_P2_U3667 = ~new_P2_U8390 | ~new_P2_U8389;
  assign new_P2_U3668 = ~new_P2_U8392 | ~new_P2_U8391;
  assign new_P2_U3669 = ~new_P2_U8394 | ~new_P2_U8393;
  assign new_P2_U3670 = ~new_P2_U8396 | ~new_P2_U8395;
  assign new_P2_U3671 = ~new_P2_U8398 | ~new_P2_U8397;
  assign new_P2_U3672 = ~new_P2_U8400 | ~new_P2_U8399;
  assign new_P2_U3673 = ~new_P2_U8402 | ~new_P2_U8401;
  assign new_P2_U3674 = ~new_P2_U8404 | ~new_P2_U8403;
  assign new_P2_U3675 = ~new_P2_U8406 | ~new_P2_U8405;
  assign new_P2_U3676 = ~new_P2_U8408 | ~new_P2_U8407;
  assign new_P2_U3677 = ~new_P2_U8410 | ~new_P2_U8409;
  assign new_P2_U3678 = ~new_P2_U8412 | ~new_P2_U8411;
  assign new_P2_U3679 = ~new_P2_U8414 | ~new_P2_U8413;
  assign new_P2_U3680 = ~new_P2_U8416 | ~new_P2_U8415;
  assign new_P2_U3681 = ~new_P2_U8418 | ~new_P2_U8417;
  assign new_P2_U3682 = ~new_P2_U8420 | ~new_P2_U8419;
  assign new_P2_U3683 = ~new_P2_U8422 | ~new_P2_U8421;
  assign new_P2_U3684 = ~new_P2_U8424 | ~new_P2_U8423;
  assign new_P2_U3685 = ~new_P2_U8426 | ~new_P2_U8425;
  assign new_P2_U3686 = ~new_P2_U8428 | ~new_P2_U8427;
  assign new_P2_U3687 = ~new_P2_U8430 | ~new_P2_U8429;
  assign new_P2_U3688 = ~new_P2_U8432 | ~new_P2_U8431;
  assign new_P2_U3689 = ~new_P2_U8434 | ~new_P2_U8433;
  assign new_P2_U3690 = new_P2_U4578 & new_P2_U3261;
  assign new_P2_U3691 = new_P2_U4583 & new_P2_U3260;
  assign new_P2_U3692 = P2_REQUESTPENDING_REG & P2_STATE_REG_0_;
  assign new_P2_U3693 = new_P2_U7751 & new_P2_U7767 & new_P2_U7799 & new_P2_U7783;
  assign new_P2_U3694 = new_P2_U7815 & new_P2_U7831 & new_P2_U7868 & new_P2_U7847;
  assign new_P2_U3695 = new_P2_U7750 & new_P2_U7766 & new_P2_U7798 & new_P2_U7782;
  assign new_P2_U3696 = new_P2_U7814 & new_P2_U7830 & new_P2_U7866 & new_P2_U7846;
  assign new_P2_U3697 = new_P2_U7749 & new_P2_U7765 & new_P2_U7797 & new_P2_U7781;
  assign new_P2_U3698 = new_P2_U7813 & new_P2_U7829 & new_P2_U7864 & new_P2_U7845;
  assign new_P2_U3699 = new_P2_U7748 & new_P2_U7764 & new_P2_U7796 & new_P2_U7780;
  assign new_P2_U3700 = new_P2_U7812 & new_P2_U7828 & new_P2_U7862 & new_P2_U7844;
  assign new_P2_U3701 = new_P2_U7747 & new_P2_U7763 & new_P2_U7795 & new_P2_U7779;
  assign new_P2_U3702 = new_P2_U7811 & new_P2_U7827 & new_P2_U7860 & new_P2_U7843;
  assign new_P2_U3703 = new_P2_U7746 & new_P2_U7762 & new_P2_U7794 & new_P2_U7778;
  assign new_P2_U3704 = new_P2_U7810 & new_P2_U7826 & new_P2_U7858 & new_P2_U7842;
  assign new_P2_U3705 = new_P2_U7753 & new_P2_U7769 & new_P2_U7801 & new_P2_U7785;
  assign new_P2_U3706 = new_P2_U7817 & new_P2_U7833 & new_P2_U7872 & new_P2_U7849;
  assign new_P2_U3707 = new_P2_U7752 & new_P2_U7768 & new_P2_U7800 & new_P2_U7784;
  assign new_P2_U3708 = new_P2_U7816 & new_P2_U7832 & new_P2_U7870 & new_P2_U7848;
  assign new_P2_U3709 = new_P2_U3710 & new_P2_U4417;
  assign new_P2_U3710 = P2_STATE2_REG_0_ & new_P2_U4595;
  assign new_P2_U3711 = new_P2_U2360 & new_P2_U3266;
  assign new_P2_U3712 = new_P2_U3521 & new_P2_U7867;
  assign new_P2_U3713 = new_P2_U4599 & new_P2_U4598;
  assign new_P2_U3714 = P2_STATE2_REG_2_ & new_P2_U3573;
  assign new_P2_U3715 = new_P2_U3714 & new_P2_U4618;
  assign new_P2_U3716 = new_P2_U4624 & new_P2_U3304;
  assign new_P2_U3717 = new_P2_U4466 & new_P2_U3265;
  assign new_P2_U3718 = P2_STATE2_REG_3_ & new_P2_U3269;
  assign new_P2_U3719 = ~P2_STATE2_REG_2_ & ~P2_STATE2_REG_1_;
  assign new_P2_U3720 = new_P2_U4465 & new_P2_U4453;
  assign new_P2_U3721 = new_P2_U3720 & new_P2_U4632;
  assign new_P2_U3722 = new_P2_U4443 & new_P2_U4661 & new_P2_U4662;
  assign new_P2_U3723 = new_P2_U4671 & new_P2_U4670 & new_P2_U4669;
  assign new_P2_U3724 = new_P2_U4676 & new_P2_U4675 & new_P2_U4674;
  assign new_P2_U3725 = new_P2_U4681 & new_P2_U4680 & new_P2_U4679;
  assign new_P2_U3726 = new_P2_U4686 & new_P2_U4685 & new_P2_U4684;
  assign new_P2_U3727 = new_P2_U4691 & new_P2_U4690 & new_P2_U4689;
  assign new_P2_U3728 = new_P2_U4696 & new_P2_U4695 & new_P2_U4694;
  assign new_P2_U3729 = new_P2_U4701 & new_P2_U4700 & new_P2_U4699;
  assign new_P2_U3730 = new_P2_U4706 & new_P2_U4705 & new_P2_U4704;
  assign new_P2_U3731 = new_P2_U4443 & new_P2_U4719 & new_P2_U4720;
  assign new_P2_U3732 = new_P2_U4729 & new_P2_U4728 & new_P2_U4727;
  assign new_P2_U3733 = new_P2_U4734 & new_P2_U4733 & new_P2_U4732;
  assign new_P2_U3734 = new_P2_U4739 & new_P2_U4738 & new_P2_U4737;
  assign new_P2_U3735 = new_P2_U4744 & new_P2_U4743 & new_P2_U4742;
  assign new_P2_U3736 = new_P2_U4749 & new_P2_U4748 & new_P2_U4747;
  assign new_P2_U3737 = new_P2_U4754 & new_P2_U4753 & new_P2_U4752;
  assign new_P2_U3738 = new_P2_U4759 & new_P2_U4758 & new_P2_U4757;
  assign new_P2_U3739 = new_P2_U4764 & new_P2_U4763 & new_P2_U4762;
  assign new_P2_U3740 = new_P2_U4443 & new_P2_U4778 & new_P2_U4779;
  assign new_P2_U3741 = new_P2_U4788 & new_P2_U4787 & new_P2_U4786;
  assign new_P2_U3742 = new_P2_U4793 & new_P2_U4792 & new_P2_U4791;
  assign new_P2_U3743 = new_P2_U4798 & new_P2_U4797 & new_P2_U4796;
  assign new_P2_U3744 = new_P2_U4803 & new_P2_U4802 & new_P2_U4801;
  assign new_P2_U3745 = new_P2_U4808 & new_P2_U4807 & new_P2_U4806;
  assign new_P2_U3746 = new_P2_U4813 & new_P2_U4812 & new_P2_U4811;
  assign new_P2_U3747 = new_P2_U4818 & new_P2_U4817 & new_P2_U4816;
  assign new_P2_U3748 = new_P2_U4823 & new_P2_U4822 & new_P2_U4821;
  assign new_P2_U3749 = new_P2_U4443 & new_P2_U4835 & new_P2_U4836;
  assign new_P2_U3750 = new_P2_U4845 & new_P2_U4844 & new_P2_U4843;
  assign new_P2_U3751 = new_P2_U4850 & new_P2_U4849 & new_P2_U4848;
  assign new_P2_U3752 = new_P2_U4855 & new_P2_U4854 & new_P2_U4853;
  assign new_P2_U3753 = new_P2_U4860 & new_P2_U4859 & new_P2_U4858;
  assign new_P2_U3754 = new_P2_U4865 & new_P2_U4864 & new_P2_U4863;
  assign new_P2_U3755 = new_P2_U4870 & new_P2_U4869 & new_P2_U4868;
  assign new_P2_U3756 = new_P2_U4875 & new_P2_U4874 & new_P2_U4873;
  assign new_P2_U3757 = new_P2_U4880 & new_P2_U4879 & new_P2_U4878;
  assign new_P2_U3758 = new_P2_U4443 & new_P2_U4893 & new_P2_U4894;
  assign new_P2_U3759 = new_P2_U4903 & new_P2_U4902 & new_P2_U4901;
  assign new_P2_U3760 = new_P2_U4908 & new_P2_U4907 & new_P2_U4906;
  assign new_P2_U3761 = new_P2_U4913 & new_P2_U4912 & new_P2_U4911;
  assign new_P2_U3762 = new_P2_U4918 & new_P2_U4917 & new_P2_U4916;
  assign new_P2_U3763 = new_P2_U4923 & new_P2_U4922 & new_P2_U4921;
  assign new_P2_U3764 = new_P2_U4928 & new_P2_U4927 & new_P2_U4926;
  assign new_P2_U3765 = new_P2_U4933 & new_P2_U4932 & new_P2_U4931;
  assign new_P2_U3766 = new_P2_U4938 & new_P2_U4937 & new_P2_U4936;
  assign new_P2_U3767 = new_P2_U4443 & new_P2_U4950 & new_P2_U4951;
  assign new_P2_U3768 = new_P2_U4960 & new_P2_U4959 & new_P2_U4958;
  assign new_P2_U3769 = new_P2_U4965 & new_P2_U4964 & new_P2_U4963;
  assign new_P2_U3770 = new_P2_U4970 & new_P2_U4969 & new_P2_U4968;
  assign new_P2_U3771 = new_P2_U4975 & new_P2_U4974 & new_P2_U4973;
  assign new_P2_U3772 = new_P2_U4980 & new_P2_U4979 & new_P2_U4978;
  assign new_P2_U3773 = new_P2_U4985 & new_P2_U4984 & new_P2_U4983;
  assign new_P2_U3774 = new_P2_U4990 & new_P2_U4989 & new_P2_U4988;
  assign new_P2_U3775 = new_P2_U4995 & new_P2_U4994 & new_P2_U4993;
  assign new_P2_U3776 = new_P2_U4443 & new_P2_U5008 & new_P2_U5009;
  assign new_P2_U3777 = new_P2_U5018 & new_P2_U5017 & new_P2_U5016;
  assign new_P2_U3778 = new_P2_U5023 & new_P2_U5022 & new_P2_U5021;
  assign new_P2_U3779 = new_P2_U5028 & new_P2_U5027 & new_P2_U5026;
  assign new_P2_U3780 = new_P2_U5033 & new_P2_U5032 & new_P2_U5031;
  assign new_P2_U3781 = new_P2_U5038 & new_P2_U5037 & new_P2_U5036;
  assign new_P2_U3782 = new_P2_U5043 & new_P2_U5042 & new_P2_U5041;
  assign new_P2_U3783 = new_P2_U5048 & new_P2_U5047 & new_P2_U5046;
  assign new_P2_U3784 = new_P2_U5053 & new_P2_U5052 & new_P2_U5051;
  assign new_P2_U3785 = new_P2_U4443 & new_P2_U5065 & new_P2_U5066;
  assign new_P2_U3786 = new_P2_U5075 & new_P2_U5074 & new_P2_U5073;
  assign new_P2_U3787 = new_P2_U5080 & new_P2_U5079 & new_P2_U5078;
  assign new_P2_U3788 = new_P2_U5085 & new_P2_U5084 & new_P2_U5083;
  assign new_P2_U3789 = new_P2_U5090 & new_P2_U5089 & new_P2_U5088;
  assign new_P2_U3790 = new_P2_U5095 & new_P2_U5094 & new_P2_U5093;
  assign new_P2_U3791 = new_P2_U5100 & new_P2_U5099 & new_P2_U5098;
  assign new_P2_U3792 = new_P2_U5105 & new_P2_U5104 & new_P2_U5103;
  assign new_P2_U3793 = new_P2_U5110 & new_P2_U5109 & new_P2_U5108;
  assign new_P2_U3794 = new_P2_U4443 & new_P2_U5121 & new_P2_U5122;
  assign new_P2_U3795 = new_P2_U5131 & new_P2_U5130 & new_P2_U5129;
  assign new_P2_U3796 = new_P2_U5136 & new_P2_U5135 & new_P2_U5134;
  assign new_P2_U3797 = new_P2_U5141 & new_P2_U5140 & new_P2_U5139;
  assign new_P2_U3798 = new_P2_U5146 & new_P2_U5145 & new_P2_U5144;
  assign new_P2_U3799 = new_P2_U5151 & new_P2_U5150 & new_P2_U5149;
  assign new_P2_U3800 = new_P2_U5156 & new_P2_U5155 & new_P2_U5154;
  assign new_P2_U3801 = new_P2_U5161 & new_P2_U5160 & new_P2_U5159;
  assign new_P2_U3802 = new_P2_U5166 & new_P2_U5165 & new_P2_U5164;
  assign new_P2_U3803 = new_P2_U4443 & new_P2_U5178 & new_P2_U5179;
  assign new_P2_U3804 = new_P2_U5188 & new_P2_U5187 & new_P2_U5186;
  assign new_P2_U3805 = new_P2_U5193 & new_P2_U5192 & new_P2_U5191;
  assign new_P2_U3806 = new_P2_U5198 & new_P2_U5197 & new_P2_U5196;
  assign new_P2_U3807 = new_P2_U5203 & new_P2_U5202 & new_P2_U5201;
  assign new_P2_U3808 = new_P2_U5208 & new_P2_U5207 & new_P2_U5206;
  assign new_P2_U3809 = new_P2_U5213 & new_P2_U5212 & new_P2_U5211;
  assign new_P2_U3810 = new_P2_U5218 & new_P2_U5217 & new_P2_U5216;
  assign new_P2_U3811 = new_P2_U5223 & new_P2_U5222 & new_P2_U5221;
  assign new_P2_U3812 = new_P2_U4443 & new_P2_U5236 & new_P2_U5237;
  assign new_P2_U3813 = new_P2_U5246 & new_P2_U5245 & new_P2_U5244;
  assign new_P2_U3814 = new_P2_U5251 & new_P2_U5250 & new_P2_U5249;
  assign new_P2_U3815 = new_P2_U5256 & new_P2_U5255 & new_P2_U5254;
  assign new_P2_U3816 = new_P2_U5261 & new_P2_U5260 & new_P2_U5259;
  assign new_P2_U3817 = new_P2_U5266 & new_P2_U5265 & new_P2_U5264;
  assign new_P2_U3818 = new_P2_U5271 & new_P2_U5270 & new_P2_U5269;
  assign new_P2_U3819 = new_P2_U5276 & new_P2_U5275 & new_P2_U5274;
  assign new_P2_U3820 = new_P2_U5281 & new_P2_U5280 & new_P2_U5279;
  assign new_P2_U3821 = new_P2_U4443 & new_P2_U5293 & new_P2_U5294;
  assign new_P2_U3822 = new_P2_U5303 & new_P2_U5302 & new_P2_U5301;
  assign new_P2_U3823 = new_P2_U5308 & new_P2_U5307 & new_P2_U5306;
  assign new_P2_U3824 = new_P2_U5313 & new_P2_U5312 & new_P2_U5311;
  assign new_P2_U3825 = new_P2_U5318 & new_P2_U5317 & new_P2_U5316;
  assign new_P2_U3826 = new_P2_U5323 & new_P2_U5322 & new_P2_U5321;
  assign new_P2_U3827 = new_P2_U5328 & new_P2_U5327 & new_P2_U5326;
  assign new_P2_U3828 = new_P2_U5333 & new_P2_U5332 & new_P2_U5331;
  assign new_P2_U3829 = new_P2_U5338 & new_P2_U5337 & new_P2_U5336;
  assign new_P2_U3830 = new_P2_U4443 & new_P2_U5351 & new_P2_U5352;
  assign new_P2_U3831 = new_P2_U5361 & new_P2_U5360 & new_P2_U5359;
  assign new_P2_U3832 = new_P2_U5366 & new_P2_U5365 & new_P2_U5364;
  assign new_P2_U3833 = new_P2_U5371 & new_P2_U5370 & new_P2_U5369;
  assign new_P2_U3834 = new_P2_U5376 & new_P2_U5375 & new_P2_U5374;
  assign new_P2_U3835 = new_P2_U5381 & new_P2_U5380 & new_P2_U5379;
  assign new_P2_U3836 = new_P2_U5386 & new_P2_U5385 & new_P2_U5384;
  assign new_P2_U3837 = new_P2_U5391 & new_P2_U5390 & new_P2_U5389;
  assign new_P2_U3838 = new_P2_U5396 & new_P2_U5395 & new_P2_U5394;
  assign new_P2_U3839 = new_P2_U4443 & new_P2_U5408 & new_P2_U5409;
  assign new_P2_U3840 = new_P2_U5418 & new_P2_U5417 & new_P2_U5416;
  assign new_P2_U3841 = new_P2_U5423 & new_P2_U5422 & new_P2_U5421;
  assign new_P2_U3842 = new_P2_U5428 & new_P2_U5427 & new_P2_U5426;
  assign new_P2_U3843 = new_P2_U5433 & new_P2_U5432 & new_P2_U5431;
  assign new_P2_U3844 = new_P2_U5438 & new_P2_U5437 & new_P2_U5436;
  assign new_P2_U3845 = new_P2_U5443 & new_P2_U5442 & new_P2_U5441;
  assign new_P2_U3846 = new_P2_U5448 & new_P2_U5447 & new_P2_U5446;
  assign new_P2_U3847 = new_P2_U5453 & new_P2_U5452 & new_P2_U5451;
  assign new_P2_U3848 = new_P2_U4443 & new_P2_U5466 & new_P2_U5467;
  assign new_P2_U3849 = new_P2_U5476 & new_P2_U5475 & new_P2_U5474;
  assign new_P2_U3850 = new_P2_U5481 & new_P2_U5480 & new_P2_U5479;
  assign new_P2_U3851 = new_P2_U5486 & new_P2_U5485 & new_P2_U5484;
  assign new_P2_U3852 = new_P2_U5491 & new_P2_U5490 & new_P2_U5489;
  assign new_P2_U3853 = new_P2_U5496 & new_P2_U5495 & new_P2_U5494;
  assign new_P2_U3854 = new_P2_U5501 & new_P2_U5500 & new_P2_U5499;
  assign new_P2_U3855 = new_P2_U5506 & new_P2_U5505 & new_P2_U5504;
  assign new_P2_U3856 = new_P2_U5511 & new_P2_U5510 & new_P2_U5509;
  assign new_P2_U3857 = new_P2_U4443 & new_P2_U5523 & new_P2_U5524;
  assign new_P2_U3858 = new_P2_U5533 & new_P2_U5532 & new_P2_U5531;
  assign new_P2_U3859 = new_P2_U5538 & new_P2_U5537 & new_P2_U5536;
  assign new_P2_U3860 = new_P2_U5543 & new_P2_U5542 & new_P2_U5541;
  assign new_P2_U3861 = new_P2_U5548 & new_P2_U5547 & new_P2_U5546;
  assign new_P2_U3862 = new_P2_U5553 & new_P2_U5552 & new_P2_U5551;
  assign new_P2_U3863 = new_P2_U5558 & new_P2_U5557 & new_P2_U5556;
  assign new_P2_U3864 = new_P2_U5563 & new_P2_U5562 & new_P2_U5561;
  assign new_P2_U3865 = new_P2_U5568 & new_P2_U5567 & new_P2_U5566;
  assign new_P2_U3866 = new_P2_R2147_U7 & new_P2_U4466;
  assign new_P2_U3867 = P2_FLUSH_REG & P2_STATE2_REG_0_;
  assign new_P2_U3868 = new_P2_U5573 & new_P2_U5571;
  assign new_P2_U3869 = new_P2_U3868 & new_P2_U5576;
  assign new_P2_U3870 = new_P2_U4460 & new_P2_U4456;
  assign new_P2_U3871 = new_P2_U2512 & new_P2_U3870 & new_P2_U8071 & new_P2_U8070;
  assign new_P2_U3872 = new_P2_U5583 & new_P2_U4455;
  assign new_P2_U3873 = new_P2_U3521 & new_P2_U7869;
  assign new_P2_U3874 = new_P2_U7861 & new_P2_U3278;
  assign new_P2_U3875 = new_P2_U3874 & new_P2_U4429;
  assign new_P2_U3876 = new_P2_U4429 & new_P2_U3279;
  assign new_P2_U3877 = new_P2_U7859 & new_P2_U5593;
  assign new_P2_U3878 = new_P2_U7863 & new_P2_U3521;
  assign new_P2_U3879 = new_P2_U3281 & new_P2_U5587 & new_P2_U5588;
  assign new_P2_U3880 = new_P2_U5599 & new_P2_U3254;
  assign new_P2_U3881 = new_P2_U3880 & new_P2_U5601 & new_P2_U5600;
  assign new_P2_U3882 = new_P2_U7897 & new_P2_U5602;
  assign new_P2_U3883 = new_P2_U5608 & new_P2_U5607;
  assign new_P2_U3884 = new_P2_U3883 & new_P2_U5609;
  assign new_P2_U3885 = new_P2_U4396 & new_P2_U5617;
  assign new_P2_U3886 = new_P2_U4601 & new_P2_U2449;
  assign new_P2_U3887 = new_P2_U3582 & new_P2_U7859;
  assign new_P2_U3888 = new_P2_U5627 & new_P2_U5626;
  assign new_P2_U3889 = new_P2_U7859 & new_P2_U3272;
  assign new_P2_U3890 = new_P2_U5635 & new_P2_U5634;
  assign new_P2_U3891 = new_P2_U5649 & new_P2_U5650;
  assign new_P2_U3892 = new_P2_U5653 & new_P2_U5654;
  assign new_P2_U3893 = new_P2_U5658 & new_P2_U5659;
  assign new_P2_U3894 = new_P2_U4456 & new_P2_U4460 & new_P2_U5668;
  assign new_P2_U3895 = new_P2_U5674 & new_P2_U3578;
  assign new_P2_U3896 = new_P2_U5681 & new_P2_U5680;
  assign new_P2_U3897 = new_P2_U5683 & new_P2_U5682;
  assign new_P2_U3898 = new_P2_U5687 & new_P2_U5686;
  assign new_P2_U3899 = new_P2_U5689 & new_P2_U5688;
  assign new_P2_U3900 = new_P2_U5691 & new_P2_U5690;
  assign new_P2_U3901 = new_P2_U5695 & new_P2_U5694;
  assign new_P2_U3902 = new_P2_U5697 & new_P2_U5696;
  assign new_P2_U3903 = new_P2_U5699 & new_P2_U5698;
  assign new_P2_U3904 = new_P2_U5703 & new_P2_U5702;
  assign new_P2_U3905 = new_P2_U5705 & new_P2_U5704;
  assign new_P2_U3906 = new_P2_U5707 & new_P2_U5706;
  assign new_P2_U3907 = new_P2_U5711 & new_P2_U5710;
  assign new_P2_U3908 = new_P2_U5713 & new_P2_U5712;
  assign new_P2_U3909 = new_P2_U5715 & new_P2_U5714;
  assign new_P2_U3910 = new_P2_U5719 & new_P2_U5718;
  assign new_P2_U3911 = new_P2_U5721 & new_P2_U5720;
  assign new_P2_U3912 = new_P2_U5723 & new_P2_U5722;
  assign new_P2_U3913 = new_P2_U5727 & new_P2_U5726;
  assign new_P2_U3914 = new_P2_U5729 & new_P2_U5728;
  assign new_P2_U3915 = new_P2_U5731 & new_P2_U5730;
  assign new_P2_U3916 = new_P2_U5735 & new_P2_U5734;
  assign new_P2_U3917 = new_P2_U5737 & new_P2_U5736;
  assign new_P2_U3918 = new_P2_U5739 & new_P2_U5738;
  assign new_P2_U3919 = new_P2_U5743 & new_P2_U5742;
  assign new_P2_U3920 = new_P2_U5745 & new_P2_U5744;
  assign new_P2_U3921 = new_P2_U5747 & new_P2_U5746;
  assign new_P2_U3922 = new_P2_U5751 & new_P2_U5750;
  assign new_P2_U3923 = new_P2_U5753 & new_P2_U5752;
  assign new_P2_U3924 = new_P2_U5755 & new_P2_U5754;
  assign new_P2_U3925 = new_P2_U5759 & new_P2_U5758;
  assign new_P2_U3926 = new_P2_U5761 & new_P2_U5760;
  assign new_P2_U3927 = new_P2_U5763 & new_P2_U5762;
  assign new_P2_U3928 = new_P2_U5767 & new_P2_U5766;
  assign new_P2_U3929 = new_P2_U5769 & new_P2_U5768;
  assign new_P2_U3930 = new_P2_U5771 & new_P2_U5770;
  assign new_P2_U3931 = new_P2_U5775 & new_P2_U5774;
  assign new_P2_U3932 = new_P2_U5777 & new_P2_U5776;
  assign new_P2_U3933 = new_P2_U5779 & new_P2_U5778;
  assign new_P2_U3934 = new_P2_U5783 & new_P2_U5782;
  assign new_P2_U3935 = new_P2_U5785 & new_P2_U5784;
  assign new_P2_U3936 = new_P2_U5787 & new_P2_U5786;
  assign new_P2_U3937 = new_P2_U5791 & new_P2_U5790;
  assign new_P2_U3938 = new_P2_U5793 & new_P2_U5792;
  assign new_P2_U3939 = new_P2_U5795 & new_P2_U5794;
  assign new_P2_U3940 = new_P2_U5799 & new_P2_U5798;
  assign new_P2_U3941 = new_P2_U5801 & new_P2_U5800;
  assign new_P2_U3942 = new_P2_U5803 & new_P2_U5802;
  assign new_P2_U3943 = new_P2_U5807 & new_P2_U5806;
  assign new_P2_U3944 = new_P2_U5809 & new_P2_U5808;
  assign new_P2_U3945 = new_P2_U5811 & new_P2_U5810;
  assign new_P2_U3946 = new_P2_U5815 & new_P2_U5814;
  assign new_P2_U3947 = new_P2_U5817 & new_P2_U5816;
  assign new_P2_U3948 = new_P2_U5819 & new_P2_U5818;
  assign new_P2_U3949 = new_P2_U5823 & new_P2_U5822;
  assign new_P2_U3950 = new_P2_U5825 & new_P2_U5824;
  assign new_P2_U3951 = new_P2_U5827 & new_P2_U5826;
  assign new_P2_U3952 = new_P2_U5831 & new_P2_U5830;
  assign new_P2_U3953 = new_P2_U5833 & new_P2_U5832;
  assign new_P2_U3954 = new_P2_U5835 & new_P2_U5834;
  assign new_P2_U3955 = new_P2_U5839 & new_P2_U5838;
  assign new_P2_U3956 = new_P2_U5841 & new_P2_U5840;
  assign new_P2_U3957 = new_P2_U5843 & new_P2_U5842;
  assign new_P2_U3958 = new_P2_U5847 & new_P2_U5846;
  assign new_P2_U3959 = new_P2_U5849 & new_P2_U5848;
  assign new_P2_U3960 = new_P2_U5851 & new_P2_U5850;
  assign new_P2_U3961 = new_P2_U5855 & new_P2_U5854;
  assign new_P2_U3962 = new_P2_U5857 & new_P2_U5856;
  assign new_P2_U3963 = new_P2_U5859 & new_P2_U5858;
  assign new_P2_U3964 = new_P2_U5863 & new_P2_U5862;
  assign new_P2_U3965 = new_P2_U5865 & new_P2_U5864;
  assign new_P2_U3966 = new_P2_U5867 & new_P2_U5866;
  assign new_P2_U3967 = new_P2_U5871 & new_P2_U5870;
  assign new_P2_U3968 = new_P2_U5873 & new_P2_U5872;
  assign new_P2_U3969 = new_P2_U5875 & new_P2_U5874;
  assign new_P2_U3970 = new_P2_U5879 & new_P2_U5878;
  assign new_P2_U3971 = new_P2_U5881 & new_P2_U5880;
  assign new_P2_U3972 = new_P2_U5883 & new_P2_U5882;
  assign new_P2_U3973 = new_P2_U5887 & new_P2_U5886;
  assign new_P2_U3974 = new_P2_U5889 & new_P2_U5888;
  assign new_P2_U3975 = new_P2_U5891 & new_P2_U5890;
  assign new_P2_U3976 = new_P2_U5895 & new_P2_U5894;
  assign new_P2_U3977 = new_P2_U5897 & new_P2_U5896;
  assign new_P2_U3978 = new_P2_U5899 & new_P2_U5898;
  assign new_P2_U3979 = new_P2_U5903 & new_P2_U5902;
  assign new_P2_U3980 = new_P2_U5905 & new_P2_U5904;
  assign new_P2_U3981 = new_P2_U5907 & new_P2_U5906;
  assign new_P2_U3982 = new_P2_U5911 & new_P2_U5910;
  assign new_P2_U3983 = new_P2_U5912 & new_P2_U5913 & new_P2_U5915 & new_P2_U5914;
  assign new_P2_U3984 = new_P2_U5919 & new_P2_U5918;
  assign new_P2_U3985 = new_P2_U5921 & new_P2_U5923 & new_P2_U5922;
  assign new_P2_U3986 = new_P2_U5927 & new_P2_U5926;
  assign new_P2_U3987 = new_P2_U5929 & new_P2_U5931 & new_P2_U5930;
  assign new_P2_U3988 = new_P2_U5935 & new_P2_U5934;
  assign new_P2_U3989 = P2_STATE2_REG_1_ & P2_STATEBS16_REG;
  assign new_P2_U3990 = ~P2_STATE2_REG_2_ & ~P2_STATE2_REG_1_;
  assign new_P2_U3991 = new_P2_U5943 & new_P2_U5942 & new_P2_U5941;
  assign new_P2_U3992 = new_P2_U5946 & new_P2_U5945 & new_P2_U5944;
  assign new_P2_U3993 = new_P2_U5949 & new_P2_U5948 & new_P2_U5947;
  assign new_P2_U3994 = new_P2_U5952 & new_P2_U5951 & new_P2_U5950;
  assign new_P2_U3995 = new_P2_U5955 & new_P2_U5954 & new_P2_U5953;
  assign new_P2_U3996 = new_P2_U5958 & new_P2_U5957 & new_P2_U5956;
  assign new_P2_U3997 = new_P2_U5961 & new_P2_U5960 & new_P2_U5959;
  assign new_P2_U3998 = new_P2_U5964 & new_P2_U5963 & new_P2_U5962;
  assign new_P2_U3999 = new_P2_U5967 & new_P2_U5966 & new_P2_U5965;
  assign new_P2_U4000 = new_P2_U5970 & new_P2_U5969 & new_P2_U5968;
  assign new_P2_U4001 = new_P2_U5973 & new_P2_U5972 & new_P2_U5971;
  assign new_P2_U4002 = new_P2_U5976 & new_P2_U5975 & new_P2_U5974;
  assign new_P2_U4003 = new_P2_U5979 & new_P2_U5978 & new_P2_U5977;
  assign new_P2_U4004 = new_P2_U5982 & new_P2_U5981 & new_P2_U5980;
  assign new_P2_U4005 = new_P2_U5985 & new_P2_U5984 & new_P2_U5983;
  assign new_P2_U4006 = new_P2_U5988 & new_P2_U5987 & new_P2_U5986;
  assign new_P2_U4007 = new_P2_U5991 & new_P2_U5990 & new_P2_U5989;
  assign new_P2_U4008 = new_P2_U5994 & new_P2_U5993 & new_P2_U5992;
  assign new_P2_U4009 = new_P2_U5997 & new_P2_U5996 & new_P2_U5995;
  assign new_P2_U4010 = new_P2_U6000 & new_P2_U5999 & new_P2_U5998;
  assign new_P2_U4011 = new_P2_U6003 & new_P2_U6002 & new_P2_U6001;
  assign new_P2_U4012 = new_P2_U6006 & new_P2_U6005 & new_P2_U6004;
  assign new_P2_U4013 = new_P2_U6009 & new_P2_U6008 & new_P2_U6007;
  assign new_P2_U4014 = new_P2_U6012 & new_P2_U6011 & new_P2_U6010;
  assign new_P2_U4015 = new_P2_U6015 & new_P2_U6014 & new_P2_U6013;
  assign new_P2_U4016 = new_P2_U6018 & new_P2_U6017 & new_P2_U6016;
  assign new_P2_U4017 = new_P2_U6021 & new_P2_U6020 & new_P2_U6019;
  assign new_P2_U4018 = new_P2_U6024 & new_P2_U6023 & new_P2_U6022;
  assign new_P2_U4019 = new_P2_U6027 & new_P2_U6026 & new_P2_U6025;
  assign new_P2_U4020 = new_P2_U6030 & new_P2_U6029 & new_P2_U6028;
  assign new_P2_U4021 = new_P2_U6033 & new_P2_U6032 & new_P2_U6031;
  assign new_P2_U4022 = new_P2_U6036 & new_P2_U6035 & new_P2_U6034;
  assign new_P2_U4023 = new_P2_U6039 & new_P2_U6038 & new_P2_U6037;
  assign new_P2_U4024 = new_P2_U6042 & new_P2_U6041 & new_P2_U6040;
  assign new_P2_U4025 = new_P2_U6045 & new_P2_U6044 & new_P2_U6043;
  assign new_P2_U4026 = new_P2_U6048 & new_P2_U6047 & new_P2_U6046;
  assign new_P2_U4027 = new_P2_U6051 & new_P2_U6050 & new_P2_U6049;
  assign new_P2_U4028 = new_P2_U6054 & new_P2_U6053 & new_P2_U6052;
  assign new_P2_U4029 = new_P2_U6057 & new_P2_U6056 & new_P2_U6055;
  assign new_P2_U4030 = new_P2_U6060 & new_P2_U6059 & new_P2_U6058;
  assign new_P2_U4031 = new_P2_U6063 & new_P2_U6062 & new_P2_U6061;
  assign new_P2_U4032 = new_P2_U6066 & new_P2_U6065 & new_P2_U6064;
  assign new_P2_U4033 = new_P2_U6069 & new_P2_U6068 & new_P2_U6067;
  assign new_P2_U4034 = new_P2_U6072 & new_P2_U6071 & new_P2_U6070;
  assign new_P2_U4035 = new_P2_U6075 & new_P2_U6074 & new_P2_U6073;
  assign new_P2_U4036 = new_P2_U6078 & new_P2_U6077 & new_P2_U6076;
  assign new_P2_U4037 = new_P2_U6081 & new_P2_U6080 & new_P2_U6079;
  assign new_P2_U4038 = new_P2_U6084 & new_P2_U6083 & new_P2_U6082;
  assign new_P2_U4039 = new_P2_U6087 & new_P2_U6086 & new_P2_U6085;
  assign new_P2_U4040 = new_P2_U6090 & new_P2_U6089 & new_P2_U6088;
  assign new_P2_U4041 = new_P2_U6093 & new_P2_U6092 & new_P2_U6091;
  assign new_P2_U4042 = new_P2_U6096 & new_P2_U6095 & new_P2_U6094;
  assign new_P2_U4043 = new_P2_U6099 & new_P2_U6098 & new_P2_U6097;
  assign new_P2_U4044 = new_P2_U6102 & new_P2_U6101 & new_P2_U6100;
  assign new_P2_U4045 = new_P2_U6105 & new_P2_U6104 & new_P2_U6103;
  assign new_P2_U4046 = new_P2_U6108 & new_P2_U6107 & new_P2_U6106;
  assign new_P2_U4047 = new_P2_U6111 & new_P2_U6110 & new_P2_U6109;
  assign new_P2_U4048 = new_P2_U6114 & new_P2_U6113 & new_P2_U6112;
  assign new_P2_U4049 = new_P2_U6117 & new_P2_U6116 & new_P2_U6115;
  assign new_P2_U4050 = new_P2_U6120 & new_P2_U6119 & new_P2_U6118;
  assign new_P2_U4051 = new_P2_U6123 & new_P2_U6122 & new_P2_U6121;
  assign new_P2_U4052 = new_P2_U6125 & new_P2_U6126 & new_P2_U6124;
  assign new_P2_U4053 = new_P2_U6129 & new_P2_U6128 & new_P2_U6127;
  assign new_P2_U4054 = new_P2_U6132 & new_P2_U6131 & new_P2_U6130;
  assign new_P2_U4055 = new_P2_U2356 & new_P2_U4468 & new_P2_U6133;
  assign new_P2_U4056 = new_P2_U7871 & new_P2_U3280 & P2_STATE2_REG_0_;
  assign new_P2_U4057 = new_P2_U2616 & new_P2_U4468;
  assign new_P2_U4058 = new_P2_U2374 & new_P2_U4417;
  assign new_P2_U4059 = new_P2_U6330 & new_P2_U6329;
  assign new_P2_U4060 = new_P2_U6334 & new_P2_U6333;
  assign new_P2_U4061 = new_P2_U6338 & new_P2_U6337;
  assign new_P2_U4062 = new_P2_U6342 & new_P2_U6341;
  assign new_P2_U4063 = new_P2_U6346 & new_P2_U6345;
  assign new_P2_U4064 = new_P2_U6350 & new_P2_U6349;
  assign new_P2_U4065 = new_P2_U6354 & new_P2_U6353;
  assign new_P2_U4066 = new_P2_U6358 & new_P2_U6357;
  assign new_P2_U4067 = new_P2_U6362 & new_P2_U6361;
  assign new_P2_U4068 = new_P2_U6366 & new_P2_U6365;
  assign new_P2_U4069 = new_P2_U6569 & new_P2_U4454 & new_P2_U4453;
  assign new_P2_U4070 = new_P2_U4071 & new_P2_U6574 & new_P2_U6573;
  assign new_P2_U4071 = new_P2_U6577 & new_P2_U6576;
  assign new_P2_U4072 = new_P2_U4073 & new_P2_U6578;
  assign new_P2_U4073 = new_P2_U6581 & new_P2_U6580;
  assign new_P2_U4074 = new_P2_U4075 & new_P2_U6583 & new_P2_U6582;
  assign new_P2_U4075 = new_P2_U6586 & new_P2_U6585;
  assign new_P2_U4076 = new_P2_U4077 & new_P2_U6587;
  assign new_P2_U4077 = new_P2_U6590 & new_P2_U6589;
  assign new_P2_U4078 = new_P2_U4079 & new_P2_U6592 & new_P2_U6591;
  assign new_P2_U4079 = new_P2_U6595 & new_P2_U6594;
  assign new_P2_U4080 = new_P2_U4081 & new_P2_U6596;
  assign new_P2_U4081 = new_P2_U6599 & new_P2_U6598;
  assign new_P2_U4082 = new_P2_U4083 & new_P2_U6601 & new_P2_U6600;
  assign new_P2_U4083 = new_P2_U6604 & new_P2_U6603;
  assign new_P2_U4084 = new_P2_U4085 & new_P2_U6605;
  assign new_P2_U4085 = new_P2_U6608 & new_P2_U6607;
  assign new_P2_U4086 = new_P2_U6610 & new_P2_U6609 & new_P2_U4446;
  assign new_P2_U4087 = new_P2_U4088 & new_P2_U6615;
  assign new_P2_U4088 = new_P2_U6617 & new_P2_U6616;
  assign new_P2_U4089 = new_P2_U6614 & new_P2_U6613 & new_P2_U4086 & new_P2_U6612 & new_P2_U6611;
  assign new_P2_U4090 = new_P2_U6619 & new_P2_U6618 & new_P2_U4446;
  assign new_P2_U4091 = new_P2_U4092 & new_P2_U6624;
  assign new_P2_U4092 = new_P2_U6626 & new_P2_U6625;
  assign new_P2_U4093 = new_P2_U6623 & new_P2_U6622 & new_P2_U4090 & new_P2_U6621 & new_P2_U6620;
  assign new_P2_U4094 = new_P2_U6628 & new_P2_U6627 & new_P2_U4446;
  assign new_P2_U4095 = new_P2_U4096 & new_P2_U6631;
  assign new_P2_U4096 = new_P2_U6634 & new_P2_U6633;
  assign new_P2_U4097 = new_P2_U6636 & new_P2_U6635 & new_P2_U4446;
  assign new_P2_U4098 = new_P2_U4099 & new_P2_U6639;
  assign new_P2_U4099 = new_P2_U6642 & new_P2_U6641;
  assign new_P2_U4100 = new_P2_U6644 & new_P2_U6643 & new_P2_U4446;
  assign new_P2_U4101 = new_P2_U4102 & new_P2_U6647;
  assign new_P2_U4102 = new_P2_U6650 & new_P2_U6649;
  assign new_P2_U4103 = new_P2_U6652 & new_P2_U6651 & new_P2_U4446;
  assign new_P2_U4104 = new_P2_U4105 & new_P2_U6655;
  assign new_P2_U4105 = new_P2_U6658 & new_P2_U6657;
  assign new_P2_U4106 = new_P2_U6660 & new_P2_U6659 & new_P2_U4446;
  assign new_P2_U4107 = new_P2_U4108 & new_P2_U6663;
  assign new_P2_U4108 = new_P2_U6666 & new_P2_U6665;
  assign new_P2_U4109 = new_P2_U6668 & new_P2_U6667 & new_P2_U4446;
  assign new_P2_U4110 = new_P2_U4111 & new_P2_U6671;
  assign new_P2_U4111 = new_P2_U6674 & new_P2_U6673;
  assign new_P2_U4112 = new_P2_U6678 & new_P2_U6675 & new_P2_U4446;
  assign new_P2_U4113 = new_P2_U4114 & new_P2_U6679;
  assign new_P2_U4114 = new_P2_U6682 & new_P2_U6681;
  assign new_P2_U4115 = new_P2_U6686 & new_P2_U6683 & new_P2_U4446;
  assign new_P2_U4116 = new_P2_U4117 & new_P2_U6687;
  assign new_P2_U4117 = new_P2_U6690 & new_P2_U6689;
  assign new_P2_U4118 = new_P2_U6694 & new_P2_U6691 & new_P2_U4446;
  assign new_P2_U4119 = new_P2_U4120 & new_P2_U6695;
  assign new_P2_U4120 = new_P2_U6698 & new_P2_U6697;
  assign new_P2_U4121 = new_P2_U6699 & new_P2_U4446;
  assign new_P2_U4122 = new_P2_U4123 & new_P2_U6703;
  assign new_P2_U4123 = new_P2_U6706 & new_P2_U6705;
  assign new_P2_U4124 = new_P2_U6704 & new_P2_U6700 & new_P2_U6702 & new_P2_U4121 & new_P2_U6701;
  assign new_P2_U4125 = new_P2_U6707 & new_P2_U4446;
  assign new_P2_U4126 = new_P2_U4127 & new_P2_U6711;
  assign new_P2_U4127 = new_P2_U6714 & new_P2_U6713;
  assign new_P2_U4128 = new_P2_U6712 & new_P2_U6708 & new_P2_U6710 & new_P2_U4125 & new_P2_U6709;
  assign new_P2_U4129 = new_P2_U6715 & new_P2_U4446;
  assign new_P2_U4130 = new_P2_U4131 & new_P2_U6719;
  assign new_P2_U4131 = new_P2_U6722 & new_P2_U6721;
  assign new_P2_U4132 = new_P2_U6720 & new_P2_U6716 & new_P2_U6718 & new_P2_U4129 & new_P2_U6717;
  assign new_P2_U4133 = new_P2_U6723 & new_P2_U4446;
  assign new_P2_U4134 = new_P2_U4135 & new_P2_U6727;
  assign new_P2_U4135 = new_P2_U6730 & new_P2_U6729;
  assign new_P2_U4136 = new_P2_U6728 & new_P2_U6724 & new_P2_U6726 & new_P2_U4133 & new_P2_U6725;
  assign new_P2_U4137 = new_P2_U6731 & new_P2_U4446;
  assign new_P2_U4138 = new_P2_U4139 & new_P2_U6735;
  assign new_P2_U4139 = new_P2_U6738 & new_P2_U6737;
  assign new_P2_U4140 = new_P2_U6736 & new_P2_U6732 & new_P2_U6734 & new_P2_U4137 & new_P2_U6733;
  assign new_P2_U4141 = new_P2_U4142 & new_P2_U6743;
  assign new_P2_U4142 = new_P2_U6746 & new_P2_U6745;
  assign new_P2_U4143 = new_P2_U6744 & new_P2_U6740 & new_P2_U6742 & new_P2_U6739 & new_P2_U6741;
  assign new_P2_U4144 = new_P2_U4145 & new_P2_U6751;
  assign new_P2_U4145 = new_P2_U6754 & new_P2_U6753;
  assign new_P2_U4146 = new_P2_U6752 & new_P2_U6748 & new_P2_U6750 & new_P2_U6747 & new_P2_U6749;
  assign new_P2_U4147 = new_P2_U6762 & new_P2_U6761;
  assign new_P2_U4148 = new_P2_U6760 & new_P2_U4147 & new_P2_U6759;
  assign new_P2_U4149 = new_P2_U4150 & new_P2_U6768 & new_P2_U6766 & new_P2_U6763 & new_P2_U6765;
  assign new_P2_U4150 = new_P2_U4151 & new_P2_U6767;
  assign new_P2_U4151 = new_P2_U6770 & new_P2_U6769;
  assign new_P2_U4152 = new_P2_U4153 & new_P2_U6776 & new_P2_U6774 & new_P2_U6771 & new_P2_U6773;
  assign new_P2_U4153 = new_P2_U4154 & new_P2_U6775;
  assign new_P2_U4154 = new_P2_U6778 & new_P2_U6777;
  assign new_P2_U4155 = new_P2_U6786 & new_P2_U6785;
  assign new_P2_U4156 = new_P2_U6784 & new_P2_U4155 & new_P2_U6783;
  assign new_P2_U4157 = new_P2_U6794 & new_P2_U6793;
  assign new_P2_U4158 = new_P2_U6792 & new_P2_U4157 & new_P2_U6791;
  assign new_P2_U4159 = new_P2_U6802 & new_P2_U6801;
  assign new_P2_U4160 = new_P2_U6800 & new_P2_U4159 & new_P2_U6799;
  assign new_P2_U4161 = new_P2_U6810 & new_P2_U6809;
  assign new_P2_U4162 = new_P2_U6808 & new_P2_U4161 & new_P2_U6807;
  assign new_P2_U4163 = new_P2_U6818 & new_P2_U6817;
  assign new_P2_U4164 = new_P2_U6816 & new_P2_U4163 & new_P2_U6815;
  assign new_P2_U4165 = new_P2_U6826 & new_P2_U6825;
  assign new_P2_U4166 = new_P2_U6824 & new_P2_U4165 & new_P2_U6823;
  assign new_P2_U4167 = new_P2_U6834 & new_P2_U6833;
  assign new_P2_U4168 = new_P2_U6832 & new_P2_U4167 & new_P2_U6831;
  assign new_P2_U4169 = ~P2_DATAWIDTH_REG_5_ & ~P2_DATAWIDTH_REG_4_ & ~P2_DATAWIDTH_REG_2_ & ~P2_DATAWIDTH_REG_3_;
  assign new_P2_U4170 = ~P2_DATAWIDTH_REG_9_ & ~P2_DATAWIDTH_REG_8_ & ~P2_DATAWIDTH_REG_6_ & ~P2_DATAWIDTH_REG_7_;
  assign new_P2_U4171 = new_P2_U4170 & new_P2_U4169;
  assign new_P2_U4172 = ~P2_DATAWIDTH_REG_13_ & ~P2_DATAWIDTH_REG_12_ & ~P2_DATAWIDTH_REG_10_ & ~P2_DATAWIDTH_REG_11_;
  assign new_P2_U4173 = ~P2_DATAWIDTH_REG_17_ & ~P2_DATAWIDTH_REG_16_ & ~P2_DATAWIDTH_REG_14_ & ~P2_DATAWIDTH_REG_15_;
  assign new_P2_U4174 = new_P2_U4173 & new_P2_U4172;
  assign new_P2_U4175 = ~P2_DATAWIDTH_REG_21_ & ~P2_DATAWIDTH_REG_20_ & ~P2_DATAWIDTH_REG_18_ & ~P2_DATAWIDTH_REG_19_;
  assign new_P2_U4176 = ~P2_DATAWIDTH_REG_25_ & ~P2_DATAWIDTH_REG_24_ & ~P2_DATAWIDTH_REG_22_ & ~P2_DATAWIDTH_REG_23_;
  assign new_P2_U4177 = new_P2_U4176 & new_P2_U4175;
  assign new_P2_U4178 = ~P2_DATAWIDTH_REG_26_ & ~P2_DATAWIDTH_REG_27_;
  assign new_P2_U4179 = ~P2_DATAWIDTH_REG_28_ & ~P2_DATAWIDTH_REG_29_;
  assign new_P2_U4180 = ~P2_DATAWIDTH_REG_30_ & ~P2_DATAWIDTH_REG_31_;
  assign new_P2_U4181 = new_P2_U4178 & new_P2_U4179 & new_P2_U4180 & new_P2_U6835;
  assign new_P2_U4182 = ~P2_DATAWIDTH_REG_0_ & ~P2_DATAWIDTH_REG_1_ & ~P2_REIP_REG_0_;
  assign new_P2_U4183 = ~P2_REIP_REG_1_ & ~P2_DATAWIDTH_REG_1_;
  assign new_P2_U4184 = new_P2_U6844 & new_P2_U7873;
  assign new_P2_U4185 = new_P2_U6848 & new_P2_U3301;
  assign new_P2_U4186 = new_P2_U4185 & new_P2_U6849;
  assign new_P2_U4187 = P2_STATE2_REG_1_ & new_P2_U3265;
  assign new_P2_U4188 = new_P2_U6841 & new_P2_U6842 & new_P2_U3313;
  assign new_P2_U4189 = new_P2_U2374 & new_P2_U3253;
  assign new_P2_U4190 = new_P2_U6860 & new_P2_U3534;
  assign new_P2_U4191 = new_P2_U6862 & new_P2_U6863 & new_P2_U6865 & new_P2_U6864;
  assign new_P2_U4192 = new_P2_U6866 & new_P2_U6867 & new_P2_U6869 & new_P2_U6868;
  assign new_P2_U4193 = new_P2_U6870 & new_P2_U6871 & new_P2_U6873 & new_P2_U6872;
  assign new_P2_U4194 = new_P2_U6874 & new_P2_U6875 & new_P2_U6877 & new_P2_U6876;
  assign new_P2_U4195 = new_P2_U6878 & new_P2_U6879 & new_P2_U6881 & new_P2_U6880;
  assign new_P2_U4196 = new_P2_U6882 & new_P2_U6883 & new_P2_U6885 & new_P2_U6884;
  assign new_P2_U4197 = new_P2_U6886 & new_P2_U6887 & new_P2_U6889 & new_P2_U6888;
  assign new_P2_U4198 = new_P2_U6890 & new_P2_U6891 & new_P2_U6893 & new_P2_U6892;
  assign new_P2_U4199 = new_P2_U6894 & new_P2_U6895 & new_P2_U6897 & new_P2_U6896;
  assign new_P2_U4200 = new_P2_U6898 & new_P2_U6899 & new_P2_U6901 & new_P2_U6900;
  assign new_P2_U4201 = new_P2_U6902 & new_P2_U6903 & new_P2_U6905 & new_P2_U6904;
  assign new_P2_U4202 = new_P2_U6906 & new_P2_U6907 & new_P2_U6909 & new_P2_U6908;
  assign new_P2_U4203 = new_P2_U6910 & new_P2_U6911 & new_P2_U6913 & new_P2_U6912;
  assign new_P2_U4204 = new_P2_U6914 & new_P2_U6915 & new_P2_U6917 & new_P2_U6916;
  assign new_P2_U4205 = new_P2_U6918 & new_P2_U6919 & new_P2_U6921 & new_P2_U6920;
  assign new_P2_U4206 = new_P2_U6922 & new_P2_U6923 & new_P2_U6925 & new_P2_U6924;
  assign new_P2_U4207 = new_P2_U6926 & new_P2_U6927 & new_P2_U6929 & new_P2_U6928;
  assign new_P2_U4208 = new_P2_U6930 & new_P2_U6931 & new_P2_U6933 & new_P2_U6932;
  assign new_P2_U4209 = new_P2_U6934 & new_P2_U6935 & new_P2_U6937 & new_P2_U6936;
  assign new_P2_U4210 = new_P2_U6938 & new_P2_U6939 & new_P2_U6941 & new_P2_U6940;
  assign new_P2_U4211 = new_P2_U6942 & new_P2_U6943 & new_P2_U6945 & new_P2_U6944;
  assign new_P2_U4212 = new_P2_U6946 & new_P2_U6947 & new_P2_U6949 & new_P2_U6948;
  assign new_P2_U4213 = new_P2_U6950 & new_P2_U6951 & new_P2_U6953 & new_P2_U6952;
  assign new_P2_U4214 = new_P2_U6954 & new_P2_U6955 & new_P2_U6957 & new_P2_U6956;
  assign new_P2_U4215 = new_P2_U6958 & new_P2_U6959 & new_P2_U6961 & new_P2_U6960;
  assign new_P2_U4216 = new_P2_U6962 & new_P2_U6963 & new_P2_U6965 & new_P2_U6964;
  assign new_P2_U4217 = new_P2_U6966 & new_P2_U6967 & new_P2_U6969 & new_P2_U6968;
  assign new_P2_U4218 = new_P2_U6970 & new_P2_U6971 & new_P2_U6973 & new_P2_U6972;
  assign new_P2_U4219 = new_P2_U6974 & new_P2_U6975 & new_P2_U6977 & new_P2_U6976;
  assign new_P2_U4220 = new_P2_U6978 & new_P2_U6979 & new_P2_U6981 & new_P2_U6980;
  assign new_P2_U4221 = new_P2_U6982 & new_P2_U6983 & new_P2_U6985 & new_P2_U6984;
  assign new_P2_U4222 = new_P2_U6986 & new_P2_U6987 & new_P2_U6989 & new_P2_U6988;
  assign new_P2_U4223 = new_P2_U6990 & new_P2_U6991 & new_P2_U6993 & new_P2_U6992;
  assign new_P2_U4224 = new_P2_U6994 & new_P2_U6995 & new_P2_U6997 & new_P2_U6996;
  assign new_P2_U4225 = new_P2_U6998 & new_P2_U6999 & new_P2_U7001 & new_P2_U7000;
  assign new_P2_U4226 = new_P2_U7002 & new_P2_U7003 & new_P2_U7005 & new_P2_U7004;
  assign new_P2_U4227 = new_P2_U7008 & new_P2_U7009 & new_P2_U7011 & new_P2_U7010;
  assign new_P2_U4228 = new_P2_U7012 & new_P2_U7013 & new_P2_U7015 & new_P2_U7014;
  assign new_P2_U4229 = new_P2_U7016 & new_P2_U7017 & new_P2_U7019 & new_P2_U7018;
  assign new_P2_U4230 = new_P2_U7020 & new_P2_U7021 & new_P2_U7023 & new_P2_U7022;
  assign new_P2_U4231 = new_P2_U7024 & new_P2_U7025 & new_P2_U7027 & new_P2_U7026;
  assign new_P2_U4232 = new_P2_U7028 & new_P2_U7029 & new_P2_U7031 & new_P2_U7030;
  assign new_P2_U4233 = new_P2_U7032 & new_P2_U7033 & new_P2_U7035 & new_P2_U7034;
  assign new_P2_U4234 = new_P2_U7036 & new_P2_U7037 & new_P2_U7039 & new_P2_U7038;
  assign new_P2_U4235 = new_P2_U7040 & new_P2_U7041 & new_P2_U7043 & new_P2_U7042;
  assign new_P2_U4236 = new_P2_U7044 & new_P2_U7045 & new_P2_U7047 & new_P2_U7046;
  assign new_P2_U4237 = new_P2_U7048 & new_P2_U7049 & new_P2_U7051 & new_P2_U7050;
  assign new_P2_U4238 = new_P2_U7052 & new_P2_U7053 & new_P2_U7055 & new_P2_U7054;
  assign new_P2_U4239 = new_P2_U7056 & new_P2_U7057 & new_P2_U7059 & new_P2_U7058;
  assign new_P2_U4240 = new_P2_U7060 & new_P2_U7061 & new_P2_U7063 & new_P2_U7062;
  assign new_P2_U4241 = new_P2_U7064 & new_P2_U7065 & new_P2_U7067 & new_P2_U7066;
  assign new_P2_U4242 = new_P2_U7068 & new_P2_U7069 & new_P2_U7071 & new_P2_U7070;
  assign new_P2_U4243 = new_P2_U7072 & new_P2_U7073 & new_P2_U7075 & new_P2_U7074;
  assign new_P2_U4244 = new_P2_U7076 & new_P2_U7077 & new_P2_U7079 & new_P2_U7078;
  assign new_P2_U4245 = new_P2_U7080 & new_P2_U7081 & new_P2_U7083 & new_P2_U7082;
  assign new_P2_U4246 = new_P2_U7084 & new_P2_U7085 & new_P2_U7087 & new_P2_U7086;
  assign new_P2_U4247 = new_P2_U7088 & new_P2_U7089 & new_P2_U7091 & new_P2_U7090;
  assign new_P2_U4248 = new_P2_U7092 & new_P2_U7093 & new_P2_U7095 & new_P2_U7094;
  assign new_P2_U4249 = new_P2_U7096 & new_P2_U7097 & new_P2_U7099 & new_P2_U7098;
  assign new_P2_U4250 = new_P2_U7100 & new_P2_U7101 & new_P2_U7103 & new_P2_U7102;
  assign new_P2_U4251 = new_P2_U7104 & new_P2_U7105 & new_P2_U7107 & new_P2_U7106;
  assign new_P2_U4252 = new_P2_U7108 & new_P2_U7109 & new_P2_U7111 & new_P2_U7110;
  assign new_P2_U4253 = new_P2_U7112 & new_P2_U7113 & new_P2_U7115 & new_P2_U7114;
  assign new_P2_U4254 = new_P2_U7116 & new_P2_U7117 & new_P2_U7119 & new_P2_U7118;
  assign new_P2_U4255 = new_P2_U7120 & new_P2_U7121 & new_P2_U7123 & new_P2_U7122;
  assign new_P2_U4256 = new_P2_U7124 & new_P2_U7125 & new_P2_U7127 & new_P2_U7126;
  assign new_P2_U4257 = new_P2_U7128 & new_P2_U7129 & new_P2_U7131 & new_P2_U7130;
  assign new_P2_U4258 = new_P2_U7132 & new_P2_U7133 & new_P2_U7135 & new_P2_U7134;
  assign new_P2_U4259 = new_P2_U7754 & new_P2_U7770 & new_P2_U7802 & new_P2_U7786;
  assign new_P2_U4260 = new_P2_U7818 & new_P2_U7834 & new_P2_U7874 & new_P2_U7850;
  assign new_P2_U4261 = new_P2_U7755 & new_P2_U7771 & new_P2_U7803 & new_P2_U7787;
  assign new_P2_U4262 = new_P2_U7819 & new_P2_U7835 & new_P2_U7875 & new_P2_U7851;
  assign new_P2_U4263 = new_P2_U7756 & new_P2_U7772 & new_P2_U7804 & new_P2_U7788;
  assign new_P2_U4264 = new_P2_U7820 & new_P2_U7836 & new_P2_U7876 & new_P2_U7852;
  assign new_P2_U4265 = new_P2_U7757 & new_P2_U7773 & new_P2_U7805 & new_P2_U7789;
  assign new_P2_U4266 = new_P2_U7821 & new_P2_U7837 & new_P2_U7877 & new_P2_U7853;
  assign new_P2_U4267 = new_P2_U7758 & new_P2_U7774 & new_P2_U7806 & new_P2_U7790;
  assign new_P2_U4268 = new_P2_U7822 & new_P2_U7838 & new_P2_U7878 & new_P2_U7854;
  assign new_P2_U4269 = new_P2_U7759 & new_P2_U7775 & new_P2_U7807 & new_P2_U7791;
  assign new_P2_U4270 = new_P2_U7823 & new_P2_U7839 & new_P2_U7879 & new_P2_U7855;
  assign new_P2_U4271 = new_P2_U7760 & new_P2_U7776 & new_P2_U7808 & new_P2_U7792;
  assign new_P2_U4272 = new_P2_U7824 & new_P2_U7840 & new_P2_U7880 & new_P2_U7856;
  assign new_P2_U4273 = new_P2_U7761 & new_P2_U7777 & new_P2_U7809 & new_P2_U7793;
  assign new_P2_U4274 = new_P2_U7825 & new_P2_U7841 & new_P2_U7881 & new_P2_U7857;
  assign new_P2_U4275 = new_P2_U7861 & new_P2_U4276;
  assign new_P2_U4276 = P2_STATE2_REG_0_ & P2_STATE2_REG_2_ & new_P2_U3300;
  assign new_P2_U4277 = new_P2_U7167 & new_P2_U7168 & new_P2_U7170 & new_P2_U7169;
  assign new_P2_U4278 = new_P2_U7171 & new_P2_U7172 & new_P2_U7174 & new_P2_U7173;
  assign new_P2_U4279 = new_P2_U7175 & new_P2_U7176 & new_P2_U7178 & new_P2_U7177;
  assign new_P2_U4280 = new_P2_U7179 & new_P2_U7180 & new_P2_U7182 & new_P2_U7181;
  assign new_P2_U4281 = new_P2_U7184 & new_P2_U7185 & new_P2_U7187 & new_P2_U7186;
  assign new_P2_U4282 = new_P2_U7188 & new_P2_U7189 & new_P2_U7191 & new_P2_U7190;
  assign new_P2_U4283 = new_P2_U7192 & new_P2_U7193 & new_P2_U7195 & new_P2_U7194;
  assign new_P2_U4284 = new_P2_U7196 & new_P2_U7197 & new_P2_U7199 & new_P2_U7198;
  assign new_P2_U4285 = new_P2_U7201 & new_P2_U7202 & new_P2_U7204 & new_P2_U7203;
  assign new_P2_U4286 = new_P2_U7205 & new_P2_U7206 & new_P2_U7208 & new_P2_U7207;
  assign new_P2_U4287 = new_P2_U7209 & new_P2_U7210 & new_P2_U7212 & new_P2_U7211;
  assign new_P2_U4288 = new_P2_U7213 & new_P2_U7214 & new_P2_U7216 & new_P2_U7215;
  assign new_P2_U4289 = new_P2_U7218 & new_P2_U7219 & new_P2_U7221 & new_P2_U7220;
  assign new_P2_U4290 = new_P2_U7222 & new_P2_U7223 & new_P2_U7225 & new_P2_U7224;
  assign new_P2_U4291 = new_P2_U7226 & new_P2_U7227 & new_P2_U7229 & new_P2_U7228;
  assign new_P2_U4292 = new_P2_U7230 & new_P2_U7231 & new_P2_U7233 & new_P2_U7232;
  assign new_P2_U4293 = new_P2_U7235 & new_P2_U7236 & new_P2_U7238 & new_P2_U7237;
  assign new_P2_U4294 = new_P2_U7239 & new_P2_U7240 & new_P2_U7242 & new_P2_U7241;
  assign new_P2_U4295 = new_P2_U7243 & new_P2_U7244 & new_P2_U7246 & new_P2_U7245;
  assign new_P2_U4296 = new_P2_U7247 & new_P2_U7248 & new_P2_U7250 & new_P2_U7249;
  assign new_P2_U4297 = new_P2_U7252 & new_P2_U7253 & new_P2_U7255 & new_P2_U7254;
  assign new_P2_U4298 = new_P2_U7256 & new_P2_U7257 & new_P2_U7259 & new_P2_U7258;
  assign new_P2_U4299 = new_P2_U7260 & new_P2_U7261 & new_P2_U7263 & new_P2_U7262;
  assign new_P2_U4300 = new_P2_U7264 & new_P2_U7265 & new_P2_U7267 & new_P2_U7266;
  assign new_P2_U4301 = new_P2_U7269 & new_P2_U7270 & new_P2_U7272 & new_P2_U7271;
  assign new_P2_U4302 = new_P2_U7273 & new_P2_U7274 & new_P2_U7276 & new_P2_U7275;
  assign new_P2_U4303 = new_P2_U7277 & new_P2_U7278 & new_P2_U7280 & new_P2_U7279;
  assign new_P2_U4304 = new_P2_U7281 & new_P2_U7282 & new_P2_U7284 & new_P2_U7283;
  assign new_P2_U4305 = new_P2_U7286 & new_P2_U7287 & new_P2_U7289 & new_P2_U7288;
  assign new_P2_U4306 = new_P2_U7290 & new_P2_U7291 & new_P2_U7293 & new_P2_U7292;
  assign new_P2_U4307 = new_P2_U7294 & new_P2_U7295 & new_P2_U7297 & new_P2_U7296;
  assign new_P2_U4308 = new_P2_U7298 & new_P2_U7299 & new_P2_U7301 & new_P2_U7300;
  assign new_P2_U4309 = new_P2_U7303 & new_P2_U7304 & new_P2_U7306 & new_P2_U7305;
  assign new_P2_U4310 = new_P2_U7307 & new_P2_U7308 & new_P2_U7310 & new_P2_U7309;
  assign new_P2_U4311 = new_P2_U7311 & new_P2_U7312 & new_P2_U7314 & new_P2_U7313;
  assign new_P2_U4312 = new_P2_U7315 & new_P2_U7316 & new_P2_U7318 & new_P2_U7317;
  assign new_P2_U4313 = new_P2_U7320 & new_P2_U7321 & new_P2_U7323 & new_P2_U7322;
  assign new_P2_U4314 = new_P2_U7324 & new_P2_U7325 & new_P2_U7327 & new_P2_U7326;
  assign new_P2_U4315 = new_P2_U7328 & new_P2_U7329 & new_P2_U7331 & new_P2_U7330;
  assign new_P2_U4316 = new_P2_U7332 & new_P2_U7333 & new_P2_U7335 & new_P2_U7334;
  assign new_P2_U4317 = new_P2_U7337 & new_P2_U7338 & new_P2_U7340 & new_P2_U7339;
  assign new_P2_U4318 = new_P2_U7341 & new_P2_U7342 & new_P2_U7344 & new_P2_U7343;
  assign new_P2_U4319 = new_P2_U7345 & new_P2_U7346 & new_P2_U7348 & new_P2_U7347;
  assign new_P2_U4320 = new_P2_U7349 & new_P2_U7350 & new_P2_U7352 & new_P2_U7351;
  assign new_P2_U4321 = new_P2_U7354 & new_P2_U7355 & new_P2_U7357 & new_P2_U7356;
  assign new_P2_U4322 = new_P2_U7358 & new_P2_U7359 & new_P2_U7361 & new_P2_U7360;
  assign new_P2_U4323 = new_P2_U7362 & new_P2_U7363 & new_P2_U7365 & new_P2_U7364;
  assign new_P2_U4324 = new_P2_U7366 & new_P2_U7367 & new_P2_U7369 & new_P2_U7368;
  assign new_P2_U4325 = new_P2_U7371 & new_P2_U7372 & new_P2_U7374 & new_P2_U7373;
  assign new_P2_U4326 = new_P2_U7375 & new_P2_U7376 & new_P2_U7378 & new_P2_U7377;
  assign new_P2_U4327 = new_P2_U7379 & new_P2_U7380 & new_P2_U7382 & new_P2_U7381;
  assign new_P2_U4328 = new_P2_U7383 & new_P2_U7384 & new_P2_U7386 & new_P2_U7385;
  assign new_P2_U4329 = new_P2_U7388 & new_P2_U7389 & new_P2_U7391 & new_P2_U7390;
  assign new_P2_U4330 = new_P2_U7392 & new_P2_U7393 & new_P2_U7395 & new_P2_U7394;
  assign new_P2_U4331 = new_P2_U7396 & new_P2_U7397 & new_P2_U7399 & new_P2_U7398;
  assign new_P2_U4332 = new_P2_U7400 & new_P2_U7401 & new_P2_U7403 & new_P2_U7402;
  assign new_P2_U4333 = new_P2_U7405 & new_P2_U7406 & new_P2_U7408 & new_P2_U7407;
  assign new_P2_U4334 = new_P2_U7409 & new_P2_U7410 & new_P2_U7412 & new_P2_U7411;
  assign new_P2_U4335 = new_P2_U7413 & new_P2_U7414 & new_P2_U7416 & new_P2_U7415;
  assign new_P2_U4336 = new_P2_U7417 & new_P2_U7418 & new_P2_U7420 & new_P2_U7419;
  assign new_P2_U4337 = new_P2_U2616 & new_P2_U3300;
  assign new_P2_U4338 = new_P2_U7425 & new_P2_U4413;
  assign new_P2_U4339 = new_P2_U4595 & new_P2_U3300;
  assign new_P2_U4340 = new_P2_U7428 & new_P2_U7426 & new_P2_U4414;
  assign new_P2_U4341 = new_P2_U7430 & new_P2_U3571;
  assign new_P2_U4342 = new_P2_U4413 & new_P2_U4341;
  assign new_P2_U4343 = new_P2_U7869 & new_P2_U7873;
  assign new_P2_U4344 = new_P2_U7436 & new_P2_U7435;
  assign new_P2_U4345 = new_P2_U7440 & new_P2_U7439;
  assign new_P2_U4346 = new_P2_U7442 & new_P2_U7443;
  assign new_P2_U4347 = new_P2_U7445 & new_P2_U7446;
  assign new_P2_U4348 = new_P2_U7448 & new_P2_U7449;
  assign new_P2_U4349 = new_P2_U7451 & new_P2_U7452;
  assign new_P2_U4350 = new_P2_U7454 & new_P2_U7455;
  assign new_P2_U4351 = new_P2_U7457 & new_P2_U7458;
  assign new_P2_U4352 = new_P2_U7460 & new_P2_U7461;
  assign new_P2_U4353 = new_P2_U7463 & new_P2_U7464;
  assign new_P2_U4354 = new_P2_U7466 & new_P2_U7467;
  assign new_P2_U4355 = new_P2_U7469 & new_P2_U7470;
  assign new_P2_U4356 = new_P2_U7472 & new_P2_U7473;
  assign new_P2_U4357 = new_P2_U7475 & new_P2_U7476;
  assign new_P2_U4358 = new_P2_U7478 & new_P2_U7479;
  assign new_P2_U4359 = new_P2_U7481 & new_P2_U7482;
  assign new_P2_U4360 = new_P2_U7484 & new_P2_U7485;
  assign new_P2_U4361 = new_P2_U7487 & new_P2_U7488;
  assign new_P2_U4362 = new_P2_U7490 & new_P2_U7491;
  assign new_P2_U4363 = new_P2_U7493 & new_P2_U7494;
  assign new_P2_U4364 = new_P2_U7496 & new_P2_U7497;
  assign new_P2_U4365 = new_P2_U7499 & new_P2_U7500;
  assign new_P2_U4366 = new_P2_U7502 & new_P2_U7503;
  assign new_P2_U4367 = new_P2_U7505 & new_P2_U7506;
  assign new_P2_U4368 = new_P2_U7510 & new_P2_U7509;
  assign new_P2_U4369 = new_P2_U7514 & new_P2_U7513;
  assign new_P2_U4370 = new_P2_U7518 & new_P2_U7517;
  assign new_P2_U4371 = new_P2_U7522 & new_P2_U7521;
  assign new_P2_U4372 = new_P2_U7526 & new_P2_U7525;
  assign new_P2_U4373 = new_P2_U7530 & new_P2_U7529;
  assign new_P2_U4374 = new_P2_U7532 & new_P2_U7533;
  assign new_P2_U4375 = new_P2_U7536 & new_P2_U7535;
  assign new_P2_U4376 = new_P2_U3255 & new_P2_U6845;
  assign new_P2_U4377 = new_P2_U7863 & new_P2_U3255;
  assign new_P2_U4378 = new_P2_U2356 & new_P2_U7873;
  assign new_P2_U4379 = new_P2_U7578 & new_P2_U7579 & new_P2_U7580;
  assign new_P2_U4380 = new_P2_U7585 & new_P2_U3269;
  assign new_P2_U4381 = new_P2_U2356 & new_P2_U4595;
  assign new_P2_U4382 = new_P2_U7586 & new_P2_U7587 & new_P2_U4472 & new_P2_U3577 & new_P2_U3539;
  assign new_P2_U4383 = new_P2_U7579 & new_P2_U4422;
  assign new_P2_U4384 = new_P2_U4383 & new_P2_U7578;
  assign new_P2_U4385 = new_P2_U7580 & new_P2_U4458;
  assign new_P2_U4386 = new_P2_U7590 & new_P2_U7589;
  assign new_P2_U4387 = P2_STATE2_REG_0_ & new_P2_U7736;
  assign new_P2_U4388 = new_P2_U3549 & new_P2_U4457 & new_P2_U3573 & new_P2_U4458;
  assign new_P2_U4389 = new_P2_U7719 & new_P2_U7718;
  assign new_P2_U4390 = new_P2_U7731 & new_P2_U3536;
  assign new_P2_U4391 = new_P2_U7735 & new_P2_U3536;
  assign new_P2_U4392 = new_P2_U7908 & new_P2_U7907;
  assign new_P2_U4393 = new_P2_U8055 & new_P2_U8054;
  assign new_P2_U4394 = ~new_P2_U3872 | ~new_P2_U5582;
  assign new_P2_U4395 = new_P2_U8079 & new_P2_U8078;
  assign new_P2_U4396 = new_P2_U8092 & new_P2_U8091;
  assign new_P2_U4397 = new_P2_U8120 & new_P2_U8119;
  assign new_P2_U4398 = new_P2_U8126 & new_P2_U8125;
  assign new_P2_U4399 = new_P2_U8132 & new_P2_U8131;
  assign new_P2_U4400 = ~new_P2_U2374 | ~new_P2_U3291;
  assign new_P2_U4401 = ~BS16;
  assign new_P2_U4402 = ~new_P2_U4462 | ~new_P2_U4188;
  assign new_P2_U4403 = ~new_P2_U3534 | ~new_P2_U4462;
  assign new_P2_U4404 = new_P2_U8146 & new_P2_U8145;
  assign new_P2_U4405 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U7006;
  assign new_P2_U4406 = ~new_P2_U2513 | ~new_P2_U3871;
  assign new_P2_U4407 = ~new_P2_R2219_U29;
  assign new_P2_U4408 = ~new_P2_R2219_U8;
  assign new_P2_U4409 = ~new_P2_U3553;
  assign new_P2_U4410 = ~HOLD | ~new_P2_U3265;
  assign new_P2_U4411 = ~new_P2_U3290;
  assign new_P2_U4412 = ~new_P2_U3571;
  assign new_P2_U4413 = ~new_P2_U4337 | ~new_P2_U4601;
  assign new_P2_U4414 = ~new_P2_U7869 | ~new_P2_U2616 | ~new_P2_U3300;
  assign new_P2_U4415 = ~new_P2_U2447 | ~new_P2_U3279;
  assign new_P2_U4416 = ~new_P2_U3576;
  assign new_P2_U4417 = ~new_P2_U3283;
  assign new_P2_U4418 = ~new_P2_U3550;
  assign new_P2_U4419 = ~new_P2_U3536;
  assign new_P2_U4420 = ~new_P2_U3288;
  assign new_P2_U4421 = ~new_P2_U3539;
  assign new_P2_U4422 = ~new_P2_U2450 | ~new_P2_U2376 | ~new_P2_U3278;
  assign new_P2_U4423 = ~new_P2_U3577;
  assign new_P2_U4424 = ~new_P2_U3282;
  assign new_P2_U4425 = ~new_P2_U3285;
  assign new_P2_U4426 = ~new_P2_U3549;
  assign new_P2_U4427 = ~new_P2_U3289;
  assign new_P2_U4428 = ~new_P2_U3286;
  assign new_P2_U4429 = ~new_P2_U3294;
  assign new_P2_U4430 = ~new_P2_U3313;
  assign new_P2_U4431 = ~new_P2_U3578;
  assign new_P2_U4432 = ~new_P2_U3254;
  assign new_P2_U4433 = ~new_P2_U3523;
  assign new_P2_U4434 = ~new_P2_U3524;
  assign new_P2_U4435 = ~new_P2_U3296;
  assign new_P2_U4436 = ~new_P2_U3522;
  assign new_P2_U4437 = ~new_P2_U3875 | ~new_P2_U2376;
  assign new_P2_U4438 = ~new_P2_U3547;
  assign new_P2_U4439 = ~new_P2_U3259;
  assign new_P2_U4440 = ~new_P2_U3543;
  assign new_P2_U4441 = ~new_P2_U3542;
  assign new_P2_U4442 = ~new_P2_U3538;
  assign new_P2_U4443 = ~new_P2_U3306;
  assign new_P2_U4444 = ~new_P2_LT_563_1260_U6;
  assign new_P2_U4445 = ~new_P2_U4430 | ~new_P2_U3302;
  assign new_P2_U4446 = ~new_P2_U4461 | ~new_P2_U3546;
  assign new_P2_U4447 = ~new_P2_R2219_U7 | ~new_P2_U2617;
  assign new_P2_U4448 = ~new_P2_U2367 | ~new_P2_U3290;
  assign new_P2_U4449 = ~new_P2_U3261;
  assign new_P2_U4450 = ~new_P2_U3260;
  assign new_P2_U4451 = ~new_P2_U3425;
  assign new_P2_U4452 = ~new_P2_U4182 | ~new_P2_U4438;
  assign new_P2_U4453 = ~new_P2_U3718 | ~new_P2_U4474;
  assign new_P2_U4454 = ~new_P2_U3284 | ~new_P2_U3270 | ~P2_STATE2_REG_1_ | ~new_P2_U3302;
  assign new_P2_U4455 = ~new_P2_U3867 | ~new_P2_U2448;
  assign new_P2_U4456 = ~new_P2_U2446 | ~new_P2_U2359;
  assign new_P2_U4457 = ~new_P2_U2356 | ~new_P2_U3280;
  assign new_P2_U4458 = ~new_P2_U4378 | ~new_P2_U7577;
  assign new_P2_U4459 = ~new_P2_U3575;
  assign new_P2_U4460 = ~new_P2_U2438 | ~new_P2_U3295;
  assign new_P2_U4461 = ~new_P2_U3534;
  assign new_P2_U4462 = ~new_P2_U2374 | ~new_P2_U6568;
  assign new_P2_U4463 = ~new_P2_U4574 | ~new_P2_U3266;
  assign new_P2_U4464 = ~new_P2_U2448 | ~new_P2_U3292;
  assign new_P2_U4465 = ~new_P2_U4474 | ~new_U211;
  assign new_P2_U4466 = ~new_P2_U3303;
  assign new_P2_U4467 = ~new_P2_U3540;
  assign new_P2_U4468 = ~new_P2_U3304;
  assign new_P2_U4469 = ~new_P2_U3305;
  assign new_P2_U4470 = ~new_P2_U3876 | ~new_P2_U2376;
  assign new_P2_U4471 = ~new_P2_U3573;
  assign new_P2_U4472 = ~new_P2_U4416 | ~new_P2_U2376 | ~new_P2_U7871;
  assign new_P2_U4473 = ~new_P2_U3262;
  assign new_P2_U4474 = ~new_P2_U3301;
  assign new_P2_U4475 = ~new_P2_U3293;
  assign new_P2_U4476 = ~new_P2_U3281;
  assign new_P2_U4477 = ~new_P2_U3548;
  assign new_P2_U4478 = ~P2_REIP_REG_31_ | ~new_P2_U4450;
  assign new_P2_U4479 = ~P2_REIP_REG_30_ | ~new_P2_U4449;
  assign new_P2_U4480 = ~P2_ADDRESS_REG_29_ | ~new_P2_U3259;
  assign new_P2_U4481 = ~P2_REIP_REG_30_ | ~new_P2_U4450;
  assign new_P2_U4482 = ~P2_REIP_REG_29_ | ~new_P2_U4449;
  assign new_P2_U4483 = ~P2_ADDRESS_REG_28_ | ~new_P2_U3259;
  assign new_P2_U4484 = ~P2_REIP_REG_29_ | ~new_P2_U4450;
  assign new_P2_U4485 = ~P2_REIP_REG_28_ | ~new_P2_U4449;
  assign new_P2_U4486 = ~P2_ADDRESS_REG_27_ | ~new_P2_U3259;
  assign new_P2_U4487 = ~P2_REIP_REG_28_ | ~new_P2_U4450;
  assign new_P2_U4488 = ~P2_REIP_REG_27_ | ~new_P2_U4449;
  assign new_P2_U4489 = ~P2_ADDRESS_REG_26_ | ~new_P2_U3259;
  assign new_P2_U4490 = ~P2_REIP_REG_27_ | ~new_P2_U4450;
  assign new_P2_U4491 = ~P2_REIP_REG_26_ | ~new_P2_U4449;
  assign new_P2_U4492 = ~P2_ADDRESS_REG_25_ | ~new_P2_U3259;
  assign new_P2_U4493 = ~P2_REIP_REG_26_ | ~new_P2_U4450;
  assign new_P2_U4494 = ~P2_REIP_REG_25_ | ~new_P2_U4449;
  assign new_P2_U4495 = ~P2_ADDRESS_REG_24_ | ~new_P2_U3259;
  assign new_P2_U4496 = ~P2_REIP_REG_25_ | ~new_P2_U4450;
  assign new_P2_U4497 = ~P2_REIP_REG_24_ | ~new_P2_U4449;
  assign new_P2_U4498 = ~P2_ADDRESS_REG_23_ | ~new_P2_U3259;
  assign new_P2_U4499 = ~P2_REIP_REG_24_ | ~new_P2_U4450;
  assign new_P2_U4500 = ~P2_REIP_REG_23_ | ~new_P2_U4449;
  assign new_P2_U4501 = ~P2_ADDRESS_REG_22_ | ~new_P2_U3259;
  assign new_P2_U4502 = ~P2_REIP_REG_23_ | ~new_P2_U4450;
  assign new_P2_U4503 = ~P2_REIP_REG_22_ | ~new_P2_U4449;
  assign new_P2_U4504 = ~P2_ADDRESS_REG_21_ | ~new_P2_U3259;
  assign new_P2_U4505 = ~P2_REIP_REG_22_ | ~new_P2_U4450;
  assign new_P2_U4506 = ~P2_REIP_REG_21_ | ~new_P2_U4449;
  assign new_P2_U4507 = ~P2_ADDRESS_REG_20_ | ~new_P2_U3259;
  assign new_P2_U4508 = ~P2_REIP_REG_21_ | ~new_P2_U4450;
  assign new_P2_U4509 = ~P2_REIP_REG_20_ | ~new_P2_U4449;
  assign new_P2_U4510 = ~P2_ADDRESS_REG_19_ | ~new_P2_U3259;
  assign new_P2_U4511 = ~P2_REIP_REG_20_ | ~new_P2_U4450;
  assign new_P2_U4512 = ~P2_REIP_REG_19_ | ~new_P2_U4449;
  assign new_P2_U4513 = ~P2_ADDRESS_REG_18_ | ~new_P2_U3259;
  assign new_P2_U4514 = ~P2_REIP_REG_19_ | ~new_P2_U4450;
  assign new_P2_U4515 = ~P2_REIP_REG_18_ | ~new_P2_U4449;
  assign new_P2_U4516 = ~P2_ADDRESS_REG_17_ | ~new_P2_U3259;
  assign new_P2_U4517 = ~P2_REIP_REG_18_ | ~new_P2_U4450;
  assign new_P2_U4518 = ~P2_REIP_REG_17_ | ~new_P2_U4449;
  assign new_P2_U4519 = ~P2_ADDRESS_REG_16_ | ~new_P2_U3259;
  assign new_P2_U4520 = ~P2_REIP_REG_17_ | ~new_P2_U4450;
  assign new_P2_U4521 = ~P2_REIP_REG_16_ | ~new_P2_U4449;
  assign new_P2_U4522 = ~P2_ADDRESS_REG_15_ | ~new_P2_U3259;
  assign new_P2_U4523 = ~P2_REIP_REG_16_ | ~new_P2_U4450;
  assign new_P2_U4524 = ~P2_REIP_REG_15_ | ~new_P2_U4449;
  assign new_P2_U4525 = ~P2_ADDRESS_REG_14_ | ~new_P2_U3259;
  assign new_P2_U4526 = ~P2_REIP_REG_15_ | ~new_P2_U4450;
  assign new_P2_U4527 = ~P2_REIP_REG_14_ | ~new_P2_U4449;
  assign new_P2_U4528 = ~P2_ADDRESS_REG_13_ | ~new_P2_U3259;
  assign new_P2_U4529 = ~P2_REIP_REG_14_ | ~new_P2_U4450;
  assign new_P2_U4530 = ~P2_REIP_REG_13_ | ~new_P2_U4449;
  assign new_P2_U4531 = ~P2_ADDRESS_REG_12_ | ~new_P2_U3259;
  assign new_P2_U4532 = ~P2_REIP_REG_13_ | ~new_P2_U4450;
  assign new_P2_U4533 = ~P2_REIP_REG_12_ | ~new_P2_U4449;
  assign new_P2_U4534 = ~P2_ADDRESS_REG_11_ | ~new_P2_U3259;
  assign new_P2_U4535 = ~P2_REIP_REG_12_ | ~new_P2_U4450;
  assign new_P2_U4536 = ~P2_REIP_REG_11_ | ~new_P2_U4449;
  assign new_P2_U4537 = ~P2_ADDRESS_REG_10_ | ~new_P2_U3259;
  assign new_P2_U4538 = ~P2_REIP_REG_11_ | ~new_P2_U4450;
  assign new_P2_U4539 = ~P2_REIP_REG_10_ | ~new_P2_U4449;
  assign new_P2_U4540 = ~P2_ADDRESS_REG_9_ | ~new_P2_U3259;
  assign new_P2_U4541 = ~P2_REIP_REG_10_ | ~new_P2_U4450;
  assign new_P2_U4542 = ~P2_REIP_REG_9_ | ~new_P2_U4449;
  assign new_P2_U4543 = ~P2_ADDRESS_REG_8_ | ~new_P2_U3259;
  assign new_P2_U4544 = ~P2_REIP_REG_9_ | ~new_P2_U4450;
  assign new_P2_U4545 = ~P2_REIP_REG_8_ | ~new_P2_U4449;
  assign new_P2_U4546 = ~P2_ADDRESS_REG_7_ | ~new_P2_U3259;
  assign new_P2_U4547 = ~P2_REIP_REG_8_ | ~new_P2_U4450;
  assign new_P2_U4548 = ~P2_REIP_REG_7_ | ~new_P2_U4449;
  assign new_P2_U4549 = ~P2_ADDRESS_REG_6_ | ~new_P2_U3259;
  assign new_P2_U4550 = ~P2_REIP_REG_7_ | ~new_P2_U4450;
  assign new_P2_U4551 = ~P2_REIP_REG_6_ | ~new_P2_U4449;
  assign new_P2_U4552 = ~P2_ADDRESS_REG_5_ | ~new_P2_U3259;
  assign new_P2_U4553 = ~P2_REIP_REG_6_ | ~new_P2_U4450;
  assign new_P2_U4554 = ~P2_REIP_REG_5_ | ~new_P2_U4449;
  assign new_P2_U4555 = ~P2_ADDRESS_REG_4_ | ~new_P2_U3259;
  assign new_P2_U4556 = ~P2_REIP_REG_5_ | ~new_P2_U4450;
  assign new_P2_U4557 = ~P2_REIP_REG_4_ | ~new_P2_U4449;
  assign new_P2_U4558 = ~P2_ADDRESS_REG_3_ | ~new_P2_U3259;
  assign new_P2_U4559 = ~P2_REIP_REG_4_ | ~new_P2_U4450;
  assign new_P2_U4560 = ~P2_REIP_REG_3_ | ~new_P2_U4449;
  assign new_P2_U4561 = ~P2_ADDRESS_REG_2_ | ~new_P2_U3259;
  assign new_P2_U4562 = ~P2_REIP_REG_3_ | ~new_P2_U4450;
  assign new_P2_U4563 = ~P2_REIP_REG_2_ | ~new_P2_U4449;
  assign new_P2_U4564 = ~P2_ADDRESS_REG_1_ | ~new_P2_U3259;
  assign new_P2_U4565 = ~P2_REIP_REG_2_ | ~new_P2_U4450;
  assign new_P2_U4566 = ~P2_REIP_REG_1_ | ~new_P2_U4449;
  assign new_P2_U4567 = ~P2_ADDRESS_REG_0_ | ~new_P2_U3259;
  assign new_P2_U4568 = ~new_P2_U3267;
  assign new_P2_U4569 = ~new_P2_U4568 | ~new_P2_U3265;
  assign new_P2_U4570 = ~NA | ~new_P2_U4473;
  assign new_P2_U4571 = ~new_P2_U3268;
  assign new_P2_U4572 = ~new_P2_U4571 | ~new_P2_U3265;
  assign new_P2_U4573 = ~new_P2_U4392 | ~new_P2_U7891;
  assign new_P2_U4574 = ~new_P2_U3263;
  assign new_P2_U4575 = ~new_P2_U4574 | ~HOLD | ~new_P2_U3256;
  assign new_P2_U4576 = ~new_U211 | ~P2_STATE_REG_1_ | ~new_P2_U3268;
  assign new_P2_U4577 = ~new_P2_U4576 | ~new_P2_U4575;
  assign new_P2_U4578 = ~new_P2_U4577 | ~P2_STATE_REG_0_ | ~new_P2_U4570;
  assign new_P2_U4579 = ~P2_STATE_REG_2_ | ~new_P2_U4573;
  assign new_P2_U4580 = ~P2_STATE_REG_0_ | ~new_P2_U4410;
  assign new_P2_U4581 = ~new_P2_U4580 | ~P2_STATE_REG_2_;
  assign new_P2_U4582 = ~new_P2_U7892 | ~new_P2_U7910 | ~new_P2_U7909;
  assign new_P2_U4583 = ~new_U211 | ~new_P2_U4439;
  assign new_P2_U4584 = ~new_P2_U3692 | ~new_P2_U7893;
  assign new_P2_U4585 = ~P2_STATE_REG_2_ | ~new_P2_U3267;
  assign new_P2_U4586 = ~NA | ~new_P2_U3266;
  assign new_P2_U4587 = ~new_P2_U4586 | ~new_P2_U4585;
  assign new_P2_U4588 = ~new_P2_U4587 | ~new_P2_U3258;
  assign new_P2_U4589 = ~new_P2_U4401 | ~new_P2_U3263;
  assign new_P2_U4590 = ~new_P2_U3277;
  assign new_P2_U4591 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U4592 = ~new_P2_U3274;
  assign new_P2_U4593 = ~new_P2_U3275;
  assign new_P2_U4594 = ~P2_STATE_REG_2_ | ~new_P2_U3258;
  assign new_P2_U4595 = ~new_P2_U3262 | ~new_P2_U4594;
  assign new_P2_U4596 = ~new_P2_U3527;
  assign new_P2_U4597 = ~new_P2_U3294 | ~new_P2_U3286;
  assign new_P2_U4598 = ~new_P2_U4597 | ~new_P2_U3265;
  assign new_P2_U4599 = ~new_P2_U2359 | ~new_P2_U3527;
  assign new_P2_U4600 = ~new_P2_U3291;
  assign new_P2_U4601 = ~new_P2_U3295;
  assign new_P2_U4602 = ~new_P2_U4424 | ~new_P2_U3253;
  assign new_P2_U4603 = ~new_P2_U3524 | ~new_P2_U4602;
  assign new_P2_U4604 = ~new_P2_U3523 | ~new_P2_U3522;
  assign new_P2_U4605 = ~new_P2_R2243_U8 | ~new_P2_U4428;
  assign new_P2_U4606 = ~new_P2_U4417 | ~new_P2_U3287;
  assign new_P2_U4607 = ~new_P2_U4606 | ~new_P2_U4605;
  assign new_P2_U4608 = ~new_P2_U4420 | ~new_P2_U4607;
  assign new_P2_U4609 = ~new_P2_U4603 | ~new_P2_U3520;
  assign new_P2_U4610 = ~new_P2_U3257;
  assign new_P2_U4611 = ~new_P2_U4428 | ~new_P2_U3292;
  assign new_P2_U4612 = ~new_P2_GTE_370_U6 | ~new_P2_U4417;
  assign new_P2_U4613 = ~new_P2_U4612 | ~new_P2_U4611;
  assign new_P2_U4614 = ~new_P2_U4420 | ~new_P2_U4613;
  assign new_P2_U4615 = P2_MORE_REG | P2_FLUSH_REG;
  assign new_P2_U4616 = ~new_P2_U3298;
  assign new_P2_U4617 = ~new_P2_U4616 | ~new_P2_U3269;
  assign new_P2_U4618 = ~new_P2_U3711 | ~new_P2_U4425;
  assign new_P2_U4619 = ~new_P2_U3715 | ~new_P2_U8057 | ~new_P2_U8056;
  assign new_P2_U4620 = ~new_P2_U3299;
  assign new_P2_U4621 = ~new_P2_U4474 | ~new_P2_U3265;
  assign new_P2_U4622 = ~P2_STATEBS16_REG | ~new_P2_U3284;
  assign new_P2_U4623 = ~new_P2_U4622 | ~new_P2_U4621;
  assign new_P2_U4624 = ~P2_STATE2_REG_1_ | ~new_P2_U4623;
  assign new_P2_U4625 = ~P2_STATE2_REG_2_ | ~new_P2_U3299;
  assign new_P2_U4626 = ~new_P2_U4619 | ~new_P2_U4465;
  assign new_P2_U4627 = ~new_P2_U3717 | ~new_P2_U4620;
  assign new_P2_U4628 = ~P2_STATE2_REG_1_ | ~new_P2_U4626;
  assign new_P2_U4629 = ~new_P2_U2374 | ~new_P2_U4619;
  assign new_P2_U4630 = ~new_P2_U3719 | ~new_P2_U4469;
  assign new_P2_U4631 = ~new_P2_U4619 | ~new_P2_U4464;
  assign new_P2_U4632 = ~new_P2_U2374 | ~new_P2_U3298;
  assign new_P2_U4633 = ~new_P2_U3337;
  assign new_P2_U4634 = ~new_P2_U3351;
  assign new_P2_U4635 = ~new_P2_U3352;
  assign new_P2_U4636 = ~new_P2_U3319;
  assign new_P2_U4637 = ~new_P2_U3318;
  assign new_P2_U4638 = ~new_P2_U3378;
  assign new_P2_U4639 = ~new_P2_R2182_U76 | ~new_P2_U3318;
  assign new_P2_U4640 = ~new_P2_U3426;
  assign new_P2_U4641 = ~new_P2_U3320;
  assign new_P2_U4642 = ~new_P2_U3311;
  assign new_P2_U4643 = ~new_P2_U3312;
  assign new_P2_U4644 = ~new_P2_U3424;
  assign new_P2_U4645 = ~new_P2_U3376;
  assign new_P2_U4646 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_U3311;
  assign new_P2_U4647 = ~new_P2_U3428;
  assign new_P2_U4648 = ~new_P2_U3349;
  assign new_P2_U4649 = ~new_P2_U3335;
  assign new_P2_U4650 = ~new_P2_U3243;
  assign new_P2_U4651 = ~new_P2_U2440 | ~new_P2_U2444;
  assign new_P2_U4652 = ~new_P2_U3325;
  assign new_P2_U4653 = ~new_P2_U3570;
  assign new_P2_U4654 = ~new_P2_U3326;
  assign new_P2_U4655 = ~P2_STATE2_REG_1_ | ~new_P2_U3270;
  assign new_P2_U4656 = ~new_P2_U3305 | ~new_P2_U4655 | ~new_P2_U3304;
  assign new_P2_U4657 = ~new_P2_U4637 | ~new_P2_U2462;
  assign new_P2_U4658 = ~new_P2_U2468 | ~new_P2_U2362;
  assign new_P2_U4659 = ~new_P2_U4445 | ~new_P2_U4658;
  assign new_P2_U4660 = ~new_P2_U4652 | ~new_P2_U4659;
  assign new_P2_U4661 = ~new_P2_U4654 | ~P2_STATE2_REG_2_;
  assign new_P2_U4662 = ~P2_STATE2_REG_3_ | ~new_P2_U3312;
  assign new_P2_U4663 = ~new_P2_U4660 | ~new_P2_U3722;
  assign new_P2_U4664 = ~new_P2_U2468 | ~new_P2_U2398;
  assign new_P2_U4665 = ~new_P2_U4445 | ~new_P2_U4664;
  assign new_P2_U4666 = ~new_P2_U4665 | ~new_P2_U3325;
  assign new_P2_U4667 = ~P2_STATE2_REG_2_ | ~new_P2_U3326;
  assign new_P2_U4668 = ~new_P2_U4667 | ~new_P2_U4666;
  assign new_P2_U4669 = ~new_P2_U2425 | ~new_P2_U4643;
  assign new_P2_U4670 = ~new_P2_U2422 | ~new_P2_U2463;
  assign new_P2_U4671 = ~new_P2_U2421 | ~new_P2_U4641;
  assign new_P2_U4672 = ~new_P2_U2406 | ~new_P2_U4668;
  assign new_P2_U4673 = ~P2_INSTQUEUE_REG_15__7_ | ~new_P2_U4663;
  assign new_P2_U4674 = ~new_P2_U2426 | ~new_P2_U4643;
  assign new_P2_U4675 = ~new_P2_U2420 | ~new_P2_U2463;
  assign new_P2_U4676 = ~new_P2_U2419 | ~new_P2_U4641;
  assign new_P2_U4677 = ~new_P2_U2405 | ~new_P2_U4668;
  assign new_P2_U4678 = ~P2_INSTQUEUE_REG_15__6_ | ~new_P2_U4663;
  assign new_P2_U4679 = ~new_P2_U2429 | ~new_P2_U4643;
  assign new_P2_U4680 = ~new_P2_U2418 | ~new_P2_U2463;
  assign new_P2_U4681 = ~new_P2_U2417 | ~new_P2_U4641;
  assign new_P2_U4682 = ~new_P2_U2404 | ~new_P2_U4668;
  assign new_P2_U4683 = ~P2_INSTQUEUE_REG_15__5_ | ~new_P2_U4663;
  assign new_P2_U4684 = ~new_P2_U2424 | ~new_P2_U4643;
  assign new_P2_U4685 = ~new_P2_U2416 | ~new_P2_U2463;
  assign new_P2_U4686 = ~new_P2_U2415 | ~new_P2_U4641;
  assign new_P2_U4687 = ~new_P2_U2403 | ~new_P2_U4668;
  assign new_P2_U4688 = ~P2_INSTQUEUE_REG_15__4_ | ~new_P2_U4663;
  assign new_P2_U4689 = ~new_P2_U2423 | ~new_P2_U4643;
  assign new_P2_U4690 = ~new_P2_U2414 | ~new_P2_U2463;
  assign new_P2_U4691 = ~new_P2_U2413 | ~new_P2_U4641;
  assign new_P2_U4692 = ~new_P2_U2402 | ~new_P2_U4668;
  assign new_P2_U4693 = ~P2_INSTQUEUE_REG_15__3_ | ~new_P2_U4663;
  assign new_P2_U4694 = ~new_P2_U2432 | ~new_P2_U4643;
  assign new_P2_U4695 = ~new_P2_U2412 | ~new_P2_U2463;
  assign new_P2_U4696 = ~new_P2_U2411 | ~new_P2_U4641;
  assign new_P2_U4697 = ~new_P2_U2401 | ~new_P2_U4668;
  assign new_P2_U4698 = ~P2_INSTQUEUE_REG_15__2_ | ~new_P2_U4663;
  assign new_P2_U4699 = ~new_P2_U2428 | ~new_P2_U4643;
  assign new_P2_U4700 = ~new_P2_U2410 | ~new_P2_U2463;
  assign new_P2_U4701 = ~new_P2_U2409 | ~new_P2_U4641;
  assign new_P2_U4702 = ~new_P2_U2400 | ~new_P2_U4668;
  assign new_P2_U4703 = ~P2_INSTQUEUE_REG_15__1_ | ~new_P2_U4663;
  assign new_P2_U4704 = ~new_P2_U2431 | ~new_P2_U4643;
  assign new_P2_U4705 = ~new_P2_U2408 | ~new_P2_U2463;
  assign new_P2_U4706 = ~new_P2_U2407 | ~new_P2_U4641;
  assign new_P2_U4707 = ~new_P2_U2399 | ~new_P2_U4668;
  assign new_P2_U4708 = ~P2_INSTQUEUE_REG_15__0_ | ~new_P2_U4663;
  assign new_P2_U4709 = ~new_P2_U3338;
  assign new_P2_U4710 = ~new_P2_U3339;
  assign new_P2_U4711 = ~new_P2_U3336;
  assign new_P2_U4712 = ~new_P2_U3245;
  assign new_P2_U4713 = ~new_P2_U3569;
  assign new_P2_U4714 = ~new_P2_U3340;
  assign new_P2_U4715 = ~new_P2_U4633 | ~new_P2_U2462;
  assign new_P2_U4716 = ~new_P2_U2471 | ~new_P2_U2362;
  assign new_P2_U4717 = ~new_P2_U4445 | ~new_P2_U4716;
  assign new_P2_U4718 = ~new_P2_U4717 | ~new_P2_U3245;
  assign new_P2_U4719 = ~new_P2_U4714 | ~P2_STATE2_REG_2_;
  assign new_P2_U4720 = ~P2_STATE2_REG_3_ | ~new_P2_U3336;
  assign new_P2_U4721 = ~new_P2_U4718 | ~new_P2_U3731;
  assign new_P2_U4722 = ~new_P2_U2471 | ~new_P2_U2398;
  assign new_P2_U4723 = ~new_P2_U4445 | ~new_P2_U4722;
  assign new_P2_U4724 = ~new_P2_U4723 | ~new_P2_U4712;
  assign new_P2_U4725 = ~P2_STATE2_REG_2_ | ~new_P2_U3340;
  assign new_P2_U4726 = ~new_P2_U4725 | ~new_P2_U4724;
  assign new_P2_U4727 = ~new_P2_U4711 | ~new_P2_U2425;
  assign new_P2_U4728 = ~new_P2_U2469 | ~new_P2_U2422;
  assign new_P2_U4729 = ~new_P2_U4710 | ~new_P2_U2421;
  assign new_P2_U4730 = ~new_P2_U2406 | ~new_P2_U4726;
  assign new_P2_U4731 = ~P2_INSTQUEUE_REG_14__7_ | ~new_P2_U4721;
  assign new_P2_U4732 = ~new_P2_U4711 | ~new_P2_U2426;
  assign new_P2_U4733 = ~new_P2_U2469 | ~new_P2_U2420;
  assign new_P2_U4734 = ~new_P2_U4710 | ~new_P2_U2419;
  assign new_P2_U4735 = ~new_P2_U2405 | ~new_P2_U4726;
  assign new_P2_U4736 = ~P2_INSTQUEUE_REG_14__6_ | ~new_P2_U4721;
  assign new_P2_U4737 = ~new_P2_U4711 | ~new_P2_U2429;
  assign new_P2_U4738 = ~new_P2_U2469 | ~new_P2_U2418;
  assign new_P2_U4739 = ~new_P2_U4710 | ~new_P2_U2417;
  assign new_P2_U4740 = ~new_P2_U2404 | ~new_P2_U4726;
  assign new_P2_U4741 = ~P2_INSTQUEUE_REG_14__5_ | ~new_P2_U4721;
  assign new_P2_U4742 = ~new_P2_U4711 | ~new_P2_U2424;
  assign new_P2_U4743 = ~new_P2_U2469 | ~new_P2_U2416;
  assign new_P2_U4744 = ~new_P2_U4710 | ~new_P2_U2415;
  assign new_P2_U4745 = ~new_P2_U2403 | ~new_P2_U4726;
  assign new_P2_U4746 = ~P2_INSTQUEUE_REG_14__4_ | ~new_P2_U4721;
  assign new_P2_U4747 = ~new_P2_U4711 | ~new_P2_U2423;
  assign new_P2_U4748 = ~new_P2_U2469 | ~new_P2_U2414;
  assign new_P2_U4749 = ~new_P2_U4710 | ~new_P2_U2413;
  assign new_P2_U4750 = ~new_P2_U2402 | ~new_P2_U4726;
  assign new_P2_U4751 = ~P2_INSTQUEUE_REG_14__3_ | ~new_P2_U4721;
  assign new_P2_U4752 = ~new_P2_U4711 | ~new_P2_U2432;
  assign new_P2_U4753 = ~new_P2_U2469 | ~new_P2_U2412;
  assign new_P2_U4754 = ~new_P2_U4710 | ~new_P2_U2411;
  assign new_P2_U4755 = ~new_P2_U2401 | ~new_P2_U4726;
  assign new_P2_U4756 = ~P2_INSTQUEUE_REG_14__2_ | ~new_P2_U4721;
  assign new_P2_U4757 = ~new_P2_U4711 | ~new_P2_U2428;
  assign new_P2_U4758 = ~new_P2_U2469 | ~new_P2_U2410;
  assign new_P2_U4759 = ~new_P2_U4710 | ~new_P2_U2409;
  assign new_P2_U4760 = ~new_P2_U2400 | ~new_P2_U4726;
  assign new_P2_U4761 = ~P2_INSTQUEUE_REG_14__1_ | ~new_P2_U4721;
  assign new_P2_U4762 = ~new_P2_U4711 | ~new_P2_U2431;
  assign new_P2_U4763 = ~new_P2_U2469 | ~new_P2_U2408;
  assign new_P2_U4764 = ~new_P2_U4710 | ~new_P2_U2407;
  assign new_P2_U4765 = ~new_P2_U2399 | ~new_P2_U4726;
  assign new_P2_U4766 = ~P2_INSTQUEUE_REG_14__0_ | ~new_P2_U4721;
  assign new_P2_U4767 = ~new_P2_U3353;
  assign new_P2_U4768 = ~new_P2_U3354;
  assign new_P2_U4769 = ~new_P2_U3350;
  assign new_P2_U4770 = ~new_P2_U2445 | ~new_P2_U2440;
  assign new_P2_U4771 = ~new_P2_U3355;
  assign new_P2_U4772 = ~new_P2_U3568;
  assign new_P2_U4773 = ~new_P2_U3356;
  assign new_P2_U4774 = ~new_P2_U4634 | ~new_P2_U2462;
  assign new_P2_U4775 = ~new_P2_U2474 | ~new_P2_U2362;
  assign new_P2_U4776 = ~new_P2_U4445 | ~new_P2_U4775;
  assign new_P2_U4777 = ~new_P2_U4771 | ~new_P2_U4776;
  assign new_P2_U4778 = ~new_P2_U4773 | ~P2_STATE2_REG_2_;
  assign new_P2_U4779 = ~P2_STATE2_REG_3_ | ~new_P2_U3350;
  assign new_P2_U4780 = ~new_P2_U4777 | ~new_P2_U3740;
  assign new_P2_U4781 = ~new_P2_U2474 | ~new_P2_U2398;
  assign new_P2_U4782 = ~new_P2_U4445 | ~new_P2_U4781;
  assign new_P2_U4783 = ~new_P2_U4782 | ~new_P2_U3355;
  assign new_P2_U4784 = ~P2_STATE2_REG_2_ | ~new_P2_U3356;
  assign new_P2_U4785 = ~new_P2_U4784 | ~new_P2_U4783;
  assign new_P2_U4786 = ~new_P2_U4769 | ~new_P2_U2425;
  assign new_P2_U4787 = ~new_P2_U2472 | ~new_P2_U2422;
  assign new_P2_U4788 = ~new_P2_U4768 | ~new_P2_U2421;
  assign new_P2_U4789 = ~new_P2_U2406 | ~new_P2_U4785;
  assign new_P2_U4790 = ~P2_INSTQUEUE_REG_13__7_ | ~new_P2_U4780;
  assign new_P2_U4791 = ~new_P2_U4769 | ~new_P2_U2426;
  assign new_P2_U4792 = ~new_P2_U2472 | ~new_P2_U2420;
  assign new_P2_U4793 = ~new_P2_U4768 | ~new_P2_U2419;
  assign new_P2_U4794 = ~new_P2_U2405 | ~new_P2_U4785;
  assign new_P2_U4795 = ~P2_INSTQUEUE_REG_13__6_ | ~new_P2_U4780;
  assign new_P2_U4796 = ~new_P2_U4769 | ~new_P2_U2429;
  assign new_P2_U4797 = ~new_P2_U2472 | ~new_P2_U2418;
  assign new_P2_U4798 = ~new_P2_U4768 | ~new_P2_U2417;
  assign new_P2_U4799 = ~new_P2_U2404 | ~new_P2_U4785;
  assign new_P2_U4800 = ~P2_INSTQUEUE_REG_13__5_ | ~new_P2_U4780;
  assign new_P2_U4801 = ~new_P2_U4769 | ~new_P2_U2424;
  assign new_P2_U4802 = ~new_P2_U2472 | ~new_P2_U2416;
  assign new_P2_U4803 = ~new_P2_U4768 | ~new_P2_U2415;
  assign new_P2_U4804 = ~new_P2_U2403 | ~new_P2_U4785;
  assign new_P2_U4805 = ~P2_INSTQUEUE_REG_13__4_ | ~new_P2_U4780;
  assign new_P2_U4806 = ~new_P2_U4769 | ~new_P2_U2423;
  assign new_P2_U4807 = ~new_P2_U2472 | ~new_P2_U2414;
  assign new_P2_U4808 = ~new_P2_U4768 | ~new_P2_U2413;
  assign new_P2_U4809 = ~new_P2_U2402 | ~new_P2_U4785;
  assign new_P2_U4810 = ~P2_INSTQUEUE_REG_13__3_ | ~new_P2_U4780;
  assign new_P2_U4811 = ~new_P2_U4769 | ~new_P2_U2432;
  assign new_P2_U4812 = ~new_P2_U2472 | ~new_P2_U2412;
  assign new_P2_U4813 = ~new_P2_U4768 | ~new_P2_U2411;
  assign new_P2_U4814 = ~new_P2_U2401 | ~new_P2_U4785;
  assign new_P2_U4815 = ~P2_INSTQUEUE_REG_13__2_ | ~new_P2_U4780;
  assign new_P2_U4816 = ~new_P2_U4769 | ~new_P2_U2428;
  assign new_P2_U4817 = ~new_P2_U2472 | ~new_P2_U2410;
  assign new_P2_U4818 = ~new_P2_U4768 | ~new_P2_U2409;
  assign new_P2_U4819 = ~new_P2_U2400 | ~new_P2_U4785;
  assign new_P2_U4820 = ~P2_INSTQUEUE_REG_13__1_ | ~new_P2_U4780;
  assign new_P2_U4821 = ~new_P2_U4769 | ~new_P2_U2431;
  assign new_P2_U4822 = ~new_P2_U2472 | ~new_P2_U2408;
  assign new_P2_U4823 = ~new_P2_U4768 | ~new_P2_U2407;
  assign new_P2_U4824 = ~new_P2_U2399 | ~new_P2_U4785;
  assign new_P2_U4825 = ~P2_INSTQUEUE_REG_13__0_ | ~new_P2_U4780;
  assign new_P2_U4826 = ~new_P2_U3366;
  assign new_P2_U4827 = ~new_P2_U3365;
  assign new_P2_U4828 = ~new_P2_U3246;
  assign new_P2_U4829 = ~new_P2_U3567;
  assign new_P2_U4830 = ~new_P2_U3367;
  assign new_P2_U4831 = ~new_P2_U2476 | ~new_P2_U2462;
  assign new_P2_U4832 = ~new_P2_U2480 | ~new_P2_U2362;
  assign new_P2_U4833 = ~new_P2_U4445 | ~new_P2_U4832;
  assign new_P2_U4834 = ~new_P2_U4833 | ~new_P2_U3246;
  assign new_P2_U4835 = ~new_P2_U4830 | ~P2_STATE2_REG_2_;
  assign new_P2_U4836 = ~P2_STATE2_REG_3_ | ~new_P2_U3365;
  assign new_P2_U4837 = ~new_P2_U4834 | ~new_P2_U3749;
  assign new_P2_U4838 = ~new_P2_U2480 | ~new_P2_U2398;
  assign new_P2_U4839 = ~new_P2_U4445 | ~new_P2_U4838;
  assign new_P2_U4840 = ~new_P2_U4839 | ~new_P2_U4828;
  assign new_P2_U4841 = ~P2_STATE2_REG_2_ | ~new_P2_U3367;
  assign new_P2_U4842 = ~new_P2_U4841 | ~new_P2_U4840;
  assign new_P2_U4843 = ~new_P2_U4827 | ~new_P2_U2425;
  assign new_P2_U4844 = ~new_P2_U2477 | ~new_P2_U2422;
  assign new_P2_U4845 = ~new_P2_U4826 | ~new_P2_U2421;
  assign new_P2_U4846 = ~new_P2_U2406 | ~new_P2_U4842;
  assign new_P2_U4847 = ~P2_INSTQUEUE_REG_12__7_ | ~new_P2_U4837;
  assign new_P2_U4848 = ~new_P2_U4827 | ~new_P2_U2426;
  assign new_P2_U4849 = ~new_P2_U2477 | ~new_P2_U2420;
  assign new_P2_U4850 = ~new_P2_U4826 | ~new_P2_U2419;
  assign new_P2_U4851 = ~new_P2_U2405 | ~new_P2_U4842;
  assign new_P2_U4852 = ~P2_INSTQUEUE_REG_12__6_ | ~new_P2_U4837;
  assign new_P2_U4853 = ~new_P2_U4827 | ~new_P2_U2429;
  assign new_P2_U4854 = ~new_P2_U2477 | ~new_P2_U2418;
  assign new_P2_U4855 = ~new_P2_U4826 | ~new_P2_U2417;
  assign new_P2_U4856 = ~new_P2_U2404 | ~new_P2_U4842;
  assign new_P2_U4857 = ~P2_INSTQUEUE_REG_12__5_ | ~new_P2_U4837;
  assign new_P2_U4858 = ~new_P2_U4827 | ~new_P2_U2424;
  assign new_P2_U4859 = ~new_P2_U2477 | ~new_P2_U2416;
  assign new_P2_U4860 = ~new_P2_U4826 | ~new_P2_U2415;
  assign new_P2_U4861 = ~new_P2_U2403 | ~new_P2_U4842;
  assign new_P2_U4862 = ~P2_INSTQUEUE_REG_12__4_ | ~new_P2_U4837;
  assign new_P2_U4863 = ~new_P2_U4827 | ~new_P2_U2423;
  assign new_P2_U4864 = ~new_P2_U2477 | ~new_P2_U2414;
  assign new_P2_U4865 = ~new_P2_U4826 | ~new_P2_U2413;
  assign new_P2_U4866 = ~new_P2_U2402 | ~new_P2_U4842;
  assign new_P2_U4867 = ~P2_INSTQUEUE_REG_12__3_ | ~new_P2_U4837;
  assign new_P2_U4868 = ~new_P2_U4827 | ~new_P2_U2432;
  assign new_P2_U4869 = ~new_P2_U2477 | ~new_P2_U2412;
  assign new_P2_U4870 = ~new_P2_U4826 | ~new_P2_U2411;
  assign new_P2_U4871 = ~new_P2_U2401 | ~new_P2_U4842;
  assign new_P2_U4872 = ~P2_INSTQUEUE_REG_12__2_ | ~new_P2_U4837;
  assign new_P2_U4873 = ~new_P2_U4827 | ~new_P2_U2428;
  assign new_P2_U4874 = ~new_P2_U2477 | ~new_P2_U2410;
  assign new_P2_U4875 = ~new_P2_U4826 | ~new_P2_U2409;
  assign new_P2_U4876 = ~new_P2_U2400 | ~new_P2_U4842;
  assign new_P2_U4877 = ~P2_INSTQUEUE_REG_12__1_ | ~new_P2_U4837;
  assign new_P2_U4878 = ~new_P2_U4827 | ~new_P2_U2431;
  assign new_P2_U4879 = ~new_P2_U2477 | ~new_P2_U2408;
  assign new_P2_U4880 = ~new_P2_U4826 | ~new_P2_U2407;
  assign new_P2_U4881 = ~new_P2_U2399 | ~new_P2_U4842;
  assign new_P2_U4882 = ~P2_INSTQUEUE_REG_12__0_ | ~new_P2_U4837;
  assign new_P2_U4883 = ~new_P2_U3379;
  assign new_P2_U4884 = ~new_P2_U3377;
  assign new_P2_U4885 = ~new_P2_U2442 | ~new_P2_U2444;
  assign new_P2_U4886 = ~new_P2_U3380;
  assign new_P2_U4887 = ~new_P2_U3566;
  assign new_P2_U4888 = ~new_P2_U3381;
  assign new_P2_U4889 = ~new_P2_U4638 | ~new_P2_U4637;
  assign new_P2_U4890 = ~new_P2_U2484 | ~new_P2_U2362;
  assign new_P2_U4891 = ~new_P2_U4445 | ~new_P2_U4890;
  assign new_P2_U4892 = ~new_P2_U4886 | ~new_P2_U4891;
  assign new_P2_U4893 = ~new_P2_U4888 | ~P2_STATE2_REG_2_;
  assign new_P2_U4894 = ~P2_STATE2_REG_3_ | ~new_P2_U3377;
  assign new_P2_U4895 = ~new_P2_U4892 | ~new_P2_U3758;
  assign new_P2_U4896 = ~new_P2_U2484 | ~new_P2_U2398;
  assign new_P2_U4897 = ~new_P2_U4445 | ~new_P2_U4896;
  assign new_P2_U4898 = ~new_P2_U4897 | ~new_P2_U3380;
  assign new_P2_U4899 = ~P2_STATE2_REG_2_ | ~new_P2_U3381;
  assign new_P2_U4900 = ~new_P2_U4899 | ~new_P2_U4898;
  assign new_P2_U4901 = ~new_P2_U4884 | ~new_P2_U2425;
  assign new_P2_U4902 = ~new_P2_U2482 | ~new_P2_U2422;
  assign new_P2_U4903 = ~new_P2_U4883 | ~new_P2_U2421;
  assign new_P2_U4904 = ~new_P2_U2406 | ~new_P2_U4900;
  assign new_P2_U4905 = ~P2_INSTQUEUE_REG_11__7_ | ~new_P2_U4895;
  assign new_P2_U4906 = ~new_P2_U4884 | ~new_P2_U2426;
  assign new_P2_U4907 = ~new_P2_U2482 | ~new_P2_U2420;
  assign new_P2_U4908 = ~new_P2_U4883 | ~new_P2_U2419;
  assign new_P2_U4909 = ~new_P2_U2405 | ~new_P2_U4900;
  assign new_P2_U4910 = ~P2_INSTQUEUE_REG_11__6_ | ~new_P2_U4895;
  assign new_P2_U4911 = ~new_P2_U4884 | ~new_P2_U2429;
  assign new_P2_U4912 = ~new_P2_U2482 | ~new_P2_U2418;
  assign new_P2_U4913 = ~new_P2_U4883 | ~new_P2_U2417;
  assign new_P2_U4914 = ~new_P2_U2404 | ~new_P2_U4900;
  assign new_P2_U4915 = ~P2_INSTQUEUE_REG_11__5_ | ~new_P2_U4895;
  assign new_P2_U4916 = ~new_P2_U4884 | ~new_P2_U2424;
  assign new_P2_U4917 = ~new_P2_U2482 | ~new_P2_U2416;
  assign new_P2_U4918 = ~new_P2_U4883 | ~new_P2_U2415;
  assign new_P2_U4919 = ~new_P2_U2403 | ~new_P2_U4900;
  assign new_P2_U4920 = ~P2_INSTQUEUE_REG_11__4_ | ~new_P2_U4895;
  assign new_P2_U4921 = ~new_P2_U4884 | ~new_P2_U2423;
  assign new_P2_U4922 = ~new_P2_U2482 | ~new_P2_U2414;
  assign new_P2_U4923 = ~new_P2_U4883 | ~new_P2_U2413;
  assign new_P2_U4924 = ~new_P2_U2402 | ~new_P2_U4900;
  assign new_P2_U4925 = ~P2_INSTQUEUE_REG_11__3_ | ~new_P2_U4895;
  assign new_P2_U4926 = ~new_P2_U4884 | ~new_P2_U2432;
  assign new_P2_U4927 = ~new_P2_U2482 | ~new_P2_U2412;
  assign new_P2_U4928 = ~new_P2_U4883 | ~new_P2_U2411;
  assign new_P2_U4929 = ~new_P2_U2401 | ~new_P2_U4900;
  assign new_P2_U4930 = ~P2_INSTQUEUE_REG_11__2_ | ~new_P2_U4895;
  assign new_P2_U4931 = ~new_P2_U4884 | ~new_P2_U2428;
  assign new_P2_U4932 = ~new_P2_U2482 | ~new_P2_U2410;
  assign new_P2_U4933 = ~new_P2_U4883 | ~new_P2_U2409;
  assign new_P2_U4934 = ~new_P2_U2400 | ~new_P2_U4900;
  assign new_P2_U4935 = ~P2_INSTQUEUE_REG_11__1_ | ~new_P2_U4895;
  assign new_P2_U4936 = ~new_P2_U4884 | ~new_P2_U2431;
  assign new_P2_U4937 = ~new_P2_U2482 | ~new_P2_U2408;
  assign new_P2_U4938 = ~new_P2_U4883 | ~new_P2_U2407;
  assign new_P2_U4939 = ~new_P2_U2399 | ~new_P2_U4900;
  assign new_P2_U4940 = ~P2_INSTQUEUE_REG_11__0_ | ~new_P2_U4895;
  assign new_P2_U4941 = ~new_P2_U3391;
  assign new_P2_U4942 = ~new_P2_U3390;
  assign new_P2_U4943 = ~new_P2_U3247;
  assign new_P2_U4944 = ~new_P2_U3565;
  assign new_P2_U4945 = ~new_P2_U3392;
  assign new_P2_U4946 = ~new_P2_U4638 | ~new_P2_U4633;
  assign new_P2_U4947 = ~new_P2_U2486 | ~new_P2_U2362;
  assign new_P2_U4948 = ~new_P2_U4445 | ~new_P2_U4947;
  assign new_P2_U4949 = ~new_P2_U4948 | ~new_P2_U3247;
  assign new_P2_U4950 = ~new_P2_U4945 | ~P2_STATE2_REG_2_;
  assign new_P2_U4951 = ~P2_STATE2_REG_3_ | ~new_P2_U3390;
  assign new_P2_U4952 = ~new_P2_U4949 | ~new_P2_U3767;
  assign new_P2_U4953 = ~new_P2_U2486 | ~new_P2_U2398;
  assign new_P2_U4954 = ~new_P2_U4445 | ~new_P2_U4953;
  assign new_P2_U4955 = ~new_P2_U4954 | ~new_P2_U4943;
  assign new_P2_U4956 = ~P2_STATE2_REG_2_ | ~new_P2_U3392;
  assign new_P2_U4957 = ~new_P2_U4956 | ~new_P2_U4955;
  assign new_P2_U4958 = ~new_P2_U4942 | ~new_P2_U2425;
  assign new_P2_U4959 = ~new_P2_U2485 | ~new_P2_U2422;
  assign new_P2_U4960 = ~new_P2_U4941 | ~new_P2_U2421;
  assign new_P2_U4961 = ~new_P2_U2406 | ~new_P2_U4957;
  assign new_P2_U4962 = ~P2_INSTQUEUE_REG_10__7_ | ~new_P2_U4952;
  assign new_P2_U4963 = ~new_P2_U4942 | ~new_P2_U2426;
  assign new_P2_U4964 = ~new_P2_U2485 | ~new_P2_U2420;
  assign new_P2_U4965 = ~new_P2_U4941 | ~new_P2_U2419;
  assign new_P2_U4966 = ~new_P2_U2405 | ~new_P2_U4957;
  assign new_P2_U4967 = ~P2_INSTQUEUE_REG_10__6_ | ~new_P2_U4952;
  assign new_P2_U4968 = ~new_P2_U4942 | ~new_P2_U2429;
  assign new_P2_U4969 = ~new_P2_U2485 | ~new_P2_U2418;
  assign new_P2_U4970 = ~new_P2_U4941 | ~new_P2_U2417;
  assign new_P2_U4971 = ~new_P2_U2404 | ~new_P2_U4957;
  assign new_P2_U4972 = ~P2_INSTQUEUE_REG_10__5_ | ~new_P2_U4952;
  assign new_P2_U4973 = ~new_P2_U4942 | ~new_P2_U2424;
  assign new_P2_U4974 = ~new_P2_U2485 | ~new_P2_U2416;
  assign new_P2_U4975 = ~new_P2_U4941 | ~new_P2_U2415;
  assign new_P2_U4976 = ~new_P2_U2403 | ~new_P2_U4957;
  assign new_P2_U4977 = ~P2_INSTQUEUE_REG_10__4_ | ~new_P2_U4952;
  assign new_P2_U4978 = ~new_P2_U4942 | ~new_P2_U2423;
  assign new_P2_U4979 = ~new_P2_U2485 | ~new_P2_U2414;
  assign new_P2_U4980 = ~new_P2_U4941 | ~new_P2_U2413;
  assign new_P2_U4981 = ~new_P2_U2402 | ~new_P2_U4957;
  assign new_P2_U4982 = ~P2_INSTQUEUE_REG_10__3_ | ~new_P2_U4952;
  assign new_P2_U4983 = ~new_P2_U4942 | ~new_P2_U2432;
  assign new_P2_U4984 = ~new_P2_U2485 | ~new_P2_U2412;
  assign new_P2_U4985 = ~new_P2_U4941 | ~new_P2_U2411;
  assign new_P2_U4986 = ~new_P2_U2401 | ~new_P2_U4957;
  assign new_P2_U4987 = ~P2_INSTQUEUE_REG_10__2_ | ~new_P2_U4952;
  assign new_P2_U4988 = ~new_P2_U4942 | ~new_P2_U2428;
  assign new_P2_U4989 = ~new_P2_U2485 | ~new_P2_U2410;
  assign new_P2_U4990 = ~new_P2_U4941 | ~new_P2_U2409;
  assign new_P2_U4991 = ~new_P2_U2400 | ~new_P2_U4957;
  assign new_P2_U4992 = ~P2_INSTQUEUE_REG_10__1_ | ~new_P2_U4952;
  assign new_P2_U4993 = ~new_P2_U4942 | ~new_P2_U2431;
  assign new_P2_U4994 = ~new_P2_U2485 | ~new_P2_U2408;
  assign new_P2_U4995 = ~new_P2_U4941 | ~new_P2_U2407;
  assign new_P2_U4996 = ~new_P2_U2399 | ~new_P2_U4957;
  assign new_P2_U4997 = ~P2_INSTQUEUE_REG_10__0_ | ~new_P2_U4952;
  assign new_P2_U4998 = ~new_P2_U3402;
  assign new_P2_U4999 = ~new_P2_U3401;
  assign new_P2_U5000 = ~new_P2_U2442 | ~new_P2_U2445;
  assign new_P2_U5001 = ~new_P2_U3403;
  assign new_P2_U5002 = ~new_P2_U3564;
  assign new_P2_U5003 = ~new_P2_U3404;
  assign new_P2_U5004 = ~new_P2_U4638 | ~new_P2_U4634;
  assign new_P2_U5005 = ~new_P2_U2488 | ~new_P2_U2362;
  assign new_P2_U5006 = ~new_P2_U4445 | ~new_P2_U5005;
  assign new_P2_U5007 = ~new_P2_U5001 | ~new_P2_U5006;
  assign new_P2_U5008 = ~new_P2_U5003 | ~P2_STATE2_REG_2_;
  assign new_P2_U5009 = ~P2_STATE2_REG_3_ | ~new_P2_U3401;
  assign new_P2_U5010 = ~new_P2_U5007 | ~new_P2_U3776;
  assign new_P2_U5011 = ~new_P2_U2488 | ~new_P2_U2398;
  assign new_P2_U5012 = ~new_P2_U4445 | ~new_P2_U5011;
  assign new_P2_U5013 = ~new_P2_U5012 | ~new_P2_U3403;
  assign new_P2_U5014 = ~P2_STATE2_REG_2_ | ~new_P2_U3404;
  assign new_P2_U5015 = ~new_P2_U5014 | ~new_P2_U5013;
  assign new_P2_U5016 = ~new_P2_U4999 | ~new_P2_U2425;
  assign new_P2_U5017 = ~new_P2_U2487 | ~new_P2_U2422;
  assign new_P2_U5018 = ~new_P2_U4998 | ~new_P2_U2421;
  assign new_P2_U5019 = ~new_P2_U2406 | ~new_P2_U5015;
  assign new_P2_U5020 = ~P2_INSTQUEUE_REG_9__7_ | ~new_P2_U5010;
  assign new_P2_U5021 = ~new_P2_U4999 | ~new_P2_U2426;
  assign new_P2_U5022 = ~new_P2_U2487 | ~new_P2_U2420;
  assign new_P2_U5023 = ~new_P2_U4998 | ~new_P2_U2419;
  assign new_P2_U5024 = ~new_P2_U2405 | ~new_P2_U5015;
  assign new_P2_U5025 = ~P2_INSTQUEUE_REG_9__6_ | ~new_P2_U5010;
  assign new_P2_U5026 = ~new_P2_U4999 | ~new_P2_U2429;
  assign new_P2_U5027 = ~new_P2_U2487 | ~new_P2_U2418;
  assign new_P2_U5028 = ~new_P2_U4998 | ~new_P2_U2417;
  assign new_P2_U5029 = ~new_P2_U2404 | ~new_P2_U5015;
  assign new_P2_U5030 = ~P2_INSTQUEUE_REG_9__5_ | ~new_P2_U5010;
  assign new_P2_U5031 = ~new_P2_U4999 | ~new_P2_U2424;
  assign new_P2_U5032 = ~new_P2_U2487 | ~new_P2_U2416;
  assign new_P2_U5033 = ~new_P2_U4998 | ~new_P2_U2415;
  assign new_P2_U5034 = ~new_P2_U2403 | ~new_P2_U5015;
  assign new_P2_U5035 = ~P2_INSTQUEUE_REG_9__4_ | ~new_P2_U5010;
  assign new_P2_U5036 = ~new_P2_U4999 | ~new_P2_U2423;
  assign new_P2_U5037 = ~new_P2_U2487 | ~new_P2_U2414;
  assign new_P2_U5038 = ~new_P2_U4998 | ~new_P2_U2413;
  assign new_P2_U5039 = ~new_P2_U2402 | ~new_P2_U5015;
  assign new_P2_U5040 = ~P2_INSTQUEUE_REG_9__3_ | ~new_P2_U5010;
  assign new_P2_U5041 = ~new_P2_U4999 | ~new_P2_U2432;
  assign new_P2_U5042 = ~new_P2_U2487 | ~new_P2_U2412;
  assign new_P2_U5043 = ~new_P2_U4998 | ~new_P2_U2411;
  assign new_P2_U5044 = ~new_P2_U2401 | ~new_P2_U5015;
  assign new_P2_U5045 = ~P2_INSTQUEUE_REG_9__2_ | ~new_P2_U5010;
  assign new_P2_U5046 = ~new_P2_U4999 | ~new_P2_U2428;
  assign new_P2_U5047 = ~new_P2_U2487 | ~new_P2_U2410;
  assign new_P2_U5048 = ~new_P2_U4998 | ~new_P2_U2409;
  assign new_P2_U5049 = ~new_P2_U2400 | ~new_P2_U5015;
  assign new_P2_U5050 = ~P2_INSTQUEUE_REG_9__1_ | ~new_P2_U5010;
  assign new_P2_U5051 = ~new_P2_U4999 | ~new_P2_U2431;
  assign new_P2_U5052 = ~new_P2_U2487 | ~new_P2_U2408;
  assign new_P2_U5053 = ~new_P2_U4998 | ~new_P2_U2407;
  assign new_P2_U5054 = ~new_P2_U2399 | ~new_P2_U5015;
  assign new_P2_U5055 = ~P2_INSTQUEUE_REG_9__0_ | ~new_P2_U5010;
  assign new_P2_U5056 = ~new_P2_U3414;
  assign new_P2_U5057 = ~new_P2_U3413;
  assign new_P2_U5058 = ~new_P2_U3248;
  assign new_P2_U5059 = ~new_P2_U3563;
  assign new_P2_U5060 = ~new_P2_U3415;
  assign new_P2_U5061 = ~new_P2_U4638 | ~new_P2_U2476;
  assign new_P2_U5062 = ~new_P2_U2490 | ~new_P2_U2362;
  assign new_P2_U5063 = ~new_P2_U4445 | ~new_P2_U5062;
  assign new_P2_U5064 = ~new_P2_U5063 | ~new_P2_U3248;
  assign new_P2_U5065 = ~new_P2_U5060 | ~P2_STATE2_REG_2_;
  assign new_P2_U5066 = ~P2_STATE2_REG_3_ | ~new_P2_U3413;
  assign new_P2_U5067 = ~new_P2_U5064 | ~new_P2_U3785;
  assign new_P2_U5068 = ~new_P2_U2490 | ~new_P2_U2398;
  assign new_P2_U5069 = ~new_P2_U4445 | ~new_P2_U5068;
  assign new_P2_U5070 = ~new_P2_U5069 | ~new_P2_U5058;
  assign new_P2_U5071 = ~P2_STATE2_REG_2_ | ~new_P2_U3415;
  assign new_P2_U5072 = ~new_P2_U5071 | ~new_P2_U5070;
  assign new_P2_U5073 = ~new_P2_U5057 | ~new_P2_U2425;
  assign new_P2_U5074 = ~new_P2_U2489 | ~new_P2_U2422;
  assign new_P2_U5075 = ~new_P2_U5056 | ~new_P2_U2421;
  assign new_P2_U5076 = ~new_P2_U2406 | ~new_P2_U5072;
  assign new_P2_U5077 = ~P2_INSTQUEUE_REG_8__7_ | ~new_P2_U5067;
  assign new_P2_U5078 = ~new_P2_U5057 | ~new_P2_U2426;
  assign new_P2_U5079 = ~new_P2_U2489 | ~new_P2_U2420;
  assign new_P2_U5080 = ~new_P2_U5056 | ~new_P2_U2419;
  assign new_P2_U5081 = ~new_P2_U2405 | ~new_P2_U5072;
  assign new_P2_U5082 = ~P2_INSTQUEUE_REG_8__6_ | ~new_P2_U5067;
  assign new_P2_U5083 = ~new_P2_U5057 | ~new_P2_U2429;
  assign new_P2_U5084 = ~new_P2_U2489 | ~new_P2_U2418;
  assign new_P2_U5085 = ~new_P2_U5056 | ~new_P2_U2417;
  assign new_P2_U5086 = ~new_P2_U2404 | ~new_P2_U5072;
  assign new_P2_U5087 = ~P2_INSTQUEUE_REG_8__5_ | ~new_P2_U5067;
  assign new_P2_U5088 = ~new_P2_U5057 | ~new_P2_U2424;
  assign new_P2_U5089 = ~new_P2_U2489 | ~new_P2_U2416;
  assign new_P2_U5090 = ~new_P2_U5056 | ~new_P2_U2415;
  assign new_P2_U5091 = ~new_P2_U2403 | ~new_P2_U5072;
  assign new_P2_U5092 = ~P2_INSTQUEUE_REG_8__4_ | ~new_P2_U5067;
  assign new_P2_U5093 = ~new_P2_U5057 | ~new_P2_U2423;
  assign new_P2_U5094 = ~new_P2_U2489 | ~new_P2_U2414;
  assign new_P2_U5095 = ~new_P2_U5056 | ~new_P2_U2413;
  assign new_P2_U5096 = ~new_P2_U2402 | ~new_P2_U5072;
  assign new_P2_U5097 = ~P2_INSTQUEUE_REG_8__3_ | ~new_P2_U5067;
  assign new_P2_U5098 = ~new_P2_U5057 | ~new_P2_U2432;
  assign new_P2_U5099 = ~new_P2_U2489 | ~new_P2_U2412;
  assign new_P2_U5100 = ~new_P2_U5056 | ~new_P2_U2411;
  assign new_P2_U5101 = ~new_P2_U2401 | ~new_P2_U5072;
  assign new_P2_U5102 = ~P2_INSTQUEUE_REG_8__2_ | ~new_P2_U5067;
  assign new_P2_U5103 = ~new_P2_U5057 | ~new_P2_U2428;
  assign new_P2_U5104 = ~new_P2_U2489 | ~new_P2_U2410;
  assign new_P2_U5105 = ~new_P2_U5056 | ~new_P2_U2409;
  assign new_P2_U5106 = ~new_P2_U2400 | ~new_P2_U5072;
  assign new_P2_U5107 = ~P2_INSTQUEUE_REG_8__1_ | ~new_P2_U5067;
  assign new_P2_U5108 = ~new_P2_U5057 | ~new_P2_U2431;
  assign new_P2_U5109 = ~new_P2_U2489 | ~new_P2_U2408;
  assign new_P2_U5110 = ~new_P2_U5056 | ~new_P2_U2407;
  assign new_P2_U5111 = ~new_P2_U2399 | ~new_P2_U5072;
  assign new_P2_U5112 = ~P2_INSTQUEUE_REG_8__0_ | ~new_P2_U5067;
  assign new_P2_U5113 = ~new_P2_U3427;
  assign new_P2_U5114 = ~new_P2_U2441 | ~new_P2_U2444;
  assign new_P2_U5115 = ~new_P2_U3429;
  assign new_P2_U5116 = ~new_P2_U3562;
  assign new_P2_U5117 = ~new_P2_U3430;
  assign new_P2_U5118 = ~new_P2_U2493 | ~new_P2_U2362;
  assign new_P2_U5119 = ~new_P2_U4445 | ~new_P2_U5118;
  assign new_P2_U5120 = ~new_P2_U5115 | ~new_P2_U5119;
  assign new_P2_U5121 = ~new_P2_U5117 | ~P2_STATE2_REG_2_;
  assign new_P2_U5122 = ~P2_STATE2_REG_3_ | ~new_P2_U3424;
  assign new_P2_U5123 = ~new_P2_U5120 | ~new_P2_U3794;
  assign new_P2_U5124 = ~new_P2_U2493 | ~new_P2_U2398;
  assign new_P2_U5125 = ~new_P2_U4445 | ~new_P2_U5124;
  assign new_P2_U5126 = ~new_P2_U5125 | ~new_P2_U3429;
  assign new_P2_U5127 = ~P2_STATE2_REG_2_ | ~new_P2_U3430;
  assign new_P2_U5128 = ~new_P2_U5127 | ~new_P2_U5126;
  assign new_P2_U5129 = ~new_P2_U4644 | ~new_P2_U2425;
  assign new_P2_U5130 = ~new_P2_U4451 | ~new_P2_U2422;
  assign new_P2_U5131 = ~new_P2_U5113 | ~new_P2_U2421;
  assign new_P2_U5132 = ~new_P2_U2406 | ~new_P2_U5128;
  assign new_P2_U5133 = ~P2_INSTQUEUE_REG_7__7_ | ~new_P2_U5123;
  assign new_P2_U5134 = ~new_P2_U4644 | ~new_P2_U2426;
  assign new_P2_U5135 = ~new_P2_U4451 | ~new_P2_U2420;
  assign new_P2_U5136 = ~new_P2_U5113 | ~new_P2_U2419;
  assign new_P2_U5137 = ~new_P2_U2405 | ~new_P2_U5128;
  assign new_P2_U5138 = ~P2_INSTQUEUE_REG_7__6_ | ~new_P2_U5123;
  assign new_P2_U5139 = ~new_P2_U4644 | ~new_P2_U2429;
  assign new_P2_U5140 = ~new_P2_U4451 | ~new_P2_U2418;
  assign new_P2_U5141 = ~new_P2_U5113 | ~new_P2_U2417;
  assign new_P2_U5142 = ~new_P2_U2404 | ~new_P2_U5128;
  assign new_P2_U5143 = ~P2_INSTQUEUE_REG_7__5_ | ~new_P2_U5123;
  assign new_P2_U5144 = ~new_P2_U4644 | ~new_P2_U2424;
  assign new_P2_U5145 = ~new_P2_U4451 | ~new_P2_U2416;
  assign new_P2_U5146 = ~new_P2_U5113 | ~new_P2_U2415;
  assign new_P2_U5147 = ~new_P2_U2403 | ~new_P2_U5128;
  assign new_P2_U5148 = ~P2_INSTQUEUE_REG_7__4_ | ~new_P2_U5123;
  assign new_P2_U5149 = ~new_P2_U4644 | ~new_P2_U2423;
  assign new_P2_U5150 = ~new_P2_U4451 | ~new_P2_U2414;
  assign new_P2_U5151 = ~new_P2_U5113 | ~new_P2_U2413;
  assign new_P2_U5152 = ~new_P2_U2402 | ~new_P2_U5128;
  assign new_P2_U5153 = ~P2_INSTQUEUE_REG_7__3_ | ~new_P2_U5123;
  assign new_P2_U5154 = ~new_P2_U4644 | ~new_P2_U2432;
  assign new_P2_U5155 = ~new_P2_U4451 | ~new_P2_U2412;
  assign new_P2_U5156 = ~new_P2_U5113 | ~new_P2_U2411;
  assign new_P2_U5157 = ~new_P2_U2401 | ~new_P2_U5128;
  assign new_P2_U5158 = ~P2_INSTQUEUE_REG_7__2_ | ~new_P2_U5123;
  assign new_P2_U5159 = ~new_P2_U4644 | ~new_P2_U2428;
  assign new_P2_U5160 = ~new_P2_U4451 | ~new_P2_U2410;
  assign new_P2_U5161 = ~new_P2_U5113 | ~new_P2_U2409;
  assign new_P2_U5162 = ~new_P2_U2400 | ~new_P2_U5128;
  assign new_P2_U5163 = ~P2_INSTQUEUE_REG_7__1_ | ~new_P2_U5123;
  assign new_P2_U5164 = ~new_P2_U4644 | ~new_P2_U2431;
  assign new_P2_U5165 = ~new_P2_U4451 | ~new_P2_U2408;
  assign new_P2_U5166 = ~new_P2_U5113 | ~new_P2_U2407;
  assign new_P2_U5167 = ~new_P2_U2399 | ~new_P2_U5128;
  assign new_P2_U5168 = ~P2_INSTQUEUE_REG_7__0_ | ~new_P2_U5123;
  assign new_P2_U5169 = ~new_P2_U3440;
  assign new_P2_U5170 = ~new_P2_U3439;
  assign new_P2_U5171 = ~new_P2_U3249;
  assign new_P2_U5172 = ~new_P2_U3561;
  assign new_P2_U5173 = ~new_P2_U3441;
  assign new_P2_U5174 = ~new_P2_U4633 | ~new_P2_U2460;
  assign new_P2_U5175 = ~new_P2_U2495 | ~new_P2_U2362;
  assign new_P2_U5176 = ~new_P2_U4445 | ~new_P2_U5175;
  assign new_P2_U5177 = ~new_P2_U5176 | ~new_P2_U3249;
  assign new_P2_U5178 = ~new_P2_U5173 | ~P2_STATE2_REG_2_;
  assign new_P2_U5179 = ~P2_STATE2_REG_3_ | ~new_P2_U3439;
  assign new_P2_U5180 = ~new_P2_U5177 | ~new_P2_U3803;
  assign new_P2_U5181 = ~new_P2_U2495 | ~new_P2_U2398;
  assign new_P2_U5182 = ~new_P2_U4445 | ~new_P2_U5181;
  assign new_P2_U5183 = ~new_P2_U5182 | ~new_P2_U5171;
  assign new_P2_U5184 = ~P2_STATE2_REG_2_ | ~new_P2_U3441;
  assign new_P2_U5185 = ~new_P2_U5184 | ~new_P2_U5183;
  assign new_P2_U5186 = ~new_P2_U5170 | ~new_P2_U2425;
  assign new_P2_U5187 = ~new_P2_U2494 | ~new_P2_U2422;
  assign new_P2_U5188 = ~new_P2_U5169 | ~new_P2_U2421;
  assign new_P2_U5189 = ~new_P2_U2406 | ~new_P2_U5185;
  assign new_P2_U5190 = ~P2_INSTQUEUE_REG_6__7_ | ~new_P2_U5180;
  assign new_P2_U5191 = ~new_P2_U5170 | ~new_P2_U2426;
  assign new_P2_U5192 = ~new_P2_U2494 | ~new_P2_U2420;
  assign new_P2_U5193 = ~new_P2_U5169 | ~new_P2_U2419;
  assign new_P2_U5194 = ~new_P2_U2405 | ~new_P2_U5185;
  assign new_P2_U5195 = ~P2_INSTQUEUE_REG_6__6_ | ~new_P2_U5180;
  assign new_P2_U5196 = ~new_P2_U5170 | ~new_P2_U2429;
  assign new_P2_U5197 = ~new_P2_U2494 | ~new_P2_U2418;
  assign new_P2_U5198 = ~new_P2_U5169 | ~new_P2_U2417;
  assign new_P2_U5199 = ~new_P2_U2404 | ~new_P2_U5185;
  assign new_P2_U5200 = ~P2_INSTQUEUE_REG_6__5_ | ~new_P2_U5180;
  assign new_P2_U5201 = ~new_P2_U5170 | ~new_P2_U2424;
  assign new_P2_U5202 = ~new_P2_U2494 | ~new_P2_U2416;
  assign new_P2_U5203 = ~new_P2_U5169 | ~new_P2_U2415;
  assign new_P2_U5204 = ~new_P2_U2403 | ~new_P2_U5185;
  assign new_P2_U5205 = ~P2_INSTQUEUE_REG_6__4_ | ~new_P2_U5180;
  assign new_P2_U5206 = ~new_P2_U5170 | ~new_P2_U2423;
  assign new_P2_U5207 = ~new_P2_U2494 | ~new_P2_U2414;
  assign new_P2_U5208 = ~new_P2_U5169 | ~new_P2_U2413;
  assign new_P2_U5209 = ~new_P2_U2402 | ~new_P2_U5185;
  assign new_P2_U5210 = ~P2_INSTQUEUE_REG_6__3_ | ~new_P2_U5180;
  assign new_P2_U5211 = ~new_P2_U5170 | ~new_P2_U2432;
  assign new_P2_U5212 = ~new_P2_U2494 | ~new_P2_U2412;
  assign new_P2_U5213 = ~new_P2_U5169 | ~new_P2_U2411;
  assign new_P2_U5214 = ~new_P2_U2401 | ~new_P2_U5185;
  assign new_P2_U5215 = ~P2_INSTQUEUE_REG_6__2_ | ~new_P2_U5180;
  assign new_P2_U5216 = ~new_P2_U5170 | ~new_P2_U2428;
  assign new_P2_U5217 = ~new_P2_U2494 | ~new_P2_U2410;
  assign new_P2_U5218 = ~new_P2_U5169 | ~new_P2_U2409;
  assign new_P2_U5219 = ~new_P2_U2400 | ~new_P2_U5185;
  assign new_P2_U5220 = ~P2_INSTQUEUE_REG_6__1_ | ~new_P2_U5180;
  assign new_P2_U5221 = ~new_P2_U5170 | ~new_P2_U2431;
  assign new_P2_U5222 = ~new_P2_U2494 | ~new_P2_U2408;
  assign new_P2_U5223 = ~new_P2_U5169 | ~new_P2_U2407;
  assign new_P2_U5224 = ~new_P2_U2399 | ~new_P2_U5185;
  assign new_P2_U5225 = ~P2_INSTQUEUE_REG_6__0_ | ~new_P2_U5180;
  assign new_P2_U5226 = ~new_P2_U3451;
  assign new_P2_U5227 = ~new_P2_U3450;
  assign new_P2_U5228 = ~new_P2_U2441 | ~new_P2_U2445;
  assign new_P2_U5229 = ~new_P2_U3452;
  assign new_P2_U5230 = ~new_P2_U3560;
  assign new_P2_U5231 = ~new_P2_U3453;
  assign new_P2_U5232 = ~new_P2_U4634 | ~new_P2_U2460;
  assign new_P2_U5233 = ~new_P2_U2497 | ~new_P2_U2362;
  assign new_P2_U5234 = ~new_P2_U4445 | ~new_P2_U5233;
  assign new_P2_U5235 = ~new_P2_U5229 | ~new_P2_U5234;
  assign new_P2_U5236 = ~new_P2_U5231 | ~P2_STATE2_REG_2_;
  assign new_P2_U5237 = ~P2_STATE2_REG_3_ | ~new_P2_U3450;
  assign new_P2_U5238 = ~new_P2_U5235 | ~new_P2_U3812;
  assign new_P2_U5239 = ~new_P2_U2497 | ~new_P2_U2398;
  assign new_P2_U5240 = ~new_P2_U4445 | ~new_P2_U5239;
  assign new_P2_U5241 = ~new_P2_U5240 | ~new_P2_U3452;
  assign new_P2_U5242 = ~P2_STATE2_REG_2_ | ~new_P2_U3453;
  assign new_P2_U5243 = ~new_P2_U5242 | ~new_P2_U5241;
  assign new_P2_U5244 = ~new_P2_U5227 | ~new_P2_U2425;
  assign new_P2_U5245 = ~new_P2_U2496 | ~new_P2_U2422;
  assign new_P2_U5246 = ~new_P2_U5226 | ~new_P2_U2421;
  assign new_P2_U5247 = ~new_P2_U2406 | ~new_P2_U5243;
  assign new_P2_U5248 = ~P2_INSTQUEUE_REG_5__7_ | ~new_P2_U5238;
  assign new_P2_U5249 = ~new_P2_U5227 | ~new_P2_U2426;
  assign new_P2_U5250 = ~new_P2_U2496 | ~new_P2_U2420;
  assign new_P2_U5251 = ~new_P2_U5226 | ~new_P2_U2419;
  assign new_P2_U5252 = ~new_P2_U2405 | ~new_P2_U5243;
  assign new_P2_U5253 = ~P2_INSTQUEUE_REG_5__6_ | ~new_P2_U5238;
  assign new_P2_U5254 = ~new_P2_U5227 | ~new_P2_U2429;
  assign new_P2_U5255 = ~new_P2_U2496 | ~new_P2_U2418;
  assign new_P2_U5256 = ~new_P2_U5226 | ~new_P2_U2417;
  assign new_P2_U5257 = ~new_P2_U2404 | ~new_P2_U5243;
  assign new_P2_U5258 = ~P2_INSTQUEUE_REG_5__5_ | ~new_P2_U5238;
  assign new_P2_U5259 = ~new_P2_U5227 | ~new_P2_U2424;
  assign new_P2_U5260 = ~new_P2_U2496 | ~new_P2_U2416;
  assign new_P2_U5261 = ~new_P2_U5226 | ~new_P2_U2415;
  assign new_P2_U5262 = ~new_P2_U2403 | ~new_P2_U5243;
  assign new_P2_U5263 = ~P2_INSTQUEUE_REG_5__4_ | ~new_P2_U5238;
  assign new_P2_U5264 = ~new_P2_U5227 | ~new_P2_U2423;
  assign new_P2_U5265 = ~new_P2_U2496 | ~new_P2_U2414;
  assign new_P2_U5266 = ~new_P2_U5226 | ~new_P2_U2413;
  assign new_P2_U5267 = ~new_P2_U2402 | ~new_P2_U5243;
  assign new_P2_U5268 = ~P2_INSTQUEUE_REG_5__3_ | ~new_P2_U5238;
  assign new_P2_U5269 = ~new_P2_U5227 | ~new_P2_U2432;
  assign new_P2_U5270 = ~new_P2_U2496 | ~new_P2_U2412;
  assign new_P2_U5271 = ~new_P2_U5226 | ~new_P2_U2411;
  assign new_P2_U5272 = ~new_P2_U2401 | ~new_P2_U5243;
  assign new_P2_U5273 = ~P2_INSTQUEUE_REG_5__2_ | ~new_P2_U5238;
  assign new_P2_U5274 = ~new_P2_U5227 | ~new_P2_U2428;
  assign new_P2_U5275 = ~new_P2_U2496 | ~new_P2_U2410;
  assign new_P2_U5276 = ~new_P2_U5226 | ~new_P2_U2409;
  assign new_P2_U5277 = ~new_P2_U2400 | ~new_P2_U5243;
  assign new_P2_U5278 = ~P2_INSTQUEUE_REG_5__1_ | ~new_P2_U5238;
  assign new_P2_U5279 = ~new_P2_U5227 | ~new_P2_U2431;
  assign new_P2_U5280 = ~new_P2_U2496 | ~new_P2_U2408;
  assign new_P2_U5281 = ~new_P2_U5226 | ~new_P2_U2407;
  assign new_P2_U5282 = ~new_P2_U2399 | ~new_P2_U5243;
  assign new_P2_U5283 = ~P2_INSTQUEUE_REG_5__0_ | ~new_P2_U5238;
  assign new_P2_U5284 = ~new_P2_U3463;
  assign new_P2_U5285 = ~new_P2_U3462;
  assign new_P2_U5286 = ~new_P2_U3250;
  assign new_P2_U5287 = ~new_P2_U3559;
  assign new_P2_U5288 = ~new_P2_U3464;
  assign new_P2_U5289 = ~new_P2_U2476 | ~new_P2_U2460;
  assign new_P2_U5290 = ~new_P2_U2499 | ~new_P2_U2362;
  assign new_P2_U5291 = ~new_P2_U4445 | ~new_P2_U5290;
  assign new_P2_U5292 = ~new_P2_U5291 | ~new_P2_U3250;
  assign new_P2_U5293 = ~new_P2_U5288 | ~P2_STATE2_REG_2_;
  assign new_P2_U5294 = ~P2_STATE2_REG_3_ | ~new_P2_U3462;
  assign new_P2_U5295 = ~new_P2_U5292 | ~new_P2_U3821;
  assign new_P2_U5296 = ~new_P2_U2499 | ~new_P2_U2398;
  assign new_P2_U5297 = ~new_P2_U4445 | ~new_P2_U5296;
  assign new_P2_U5298 = ~new_P2_U5297 | ~new_P2_U5286;
  assign new_P2_U5299 = ~P2_STATE2_REG_2_ | ~new_P2_U3464;
  assign new_P2_U5300 = ~new_P2_U5299 | ~new_P2_U5298;
  assign new_P2_U5301 = ~new_P2_U5285 | ~new_P2_U2425;
  assign new_P2_U5302 = ~new_P2_U2498 | ~new_P2_U2422;
  assign new_P2_U5303 = ~new_P2_U5284 | ~new_P2_U2421;
  assign new_P2_U5304 = ~new_P2_U2406 | ~new_P2_U5300;
  assign new_P2_U5305 = ~P2_INSTQUEUE_REG_4__7_ | ~new_P2_U5295;
  assign new_P2_U5306 = ~new_P2_U5285 | ~new_P2_U2426;
  assign new_P2_U5307 = ~new_P2_U2498 | ~new_P2_U2420;
  assign new_P2_U5308 = ~new_P2_U5284 | ~new_P2_U2419;
  assign new_P2_U5309 = ~new_P2_U2405 | ~new_P2_U5300;
  assign new_P2_U5310 = ~P2_INSTQUEUE_REG_4__6_ | ~new_P2_U5295;
  assign new_P2_U5311 = ~new_P2_U5285 | ~new_P2_U2429;
  assign new_P2_U5312 = ~new_P2_U2498 | ~new_P2_U2418;
  assign new_P2_U5313 = ~new_P2_U5284 | ~new_P2_U2417;
  assign new_P2_U5314 = ~new_P2_U2404 | ~new_P2_U5300;
  assign new_P2_U5315 = ~P2_INSTQUEUE_REG_4__5_ | ~new_P2_U5295;
  assign new_P2_U5316 = ~new_P2_U5285 | ~new_P2_U2424;
  assign new_P2_U5317 = ~new_P2_U2498 | ~new_P2_U2416;
  assign new_P2_U5318 = ~new_P2_U5284 | ~new_P2_U2415;
  assign new_P2_U5319 = ~new_P2_U2403 | ~new_P2_U5300;
  assign new_P2_U5320 = ~P2_INSTQUEUE_REG_4__4_ | ~new_P2_U5295;
  assign new_P2_U5321 = ~new_P2_U5285 | ~new_P2_U2423;
  assign new_P2_U5322 = ~new_P2_U2498 | ~new_P2_U2414;
  assign new_P2_U5323 = ~new_P2_U5284 | ~new_P2_U2413;
  assign new_P2_U5324 = ~new_P2_U2402 | ~new_P2_U5300;
  assign new_P2_U5325 = ~P2_INSTQUEUE_REG_4__3_ | ~new_P2_U5295;
  assign new_P2_U5326 = ~new_P2_U5285 | ~new_P2_U2432;
  assign new_P2_U5327 = ~new_P2_U2498 | ~new_P2_U2412;
  assign new_P2_U5328 = ~new_P2_U5284 | ~new_P2_U2411;
  assign new_P2_U5329 = ~new_P2_U2401 | ~new_P2_U5300;
  assign new_P2_U5330 = ~P2_INSTQUEUE_REG_4__2_ | ~new_P2_U5295;
  assign new_P2_U5331 = ~new_P2_U5285 | ~new_P2_U2428;
  assign new_P2_U5332 = ~new_P2_U2498 | ~new_P2_U2410;
  assign new_P2_U5333 = ~new_P2_U5284 | ~new_P2_U2409;
  assign new_P2_U5334 = ~new_P2_U2400 | ~new_P2_U5300;
  assign new_P2_U5335 = ~P2_INSTQUEUE_REG_4__1_ | ~new_P2_U5295;
  assign new_P2_U5336 = ~new_P2_U5285 | ~new_P2_U2431;
  assign new_P2_U5337 = ~new_P2_U2498 | ~new_P2_U2408;
  assign new_P2_U5338 = ~new_P2_U5284 | ~new_P2_U2407;
  assign new_P2_U5339 = ~new_P2_U2399 | ~new_P2_U5300;
  assign new_P2_U5340 = ~P2_INSTQUEUE_REG_4__0_ | ~new_P2_U5295;
  assign new_P2_U5341 = ~new_P2_U3474;
  assign new_P2_U5342 = ~new_P2_U3473;
  assign new_P2_U5343 = ~new_P2_U2443 | ~new_P2_U2444;
  assign new_P2_U5344 = ~new_P2_U3475;
  assign new_P2_U5345 = ~new_P2_U3558;
  assign new_P2_U5346 = ~new_P2_U3476;
  assign new_P2_U5347 = ~new_P2_U2501 | ~new_P2_U4637;
  assign new_P2_U5348 = ~new_P2_U2505 | ~new_P2_U2362;
  assign new_P2_U5349 = ~new_P2_U4445 | ~new_P2_U5348;
  assign new_P2_U5350 = ~new_P2_U5344 | ~new_P2_U5349;
  assign new_P2_U5351 = ~new_P2_U5346 | ~P2_STATE2_REG_2_;
  assign new_P2_U5352 = ~P2_STATE2_REG_3_ | ~new_P2_U3473;
  assign new_P2_U5353 = ~new_P2_U5350 | ~new_P2_U3830;
  assign new_P2_U5354 = ~new_P2_U2505 | ~new_P2_U2398;
  assign new_P2_U5355 = ~new_P2_U4445 | ~new_P2_U5354;
  assign new_P2_U5356 = ~new_P2_U5355 | ~new_P2_U3475;
  assign new_P2_U5357 = ~P2_STATE2_REG_2_ | ~new_P2_U3476;
  assign new_P2_U5358 = ~new_P2_U5357 | ~new_P2_U5356;
  assign new_P2_U5359 = ~new_P2_U5342 | ~new_P2_U2425;
  assign new_P2_U5360 = ~new_P2_U2502 | ~new_P2_U2422;
  assign new_P2_U5361 = ~new_P2_U5341 | ~new_P2_U2421;
  assign new_P2_U5362 = ~new_P2_U2406 | ~new_P2_U5358;
  assign new_P2_U5363 = ~P2_INSTQUEUE_REG_3__7_ | ~new_P2_U5353;
  assign new_P2_U5364 = ~new_P2_U5342 | ~new_P2_U2426;
  assign new_P2_U5365 = ~new_P2_U2502 | ~new_P2_U2420;
  assign new_P2_U5366 = ~new_P2_U5341 | ~new_P2_U2419;
  assign new_P2_U5367 = ~new_P2_U2405 | ~new_P2_U5358;
  assign new_P2_U5368 = ~P2_INSTQUEUE_REG_3__6_ | ~new_P2_U5353;
  assign new_P2_U5369 = ~new_P2_U5342 | ~new_P2_U2429;
  assign new_P2_U5370 = ~new_P2_U2502 | ~new_P2_U2418;
  assign new_P2_U5371 = ~new_P2_U5341 | ~new_P2_U2417;
  assign new_P2_U5372 = ~new_P2_U2404 | ~new_P2_U5358;
  assign new_P2_U5373 = ~P2_INSTQUEUE_REG_3__5_ | ~new_P2_U5353;
  assign new_P2_U5374 = ~new_P2_U5342 | ~new_P2_U2424;
  assign new_P2_U5375 = ~new_P2_U2502 | ~new_P2_U2416;
  assign new_P2_U5376 = ~new_P2_U5341 | ~new_P2_U2415;
  assign new_P2_U5377 = ~new_P2_U2403 | ~new_P2_U5358;
  assign new_P2_U5378 = ~P2_INSTQUEUE_REG_3__4_ | ~new_P2_U5353;
  assign new_P2_U5379 = ~new_P2_U5342 | ~new_P2_U2423;
  assign new_P2_U5380 = ~new_P2_U2502 | ~new_P2_U2414;
  assign new_P2_U5381 = ~new_P2_U5341 | ~new_P2_U2413;
  assign new_P2_U5382 = ~new_P2_U2402 | ~new_P2_U5358;
  assign new_P2_U5383 = ~P2_INSTQUEUE_REG_3__3_ | ~new_P2_U5353;
  assign new_P2_U5384 = ~new_P2_U5342 | ~new_P2_U2432;
  assign new_P2_U5385 = ~new_P2_U2502 | ~new_P2_U2412;
  assign new_P2_U5386 = ~new_P2_U5341 | ~new_P2_U2411;
  assign new_P2_U5387 = ~new_P2_U2401 | ~new_P2_U5358;
  assign new_P2_U5388 = ~P2_INSTQUEUE_REG_3__2_ | ~new_P2_U5353;
  assign new_P2_U5389 = ~new_P2_U5342 | ~new_P2_U2428;
  assign new_P2_U5390 = ~new_P2_U2502 | ~new_P2_U2410;
  assign new_P2_U5391 = ~new_P2_U5341 | ~new_P2_U2409;
  assign new_P2_U5392 = ~new_P2_U2400 | ~new_P2_U5358;
  assign new_P2_U5393 = ~P2_INSTQUEUE_REG_3__1_ | ~new_P2_U5353;
  assign new_P2_U5394 = ~new_P2_U5342 | ~new_P2_U2431;
  assign new_P2_U5395 = ~new_P2_U2502 | ~new_P2_U2408;
  assign new_P2_U5396 = ~new_P2_U5341 | ~new_P2_U2407;
  assign new_P2_U5397 = ~new_P2_U2399 | ~new_P2_U5358;
  assign new_P2_U5398 = ~P2_INSTQUEUE_REG_3__0_ | ~new_P2_U5353;
  assign new_P2_U5399 = ~new_P2_U3486;
  assign new_P2_U5400 = ~new_P2_U3485;
  assign new_P2_U5401 = ~new_P2_U3251;
  assign new_P2_U5402 = ~new_P2_U3557;
  assign new_P2_U5403 = ~new_P2_U3487;
  assign new_P2_U5404 = ~new_P2_U2501 | ~new_P2_U4633;
  assign new_P2_U5405 = ~new_P2_U2507 | ~new_P2_U2362;
  assign new_P2_U5406 = ~new_P2_U4445 | ~new_P2_U5405;
  assign new_P2_U5407 = ~new_P2_U5406 | ~new_P2_U3251;
  assign new_P2_U5408 = ~new_P2_U5403 | ~P2_STATE2_REG_2_;
  assign new_P2_U5409 = ~P2_STATE2_REG_3_ | ~new_P2_U3485;
  assign new_P2_U5410 = ~new_P2_U5407 | ~new_P2_U3839;
  assign new_P2_U5411 = ~new_P2_U2507 | ~new_P2_U2398;
  assign new_P2_U5412 = ~new_P2_U4445 | ~new_P2_U5411;
  assign new_P2_U5413 = ~new_P2_U5412 | ~new_P2_U5401;
  assign new_P2_U5414 = ~P2_STATE2_REG_2_ | ~new_P2_U3487;
  assign new_P2_U5415 = ~new_P2_U5414 | ~new_P2_U5413;
  assign new_P2_U5416 = ~new_P2_U5400 | ~new_P2_U2425;
  assign new_P2_U5417 = ~new_P2_U2506 | ~new_P2_U2422;
  assign new_P2_U5418 = ~new_P2_U5399 | ~new_P2_U2421;
  assign new_P2_U5419 = ~new_P2_U2406 | ~new_P2_U5415;
  assign new_P2_U5420 = ~P2_INSTQUEUE_REG_2__7_ | ~new_P2_U5410;
  assign new_P2_U5421 = ~new_P2_U5400 | ~new_P2_U2426;
  assign new_P2_U5422 = ~new_P2_U2506 | ~new_P2_U2420;
  assign new_P2_U5423 = ~new_P2_U5399 | ~new_P2_U2419;
  assign new_P2_U5424 = ~new_P2_U2405 | ~new_P2_U5415;
  assign new_P2_U5425 = ~P2_INSTQUEUE_REG_2__6_ | ~new_P2_U5410;
  assign new_P2_U5426 = ~new_P2_U5400 | ~new_P2_U2429;
  assign new_P2_U5427 = ~new_P2_U2506 | ~new_P2_U2418;
  assign new_P2_U5428 = ~new_P2_U5399 | ~new_P2_U2417;
  assign new_P2_U5429 = ~new_P2_U2404 | ~new_P2_U5415;
  assign new_P2_U5430 = ~P2_INSTQUEUE_REG_2__5_ | ~new_P2_U5410;
  assign new_P2_U5431 = ~new_P2_U5400 | ~new_P2_U2424;
  assign new_P2_U5432 = ~new_P2_U2506 | ~new_P2_U2416;
  assign new_P2_U5433 = ~new_P2_U5399 | ~new_P2_U2415;
  assign new_P2_U5434 = ~new_P2_U2403 | ~new_P2_U5415;
  assign new_P2_U5435 = ~P2_INSTQUEUE_REG_2__4_ | ~new_P2_U5410;
  assign new_P2_U5436 = ~new_P2_U5400 | ~new_P2_U2423;
  assign new_P2_U5437 = ~new_P2_U2506 | ~new_P2_U2414;
  assign new_P2_U5438 = ~new_P2_U5399 | ~new_P2_U2413;
  assign new_P2_U5439 = ~new_P2_U2402 | ~new_P2_U5415;
  assign new_P2_U5440 = ~P2_INSTQUEUE_REG_2__3_ | ~new_P2_U5410;
  assign new_P2_U5441 = ~new_P2_U5400 | ~new_P2_U2432;
  assign new_P2_U5442 = ~new_P2_U2506 | ~new_P2_U2412;
  assign new_P2_U5443 = ~new_P2_U5399 | ~new_P2_U2411;
  assign new_P2_U5444 = ~new_P2_U2401 | ~new_P2_U5415;
  assign new_P2_U5445 = ~P2_INSTQUEUE_REG_2__2_ | ~new_P2_U5410;
  assign new_P2_U5446 = ~new_P2_U5400 | ~new_P2_U2428;
  assign new_P2_U5447 = ~new_P2_U2506 | ~new_P2_U2410;
  assign new_P2_U5448 = ~new_P2_U5399 | ~new_P2_U2409;
  assign new_P2_U5449 = ~new_P2_U2400 | ~new_P2_U5415;
  assign new_P2_U5450 = ~P2_INSTQUEUE_REG_2__1_ | ~new_P2_U5410;
  assign new_P2_U5451 = ~new_P2_U5400 | ~new_P2_U2431;
  assign new_P2_U5452 = ~new_P2_U2506 | ~new_P2_U2408;
  assign new_P2_U5453 = ~new_P2_U5399 | ~new_P2_U2407;
  assign new_P2_U5454 = ~new_P2_U2399 | ~new_P2_U5415;
  assign new_P2_U5455 = ~P2_INSTQUEUE_REG_2__0_ | ~new_P2_U5410;
  assign new_P2_U5456 = ~new_P2_U3497;
  assign new_P2_U5457 = ~new_P2_U3496;
  assign new_P2_U5458 = ~new_P2_U2443 | ~new_P2_U2445;
  assign new_P2_U5459 = ~new_P2_U3498;
  assign new_P2_U5460 = ~new_P2_U3556;
  assign new_P2_U5461 = ~new_P2_U3499;
  assign new_P2_U5462 = ~new_P2_U2501 | ~new_P2_U4634;
  assign new_P2_U5463 = ~new_P2_U2509 | ~new_P2_U2362;
  assign new_P2_U5464 = ~new_P2_U4445 | ~new_P2_U5463;
  assign new_P2_U5465 = ~new_P2_U5459 | ~new_P2_U5464;
  assign new_P2_U5466 = ~new_P2_U5461 | ~P2_STATE2_REG_2_;
  assign new_P2_U5467 = ~P2_STATE2_REG_3_ | ~new_P2_U3496;
  assign new_P2_U5468 = ~new_P2_U5465 | ~new_P2_U3848;
  assign new_P2_U5469 = ~new_P2_U2509 | ~new_P2_U2398;
  assign new_P2_U5470 = ~new_P2_U4445 | ~new_P2_U5469;
  assign new_P2_U5471 = ~new_P2_U5470 | ~new_P2_U3498;
  assign new_P2_U5472 = ~P2_STATE2_REG_2_ | ~new_P2_U3499;
  assign new_P2_U5473 = ~new_P2_U5472 | ~new_P2_U5471;
  assign new_P2_U5474 = ~new_P2_U5457 | ~new_P2_U2425;
  assign new_P2_U5475 = ~new_P2_U2508 | ~new_P2_U2422;
  assign new_P2_U5476 = ~new_P2_U5456 | ~new_P2_U2421;
  assign new_P2_U5477 = ~new_P2_U2406 | ~new_P2_U5473;
  assign new_P2_U5478 = ~P2_INSTQUEUE_REG_1__7_ | ~new_P2_U5468;
  assign new_P2_U5479 = ~new_P2_U5457 | ~new_P2_U2426;
  assign new_P2_U5480 = ~new_P2_U2508 | ~new_P2_U2420;
  assign new_P2_U5481 = ~new_P2_U5456 | ~new_P2_U2419;
  assign new_P2_U5482 = ~new_P2_U2405 | ~new_P2_U5473;
  assign new_P2_U5483 = ~P2_INSTQUEUE_REG_1__6_ | ~new_P2_U5468;
  assign new_P2_U5484 = ~new_P2_U5457 | ~new_P2_U2429;
  assign new_P2_U5485 = ~new_P2_U2508 | ~new_P2_U2418;
  assign new_P2_U5486 = ~new_P2_U5456 | ~new_P2_U2417;
  assign new_P2_U5487 = ~new_P2_U2404 | ~new_P2_U5473;
  assign new_P2_U5488 = ~P2_INSTQUEUE_REG_1__5_ | ~new_P2_U5468;
  assign new_P2_U5489 = ~new_P2_U5457 | ~new_P2_U2424;
  assign new_P2_U5490 = ~new_P2_U2508 | ~new_P2_U2416;
  assign new_P2_U5491 = ~new_P2_U5456 | ~new_P2_U2415;
  assign new_P2_U5492 = ~new_P2_U2403 | ~new_P2_U5473;
  assign new_P2_U5493 = ~P2_INSTQUEUE_REG_1__4_ | ~new_P2_U5468;
  assign new_P2_U5494 = ~new_P2_U5457 | ~new_P2_U2423;
  assign new_P2_U5495 = ~new_P2_U2508 | ~new_P2_U2414;
  assign new_P2_U5496 = ~new_P2_U5456 | ~new_P2_U2413;
  assign new_P2_U5497 = ~new_P2_U2402 | ~new_P2_U5473;
  assign new_P2_U5498 = ~P2_INSTQUEUE_REG_1__3_ | ~new_P2_U5468;
  assign new_P2_U5499 = ~new_P2_U5457 | ~new_P2_U2432;
  assign new_P2_U5500 = ~new_P2_U2508 | ~new_P2_U2412;
  assign new_P2_U5501 = ~new_P2_U5456 | ~new_P2_U2411;
  assign new_P2_U5502 = ~new_P2_U2401 | ~new_P2_U5473;
  assign new_P2_U5503 = ~P2_INSTQUEUE_REG_1__2_ | ~new_P2_U5468;
  assign new_P2_U5504 = ~new_P2_U5457 | ~new_P2_U2428;
  assign new_P2_U5505 = ~new_P2_U2508 | ~new_P2_U2410;
  assign new_P2_U5506 = ~new_P2_U5456 | ~new_P2_U2409;
  assign new_P2_U5507 = ~new_P2_U2400 | ~new_P2_U5473;
  assign new_P2_U5508 = ~P2_INSTQUEUE_REG_1__1_ | ~new_P2_U5468;
  assign new_P2_U5509 = ~new_P2_U5457 | ~new_P2_U2431;
  assign new_P2_U5510 = ~new_P2_U2508 | ~new_P2_U2408;
  assign new_P2_U5511 = ~new_P2_U5456 | ~new_P2_U2407;
  assign new_P2_U5512 = ~new_P2_U2399 | ~new_P2_U5473;
  assign new_P2_U5513 = ~P2_INSTQUEUE_REG_1__0_ | ~new_P2_U5468;
  assign new_P2_U5514 = ~new_P2_U3509;
  assign new_P2_U5515 = ~new_P2_U3508;
  assign new_P2_U5516 = ~new_P2_U3252;
  assign new_P2_U5517 = ~new_P2_U3555;
  assign new_P2_U5518 = ~new_P2_U3510;
  assign new_P2_U5519 = ~new_P2_U2501 | ~new_P2_U2476;
  assign new_P2_U5520 = ~new_P2_U2511 | ~new_P2_U2362;
  assign new_P2_U5521 = ~new_P2_U4445 | ~new_P2_U5520;
  assign new_P2_U5522 = ~new_P2_U5521 | ~new_P2_U3252;
  assign new_P2_U5523 = ~new_P2_U5518 | ~P2_STATE2_REG_2_;
  assign new_P2_U5524 = ~P2_STATE2_REG_3_ | ~new_P2_U3508;
  assign new_P2_U5525 = ~new_P2_U5522 | ~new_P2_U3857;
  assign new_P2_U5526 = ~new_P2_U2511 | ~new_P2_U2398;
  assign new_P2_U5527 = ~new_P2_U4445 | ~new_P2_U5526;
  assign new_P2_U5528 = ~new_P2_U5527 | ~new_P2_U5516;
  assign new_P2_U5529 = ~P2_STATE2_REG_2_ | ~new_P2_U3510;
  assign new_P2_U5530 = ~new_P2_U5529 | ~new_P2_U5528;
  assign new_P2_U5531 = ~new_P2_U5515 | ~new_P2_U2425;
  assign new_P2_U5532 = ~new_P2_U2510 | ~new_P2_U2422;
  assign new_P2_U5533 = ~new_P2_U5514 | ~new_P2_U2421;
  assign new_P2_U5534 = ~new_P2_U2406 | ~new_P2_U5530;
  assign new_P2_U5535 = ~P2_INSTQUEUE_REG_0__7_ | ~new_P2_U5525;
  assign new_P2_U5536 = ~new_P2_U5515 | ~new_P2_U2426;
  assign new_P2_U5537 = ~new_P2_U2510 | ~new_P2_U2420;
  assign new_P2_U5538 = ~new_P2_U5514 | ~new_P2_U2419;
  assign new_P2_U5539 = ~new_P2_U2405 | ~new_P2_U5530;
  assign new_P2_U5540 = ~P2_INSTQUEUE_REG_0__6_ | ~new_P2_U5525;
  assign new_P2_U5541 = ~new_P2_U5515 | ~new_P2_U2429;
  assign new_P2_U5542 = ~new_P2_U2510 | ~new_P2_U2418;
  assign new_P2_U5543 = ~new_P2_U5514 | ~new_P2_U2417;
  assign new_P2_U5544 = ~new_P2_U2404 | ~new_P2_U5530;
  assign new_P2_U5545 = ~P2_INSTQUEUE_REG_0__5_ | ~new_P2_U5525;
  assign new_P2_U5546 = ~new_P2_U5515 | ~new_P2_U2424;
  assign new_P2_U5547 = ~new_P2_U2510 | ~new_P2_U2416;
  assign new_P2_U5548 = ~new_P2_U5514 | ~new_P2_U2415;
  assign new_P2_U5549 = ~new_P2_U2403 | ~new_P2_U5530;
  assign new_P2_U5550 = ~P2_INSTQUEUE_REG_0__4_ | ~new_P2_U5525;
  assign new_P2_U5551 = ~new_P2_U5515 | ~new_P2_U2423;
  assign new_P2_U5552 = ~new_P2_U2510 | ~new_P2_U2414;
  assign new_P2_U5553 = ~new_P2_U5514 | ~new_P2_U2413;
  assign new_P2_U5554 = ~new_P2_U2402 | ~new_P2_U5530;
  assign new_P2_U5555 = ~P2_INSTQUEUE_REG_0__3_ | ~new_P2_U5525;
  assign new_P2_U5556 = ~new_P2_U5515 | ~new_P2_U2432;
  assign new_P2_U5557 = ~new_P2_U2510 | ~new_P2_U2412;
  assign new_P2_U5558 = ~new_P2_U5514 | ~new_P2_U2411;
  assign new_P2_U5559 = ~new_P2_U2401 | ~new_P2_U5530;
  assign new_P2_U5560 = ~P2_INSTQUEUE_REG_0__2_ | ~new_P2_U5525;
  assign new_P2_U5561 = ~new_P2_U5515 | ~new_P2_U2428;
  assign new_P2_U5562 = ~new_P2_U2510 | ~new_P2_U2410;
  assign new_P2_U5563 = ~new_P2_U5514 | ~new_P2_U2409;
  assign new_P2_U5564 = ~new_P2_U2400 | ~new_P2_U5530;
  assign new_P2_U5565 = ~P2_INSTQUEUE_REG_0__1_ | ~new_P2_U5525;
  assign new_P2_U5566 = ~new_P2_U5515 | ~new_P2_U2431;
  assign new_P2_U5567 = ~new_P2_U2510 | ~new_P2_U2408;
  assign new_P2_U5568 = ~new_P2_U5514 | ~new_P2_U2407;
  assign new_P2_U5569 = ~new_P2_U2399 | ~new_P2_U5530;
  assign new_P2_U5570 = ~P2_INSTQUEUE_REG_0__0_ | ~new_P2_U5525;
  assign new_P2_U5571 = ~new_P2_U3279 | ~new_P2_U7869;
  assign new_P2_U5572 = ~new_P2_U3574;
  assign new_P2_U5573 = ~new_P2_U7861 | ~new_P2_U7863 | ~new_P2_U2617;
  assign new_P2_U5574 = ~new_P2_U3289 | ~new_P2_U3255 | ~new_P2_U7895 | ~new_P2_U3521;
  assign new_P2_U5575 = ~new_P2_U2357 | ~new_P2_U7871;
  assign new_P2_U5576 = ~new_P2_U4417 | ~new_P2_U3574;
  assign new_P2_U5577 = ~new_P2_U4428 | ~new_P2_U4424;
  assign new_P2_U5578 = ~new_P2_U3524 | ~new_P2_U5577;
  assign new_P2_U5579 = ~new_P2_R2088_U6 | ~new_P2_U5578 | ~new_P2_U3265;
  assign new_P2_U5580 = ~new_P2_U4436 | ~new_P2_R2167_U6;
  assign new_P2_U5581 = ~new_P2_U4406;
  assign new_P2_U5582 = ~new_P2_U2374 | ~new_P2_U4406;
  assign new_P2_U5583 = ~P2_STATE2_REG_3_ | ~new_P2_U3284;
  assign new_P2_U5584 = ~new_P2_U4394;
  assign new_P2_U5585 = ~new_P2_U4591 | ~new_P2_U3276;
  assign new_P2_U5586 = ~new_P2_U3878 | ~new_P2_U2617 | ~new_P2_U3295;
  assign new_P2_U5587 = ~new_P2_U3295 | ~new_P2_U3255;
  assign new_P2_U5588 = ~new_P2_U7865 | ~new_P2_U3278;
  assign new_P2_U5589 = ~new_P2_U3879 | ~new_P2_U8075 | ~new_P2_U8074;
  assign new_P2_U5590 = ~new_P2_U3525;
  assign new_P2_U5591 = ~new_P2_U7738 | ~new_P2_U3278;
  assign new_P2_U5592 = ~new_P2_U5571 | ~new_P2_U5573 | ~new_P2_U3521 | ~new_P2_U5591;
  assign new_P2_U5593 = ~new_P2_U4417 | ~new_P2_U3574;
  assign new_P2_U5594 = ~new_P2_U5592 | ~new_P2_U2616;
  assign new_P2_U5595 = ~new_P2_U3877 | ~new_P2_U5594;
  assign new_P2_U5596 = ~new_P2_U3295 | ~new_P2_U7873;
  assign new_P2_U5597 = ~new_P2_U3279 | ~new_P2_U7871;
  assign new_P2_U5598 = ~new_P2_U2617 | ~new_P2_U3521;
  assign new_P2_U5599 = ~new_P2_U4427 | ~new_P2_U5598;
  assign new_P2_U5600 = ~new_P2_U5597 | ~new_P2_U3280;
  assign new_P2_U5601 = ~new_P2_U2436 | ~new_P2_U7884;
  assign new_P2_U5602 = ~new_P2_U3527 | ~new_P2_U3278;
  assign new_P2_U5603 = ~new_P2_U2514 | ~new_P2_U3288;
  assign new_P2_U5604 = ~new_P2_U4470 | ~new_P2_U8077 | ~new_P2_U8076;
  assign new_P2_U5605 = ~new_P2_U3296 | ~new_P2_U3522;
  assign new_P2_U5606 = ~new_P2_U3578 | ~new_P2_U4437;
  assign new_P2_U5607 = ~new_P2_U4395 | ~new_P2_U5605;
  assign new_P2_U5608 = ~new_P2_U3581 | ~new_P2_U5606;
  assign new_P2_U5609 = ~new_P2_R2147_U8 | ~new_P2_U5604;
  assign new_P2_U5610 = ~new_P2_R2099_U95 | ~new_P2_U5603;
  assign new_P2_U5611 = ~new_P2_U3884 | ~new_P2_U5610;
  assign new_P2_U5612 = ~new_P2_R2182_U76 | ~new_P2_U4469;
  assign new_P2_U5613 = ~new_P2_U4466 | ~new_P2_U5611;
  assign new_P2_U5614 = ~new_P2_U5613 | ~new_P2_U5612;
  assign new_P2_U5615 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U4591;
  assign new_P2_U5616 = ~new_P2_U3530;
  assign new_P2_U5617 = ~new_P2_R2147_U9 | ~new_P2_U5604;
  assign new_P2_U5618 = ~new_P2_R2099_U96 | ~new_P2_U5603;
  assign new_P2_U5619 = ~new_P2_U3885 | ~new_P2_U5618;
  assign new_P2_U5620 = ~P2_STATE2_REG_1_ | ~new_P2_U3598 | ~new_P2_U3597;
  assign new_P2_U5621 = ~new_P2_R2182_U40 | ~new_P2_U4469;
  assign new_P2_U5622 = ~new_P2_U4466 | ~new_P2_U5619;
  assign new_P2_U5623 = ~new_P2_U5620 | ~new_P2_U5621 | ~new_P2_U5622;
  assign new_P2_U5624 = ~new_P2_U4429 | ~new_P2_U2449 | ~new_P2_U7861;
  assign new_P2_U5625 = ~new_P2_U7882 | ~new_P2_U5624;
  assign new_P2_U5626 = ~new_P2_U3887 | ~new_P2_U8097;
  assign new_P2_U5627 = ~new_P2_R2147_U4 | ~new_P2_U5604;
  assign new_P2_U5628 = ~new_P2_R2099_U5 | ~new_P2_U5603;
  assign new_P2_U5629 = ~new_P2_U3888 | ~new_P2_U5628;
  assign new_P2_U5630 = ~new_P2_U3597 | ~P2_STATE2_REG_1_ | ~new_P2_U8090;
  assign new_P2_U5631 = ~new_P2_R2182_U68 | ~new_P2_U4469;
  assign new_P2_U5632 = ~new_P2_U4466 | ~new_P2_U5629;
  assign new_P2_U5633 = ~new_P2_U5630 | ~new_P2_U5631 | ~new_P2_U5632;
  assign new_P2_U5634 = ~new_P2_U3889 | ~new_P2_U8097;
  assign new_P2_U5635 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_U5604;
  assign new_P2_U5636 = ~new_P2_R2099_U94 | ~new_P2_U5603;
  assign new_P2_U5637 = ~new_P2_U3890 | ~new_P2_U5636;
  assign new_P2_U5638 = ~new_P2_R2182_U69 | ~new_P2_U4469;
  assign new_P2_U5639 = ~new_P2_U4466 | ~new_P2_U5637;
  assign new_P2_U5640 = ~new_P2_U8087 | ~P2_STATE2_REG_1_;
  assign new_P2_U5641 = ~new_P2_U5640 | ~new_P2_U5639 | ~new_P2_U5638;
  assign new_P2_U5642 = ~new_P2_R2243_U8 | ~new_P2_U2448 | ~P2_STATE2_REG_0_;
  assign new_P2_U5643 = ~new_P2_U3533;
  assign new_P2_U5644 = ~new_P2_U4445 | ~new_P2_U3303;
  assign new_P2_U5645 = ~new_P2_U4636 | ~new_P2_U3579;
  assign new_P2_U5646 = ~new_P2_U3426 | ~new_P2_U5645;
  assign new_P2_U5647 = ~new_P2_U3427 | ~new_P2_U5646;
  assign new_P2_U5648 = ~new_P2_U2398 | ~new_P2_U5647;
  assign new_P2_U5649 = ~new_P2_R2182_U76 | ~new_P2_U5644;
  assign new_P2_U5650 = ~new_P2_R2096_U75 | ~P2_STATE2_REG_3_;
  assign new_P2_U5651 = ~new_P2_U3891 | ~new_P2_U5648;
  assign new_P2_U5652 = ~new_P2_U2398 | ~new_P2_U8109;
  assign new_P2_U5653 = ~new_P2_R2182_U40 | ~new_P2_U5644;
  assign new_P2_U5654 = ~new_P2_R2096_U77 | ~P2_STATE2_REG_3_;
  assign new_P2_U5655 = ~new_P2_U3892 | ~new_P2_U5652;
  assign new_P2_U5656 = ~new_P2_U3338 | ~new_P2_U3353;
  assign new_P2_U5657 = ~new_P2_U2398 | ~new_P2_U5656;
  assign new_P2_U5658 = ~new_P2_R2182_U68 | ~new_P2_U5644;
  assign new_P2_U5659 = ~new_P2_R2096_U51 | ~P2_STATE2_REG_3_;
  assign new_P2_U5660 = ~new_P2_U3893 | ~new_P2_U5657;
  assign new_P2_U5661 = ~new_P2_U3313 | ~new_P2_U3303;
  assign new_P2_U5662 = ~new_P2_R2182_U69 | ~new_P2_U5661;
  assign new_P2_U5663 = ~new_P2_R2096_U68 | ~P2_STATE2_REG_3_;
  assign new_P2_U5664 = ~new_P2_U4464 | ~new_P2_U5662 | ~new_P2_U5663;
  assign new_P2_U5665 = ~new_P2_U2616 | ~new_P2_U3292;
  assign new_P2_U5666 = ~new_P2_GTE_370_U6 | ~new_P2_U4417;
  assign new_P2_U5667 = ~new_P2_U5666 | ~new_P2_U5665;
  assign new_P2_U5668 = ~new_P2_R2088_U6 | ~new_P2_U3265 | ~new_P2_U8122 | ~new_P2_U8121;
  assign new_P2_U5669 = ~new_P2_U4420 | ~new_P2_U5667;
  assign new_P2_U5670 = ~new_P2_U5669 | ~new_P2_U4397 | ~new_P2_U2512 | ~new_P2_U3894;
  assign new_P2_U5671 = ~new_P2_U2374 | ~new_P2_U5670;
  assign new_P2_U5672 = ~new_P2_U4461 | ~new_P2_U3284;
  assign new_P2_U5673 = ~new_P2_U3535;
  assign new_P2_U5674 = ~new_P2_U4427 | ~new_P2_U4420;
  assign new_P2_U5675 = ~new_P2_U3895 | ~new_P2_U2514;
  assign new_P2_U5676 = ~new_P2_U4417 | ~new_P2_U4424;
  assign new_P2_U5677 = ~new_P2_U3524 | ~new_P2_U4437 | ~new_P2_U5676 | ~new_P2_U4470;
  assign new_P2_U5678 = ~new_P2_U4428 | ~new_P2_U4424;
  assign new_P2_U5679 = ~new_P2_U3523 | ~new_P2_U3296 | ~new_P2_U5678;
  assign new_P2_U5680 = ~new_P2_U2390 | ~new_P2_R2096_U68;
  assign new_P2_U5681 = ~new_P2_U2389 | ~new_P2_R2099_U94;
  assign new_P2_U5682 = ~new_P2_R2027_U5 | ~new_P2_U2388;
  assign new_P2_U5683 = ~new_P2_ADD_394_U4 | ~new_P2_U2386;
  assign new_P2_U5684 = ~new_P2_R2278_U83 | ~new_P2_U2385;
  assign new_P2_U5685 = ~new_P2_ADD_371_1212_U68 | ~new_P2_U2384;
  assign new_P2_U5686 = ~P2_REIP_REG_0_ | ~new_P2_U2381;
  assign new_P2_U5687 = ~new_P2_U5673 | ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_U5688 = ~new_P2_U2390 | ~new_P2_R2096_U51;
  assign new_P2_U5689 = ~new_P2_U2389 | ~new_P2_R2099_U5;
  assign new_P2_U5690 = ~new_P2_R2027_U85 | ~new_P2_U2388;
  assign new_P2_U5691 = ~new_P2_ADD_394_U85 | ~new_P2_U2386;
  assign new_P2_U5692 = ~new_P2_R2278_U6 | ~new_P2_U2385;
  assign new_P2_U5693 = ~new_P2_ADD_371_1212_U25 | ~new_P2_U2384;
  assign new_P2_U5694 = ~new_P2_U2381 | ~P2_REIP_REG_1_;
  assign new_P2_U5695 = ~new_P2_U5673 | ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_U5696 = ~new_P2_U2390 | ~new_P2_R2096_U77;
  assign new_P2_U5697 = ~new_P2_U2389 | ~new_P2_R2099_U96;
  assign new_P2_U5698 = ~new_P2_R2027_U74 | ~new_P2_U2388;
  assign new_P2_U5699 = ~new_P2_ADD_394_U5 | ~new_P2_U2386;
  assign new_P2_U5700 = ~new_P2_R2278_U92 | ~new_P2_U2385;
  assign new_P2_U5701 = ~new_P2_ADD_371_1212_U79 | ~new_P2_U2384;
  assign new_P2_U5702 = ~new_P2_U2381 | ~P2_REIP_REG_2_;
  assign new_P2_U5703 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_U5673;
  assign new_P2_U5704 = ~new_P2_U2390 | ~new_P2_R2096_U75;
  assign new_P2_U5705 = ~new_P2_U2389 | ~new_P2_R2099_U95;
  assign new_P2_U5706 = ~new_P2_R2027_U71 | ~new_P2_U2388;
  assign new_P2_U5707 = ~new_P2_ADD_394_U95 | ~new_P2_U2386;
  assign new_P2_U5708 = ~new_P2_R2278_U90 | ~new_P2_U2385;
  assign new_P2_U5709 = ~new_P2_ADD_371_1212_U84 | ~new_P2_U2384;
  assign new_P2_U5710 = ~new_P2_U2381 | ~P2_REIP_REG_3_;
  assign new_P2_U5711 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_U5673;
  assign new_P2_U5712 = ~new_P2_R2096_U74 | ~new_P2_U2390;
  assign new_P2_U5713 = ~new_P2_R2099_U98 | ~new_P2_U2389;
  assign new_P2_U5714 = ~new_P2_R2027_U70 | ~new_P2_U2388;
  assign new_P2_U5715 = ~new_P2_ADD_394_U76 | ~new_P2_U2386;
  assign new_P2_U5716 = ~new_P2_R2278_U89 | ~new_P2_U2385;
  assign new_P2_U5717 = ~new_P2_ADD_371_1212_U80 | ~new_P2_U2384;
  assign new_P2_U5718 = ~new_P2_U2381 | ~P2_REIP_REG_4_;
  assign new_P2_U5719 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_U5673;
  assign new_P2_U5720 = ~new_P2_R2096_U73 | ~new_P2_U2390;
  assign new_P2_U5721 = ~new_P2_R2099_U71 | ~new_P2_U2389;
  assign new_P2_U5722 = ~new_P2_R2027_U69 | ~new_P2_U2388;
  assign new_P2_U5723 = ~new_P2_ADD_394_U79 | ~new_P2_U2386;
  assign new_P2_U5724 = ~new_P2_R2278_U88 | ~new_P2_U2385;
  assign new_P2_U5725 = ~new_P2_ADD_371_1212_U81 | ~new_P2_U2384;
  assign new_P2_U5726 = ~new_P2_U2381 | ~P2_REIP_REG_5_;
  assign new_P2_U5727 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_U5673;
  assign new_P2_U5728 = ~new_P2_R2096_U72 | ~new_P2_U2390;
  assign new_P2_U5729 = ~new_P2_R2099_U70 | ~new_P2_U2389;
  assign new_P2_U5730 = ~new_P2_R2027_U68 | ~new_P2_U2388;
  assign new_P2_U5731 = ~new_P2_ADD_394_U63 | ~new_P2_U2386;
  assign new_P2_U5732 = ~new_P2_R2278_U87 | ~new_P2_U2385;
  assign new_P2_U5733 = ~new_P2_ADD_371_1212_U78 | ~new_P2_U2384;
  assign new_P2_U5734 = ~new_P2_U2381 | ~P2_REIP_REG_6_;
  assign new_P2_U5735 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_U5673;
  assign new_P2_U5736 = ~new_P2_R2096_U71 | ~new_P2_U2390;
  assign new_P2_U5737 = ~new_P2_R2099_U69 | ~new_P2_U2389;
  assign new_P2_U5738 = ~new_P2_R2027_U67 | ~new_P2_U2388;
  assign new_P2_U5739 = ~new_P2_ADD_394_U89 | ~new_P2_U2386;
  assign new_P2_U5740 = ~new_P2_R2278_U86 | ~new_P2_U2385;
  assign new_P2_U5741 = ~new_P2_ADD_371_1212_U85 | ~new_P2_U2384;
  assign new_P2_U5742 = ~new_P2_U2381 | ~P2_REIP_REG_7_;
  assign new_P2_U5743 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_U5673;
  assign new_P2_U5744 = ~new_P2_R2096_U70 | ~new_P2_U2390;
  assign new_P2_U5745 = ~new_P2_R2099_U68 | ~new_P2_U2389;
  assign new_P2_U5746 = ~new_P2_R2027_U66 | ~new_P2_U2388;
  assign new_P2_U5747 = ~new_P2_ADD_394_U80 | ~new_P2_U2386;
  assign new_P2_U5748 = ~new_P2_R2278_U85 | ~new_P2_U2385;
  assign new_P2_U5749 = ~new_P2_ADD_371_1212_U82 | ~new_P2_U2384;
  assign new_P2_U5750 = ~new_P2_U2381 | ~P2_REIP_REG_8_;
  assign new_P2_U5751 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_U5673;
  assign new_P2_U5752 = ~new_P2_R2096_U69 | ~new_P2_U2390;
  assign new_P2_U5753 = ~new_P2_R2099_U67 | ~new_P2_U2389;
  assign new_P2_U5754 = ~new_P2_R2027_U65 | ~new_P2_U2388;
  assign new_P2_U5755 = ~new_P2_ADD_394_U70 | ~new_P2_U2386;
  assign new_P2_U5756 = ~new_P2_R2278_U84 | ~new_P2_U2385;
  assign new_P2_U5757 = ~new_P2_ADD_371_1212_U118 | ~new_P2_U2384;
  assign new_P2_U5758 = ~new_P2_U2381 | ~P2_REIP_REG_9_;
  assign new_P2_U5759 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_U5673;
  assign new_P2_U5760 = ~new_P2_R2096_U97 | ~new_P2_U2390;
  assign new_P2_U5761 = ~new_P2_R2099_U93 | ~new_P2_U2389;
  assign new_P2_U5762 = ~new_P2_R2027_U95 | ~new_P2_U2388;
  assign new_P2_U5763 = ~new_P2_ADD_394_U83 | ~new_P2_U2386;
  assign new_P2_U5764 = ~new_P2_R2278_U112 | ~new_P2_U2385;
  assign new_P2_U5765 = ~new_P2_ADD_371_1212_U13 | ~new_P2_U2384;
  assign new_P2_U5766 = ~new_P2_U2381 | ~P2_REIP_REG_10_;
  assign new_P2_U5767 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_U5673;
  assign new_P2_U5768 = ~new_P2_R2096_U96 | ~new_P2_U2390;
  assign new_P2_U5769 = ~new_P2_R2099_U92 | ~new_P2_U2389;
  assign new_P2_U5770 = ~new_P2_R2027_U94 | ~new_P2_U2388;
  assign new_P2_U5771 = ~new_P2_ADD_394_U73 | ~new_P2_U2386;
  assign new_P2_U5772 = ~new_P2_R2278_U111 | ~new_P2_U2385;
  assign new_P2_U5773 = ~new_P2_ADD_371_1212_U14 | ~new_P2_U2384;
  assign new_P2_U5774 = ~new_P2_U2381 | ~P2_REIP_REG_11_;
  assign new_P2_U5775 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_U5673;
  assign new_P2_U5776 = ~new_P2_R2096_U95 | ~new_P2_U2390;
  assign new_P2_U5777 = ~new_P2_R2099_U91 | ~new_P2_U2389;
  assign new_P2_U5778 = ~new_P2_R2027_U93 | ~new_P2_U2388;
  assign new_P2_U5779 = ~new_P2_ADD_394_U88 | ~new_P2_U2386;
  assign new_P2_U5780 = ~new_P2_R2278_U110 | ~new_P2_U2385;
  assign new_P2_U5781 = ~new_P2_ADD_371_1212_U76 | ~new_P2_U2384;
  assign new_P2_U5782 = ~new_P2_U2381 | ~P2_REIP_REG_12_;
  assign new_P2_U5783 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_U5673;
  assign new_P2_U5784 = ~new_P2_R2096_U94 | ~new_P2_U2390;
  assign new_P2_U5785 = ~new_P2_R2099_U90 | ~new_P2_U2389;
  assign new_P2_U5786 = ~new_P2_R2027_U92 | ~new_P2_U2388;
  assign new_P2_U5787 = ~new_P2_ADD_394_U69 | ~new_P2_U2386;
  assign new_P2_U5788 = ~new_P2_R2278_U109 | ~new_P2_U2385;
  assign new_P2_U5789 = ~new_P2_ADD_371_1212_U15 | ~new_P2_U2384;
  assign new_P2_U5790 = ~new_P2_U2381 | ~P2_REIP_REG_13_;
  assign new_P2_U5791 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_U5673;
  assign new_P2_U5792 = ~new_P2_R2096_U93 | ~new_P2_U2390;
  assign new_P2_U5793 = ~new_P2_R2099_U89 | ~new_P2_U2389;
  assign new_P2_U5794 = ~new_P2_R2027_U91 | ~new_P2_U2388;
  assign new_P2_U5795 = ~new_P2_ADD_394_U78 | ~new_P2_U2386;
  assign new_P2_U5796 = ~new_P2_R2278_U108 | ~new_P2_U2385;
  assign new_P2_U5797 = ~new_P2_ADD_371_1212_U16 | ~new_P2_U2384;
  assign new_P2_U5798 = ~new_P2_U2381 | ~P2_REIP_REG_14_;
  assign new_P2_U5799 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_U5673;
  assign new_P2_U5800 = ~new_P2_R2096_U92 | ~new_P2_U2390;
  assign new_P2_U5801 = ~new_P2_R2099_U88 | ~new_P2_U2389;
  assign new_P2_U5802 = ~new_P2_R2027_U90 | ~new_P2_U2388;
  assign new_P2_U5803 = ~new_P2_ADD_394_U75 | ~new_P2_U2386;
  assign new_P2_U5804 = ~new_P2_R2278_U107 | ~new_P2_U2385;
  assign new_P2_U5805 = ~new_P2_ADD_371_1212_U73 | ~new_P2_U2384;
  assign new_P2_U5806 = ~new_P2_U2381 | ~P2_REIP_REG_15_;
  assign new_P2_U5807 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_U5673;
  assign new_P2_U5808 = ~new_P2_R2096_U91 | ~new_P2_U2390;
  assign new_P2_U5809 = ~new_P2_R2099_U87 | ~new_P2_U2389;
  assign new_P2_U5810 = ~new_P2_R2027_U89 | ~new_P2_U2388;
  assign new_P2_U5811 = ~new_P2_ADD_394_U91 | ~new_P2_U2386;
  assign new_P2_U5812 = ~new_P2_R2278_U106 | ~new_P2_U2385;
  assign new_P2_U5813 = ~new_P2_ADD_371_1212_U17 | ~new_P2_U2384;
  assign new_P2_U5814 = ~new_P2_U2381 | ~P2_REIP_REG_16_;
  assign new_P2_U5815 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_U5673;
  assign new_P2_U5816 = ~new_P2_R2096_U90 | ~new_P2_U2390;
  assign new_P2_U5817 = ~new_P2_R2099_U86 | ~new_P2_U2389;
  assign new_P2_U5818 = ~new_P2_R2027_U88 | ~new_P2_U2388;
  assign new_P2_U5819 = ~new_P2_ADD_394_U67 | ~new_P2_U2386;
  assign new_P2_U5820 = ~new_P2_R2278_U105 | ~new_P2_U2385;
  assign new_P2_U5821 = ~new_P2_ADD_371_1212_U71 | ~new_P2_U2384;
  assign new_P2_U5822 = ~new_P2_U2381 | ~P2_REIP_REG_17_;
  assign new_P2_U5823 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_U5673;
  assign new_P2_U5824 = ~new_P2_R2096_U89 | ~new_P2_U2390;
  assign new_P2_U5825 = ~new_P2_R2099_U85 | ~new_P2_U2389;
  assign new_P2_U5826 = ~new_P2_R2027_U87 | ~new_P2_U2388;
  assign new_P2_U5827 = ~new_P2_ADD_394_U72 | ~new_P2_U2386;
  assign new_P2_U5828 = ~new_P2_R2278_U104 | ~new_P2_U2385;
  assign new_P2_U5829 = ~new_P2_ADD_371_1212_U72 | ~new_P2_U2384;
  assign new_P2_U5830 = ~new_P2_U2381 | ~P2_REIP_REG_18_;
  assign new_P2_U5831 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_U5673;
  assign new_P2_U5832 = ~new_P2_R2096_U88 | ~new_P2_U2390;
  assign new_P2_U5833 = ~new_P2_R2099_U84 | ~new_P2_U2389;
  assign new_P2_U5834 = ~new_P2_R2027_U86 | ~new_P2_U2388;
  assign new_P2_U5835 = ~new_P2_ADD_394_U82 | ~new_P2_U2386;
  assign new_P2_U5836 = ~new_P2_R2278_U103 | ~new_P2_U2385;
  assign new_P2_U5837 = ~new_P2_ADD_371_1212_U18 | ~new_P2_U2384;
  assign new_P2_U5838 = ~new_P2_U2381 | ~P2_REIP_REG_19_;
  assign new_P2_U5839 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_U5673;
  assign new_P2_U5840 = ~new_P2_R2096_U87 | ~new_P2_U2390;
  assign new_P2_U5841 = ~new_P2_R2099_U83 | ~new_P2_U2389;
  assign new_P2_U5842 = ~new_P2_R2027_U84 | ~new_P2_U2388;
  assign new_P2_U5843 = ~new_P2_ADD_394_U68 | ~new_P2_U2386;
  assign new_P2_U5844 = ~new_P2_R2278_U102 | ~new_P2_U2385;
  assign new_P2_U5845 = ~new_P2_ADD_371_1212_U19 | ~new_P2_U2384;
  assign new_P2_U5846 = ~new_P2_U2381 | ~P2_REIP_REG_20_;
  assign new_P2_U5847 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_U5673;
  assign new_P2_U5848 = ~new_P2_R2096_U86 | ~new_P2_U2390;
  assign new_P2_U5849 = ~new_P2_R2099_U82 | ~new_P2_U2389;
  assign new_P2_U5850 = ~new_P2_R2027_U83 | ~new_P2_U2388;
  assign new_P2_U5851 = ~new_P2_ADD_394_U87 | ~new_P2_U2386;
  assign new_P2_U5852 = ~new_P2_R2278_U101 | ~new_P2_U2385;
  assign new_P2_U5853 = ~new_P2_ADD_371_1212_U75 | ~new_P2_U2384;
  assign new_P2_U5854 = ~new_P2_U2381 | ~P2_REIP_REG_21_;
  assign new_P2_U5855 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_U5673;
  assign new_P2_U5856 = ~new_P2_R2096_U85 | ~new_P2_U2390;
  assign new_P2_U5857 = ~new_P2_R2099_U81 | ~new_P2_U2389;
  assign new_P2_U5858 = ~new_P2_R2027_U82 | ~new_P2_U2388;
  assign new_P2_U5859 = ~new_P2_ADD_394_U71 | ~new_P2_U2386;
  assign new_P2_U5860 = ~new_P2_R2278_U100 | ~new_P2_U2385;
  assign new_P2_U5861 = ~new_P2_ADD_371_1212_U20 | ~new_P2_U2384;
  assign new_P2_U5862 = ~new_P2_U2381 | ~P2_REIP_REG_22_;
  assign new_P2_U5863 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_U5673;
  assign new_P2_U5864 = ~new_P2_R2096_U84 | ~new_P2_U2390;
  assign new_P2_U5865 = ~new_P2_R2099_U80 | ~new_P2_U2389;
  assign new_P2_U5866 = ~new_P2_R2027_U81 | ~new_P2_U2388;
  assign new_P2_U5867 = ~new_P2_ADD_394_U81 | ~new_P2_U2386;
  assign new_P2_U5868 = ~new_P2_R2278_U99 | ~new_P2_U2385;
  assign new_P2_U5869 = ~new_P2_ADD_371_1212_U21 | ~new_P2_U2384;
  assign new_P2_U5870 = ~new_P2_U2381 | ~P2_REIP_REG_23_;
  assign new_P2_U5871 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_U5673;
  assign new_P2_U5872 = ~new_P2_R2096_U83 | ~new_P2_U2390;
  assign new_P2_U5873 = ~new_P2_R2099_U79 | ~new_P2_U2389;
  assign new_P2_U5874 = ~new_P2_R2027_U80 | ~new_P2_U2388;
  assign new_P2_U5875 = ~new_P2_ADD_394_U66 | ~new_P2_U2386;
  assign new_P2_U5876 = ~new_P2_R2278_U98 | ~new_P2_U2385;
  assign new_P2_U5877 = ~new_P2_ADD_371_1212_U70 | ~new_P2_U2384;
  assign new_P2_U5878 = ~new_P2_U2381 | ~P2_REIP_REG_24_;
  assign new_P2_U5879 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_U5673;
  assign new_P2_U5880 = ~new_P2_R2096_U82 | ~new_P2_U2390;
  assign new_P2_U5881 = ~new_P2_R2099_U78 | ~new_P2_U2389;
  assign new_P2_U5882 = ~new_P2_R2027_U79 | ~new_P2_U2388;
  assign new_P2_U5883 = ~new_P2_ADD_394_U90 | ~new_P2_U2386;
  assign new_P2_U5884 = ~new_P2_R2278_U97 | ~new_P2_U2385;
  assign new_P2_U5885 = ~new_P2_ADD_371_1212_U77 | ~new_P2_U2384;
  assign new_P2_U5886 = ~new_P2_U2381 | ~P2_REIP_REG_25_;
  assign new_P2_U5887 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_U5673;
  assign new_P2_U5888 = ~new_P2_R2096_U81 | ~new_P2_U2390;
  assign new_P2_U5889 = ~new_P2_R2099_U77 | ~new_P2_U2389;
  assign new_P2_U5890 = ~new_P2_R2027_U78 | ~new_P2_U2388;
  assign new_P2_U5891 = ~new_P2_ADD_394_U74 | ~new_P2_U2386;
  assign new_P2_U5892 = ~new_P2_R2278_U96 | ~new_P2_U2385;
  assign new_P2_U5893 = ~new_P2_ADD_371_1212_U22 | ~new_P2_U2384;
  assign new_P2_U5894 = ~new_P2_U2381 | ~P2_REIP_REG_26_;
  assign new_P2_U5895 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_U5673;
  assign new_P2_U5896 = ~new_P2_R2096_U80 | ~new_P2_U2390;
  assign new_P2_U5897 = ~new_P2_R2099_U76 | ~new_P2_U2389;
  assign new_P2_U5898 = ~new_P2_R2027_U77 | ~new_P2_U2388;
  assign new_P2_U5899 = ~new_P2_ADD_394_U77 | ~new_P2_U2386;
  assign new_P2_U5900 = ~new_P2_R2278_U95 | ~new_P2_U2385;
  assign new_P2_U5901 = ~new_P2_ADD_371_1212_U74 | ~new_P2_U2384;
  assign new_P2_U5902 = ~new_P2_U2381 | ~P2_REIP_REG_27_;
  assign new_P2_U5903 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_U5673;
  assign new_P2_U5904 = ~new_P2_R2096_U79 | ~new_P2_U2390;
  assign new_P2_U5905 = ~new_P2_R2099_U75 | ~new_P2_U2389;
  assign new_P2_U5906 = ~new_P2_R2027_U76 | ~new_P2_U2388;
  assign new_P2_U5907 = ~new_P2_ADD_394_U86 | ~new_P2_U2386;
  assign new_P2_U5908 = ~new_P2_R2278_U94 | ~new_P2_U2385;
  assign new_P2_U5909 = ~new_P2_ADD_371_1212_U23 | ~new_P2_U2384;
  assign new_P2_U5910 = ~new_P2_U2381 | ~P2_REIP_REG_28_;
  assign new_P2_U5911 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_U5673;
  assign new_P2_U5912 = ~new_P2_R2096_U78 | ~new_P2_U2390;
  assign new_P2_U5913 = ~new_P2_R2099_U74 | ~new_P2_U2389;
  assign new_P2_U5914 = ~new_P2_R2027_U75 | ~new_P2_U2388;
  assign new_P2_U5915 = ~new_P2_ADD_394_U65 | ~new_P2_U2386;
  assign new_P2_U5916 = ~new_P2_R2278_U93 | ~new_P2_U2385;
  assign new_P2_U5917 = ~new_P2_ADD_371_1212_U24 | ~new_P2_U2384;
  assign new_P2_U5918 = ~new_P2_U2381 | ~P2_REIP_REG_29_;
  assign new_P2_U5919 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_U5673;
  assign new_P2_U5920 = ~new_P2_R2096_U76 | ~new_P2_U2390;
  assign new_P2_U5921 = ~new_P2_R2099_U73 | ~new_P2_U2389;
  assign new_P2_U5922 = ~new_P2_R2027_U73 | ~new_P2_U2388;
  assign new_P2_U5923 = ~new_P2_ADD_394_U64 | ~new_P2_U2386;
  assign new_P2_U5924 = ~new_P2_R2278_U91 | ~new_P2_U2385;
  assign new_P2_U5925 = ~new_P2_ADD_371_1212_U69 | ~new_P2_U2384;
  assign new_P2_U5926 = ~new_P2_U2381 | ~P2_REIP_REG_30_;
  assign new_P2_U5927 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_U5673;
  assign new_P2_U5928 = ~new_P2_R2096_U50 | ~new_P2_U2390;
  assign new_P2_U5929 = ~new_P2_R2099_U72 | ~new_P2_U2389;
  assign new_P2_U5930 = ~new_P2_R2027_U72 | ~new_P2_U2388;
  assign new_P2_U5931 = ~new_P2_ADD_394_U84 | ~new_P2_U2386;
  assign new_P2_U5932 = ~new_P2_R2278_U5 | ~new_P2_U2385;
  assign new_P2_U5933 = ~new_P2_ADD_371_1212_U83 | ~new_P2_U2384;
  assign new_P2_U5934 = ~new_P2_U2381 | ~P2_REIP_REG_31_;
  assign new_P2_U5935 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_U5673;
  assign new_P2_U5936 = ~new_P2_U4613 | ~new_P2_U4420 | ~new_P2_U2374;
  assign new_P2_U5937 = ~new_P2_U5661 | ~new_P2_U3284;
  assign new_P2_U5938 = ~new_P2_U3537;
  assign new_P2_U5939 = ~P2_STATE2_REG_1_ | ~new_P2_U3302;
  assign new_P2_U5940 = ~new_P2_U3540 | ~new_P2_U5939;
  assign new_P2_U5941 = ~P2_PHYADDRPOINTER_REG_0_ | ~new_P2_U2387;
  assign new_P2_U5942 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U68;
  assign new_P2_U5943 = ~new_P2_U2372 | ~new_P2_R2099_U94;
  assign new_P2_U5944 = ~new_P2_U2371 | ~P2_REIP_REG_0_;
  assign new_P2_U5945 = ~new_P2_U2370 | ~new_P2_R2278_U83;
  assign new_P2_U5946 = ~P2_PHYADDRPOINTER_REG_0_ | ~new_P2_U5938;
  assign new_P2_U5947 = ~new_P2_R2337_U4 | ~new_P2_U2387;
  assign new_P2_U5948 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U25;
  assign new_P2_U5949 = ~new_P2_U2372 | ~new_P2_R2099_U5;
  assign new_P2_U5950 = ~new_P2_U2371 | ~P2_REIP_REG_1_;
  assign new_P2_U5951 = ~new_P2_U2370 | ~new_P2_R2278_U6;
  assign new_P2_U5952 = ~P2_PHYADDRPOINTER_REG_1_ | ~new_P2_U5938;
  assign new_P2_U5953 = ~new_P2_R2337_U70 | ~new_P2_U2387;
  assign new_P2_U5954 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U79;
  assign new_P2_U5955 = ~new_P2_U2372 | ~new_P2_R2099_U96;
  assign new_P2_U5956 = ~new_P2_U2371 | ~P2_REIP_REG_2_;
  assign new_P2_U5957 = ~new_P2_U2370 | ~new_P2_R2278_U92;
  assign new_P2_U5958 = ~P2_PHYADDRPOINTER_REG_2_ | ~new_P2_U5938;
  assign new_P2_U5959 = ~new_P2_R2337_U67 | ~new_P2_U2387;
  assign new_P2_U5960 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U84;
  assign new_P2_U5961 = ~new_P2_U2372 | ~new_P2_R2099_U95;
  assign new_P2_U5962 = ~new_P2_U2371 | ~P2_REIP_REG_3_;
  assign new_P2_U5963 = ~new_P2_U2370 | ~new_P2_R2278_U90;
  assign new_P2_U5964 = ~P2_PHYADDRPOINTER_REG_3_ | ~new_P2_U5938;
  assign new_P2_U5965 = ~new_P2_R2337_U66 | ~new_P2_U2387;
  assign new_P2_U5966 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U80;
  assign new_P2_U5967 = ~new_P2_U2372 | ~new_P2_R2099_U98;
  assign new_P2_U5968 = ~new_P2_U2371 | ~P2_REIP_REG_4_;
  assign new_P2_U5969 = ~new_P2_U2370 | ~new_P2_R2278_U89;
  assign new_P2_U5970 = ~P2_PHYADDRPOINTER_REG_4_ | ~new_P2_U5938;
  assign new_P2_U5971 = ~new_P2_R2337_U65 | ~new_P2_U2387;
  assign new_P2_U5972 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U81;
  assign new_P2_U5973 = ~new_P2_U2372 | ~new_P2_R2099_U71;
  assign new_P2_U5974 = ~new_P2_U2371 | ~P2_REIP_REG_5_;
  assign new_P2_U5975 = ~new_P2_U2370 | ~new_P2_R2278_U88;
  assign new_P2_U5976 = ~P2_PHYADDRPOINTER_REG_5_ | ~new_P2_U5938;
  assign new_P2_U5977 = ~new_P2_R2337_U64 | ~new_P2_U2387;
  assign new_P2_U5978 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U78;
  assign new_P2_U5979 = ~new_P2_U2372 | ~new_P2_R2099_U70;
  assign new_P2_U5980 = ~new_P2_U2371 | ~P2_REIP_REG_6_;
  assign new_P2_U5981 = ~new_P2_U2370 | ~new_P2_R2278_U87;
  assign new_P2_U5982 = ~P2_PHYADDRPOINTER_REG_6_ | ~new_P2_U5938;
  assign new_P2_U5983 = ~new_P2_R2337_U63 | ~new_P2_U2387;
  assign new_P2_U5984 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U85;
  assign new_P2_U5985 = ~new_P2_U2372 | ~new_P2_R2099_U69;
  assign new_P2_U5986 = ~new_P2_U2371 | ~P2_REIP_REG_7_;
  assign new_P2_U5987 = ~new_P2_U2370 | ~new_P2_R2278_U86;
  assign new_P2_U5988 = ~P2_PHYADDRPOINTER_REG_7_ | ~new_P2_U5938;
  assign new_P2_U5989 = ~new_P2_R2337_U62 | ~new_P2_U2387;
  assign new_P2_U5990 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U82;
  assign new_P2_U5991 = ~new_P2_U2372 | ~new_P2_R2099_U68;
  assign new_P2_U5992 = ~new_P2_U2371 | ~P2_REIP_REG_8_;
  assign new_P2_U5993 = ~new_P2_U2370 | ~new_P2_R2278_U85;
  assign new_P2_U5994 = ~P2_PHYADDRPOINTER_REG_8_ | ~new_P2_U5938;
  assign new_P2_U5995 = ~new_P2_R2337_U61 | ~new_P2_U2387;
  assign new_P2_U5996 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U118;
  assign new_P2_U5997 = ~new_P2_U2372 | ~new_P2_R2099_U67;
  assign new_P2_U5998 = ~new_P2_U2371 | ~P2_REIP_REG_9_;
  assign new_P2_U5999 = ~new_P2_U2370 | ~new_P2_R2278_U84;
  assign new_P2_U6000 = ~P2_PHYADDRPOINTER_REG_9_ | ~new_P2_U5938;
  assign new_P2_U6001 = ~new_P2_R2337_U90 | ~new_P2_U2387;
  assign new_P2_U6002 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U13;
  assign new_P2_U6003 = ~new_P2_U2372 | ~new_P2_R2099_U93;
  assign new_P2_U6004 = ~new_P2_U2371 | ~P2_REIP_REG_10_;
  assign new_P2_U6005 = ~new_P2_U2370 | ~new_P2_R2278_U112;
  assign new_P2_U6006 = ~P2_PHYADDRPOINTER_REG_10_ | ~new_P2_U5938;
  assign new_P2_U6007 = ~new_P2_R2337_U89 | ~new_P2_U2387;
  assign new_P2_U6008 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U14;
  assign new_P2_U6009 = ~new_P2_U2372 | ~new_P2_R2099_U92;
  assign new_P2_U6010 = ~new_P2_U2371 | ~P2_REIP_REG_11_;
  assign new_P2_U6011 = ~new_P2_U2370 | ~new_P2_R2278_U111;
  assign new_P2_U6012 = ~P2_PHYADDRPOINTER_REG_11_ | ~new_P2_U5938;
  assign new_P2_U6013 = ~new_P2_R2337_U88 | ~new_P2_U2387;
  assign new_P2_U6014 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U76;
  assign new_P2_U6015 = ~new_P2_U2372 | ~new_P2_R2099_U91;
  assign new_P2_U6016 = ~new_P2_U2371 | ~P2_REIP_REG_12_;
  assign new_P2_U6017 = ~new_P2_U2370 | ~new_P2_R2278_U110;
  assign new_P2_U6018 = ~P2_PHYADDRPOINTER_REG_12_ | ~new_P2_U5938;
  assign new_P2_U6019 = ~new_P2_R2337_U87 | ~new_P2_U2387;
  assign new_P2_U6020 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U15;
  assign new_P2_U6021 = ~new_P2_U2372 | ~new_P2_R2099_U90;
  assign new_P2_U6022 = ~new_P2_U2371 | ~P2_REIP_REG_13_;
  assign new_P2_U6023 = ~new_P2_U2370 | ~new_P2_R2278_U109;
  assign new_P2_U6024 = ~P2_PHYADDRPOINTER_REG_13_ | ~new_P2_U5938;
  assign new_P2_U6025 = ~new_P2_R2337_U86 | ~new_P2_U2387;
  assign new_P2_U6026 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U16;
  assign new_P2_U6027 = ~new_P2_U2372 | ~new_P2_R2099_U89;
  assign new_P2_U6028 = ~new_P2_U2371 | ~P2_REIP_REG_14_;
  assign new_P2_U6029 = ~new_P2_U2370 | ~new_P2_R2278_U108;
  assign new_P2_U6030 = ~P2_PHYADDRPOINTER_REG_14_ | ~new_P2_U5938;
  assign new_P2_U6031 = ~new_P2_R2337_U85 | ~new_P2_U2387;
  assign new_P2_U6032 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U73;
  assign new_P2_U6033 = ~new_P2_U2372 | ~new_P2_R2099_U88;
  assign new_P2_U6034 = ~new_P2_U2371 | ~P2_REIP_REG_15_;
  assign new_P2_U6035 = ~new_P2_U2370 | ~new_P2_R2278_U107;
  assign new_P2_U6036 = ~P2_PHYADDRPOINTER_REG_15_ | ~new_P2_U5938;
  assign new_P2_U6037 = ~new_P2_R2337_U84 | ~new_P2_U2387;
  assign new_P2_U6038 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U17;
  assign new_P2_U6039 = ~new_P2_U2372 | ~new_P2_R2099_U87;
  assign new_P2_U6040 = ~new_P2_U2371 | ~P2_REIP_REG_16_;
  assign new_P2_U6041 = ~new_P2_U2370 | ~new_P2_R2278_U106;
  assign new_P2_U6042 = ~P2_PHYADDRPOINTER_REG_16_ | ~new_P2_U5938;
  assign new_P2_U6043 = ~new_P2_R2337_U83 | ~new_P2_U2387;
  assign new_P2_U6044 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U71;
  assign new_P2_U6045 = ~new_P2_U2372 | ~new_P2_R2099_U86;
  assign new_P2_U6046 = ~new_P2_U2371 | ~P2_REIP_REG_17_;
  assign new_P2_U6047 = ~new_P2_U2370 | ~new_P2_R2278_U105;
  assign new_P2_U6048 = ~P2_PHYADDRPOINTER_REG_17_ | ~new_P2_U5938;
  assign new_P2_U6049 = ~new_P2_R2337_U82 | ~new_P2_U2387;
  assign new_P2_U6050 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U72;
  assign new_P2_U6051 = ~new_P2_U2372 | ~new_P2_R2099_U85;
  assign new_P2_U6052 = ~new_P2_U2371 | ~P2_REIP_REG_18_;
  assign new_P2_U6053 = ~new_P2_U2370 | ~new_P2_R2278_U104;
  assign new_P2_U6054 = ~P2_PHYADDRPOINTER_REG_18_ | ~new_P2_U5938;
  assign new_P2_U6055 = ~new_P2_R2337_U81 | ~new_P2_U2387;
  assign new_P2_U6056 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U18;
  assign new_P2_U6057 = ~new_P2_U2372 | ~new_P2_R2099_U84;
  assign new_P2_U6058 = ~new_P2_U2371 | ~P2_REIP_REG_19_;
  assign new_P2_U6059 = ~new_P2_U2370 | ~new_P2_R2278_U103;
  assign new_P2_U6060 = ~P2_PHYADDRPOINTER_REG_19_ | ~new_P2_U5938;
  assign new_P2_U6061 = ~new_P2_R2337_U80 | ~new_P2_U2387;
  assign new_P2_U6062 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U19;
  assign new_P2_U6063 = ~new_P2_U2372 | ~new_P2_R2099_U83;
  assign new_P2_U6064 = ~new_P2_U2371 | ~P2_REIP_REG_20_;
  assign new_P2_U6065 = ~new_P2_U2370 | ~new_P2_R2278_U102;
  assign new_P2_U6066 = ~P2_PHYADDRPOINTER_REG_20_ | ~new_P2_U5938;
  assign new_P2_U6067 = ~new_P2_R2337_U79 | ~new_P2_U2387;
  assign new_P2_U6068 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U75;
  assign new_P2_U6069 = ~new_P2_U2372 | ~new_P2_R2099_U82;
  assign new_P2_U6070 = ~new_P2_U2371 | ~P2_REIP_REG_21_;
  assign new_P2_U6071 = ~new_P2_U2370 | ~new_P2_R2278_U101;
  assign new_P2_U6072 = ~P2_PHYADDRPOINTER_REG_21_ | ~new_P2_U5938;
  assign new_P2_U6073 = ~new_P2_R2337_U78 | ~new_P2_U2387;
  assign new_P2_U6074 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U20;
  assign new_P2_U6075 = ~new_P2_U2372 | ~new_P2_R2099_U81;
  assign new_P2_U6076 = ~new_P2_U2371 | ~P2_REIP_REG_22_;
  assign new_P2_U6077 = ~new_P2_U2370 | ~new_P2_R2278_U100;
  assign new_P2_U6078 = ~P2_PHYADDRPOINTER_REG_22_ | ~new_P2_U5938;
  assign new_P2_U6079 = ~new_P2_R2337_U77 | ~new_P2_U2387;
  assign new_P2_U6080 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U21;
  assign new_P2_U6081 = ~new_P2_U2372 | ~new_P2_R2099_U80;
  assign new_P2_U6082 = ~new_P2_U2371 | ~P2_REIP_REG_23_;
  assign new_P2_U6083 = ~new_P2_U2370 | ~new_P2_R2278_U99;
  assign new_P2_U6084 = ~P2_PHYADDRPOINTER_REG_23_ | ~new_P2_U5938;
  assign new_P2_U6085 = ~new_P2_R2337_U76 | ~new_P2_U2387;
  assign new_P2_U6086 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U70;
  assign new_P2_U6087 = ~new_P2_U2372 | ~new_P2_R2099_U79;
  assign new_P2_U6088 = ~new_P2_U2371 | ~P2_REIP_REG_24_;
  assign new_P2_U6089 = ~new_P2_U2370 | ~new_P2_R2278_U98;
  assign new_P2_U6090 = ~P2_PHYADDRPOINTER_REG_24_ | ~new_P2_U5938;
  assign new_P2_U6091 = ~new_P2_R2337_U75 | ~new_P2_U2387;
  assign new_P2_U6092 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U77;
  assign new_P2_U6093 = ~new_P2_U2372 | ~new_P2_R2099_U78;
  assign new_P2_U6094 = ~new_P2_U2371 | ~P2_REIP_REG_25_;
  assign new_P2_U6095 = ~new_P2_U2370 | ~new_P2_R2278_U97;
  assign new_P2_U6096 = ~P2_PHYADDRPOINTER_REG_25_ | ~new_P2_U5938;
  assign new_P2_U6097 = ~new_P2_R2337_U74 | ~new_P2_U2387;
  assign new_P2_U6098 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U22;
  assign new_P2_U6099 = ~new_P2_U2372 | ~new_P2_R2099_U77;
  assign new_P2_U6100 = ~new_P2_U2371 | ~P2_REIP_REG_26_;
  assign new_P2_U6101 = ~new_P2_U2370 | ~new_P2_R2278_U96;
  assign new_P2_U6102 = ~P2_PHYADDRPOINTER_REG_26_ | ~new_P2_U5938;
  assign new_P2_U6103 = ~new_P2_R2337_U73 | ~new_P2_U2387;
  assign new_P2_U6104 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U74;
  assign new_P2_U6105 = ~new_P2_U2372 | ~new_P2_R2099_U76;
  assign new_P2_U6106 = ~new_P2_U2371 | ~P2_REIP_REG_27_;
  assign new_P2_U6107 = ~new_P2_U2370 | ~new_P2_R2278_U95;
  assign new_P2_U6108 = ~P2_PHYADDRPOINTER_REG_27_ | ~new_P2_U5938;
  assign new_P2_U6109 = ~new_P2_R2337_U72 | ~new_P2_U2387;
  assign new_P2_U6110 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U23;
  assign new_P2_U6111 = ~new_P2_U2372 | ~new_P2_R2099_U75;
  assign new_P2_U6112 = ~new_P2_U2371 | ~P2_REIP_REG_28_;
  assign new_P2_U6113 = ~new_P2_U2370 | ~new_P2_R2278_U94;
  assign new_P2_U6114 = ~P2_PHYADDRPOINTER_REG_28_ | ~new_P2_U5938;
  assign new_P2_U6115 = ~new_P2_R2337_U71 | ~new_P2_U2387;
  assign new_P2_U6116 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U24;
  assign new_P2_U6117 = ~new_P2_U2372 | ~new_P2_R2099_U74;
  assign new_P2_U6118 = ~new_P2_U2371 | ~P2_REIP_REG_29_;
  assign new_P2_U6119 = ~new_P2_U2370 | ~new_P2_R2278_U93;
  assign new_P2_U6120 = ~P2_PHYADDRPOINTER_REG_29_ | ~new_P2_U5938;
  assign new_P2_U6121 = ~new_P2_R2337_U69 | ~new_P2_U2387;
  assign new_P2_U6122 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U69;
  assign new_P2_U6123 = ~new_P2_U2372 | ~new_P2_R2099_U73;
  assign new_P2_U6124 = ~new_P2_U2371 | ~P2_REIP_REG_30_;
  assign new_P2_U6125 = ~new_P2_U2370 | ~new_P2_R2278_U91;
  assign new_P2_U6126 = ~P2_PHYADDRPOINTER_REG_30_ | ~new_P2_U5938;
  assign new_P2_U6127 = ~new_P2_R2337_U68 | ~new_P2_U2387;
  assign new_P2_U6128 = ~new_P2_U2373 | ~new_P2_ADD_371_1212_U83;
  assign new_P2_U6129 = ~new_P2_U2372 | ~new_P2_R2099_U72;
  assign new_P2_U6130 = ~new_P2_U2371 | ~P2_REIP_REG_31_;
  assign new_P2_U6131 = ~new_P2_U2370 | ~new_P2_R2278_U5;
  assign new_P2_U6132 = ~P2_PHYADDRPOINTER_REG_31_ | ~new_P2_U5938;
  assign new_P2_U6133 = ~new_U211 | ~new_P2_U2616;
  assign new_P2_U6134 = ~P2_EAX_REG_15_ | ~new_P2_U2395;
  assign new_P2_U6135 = ~new_U308 | ~new_P2_U2394;
  assign new_P2_U6136 = ~P2_LWORD_REG_15_ | ~new_P2_U3538;
  assign new_P2_U6137 = ~P2_EAX_REG_14_ | ~new_P2_U2395;
  assign new_P2_U6138 = ~new_U309 | ~new_P2_U2394;
  assign new_P2_U6139 = ~P2_LWORD_REG_14_ | ~new_P2_U3538;
  assign new_P2_U6140 = ~P2_EAX_REG_13_ | ~new_P2_U2395;
  assign new_P2_U6141 = ~new_U310 | ~new_P2_U2394;
  assign new_P2_U6142 = ~P2_LWORD_REG_13_ | ~new_P2_U3538;
  assign new_P2_U6143 = ~P2_EAX_REG_12_ | ~new_P2_U2395;
  assign new_P2_U6144 = ~new_U311 | ~new_P2_U2394;
  assign new_P2_U6145 = ~P2_LWORD_REG_12_ | ~new_P2_U3538;
  assign new_P2_U6146 = ~P2_EAX_REG_11_ | ~new_P2_U2395;
  assign new_P2_U6147 = ~new_U312 | ~new_P2_U2394;
  assign new_P2_U6148 = ~P2_LWORD_REG_11_ | ~new_P2_U3538;
  assign new_P2_U6149 = ~P2_EAX_REG_10_ | ~new_P2_U2395;
  assign new_P2_U6150 = ~new_U313 | ~new_P2_U2394;
  assign new_P2_U6151 = ~P2_LWORD_REG_10_ | ~new_P2_U3538;
  assign new_P2_U6152 = ~P2_EAX_REG_9_ | ~new_P2_U2395;
  assign new_P2_U6153 = ~new_U283 | ~new_P2_U2394;
  assign new_P2_U6154 = ~P2_LWORD_REG_9_ | ~new_P2_U3538;
  assign new_P2_U6155 = ~P2_EAX_REG_8_ | ~new_P2_U2395;
  assign new_P2_U6156 = ~new_U284 | ~new_P2_U2394;
  assign new_P2_U6157 = ~P2_LWORD_REG_8_ | ~new_P2_U3538;
  assign new_P2_U6158 = ~P2_EAX_REG_7_ | ~new_P2_U2395;
  assign new_P2_U6159 = ~new_P2_U2394 | ~new_U285;
  assign new_P2_U6160 = ~P2_LWORD_REG_7_ | ~new_P2_U3538;
  assign new_P2_U6161 = ~P2_EAX_REG_6_ | ~new_P2_U2395;
  assign new_P2_U6162 = ~new_P2_U2394 | ~new_U286;
  assign new_P2_U6163 = ~P2_LWORD_REG_6_ | ~new_P2_U3538;
  assign new_P2_U6164 = ~P2_EAX_REG_5_ | ~new_P2_U2395;
  assign new_P2_U6165 = ~new_P2_U2394 | ~new_U287;
  assign new_P2_U6166 = ~P2_LWORD_REG_5_ | ~new_P2_U3538;
  assign new_P2_U6167 = ~P2_EAX_REG_4_ | ~new_P2_U2395;
  assign new_P2_U6168 = ~new_P2_U2394 | ~new_U288;
  assign new_P2_U6169 = ~P2_LWORD_REG_4_ | ~new_P2_U3538;
  assign new_P2_U6170 = ~P2_EAX_REG_3_ | ~new_P2_U2395;
  assign new_P2_U6171 = ~new_P2_U2394 | ~new_U289;
  assign new_P2_U6172 = ~P2_LWORD_REG_3_ | ~new_P2_U3538;
  assign new_P2_U6173 = ~P2_EAX_REG_2_ | ~new_P2_U2395;
  assign new_P2_U6174 = ~new_P2_U2394 | ~new_U292;
  assign new_P2_U6175 = ~P2_LWORD_REG_2_ | ~new_P2_U3538;
  assign new_P2_U6176 = ~P2_EAX_REG_1_ | ~new_P2_U2395;
  assign new_P2_U6177 = ~new_P2_U2394 | ~new_U303;
  assign new_P2_U6178 = ~P2_LWORD_REG_1_ | ~new_P2_U3538;
  assign new_P2_U6179 = ~P2_EAX_REG_0_ | ~new_P2_U2395;
  assign new_P2_U6180 = ~new_P2_U2394 | ~new_U314;
  assign new_P2_U6181 = ~P2_LWORD_REG_0_ | ~new_P2_U3538;
  assign new_P2_U6182 = ~P2_EAX_REG_30_ | ~new_P2_U2395;
  assign new_P2_U6183 = ~new_U309 | ~new_P2_U2394;
  assign new_P2_U6184 = ~P2_UWORD_REG_14_ | ~new_P2_U3538;
  assign new_P2_U6185 = ~P2_EAX_REG_29_ | ~new_P2_U2395;
  assign new_P2_U6186 = ~new_U310 | ~new_P2_U2394;
  assign new_P2_U6187 = ~P2_UWORD_REG_13_ | ~new_P2_U3538;
  assign new_P2_U6188 = ~P2_EAX_REG_28_ | ~new_P2_U2395;
  assign new_P2_U6189 = ~new_U311 | ~new_P2_U2394;
  assign new_P2_U6190 = ~P2_UWORD_REG_12_ | ~new_P2_U3538;
  assign new_P2_U6191 = ~P2_EAX_REG_27_ | ~new_P2_U2395;
  assign new_P2_U6192 = ~new_U312 | ~new_P2_U2394;
  assign new_P2_U6193 = ~P2_UWORD_REG_11_ | ~new_P2_U3538;
  assign new_P2_U6194 = ~P2_EAX_REG_26_ | ~new_P2_U2395;
  assign new_P2_U6195 = ~new_U313 | ~new_P2_U2394;
  assign new_P2_U6196 = ~P2_UWORD_REG_10_ | ~new_P2_U3538;
  assign new_P2_U6197 = ~P2_EAX_REG_25_ | ~new_P2_U2395;
  assign new_P2_U6198 = ~new_U283 | ~new_P2_U2394;
  assign new_P2_U6199 = ~P2_UWORD_REG_9_ | ~new_P2_U3538;
  assign new_P2_U6200 = ~P2_EAX_REG_24_ | ~new_P2_U2395;
  assign new_P2_U6201 = ~new_U284 | ~new_P2_U2394;
  assign new_P2_U6202 = ~P2_UWORD_REG_8_ | ~new_P2_U3538;
  assign new_P2_U6203 = ~P2_EAX_REG_23_ | ~new_P2_U2395;
  assign new_P2_U6204 = ~new_P2_U2394 | ~new_U285;
  assign new_P2_U6205 = ~P2_UWORD_REG_7_ | ~new_P2_U3538;
  assign new_P2_U6206 = ~P2_EAX_REG_22_ | ~new_P2_U2395;
  assign new_P2_U6207 = ~new_P2_U2394 | ~new_U286;
  assign new_P2_U6208 = ~P2_UWORD_REG_6_ | ~new_P2_U3538;
  assign new_P2_U6209 = ~P2_EAX_REG_21_ | ~new_P2_U2395;
  assign new_P2_U6210 = ~new_P2_U2394 | ~new_U287;
  assign new_P2_U6211 = ~P2_UWORD_REG_5_ | ~new_P2_U3538;
  assign new_P2_U6212 = ~P2_EAX_REG_20_ | ~new_P2_U2395;
  assign new_P2_U6213 = ~new_P2_U2394 | ~new_U288;
  assign new_P2_U6214 = ~P2_UWORD_REG_4_ | ~new_P2_U3538;
  assign new_P2_U6215 = ~P2_EAX_REG_19_ | ~new_P2_U2395;
  assign new_P2_U6216 = ~new_P2_U2394 | ~new_U289;
  assign new_P2_U6217 = ~P2_UWORD_REG_3_ | ~new_P2_U3538;
  assign new_P2_U6218 = ~P2_EAX_REG_18_ | ~new_P2_U2395;
  assign new_P2_U6219 = ~new_P2_U2394 | ~new_U292;
  assign new_P2_U6220 = ~P2_UWORD_REG_2_ | ~new_P2_U3538;
  assign new_P2_U6221 = ~P2_EAX_REG_17_ | ~new_P2_U2395;
  assign new_P2_U6222 = ~new_P2_U2394 | ~new_U303;
  assign new_P2_U6223 = ~P2_UWORD_REG_1_ | ~new_P2_U3538;
  assign new_P2_U6224 = ~P2_EAX_REG_16_ | ~new_P2_U2395;
  assign new_P2_U6225 = ~new_P2_U2394 | ~new_U314;
  assign new_P2_U6226 = ~P2_UWORD_REG_0_ | ~new_P2_U3538;
  assign new_P2_U6227 = ~new_P2_R2167_U6 | ~new_P2_U4057 | ~new_P2_U4421;
  assign new_P2_U6228 = ~new_P2_U4058 | ~new_P2_U2446;
  assign new_P2_U6229 = ~new_P2_U6228 | ~new_P2_U6227;
  assign new_P2_U6230 = ~new_P2_U4411 | ~new_P2_U6229;
  assign new_P2_U6231 = ~new_P2_U4467 | ~P2_STATE2_REG_1_;
  assign new_P2_U6232 = ~new_P2_U3541;
  assign new_P2_U6233 = ~new_P2_U2430 | ~P2_EAX_REG_0_;
  assign new_P2_U6234 = ~new_P2_U2396 | ~P2_LWORD_REG_0_;
  assign new_P2_U6235 = ~P2_DATAO_REG_0_ | ~new_P2_U6232;
  assign new_P2_U6236 = ~new_P2_U2430 | ~P2_EAX_REG_1_;
  assign new_P2_U6237 = ~new_P2_U2396 | ~P2_LWORD_REG_1_;
  assign new_P2_U6238 = ~P2_DATAO_REG_1_ | ~new_P2_U6232;
  assign new_P2_U6239 = ~new_P2_U2430 | ~P2_EAX_REG_2_;
  assign new_P2_U6240 = ~new_P2_U2396 | ~P2_LWORD_REG_2_;
  assign new_P2_U6241 = ~P2_DATAO_REG_2_ | ~new_P2_U6232;
  assign new_P2_U6242 = ~new_P2_U2430 | ~P2_EAX_REG_3_;
  assign new_P2_U6243 = ~new_P2_U2396 | ~P2_LWORD_REG_3_;
  assign new_P2_U6244 = ~P2_DATAO_REG_3_ | ~new_P2_U6232;
  assign new_P2_U6245 = ~new_P2_U2430 | ~P2_EAX_REG_4_;
  assign new_P2_U6246 = ~new_P2_U2396 | ~P2_LWORD_REG_4_;
  assign new_P2_U6247 = ~P2_DATAO_REG_4_ | ~new_P2_U6232;
  assign new_P2_U6248 = ~new_P2_U2430 | ~P2_EAX_REG_5_;
  assign new_P2_U6249 = ~new_P2_U2396 | ~P2_LWORD_REG_5_;
  assign new_P2_U6250 = ~P2_DATAO_REG_5_ | ~new_P2_U6232;
  assign new_P2_U6251 = ~new_P2_U2430 | ~P2_EAX_REG_6_;
  assign new_P2_U6252 = ~new_P2_U2396 | ~P2_LWORD_REG_6_;
  assign new_P2_U6253 = ~P2_DATAO_REG_6_ | ~new_P2_U6232;
  assign new_P2_U6254 = ~new_P2_U2430 | ~P2_EAX_REG_7_;
  assign new_P2_U6255 = ~new_P2_U2396 | ~P2_LWORD_REG_7_;
  assign new_P2_U6256 = ~P2_DATAO_REG_7_ | ~new_P2_U6232;
  assign new_P2_U6257 = ~new_P2_U2430 | ~P2_EAX_REG_8_;
  assign new_P2_U6258 = ~new_P2_U2396 | ~P2_LWORD_REG_8_;
  assign new_P2_U6259 = ~P2_DATAO_REG_8_ | ~new_P2_U6232;
  assign new_P2_U6260 = ~new_P2_U2430 | ~P2_EAX_REG_9_;
  assign new_P2_U6261 = ~new_P2_U2396 | ~P2_LWORD_REG_9_;
  assign new_P2_U6262 = ~P2_DATAO_REG_9_ | ~new_P2_U6232;
  assign new_P2_U6263 = ~new_P2_U2430 | ~P2_EAX_REG_10_;
  assign new_P2_U6264 = ~new_P2_U2396 | ~P2_LWORD_REG_10_;
  assign new_P2_U6265 = ~P2_DATAO_REG_10_ | ~new_P2_U6232;
  assign new_P2_U6266 = ~new_P2_U2430 | ~P2_EAX_REG_11_;
  assign new_P2_U6267 = ~new_P2_U2396 | ~P2_LWORD_REG_11_;
  assign new_P2_U6268 = ~P2_DATAO_REG_11_ | ~new_P2_U6232;
  assign new_P2_U6269 = ~new_P2_U2430 | ~P2_EAX_REG_12_;
  assign new_P2_U6270 = ~new_P2_U2396 | ~P2_LWORD_REG_12_;
  assign new_P2_U6271 = ~P2_DATAO_REG_12_ | ~new_P2_U6232;
  assign new_P2_U6272 = ~new_P2_U2430 | ~P2_EAX_REG_13_;
  assign new_P2_U6273 = ~new_P2_U2396 | ~P2_LWORD_REG_13_;
  assign new_P2_U6274 = ~P2_DATAO_REG_13_ | ~new_P2_U6232;
  assign new_P2_U6275 = ~new_P2_U2430 | ~P2_EAX_REG_14_;
  assign new_P2_U6276 = ~new_P2_U2396 | ~P2_LWORD_REG_14_;
  assign new_P2_U6277 = ~P2_DATAO_REG_14_ | ~new_P2_U6232;
  assign new_P2_U6278 = ~new_P2_U2430 | ~P2_EAX_REG_15_;
  assign new_P2_U6279 = ~new_P2_U2396 | ~P2_LWORD_REG_15_;
  assign new_P2_U6280 = ~P2_DATAO_REG_15_ | ~new_P2_U6232;
  assign new_P2_U6281 = ~new_P2_U2435 | ~P2_EAX_REG_16_;
  assign new_P2_U6282 = ~new_P2_U2396 | ~P2_UWORD_REG_0_;
  assign new_P2_U6283 = ~P2_DATAO_REG_16_ | ~new_P2_U6232;
  assign new_P2_U6284 = ~new_P2_U2435 | ~P2_EAX_REG_17_;
  assign new_P2_U6285 = ~new_P2_U2396 | ~P2_UWORD_REG_1_;
  assign new_P2_U6286 = ~P2_DATAO_REG_17_ | ~new_P2_U6232;
  assign new_P2_U6287 = ~new_P2_U2435 | ~P2_EAX_REG_18_;
  assign new_P2_U6288 = ~new_P2_U2396 | ~P2_UWORD_REG_2_;
  assign new_P2_U6289 = ~P2_DATAO_REG_18_ | ~new_P2_U6232;
  assign new_P2_U6290 = ~new_P2_U2435 | ~P2_EAX_REG_19_;
  assign new_P2_U6291 = ~new_P2_U2396 | ~P2_UWORD_REG_3_;
  assign new_P2_U6292 = ~P2_DATAO_REG_19_ | ~new_P2_U6232;
  assign new_P2_U6293 = ~new_P2_U2435 | ~P2_EAX_REG_20_;
  assign new_P2_U6294 = ~new_P2_U2396 | ~P2_UWORD_REG_4_;
  assign new_P2_U6295 = ~P2_DATAO_REG_20_ | ~new_P2_U6232;
  assign new_P2_U6296 = ~new_P2_U2435 | ~P2_EAX_REG_21_;
  assign new_P2_U6297 = ~new_P2_U2396 | ~P2_UWORD_REG_5_;
  assign new_P2_U6298 = ~P2_DATAO_REG_21_ | ~new_P2_U6232;
  assign new_P2_U6299 = ~new_P2_U2435 | ~P2_EAX_REG_22_;
  assign new_P2_U6300 = ~new_P2_U2396 | ~P2_UWORD_REG_6_;
  assign new_P2_U6301 = ~P2_DATAO_REG_22_ | ~new_P2_U6232;
  assign new_P2_U6302 = ~new_P2_U2435 | ~P2_EAX_REG_23_;
  assign new_P2_U6303 = ~new_P2_U2396 | ~P2_UWORD_REG_7_;
  assign new_P2_U6304 = ~P2_DATAO_REG_23_ | ~new_P2_U6232;
  assign new_P2_U6305 = ~new_P2_U2435 | ~P2_EAX_REG_24_;
  assign new_P2_U6306 = ~new_P2_U2396 | ~P2_UWORD_REG_8_;
  assign new_P2_U6307 = ~P2_DATAO_REG_24_ | ~new_P2_U6232;
  assign new_P2_U6308 = ~new_P2_U2435 | ~P2_EAX_REG_25_;
  assign new_P2_U6309 = ~new_P2_U2396 | ~P2_UWORD_REG_9_;
  assign new_P2_U6310 = ~P2_DATAO_REG_25_ | ~new_P2_U6232;
  assign new_P2_U6311 = ~new_P2_U2435 | ~P2_EAX_REG_26_;
  assign new_P2_U6312 = ~new_P2_U2396 | ~P2_UWORD_REG_10_;
  assign new_P2_U6313 = ~P2_DATAO_REG_26_ | ~new_P2_U6232;
  assign new_P2_U6314 = ~new_P2_U2435 | ~P2_EAX_REG_27_;
  assign new_P2_U6315 = ~new_P2_U2396 | ~P2_UWORD_REG_11_;
  assign new_P2_U6316 = ~P2_DATAO_REG_27_ | ~new_P2_U6232;
  assign new_P2_U6317 = ~new_P2_U2435 | ~P2_EAX_REG_28_;
  assign new_P2_U6318 = ~new_P2_U2396 | ~P2_UWORD_REG_12_;
  assign new_P2_U6319 = ~P2_DATAO_REG_28_ | ~new_P2_U6232;
  assign new_P2_U6320 = ~new_P2_U2435 | ~P2_EAX_REG_29_;
  assign new_P2_U6321 = ~new_P2_U2396 | ~P2_UWORD_REG_13_;
  assign new_P2_U6322 = ~P2_DATAO_REG_29_ | ~new_P2_U6232;
  assign new_P2_U6323 = ~new_P2_U2435 | ~P2_EAX_REG_30_;
  assign new_P2_U6324 = ~new_P2_U2396 | ~P2_UWORD_REG_14_;
  assign new_P2_U6325 = ~P2_DATAO_REG_30_ | ~new_P2_U6232;
  assign new_P2_U6326 = ~new_P2_U2513 | ~new_P2_U3254;
  assign new_P2_U6327 = ~new_P2_U2433 | ~new_U314;
  assign new_P2_U6328 = ~new_P2_ADD_391_1196_U87 | ~new_P2_U2397;
  assign new_P2_U6329 = ~new_P2_U2380 | ~new_P2_R2096_U68;
  assign new_P2_U6330 = ~P2_EAX_REG_0_ | ~new_P2_U3542;
  assign new_P2_U6331 = ~new_P2_U2433 | ~new_U303;
  assign new_P2_U6332 = ~new_P2_ADD_391_1196_U12 | ~new_P2_U2397;
  assign new_P2_U6333 = ~new_P2_U2380 | ~new_P2_R2096_U51;
  assign new_P2_U6334 = ~P2_EAX_REG_1_ | ~new_P2_U3542;
  assign new_P2_U6335 = ~new_P2_U2433 | ~new_U292;
  assign new_P2_U6336 = ~new_P2_ADD_391_1196_U92 | ~new_P2_U2397;
  assign new_P2_U6337 = ~new_P2_U2380 | ~new_P2_R2096_U77;
  assign new_P2_U6338 = ~P2_EAX_REG_2_ | ~new_P2_U3542;
  assign new_P2_U6339 = ~new_P2_U2433 | ~new_U289;
  assign new_P2_U6340 = ~new_P2_ADD_391_1196_U91 | ~new_P2_U2397;
  assign new_P2_U6341 = ~new_P2_U2380 | ~new_P2_R2096_U75;
  assign new_P2_U6342 = ~P2_EAX_REG_3_ | ~new_P2_U3542;
  assign new_P2_U6343 = ~new_P2_U2433 | ~new_U288;
  assign new_P2_U6344 = ~new_P2_ADD_391_1196_U90 | ~new_P2_U2397;
  assign new_P2_U6345 = ~new_P2_U2380 | ~new_P2_R2096_U74;
  assign new_P2_U6346 = ~P2_EAX_REG_4_ | ~new_P2_U3542;
  assign new_P2_U6347 = ~new_P2_U2433 | ~new_U287;
  assign new_P2_U6348 = ~new_P2_ADD_391_1196_U9 | ~new_P2_U2397;
  assign new_P2_U6349 = ~new_P2_U2380 | ~new_P2_R2096_U73;
  assign new_P2_U6350 = ~P2_EAX_REG_5_ | ~new_P2_U3542;
  assign new_P2_U6351 = ~new_P2_U2433 | ~new_U286;
  assign new_P2_U6352 = ~new_P2_ADD_391_1196_U89 | ~new_P2_U2397;
  assign new_P2_U6353 = ~new_P2_U2380 | ~new_P2_R2096_U72;
  assign new_P2_U6354 = ~P2_EAX_REG_6_ | ~new_P2_U3542;
  assign new_P2_U6355 = ~new_P2_U2433 | ~new_U285;
  assign new_P2_U6356 = ~new_P2_ADD_391_1196_U10 | ~new_P2_U2397;
  assign new_P2_U6357 = ~new_P2_U2380 | ~new_P2_R2096_U71;
  assign new_P2_U6358 = ~P2_EAX_REG_7_ | ~new_P2_U3542;
  assign new_P2_U6359 = ~new_P2_U2433 | ~new_U284;
  assign new_P2_U6360 = ~new_P2_ADD_391_1196_U88 | ~new_P2_U2397;
  assign new_P2_U6361 = ~new_P2_U2380 | ~new_P2_R2096_U70;
  assign new_P2_U6362 = ~P2_EAX_REG_8_ | ~new_P2_U3542;
  assign new_P2_U6363 = ~new_P2_U2433 | ~new_U283;
  assign new_P2_U6364 = ~new_P2_ADD_391_1196_U11 | ~new_P2_U2397;
  assign new_P2_U6365 = ~new_P2_U2380 | ~new_P2_R2096_U69;
  assign new_P2_U6366 = ~P2_EAX_REG_9_ | ~new_P2_U3542;
  assign new_P2_U6367 = ~new_P2_U2433 | ~new_U313;
  assign new_P2_U6368 = ~new_P2_ADD_391_1196_U109 | ~new_P2_U2397;
  assign new_P2_U6369 = ~new_P2_U2380 | ~new_P2_R2096_U97;
  assign new_P2_U6370 = ~P2_EAX_REG_10_ | ~new_P2_U3542;
  assign new_P2_U6371 = ~new_P2_U2433 | ~new_U312;
  assign new_P2_U6372 = ~new_P2_ADD_391_1196_U5 | ~new_P2_U2397;
  assign new_P2_U6373 = ~new_P2_U2380 | ~new_P2_R2096_U96;
  assign new_P2_U6374 = ~P2_EAX_REG_11_ | ~new_P2_U3542;
  assign new_P2_U6375 = ~new_P2_U2433 | ~new_U311;
  assign new_P2_U6376 = ~new_P2_ADD_391_1196_U108 | ~new_P2_U2397;
  assign new_P2_U6377 = ~new_P2_U2380 | ~new_P2_R2096_U95;
  assign new_P2_U6378 = ~P2_EAX_REG_12_ | ~new_P2_U3542;
  assign new_P2_U6379 = ~new_P2_U2433 | ~new_U310;
  assign new_P2_U6380 = ~new_P2_ADD_391_1196_U6 | ~new_P2_U2397;
  assign new_P2_U6381 = ~new_P2_U2380 | ~new_P2_R2096_U94;
  assign new_P2_U6382 = ~P2_EAX_REG_13_ | ~new_P2_U3542;
  assign new_P2_U6383 = ~new_P2_U2433 | ~new_U309;
  assign new_P2_U6384 = ~new_P2_ADD_391_1196_U107 | ~new_P2_U2397;
  assign new_P2_U6385 = ~new_P2_U2380 | ~new_P2_R2096_U93;
  assign new_P2_U6386 = ~P2_EAX_REG_14_ | ~new_P2_U3542;
  assign new_P2_U6387 = ~new_P2_U2433 | ~new_U308;
  assign new_P2_U6388 = ~new_P2_ADD_391_1196_U7 | ~new_P2_U2397;
  assign new_P2_U6389 = ~new_P2_U2380 | ~new_P2_R2096_U92;
  assign new_P2_U6390 = ~P2_EAX_REG_15_ | ~new_P2_U3542;
  assign new_P2_U6391 = ~new_P2_U2434 | ~new_U314;
  assign new_P2_U6392 = ~new_P2_U2427 | ~new_U307;
  assign new_P2_U6393 = ~new_P2_ADD_391_1196_U106 | ~new_P2_U2397;
  assign new_P2_U6394 = ~new_P2_U2380 | ~new_P2_R2096_U91;
  assign new_P2_U6395 = ~P2_EAX_REG_16_ | ~new_P2_U3542;
  assign new_P2_U6396 = ~new_P2_U2434 | ~new_U303;
  assign new_P2_U6397 = ~new_P2_U2427 | ~new_U306;
  assign new_P2_U6398 = ~new_P2_ADD_391_1196_U105 | ~new_P2_U2397;
  assign new_P2_U6399 = ~new_P2_U2380 | ~new_P2_R2096_U90;
  assign new_P2_U6400 = ~P2_EAX_REG_17_ | ~new_P2_U3542;
  assign new_P2_U6401 = ~new_P2_U2434 | ~new_U292;
  assign new_P2_U6402 = ~new_P2_U2427 | ~new_U305;
  assign new_P2_U6403 = ~new_P2_ADD_391_1196_U104 | ~new_P2_U2397;
  assign new_P2_U6404 = ~new_P2_U2380 | ~new_P2_R2096_U89;
  assign new_P2_U6405 = ~P2_EAX_REG_18_ | ~new_P2_U3542;
  assign new_P2_U6406 = ~new_P2_U2434 | ~new_U289;
  assign new_P2_U6407 = ~new_P2_U2427 | ~new_U304;
  assign new_P2_U6408 = ~new_P2_ADD_391_1196_U103 | ~new_P2_U2397;
  assign new_P2_U6409 = ~new_P2_U2380 | ~new_P2_R2096_U88;
  assign new_P2_U6410 = ~P2_EAX_REG_19_ | ~new_P2_U3542;
  assign new_P2_U6411 = ~new_P2_U2434 | ~new_U288;
  assign new_P2_U6412 = ~new_P2_U2427 | ~new_U302;
  assign new_P2_U6413 = ~new_P2_ADD_391_1196_U102 | ~new_P2_U2397;
  assign new_P2_U6414 = ~new_P2_U2380 | ~new_P2_R2096_U87;
  assign new_P2_U6415 = ~P2_EAX_REG_20_ | ~new_P2_U3542;
  assign new_P2_U6416 = ~new_P2_U2434 | ~new_U287;
  assign new_P2_U6417 = ~new_P2_U2427 | ~new_U301;
  assign new_P2_U6418 = ~new_P2_ADD_391_1196_U101 | ~new_P2_U2397;
  assign new_P2_U6419 = ~new_P2_U2380 | ~new_P2_R2096_U86;
  assign new_P2_U6420 = ~P2_EAX_REG_21_ | ~new_P2_U3542;
  assign new_P2_U6421 = ~new_P2_U2434 | ~new_U286;
  assign new_P2_U6422 = ~new_P2_U2427 | ~new_U300;
  assign new_P2_U6423 = ~new_P2_ADD_391_1196_U100 | ~new_P2_U2397;
  assign new_P2_U6424 = ~new_P2_U2380 | ~new_P2_R2096_U85;
  assign new_P2_U6425 = ~P2_EAX_REG_22_ | ~new_P2_U3542;
  assign new_P2_U6426 = ~new_P2_U2434 | ~new_U285;
  assign new_P2_U6427 = ~new_P2_U2427 | ~new_U299;
  assign new_P2_U6428 = ~new_P2_ADD_391_1196_U99 | ~new_P2_U2397;
  assign new_P2_U6429 = ~new_P2_U2380 | ~new_P2_R2096_U84;
  assign new_P2_U6430 = ~P2_EAX_REG_23_ | ~new_P2_U3542;
  assign new_P2_U6431 = ~new_P2_U2434 | ~new_U284;
  assign new_P2_U6432 = ~new_P2_U2427 | ~new_U298;
  assign new_P2_U6433 = ~new_P2_ADD_391_1196_U98 | ~new_P2_U2397;
  assign new_P2_U6434 = ~new_P2_U2380 | ~new_P2_R2096_U83;
  assign new_P2_U6435 = ~P2_EAX_REG_24_ | ~new_P2_U3542;
  assign new_P2_U6436 = ~new_P2_U2434 | ~new_U283;
  assign new_P2_U6437 = ~new_P2_U2427 | ~new_U297;
  assign new_P2_U6438 = ~new_P2_ADD_391_1196_U97 | ~new_P2_U2397;
  assign new_P2_U6439 = ~new_P2_U2380 | ~new_P2_R2096_U82;
  assign new_P2_U6440 = ~P2_EAX_REG_25_ | ~new_P2_U3542;
  assign new_P2_U6441 = ~new_P2_U2434 | ~new_U313;
  assign new_P2_U6442 = ~new_P2_U2427 | ~new_U296;
  assign new_P2_U6443 = ~new_P2_ADD_391_1196_U96 | ~new_P2_U2397;
  assign new_P2_U6444 = ~new_P2_U2380 | ~new_P2_R2096_U81;
  assign new_P2_U6445 = ~P2_EAX_REG_26_ | ~new_P2_U3542;
  assign new_P2_U6446 = ~new_P2_U2434 | ~new_U312;
  assign new_P2_U6447 = ~new_P2_U2427 | ~new_U295;
  assign new_P2_U6448 = ~new_P2_ADD_391_1196_U95 | ~new_P2_U2397;
  assign new_P2_U6449 = ~new_P2_U2380 | ~new_P2_R2096_U80;
  assign new_P2_U6450 = ~P2_EAX_REG_27_ | ~new_P2_U3542;
  assign new_P2_U6451 = ~new_P2_U2434 | ~new_U311;
  assign new_P2_U6452 = ~new_P2_U2427 | ~new_U294;
  assign new_P2_U6453 = ~new_P2_ADD_391_1196_U94 | ~new_P2_U2397;
  assign new_P2_U6454 = ~new_P2_U2380 | ~new_P2_R2096_U79;
  assign new_P2_U6455 = ~P2_EAX_REG_28_ | ~new_P2_U3542;
  assign new_P2_U6456 = ~new_P2_U2434 | ~new_U310;
  assign new_P2_U6457 = ~new_P2_U2427 | ~new_U293;
  assign new_P2_U6458 = ~new_P2_ADD_391_1196_U93 | ~new_P2_U2397;
  assign new_P2_U6459 = ~new_P2_U2380 | ~new_P2_R2096_U78;
  assign new_P2_U6460 = ~P2_EAX_REG_29_ | ~new_P2_U3542;
  assign new_P2_U6461 = ~new_P2_U2434 | ~new_U309;
  assign new_P2_U6462 = ~new_P2_U2427 | ~new_U291;
  assign new_P2_U6463 = ~new_P2_ADD_391_1196_U8 | ~new_P2_U2397;
  assign new_P2_U6464 = ~new_P2_U2380 | ~new_P2_R2096_U76;
  assign new_P2_U6465 = ~P2_EAX_REG_30_ | ~new_P2_U3542;
  assign new_P2_U6466 = ~new_P2_U2427 | ~new_U290;
  assign new_P2_U6467 = ~new_P2_U2380 | ~new_P2_R2096_U50;
  assign new_P2_U6468 = ~P2_EAX_REG_31_ | ~new_P2_U3542;
  assign new_P2_U6469 = ~new_P2_U4435 | ~new_P2_U3297;
  assign new_P2_U6470 = ~new_P2_U3578 | ~new_P2_U6469;
  assign new_P2_U6471 = ~new_P2_U2393 | ~new_P2_R2182_U69;
  assign new_P2_U6472 = ~new_P2_U2379 | ~new_P2_R2099_U94;
  assign new_P2_U6473 = ~P2_EBX_REG_0_ | ~new_P2_U3543;
  assign new_P2_U6474 = ~new_P2_U2393 | ~new_P2_R2182_U68;
  assign new_P2_U6475 = ~new_P2_U2379 | ~new_P2_R2099_U5;
  assign new_P2_U6476 = ~P2_EBX_REG_1_ | ~new_P2_U3543;
  assign new_P2_U6477 = ~new_P2_U2393 | ~new_P2_R2182_U40;
  assign new_P2_U6478 = ~new_P2_U2379 | ~new_P2_R2099_U96;
  assign new_P2_U6479 = ~P2_EBX_REG_2_ | ~new_P2_U3543;
  assign new_P2_U6480 = ~new_P2_U2393 | ~new_P2_R2182_U76;
  assign new_P2_U6481 = ~new_P2_U2379 | ~new_P2_R2099_U95;
  assign new_P2_U6482 = ~P2_EBX_REG_3_ | ~new_P2_U3543;
  assign new_P2_U6483 = ~new_P2_R2182_U75 | ~new_P2_U2393;
  assign new_P2_U6484 = ~new_P2_U2379 | ~new_P2_R2099_U98;
  assign new_P2_U6485 = ~P2_EBX_REG_4_ | ~new_P2_U3543;
  assign new_P2_U6486 = ~new_P2_R2182_U74 | ~new_P2_U2393;
  assign new_P2_U6487 = ~new_P2_U2379 | ~new_P2_R2099_U71;
  assign new_P2_U6488 = ~P2_EBX_REG_5_ | ~new_P2_U3543;
  assign new_P2_U6489 = ~new_P2_R2182_U73 | ~new_P2_U2393;
  assign new_P2_U6490 = ~new_P2_U2379 | ~new_P2_R2099_U70;
  assign new_P2_U6491 = ~P2_EBX_REG_6_ | ~new_P2_U3543;
  assign new_P2_U6492 = ~new_P2_R2182_U72 | ~new_P2_U2393;
  assign new_P2_U6493 = ~new_P2_U2379 | ~new_P2_R2099_U69;
  assign new_P2_U6494 = ~P2_EBX_REG_7_ | ~new_P2_U3543;
  assign new_P2_U6495 = ~new_P2_R2182_U71 | ~new_P2_U2393;
  assign new_P2_U6496 = ~new_P2_U2379 | ~new_P2_R2099_U68;
  assign new_P2_U6497 = ~P2_EBX_REG_8_ | ~new_P2_U3543;
  assign new_P2_U6498 = ~new_P2_R2182_U70 | ~new_P2_U2393;
  assign new_P2_U6499 = ~new_P2_U2379 | ~new_P2_R2099_U67;
  assign new_P2_U6500 = ~P2_EBX_REG_9_ | ~new_P2_U3543;
  assign new_P2_U6501 = ~new_P2_R2182_U96 | ~new_P2_U2393;
  assign new_P2_U6502 = ~new_P2_U2379 | ~new_P2_R2099_U93;
  assign new_P2_U6503 = ~P2_EBX_REG_10_ | ~new_P2_U3543;
  assign new_P2_U6504 = ~new_P2_R2182_U95 | ~new_P2_U2393;
  assign new_P2_U6505 = ~new_P2_U2379 | ~new_P2_R2099_U92;
  assign new_P2_U6506 = ~P2_EBX_REG_11_ | ~new_P2_U3543;
  assign new_P2_U6507 = ~new_P2_R2182_U94 | ~new_P2_U2393;
  assign new_P2_U6508 = ~new_P2_U2379 | ~new_P2_R2099_U91;
  assign new_P2_U6509 = ~P2_EBX_REG_12_ | ~new_P2_U3543;
  assign new_P2_U6510 = ~new_P2_R2182_U93 | ~new_P2_U2393;
  assign new_P2_U6511 = ~new_P2_U2379 | ~new_P2_R2099_U90;
  assign new_P2_U6512 = ~P2_EBX_REG_13_ | ~new_P2_U3543;
  assign new_P2_U6513 = ~new_P2_R2182_U92 | ~new_P2_U2393;
  assign new_P2_U6514 = ~new_P2_U2379 | ~new_P2_R2099_U89;
  assign new_P2_U6515 = ~P2_EBX_REG_14_ | ~new_P2_U3543;
  assign new_P2_U6516 = ~new_P2_R2182_U91 | ~new_P2_U2393;
  assign new_P2_U6517 = ~new_P2_U2379 | ~new_P2_R2099_U88;
  assign new_P2_U6518 = ~P2_EBX_REG_15_ | ~new_P2_U3543;
  assign new_P2_U6519 = ~new_P2_R2182_U90 | ~new_P2_U2393;
  assign new_P2_U6520 = ~new_P2_U2379 | ~new_P2_R2099_U87;
  assign new_P2_U6521 = ~P2_EBX_REG_16_ | ~new_P2_U3543;
  assign new_P2_U6522 = ~new_P2_R2182_U89 | ~new_P2_U2393;
  assign new_P2_U6523 = ~new_P2_U2379 | ~new_P2_R2099_U86;
  assign new_P2_U6524 = ~P2_EBX_REG_17_ | ~new_P2_U3543;
  assign new_P2_U6525 = ~new_P2_R2182_U88 | ~new_P2_U2393;
  assign new_P2_U6526 = ~new_P2_U2379 | ~new_P2_R2099_U85;
  assign new_P2_U6527 = ~P2_EBX_REG_18_ | ~new_P2_U3543;
  assign new_P2_U6528 = ~new_P2_R2182_U87 | ~new_P2_U2393;
  assign new_P2_U6529 = ~new_P2_U2379 | ~new_P2_R2099_U84;
  assign new_P2_U6530 = ~P2_EBX_REG_19_ | ~new_P2_U3543;
  assign new_P2_U6531 = ~new_P2_R2182_U86 | ~new_P2_U2393;
  assign new_P2_U6532 = ~new_P2_U2379 | ~new_P2_R2099_U83;
  assign new_P2_U6533 = ~P2_EBX_REG_20_ | ~new_P2_U3543;
  assign new_P2_U6534 = ~new_P2_R2182_U85 | ~new_P2_U2393;
  assign new_P2_U6535 = ~new_P2_U2379 | ~new_P2_R2099_U82;
  assign new_P2_U6536 = ~P2_EBX_REG_21_ | ~new_P2_U3543;
  assign new_P2_U6537 = ~new_P2_R2182_U84 | ~new_P2_U2393;
  assign new_P2_U6538 = ~new_P2_U2379 | ~new_P2_R2099_U81;
  assign new_P2_U6539 = ~P2_EBX_REG_22_ | ~new_P2_U3543;
  assign new_P2_U6540 = ~new_P2_R2182_U83 | ~new_P2_U2393;
  assign new_P2_U6541 = ~new_P2_U2379 | ~new_P2_R2099_U80;
  assign new_P2_U6542 = ~P2_EBX_REG_23_ | ~new_P2_U3543;
  assign new_P2_U6543 = ~new_P2_R2182_U82 | ~new_P2_U2393;
  assign new_P2_U6544 = ~new_P2_U2379 | ~new_P2_R2099_U79;
  assign new_P2_U6545 = ~P2_EBX_REG_24_ | ~new_P2_U3543;
  assign new_P2_U6546 = ~new_P2_R2182_U81 | ~new_P2_U2393;
  assign new_P2_U6547 = ~new_P2_U2379 | ~new_P2_R2099_U78;
  assign new_P2_U6548 = ~P2_EBX_REG_25_ | ~new_P2_U3543;
  assign new_P2_U6549 = ~new_P2_R2182_U80 | ~new_P2_U2393;
  assign new_P2_U6550 = ~new_P2_U2379 | ~new_P2_R2099_U77;
  assign new_P2_U6551 = ~P2_EBX_REG_26_ | ~new_P2_U3543;
  assign new_P2_U6552 = ~new_P2_R2182_U79 | ~new_P2_U2393;
  assign new_P2_U6553 = ~new_P2_U2379 | ~new_P2_R2099_U76;
  assign new_P2_U6554 = ~P2_EBX_REG_27_ | ~new_P2_U3543;
  assign new_P2_U6555 = ~new_P2_R2182_U78 | ~new_P2_U2393;
  assign new_P2_U6556 = ~new_P2_U2379 | ~new_P2_R2099_U75;
  assign new_P2_U6557 = ~P2_EBX_REG_28_ | ~new_P2_U3543;
  assign new_P2_U6558 = ~new_P2_R2182_U77 | ~new_P2_U2393;
  assign new_P2_U6559 = ~new_P2_U2379 | ~new_P2_R2099_U74;
  assign new_P2_U6560 = ~P2_EBX_REG_29_ | ~new_P2_U3543;
  assign new_P2_U6561 = ~new_P2_R2182_U41 | ~new_P2_U2393;
  assign new_P2_U6562 = ~new_P2_U2379 | ~new_P2_R2099_U73;
  assign new_P2_U6563 = ~P2_EBX_REG_30_ | ~new_P2_U3543;
  assign new_P2_U6564 = ~new_P2_U2379 | ~new_P2_R2099_U72;
  assign new_P2_U6565 = ~P2_EBX_REG_31_ | ~new_P2_U3543;
  assign new_P2_U6566 = ~new_P2_R2088_U6 | ~new_P2_U4603;
  assign new_P2_U6567 = ~new_P2_U4433 | ~new_P2_R2167_U6;
  assign new_P2_U6568 = ~new_P2_U6567 | ~new_P2_U6566;
  assign new_P2_U6569 = ~new_P2_U4461 | ~new_P2_U3284;
  assign new_P2_U6570 = ~new_P2_U3546;
  assign new_P2_U6571 = ~new_P2_U3545;
  assign new_P2_U6572 = P2_STATEBS16_REG | new_U211;
  assign new_P2_U6573 = ~new_P2_R2267_U21 | ~new_P2_U2587;
  assign new_P2_U6574 = ~new_P2_U2588 | ~new_P2_R2096_U68;
  assign new_P2_U6575 = ~P2_EBX_REG_0_ | ~new_P2_U7743;
  assign new_P2_U6576 = ~new_P2_U2437 | ~new_P2_R2182_U69;
  assign new_P2_U6577 = ~new_P2_U2392 | ~new_P2_R2099_U94;
  assign new_P2_U6578 = ~new_P2_U2383 | ~P2_PHYADDRPOINTER_REG_0_;
  assign new_P2_U6579 = ~new_P2_U2382 | ~new_P2_U3683;
  assign new_P2_U6580 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_0_;
  assign new_P2_U6581 = ~new_P2_U6570 | ~P2_REIP_REG_0_;
  assign new_P2_U6582 = ~new_P2_R2267_U43 | ~new_P2_U2587;
  assign new_P2_U6583 = ~new_P2_U2588 | ~new_P2_R2096_U51;
  assign new_P2_U6584 = ~P2_EBX_REG_1_ | ~new_P2_U7743;
  assign new_P2_U6585 = ~new_P2_U2437 | ~new_P2_R2182_U68;
  assign new_P2_U6586 = ~new_P2_U2392 | ~new_P2_R2099_U5;
  assign new_P2_U6587 = ~new_P2_U2383 | ~new_P2_R2337_U4;
  assign new_P2_U6588 = ~new_P2_U2382 | ~new_P2_R1957_U49;
  assign new_P2_U6589 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_1_;
  assign new_P2_U6590 = ~new_P2_U6570 | ~P2_REIP_REG_1_;
  assign new_P2_U6591 = ~new_P2_R2267_U65 | ~new_P2_U2587;
  assign new_P2_U6592 = ~new_P2_U2588 | ~new_P2_R2096_U77;
  assign new_P2_U6593 = ~P2_EBX_REG_2_ | ~new_P2_U7743;
  assign new_P2_U6594 = ~new_P2_U2437 | ~new_P2_R2182_U40;
  assign new_P2_U6595 = ~new_P2_U2392 | ~new_P2_R2099_U96;
  assign new_P2_U6596 = ~new_P2_U2383 | ~new_P2_R2337_U70;
  assign new_P2_U6597 = ~new_P2_R1957_U17 | ~new_P2_U2382;
  assign new_P2_U6598 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_2_;
  assign new_P2_U6599 = ~new_P2_U6570 | ~P2_REIP_REG_2_;
  assign new_P2_U6600 = ~new_P2_R2267_U17 | ~new_P2_U2587;
  assign new_P2_U6601 = ~new_P2_U2588 | ~new_P2_R2096_U75;
  assign new_P2_U6602 = ~P2_EBX_REG_3_ | ~new_P2_U7743;
  assign new_P2_U6603 = ~new_P2_U2437 | ~new_P2_R2182_U76;
  assign new_P2_U6604 = ~new_P2_U2392 | ~new_P2_R2099_U95;
  assign new_P2_U6605 = ~new_P2_U2383 | ~new_P2_R2337_U67;
  assign new_P2_U6606 = ~new_P2_R1957_U59 | ~new_P2_U2382;
  assign new_P2_U6607 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_3_;
  assign new_P2_U6608 = ~new_P2_U6570 | ~P2_REIP_REG_3_;
  assign new_P2_U6609 = ~new_P2_R2267_U60 | ~new_P2_U2587;
  assign new_P2_U6610 = ~new_P2_U2588 | ~new_P2_R2096_U74;
  assign new_P2_U6611 = ~P2_EBX_REG_4_ | ~new_P2_U7743;
  assign new_P2_U6612 = ~new_P2_U2437 | ~new_P2_R2182_U75;
  assign new_P2_U6613 = ~new_P2_U2392 | ~new_P2_R2099_U98;
  assign new_P2_U6614 = ~new_P2_U2383 | ~new_P2_R2337_U66;
  assign new_P2_U6615 = ~new_P2_R1957_U18 | ~new_P2_U2382;
  assign new_P2_U6616 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_4_;
  assign new_P2_U6617 = ~new_P2_U6570 | ~P2_REIP_REG_4_;
  assign new_P2_U6618 = ~new_P2_R2267_U18 | ~new_P2_U2587;
  assign new_P2_U6619 = ~new_P2_U2588 | ~new_P2_R2096_U73;
  assign new_P2_U6620 = ~P2_EBX_REG_5_ | ~new_P2_U7743;
  assign new_P2_U6621 = ~new_P2_U2437 | ~new_P2_R2182_U74;
  assign new_P2_U6622 = ~new_P2_U2392 | ~new_P2_R2099_U71;
  assign new_P2_U6623 = ~new_P2_U2383 | ~new_P2_R2337_U65;
  assign new_P2_U6624 = ~new_P2_R1957_U57 | ~new_P2_U2382;
  assign new_P2_U6625 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_5_;
  assign new_P2_U6626 = ~new_P2_U6570 | ~P2_REIP_REG_5_;
  assign new_P2_U6627 = ~new_P2_R2267_U58 | ~new_P2_U2587;
  assign new_P2_U6628 = ~new_P2_U2588 | ~new_P2_R2096_U72;
  assign new_P2_U6629 = ~P2_EBX_REG_6_ | ~new_P2_U7743;
  assign new_P2_U6630 = ~new_P2_U2392 | ~new_P2_R2099_U70;
  assign new_P2_U6631 = ~new_P2_U2383 | ~new_P2_R2337_U64;
  assign new_P2_U6632 = ~new_P2_R1957_U19 | ~new_P2_U2382;
  assign new_P2_U6633 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_6_;
  assign new_P2_U6634 = ~new_P2_U6570 | ~P2_REIP_REG_6_;
  assign new_P2_U6635 = ~new_P2_R2267_U19 | ~new_P2_U2587;
  assign new_P2_U6636 = ~new_P2_U2588 | ~new_P2_R2096_U71;
  assign new_P2_U6637 = ~P2_EBX_REG_7_ | ~new_P2_U7743;
  assign new_P2_U6638 = ~new_P2_U2392 | ~new_P2_R2099_U69;
  assign new_P2_U6639 = ~new_P2_U2383 | ~new_P2_R2337_U63;
  assign new_P2_U6640 = ~new_P2_R1957_U55 | ~new_P2_U2382;
  assign new_P2_U6641 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_7_;
  assign new_P2_U6642 = ~new_P2_U6570 | ~P2_REIP_REG_7_;
  assign new_P2_U6643 = ~new_P2_R2267_U56 | ~new_P2_U2587;
  assign new_P2_U6644 = ~new_P2_U2588 | ~new_P2_R2096_U70;
  assign new_P2_U6645 = ~P2_EBX_REG_8_ | ~new_P2_U7743;
  assign new_P2_U6646 = ~new_P2_U2392 | ~new_P2_R2099_U68;
  assign new_P2_U6647 = ~new_P2_U2383 | ~new_P2_R2337_U62;
  assign new_P2_U6648 = ~new_P2_R1957_U20 | ~new_P2_U2382;
  assign new_P2_U6649 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_8_;
  assign new_P2_U6650 = ~new_P2_U6570 | ~P2_REIP_REG_8_;
  assign new_P2_U6651 = ~new_P2_R2267_U20 | ~new_P2_U2587;
  assign new_P2_U6652 = ~new_P2_U2588 | ~new_P2_R2096_U69;
  assign new_P2_U6653 = ~P2_EBX_REG_9_ | ~new_P2_U7743;
  assign new_P2_U6654 = ~new_P2_U2392 | ~new_P2_R2099_U67;
  assign new_P2_U6655 = ~new_P2_U2383 | ~new_P2_R2337_U61;
  assign new_P2_U6656 = ~new_P2_R1957_U53 | ~new_P2_U2382;
  assign new_P2_U6657 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_9_;
  assign new_P2_U6658 = ~new_P2_U6570 | ~P2_REIP_REG_9_;
  assign new_P2_U6659 = ~new_P2_R2267_U87 | ~new_P2_U2587;
  assign new_P2_U6660 = ~new_P2_U2588 | ~new_P2_R2096_U97;
  assign new_P2_U6661 = ~P2_EBX_REG_10_ | ~new_P2_U7743;
  assign new_P2_U6662 = ~new_P2_U2392 | ~new_P2_R2099_U93;
  assign new_P2_U6663 = ~new_P2_U2383 | ~new_P2_R2337_U90;
  assign new_P2_U6664 = ~new_P2_R1957_U6 | ~new_P2_U2382;
  assign new_P2_U6665 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_10_;
  assign new_P2_U6666 = ~new_P2_U6570 | ~P2_REIP_REG_10_;
  assign new_P2_U6667 = ~new_P2_R2267_U6 | ~new_P2_U2587;
  assign new_P2_U6668 = ~new_P2_U2588 | ~new_P2_R2096_U96;
  assign new_P2_U6669 = ~P2_EBX_REG_11_ | ~new_P2_U7743;
  assign new_P2_U6670 = ~new_P2_U2392 | ~new_P2_R2099_U92;
  assign new_P2_U6671 = ~new_P2_U2383 | ~new_P2_R2337_U89;
  assign new_P2_U6672 = ~new_P2_R1957_U82 | ~new_P2_U2382;
  assign new_P2_U6673 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_11_;
  assign new_P2_U6674 = ~new_P2_U6570 | ~P2_REIP_REG_11_;
  assign new_P2_U6675 = ~new_P2_R2267_U85 | ~new_P2_U2587;
  assign new_P2_U6676 = ~new_P2_U2588 | ~new_P2_R2096_U95;
  assign new_P2_U6677 = ~P2_EBX_REG_12_ | ~new_P2_U7743;
  assign new_P2_U6678 = ~new_P2_U2392 | ~new_P2_R2099_U91;
  assign new_P2_U6679 = ~new_P2_U2383 | ~new_P2_R2337_U88;
  assign new_P2_U6680 = ~new_P2_R1957_U7 | ~new_P2_U2382;
  assign new_P2_U6681 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_12_;
  assign new_P2_U6682 = ~new_P2_U6570 | ~P2_REIP_REG_12_;
  assign new_P2_U6683 = ~new_P2_R2267_U7 | ~new_P2_U2587;
  assign new_P2_U6684 = ~new_P2_U2588 | ~new_P2_R2096_U94;
  assign new_P2_U6685 = ~P2_EBX_REG_13_ | ~new_P2_U7743;
  assign new_P2_U6686 = ~new_P2_U2392 | ~new_P2_R2099_U90;
  assign new_P2_U6687 = ~new_P2_U2383 | ~new_P2_R2337_U87;
  assign new_P2_U6688 = ~new_P2_R1957_U80 | ~new_P2_U2382;
  assign new_P2_U6689 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_13_;
  assign new_P2_U6690 = ~new_P2_U6570 | ~P2_REIP_REG_13_;
  assign new_P2_U6691 = ~new_P2_R2267_U83 | ~new_P2_U2587;
  assign new_P2_U6692 = ~new_P2_U2588 | ~new_P2_R2096_U93;
  assign new_P2_U6693 = ~P2_EBX_REG_14_ | ~new_P2_U7743;
  assign new_P2_U6694 = ~new_P2_U2392 | ~new_P2_R2099_U89;
  assign new_P2_U6695 = ~new_P2_U2383 | ~new_P2_R2337_U86;
  assign new_P2_U6696 = ~new_P2_R1957_U8 | ~new_P2_U2382;
  assign new_P2_U6697 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_14_;
  assign new_P2_U6698 = ~new_P2_U6570 | ~P2_REIP_REG_14_;
  assign new_P2_U6699 = ~new_P2_R2267_U8 | ~new_P2_U2587;
  assign new_P2_U6700 = ~new_P2_U2588 | ~new_P2_R2096_U92;
  assign new_P2_U6701 = ~P2_EBX_REG_15_ | ~new_P2_U7743;
  assign new_P2_U6702 = ~new_P2_U2392 | ~new_P2_R2099_U88;
  assign new_P2_U6703 = ~new_P2_U2383 | ~new_P2_R2337_U85;
  assign new_P2_U6704 = ~new_P2_R1957_U78 | ~new_P2_U2382;
  assign new_P2_U6705 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_15_;
  assign new_P2_U6706 = ~new_P2_U6570 | ~P2_REIP_REG_15_;
  assign new_P2_U6707 = ~new_P2_R2267_U81 | ~new_P2_U2587;
  assign new_P2_U6708 = ~new_P2_U2588 | ~new_P2_R2096_U91;
  assign new_P2_U6709 = ~P2_EBX_REG_16_ | ~new_P2_U7743;
  assign new_P2_U6710 = ~new_P2_U2392 | ~new_P2_R2099_U87;
  assign new_P2_U6711 = ~new_P2_U2383 | ~new_P2_R2337_U84;
  assign new_P2_U6712 = ~new_P2_R1957_U9 | ~new_P2_U2382;
  assign new_P2_U6713 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_16_;
  assign new_P2_U6714 = ~new_P2_U6570 | ~P2_REIP_REG_16_;
  assign new_P2_U6715 = ~new_P2_R2267_U9 | ~new_P2_U2587;
  assign new_P2_U6716 = ~new_P2_U2588 | ~new_P2_R2096_U90;
  assign new_P2_U6717 = ~P2_EBX_REG_17_ | ~new_P2_U7743;
  assign new_P2_U6718 = ~new_P2_U2392 | ~new_P2_R2099_U86;
  assign new_P2_U6719 = ~new_P2_U2383 | ~new_P2_R2337_U83;
  assign new_P2_U6720 = ~new_P2_R1957_U76 | ~new_P2_U2382;
  assign new_P2_U6721 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_17_;
  assign new_P2_U6722 = ~new_P2_U6570 | ~P2_REIP_REG_17_;
  assign new_P2_U6723 = ~new_P2_R2267_U79 | ~new_P2_U2587;
  assign new_P2_U6724 = ~new_P2_U2588 | ~new_P2_R2096_U89;
  assign new_P2_U6725 = ~P2_EBX_REG_18_ | ~new_P2_U7743;
  assign new_P2_U6726 = ~new_P2_U2392 | ~new_P2_R2099_U85;
  assign new_P2_U6727 = ~new_P2_U2383 | ~new_P2_R2337_U82;
  assign new_P2_U6728 = ~new_P2_R1957_U10 | ~new_P2_U2382;
  assign new_P2_U6729 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_18_;
  assign new_P2_U6730 = ~new_P2_U6570 | ~P2_REIP_REG_18_;
  assign new_P2_U6731 = ~new_P2_R2267_U10 | ~new_P2_U2587;
  assign new_P2_U6732 = ~new_P2_U2588 | ~new_P2_R2096_U88;
  assign new_P2_U6733 = ~P2_EBX_REG_19_ | ~new_P2_U7743;
  assign new_P2_U6734 = ~new_P2_U2392 | ~new_P2_R2099_U84;
  assign new_P2_U6735 = ~new_P2_U2383 | ~new_P2_R2337_U81;
  assign new_P2_U6736 = ~new_P2_R1957_U74 | ~new_P2_U2382;
  assign new_P2_U6737 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_19_;
  assign new_P2_U6738 = ~new_P2_U6570 | ~P2_REIP_REG_19_;
  assign new_P2_U6739 = ~new_P2_R2267_U75 | ~new_P2_U2587;
  assign new_P2_U6740 = ~new_P2_U2588 | ~new_P2_R2096_U87;
  assign new_P2_U6741 = ~P2_EBX_REG_20_ | ~new_P2_U7743;
  assign new_P2_U6742 = ~new_P2_U2392 | ~new_P2_R2099_U83;
  assign new_P2_U6743 = ~new_P2_U2383 | ~new_P2_R2337_U80;
  assign new_P2_U6744 = ~new_P2_R1957_U11 | ~new_P2_U2382;
  assign new_P2_U6745 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_20_;
  assign new_P2_U6746 = ~new_P2_U6570 | ~P2_REIP_REG_20_;
  assign new_P2_U6747 = ~new_P2_R2267_U11 | ~new_P2_U2587;
  assign new_P2_U6748 = ~new_P2_U2588 | ~new_P2_R2096_U86;
  assign new_P2_U6749 = ~P2_EBX_REG_21_ | ~new_P2_U7743;
  assign new_P2_U6750 = ~new_P2_U2392 | ~new_P2_R2099_U82;
  assign new_P2_U6751 = ~new_P2_U2383 | ~new_P2_R2337_U79;
  assign new_P2_U6752 = ~new_P2_R1957_U70 | ~new_P2_U2382;
  assign new_P2_U6753 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_21_;
  assign new_P2_U6754 = ~new_P2_U6570 | ~P2_REIP_REG_21_;
  assign new_P2_U6755 = ~new_P2_R2267_U73 | ~new_P2_U2587;
  assign new_P2_U6756 = ~new_P2_U2588 | ~new_P2_R2096_U85;
  assign new_P2_U6757 = ~P2_EBX_REG_22_ | ~new_P2_U7743;
  assign new_P2_U6758 = ~new_P2_U2392 | ~new_P2_R2099_U81;
  assign new_P2_U6759 = ~new_P2_U2383 | ~new_P2_R2337_U78;
  assign new_P2_U6760 = ~new_P2_R1957_U12 | ~new_P2_U2382;
  assign new_P2_U6761 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_22_;
  assign new_P2_U6762 = ~new_P2_U6570 | ~P2_REIP_REG_22_;
  assign new_P2_U6763 = ~new_P2_R2267_U12 | ~new_P2_U2587;
  assign new_P2_U6764 = ~new_P2_U2588 | ~new_P2_R2096_U84;
  assign new_P2_U6765 = ~P2_EBX_REG_23_ | ~new_P2_U7743;
  assign new_P2_U6766 = ~new_P2_U2392 | ~new_P2_R2099_U80;
  assign new_P2_U6767 = ~new_P2_U2383 | ~new_P2_R2337_U77;
  assign new_P2_U6768 = ~new_P2_R1957_U68 | ~new_P2_U2382;
  assign new_P2_U6769 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_23_;
  assign new_P2_U6770 = ~new_P2_U6570 | ~P2_REIP_REG_23_;
  assign new_P2_U6771 = ~new_P2_R2267_U71 | ~new_P2_U2587;
  assign new_P2_U6772 = ~new_P2_U2588 | ~new_P2_R2096_U83;
  assign new_P2_U6773 = ~P2_EBX_REG_24_ | ~new_P2_U7743;
  assign new_P2_U6774 = ~new_P2_U2392 | ~new_P2_R2099_U79;
  assign new_P2_U6775 = ~new_P2_U2383 | ~new_P2_R2337_U76;
  assign new_P2_U6776 = ~new_P2_R1957_U13 | ~new_P2_U2382;
  assign new_P2_U6777 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_24_;
  assign new_P2_U6778 = ~new_P2_U6570 | ~P2_REIP_REG_24_;
  assign new_P2_U6779 = ~new_P2_R2267_U13 | ~new_P2_U2587;
  assign new_P2_U6780 = ~new_P2_U2588 | ~new_P2_R2096_U82;
  assign new_P2_U6781 = ~P2_EBX_REG_25_ | ~new_P2_U7743;
  assign new_P2_U6782 = ~new_P2_U2392 | ~new_P2_R2099_U78;
  assign new_P2_U6783 = ~new_P2_U2383 | ~new_P2_R2337_U75;
  assign new_P2_U6784 = ~new_P2_R1957_U66 | ~new_P2_U2382;
  assign new_P2_U6785 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_25_;
  assign new_P2_U6786 = ~new_P2_U6570 | ~P2_REIP_REG_25_;
  assign new_P2_U6787 = ~new_P2_R2267_U69 | ~new_P2_U2587;
  assign new_P2_U6788 = ~new_P2_U2588 | ~new_P2_R2096_U81;
  assign new_P2_U6789 = ~P2_EBX_REG_26_ | ~new_P2_U7743;
  assign new_P2_U6790 = ~new_P2_U2392 | ~new_P2_R2099_U77;
  assign new_P2_U6791 = ~new_P2_U2383 | ~new_P2_R2337_U74;
  assign new_P2_U6792 = ~new_P2_R1957_U14 | ~new_P2_U2382;
  assign new_P2_U6793 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_26_;
  assign new_P2_U6794 = ~new_P2_U6570 | ~P2_REIP_REG_26_;
  assign new_P2_U6795 = ~new_P2_R2267_U14 | ~new_P2_U2587;
  assign new_P2_U6796 = ~new_P2_U2588 | ~new_P2_R2096_U80;
  assign new_P2_U6797 = ~P2_EBX_REG_27_ | ~new_P2_U7743;
  assign new_P2_U6798 = ~new_P2_U2392 | ~new_P2_R2099_U76;
  assign new_P2_U6799 = ~new_P2_U2383 | ~new_P2_R2337_U73;
  assign new_P2_U6800 = ~new_P2_R1957_U64 | ~new_P2_U2382;
  assign new_P2_U6801 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_27_;
  assign new_P2_U6802 = ~new_P2_U6570 | ~P2_REIP_REG_27_;
  assign new_P2_U6803 = ~new_P2_R2267_U67 | ~new_P2_U2587;
  assign new_P2_U6804 = ~new_P2_U2588 | ~new_P2_R2096_U79;
  assign new_P2_U6805 = ~P2_EBX_REG_28_ | ~new_P2_U7743;
  assign new_P2_U6806 = ~new_P2_U2392 | ~new_P2_R2099_U75;
  assign new_P2_U6807 = ~new_P2_U2383 | ~new_P2_R2337_U72;
  assign new_P2_U6808 = ~new_P2_R1957_U15 | ~new_P2_U2382;
  assign new_P2_U6809 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_28_;
  assign new_P2_U6810 = ~new_P2_U6570 | ~P2_REIP_REG_28_;
  assign new_P2_U6811 = ~new_P2_R2267_U15 | ~new_P2_U2587;
  assign new_P2_U6812 = ~new_P2_U2588 | ~new_P2_R2096_U78;
  assign new_P2_U6813 = ~P2_EBX_REG_29_ | ~new_P2_U7743;
  assign new_P2_U6814 = ~new_P2_U2392 | ~new_P2_R2099_U74;
  assign new_P2_U6815 = ~new_P2_U2383 | ~new_P2_R2337_U71;
  assign new_P2_U6816 = ~new_P2_R1957_U16 | ~new_P2_U2382;
  assign new_P2_U6817 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_29_;
  assign new_P2_U6818 = ~new_P2_U6570 | ~P2_REIP_REG_29_;
  assign new_P2_U6819 = ~new_P2_R2267_U16 | ~new_P2_U2587;
  assign new_P2_U6820 = ~new_P2_U2588 | ~new_P2_R2096_U76;
  assign new_P2_U6821 = ~P2_EBX_REG_30_ | ~new_P2_U7743;
  assign new_P2_U6822 = ~new_P2_U2392 | ~new_P2_R2099_U73;
  assign new_P2_U6823 = ~new_P2_U2383 | ~new_P2_R2337_U69;
  assign new_P2_U6824 = ~new_P2_R1957_U62 | ~new_P2_U2382;
  assign new_P2_U6825 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_30_;
  assign new_P2_U6826 = ~new_P2_U6570 | ~P2_REIP_REG_30_;
  assign new_P2_U6827 = ~new_P2_R2267_U63 | ~new_P2_U2587;
  assign new_P2_U6828 = ~new_P2_U2588 | ~new_P2_R2096_U50;
  assign new_P2_U6829 = ~P2_EBX_REG_31_ | ~new_P2_U7743;
  assign new_P2_U6830 = ~new_P2_U2392 | ~new_P2_R2099_U72;
  assign new_P2_U6831 = ~new_P2_U2383 | ~new_P2_R2337_U68;
  assign new_P2_U6832 = ~new_P2_R1957_U50 | ~new_P2_U2382;
  assign new_P2_U6833 = ~new_P2_U2378 | ~P2_PHYADDRPOINTER_REG_31_;
  assign new_P2_U6834 = ~new_P2_U6570 | ~P2_REIP_REG_31_;
  assign new_P2_U6835 = ~P2_DATAWIDTH_REG_1_ | ~P2_DATAWIDTH_REG_0_;
  assign new_P2_U6836 = ~new_P2_U4477 | ~P2_REIP_REG_0_;
  assign new_P2_U6837 = ~P2_BYTEENABLE_REG_1_ | ~new_P2_U3547;
  assign new_P2_U6838 = ~new_P2_U4400;
  assign new_P2_U6839 = ~new_P2_U4399 | ~new_P2_U4426 | ~new_P2_U4468;
  assign new_P2_U6840 = ~P2_FLUSH_REG | ~new_P2_U4400;
  assign new_P2_U6841 = ~new_P2_U4187 | ~new_P2_U4467;
  assign new_P2_U6842 = ~new_P2_U4466 | ~new_P2_U3284;
  assign new_P2_U6843 = ~new_P2_U4402;
  assign new_P2_U6844 = ~new_P2_U4411 | ~P2_STATEBS16_REG;
  assign new_P2_U6845 = ~new_P2_U2715;
  assign new_P2_U6846 = ~new_P2_U2715 | ~new_P2_U3536;
  assign new_P2_U6847 = ~new_P2_U4411 | ~new_P2_U3265;
  assign new_P2_U6848 = ~new_P2_U4184 | ~new_P2_U2356;
  assign new_P2_U6849 = ~new_P2_U4418 | ~new_P2_U6847;
  assign new_P2_U6850 = ~new_U211 | ~new_P2_U6846;
  assign new_P2_U6851 = P2_STATE2_REG_2_ | P2_STATE2_REG_1_;
  assign new_P2_U6852 = ~new_P2_U4186 | ~new_P2_U6851 | ~new_P2_U6850;
  assign new_P2_U6853 = ~new_P2_U2374 | ~new_P2_U2459;
  assign new_P2_U6854 = ~P2_CODEFETCH_REG | ~new_P2_U6853;
  assign new_P2_U6855 = ~new_P2_U4461 | ~P2_STATE2_REG_0_;
  assign new_P2_U6856 = ~P2_ADS_N_REG | ~P2_STATE_REG_0_;
  assign new_P2_U6857 = ~new_P2_U4403;
  assign new_P2_U6858 = ~new_P2_U3294 | ~P2_STATE2_REG_2_ | ~new_P2_U3286;
  assign new_P2_U6859 = ~new_P2_U4404 | ~new_P2_U4421 | ~new_P2_U4468;
  assign new_P2_U6860 = ~new_P2_U4189 | ~new_P2_U2446;
  assign new_P2_U6861 = ~P2_MEMORYFETCH_REG | ~new_P2_U6859;
  assign new_P2_U6862 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__7_;
  assign new_P2_U6863 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__7_;
  assign new_P2_U6864 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__7_;
  assign new_P2_U6865 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__7_;
  assign new_P2_U6866 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__7_;
  assign new_P2_U6867 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__7_;
  assign new_P2_U6868 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__7_;
  assign new_P2_U6869 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__7_;
  assign new_P2_U6870 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__7_;
  assign new_P2_U6871 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__7_;
  assign new_P2_U6872 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__7_;
  assign new_P2_U6873 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__7_;
  assign new_P2_U6874 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__7_;
  assign new_P2_U6875 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__7_;
  assign new_P2_U6876 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__7_;
  assign new_P2_U6877 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__7_;
  assign new_P2_U6878 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__7_;
  assign new_P2_U6879 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__7_;
  assign new_P2_U6880 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__7_;
  assign new_P2_U6881 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__7_;
  assign new_P2_U6882 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__7_;
  assign new_P2_U6883 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__7_;
  assign new_P2_U6884 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__7_;
  assign new_P2_U6885 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__7_;
  assign new_P2_U6886 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__7_;
  assign new_P2_U6887 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__7_;
  assign new_P2_U6888 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__7_;
  assign new_P2_U6889 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__7_;
  assign new_P2_U6890 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__7_;
  assign new_P2_U6891 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__7_;
  assign new_P2_U6892 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__7_;
  assign new_P2_U6893 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__7_;
  assign new_P2_U6894 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__6_;
  assign new_P2_U6895 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__6_;
  assign new_P2_U6896 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__6_;
  assign new_P2_U6897 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__6_;
  assign new_P2_U6898 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__6_;
  assign new_P2_U6899 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__6_;
  assign new_P2_U6900 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__6_;
  assign new_P2_U6901 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__6_;
  assign new_P2_U6902 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__6_;
  assign new_P2_U6903 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__6_;
  assign new_P2_U6904 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__6_;
  assign new_P2_U6905 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__6_;
  assign new_P2_U6906 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__6_;
  assign new_P2_U6907 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__6_;
  assign new_P2_U6908 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__6_;
  assign new_P2_U6909 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__6_;
  assign new_P2_U6910 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__5_;
  assign new_P2_U6911 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__5_;
  assign new_P2_U6912 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__5_;
  assign new_P2_U6913 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__5_;
  assign new_P2_U6914 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__5_;
  assign new_P2_U6915 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__5_;
  assign new_P2_U6916 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__5_;
  assign new_P2_U6917 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__5_;
  assign new_P2_U6918 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__5_;
  assign new_P2_U6919 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__5_;
  assign new_P2_U6920 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__5_;
  assign new_P2_U6921 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__5_;
  assign new_P2_U6922 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__5_;
  assign new_P2_U6923 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__5_;
  assign new_P2_U6924 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__5_;
  assign new_P2_U6925 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__5_;
  assign new_P2_U6926 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__4_;
  assign new_P2_U6927 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__4_;
  assign new_P2_U6928 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__4_;
  assign new_P2_U6929 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__4_;
  assign new_P2_U6930 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__4_;
  assign new_P2_U6931 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__4_;
  assign new_P2_U6932 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__4_;
  assign new_P2_U6933 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__4_;
  assign new_P2_U6934 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__4_;
  assign new_P2_U6935 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__4_;
  assign new_P2_U6936 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__4_;
  assign new_P2_U6937 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__4_;
  assign new_P2_U6938 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__4_;
  assign new_P2_U6939 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__4_;
  assign new_P2_U6940 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__4_;
  assign new_P2_U6941 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__4_;
  assign new_P2_U6942 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__3_;
  assign new_P2_U6943 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__3_;
  assign new_P2_U6944 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__3_;
  assign new_P2_U6945 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__3_;
  assign new_P2_U6946 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__3_;
  assign new_P2_U6947 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__3_;
  assign new_P2_U6948 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__3_;
  assign new_P2_U6949 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__3_;
  assign new_P2_U6950 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__3_;
  assign new_P2_U6951 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__3_;
  assign new_P2_U6952 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__3_;
  assign new_P2_U6953 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__3_;
  assign new_P2_U6954 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__3_;
  assign new_P2_U6955 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__3_;
  assign new_P2_U6956 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__3_;
  assign new_P2_U6957 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__3_;
  assign new_P2_U6958 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__2_;
  assign new_P2_U6959 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__2_;
  assign new_P2_U6960 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__2_;
  assign new_P2_U6961 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__2_;
  assign new_P2_U6962 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__2_;
  assign new_P2_U6963 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__2_;
  assign new_P2_U6964 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__2_;
  assign new_P2_U6965 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__2_;
  assign new_P2_U6966 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__2_;
  assign new_P2_U6967 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__2_;
  assign new_P2_U6968 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__2_;
  assign new_P2_U6969 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__2_;
  assign new_P2_U6970 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__2_;
  assign new_P2_U6971 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__2_;
  assign new_P2_U6972 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__2_;
  assign new_P2_U6973 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__2_;
  assign new_P2_U6974 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__1_;
  assign new_P2_U6975 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__1_;
  assign new_P2_U6976 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__1_;
  assign new_P2_U6977 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__1_;
  assign new_P2_U6978 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__1_;
  assign new_P2_U6979 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__1_;
  assign new_P2_U6980 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__1_;
  assign new_P2_U6981 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__1_;
  assign new_P2_U6982 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__1_;
  assign new_P2_U6983 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__1_;
  assign new_P2_U6984 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__1_;
  assign new_P2_U6985 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__1_;
  assign new_P2_U6986 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__1_;
  assign new_P2_U6987 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__1_;
  assign new_P2_U6988 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__1_;
  assign new_P2_U6989 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__1_;
  assign new_P2_U6990 = ~new_P2_U2562 | ~P2_INSTQUEUE_REG_15__0_;
  assign new_P2_U6991 = ~new_P2_U2561 | ~P2_INSTQUEUE_REG_14__0_;
  assign new_P2_U6992 = ~new_P2_U2560 | ~P2_INSTQUEUE_REG_13__0_;
  assign new_P2_U6993 = ~new_P2_U2559 | ~P2_INSTQUEUE_REG_12__0_;
  assign new_P2_U6994 = ~new_P2_U2558 | ~P2_INSTQUEUE_REG_11__0_;
  assign new_P2_U6995 = ~new_P2_U2557 | ~P2_INSTQUEUE_REG_10__0_;
  assign new_P2_U6996 = ~new_P2_U2555 | ~P2_INSTQUEUE_REG_9__0_;
  assign new_P2_U6997 = ~new_P2_U2554 | ~P2_INSTQUEUE_REG_8__0_;
  assign new_P2_U6998 = ~new_P2_U2552 | ~P2_INSTQUEUE_REG_7__0_;
  assign new_P2_U6999 = ~new_P2_U2551 | ~P2_INSTQUEUE_REG_6__0_;
  assign new_P2_U7000 = ~new_P2_U2550 | ~P2_INSTQUEUE_REG_5__0_;
  assign new_P2_U7001 = ~new_P2_U2548 | ~P2_INSTQUEUE_REG_4__0_;
  assign new_P2_U7002 = ~new_P2_U2546 | ~P2_INSTQUEUE_REG_3__0_;
  assign new_P2_U7003 = ~new_P2_U2545 | ~P2_INSTQUEUE_REG_2__0_;
  assign new_P2_U7004 = ~new_P2_U2543 | ~P2_INSTQUEUE_REG_1__0_;
  assign new_P2_U7005 = ~new_P2_U2541 | ~P2_INSTQUEUE_REG_0__0_;
  assign new_P2_U7006 = P2_INSTQUEUERD_ADDR_REG_0_ | P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U7007 = ~new_P2_U4405;
  assign new_P2_U7008 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__7_;
  assign new_P2_U7009 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__7_;
  assign new_P2_U7010 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__7_;
  assign new_P2_U7011 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__7_;
  assign new_P2_U7012 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__7_;
  assign new_P2_U7013 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__7_;
  assign new_P2_U7014 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__7_;
  assign new_P2_U7015 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__7_;
  assign new_P2_U7016 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__7_;
  assign new_P2_U7017 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__7_;
  assign new_P2_U7018 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__7_;
  assign new_P2_U7019 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__7_;
  assign new_P2_U7020 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__7_;
  assign new_P2_U7021 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__7_;
  assign new_P2_U7022 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__7_;
  assign new_P2_U7023 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__7_;
  assign new_P2_U7024 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__6_;
  assign new_P2_U7025 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__6_;
  assign new_P2_U7026 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__6_;
  assign new_P2_U7027 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__6_;
  assign new_P2_U7028 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__6_;
  assign new_P2_U7029 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__6_;
  assign new_P2_U7030 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__6_;
  assign new_P2_U7031 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__6_;
  assign new_P2_U7032 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__6_;
  assign new_P2_U7033 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__6_;
  assign new_P2_U7034 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__6_;
  assign new_P2_U7035 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__6_;
  assign new_P2_U7036 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__6_;
  assign new_P2_U7037 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__6_;
  assign new_P2_U7038 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__6_;
  assign new_P2_U7039 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__6_;
  assign new_P2_U7040 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__5_;
  assign new_P2_U7041 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__5_;
  assign new_P2_U7042 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__5_;
  assign new_P2_U7043 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__5_;
  assign new_P2_U7044 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__5_;
  assign new_P2_U7045 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__5_;
  assign new_P2_U7046 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__5_;
  assign new_P2_U7047 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__5_;
  assign new_P2_U7048 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__5_;
  assign new_P2_U7049 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__5_;
  assign new_P2_U7050 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__5_;
  assign new_P2_U7051 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__5_;
  assign new_P2_U7052 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__5_;
  assign new_P2_U7053 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__5_;
  assign new_P2_U7054 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__5_;
  assign new_P2_U7055 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__5_;
  assign new_P2_U7056 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__4_;
  assign new_P2_U7057 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__4_;
  assign new_P2_U7058 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__4_;
  assign new_P2_U7059 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__4_;
  assign new_P2_U7060 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__4_;
  assign new_P2_U7061 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__4_;
  assign new_P2_U7062 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__4_;
  assign new_P2_U7063 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__4_;
  assign new_P2_U7064 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__4_;
  assign new_P2_U7065 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__4_;
  assign new_P2_U7066 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__4_;
  assign new_P2_U7067 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__4_;
  assign new_P2_U7068 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__4_;
  assign new_P2_U7069 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__4_;
  assign new_P2_U7070 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__4_;
  assign new_P2_U7071 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__4_;
  assign new_P2_U7072 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__3_;
  assign new_P2_U7073 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__3_;
  assign new_P2_U7074 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__3_;
  assign new_P2_U7075 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__3_;
  assign new_P2_U7076 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__3_;
  assign new_P2_U7077 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__3_;
  assign new_P2_U7078 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__3_;
  assign new_P2_U7079 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__3_;
  assign new_P2_U7080 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__3_;
  assign new_P2_U7081 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__3_;
  assign new_P2_U7082 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__3_;
  assign new_P2_U7083 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__3_;
  assign new_P2_U7084 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__3_;
  assign new_P2_U7085 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__3_;
  assign new_P2_U7086 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__3_;
  assign new_P2_U7087 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__3_;
  assign new_P2_U7088 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__2_;
  assign new_P2_U7089 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__2_;
  assign new_P2_U7090 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__2_;
  assign new_P2_U7091 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__2_;
  assign new_P2_U7092 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__2_;
  assign new_P2_U7093 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__2_;
  assign new_P2_U7094 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__2_;
  assign new_P2_U7095 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__2_;
  assign new_P2_U7096 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__2_;
  assign new_P2_U7097 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__2_;
  assign new_P2_U7098 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__2_;
  assign new_P2_U7099 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__2_;
  assign new_P2_U7100 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__2_;
  assign new_P2_U7101 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__2_;
  assign new_P2_U7102 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__2_;
  assign new_P2_U7103 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__2_;
  assign new_P2_U7104 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__1_;
  assign new_P2_U7105 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__1_;
  assign new_P2_U7106 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__1_;
  assign new_P2_U7107 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__1_;
  assign new_P2_U7108 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__1_;
  assign new_P2_U7109 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__1_;
  assign new_P2_U7110 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__1_;
  assign new_P2_U7111 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__1_;
  assign new_P2_U7112 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__1_;
  assign new_P2_U7113 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__1_;
  assign new_P2_U7114 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__1_;
  assign new_P2_U7115 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__1_;
  assign new_P2_U7116 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__1_;
  assign new_P2_U7117 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__1_;
  assign new_P2_U7118 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__1_;
  assign new_P2_U7119 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__1_;
  assign new_P2_U7120 = ~new_P2_U2586 | ~P2_INSTQUEUE_REG_0__0_;
  assign new_P2_U7121 = ~new_P2_U2585 | ~P2_INSTQUEUE_REG_1__0_;
  assign new_P2_U7122 = ~new_P2_U2584 | ~P2_INSTQUEUE_REG_2__0_;
  assign new_P2_U7123 = ~new_P2_U2583 | ~P2_INSTQUEUE_REG_3__0_;
  assign new_P2_U7124 = ~new_P2_U2581 | ~P2_INSTQUEUE_REG_4__0_;
  assign new_P2_U7125 = ~new_P2_U2580 | ~P2_INSTQUEUE_REG_5__0_;
  assign new_P2_U7126 = ~new_P2_U2579 | ~P2_INSTQUEUE_REG_6__0_;
  assign new_P2_U7127 = ~new_P2_U2578 | ~P2_INSTQUEUE_REG_7__0_;
  assign new_P2_U7128 = ~new_P2_U2576 | ~P2_INSTQUEUE_REG_8__0_;
  assign new_P2_U7129 = ~new_P2_U2575 | ~P2_INSTQUEUE_REG_9__0_;
  assign new_P2_U7130 = ~new_P2_U2574 | ~P2_INSTQUEUE_REG_10__0_;
  assign new_P2_U7131 = ~new_P2_U2573 | ~P2_INSTQUEUE_REG_11__0_;
  assign new_P2_U7132 = ~new_P2_U2571 | ~P2_INSTQUEUE_REG_12__0_;
  assign new_P2_U7133 = ~new_P2_U2569 | ~P2_INSTQUEUE_REG_13__0_;
  assign new_P2_U7134 = ~new_P2_U2567 | ~P2_INSTQUEUE_REG_14__0_;
  assign new_P2_U7135 = ~new_P2_U2565 | ~P2_INSTQUEUE_REG_15__0_;
  assign new_P2_U7136 = ~new_P2_U3554;
  assign new_P2_U7137 = ~new_P2_U7136 | ~new_P2_U3300;
  assign new_P2_U7138 = ~new_P2_U4467 | ~new_P2_R2099_U95;
  assign new_P2_U7139 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U7137;
  assign new_P2_U7140 = ~new_P2_U4430 | ~new_P2_U3428;
  assign new_P2_U7141 = ~new_P2_ADD_402_1132_U23 | ~new_P2_U2355;
  assign new_P2_U7142 = ~new_P2_U2354 | ~new_P2_U2606;
  assign new_P2_U7143 = ~new_P2_U2605 | ~new_P2_U2355;
  assign new_P2_U7144 = ~new_P2_U2354 | ~new_P2_U2605;
  assign new_P2_U7145 = ~new_P2_U2604 | ~new_P2_U2355;
  assign new_P2_U7146 = ~new_P2_U2354 | ~new_P2_U2604;
  assign new_P2_U7147 = ~new_P2_U2603 | ~new_P2_U2355;
  assign new_P2_U7148 = ~new_P2_U2354 | ~new_P2_U2603;
  assign new_P2_U7149 = ~new_P2_U4467 | ~new_P2_R2099_U96;
  assign new_P2_U7150 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U7137;
  assign new_P2_U7151 = ~new_P2_U4430 | ~new_P2_U3580;
  assign new_P2_U7152 = ~new_P2_U2602 | ~new_P2_U2355;
  assign new_P2_U7153 = ~new_P2_U2354 | ~new_P2_U2602;
  assign new_P2_U7154 = ~new_P2_U2601 | ~new_P2_U2355;
  assign new_P2_U7155 = ~new_P2_U2354 | ~new_P2_U2601;
  assign new_P2_U7156 = ~new_P2_U2600 | ~new_P2_U2355;
  assign new_P2_U7157 = ~new_P2_U2354 | ~new_P2_U2600;
  assign new_P2_U7158 = ~new_P2_U2599 | ~new_P2_U2355;
  assign new_P2_U7159 = ~new_P2_U2354 | ~new_P2_U2599;
  assign new_P2_U7160 = ~new_P2_U4467 | ~new_P2_R2099_U5;
  assign new_P2_U7161 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U7137;
  assign new_P2_U7162 = ~new_P2_U4430 | ~new_P2_U3243;
  assign new_P2_U7163 = ~new_P2_U4467 | ~new_P2_R2099_U94;
  assign new_P2_U7164 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_U7137;
  assign new_P2_U7165 = ~new_P2_U4430 | ~new_P2_U3307;
  assign new_P2_U7166 = ~P2_INSTQUEUE_REG_0__0_ | ~new_P2_U2355;
  assign new_P2_U7167 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__7_;
  assign new_P2_U7168 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__7_;
  assign new_P2_U7169 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__7_;
  assign new_P2_U7170 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__7_;
  assign new_P2_U7171 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__7_;
  assign new_P2_U7172 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__7_;
  assign new_P2_U7173 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__7_;
  assign new_P2_U7174 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__7_;
  assign new_P2_U7175 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__7_;
  assign new_P2_U7176 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__7_;
  assign new_P2_U7177 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__7_;
  assign new_P2_U7178 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__7_;
  assign new_P2_U7179 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__7_;
  assign new_P2_U7180 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__7_;
  assign new_P2_U7181 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__7_;
  assign new_P2_U7182 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__7_;
  assign new_P2_U7183 = ~new_P2_U4277 | ~new_P2_U4278 | ~new_P2_U4280 | ~new_P2_U4279;
  assign new_P2_U7184 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__6_;
  assign new_P2_U7185 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__6_;
  assign new_P2_U7186 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__6_;
  assign new_P2_U7187 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__6_;
  assign new_P2_U7188 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__6_;
  assign new_P2_U7189 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__6_;
  assign new_P2_U7190 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__6_;
  assign new_P2_U7191 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__6_;
  assign new_P2_U7192 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__6_;
  assign new_P2_U7193 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__6_;
  assign new_P2_U7194 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__6_;
  assign new_P2_U7195 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__6_;
  assign new_P2_U7196 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__6_;
  assign new_P2_U7197 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__6_;
  assign new_P2_U7198 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__6_;
  assign new_P2_U7199 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__6_;
  assign new_P2_U7200 = ~new_P2_U4281 | ~new_P2_U4282 | ~new_P2_U4284 | ~new_P2_U4283;
  assign new_P2_U7201 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__6_;
  assign new_P2_U7202 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__6_;
  assign new_P2_U7203 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__6_;
  assign new_P2_U7204 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__6_;
  assign new_P2_U7205 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__6_;
  assign new_P2_U7206 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__6_;
  assign new_P2_U7207 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__6_;
  assign new_P2_U7208 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__6_;
  assign new_P2_U7209 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__6_;
  assign new_P2_U7210 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__6_;
  assign new_P2_U7211 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__6_;
  assign new_P2_U7212 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__6_;
  assign new_P2_U7213 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__6_;
  assign new_P2_U7214 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__6_;
  assign new_P2_U7215 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__6_;
  assign new_P2_U7216 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__6_;
  assign new_P2_U7217 = ~new_P2_U4285 | ~new_P2_U4286 | ~new_P2_U4288 | ~new_P2_U4287;
  assign new_P2_U7218 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__5_;
  assign new_P2_U7219 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__5_;
  assign new_P2_U7220 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__5_;
  assign new_P2_U7221 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__5_;
  assign new_P2_U7222 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__5_;
  assign new_P2_U7223 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__5_;
  assign new_P2_U7224 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__5_;
  assign new_P2_U7225 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__5_;
  assign new_P2_U7226 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__5_;
  assign new_P2_U7227 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__5_;
  assign new_P2_U7228 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__5_;
  assign new_P2_U7229 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__5_;
  assign new_P2_U7230 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__5_;
  assign new_P2_U7231 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__5_;
  assign new_P2_U7232 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__5_;
  assign new_P2_U7233 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__5_;
  assign new_P2_U7234 = ~new_P2_U4289 | ~new_P2_U4290 | ~new_P2_U4292 | ~new_P2_U4291;
  assign new_P2_U7235 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__5_;
  assign new_P2_U7236 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__5_;
  assign new_P2_U7237 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__5_;
  assign new_P2_U7238 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__5_;
  assign new_P2_U7239 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__5_;
  assign new_P2_U7240 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__5_;
  assign new_P2_U7241 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__5_;
  assign new_P2_U7242 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__5_;
  assign new_P2_U7243 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__5_;
  assign new_P2_U7244 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__5_;
  assign new_P2_U7245 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__5_;
  assign new_P2_U7246 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__5_;
  assign new_P2_U7247 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__5_;
  assign new_P2_U7248 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__5_;
  assign new_P2_U7249 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__5_;
  assign new_P2_U7250 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__5_;
  assign new_P2_U7251 = ~new_P2_U4293 | ~new_P2_U4294 | ~new_P2_U4296 | ~new_P2_U4295;
  assign new_P2_U7252 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__4_;
  assign new_P2_U7253 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__4_;
  assign new_P2_U7254 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__4_;
  assign new_P2_U7255 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__4_;
  assign new_P2_U7256 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__4_;
  assign new_P2_U7257 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__4_;
  assign new_P2_U7258 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__4_;
  assign new_P2_U7259 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__4_;
  assign new_P2_U7260 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__4_;
  assign new_P2_U7261 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__4_;
  assign new_P2_U7262 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__4_;
  assign new_P2_U7263 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__4_;
  assign new_P2_U7264 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__4_;
  assign new_P2_U7265 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__4_;
  assign new_P2_U7266 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__4_;
  assign new_P2_U7267 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__4_;
  assign new_P2_U7268 = ~new_P2_U4297 | ~new_P2_U4298 | ~new_P2_U4300 | ~new_P2_U4299;
  assign new_P2_U7269 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__4_;
  assign new_P2_U7270 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__4_;
  assign new_P2_U7271 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__4_;
  assign new_P2_U7272 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__4_;
  assign new_P2_U7273 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__4_;
  assign new_P2_U7274 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__4_;
  assign new_P2_U7275 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__4_;
  assign new_P2_U7276 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__4_;
  assign new_P2_U7277 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__4_;
  assign new_P2_U7278 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__4_;
  assign new_P2_U7279 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__4_;
  assign new_P2_U7280 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__4_;
  assign new_P2_U7281 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__4_;
  assign new_P2_U7282 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__4_;
  assign new_P2_U7283 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__4_;
  assign new_P2_U7284 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__4_;
  assign new_P2_U7285 = ~new_P2_U4301 | ~new_P2_U4302 | ~new_P2_U4304 | ~new_P2_U4303;
  assign new_P2_U7286 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__3_;
  assign new_P2_U7287 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__3_;
  assign new_P2_U7288 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__3_;
  assign new_P2_U7289 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__3_;
  assign new_P2_U7290 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__3_;
  assign new_P2_U7291 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__3_;
  assign new_P2_U7292 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__3_;
  assign new_P2_U7293 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__3_;
  assign new_P2_U7294 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__3_;
  assign new_P2_U7295 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__3_;
  assign new_P2_U7296 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__3_;
  assign new_P2_U7297 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__3_;
  assign new_P2_U7298 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__3_;
  assign new_P2_U7299 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__3_;
  assign new_P2_U7300 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__3_;
  assign new_P2_U7301 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__3_;
  assign new_P2_U7302 = ~new_P2_U4305 | ~new_P2_U4306 | ~new_P2_U4308 | ~new_P2_U4307;
  assign new_P2_U7303 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__3_;
  assign new_P2_U7304 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__3_;
  assign new_P2_U7305 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__3_;
  assign new_P2_U7306 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__3_;
  assign new_P2_U7307 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__3_;
  assign new_P2_U7308 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__3_;
  assign new_P2_U7309 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__3_;
  assign new_P2_U7310 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__3_;
  assign new_P2_U7311 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__3_;
  assign new_P2_U7312 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__3_;
  assign new_P2_U7313 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__3_;
  assign new_P2_U7314 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__3_;
  assign new_P2_U7315 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__3_;
  assign new_P2_U7316 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__3_;
  assign new_P2_U7317 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__3_;
  assign new_P2_U7318 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__3_;
  assign new_P2_U7319 = ~new_P2_U4309 | ~new_P2_U4310 | ~new_P2_U4312 | ~new_P2_U4311;
  assign new_P2_U7320 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__2_;
  assign new_P2_U7321 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__2_;
  assign new_P2_U7322 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__2_;
  assign new_P2_U7323 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__2_;
  assign new_P2_U7324 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__2_;
  assign new_P2_U7325 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__2_;
  assign new_P2_U7326 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__2_;
  assign new_P2_U7327 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__2_;
  assign new_P2_U7328 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__2_;
  assign new_P2_U7329 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__2_;
  assign new_P2_U7330 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__2_;
  assign new_P2_U7331 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__2_;
  assign new_P2_U7332 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__2_;
  assign new_P2_U7333 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__2_;
  assign new_P2_U7334 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__2_;
  assign new_P2_U7335 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__2_;
  assign new_P2_U7336 = ~new_P2_U4313 | ~new_P2_U4314 | ~new_P2_U4316 | ~new_P2_U4315;
  assign new_P2_U7337 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__2_;
  assign new_P2_U7338 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__2_;
  assign new_P2_U7339 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__2_;
  assign new_P2_U7340 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__2_;
  assign new_P2_U7341 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__2_;
  assign new_P2_U7342 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__2_;
  assign new_P2_U7343 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__2_;
  assign new_P2_U7344 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__2_;
  assign new_P2_U7345 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__2_;
  assign new_P2_U7346 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__2_;
  assign new_P2_U7347 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__2_;
  assign new_P2_U7348 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__2_;
  assign new_P2_U7349 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__2_;
  assign new_P2_U7350 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__2_;
  assign new_P2_U7351 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__2_;
  assign new_P2_U7352 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__2_;
  assign new_P2_U7353 = ~new_P2_U4317 | ~new_P2_U4318 | ~new_P2_U4320 | ~new_P2_U4319;
  assign new_P2_U7354 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__1_;
  assign new_P2_U7355 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__1_;
  assign new_P2_U7356 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__1_;
  assign new_P2_U7357 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__1_;
  assign new_P2_U7358 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__1_;
  assign new_P2_U7359 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__1_;
  assign new_P2_U7360 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__1_;
  assign new_P2_U7361 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__1_;
  assign new_P2_U7362 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__1_;
  assign new_P2_U7363 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__1_;
  assign new_P2_U7364 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__1_;
  assign new_P2_U7365 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__1_;
  assign new_P2_U7366 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__1_;
  assign new_P2_U7367 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__1_;
  assign new_P2_U7368 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__1_;
  assign new_P2_U7369 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__1_;
  assign new_P2_U7370 = ~new_P2_U4321 | ~new_P2_U4322 | ~new_P2_U4324 | ~new_P2_U4323;
  assign new_P2_U7371 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__1_;
  assign new_P2_U7372 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__1_;
  assign new_P2_U7373 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__1_;
  assign new_P2_U7374 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__1_;
  assign new_P2_U7375 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__1_;
  assign new_P2_U7376 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__1_;
  assign new_P2_U7377 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__1_;
  assign new_P2_U7378 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__1_;
  assign new_P2_U7379 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__1_;
  assign new_P2_U7380 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__1_;
  assign new_P2_U7381 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__1_;
  assign new_P2_U7382 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__1_;
  assign new_P2_U7383 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__1_;
  assign new_P2_U7384 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__1_;
  assign new_P2_U7385 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__1_;
  assign new_P2_U7386 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__1_;
  assign new_P2_U7387 = ~new_P2_U4325 | ~new_P2_U4326 | ~new_P2_U4328 | ~new_P2_U4327;
  assign new_P2_U7388 = ~new_P2_U5517 | ~P2_INSTQUEUE_REG_0__0_;
  assign new_P2_U7389 = ~new_P2_U5460 | ~P2_INSTQUEUE_REG_1__0_;
  assign new_P2_U7390 = ~new_P2_U5402 | ~P2_INSTQUEUE_REG_2__0_;
  assign new_P2_U7391 = ~new_P2_U5345 | ~P2_INSTQUEUE_REG_3__0_;
  assign new_P2_U7392 = ~new_P2_U5287 | ~P2_INSTQUEUE_REG_4__0_;
  assign new_P2_U7393 = ~new_P2_U5230 | ~P2_INSTQUEUE_REG_5__0_;
  assign new_P2_U7394 = ~new_P2_U5172 | ~P2_INSTQUEUE_REG_6__0_;
  assign new_P2_U7395 = ~new_P2_U5116 | ~P2_INSTQUEUE_REG_7__0_;
  assign new_P2_U7396 = ~new_P2_U5059 | ~P2_INSTQUEUE_REG_8__0_;
  assign new_P2_U7397 = ~new_P2_U5002 | ~P2_INSTQUEUE_REG_9__0_;
  assign new_P2_U7398 = ~new_P2_U4944 | ~P2_INSTQUEUE_REG_10__0_;
  assign new_P2_U7399 = ~new_P2_U4887 | ~P2_INSTQUEUE_REG_11__0_;
  assign new_P2_U7400 = ~new_P2_U4829 | ~P2_INSTQUEUE_REG_12__0_;
  assign new_P2_U7401 = ~new_P2_U4772 | ~P2_INSTQUEUE_REG_13__0_;
  assign new_P2_U7402 = ~new_P2_U4713 | ~P2_INSTQUEUE_REG_14__0_;
  assign new_P2_U7403 = ~new_P2_U4653 | ~P2_INSTQUEUE_REG_15__0_;
  assign new_P2_U7404 = ~new_P2_U4329 | ~new_P2_U4330 | ~new_P2_U4332 | ~new_P2_U4331;
  assign new_P2_U7405 = ~new_P2_U2538 | ~P2_INSTQUEUE_REG_8__0_;
  assign new_P2_U7406 = ~new_P2_U2537 | ~P2_INSTQUEUE_REG_9__0_;
  assign new_P2_U7407 = ~new_P2_U2536 | ~P2_INSTQUEUE_REG_10__0_;
  assign new_P2_U7408 = ~new_P2_U2535 | ~P2_INSTQUEUE_REG_11__0_;
  assign new_P2_U7409 = ~new_P2_U2534 | ~P2_INSTQUEUE_REG_12__0_;
  assign new_P2_U7410 = ~new_P2_U2533 | ~P2_INSTQUEUE_REG_13__0_;
  assign new_P2_U7411 = ~new_P2_U2531 | ~P2_INSTQUEUE_REG_14__0_;
  assign new_P2_U7412 = ~new_P2_U2530 | ~P2_INSTQUEUE_REG_15__0_;
  assign new_P2_U7413 = ~new_P2_U2528 | ~P2_INSTQUEUE_REG_7__0_;
  assign new_P2_U7414 = ~new_P2_U2527 | ~P2_INSTQUEUE_REG_6__0_;
  assign new_P2_U7415 = ~new_P2_U2526 | ~P2_INSTQUEUE_REG_5__0_;
  assign new_P2_U7416 = ~new_P2_U2524 | ~P2_INSTQUEUE_REG_4__0_;
  assign new_P2_U7417 = ~new_P2_U2522 | ~P2_INSTQUEUE_REG_3__0_;
  assign new_P2_U7418 = ~new_P2_U2521 | ~P2_INSTQUEUE_REG_2__0_;
  assign new_P2_U7419 = ~new_P2_U2519 | ~P2_INSTQUEUE_REG_1__0_;
  assign new_P2_U7420 = ~new_P2_U2517 | ~P2_INSTQUEUE_REG_0__0_;
  assign new_P2_U7421 = ~new_P2_U4333 | ~new_P2_U4334 | ~new_P2_U4336 | ~new_P2_U4335;
  assign new_P2_U7422 = ~new_P2_U2352 | ~new_P2_U7319;
  assign new_P2_U7423 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~P2_STATE2_REG_3_;
  assign new_P2_U7424 = ~new_P2_U2352 | ~new_P2_U7353;
  assign new_P2_U7425 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~P2_STATE2_REG_3_;
  assign new_P2_U7426 = ~new_P2_U2439 | ~new_P2_U3295;
  assign new_P2_U7427 = ~new_P2_U2352 | ~new_P2_U7387;
  assign new_P2_U7428 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~P2_STATE2_REG_3_;
  assign new_P2_U7429 = ~new_P2_U2352 | ~new_P2_U7421;
  assign new_P2_U7430 = ~P2_INSTQUEUEWR_ADDR_REG_0_ | ~P2_STATE2_REG_3_;
  assign new_P2_U7431 = ~new_P2_U2439 | ~new_P2_U3279;
  assign new_P2_U7432 = ~new_P2_U4413 | ~new_P2_U4414 | ~new_P2_U7431;
  assign new_P2_U7433 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_U7432;
  assign new_P2_U7434 = ~new_P2_U2353 | ~P2_REIP_REG_9_;
  assign new_P2_U7435 = ~new_P2_U4412 | ~P2_EAX_REG_9_;
  assign new_P2_U7436 = ~new_P2_U2352 | ~new_P2_U2608;
  assign new_P2_U7437 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_U7432;
  assign new_P2_U7438 = ~new_P2_U2353 | ~P2_REIP_REG_8_;
  assign new_P2_U7439 = ~new_P2_U4412 | ~P2_EAX_REG_8_;
  assign new_P2_U7440 = ~new_P2_U2352 | ~new_P2_U2607;
  assign new_P2_U7441 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_U7432;
  assign new_P2_U7442 = ~new_P2_U2353 | ~P2_REIP_REG_7_;
  assign new_P2_U7443 = ~new_P2_U4412 | ~P2_EAX_REG_7_;
  assign new_P2_U7444 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_U7432;
  assign new_P2_U7445 = ~new_P2_U2353 | ~P2_REIP_REG_6_;
  assign new_P2_U7446 = ~new_P2_U4412 | ~P2_EAX_REG_6_;
  assign new_P2_U7447 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_U7432;
  assign new_P2_U7448 = ~new_P2_U2353 | ~P2_REIP_REG_5_;
  assign new_P2_U7449 = ~new_P2_U4412 | ~P2_EAX_REG_5_;
  assign new_P2_U7450 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_U7432;
  assign new_P2_U7451 = ~new_P2_U2353 | ~P2_REIP_REG_4_;
  assign new_P2_U7452 = ~new_P2_U4412 | ~P2_EAX_REG_4_;
  assign new_P2_U7453 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_U7432;
  assign new_P2_U7454 = ~new_P2_U2353 | ~P2_REIP_REG_31_;
  assign new_P2_U7455 = ~new_P2_U4412 | ~P2_EAX_REG_31_;
  assign new_P2_U7456 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_U7432;
  assign new_P2_U7457 = ~new_P2_U2353 | ~P2_REIP_REG_30_;
  assign new_P2_U7458 = ~new_P2_U4412 | ~P2_EAX_REG_30_;
  assign new_P2_U7459 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_U7432;
  assign new_P2_U7460 = ~new_P2_U2353 | ~P2_REIP_REG_3_;
  assign new_P2_U7461 = ~new_P2_U4412 | ~P2_EAX_REG_3_;
  assign new_P2_U7462 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_U7432;
  assign new_P2_U7463 = ~new_P2_U2353 | ~P2_REIP_REG_29_;
  assign new_P2_U7464 = ~new_P2_U4412 | ~P2_EAX_REG_29_;
  assign new_P2_U7465 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_U7432;
  assign new_P2_U7466 = ~new_P2_U2353 | ~P2_REIP_REG_28_;
  assign new_P2_U7467 = ~new_P2_U4412 | ~P2_EAX_REG_28_;
  assign new_P2_U7468 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_U7432;
  assign new_P2_U7469 = ~new_P2_U2353 | ~P2_REIP_REG_27_;
  assign new_P2_U7470 = ~new_P2_U4412 | ~P2_EAX_REG_27_;
  assign new_P2_U7471 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_U7432;
  assign new_P2_U7472 = ~new_P2_U2353 | ~P2_REIP_REG_26_;
  assign new_P2_U7473 = ~new_P2_U4412 | ~P2_EAX_REG_26_;
  assign new_P2_U7474 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_U7432;
  assign new_P2_U7475 = ~new_P2_U2353 | ~P2_REIP_REG_25_;
  assign new_P2_U7476 = ~new_P2_U4412 | ~P2_EAX_REG_25_;
  assign new_P2_U7477 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_U7432;
  assign new_P2_U7478 = ~new_P2_U2353 | ~P2_REIP_REG_24_;
  assign new_P2_U7479 = ~new_P2_U4412 | ~P2_EAX_REG_24_;
  assign new_P2_U7480 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_U7432;
  assign new_P2_U7481 = ~new_P2_U2353 | ~P2_REIP_REG_23_;
  assign new_P2_U7482 = ~new_P2_U4412 | ~P2_EAX_REG_23_;
  assign new_P2_U7483 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_U7432;
  assign new_P2_U7484 = ~new_P2_U2353 | ~P2_REIP_REG_22_;
  assign new_P2_U7485 = ~new_P2_U4412 | ~P2_EAX_REG_22_;
  assign new_P2_U7486 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_U7432;
  assign new_P2_U7487 = ~new_P2_U2353 | ~P2_REIP_REG_21_;
  assign new_P2_U7488 = ~new_P2_U4412 | ~P2_EAX_REG_21_;
  assign new_P2_U7489 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_U7432;
  assign new_P2_U7490 = ~new_P2_U2353 | ~P2_REIP_REG_20_;
  assign new_P2_U7491 = ~new_P2_U4412 | ~P2_EAX_REG_20_;
  assign new_P2_U7492 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_U7432;
  assign new_P2_U7493 = ~new_P2_U2353 | ~P2_REIP_REG_2_;
  assign new_P2_U7494 = ~new_P2_U4412 | ~P2_EAX_REG_2_;
  assign new_P2_U7495 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_U7432;
  assign new_P2_U7496 = ~new_P2_U2353 | ~P2_REIP_REG_19_;
  assign new_P2_U7497 = ~new_P2_U4412 | ~P2_EAX_REG_19_;
  assign new_P2_U7498 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_U7432;
  assign new_P2_U7499 = ~new_P2_U2353 | ~P2_REIP_REG_18_;
  assign new_P2_U7500 = ~new_P2_U4412 | ~P2_EAX_REG_18_;
  assign new_P2_U7501 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_U7432;
  assign new_P2_U7502 = ~new_P2_U2353 | ~P2_REIP_REG_17_;
  assign new_P2_U7503 = ~new_P2_U4412 | ~P2_EAX_REG_17_;
  assign new_P2_U7504 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_U7432;
  assign new_P2_U7505 = ~new_P2_U2353 | ~P2_REIP_REG_16_;
  assign new_P2_U7506 = ~new_P2_U4412 | ~P2_EAX_REG_16_;
  assign new_P2_U7507 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_U7432;
  assign new_P2_U7508 = ~new_P2_U2353 | ~P2_REIP_REG_15_;
  assign new_P2_U7509 = ~new_P2_U4412 | ~P2_EAX_REG_15_;
  assign new_P2_U7510 = ~new_P2_U2352 | ~new_P2_U2614;
  assign new_P2_U7511 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_U7432;
  assign new_P2_U7512 = ~new_P2_U2353 | ~P2_REIP_REG_14_;
  assign new_P2_U7513 = ~new_P2_U4412 | ~P2_EAX_REG_14_;
  assign new_P2_U7514 = ~new_P2_U2352 | ~new_P2_U2613;
  assign new_P2_U7515 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_U7432;
  assign new_P2_U7516 = ~new_P2_U2353 | ~P2_REIP_REG_13_;
  assign new_P2_U7517 = ~new_P2_U4412 | ~P2_EAX_REG_13_;
  assign new_P2_U7518 = ~new_P2_U2352 | ~new_P2_U2612;
  assign new_P2_U7519 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_U7432;
  assign new_P2_U7520 = ~new_P2_U2353 | ~P2_REIP_REG_12_;
  assign new_P2_U7521 = ~new_P2_U4412 | ~P2_EAX_REG_12_;
  assign new_P2_U7522 = ~new_P2_U2352 | ~new_P2_U2611;
  assign new_P2_U7523 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_U7432;
  assign new_P2_U7524 = ~new_P2_U2353 | ~P2_REIP_REG_11_;
  assign new_P2_U7525 = ~new_P2_U4412 | ~P2_EAX_REG_11_;
  assign new_P2_U7526 = ~new_P2_U2352 | ~new_P2_U2610;
  assign new_P2_U7527 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_U7432;
  assign new_P2_U7528 = ~new_P2_U2353 | ~P2_REIP_REG_10_;
  assign new_P2_U7529 = ~new_P2_U4412 | ~P2_EAX_REG_10_;
  assign new_P2_U7530 = ~new_P2_U2352 | ~new_P2_U2609;
  assign new_P2_U7531 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_U7432;
  assign new_P2_U7532 = ~new_P2_U2353 | ~P2_REIP_REG_1_;
  assign new_P2_U7533 = ~new_P2_U4412 | ~P2_EAX_REG_1_;
  assign new_P2_U7534 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_U7432;
  assign new_P2_U7535 = ~new_P2_U2353 | ~P2_REIP_REG_0_;
  assign new_P2_U7536 = ~new_P2_U4412 | ~P2_EAX_REG_0_;
  assign new_P2_U7537 = ~P2_EBX_REG_9_ | ~new_P2_U7869;
  assign new_P2_U7538 = ~P2_EBX_REG_8_ | ~new_P2_U7869;
  assign new_P2_U7539 = ~P2_EBX_REG_31_ | ~new_P2_U7869;
  assign new_P2_U7540 = ~P2_EBX_REG_30_ | ~new_P2_U7869;
  assign new_P2_U7541 = ~P2_EBX_REG_29_ | ~new_P2_U7869;
  assign new_P2_U7542 = ~P2_EBX_REG_28_ | ~new_P2_U7869;
  assign new_P2_U7543 = ~P2_EBX_REG_27_ | ~new_P2_U7869;
  assign new_P2_U7544 = ~P2_EBX_REG_26_ | ~new_P2_U7869;
  assign new_P2_U7545 = ~P2_EBX_REG_25_ | ~new_P2_U7869;
  assign new_P2_U7546 = ~P2_EBX_REG_24_ | ~new_P2_U7869;
  assign new_P2_U7547 = ~P2_EBX_REG_23_ | ~new_P2_U7869;
  assign new_P2_U7548 = ~P2_EBX_REG_22_ | ~new_P2_U7869;
  assign new_P2_U7549 = ~P2_EBX_REG_21_ | ~new_P2_U7869;
  assign new_P2_U7550 = ~P2_EBX_REG_20_ | ~new_P2_U7869;
  assign new_P2_U7551 = ~P2_EBX_REG_19_ | ~new_P2_U7869;
  assign new_P2_U7552 = ~P2_EBX_REG_18_ | ~new_P2_U7869;
  assign new_P2_U7553 = ~P2_EBX_REG_17_ | ~new_P2_U7869;
  assign new_P2_U7554 = ~P2_EBX_REG_16_ | ~new_P2_U7869;
  assign new_P2_U7555 = ~P2_EBX_REG_15_ | ~new_P2_U7869;
  assign new_P2_U7556 = ~P2_EBX_REG_14_ | ~new_P2_U7869;
  assign new_P2_U7557 = ~P2_EBX_REG_13_ | ~new_P2_U7869;
  assign new_P2_U7558 = ~P2_EBX_REG_12_ | ~new_P2_U7869;
  assign new_P2_U7559 = ~P2_EBX_REG_11_ | ~new_P2_U7869;
  assign new_P2_U7560 = ~P2_EBX_REG_10_ | ~new_P2_U7869;
  assign new_P2_U7561 = ~new_P2_U4596 | ~new_P2_U3294;
  assign new_P2_U7562 = ~new_P2_U4428 | ~new_P2_U7285;
  assign new_P2_U7563 = ~P2_INSTQUEUERD_ADDR_REG_4_ | ~new_P2_U7561;
  assign new_P2_U7564 = ~new_P2_U4428 | ~new_P2_U7319;
  assign new_P2_U7565 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U7561;
  assign new_P2_U7566 = ~new_P2_U4428 | ~new_P2_U7353;
  assign new_P2_U7567 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U7561;
  assign new_P2_U7568 = ~new_P2_U4428 | ~new_P2_U7387;
  assign new_P2_U7569 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U7561;
  assign new_P2_U7570 = ~new_P2_U4428 | ~new_P2_U7421;
  assign new_P2_U7571 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_U7561;
  assign new_P2_U7572 = ~P2_INSTQUEUEWR_ADDR_REG_4_ | ~new_P2_U7561;
  assign new_P2_U7573 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_U7561;
  assign new_P2_U7574 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_U7561;
  assign new_P2_U7575 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_U7561;
  assign new_P2_U7576 = ~P2_INSTQUEUEWR_ADDR_REG_0_ | ~new_P2_U7561;
  assign new_P2_U7577 = ~new_P2_U4377 | ~new_P2_U5572;
  assign new_P2_U7578 = ~P2_STATE2_REG_0_ | ~new_P2_U4432;
  assign new_P2_U7579 = ~new_P2_U2617 | ~new_P2_U2450;
  assign new_P2_U7580 = ~new_P2_U4376 | ~new_P2_U5592;
  assign new_P2_U7581 = ~new_P2_U7867 | ~new_P2_U3525 | ~new_P2_U6845;
  assign new_P2_U7582 = ~new_P2_U4471 | ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_U7583 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U7890;
  assign new_P2_U7584 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U7890;
  assign new_P2_U7585 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_U3284;
  assign new_P2_U7586 = ~new_P2_U4381 | ~new_P2_U4424;
  assign new_P2_U7587 = ~new_P2_U4471 | ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_U7588 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U7890;
  assign new_P2_U7589 = ~new_P2_U2590 | ~new_P2_U6845;
  assign new_P2_U7590 = ~new_P2_U4471 | ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P2_U7591 = ~new_P2_U4416 | ~new_P2_U2376 | ~new_P2_U7871;
  assign new_P2_U7592 = ~new_P2_U3539 | ~new_P2_U4422 | ~new_P2_U7591 | ~new_P2_U3285;
  assign new_P2_U7593 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_U7592;
  assign new_P2_U7594 = ~P2_PHYADDRPOINTER_REG_9_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7595 = ~new_P2_U4423 | ~P2_REIP_REG_9_;
  assign new_P2_U7596 = ~new_P2_U2358 | ~P2_EBX_REG_9_;
  assign new_P2_U7597 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_U7592;
  assign new_P2_U7598 = ~P2_PHYADDRPOINTER_REG_8_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7599 = ~new_P2_U4423 | ~P2_REIP_REG_8_;
  assign new_P2_U7600 = ~new_P2_U2358 | ~P2_EBX_REG_8_;
  assign new_P2_U7601 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_U7592;
  assign new_P2_U7602 = ~P2_PHYADDRPOINTER_REG_7_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7603 = ~new_P2_U4423 | ~P2_REIP_REG_7_;
  assign new_P2_U7604 = ~new_P2_U2358 | ~P2_EBX_REG_7_;
  assign new_P2_U7605 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_U7592;
  assign new_P2_U7606 = ~P2_PHYADDRPOINTER_REG_6_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7607 = ~new_P2_U4423 | ~P2_REIP_REG_6_;
  assign new_P2_U7608 = ~new_P2_U2358 | ~P2_EBX_REG_6_;
  assign new_P2_U7609 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_U7592;
  assign new_P2_U7610 = ~P2_PHYADDRPOINTER_REG_5_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7611 = ~new_P2_U4423 | ~P2_REIP_REG_5_;
  assign new_P2_U7612 = ~new_P2_U2358 | ~P2_EBX_REG_5_;
  assign new_P2_U7613 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_U7592;
  assign new_P2_U7614 = ~P2_PHYADDRPOINTER_REG_4_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7615 = ~new_P2_U4423 | ~P2_REIP_REG_4_;
  assign new_P2_U7616 = ~new_P2_U2358 | ~P2_EBX_REG_4_;
  assign new_P2_U7617 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_U7592;
  assign new_P2_U7618 = ~P2_PHYADDRPOINTER_REG_31_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7619 = ~new_P2_U4423 | ~P2_REIP_REG_31_;
  assign new_P2_U7620 = ~new_P2_U2358 | ~P2_EBX_REG_31_;
  assign new_P2_U7621 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_U7592;
  assign new_P2_U7622 = ~P2_PHYADDRPOINTER_REG_30_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7623 = ~new_P2_U4423 | ~P2_REIP_REG_30_;
  assign new_P2_U7624 = ~new_P2_U2358 | ~P2_EBX_REG_30_;
  assign new_P2_U7625 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_U7592;
  assign new_P2_U7626 = ~P2_PHYADDRPOINTER_REG_3_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7627 = ~new_P2_U4423 | ~P2_REIP_REG_3_;
  assign new_P2_U7628 = ~new_P2_U2358 | ~P2_EBX_REG_3_;
  assign new_P2_U7629 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_U7592;
  assign new_P2_U7630 = ~P2_PHYADDRPOINTER_REG_29_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7631 = ~new_P2_U4423 | ~P2_REIP_REG_29_;
  assign new_P2_U7632 = ~new_P2_U2358 | ~P2_EBX_REG_29_;
  assign new_P2_U7633 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_U7592;
  assign new_P2_U7634 = ~P2_PHYADDRPOINTER_REG_28_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7635 = ~new_P2_U4423 | ~P2_REIP_REG_28_;
  assign new_P2_U7636 = ~new_P2_U2358 | ~P2_EBX_REG_28_;
  assign new_P2_U7637 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_U7592;
  assign new_P2_U7638 = ~P2_PHYADDRPOINTER_REG_27_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7639 = ~new_P2_U4423 | ~P2_REIP_REG_27_;
  assign new_P2_U7640 = ~new_P2_U2358 | ~P2_EBX_REG_27_;
  assign new_P2_U7641 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_U7592;
  assign new_P2_U7642 = ~P2_PHYADDRPOINTER_REG_26_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7643 = ~new_P2_U4423 | ~P2_REIP_REG_26_;
  assign new_P2_U7644 = ~new_P2_U2358 | ~P2_EBX_REG_26_;
  assign new_P2_U7645 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_U7592;
  assign new_P2_U7646 = ~P2_PHYADDRPOINTER_REG_25_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7647 = ~new_P2_U4423 | ~P2_REIP_REG_25_;
  assign new_P2_U7648 = ~new_P2_U2358 | ~P2_EBX_REG_25_;
  assign new_P2_U7649 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_U7592;
  assign new_P2_U7650 = ~P2_PHYADDRPOINTER_REG_24_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7651 = ~new_P2_U4423 | ~P2_REIP_REG_24_;
  assign new_P2_U7652 = ~new_P2_U2358 | ~P2_EBX_REG_24_;
  assign new_P2_U7653 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_U7592;
  assign new_P2_U7654 = ~P2_PHYADDRPOINTER_REG_23_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7655 = ~new_P2_U4423 | ~P2_REIP_REG_23_;
  assign new_P2_U7656 = ~new_P2_U2358 | ~P2_EBX_REG_23_;
  assign new_P2_U7657 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_U7592;
  assign new_P2_U7658 = ~P2_PHYADDRPOINTER_REG_22_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7659 = ~new_P2_U4423 | ~P2_REIP_REG_22_;
  assign new_P2_U7660 = ~new_P2_U2358 | ~P2_EBX_REG_22_;
  assign new_P2_U7661 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_U7592;
  assign new_P2_U7662 = ~P2_PHYADDRPOINTER_REG_21_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7663 = ~new_P2_U4423 | ~P2_REIP_REG_21_;
  assign new_P2_U7664 = ~new_P2_U2358 | ~P2_EBX_REG_21_;
  assign new_P2_U7665 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_U7592;
  assign new_P2_U7666 = ~P2_PHYADDRPOINTER_REG_20_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7667 = ~new_P2_U4423 | ~P2_REIP_REG_20_;
  assign new_P2_U7668 = ~new_P2_U2358 | ~P2_EBX_REG_20_;
  assign new_P2_U7669 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_U7592;
  assign new_P2_U7670 = ~P2_PHYADDRPOINTER_REG_2_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7671 = ~new_P2_U4423 | ~P2_REIP_REG_2_;
  assign new_P2_U7672 = ~new_P2_U2358 | ~P2_EBX_REG_2_;
  assign new_P2_U7673 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_U7592;
  assign new_P2_U7674 = ~P2_PHYADDRPOINTER_REG_19_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7675 = ~new_P2_U4423 | ~P2_REIP_REG_19_;
  assign new_P2_U7676 = ~new_P2_U2358 | ~P2_EBX_REG_19_;
  assign new_P2_U7677 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_U7592;
  assign new_P2_U7678 = ~P2_PHYADDRPOINTER_REG_18_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7679 = ~new_P2_U4423 | ~P2_REIP_REG_18_;
  assign new_P2_U7680 = ~new_P2_U2358 | ~P2_EBX_REG_18_;
  assign new_P2_U7681 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_U7592;
  assign new_P2_U7682 = ~P2_PHYADDRPOINTER_REG_17_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7683 = ~new_P2_U4423 | ~P2_REIP_REG_17_;
  assign new_P2_U7684 = ~new_P2_U2358 | ~P2_EBX_REG_17_;
  assign new_P2_U7685 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_U7592;
  assign new_P2_U7686 = ~P2_PHYADDRPOINTER_REG_16_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7687 = ~new_P2_U4423 | ~P2_REIP_REG_16_;
  assign new_P2_U7688 = ~new_P2_U2358 | ~P2_EBX_REG_16_;
  assign new_P2_U7689 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_U7592;
  assign new_P2_U7690 = ~P2_PHYADDRPOINTER_REG_15_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7691 = ~new_P2_U4423 | ~P2_REIP_REG_15_;
  assign new_P2_U7692 = ~new_P2_U2358 | ~P2_EBX_REG_15_;
  assign new_P2_U7693 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_U7592;
  assign new_P2_U7694 = ~P2_PHYADDRPOINTER_REG_14_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7695 = ~new_P2_U4423 | ~P2_REIP_REG_14_;
  assign new_P2_U7696 = ~new_P2_U2358 | ~P2_EBX_REG_14_;
  assign new_P2_U7697 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_U7592;
  assign new_P2_U7698 = ~P2_PHYADDRPOINTER_REG_13_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7699 = ~new_P2_U4423 | ~P2_REIP_REG_13_;
  assign new_P2_U7700 = ~new_P2_U2358 | ~P2_EBX_REG_13_;
  assign new_P2_U7701 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_U7592;
  assign new_P2_U7702 = ~P2_PHYADDRPOINTER_REG_12_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7703 = ~new_P2_U4423 | ~P2_REIP_REG_12_;
  assign new_P2_U7704 = ~new_P2_U2358 | ~P2_EBX_REG_12_;
  assign new_P2_U7705 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_U7592;
  assign new_P2_U7706 = ~P2_PHYADDRPOINTER_REG_11_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7707 = ~new_P2_U4423 | ~P2_REIP_REG_11_;
  assign new_P2_U7708 = ~new_P2_U2358 | ~P2_EBX_REG_11_;
  assign new_P2_U7709 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_U7592;
  assign new_P2_U7710 = ~P2_PHYADDRPOINTER_REG_10_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7711 = ~new_P2_U4423 | ~P2_REIP_REG_10_;
  assign new_P2_U7712 = ~new_P2_U2358 | ~P2_EBX_REG_10_;
  assign new_P2_U7713 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_U7592;
  assign new_P2_U7714 = ~P2_PHYADDRPOINTER_REG_1_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7715 = ~new_P2_U4423 | ~P2_REIP_REG_1_;
  assign new_P2_U7716 = ~new_P2_U2358 | ~P2_EBX_REG_1_;
  assign new_P2_U7717 = ~new_P2_U4387 | ~new_P2_U7885;
  assign new_P2_U7718 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_U7739;
  assign new_P2_U7719 = ~P2_PHYADDRPOINTER_REG_0_ | ~P2_STATE2_REG_1_;
  assign new_P2_U7720 = ~new_P2_U4423 | ~P2_REIP_REG_0_;
  assign new_P2_U7721 = ~new_P2_U2358 | ~P2_EBX_REG_0_;
  assign new_P2_U7722 = ~new_P2_U7720 | ~new_P2_U3575;
  assign new_P2_U7723 = ~new_P2_U3550 | ~new_P2_U3536;
  assign new_P2_U7724 = ~new_P2_R2219_U28 | ~new_P2_U7723;
  assign new_P2_U7725 = ~new_P2_R2219_U30 | ~new_P2_U7723;
  assign new_P2_U7726 = ~new_P2_R2238_U19 | ~new_P2_U2356;
  assign new_P2_U7727 = ~P2_INSTQUEUERD_ADDR_REG_4_ | ~new_P2_U3284;
  assign new_P2_U7728 = ~new_P2_R2238_U20 | ~new_P2_U2356;
  assign new_P2_U7729 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3284;
  assign new_P2_U7730 = ~new_P2_R2238_U21 | ~new_P2_U2356;
  assign new_P2_U7731 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U3284;
  assign new_P2_U7732 = ~new_P2_R2238_U22 | ~new_P2_U2356;
  assign new_P2_U7733 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U3284;
  assign new_P2_U7734 = ~new_P2_R2238_U7 | ~new_P2_U2356;
  assign new_P2_U7735 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_U3284;
  assign new_P2_U7736 = ~new_P2_U3525 | ~new_P2_U3295 | ~new_P2_U7873;
  assign new_P2_U7737 = ~new_P2_U3272 | ~new_P2_U4422 | ~new_P2_U7590 | ~new_P2_U7589;
  assign new_P2_U7738 = ~new_P2_U7861 | ~new_P2_U2617;
  assign new_P2_U7739 = ~new_P2_U3539 | ~new_P2_U4422 | ~new_P2_U7591 | ~new_P2_U3285;
  assign new_P2_U7740 = ~new_P2_U5571 | ~new_P2_U5573 | ~new_P2_U3521 | ~new_P2_U7744;
  assign new_P2_U7741 = ~new_P2_U2391 | ~new_P2_U3544;
  assign new_P2_U7742 = ~new_P2_U2377 | ~new_P2_U6572;
  assign new_P2_U7743 = ~new_P2_U7742 | ~new_P2_U7741 | ~new_P2_U4448;
  assign new_P2_U7744 = ~new_P2_U7745 | ~new_P2_U3278;
  assign new_P2_U7745 = ~new_P2_U7861 | ~new_P2_U2617;
  assign new_P2_U7746 = ~new_P2_U4592 | ~new_P2_U8003 | ~new_P2_U8002;
  assign new_P2_U7747 = ~new_P2_U4592 | ~new_P2_U7971 | ~new_P2_U7970;
  assign new_P2_U7748 = ~new_P2_U4592 | ~new_P2_U7955 | ~new_P2_U7954;
  assign new_P2_U7749 = ~new_P2_U4592 | ~new_P2_U8035 | ~new_P2_U8034;
  assign new_P2_U7750 = ~new_P2_U4592 | ~new_P2_U8019 | ~new_P2_U8018;
  assign new_P2_U7751 = ~new_P2_U4592 | ~new_P2_U7987 | ~new_P2_U7986;
  assign new_P2_U7752 = ~new_P2_U4592 | ~new_P2_U7939 | ~new_P2_U7938;
  assign new_P2_U7753 = ~new_P2_U4592 | ~new_P2_U7923 | ~new_P2_U7922;
  assign new_P2_U7754 = ~new_P2_U4592 | ~new_P2_U8154 | ~new_P2_U8153;
  assign new_P2_U7755 = ~new_P2_U4592 | ~new_P2_U8170 | ~new_P2_U8169;
  assign new_P2_U7756 = ~new_P2_U4592 | ~new_P2_U8186 | ~new_P2_U8185;
  assign new_P2_U7757 = ~new_P2_U4592 | ~new_P2_U8202 | ~new_P2_U8201;
  assign new_P2_U7758 = ~new_P2_U4592 | ~new_P2_U8218 | ~new_P2_U8217;
  assign new_P2_U7759 = ~new_P2_U4592 | ~new_P2_U8234 | ~new_P2_U8233;
  assign new_P2_U7760 = ~new_P2_U4592 | ~new_P2_U8250 | ~new_P2_U8249;
  assign new_P2_U7761 = ~new_P2_U4592 | ~new_P2_U8266 | ~new_P2_U8265;
  assign new_P2_U7762 = ~new_P2_U4593 | ~new_P2_U8005 | ~new_P2_U8004;
  assign new_P2_U7763 = ~new_P2_U4593 | ~new_P2_U7973 | ~new_P2_U7972;
  assign new_P2_U7764 = ~new_P2_U4593 | ~new_P2_U7957 | ~new_P2_U7956;
  assign new_P2_U7765 = ~new_P2_U4593 | ~new_P2_U8037 | ~new_P2_U8036;
  assign new_P2_U7766 = ~new_P2_U4593 | ~new_P2_U8021 | ~new_P2_U8020;
  assign new_P2_U7767 = ~new_P2_U4593 | ~new_P2_U7989 | ~new_P2_U7988;
  assign new_P2_U7768 = ~new_P2_U4593 | ~new_P2_U7941 | ~new_P2_U7940;
  assign new_P2_U7769 = ~new_P2_U4593 | ~new_P2_U7925 | ~new_P2_U7924;
  assign new_P2_U7770 = ~new_P2_U4593 | ~new_P2_U8156 | ~new_P2_U8155;
  assign new_P2_U7771 = ~new_P2_U4593 | ~new_P2_U8172 | ~new_P2_U8171;
  assign new_P2_U7772 = ~new_P2_U4593 | ~new_P2_U8188 | ~new_P2_U8187;
  assign new_P2_U7773 = ~new_P2_U4593 | ~new_P2_U8204 | ~new_P2_U8203;
  assign new_P2_U7774 = ~new_P2_U4593 | ~new_P2_U8220 | ~new_P2_U8219;
  assign new_P2_U7775 = ~new_P2_U4593 | ~new_P2_U8236 | ~new_P2_U8235;
  assign new_P2_U7776 = ~new_P2_U4593 | ~new_P2_U8252 | ~new_P2_U8251;
  assign new_P2_U7777 = ~new_P2_U4593 | ~new_P2_U8268 | ~new_P2_U8267;
  assign new_P2_U7778 = ~new_P2_U2456 | ~new_P2_U8007 | ~new_P2_U8006;
  assign new_P2_U7779 = ~new_P2_U2456 | ~new_P2_U7975 | ~new_P2_U7974;
  assign new_P2_U7780 = ~new_P2_U2456 | ~new_P2_U7959 | ~new_P2_U7958;
  assign new_P2_U7781 = ~new_P2_U2456 | ~new_P2_U8039 | ~new_P2_U8038;
  assign new_P2_U7782 = ~new_P2_U2456 | ~new_P2_U8023 | ~new_P2_U8022;
  assign new_P2_U7783 = ~new_P2_U2456 | ~new_P2_U7991 | ~new_P2_U7990;
  assign new_P2_U7784 = ~new_P2_U2456 | ~new_P2_U7943 | ~new_P2_U7942;
  assign new_P2_U7785 = ~new_P2_U2456 | ~new_P2_U7927 | ~new_P2_U7926;
  assign new_P2_U7786 = ~new_P2_U2456 | ~new_P2_U8158 | ~new_P2_U8157;
  assign new_P2_U7787 = ~new_P2_U2456 | ~new_P2_U8174 | ~new_P2_U8173;
  assign new_P2_U7788 = ~new_P2_U2456 | ~new_P2_U8190 | ~new_P2_U8189;
  assign new_P2_U7789 = ~new_P2_U2456 | ~new_P2_U8206 | ~new_P2_U8205;
  assign new_P2_U7790 = ~new_P2_U2456 | ~new_P2_U8222 | ~new_P2_U8221;
  assign new_P2_U7791 = ~new_P2_U2456 | ~new_P2_U8238 | ~new_P2_U8237;
  assign new_P2_U7792 = ~new_P2_U2456 | ~new_P2_U8254 | ~new_P2_U8253;
  assign new_P2_U7793 = ~new_P2_U2456 | ~new_P2_U8270 | ~new_P2_U8269;
  assign new_P2_U7794 = ~new_P2_U2454 | ~new_P2_U8009 | ~new_P2_U8008;
  assign new_P2_U7795 = ~new_P2_U2454 | ~new_P2_U7977 | ~new_P2_U7976;
  assign new_P2_U7796 = ~new_P2_U2454 | ~new_P2_U7961 | ~new_P2_U7960;
  assign new_P2_U7797 = ~new_P2_U2454 | ~new_P2_U8041 | ~new_P2_U8040;
  assign new_P2_U7798 = ~new_P2_U2454 | ~new_P2_U8025 | ~new_P2_U8024;
  assign new_P2_U7799 = ~new_P2_U2454 | ~new_P2_U7993 | ~new_P2_U7992;
  assign new_P2_U7800 = ~new_P2_U2454 | ~new_P2_U7945 | ~new_P2_U7944;
  assign new_P2_U7801 = ~new_P2_U2454 | ~new_P2_U7929 | ~new_P2_U7928;
  assign new_P2_U7802 = ~new_P2_U2454 | ~new_P2_U8160 | ~new_P2_U8159;
  assign new_P2_U7803 = ~new_P2_U2454 | ~new_P2_U8176 | ~new_P2_U8175;
  assign new_P2_U7804 = ~new_P2_U2454 | ~new_P2_U8192 | ~new_P2_U8191;
  assign new_P2_U7805 = ~new_P2_U2454 | ~new_P2_U8208 | ~new_P2_U8207;
  assign new_P2_U7806 = ~new_P2_U2454 | ~new_P2_U8224 | ~new_P2_U8223;
  assign new_P2_U7807 = ~new_P2_U2454 | ~new_P2_U8240 | ~new_P2_U8239;
  assign new_P2_U7808 = ~new_P2_U2454 | ~new_P2_U8256 | ~new_P2_U8255;
  assign new_P2_U7809 = ~new_P2_U2454 | ~new_P2_U8272 | ~new_P2_U8271;
  assign new_P2_U7810 = ~new_P2_U4590 | ~new_P2_U8011 | ~new_P2_U8010;
  assign new_P2_U7811 = ~new_P2_U4590 | ~new_P2_U7979 | ~new_P2_U7978;
  assign new_P2_U7812 = ~new_P2_U4590 | ~new_P2_U7963 | ~new_P2_U7962;
  assign new_P2_U7813 = ~new_P2_U4590 | ~new_P2_U8043 | ~new_P2_U8042;
  assign new_P2_U7814 = ~new_P2_U4590 | ~new_P2_U8027 | ~new_P2_U8026;
  assign new_P2_U7815 = ~new_P2_U4590 | ~new_P2_U7995 | ~new_P2_U7994;
  assign new_P2_U7816 = ~new_P2_U4590 | ~new_P2_U7947 | ~new_P2_U7946;
  assign new_P2_U7817 = ~new_P2_U4590 | ~new_P2_U7931 | ~new_P2_U7930;
  assign new_P2_U7818 = ~new_P2_U4590 | ~new_P2_U8162 | ~new_P2_U8161;
  assign new_P2_U7819 = ~new_P2_U4590 | ~new_P2_U8178 | ~new_P2_U8177;
  assign new_P2_U7820 = ~new_P2_U4590 | ~new_P2_U8194 | ~new_P2_U8193;
  assign new_P2_U7821 = ~new_P2_U4590 | ~new_P2_U8210 | ~new_P2_U8209;
  assign new_P2_U7822 = ~new_P2_U4590 | ~new_P2_U8226 | ~new_P2_U8225;
  assign new_P2_U7823 = ~new_P2_U4590 | ~new_P2_U8242 | ~new_P2_U8241;
  assign new_P2_U7824 = ~new_P2_U4590 | ~new_P2_U8258 | ~new_P2_U8257;
  assign new_P2_U7825 = ~new_P2_U4590 | ~new_P2_U8274 | ~new_P2_U8273;
  assign new_P2_U7826 = ~new_P2_U2453 | ~new_P2_U8013 | ~new_P2_U8012;
  assign new_P2_U7827 = ~new_P2_U2453 | ~new_P2_U7981 | ~new_P2_U7980;
  assign new_P2_U7828 = ~new_P2_U2453 | ~new_P2_U7965 | ~new_P2_U7964;
  assign new_P2_U7829 = ~new_P2_U2453 | ~new_P2_U8045 | ~new_P2_U8044;
  assign new_P2_U7830 = ~new_P2_U2453 | ~new_P2_U8029 | ~new_P2_U8028;
  assign new_P2_U7831 = ~new_P2_U2453 | ~new_P2_U7997 | ~new_P2_U7996;
  assign new_P2_U7832 = ~new_P2_U2453 | ~new_P2_U7949 | ~new_P2_U7948;
  assign new_P2_U7833 = ~new_P2_U2453 | ~new_P2_U7933 | ~new_P2_U7932;
  assign new_P2_U7834 = ~new_P2_U2453 | ~new_P2_U8164 | ~new_P2_U8163;
  assign new_P2_U7835 = ~new_P2_U2453 | ~new_P2_U8180 | ~new_P2_U8179;
  assign new_P2_U7836 = ~new_P2_U2453 | ~new_P2_U8196 | ~new_P2_U8195;
  assign new_P2_U7837 = ~new_P2_U2453 | ~new_P2_U8212 | ~new_P2_U8211;
  assign new_P2_U7838 = ~new_P2_U2453 | ~new_P2_U8228 | ~new_P2_U8227;
  assign new_P2_U7839 = ~new_P2_U2453 | ~new_P2_U8244 | ~new_P2_U8243;
  assign new_P2_U7840 = ~new_P2_U2453 | ~new_P2_U8260 | ~new_P2_U8259;
  assign new_P2_U7841 = ~new_P2_U2453 | ~new_P2_U8276 | ~new_P2_U8275;
  assign new_P2_U7842 = ~new_P2_U2452 | ~new_P2_U8015 | ~new_P2_U8014;
  assign new_P2_U7843 = ~new_P2_U2452 | ~new_P2_U7983 | ~new_P2_U7982;
  assign new_P2_U7844 = ~new_P2_U2452 | ~new_P2_U7967 | ~new_P2_U7966;
  assign new_P2_U7845 = ~new_P2_U2452 | ~new_P2_U8047 | ~new_P2_U8046;
  assign new_P2_U7846 = ~new_P2_U2452 | ~new_P2_U8031 | ~new_P2_U8030;
  assign new_P2_U7847 = ~new_P2_U2452 | ~new_P2_U7999 | ~new_P2_U7998;
  assign new_P2_U7848 = ~new_P2_U2452 | ~new_P2_U7951 | ~new_P2_U7950;
  assign new_P2_U7849 = ~new_P2_U2452 | ~new_P2_U7935 | ~new_P2_U7934;
  assign new_P2_U7850 = ~new_P2_U2452 | ~new_P2_U8166 | ~new_P2_U8165;
  assign new_P2_U7851 = ~new_P2_U2452 | ~new_P2_U8182 | ~new_P2_U8181;
  assign new_P2_U7852 = ~new_P2_U2452 | ~new_P2_U8198 | ~new_P2_U8197;
  assign new_P2_U7853 = ~new_P2_U2452 | ~new_P2_U8214 | ~new_P2_U8213;
  assign new_P2_U7854 = ~new_P2_U2452 | ~new_P2_U8230 | ~new_P2_U8229;
  assign new_P2_U7855 = ~new_P2_U2452 | ~new_P2_U8246 | ~new_P2_U8245;
  assign new_P2_U7856 = ~new_P2_U2452 | ~new_P2_U8262 | ~new_P2_U8261;
  assign new_P2_U7857 = ~new_P2_U2452 | ~new_P2_U8278 | ~new_P2_U8277;
  assign new_P2_U7858 = ~new_P2_U2455 | ~new_P2_U8017 | ~new_P2_U8016;
  assign new_P2_U7859 = ~new_P2_U3280;
  assign new_P2_U7860 = ~new_P2_U2455 | ~new_P2_U7985 | ~new_P2_U7984;
  assign new_P2_U7861 = ~new_P2_U3279;
  assign new_P2_U7862 = ~new_P2_U2455 | ~new_P2_U7969 | ~new_P2_U7968;
  assign new_P2_U7863 = ~new_P2_U3278;
  assign new_P2_U7864 = ~new_P2_U2455 | ~new_P2_U8049 | ~new_P2_U8048;
  assign new_P2_U7865 = ~new_P2_U3521;
  assign new_P2_U7866 = ~new_P2_U2455 | ~new_P2_U8033 | ~new_P2_U8032;
  assign new_P2_U7867 = ~new_P2_U3255;
  assign new_P2_U7868 = ~new_P2_U2455 | ~new_P2_U8001 | ~new_P2_U8000;
  assign new_P2_U7869 = ~new_P2_U2617;
  assign new_P2_U7870 = ~new_P2_U2455 | ~new_P2_U7953 | ~new_P2_U7952;
  assign new_P2_U7871 = ~new_P2_U3253;
  assign new_P2_U7872 = ~new_P2_U2455 | ~new_P2_U7937 | ~new_P2_U7936;
  assign new_P2_U7873 = ~new_P2_U2616;
  assign new_P2_U7874 = ~new_P2_U2455 | ~new_P2_U8168 | ~new_P2_U8167;
  assign new_P2_U7875 = ~new_P2_U2455 | ~new_P2_U8184 | ~new_P2_U8183;
  assign new_P2_U7876 = ~new_P2_U2455 | ~new_P2_U8200 | ~new_P2_U8199;
  assign new_P2_U7877 = ~new_P2_U2455 | ~new_P2_U8216 | ~new_P2_U8215;
  assign new_P2_U7878 = ~new_P2_U2455 | ~new_P2_U8232 | ~new_P2_U8231;
  assign new_P2_U7879 = ~new_P2_U2455 | ~new_P2_U8248 | ~new_P2_U8247;
  assign new_P2_U7880 = ~new_P2_U2455 | ~new_P2_U8264 | ~new_P2_U8263;
  assign new_P2_U7881 = ~new_P2_U2455 | ~new_P2_U8280 | ~new_P2_U8279;
  assign new_P2_U7882 = ~new_P2_U5590 | ~new_P2_U4428;
  assign new_P2_U7883 = ~new_P2_U5596 | ~new_P2_U3525;
  assign new_P2_U7884 = ~new_P2_U4596 | ~new_P2_U7883;
  assign new_P2_U7885 = ~new_P2_U3253 | ~new_P2_U8348 | ~new_P2_U8347;
  assign new_P2_U7886 = ~new_P2_U7722 | ~new_P2_U5589;
  assign new_P2_U7887 = ~new_P2_U4459 | ~new_P2_U5589;
  assign new_P2_U7888 = ~new_P2_U4384 | ~new_P2_U4385 | ~new_P2_U2589 | ~new_P2_U4386 | ~new_P2_U7887;
  assign new_P2_U7889 = ~new_P2_U4459 | ~new_P2_U5589;
  assign new_P2_U7890 = ~new_P2_U4379 | ~new_P2_U2589 | ~new_P2_U7889 | ~new_P2_U4458;
  assign new_P2_U7891 = ~new_P2_U4569 | ~new_P2_U4572 | ~P2_STATE_REG_1_;
  assign new_P2_U7892 = ~P2_STATE_REG_0_ | ~P2_REQUESTPENDING_REG | ~new_P2_U3244;
  assign new_P2_U7893 = ~P2_STATE_REG_1_ | ~new_P2_U4569;
  assign new_P2_U7894 = ~new_P2_U4600 | ~new_P2_U4615;
  assign new_P2_U7895 = ~new_P2_U7863 | ~new_P2_U7871;
  assign new_P2_U7896 = ~new_P2_U3255 | ~new_P2_U5595;
  assign new_P2_U7897 = ~new_P2_U4429 | ~new_P2_U5589;
  assign new_P2_U7898 = ~P2_REIP_REG_0_ | ~P2_DATAWIDTH_REG_0_;
  assign new_P2_U7899 = ~P2_BE_N_REG_3_ | ~new_P2_U3259;
  assign new_P2_U7900 = ~P2_BYTEENABLE_REG_3_ | ~new_P2_U4439;
  assign new_P2_U7901 = ~P2_BE_N_REG_2_ | ~new_P2_U3259;
  assign new_P2_U7902 = ~P2_BYTEENABLE_REG_2_ | ~new_P2_U4439;
  assign new_P2_U7903 = ~P2_BE_N_REG_1_ | ~new_P2_U3259;
  assign new_P2_U7904 = ~P2_BYTEENABLE_REG_1_ | ~new_P2_U4439;
  assign new_P2_U7905 = ~P2_BE_N_REG_0_ | ~new_P2_U3259;
  assign new_P2_U7906 = ~P2_BYTEENABLE_REG_0_ | ~new_P2_U4439;
  assign new_P2_U7907 = ~P2_STATE_REG_0_ | ~new_P2_U3268 | ~new_P2_U3267;
  assign new_P2_U7908 = NA | P2_STATE_REG_0_;
  assign new_P2_U7909 = ~P2_STATE_REG_2_ | ~new_P2_U3266;
  assign new_P2_U7910 = ~new_P2_U4568 | ~P2_STATE_REG_0_;
  assign new_P2_U7911 = ~P2_STATE_REG_1_ | ~new_P2_U4581 | ~new_P2_U4572;
  assign new_P2_U7912 = ~new_P2_U4582 | ~new_P2_U3258;
  assign new_P2_U7913 = ~P2_STATE_REG_2_ | ~P2_STATE_REG_0_ | ~new_P2_U3267;
  assign new_P2_U7914 = ~new_P2_U4584 | ~new_P2_U3244;
  assign new_P2_U7915 = P2_STATE_REG_0_ | P2_STATE_REG_1_;
  assign new_P2_U7916 = ~P2_STATE_REG_0_ | ~new_P2_U4473;
  assign new_P2_U7917 = ~new_P2_U3589;
  assign new_P2_U7918 = ~new_P2_U7917 | ~P2_DATAWIDTH_REG_0_;
  assign new_P2_U7919 = ~new_P2_U3590 | ~new_P2_U3589;
  assign new_P2_U7920 = ~new_P2_U3589 | ~new_P2_U4589;
  assign new_P2_U7921 = ~new_P2_U7917 | ~P2_DATAWIDTH_REG_1_;
  assign new_P2_U7922 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3388;
  assign new_P2_U7923 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__1_;
  assign new_P2_U7924 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__1_;
  assign new_P2_U7925 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3422;
  assign new_P2_U7926 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__1_;
  assign new_P2_U7927 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3411;
  assign new_P2_U7928 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3374;
  assign new_P2_U7929 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__1_;
  assign new_P2_U7930 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3333;
  assign new_P2_U7931 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__1_;
  assign new_P2_U7932 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3363;
  assign new_P2_U7933 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__1_;
  assign new_P2_U7934 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3347;
  assign new_P2_U7935 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__1_;
  assign new_P2_U7936 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3399;
  assign new_P2_U7937 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__1_;
  assign new_P2_U7938 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3389;
  assign new_P2_U7939 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__0_;
  assign new_P2_U7940 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__0_;
  assign new_P2_U7941 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3423;
  assign new_P2_U7942 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__0_;
  assign new_P2_U7943 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3412;
  assign new_P2_U7944 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3375;
  assign new_P2_U7945 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__0_;
  assign new_P2_U7946 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3334;
  assign new_P2_U7947 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__0_;
  assign new_P2_U7948 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3364;
  assign new_P2_U7949 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__0_;
  assign new_P2_U7950 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3348;
  assign new_P2_U7951 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__0_;
  assign new_P2_U7952 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3400;
  assign new_P2_U7953 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__0_;
  assign new_P2_U7954 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3385;
  assign new_P2_U7955 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__4_;
  assign new_P2_U7956 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__4_;
  assign new_P2_U7957 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3419;
  assign new_P2_U7958 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__4_;
  assign new_P2_U7959 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3408;
  assign new_P2_U7960 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3371;
  assign new_P2_U7961 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__4_;
  assign new_P2_U7962 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3330;
  assign new_P2_U7963 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__4_;
  assign new_P2_U7964 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3360;
  assign new_P2_U7965 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__4_;
  assign new_P2_U7966 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3344;
  assign new_P2_U7967 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__4_;
  assign new_P2_U7968 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3396;
  assign new_P2_U7969 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__4_;
  assign new_P2_U7970 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3383;
  assign new_P2_U7971 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__6_;
  assign new_P2_U7972 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__6_;
  assign new_P2_U7973 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3417;
  assign new_P2_U7974 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__6_;
  assign new_P2_U7975 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3406;
  assign new_P2_U7976 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3369;
  assign new_P2_U7977 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__6_;
  assign new_P2_U7978 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3328;
  assign new_P2_U7979 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__6_;
  assign new_P2_U7980 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3358;
  assign new_P2_U7981 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__6_;
  assign new_P2_U7982 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3342;
  assign new_P2_U7983 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__6_;
  assign new_P2_U7984 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3394;
  assign new_P2_U7985 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__6_;
  assign new_P2_U7986 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3384;
  assign new_P2_U7987 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__5_;
  assign new_P2_U7988 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__5_;
  assign new_P2_U7989 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3418;
  assign new_P2_U7990 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__5_;
  assign new_P2_U7991 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3407;
  assign new_P2_U7992 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3370;
  assign new_P2_U7993 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__5_;
  assign new_P2_U7994 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3329;
  assign new_P2_U7995 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__5_;
  assign new_P2_U7996 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3359;
  assign new_P2_U7997 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__5_;
  assign new_P2_U7998 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3343;
  assign new_P2_U7999 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__5_;
  assign new_P2_U8000 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3395;
  assign new_P2_U8001 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__5_;
  assign new_P2_U8002 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3387;
  assign new_P2_U8003 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__2_;
  assign new_P2_U8004 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__2_;
  assign new_P2_U8005 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3421;
  assign new_P2_U8006 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__2_;
  assign new_P2_U8007 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3410;
  assign new_P2_U8008 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3373;
  assign new_P2_U8009 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__2_;
  assign new_P2_U8010 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3332;
  assign new_P2_U8011 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__2_;
  assign new_P2_U8012 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3362;
  assign new_P2_U8013 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__2_;
  assign new_P2_U8014 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3346;
  assign new_P2_U8015 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__2_;
  assign new_P2_U8016 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3398;
  assign new_P2_U8017 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__2_;
  assign new_P2_U8018 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3386;
  assign new_P2_U8019 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__3_;
  assign new_P2_U8020 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__3_;
  assign new_P2_U8021 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3420;
  assign new_P2_U8022 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__3_;
  assign new_P2_U8023 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3409;
  assign new_P2_U8024 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3372;
  assign new_P2_U8025 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__3_;
  assign new_P2_U8026 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3331;
  assign new_P2_U8027 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__3_;
  assign new_P2_U8028 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3361;
  assign new_P2_U8029 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__3_;
  assign new_P2_U8030 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3345;
  assign new_P2_U8031 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__3_;
  assign new_P2_U8032 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3397;
  assign new_P2_U8033 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__3_;
  assign new_P2_U8034 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3382;
  assign new_P2_U8035 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_3__7_;
  assign new_P2_U8036 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_0__7_;
  assign new_P2_U8037 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3416;
  assign new_P2_U8038 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_1__7_;
  assign new_P2_U8039 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3405;
  assign new_P2_U8040 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3368;
  assign new_P2_U8041 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_4__7_;
  assign new_P2_U8042 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3327;
  assign new_P2_U8043 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_7__7_;
  assign new_P2_U8044 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3357;
  assign new_P2_U8045 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_5__7_;
  assign new_P2_U8046 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3341;
  assign new_P2_U8047 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_6__7_;
  assign new_P2_U8048 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3393;
  assign new_P2_U8049 = P2_INSTQUEUERD_ADDR_REG_3_ | P2_INSTQUEUE_REG_2__7_;
  assign new_P2_U8050 = ~new_P2_R2167_U6 | ~new_P2_U4435;
  assign new_P2_U8051 = ~new_P2_U4604 | ~new_P2_U3297;
  assign new_P2_U8052 = ~new_P2_U7871 | ~new_P2_U3293;
  assign new_P2_U8053 = ~new_P2_U3253 | ~new_P2_U3282;
  assign new_P2_U8054 = ~new_P2_U4427 | ~new_P2_U3297;
  assign new_P2_U8055 = ~new_P2_U3289 | ~new_P2_U3520;
  assign new_P2_U8056 = new_U211 | P2_STATE2_REG_0_;
  assign new_P2_U8057 = ~P2_STATE2_REG_0_ | ~new_P2_U4617;
  assign new_P2_U8058 = ~P2_STATE2_REG_3_ | ~new_P2_U3299;
  assign new_P2_U8059 = ~new_P2_U2448 | ~new_P2_U4620;
  assign new_P2_U8060 = ~P2_STATE2_REG_0_ | ~new_P2_U4631;
  assign new_P2_U8061 = ~new_P2_U3284 | ~new_P2_U4630 | ~new_P2_U4619;
  assign new_P2_U8062 = ~new_P2_R2182_U40 | ~new_P2_U3318;
  assign new_P2_U8063 = ~new_P2_U4637 | ~new_P2_U3316;
  assign new_P2_U8064 = ~new_P2_U3579;
  assign new_P2_U8065 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_U3311;
  assign new_P2_U8066 = ~new_P2_U4642 | ~new_P2_U3310;
  assign new_P2_U8067 = ~new_P2_U3580;
  assign new_P2_U8068 = ~new_P2_U7859 | ~new_P2_U5574;
  assign new_P2_U8069 = ~new_P2_U3280 | ~new_P2_U5575;
  assign new_P2_U8070 = ~new_P2_U4435 | ~new_P2_U3297;
  assign new_P2_U8071 = ~new_P2_R2167_U6 | ~new_P2_U4433 | ~new_P2_U2359;
  assign new_P2_U8072 = ~new_P2_U3594 | ~new_P2_U4394;
  assign new_P2_U8073 = ~new_P2_U5584 | ~P2_INSTQUEUERD_ADDR_REG_4_;
  assign new_P2_U8074 = ~new_P2_U3280 | ~new_P2_U5586;
  assign new_P2_U8075 = ~new_P2_U7859 | ~new_P2_U2617 | ~new_P2_U3279;
  assign new_P2_U8076 = ~new_P2_U4424 | ~new_P2_U3253;
  assign new_P2_U8077 = ~new_P2_U4475 | ~new_P2_U7871;
  assign new_P2_U8078 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U5585;
  assign new_P2_U8079 = ~new_P2_U3273 | ~new_P2_U4591 | ~new_P2_U3276;
  assign new_P2_U8080 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3277;
  assign new_P2_U8081 = ~new_P2_U4590 | ~new_P2_U3273;
  assign new_P2_U8082 = ~new_P2_U3581;
  assign new_P2_U8083 = ~new_P2_U5584 | ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign new_P2_U8084 = ~new_P2_U5614 | ~new_P2_U4394;
  assign new_P2_U8085 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_U3528;
  assign new_P2_U8086 = ~new_P2_U3647 | ~new_P2_U3683;
  assign new_P2_U8087 = ~new_P2_U3597;
  assign new_P2_U8088 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_U3528;
  assign new_P2_U8089 = ~new_P2_R1957_U49 | ~new_P2_U3647;
  assign new_P2_U8090 = ~new_P2_U3598;
  assign new_P2_U8091 = ~new_P2_U5616 | ~new_P2_U5605;
  assign new_P2_U8092 = ~new_P2_U3530 | ~new_P2_U5606;
  assign new_P2_U8093 = ~new_P2_U5584 | ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign new_P2_U8094 = ~new_P2_U5623 | ~new_P2_U4394;
  assign new_P2_U8095 = ~new_P2_U3255 | ~new_P2_U3886 | ~new_P2_U4597;
  assign new_P2_U8096 = ~new_P2_U7867 | ~new_P2_U7869 | ~new_P2_U5625;
  assign new_P2_U8097 = ~new_P2_U8096 | ~new_P2_U8095;
  assign new_P2_U8098 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_U3271;
  assign new_P2_U8099 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U3272;
  assign new_P2_U8100 = ~new_P2_U3582;
  assign new_P2_U8101 = ~new_P2_U5584 | ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U8102 = ~new_P2_U5633 | ~new_P2_U4394;
  assign new_P2_U8103 = ~new_P2_U5584 | ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_U8104 = ~new_P2_U5641 | ~new_P2_U4394;
  assign new_P2_U8105 = ~new_P2_U5643 | ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_U8106 = ~new_P2_U5651 | ~new_P2_U3533;
  assign new_P2_U8107 = ~new_P2_U8064 | ~new_P2_U4636;
  assign new_P2_U8108 = ~new_P2_U3579 | ~new_P2_U3319;
  assign new_P2_U8109 = ~new_P2_U8108 | ~new_P2_U8107;
  assign new_P2_U8110 = ~new_P2_U5643 | ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P2_U8111 = ~new_P2_U5655 | ~new_P2_U3533;
  assign new_P2_U8112 = ~new_P2_U5643 | ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_U8113 = ~new_P2_U5660 | ~new_P2_U3533;
  assign new_P2_U8114 = ~new_P2_U5643 | ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P2_U8115 = ~new_P2_U5664 | ~new_P2_U3533;
  assign new_P2_U8116 = ~new_P2_U2616 | ~new_P2_U2359 | ~new_P2_U3280;
  assign new_P2_U8117 = ~new_P2_U2438 | ~new_P2_U7873;
  assign new_P2_U8118 = ~new_P2_U8117 | ~new_P2_U8116;
  assign new_P2_U8119 = ~new_P2_U3297 | ~new_P2_U3253 | ~new_P2_U3278;
  assign new_P2_U8120 = ~new_P2_U8118 | ~new_P2_R2167_U6;
  assign new_P2_U8121 = ~new_P2_U7859 | ~new_P2_U7873;
  assign new_P2_U8122 = ~new_P2_U2616 | ~new_P2_U3282;
  assign new_P2_U8123 = ~P2_BYTEENABLE_REG_3_ | ~new_P2_U3547;
  assign new_P2_U8124 = ~new_P2_U3606 | ~new_P2_U4438;
  assign new_P2_U8125 = ~P2_BYTEENABLE_REG_2_ | ~new_P2_U3547;
  assign new_P2_U8126 = ~new_P2_U3607 | ~new_P2_U4438;
  assign new_P2_U8127 = ~P2_BYTEENABLE_REG_0_ | ~new_P2_U3547;
  assign new_P2_U8128 = ~new_P2_U4438 | ~P2_REIP_REG_0_;
  assign new_P2_U8129 = ~new_P2_U4439 | ~new_P2_U3552;
  assign new_P2_U8130 = ~P2_W_R_N_REG | ~new_P2_U3259;
  assign new_P2_U8131 = ~new_P2_U3287 | ~new_P2_U7873;
  assign new_P2_U8132 = ~new_P2_R2243_U8 | ~new_P2_U2616;
  assign new_P2_U8133 = ~new_P2_U6838 | ~new_P2_U3257;
  assign new_P2_U8134 = ~P2_MORE_REG | ~new_P2_U4400;
  assign new_P2_U8135 = ~new_P2_U7917 | ~P2_STATEBS16_REG;
  assign new_P2_U8136 = ~BS16 | ~new_P2_U3589;
  assign new_P2_U8137 = ~new_P2_U6843 | ~P2_REQUESTPENDING_REG;
  assign new_P2_U8138 = ~new_P2_U6852 | ~new_P2_U4402;
  assign new_P2_U8139 = ~new_P2_U4439 | ~new_P2_U3551;
  assign new_P2_U8140 = ~P2_D_C_N_REG | ~new_P2_U3259;
  assign new_P2_U8141 = ~P2_M_IO_N_REG | ~new_P2_U3259;
  assign new_P2_U8142 = ~P2_MEMORYFETCH_REG | ~new_P2_U4439;
  assign new_P2_U8143 = ~new_P2_U6857 | ~P2_READREQUEST_REG;
  assign new_P2_U8144 = ~new_P2_U6858 | ~new_P2_U4403;
  assign new_P2_U8145 = ~new_P2_U7873 | ~new_P2_U3520;
  assign new_P2_U8146 = ~new_P2_U2616 | ~new_P2_U3297;
  assign new_P2_U8147 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U4405;
  assign new_P2_U8148 = ~new_P2_U7007 | ~new_P2_U3273;
  assign new_P2_U8149 = ~new_P2_U3583;
  assign new_P2_U8150 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U3273;
  assign new_P2_U8151 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_U3276;
  assign new_P2_U8152 = ~new_P2_U3584;
  assign new_P2_U8153 = ~new_P2_U3584 | ~new_P2_U3327;
  assign new_P2_U8154 = ~new_P2_U8152 | ~new_P2_U3431;
  assign new_P2_U8155 = ~new_P2_U3584 | ~new_P2_U3368;
  assign new_P2_U8156 = ~new_P2_U8152 | ~new_P2_U3465;
  assign new_P2_U8157 = ~new_P2_U3584 | ~new_P2_U3357;
  assign new_P2_U8158 = ~new_P2_U8152 | ~new_P2_U3454;
  assign new_P2_U8159 = ~new_P2_U3584 | ~new_P2_U3416;
  assign new_P2_U8160 = ~new_P2_U8152 | ~new_P2_U3511;
  assign new_P2_U8161 = ~new_P2_U3584 | ~new_P2_U3382;
  assign new_P2_U8162 = ~new_P2_U8152 | ~new_P2_U3477;
  assign new_P2_U8163 = ~new_P2_U3584 | ~new_P2_U3405;
  assign new_P2_U8164 = ~new_P2_U8152 | ~new_P2_U3500;
  assign new_P2_U8165 = ~new_P2_U3584 | ~new_P2_U3393;
  assign new_P2_U8166 = ~new_P2_U8152 | ~new_P2_U3488;
  assign new_P2_U8167 = ~new_P2_U3584 | ~new_P2_U3341;
  assign new_P2_U8168 = ~new_P2_U8152 | ~new_P2_U3442;
  assign new_P2_U8169 = ~new_P2_U3584 | ~new_P2_U3328;
  assign new_P2_U8170 = ~new_P2_U8152 | ~new_P2_U3432;
  assign new_P2_U8171 = ~new_P2_U3584 | ~new_P2_U3369;
  assign new_P2_U8172 = ~new_P2_U8152 | ~new_P2_U3466;
  assign new_P2_U8173 = ~new_P2_U3584 | ~new_P2_U3358;
  assign new_P2_U8174 = ~new_P2_U8152 | ~new_P2_U3455;
  assign new_P2_U8175 = ~new_P2_U3584 | ~new_P2_U3417;
  assign new_P2_U8176 = ~new_P2_U8152 | ~new_P2_U3512;
  assign new_P2_U8177 = ~new_P2_U3584 | ~new_P2_U3383;
  assign new_P2_U8178 = ~new_P2_U8152 | ~new_P2_U3478;
  assign new_P2_U8179 = ~new_P2_U3584 | ~new_P2_U3406;
  assign new_P2_U8180 = ~new_P2_U8152 | ~new_P2_U3501;
  assign new_P2_U8181 = ~new_P2_U3584 | ~new_P2_U3394;
  assign new_P2_U8182 = ~new_P2_U8152 | ~new_P2_U3489;
  assign new_P2_U8183 = ~new_P2_U3584 | ~new_P2_U3342;
  assign new_P2_U8184 = ~new_P2_U8152 | ~new_P2_U3443;
  assign new_P2_U8185 = ~new_P2_U3584 | ~new_P2_U3329;
  assign new_P2_U8186 = ~new_P2_U8152 | ~new_P2_U3433;
  assign new_P2_U8187 = ~new_P2_U3584 | ~new_P2_U3370;
  assign new_P2_U8188 = ~new_P2_U8152 | ~new_P2_U3467;
  assign new_P2_U8189 = ~new_P2_U3584 | ~new_P2_U3359;
  assign new_P2_U8190 = ~new_P2_U8152 | ~new_P2_U3456;
  assign new_P2_U8191 = ~new_P2_U3584 | ~new_P2_U3418;
  assign new_P2_U8192 = ~new_P2_U8152 | ~new_P2_U3513;
  assign new_P2_U8193 = ~new_P2_U3584 | ~new_P2_U3384;
  assign new_P2_U8194 = ~new_P2_U8152 | ~new_P2_U3479;
  assign new_P2_U8195 = ~new_P2_U3584 | ~new_P2_U3407;
  assign new_P2_U8196 = ~new_P2_U8152 | ~new_P2_U3502;
  assign new_P2_U8197 = ~new_P2_U3584 | ~new_P2_U3395;
  assign new_P2_U8198 = ~new_P2_U8152 | ~new_P2_U3490;
  assign new_P2_U8199 = ~new_P2_U3584 | ~new_P2_U3343;
  assign new_P2_U8200 = ~new_P2_U8152 | ~new_P2_U3444;
  assign new_P2_U8201 = ~new_P2_U3584 | ~new_P2_U3330;
  assign new_P2_U8202 = ~new_P2_U8152 | ~new_P2_U3434;
  assign new_P2_U8203 = ~new_P2_U3584 | ~new_P2_U3371;
  assign new_P2_U8204 = ~new_P2_U8152 | ~new_P2_U3468;
  assign new_P2_U8205 = ~new_P2_U3584 | ~new_P2_U3360;
  assign new_P2_U8206 = ~new_P2_U8152 | ~new_P2_U3457;
  assign new_P2_U8207 = ~new_P2_U3584 | ~new_P2_U3419;
  assign new_P2_U8208 = ~new_P2_U8152 | ~new_P2_U3514;
  assign new_P2_U8209 = ~new_P2_U3584 | ~new_P2_U3385;
  assign new_P2_U8210 = ~new_P2_U8152 | ~new_P2_U3480;
  assign new_P2_U8211 = ~new_P2_U3584 | ~new_P2_U3408;
  assign new_P2_U8212 = ~new_P2_U8152 | ~new_P2_U3503;
  assign new_P2_U8213 = ~new_P2_U3584 | ~new_P2_U3396;
  assign new_P2_U8214 = ~new_P2_U8152 | ~new_P2_U3491;
  assign new_P2_U8215 = ~new_P2_U3584 | ~new_P2_U3344;
  assign new_P2_U8216 = ~new_P2_U8152 | ~new_P2_U3445;
  assign new_P2_U8217 = ~new_P2_U3584 | ~new_P2_U3331;
  assign new_P2_U8218 = ~new_P2_U8152 | ~new_P2_U3435;
  assign new_P2_U8219 = ~new_P2_U3584 | ~new_P2_U3372;
  assign new_P2_U8220 = ~new_P2_U8152 | ~new_P2_U3469;
  assign new_P2_U8221 = ~new_P2_U3584 | ~new_P2_U3361;
  assign new_P2_U8222 = ~new_P2_U8152 | ~new_P2_U3458;
  assign new_P2_U8223 = ~new_P2_U3584 | ~new_P2_U3420;
  assign new_P2_U8224 = ~new_P2_U8152 | ~new_P2_U3515;
  assign new_P2_U8225 = ~new_P2_U3584 | ~new_P2_U3386;
  assign new_P2_U8226 = ~new_P2_U8152 | ~new_P2_U3481;
  assign new_P2_U8227 = ~new_P2_U3584 | ~new_P2_U3409;
  assign new_P2_U8228 = ~new_P2_U8152 | ~new_P2_U3504;
  assign new_P2_U8229 = ~new_P2_U3584 | ~new_P2_U3397;
  assign new_P2_U8230 = ~new_P2_U8152 | ~new_P2_U3492;
  assign new_P2_U8231 = ~new_P2_U3584 | ~new_P2_U3345;
  assign new_P2_U8232 = ~new_P2_U8152 | ~new_P2_U3446;
  assign new_P2_U8233 = ~new_P2_U3584 | ~new_P2_U3332;
  assign new_P2_U8234 = ~new_P2_U8152 | ~new_P2_U3436;
  assign new_P2_U8235 = ~new_P2_U3584 | ~new_P2_U3373;
  assign new_P2_U8236 = ~new_P2_U8152 | ~new_P2_U3470;
  assign new_P2_U8237 = ~new_P2_U3584 | ~new_P2_U3362;
  assign new_P2_U8238 = ~new_P2_U8152 | ~new_P2_U3459;
  assign new_P2_U8239 = ~new_P2_U3584 | ~new_P2_U3421;
  assign new_P2_U8240 = ~new_P2_U8152 | ~new_P2_U3516;
  assign new_P2_U8241 = ~new_P2_U3584 | ~new_P2_U3387;
  assign new_P2_U8242 = ~new_P2_U8152 | ~new_P2_U3482;
  assign new_P2_U8243 = ~new_P2_U3584 | ~new_P2_U3410;
  assign new_P2_U8244 = ~new_P2_U8152 | ~new_P2_U3505;
  assign new_P2_U8245 = ~new_P2_U3584 | ~new_P2_U3398;
  assign new_P2_U8246 = ~new_P2_U8152 | ~new_P2_U3493;
  assign new_P2_U8247 = ~new_P2_U3584 | ~new_P2_U3346;
  assign new_P2_U8248 = ~new_P2_U8152 | ~new_P2_U3447;
  assign new_P2_U8249 = ~new_P2_U3584 | ~new_P2_U3333;
  assign new_P2_U8250 = ~new_P2_U8152 | ~new_P2_U3437;
  assign new_P2_U8251 = ~new_P2_U3584 | ~new_P2_U3374;
  assign new_P2_U8252 = ~new_P2_U8152 | ~new_P2_U3471;
  assign new_P2_U8253 = ~new_P2_U3584 | ~new_P2_U3363;
  assign new_P2_U8254 = ~new_P2_U8152 | ~new_P2_U3460;
  assign new_P2_U8255 = ~new_P2_U3584 | ~new_P2_U3422;
  assign new_P2_U8256 = ~new_P2_U8152 | ~new_P2_U3517;
  assign new_P2_U8257 = ~new_P2_U3584 | ~new_P2_U3388;
  assign new_P2_U8258 = ~new_P2_U8152 | ~new_P2_U3483;
  assign new_P2_U8259 = ~new_P2_U3584 | ~new_P2_U3411;
  assign new_P2_U8260 = ~new_P2_U8152 | ~new_P2_U3506;
  assign new_P2_U8261 = ~new_P2_U3584 | ~new_P2_U3399;
  assign new_P2_U8262 = ~new_P2_U8152 | ~new_P2_U3494;
  assign new_P2_U8263 = ~new_P2_U3584 | ~new_P2_U3347;
  assign new_P2_U8264 = ~new_P2_U8152 | ~new_P2_U3448;
  assign new_P2_U8265 = ~new_P2_U3584 | ~new_P2_U3334;
  assign new_P2_U8266 = ~new_P2_U8152 | ~new_P2_U3438;
  assign new_P2_U8267 = ~new_P2_U3584 | ~new_P2_U3375;
  assign new_P2_U8268 = ~new_P2_U8152 | ~new_P2_U3472;
  assign new_P2_U8269 = ~new_P2_U3584 | ~new_P2_U3364;
  assign new_P2_U8270 = ~new_P2_U8152 | ~new_P2_U3461;
  assign new_P2_U8271 = ~new_P2_U3584 | ~new_P2_U3423;
  assign new_P2_U8272 = ~new_P2_U8152 | ~new_P2_U3518;
  assign new_P2_U8273 = ~new_P2_U3584 | ~new_P2_U3389;
  assign new_P2_U8274 = ~new_P2_U8152 | ~new_P2_U3484;
  assign new_P2_U8275 = ~new_P2_U3584 | ~new_P2_U3412;
  assign new_P2_U8276 = ~new_P2_U8152 | ~new_P2_U3507;
  assign new_P2_U8277 = ~new_P2_U3584 | ~new_P2_U3400;
  assign new_P2_U8278 = ~new_P2_U8152 | ~new_P2_U3495;
  assign new_P2_U8279 = ~new_P2_U3584 | ~new_P2_U3348;
  assign new_P2_U8280 = ~new_P2_U8152 | ~new_P2_U3449;
  assign new_P2_U8281 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_U3519;
  assign new_P2_U8282 = ~P2_FLUSH_REG | ~new_P2_U3598 | ~new_P2_U3597;
  assign new_P2_U8283 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_U3519;
  assign new_P2_U8284 = ~P2_FLUSH_REG | ~new_P2_U3597 | ~new_P2_U8090;
  assign new_P2_U8285 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_U3519;
  assign new_P2_U8286 = ~new_P2_U8087 | ~P2_FLUSH_REG;
  assign new_P2_U8287 = ~new_P2_U3616 | ~new_P2_U4406;
  assign new_P2_U8288 = ~new_P2_U5581 | ~P2_INSTQUEUERD_ADDR_REG_4_;
  assign new_P2_U8289 = ~new_P2_U5581 | ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign new_P2_U8290 = ~new_P2_U5611 | ~new_P2_U4406;
  assign new_P2_U8291 = ~new_P2_U5581 | ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign new_P2_U8292 = ~new_P2_U5619 | ~new_P2_U4406;
  assign new_P2_U8293 = ~new_P2_U5581 | ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_U8294 = ~new_P2_U5629 | ~new_P2_U4406;
  assign new_P2_U8295 = ~new_P2_U5581 | ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_U8296 = ~new_P2_U5637 | ~new_P2_U4406;
  assign new_P2_U8297 = ~new_P2_U3242 | ~new_P2_U7873;
  assign new_P2_U8298 = ~new_P2_U2616 | ~new_P2_U7183;
  assign new_P2_U8299 = ~new_P2_U7217 | ~new_P2_U7873;
  assign new_P2_U8300 = ~new_P2_U2616 | ~new_P2_U7200;
  assign new_P2_U8301 = ~new_P2_U7251 | ~new_P2_U7873;
  assign new_P2_U8302 = ~new_P2_U2616 | ~new_P2_U7234;
  assign new_P2_U8303 = ~new_P2_U7285 | ~new_P2_U7873;
  assign new_P2_U8304 = ~new_P2_U2616 | ~new_P2_U7268;
  assign new_P2_U8305 = ~new_P2_U7319 | ~new_P2_U7873;
  assign new_P2_U8306 = ~new_P2_U2616 | ~new_P2_U7302;
  assign new_P2_U8307 = ~new_P2_U7353 | ~new_P2_U7873;
  assign new_P2_U8308 = ~new_P2_U2616 | ~new_P2_U7336;
  assign new_P2_U8309 = ~new_P2_U7387 | ~new_P2_U7873;
  assign new_P2_U8310 = ~new_P2_U2616 | ~new_P2_U7370;
  assign new_P2_U8311 = ~new_P2_U7421 | ~new_P2_U7873;
  assign new_P2_U8312 = ~new_P2_U2616 | ~new_P2_U7404;
  assign new_P2_U8313 = ~new_P2_R2256_U5 | ~new_P2_U3572;
  assign new_P2_U8314 = ~new_P2_U3242 | ~new_P2_R2267_U56;
  assign new_P2_U8315 = ~new_P2_R2256_U17 | ~new_P2_U3572;
  assign new_P2_U8316 = ~new_P2_U3242 | ~new_P2_R2267_U19;
  assign new_P2_U8317 = ~new_P2_R2256_U18 | ~new_P2_U3572;
  assign new_P2_U8318 = ~new_P2_U3242 | ~new_P2_R2267_U58;
  assign new_P2_U8319 = ~new_P2_R2256_U19 | ~new_P2_U3572;
  assign new_P2_U8320 = ~new_P2_U3242 | ~new_P2_R2267_U18;
  assign new_P2_U8321 = ~new_P2_R2256_U20 | ~new_P2_U3572;
  assign new_P2_U8322 = ~new_P2_U3242 | ~new_P2_R2267_U60;
  assign new_P2_U8323 = ~new_P2_R2256_U26 | ~new_P2_U3572;
  assign new_P2_U8324 = ~new_P2_U3242 | ~new_P2_R2267_U17;
  assign new_P2_U8325 = ~new_P2_R2256_U22 | ~new_P2_U3572;
  assign new_P2_U8326 = ~new_P2_U3242 | ~new_P2_R2267_U65;
  assign new_P2_U8327 = ~new_P2_R2256_U4 | ~new_P2_U3572;
  assign new_P2_U8328 = ~new_P2_U3242 | ~new_P2_R2267_U43;
  assign new_P2_U8329 = ~new_P2_R2256_U21 | ~new_P2_U3572;
  assign new_P2_U8330 = ~new_P2_U3242 | ~new_P2_R2267_U21;
  assign new_P2_U8331 = ~new_P2_R2219_U24 | ~new_P2_U2617;
  assign new_P2_U8332 = ~P2_EBX_REG_7_ | ~new_P2_U7869;
  assign new_P2_U8333 = ~new_P2_R2219_U25 | ~new_P2_U2617;
  assign new_P2_U8334 = ~P2_EBX_REG_6_ | ~new_P2_U7869;
  assign new_P2_U8335 = ~new_P2_R2219_U26 | ~new_P2_U2617;
  assign new_P2_U8336 = ~P2_EBX_REG_5_ | ~new_P2_U7869;
  assign new_P2_U8337 = ~new_P2_R2219_U27 | ~new_P2_U2617;
  assign new_P2_U8338 = ~P2_EBX_REG_4_ | ~new_P2_U7869;
  assign new_P2_U8339 = ~new_P2_R2219_U28 | ~new_P2_U2617;
  assign new_P2_U8340 = ~P2_EBX_REG_3_ | ~new_P2_U7869;
  assign new_P2_U8341 = ~new_P2_R2219_U29 | ~new_P2_U2617;
  assign new_P2_U8342 = ~P2_EBX_REG_2_ | ~new_P2_U7869;
  assign new_P2_U8343 = ~new_P2_R2219_U30 | ~new_P2_U2617;
  assign new_P2_U8344 = ~P2_EBX_REG_1_ | ~new_P2_U7869;
  assign new_P2_U8345 = ~new_P2_R2219_U8 | ~new_P2_U2617;
  assign new_P2_U8346 = ~P2_EBX_REG_0_ | ~new_P2_U7869;
  assign new_P2_U8347 = ~new_P2_U3255 | ~new_P2_U7740;
  assign new_P2_U8348 = ~new_P2_U7867 | ~new_P2_U3525;
  assign new_P2_U8349 = ~new_P2_R2337_U68 | ~new_P2_U3284;
  assign new_P2_U8350 = ~P2_INSTADDRPOINTER_REG_31_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8351 = ~new_P2_R2238_U6 | ~new_P2_U3283;
  assign new_P2_U8352 = ~new_P2_SUB_450_U6 | ~new_P2_U4417;
  assign new_P2_U8353 = ~new_P2_R2238_U19 | ~new_P2_U3283;
  assign new_P2_U8354 = ~new_P2_SUB_450_U17 | ~new_P2_U4417;
  assign new_P2_U8355 = ~new_P2_R2238_U20 | ~new_P2_U3283;
  assign new_P2_U8356 = ~new_P2_SUB_450_U18 | ~new_P2_U4417;
  assign new_P2_U8357 = ~new_P2_R2238_U21 | ~new_P2_U3283;
  assign new_P2_U8358 = ~new_P2_SUB_450_U19 | ~new_P2_U4417;
  assign new_P2_U8359 = ~new_P2_R2238_U22 | ~new_P2_U3283;
  assign new_P2_U8360 = ~new_P2_SUB_450_U20 | ~new_P2_U4417;
  assign new_P2_U8361 = ~new_P2_R2337_U61 | ~new_P2_U3284;
  assign new_P2_U8362 = ~P2_INSTADDRPOINTER_REG_9_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8363 = ~new_P2_R2337_U62 | ~new_P2_U3284;
  assign new_P2_U8364 = ~P2_INSTADDRPOINTER_REG_8_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8365 = ~new_P2_R2337_U63 | ~new_P2_U3284;
  assign new_P2_U8366 = ~P2_INSTADDRPOINTER_REG_7_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8367 = ~new_P2_R2337_U64 | ~new_P2_U3284;
  assign new_P2_U8368 = ~P2_INSTADDRPOINTER_REG_6_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8369 = ~new_P2_R2337_U65 | ~new_P2_U3284;
  assign new_P2_U8370 = ~P2_INSTADDRPOINTER_REG_5_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8371 = ~new_P2_R2337_U66 | ~new_P2_U3284;
  assign new_P2_U8372 = ~P2_INSTADDRPOINTER_REG_4_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8373 = ~new_P2_R2337_U69 | ~new_P2_U3284;
  assign new_P2_U8374 = ~P2_INSTADDRPOINTER_REG_30_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8375 = ~new_P2_R2337_U67 | ~new_P2_U3284;
  assign new_P2_U8376 = ~P2_INSTADDRPOINTER_REG_3_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8377 = ~new_P2_R2337_U71 | ~new_P2_U3284;
  assign new_P2_U8378 = ~P2_INSTADDRPOINTER_REG_29_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8379 = ~new_P2_R2337_U72 | ~new_P2_U3284;
  assign new_P2_U8380 = ~P2_INSTADDRPOINTER_REG_28_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8381 = ~new_P2_R2337_U73 | ~new_P2_U3284;
  assign new_P2_U8382 = ~P2_INSTADDRPOINTER_REG_27_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8383 = ~new_P2_R2337_U74 | ~new_P2_U3284;
  assign new_P2_U8384 = ~P2_INSTADDRPOINTER_REG_26_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8385 = ~new_P2_R2337_U75 | ~new_P2_U3284;
  assign new_P2_U8386 = ~P2_INSTADDRPOINTER_REG_25_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8387 = ~new_P2_R2337_U76 | ~new_P2_U3284;
  assign new_P2_U8388 = ~P2_INSTADDRPOINTER_REG_24_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8389 = ~new_P2_R2337_U77 | ~new_P2_U3284;
  assign new_P2_U8390 = ~P2_INSTADDRPOINTER_REG_23_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8391 = ~new_P2_R2337_U78 | ~new_P2_U3284;
  assign new_P2_U8392 = ~P2_INSTADDRPOINTER_REG_22_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8393 = ~new_P2_R2337_U79 | ~new_P2_U3284;
  assign new_P2_U8394 = ~P2_INSTADDRPOINTER_REG_21_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8395 = ~new_P2_R2337_U80 | ~new_P2_U3284;
  assign new_P2_U8396 = ~P2_INSTADDRPOINTER_REG_20_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8397 = ~new_P2_R2337_U70 | ~new_P2_U3284;
  assign new_P2_U8398 = ~P2_INSTADDRPOINTER_REG_2_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8399 = ~new_P2_R2337_U81 | ~new_P2_U3284;
  assign new_P2_U8400 = ~P2_INSTADDRPOINTER_REG_19_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8401 = ~new_P2_R2337_U82 | ~new_P2_U3284;
  assign new_P2_U8402 = ~P2_INSTADDRPOINTER_REG_18_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8403 = ~new_P2_R2337_U83 | ~new_P2_U3284;
  assign new_P2_U8404 = ~P2_INSTADDRPOINTER_REG_17_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8405 = ~new_P2_R2337_U84 | ~new_P2_U3284;
  assign new_P2_U8406 = ~P2_INSTADDRPOINTER_REG_16_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8407 = ~new_P2_R2337_U85 | ~new_P2_U3284;
  assign new_P2_U8408 = ~P2_INSTADDRPOINTER_REG_15_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8409 = ~new_P2_R2337_U86 | ~new_P2_U3284;
  assign new_P2_U8410 = ~P2_INSTADDRPOINTER_REG_14_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8411 = ~new_P2_R2337_U87 | ~new_P2_U3284;
  assign new_P2_U8412 = ~P2_INSTADDRPOINTER_REG_13_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8413 = ~new_P2_R2337_U88 | ~new_P2_U3284;
  assign new_P2_U8414 = ~P2_INSTADDRPOINTER_REG_12_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8415 = ~new_P2_R2337_U89 | ~new_P2_U3284;
  assign new_P2_U8416 = ~P2_INSTADDRPOINTER_REG_11_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8417 = ~new_P2_R2337_U90 | ~new_P2_U3284;
  assign new_P2_U8418 = ~P2_INSTADDRPOINTER_REG_10_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8419 = ~new_P2_R2337_U4 | ~new_P2_U3284;
  assign new_P2_U8420 = ~P2_INSTADDRPOINTER_REG_1_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8421 = ~P2_PHYADDRPOINTER_REG_0_ | ~new_P2_U3284;
  assign new_P2_U8422 = ~P2_INSTADDRPOINTER_REG_0_ | ~P2_STATE2_REG_0_;
  assign new_P2_U8423 = ~new_P2_R2238_U6 | ~new_P2_U3269;
  assign new_P2_U8424 = ~new_P2_U2615 | ~P2_STATE2_REG_1_;
  assign new_P2_U8425 = ~new_P2_R2238_U19 | ~new_P2_U3269;
  assign new_P2_U8426 = ~new_P2_U2615 | ~P2_STATE2_REG_1_;
  assign new_P2_U8427 = ~new_P2_R2238_U20 | ~new_P2_U3269;
  assign new_P2_U8428 = ~new_P2_SUB_589_U8 | ~P2_STATE2_REG_1_;
  assign new_P2_U8429 = ~new_P2_R2238_U21 | ~new_P2_U3269;
  assign new_P2_U8430 = ~new_P2_SUB_589_U9 | ~P2_STATE2_REG_1_;
  assign new_P2_U8431 = ~new_P2_R2238_U22 | ~new_P2_U3269;
  assign new_P2_U8432 = ~new_P2_SUB_589_U6 | ~P2_STATE2_REG_1_;
  assign new_P2_U8433 = ~new_P2_R2238_U7 | ~new_P2_U3269;
  assign new_P2_U8434 = ~new_P2_SUB_589_U7 | ~P2_STATE2_REG_1_;
  assign new_P1_ADD_405_U171 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_ADD_405_U94;
  assign new_P1_ADD_405_U170 = ~new_P1_ADD_405_U126 | ~new_P1_ADD_405_U92;
  assign new_P1_ADD_405_U169 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_ADD_405_U93;
  assign new_P1_ADD_405_U168 = ~new_P1_ADD_405_U104 | ~new_P1_ADD_405_U21;
  assign new_P1_ADD_405_U167 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_ADD_405_U20;
  assign new_P1_ADD_405_U166 = ~new_P1_ADD_405_U113 | ~new_P1_ADD_405_U39;
  assign new_P1_ADD_405_U165 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_ADD_405_U38;
  assign new_P1_ADD_405_U164 = ~new_P1_ADD_405_U117 | ~new_P1_ADD_405_U47;
  assign new_P1_ADD_405_U163 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_ADD_405_U46;
  assign new_P1_ADD_405_U162 = ~new_P1_ADD_405_U102 | ~new_P1_ADD_405_U17;
  assign new_P1_ADD_405_U161 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_ADD_405_U16;
  assign new_P1_ADD_405_U160 = ~new_P1_ADD_405_U99 | ~new_P1_ADD_405_U11;
  assign new_P1_ADD_405_U159 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_ADD_405_U10;
  assign new_P1_ADD_405_U158 = ~new_P1_ADD_405_U108 | ~new_P1_ADD_405_U29;
  assign new_P1_ADD_405_U157 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_ADD_405_U28;
  assign new_P1_ADD_405_U156 = ~new_P1_ADD_405_U121 | ~new_P1_ADD_405_U55;
  assign new_P1_ADD_405_U155 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_ADD_405_U54;
  assign new_P1_ADD_405_U154 = ~new_P1_ADD_405_U98 | ~new_P1_ADD_405_U9;
  assign new_P1_ADD_405_U153 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_ADD_405_U8;
  assign new_P1_ADD_405_U152 = ~new_P1_ADD_405_U109 | ~new_P1_ADD_405_U31;
  assign new_P1_ADD_405_U151 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_ADD_405_U30;
  assign new_P1_ADD_405_U150 = ~new_P1_ADD_405_U120 | ~new_P1_ADD_405_U53;
  assign new_P1_ADD_405_U149 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_ADD_405_U52;
  assign new_P1_ADD_405_U148 = ~new_P1_ADD_405_U105 | ~new_P1_ADD_405_U23;
  assign new_P1_ADD_405_U147 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_ADD_405_U22;
  assign new_P1_ADD_405_U146 = ~new_P1_ADD_405_U112 | ~new_P1_ADD_405_U37;
  assign new_P1_ADD_405_U145 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_ADD_405_U36;
  assign new_P1_ADD_405_U144 = ~new_P1_ADD_405_U116 | ~new_P1_ADD_405_U45;
  assign new_P1_ADD_405_U143 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_ADD_405_U44;
  assign new_P1_ADD_405_U142 = ~new_P1_ADD_405_U103 | ~new_P1_ADD_405_U19;
  assign new_P1_ADD_405_U141 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_ADD_405_U18;
  assign new_P1_ADD_405_U140 = ~new_P1_ADD_405_U107 | ~new_P1_ADD_405_U27;
  assign new_P1_ADD_405_U139 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_ADD_405_U26;
  assign new_P1_ADD_405_U138 = ~new_P1_ADD_405_U114 | ~new_P1_ADD_405_U41;
  assign new_P1_ADD_405_U137 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_ADD_405_U40;
  assign new_P1_ADD_405_U136 = ~new_P1_ADD_405_U111 | ~new_P1_ADD_405_U35;
  assign new_P1_ADD_405_U135 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_ADD_405_U34;
  assign new_P1_ADD_405_U134 = ~new_P1_ADD_405_U118 | ~new_P1_ADD_405_U49;
  assign new_P1_ADD_405_U133 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_ADD_405_U48;
  assign new_P1_ADD_405_U132 = ~new_P1_ADD_405_U123 | ~new_P1_ADD_405_U59;
  assign new_P1_ADD_405_U131 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_ADD_405_U58;
  assign new_P1_ADD_405_U130 = ~new_P1_ADD_405_U124 | ~new_P1_ADD_405_U60;
  assign new_P1_ADD_405_U129 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_ADD_405_U61;
  assign new_P1_ADD_405_U128 = ~new_P1_ADD_405_U100 | ~new_P1_ADD_405_U12;
  assign new_P1_ADD_405_U127 = ~P1_INSTADDRPOINTER_REG_6_ | ~new_P1_ADD_405_U13;
  assign new_P1_ADD_405_U126 = ~new_P1_ADD_405_U93;
  assign new_P1_ADD_405_U125 = ~P1_INSTADDRPOINTER_REG_2_ | ~P1_INSTADDRPOINTER_REG_1_ | ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_ADD_405_U124 = ~new_P1_ADD_405_U61;
  assign new_P1_ADD_405_U123 = ~new_P1_ADD_405_U58;
  assign new_P1_ADD_405_U122 = ~new_P1_ADD_405_U56;
  assign new_P1_ADD_405_U121 = ~new_P1_ADD_405_U54;
  assign new_P1_ADD_405_U120 = ~new_P1_ADD_405_U52;
  assign new_P1_ADD_405_U119 = ~new_P1_ADD_405_U50;
  assign new_P1_ADD_405_U118 = ~new_P1_ADD_405_U48;
  assign new_P1_ADD_405_U117 = ~new_P1_ADD_405_U46;
  assign new_P1_ADD_405_U116 = ~new_P1_ADD_405_U44;
  assign new_P1_ADD_405_U115 = ~new_P1_ADD_405_U42;
  assign new_P1_U2352 = ~P1_STATEBS16_REG & ~P1_STATE2_REG_2_;
  assign new_P1_U2353 = new_P1_U4231 & P1_STATE2_REG_2_;
  assign new_P1_U2354 = new_P1_U4265 & new_P1_U4477;
  assign new_P1_U2355 = new_P1_U3234 & new_P1_U2450;
  assign new_P1_U2356 = new_P1_R2238_U6 & new_P1_U4192;
  assign new_P1_U2357 = new_P1_R2167_U17 & new_P1_U5959 & new_P1_U3865;
  assign new_P1_U2358 = new_P1_U2388 & new_P1_U4224;
  assign new_P1_U2359 = P1_STATE2_REG_2_ & new_P1_U3431;
  assign new_P1_U2360 = P1_STATE2_REG_2_ & new_P1_U3414;
  assign new_P1_U2361 = new_P1_U4224 & P1_STATE2_REG_3_;
  assign new_P1_U2362 = new_P1_U2359 & new_P1_U4208;
  assign new_P1_U2363 = new_P1_U2359 & new_P1_U4210;
  assign new_P1_U2364 = new_P1_U3864 & new_P1_U3416;
  assign new_P1_U2365 = new_P1_U4261 & new_P1_U3416;
  assign new_P1_U2366 = new_P1_U3430 & new_P1_U3431 & P1_STATE2_REG_1_;
  assign new_P1_U2367 = new_P1_R2337_U69 & P1_STATE2_REG_1_ & new_P1_U3431;
  assign new_P1_U2368 = new_P1_U4235 & P1_STATE2_REG_0_;
  assign new_P1_U2369 = new_P1_U2362 & new_P1_U4497;
  assign new_P1_U2370 = new_P1_U3414 & new_P1_U3263;
  assign new_P1_U2371 = new_P1_U4222 & new_P1_U4449;
  assign new_P1_U2372 = P1_STATE2_REG_0_ & new_P1_U3416;
  assign new_P1_U2373 = P1_STATE2_REG_3_ & new_P1_U3431;
  assign new_P1_U2374 = new_P1_U2360 & new_P1_U4214;
  assign new_P1_U2375 = new_P1_U2360 & new_P1_U4216;
  assign new_P1_U2376 = new_P1_U5798 & new_P1_U3416;
  assign new_P1_U2377 = new_P1_U3762 & new_P1_U3414;
  assign new_P1_U2378 = new_P1_U2360 & new_P1_U5569;
  assign new_P1_U2379 = new_P1_U2363 & new_P1_U3280;
  assign new_P1_U2380 = new_P1_U2360 & new_P1_U7608;
  assign new_P1_U2381 = new_P1_U2357 & new_P1_U3271;
  assign new_P1_U2382 = new_P1_U2357 & new_P1_U4477;
  assign new_P1_U2383 = new_P1_U4222 & new_P1_U3391;
  assign new_P1_U2384 = P1_STATE2_REG_0_ & new_P1_U3417;
  assign new_P1_U2385 = new_P1_U3417 & new_P1_U3294;
  assign new_P1_U2386 = new_P1_U4223 & new_P1_U3423;
  assign new_P1_U2387 = new_P1_U3884 & new_P1_U4223;
  assign new_P1_U2388 = P1_STATEBS16_REG & new_P1_U4209;
  assign new_P1_U2389 = new_P1_U2452 & new_P1_U7494;
  assign new_P1_U2390 = new_U346 & new_P1_U4224;
  assign new_P1_U2391 = new_U335 & new_P1_U4224;
  assign new_P1_U2392 = new_U324 & new_P1_U4224;
  assign new_P1_U2393 = new_U321 & new_P1_U4224;
  assign new_P1_U2394 = new_U320 & new_P1_U4224;
  assign new_P1_U2395 = new_U319 & new_P1_U4224;
  assign new_P1_U2396 = new_U318 & new_P1_U4224;
  assign new_P1_U2397 = new_U317 & new_P1_U4224;
  assign new_P1_U2398 = new_U330 & new_P1_U2358;
  assign new_P1_U2399 = new_U339 & new_P1_U2358;
  assign new_P1_U2400 = new_U329 & new_P1_U2358;
  assign new_P1_U2401 = new_U338 & new_P1_U2358;
  assign new_P1_U2402 = new_U328 & new_P1_U2358;
  assign new_P1_U2403 = new_U337 & new_P1_U2358;
  assign new_P1_U2404 = new_U327 & new_P1_U2358;
  assign new_P1_U2405 = new_U336 & new_P1_U2358;
  assign new_P1_U2406 = new_U326 & new_P1_U2358;
  assign new_P1_U2407 = new_U334 & new_P1_U2358;
  assign new_P1_U2408 = new_U325 & new_P1_U2358;
  assign new_P1_U2409 = new_U333 & new_P1_U2358;
  assign new_P1_U2410 = new_U323 & new_P1_U2358;
  assign new_P1_U2411 = new_U332 & new_P1_U2358;
  assign new_P1_U2412 = new_U322 & new_P1_U2358;
  assign new_P1_U2413 = new_U331 & new_P1_U2358;
  assign new_P1_U2414 = new_P1_U2361 & new_P1_U3271;
  assign new_P1_U2415 = new_P1_U2361 & new_P1_U3391;
  assign new_P1_U2416 = new_P1_U2361 & new_P1_U3277;
  assign new_P1_U2417 = new_P1_U2361 & new_P1_U3284;
  assign new_P1_U2418 = new_P1_U2361 & new_P1_U3283;
  assign new_P1_U2419 = new_P1_U2361 & new_P1_U3278;
  assign new_P1_U2420 = new_P1_U2361 & new_P1_U4173;
  assign new_P1_U2421 = new_P1_U2361 & new_P1_U4171;
  assign new_P1_U2422 = new_P1_U4223 & new_P1_U5461;
  assign new_P1_U2423 = new_P1_U4223 & new_P1_U4231;
  assign new_P1_U2424 = new_P1_U2384 & new_P1_U3284;
  assign new_P1_U2425 = new_P1_U2368 & new_P1_U2448;
  assign new_P1_U2426 = new_P1_U3889 & new_P1_U3431;
  assign new_P1_U2427 = ~P1_STATE2_REG_1_ & ~P1_STATE2_REG_3_;
  assign new_P1_U2428 = P1_STATE2_REG_2_ & P1_STATE2_REG_1_;
  assign new_P1_U2429 = new_P1_U6366 & new_P1_U3431;
  assign new_P1_U2430 = P1_STATE2_REG_1_ & new_P1_U3387;
  assign new_P1_U2431 = new_P1_U4199 & new_P1_U7494;
  assign new_P1_U2432 = new_P1_U3455 & new_P1_U3360;
  assign new_P1_U2433 = new_P1_U4540 & new_P1_U3455;
  assign new_P1_U2434 = new_P1_U7696 & new_P1_U3360;
  assign new_P1_U2435 = new_P1_U4540 & new_P1_U7696;
  assign new_P1_U2436 = new_P1_U3235 & new_P1_U3301;
  assign new_P1_U2437 = new_P1_U4543 & new_P1_U3301;
  assign new_P1_U2438 = new_P1_R2182_U42 & new_P1_R2182_U25;
  assign new_P1_U2439 = new_P1_R2182_U42 & new_P1_U3316;
  assign new_P1_U2440 = new_P1_R2182_U25 & new_P1_U3317;
  assign new_P1_U2441 = ~new_P1_R2182_U42 & ~new_P1_R2182_U25;
  assign new_P1_U2442 = new_P1_R2182_U33 & new_P1_R2182_U34;
  assign new_P1_U2443 = new_P1_R2182_U33 & new_P1_U3318;
  assign new_P1_U2444 = new_P1_R2182_U34 & new_P1_U3319;
  assign new_P1_U2445 = ~new_P1_R2182_U33 & ~new_P1_R2182_U34;
  assign new_P1_U2446 = P1_STATE2_REG_1_ & new_P1_U3471;
  assign new_P1_U2447 = new_P1_U3577 & new_P1_U2452;
  assign new_P1_U2448 = new_P1_R2167_U17 & new_P1_U3284;
  assign new_P1_U2449 = new_P1_U4494 & new_P1_U3271;
  assign new_P1_U2450 = P1_STATE2_REG_0_ & new_P1_U4400;
  assign new_P1_U2451 = new_P1_U4251 & P1_STATE2_REG_0_;
  assign new_P1_U2452 = new_P1_U4173 & new_P1_U3391 & new_P1_U4400 & new_P1_U3277;
  assign new_P1_U2453 = P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U2454 = P1_INSTQUEUERD_ADDR_REG_1_ & new_P1_U3266;
  assign new_P1_U2455 = new_P1_U3266 & P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U2456 = P1_INSTQUEUERD_ADDR_REG_0_ & new_P1_U3265;
  assign new_P1_U2457 = new_P1_U3265 & P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U2458 = new_P1_U3507 & new_P1_U4378;
  assign new_P1_U2459 = new_P1_U3264 & P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U2460 = P1_INSTQUEUERD_ADDR_REG_1_ & new_P1_U3264 & new_P1_U3266;
  assign new_P1_U2461 = new_P1_U3506 & new_P1_U3505;
  assign new_P1_U2462 = P1_INSTQUEUERD_ADDR_REG_0_ & new_P1_U3264 & new_P1_U3265;
  assign new_P1_U2463 = new_P1_U3504 & new_P1_U3503;
  assign new_P1_U2464 = P1_INSTQUEUERD_ADDR_REG_3_ & new_P1_U4380;
  assign new_P1_U2465 = new_P1_U3502 & new_P1_U3501;
  assign new_P1_U2466 = new_P1_U3500 & new_P1_U3499;
  assign new_P1_U2467 = new_P1_U4378 & P1_INSTQUEUERD_ADDR_REG_2_ & new_P1_U3270;
  assign new_P1_U2468 = new_P1_U3498 & new_P1_U3497;
  assign new_P1_U2469 = ~P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U2470 = new_P1_U2469 & P1_INSTQUEUERD_ADDR_REG_1_ & new_P1_U3266;
  assign new_P1_U2471 = new_P1_U2469 & P1_INSTQUEUERD_ADDR_REG_0_ & new_P1_U3265;
  assign new_P1_U2472 = new_P1_U4380 & new_P1_U3270;
  assign new_P1_U2473 = new_P1_U3406 & new_P1_U7680 & new_P1_U7679;
  assign new_P1_U2474 = new_P1_R2144_U49 & new_P1_U3312;
  assign new_P1_U2475 = new_P1_U3454 & new_P1_U3358;
  assign new_P1_U2476 = new_P1_R2144_U8 & new_P1_R2144_U49;
  assign new_P1_U2477 = new_P1_U4528 & new_P1_U2476;
  assign new_P1_U2478 = P1_INSTQUEUEWR_ADDR_REG_2_ & P1_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P1_U2479 = P1_INSTQUEUEWR_ADDR_REG_2_ & new_P1_U3303;
  assign new_P1_U2480 = new_P1_U3315 & new_P1_U4548;
  assign new_P1_U2481 = new_P1_U4524 & new_P1_U2476;
  assign new_P1_U2482 = new_P1_U3327 & new_P1_U4606;
  assign new_P1_U2483 = new_P1_U4525 & new_P1_U2476;
  assign new_P1_U2484 = new_P1_U3334 & new_P1_U4665;
  assign new_P1_U2485 = new_P1_U4526 & new_P1_R2144_U43;
  assign new_P1_U2486 = ~new_P1_R2144_U43 & ~new_P1_R2144_U50;
  assign new_P1_U2487 = new_P1_U2486 & new_P1_U2476;
  assign new_P1_U2488 = ~P1_INSTQUEUEWR_ADDR_REG_0_ & ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P1_U2489 = new_P1_U3338 & new_P1_U4722;
  assign new_P1_U2490 = new_P1_U7693 & new_P1_U3358;
  assign new_P1_U2491 = new_P1_U4529 & new_P1_U4528;
  assign new_P1_U2492 = new_P1_U3343 & new_P1_U4780;
  assign new_P1_U2493 = new_P1_U4529 & new_P1_U4524;
  assign new_P1_U2494 = new_P1_U3347 & new_P1_U4837;
  assign new_P1_U2495 = new_P1_U4529 & new_P1_U4525;
  assign new_P1_U2496 = new_P1_U3350 & new_P1_U4895;
  assign new_P1_U2497 = new_P1_U4529 & new_P1_U2486;
  assign new_P1_U2498 = new_P1_U3354 & new_P1_U4952;
  assign new_P1_U2499 = new_P1_U4531 & new_P1_U3454;
  assign new_P1_U2500 = new_P1_U3359 & new_P1_U3357;
  assign new_P1_U2501 = new_P1_U4524 & new_P1_U2474;
  assign new_P1_U2502 = new_P1_U3364 & new_P1_U5065;
  assign new_P1_U2503 = new_P1_U4525 & new_P1_U2474;
  assign new_P1_U2504 = new_P1_U3367 & new_P1_U5123;
  assign new_P1_U2505 = new_P1_U2486 & new_P1_U2474;
  assign new_P1_U2506 = new_P1_U3371 & new_P1_U5180;
  assign new_P1_U2507 = new_P1_U4531 & new_P1_U7693;
  assign new_P1_U2508 = ~new_P1_R2144_U49 & ~new_P1_R2144_U8;
  assign new_P1_U2509 = new_P1_U2508 & new_P1_U4528;
  assign new_P1_U2510 = ~P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P1_U2511 = new_P1_U3374 & new_P1_U5238;
  assign new_P1_U2512 = new_P1_U2508 & new_P1_U4524;
  assign new_P1_U2513 = new_P1_U3378 & new_P1_U5295;
  assign new_P1_U2514 = new_P1_U2508 & new_P1_U4525;
  assign new_P1_U2515 = new_P1_U3381 & new_P1_U5353;
  assign new_P1_U2516 = new_P1_U2508 & new_P1_U2486;
  assign new_P1_U2517 = new_P1_U3385 & new_P1_U5410;
  assign new_P1_U2518 = new_P1_U5468 & new_P1_U7700 & new_P1_U7699;
  assign new_P1_U2519 = new_P1_U3744 & new_P1_U5499;
  assign new_P1_U2520 = new_P1_U4219 & new_P1_U3446;
  assign new_P1_U2521 = P1_INSTQUEUERD_ADDR_REG_0_ & new_P1_U3402;
  assign new_P1_U2522 = new_P1_U5483 & new_P1_U5511;
  assign new_P1_U2523 = new_P1_U2522 & new_P1_U2521;
  assign new_P1_U2524 = new_P1_U3266 & new_P1_U3402;
  assign new_P1_U2525 = new_P1_U2522 & new_P1_U2524;
  assign new_P1_U2526 = new_P1_U5519 & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U2527 = new_P1_U2522 & new_P1_U2526;
  assign new_P1_U2528 = new_P1_U5519 & new_P1_U3266;
  assign new_P1_U2529 = new_P1_U2522 & new_P1_U2528;
  assign new_P1_U2530 = new_P1_U5483 & new_P1_U3401;
  assign new_P1_U2531 = new_P1_U2530 & new_P1_U2521;
  assign new_P1_U2532 = new_P1_U2530 & new_P1_U2524;
  assign new_P1_U2533 = new_P1_U2530 & new_P1_U2526;
  assign new_P1_U2534 = new_P1_U2530 & new_P1_U2528;
  assign new_P1_U2535 = new_P1_U5511 & new_P1_U3438;
  assign new_P1_U2536 = new_P1_U2535 & new_P1_U2521;
  assign new_P1_U2537 = new_P1_U2535 & new_P1_U2524;
  assign new_P1_U2538 = new_P1_U2535 & new_P1_U2526;
  assign new_P1_U2539 = new_P1_U2535 & new_P1_U2528;
  assign new_P1_U2540 = new_P1_U3438 & new_P1_U3401;
  assign new_P1_U2541 = new_P1_U2521 & new_P1_U2540;
  assign new_P1_U2542 = new_P1_U2524 & new_P1_U2540;
  assign new_P1_U2543 = new_P1_U2526 & new_P1_U2540;
  assign new_P1_U2544 = new_P1_U2528 & new_P1_U2540;
  assign new_P1_U2545 = new_P1_U5480 & new_P1_U7720;
  assign new_P1_U2546 = new_P1_U2545 & new_P1_U2454;
  assign new_P1_U2547 = new_P1_U2545 & new_P1_U3498;
  assign new_P1_U2548 = new_P1_U2545 & new_P1_U4378;
  assign new_P1_U2549 = new_P1_U2545 & new_P1_U2456;
  assign new_P1_U2550 = new_P1_U5480 & new_P1_U3456;
  assign new_P1_U2551 = new_P1_U2550 & new_P1_U2454;
  assign new_P1_U2552 = new_P1_U2550 & new_P1_U3498;
  assign new_P1_U2553 = new_P1_U2550 & new_P1_U4378;
  assign new_P1_U2554 = new_P1_U2550 & new_P1_U2456;
  assign new_P1_U2555 = new_P1_U7720 & new_P1_U3442;
  assign new_P1_U2556 = new_P1_U2555 & new_P1_U2454;
  assign new_P1_U2557 = new_P1_U2555 & new_P1_U3498;
  assign new_P1_U2558 = new_P1_U2555 & new_P1_U4378;
  assign new_P1_U2559 = new_P1_U2555 & new_P1_U2456;
  assign new_P1_U2560 = new_P1_U3456 & new_P1_U3442;
  assign new_P1_U2561 = new_P1_U2560 & new_P1_U2454;
  assign new_P1_U2562 = new_P1_U2560 & new_P1_U3498;
  assign new_P1_U2563 = new_P1_U2560 & new_P1_U4378;
  assign new_P1_U2564 = new_P1_U2560 & new_P1_U2456;
  assign new_P1_U2565 = new_P1_U7065 & new_P1_U4379;
  assign new_P1_U2566 = new_P1_U7065 & new_P1_U2460;
  assign new_P1_U2567 = new_P1_U7065 & new_P1_U2462;
  assign new_P1_U2568 = new_P1_U7065 & new_P1_U4380;
  assign new_P1_U2569 = new_P1_U7065 & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U2570 = new_P1_U2569 & new_P1_U3498;
  assign new_P1_U2571 = new_P1_U2569 & new_P1_U2454;
  assign new_P1_U2572 = new_P1_U2569 & new_P1_U2456;
  assign new_P1_U2573 = new_P1_U2569 & new_P1_U4378;
  assign new_P1_U2574 = new_P1_U4379 & new_P1_U3445;
  assign new_P1_U2575 = new_P1_U2460 & new_P1_U3445;
  assign new_P1_U2576 = new_P1_U2462 & new_P1_U3445;
  assign new_P1_U2577 = new_P1_U4380 & new_P1_U3445;
  assign new_P1_U2578 = P1_INSTQUEUERD_ADDR_REG_2_ & new_P1_U3445;
  assign new_P1_U2579 = new_P1_U2578 & new_P1_U3498;
  assign new_P1_U2580 = new_P1_U2578 & new_P1_U2454;
  assign new_P1_U2581 = new_P1_U2578 & new_P1_U2456;
  assign new_P1_U2582 = new_P1_U2578 & new_P1_U4378;
  assign new_P1_U2583 = new_P1_U7790 & new_P1_U4184;
  assign new_P1_U2584 = new_P1_U2583 & new_P1_U2524;
  assign new_P1_U2585 = new_P1_U2583 & new_P1_U2521;
  assign new_P1_U2586 = new_P1_U2583 & new_P1_U2528;
  assign new_P1_U2587 = new_P1_U2583 & new_P1_U2526;
  assign new_P1_U2588 = new_P1_U7790 & new_P1_U3452;
  assign new_P1_U2589 = new_P1_U2588 & new_P1_U2524;
  assign new_P1_U2590 = new_P1_U2588 & new_P1_U2521;
  assign new_P1_U2591 = new_P1_U2588 & new_P1_U2528;
  assign new_P1_U2592 = new_P1_U2588 & new_P1_U2526;
  assign new_P1_U2593 = new_P1_U4184 & new_P1_U3457;
  assign new_P1_U2594 = new_P1_U2593 & new_P1_U2524;
  assign new_P1_U2595 = new_P1_U2593 & new_P1_U2521;
  assign new_P1_U2596 = new_P1_U2593 & new_P1_U2528;
  assign new_P1_U2597 = new_P1_U2593 & new_P1_U2526;
  assign new_P1_U2598 = new_P1_U3457 & new_P1_U3452;
  assign new_P1_U2599 = new_P1_U2598 & new_P1_U2524;
  assign new_P1_U2600 = new_P1_U2598 & new_P1_U2521;
  assign new_P1_U2601 = new_P1_U2598 & new_P1_U2528;
  assign new_P1_U2602 = new_P1_U2598 & new_P1_U2526;
  assign new_P1_U2603 = P1_STATE2_REG_0_ & new_P1_U3389;
  assign new_P1_U2604 = P1_EBX_REG_31_ & new_P1_U2379;
  assign new_P1_U2605 = new_P1_U3530 & new_P1_U3531 & new_P1_U3532 & new_P1_U3533 & new_P1_U2607;
  assign new_P1_U2606 = new_P1_U7504 & new_P1_U3427;
  assign new_P1_U2607 = new_P1_U7672 & new_P1_U7671;
  assign new_P1_U2608 = new_P1_U7787 & new_P1_U7786;
  assign new_P1_U2609 = ~new_P1_U6855 | ~new_P1_U6853 | ~new_P1_U6854;
  assign new_P1_U2610 = ~new_P1_U6856 | ~new_P1_U4026;
  assign new_P1_U2611 = ~new_P1_U6843 | ~new_P1_U6841 | ~new_P1_U6842;
  assign new_P1_U2612 = ~new_P1_U6846 | ~new_P1_U6844 | ~new_P1_U6845;
  assign new_P1_U2613 = ~new_P1_U6849 | ~new_P1_U6847 | ~new_P1_U6848;
  assign new_P1_U2614 = ~new_P1_U6756 | ~new_P1_U4005;
  assign new_P1_U2615 = ~new_P1_U6753 | ~new_P1_U4004;
  assign new_P1_U2616 = ~new_P1_U6852 | ~new_P1_U6850 | ~new_P1_U6851;
  assign new_P1_U2617 = ~new_P1_U6750 | ~new_P1_U4003;
  assign new_P1_U2618 = ~new_P1_U6747 | ~new_P1_U4002;
  assign new_P1_ADD_405_U114 = ~new_P1_ADD_405_U40;
  assign new_P1_U2620 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2621 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2622 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2623 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2624 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2625 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2626 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2627 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2628 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2629 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2630 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2631 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2632 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2633 = new_P1_R2144_U145 & new_P1_U6746;
  assign new_P1_U2634 = new_P1_R2144_U11 & new_P1_U6746;
  assign new_P1_U2635 = new_P1_R2144_U37 & new_P1_U6746;
  assign new_P1_U2636 = new_P1_R2144_U38 & new_P1_U6746;
  assign new_P1_U2637 = new_P1_R2144_U39 & new_P1_U6746;
  assign new_P1_U2638 = new_P1_R2144_U40 & new_P1_U6746;
  assign new_P1_U2639 = new_P1_R2144_U41 & new_P1_U6746;
  assign new_P1_U2640 = new_P1_R2144_U42 & new_P1_U6746;
  assign new_P1_U2641 = new_P1_R2144_U30 & new_P1_U6746;
  assign new_P1_U2642 = new_P1_R2144_U80 & new_P1_U6746;
  assign new_P1_U2643 = new_P1_R2144_U10 & new_P1_U6746;
  assign new_P1_U2644 = new_P1_R2144_U9 & new_P1_U6746;
  assign new_P1_U2645 = new_P1_R2144_U45 & new_P1_U6746;
  assign new_P1_U2646 = new_P1_R2144_U47 & new_P1_U6746;
  assign new_P1_U2647 = new_P1_R2144_U8 & new_P1_U6746;
  assign new_P1_U2648 = ~new_P1_U3440 | ~new_P1_U6869;
  assign new_P1_U2649 = new_P1_R2144_U50 & new_P1_U6746;
  assign new_P1_U2650 = P1_STATE2_REG_2_ & new_P1_U6870;
  assign new_P1_U2651 = ~new_P1_U6770 | ~new_P1_U6769 | ~new_P1_U6768;
  assign new_P1_U2652 = ~new_P1_U6771 | ~new_P1_U4009;
  assign new_P1_U2653 = ~new_P1_U6780 | ~new_P1_U4011;
  assign new_P1_U2654 = ~new_P1_U6784 | ~new_P1_U4012;
  assign new_P1_U2655 = ~new_P1_U6788 | ~new_P1_U4013;
  assign new_P1_U2656 = ~new_P1_U6792 | ~new_P1_U4014;
  assign new_P1_U2657 = ~new_P1_U6796 | ~new_P1_U4015;
  assign new_P1_U2658 = ~new_P1_U6800 | ~new_P1_U4016;
  assign new_P1_U2659 = ~new_P1_U6804 | ~new_P1_U4017;
  assign new_P1_U2660 = ~new_P1_U6808 | ~new_P1_U4018;
  assign new_P1_U2661 = ~new_P1_U6812 | ~new_P1_U4019;
  assign new_P1_U2662 = ~new_P1_U6816 | ~new_P1_U4020;
  assign new_P1_U2663 = ~new_P1_U6825 | ~new_P1_U4022;
  assign new_P1_U2664 = ~new_P1_U6829 | ~new_P1_U4023;
  assign new_P1_U2665 = ~new_P1_U6833 | ~new_P1_U4024;
  assign new_P1_U2666 = ~new_P1_U6837 | ~new_P1_U4025;
  assign new_P1_U2667 = ~new_P1_U6759 | ~new_P1_U4006;
  assign new_P1_U2668 = ~new_P1_U6763 | ~new_P1_U4008 | ~new_P1_U6767 | ~new_P1_U6766;
  assign new_P1_U2669 = ~new_P1_U6775 | ~new_P1_U4010 | ~new_P1_U6779 | ~new_P1_U6778;
  assign new_P1_U2670 = ~new_P1_U6820 | ~new_P1_U4021 | ~new_P1_U6824 | ~new_P1_U6823;
  assign new_P1_U2671 = ~new_P1_U6859 | ~new_P1_U4027 | ~new_P1_U6863 | ~new_P1_U6862;
  assign new_P1_U2672 = ~new_P1_U6867 | ~new_P1_U6868 | ~new_P1_U6865 | ~new_P1_U6866 | ~new_P1_U6864;
  assign new_P1_U2673 = ~new_P1_U7458 | ~new_P1_U7457;
  assign new_P1_U2674 = ~new_P1_U7460 | ~new_P1_U7459;
  assign new_P1_U2675 = ~new_P1_U4168 | ~new_P1_U7463;
  assign new_P1_U2676 = ~new_P1_U4169 | ~new_P1_U7466;
  assign new_P1_U2677 = ~new_P1_U7467 | ~new_P1_U7794 | ~new_P1_U7793;
  assign new_P1_U2678 = ~new_P1_U7456 | ~new_P1_U3284;
  assign new_P1_U2679 = ~new_P1_U7405 | ~new_P1_U7404;
  assign new_P1_U2680 = ~new_P1_U7407 | ~new_P1_U7406;
  assign new_P1_U2681 = ~new_P1_U7411 | ~new_P1_U7410;
  assign new_P1_U2682 = ~new_P1_U7413 | ~new_P1_U7412;
  assign new_P1_U2683 = ~new_P1_U7415 | ~new_P1_U7414;
  assign new_P1_U2684 = ~new_P1_U7417 | ~new_P1_U7416;
  assign new_P1_U2685 = ~new_P1_U7419 | ~new_P1_U7418;
  assign new_P1_U2686 = ~new_P1_U7421 | ~new_P1_U7420;
  assign new_P1_U2687 = ~new_P1_U7423 | ~new_P1_U7422;
  assign new_P1_U2688 = ~new_P1_U7425 | ~new_P1_U7424;
  assign new_P1_U2689 = ~new_P1_U7427 | ~new_P1_U7426;
  assign new_P1_U2690 = ~new_P1_U7429 | ~new_P1_U7428;
  assign new_P1_U2691 = ~new_P1_U7433 | ~new_P1_U7432;
  assign new_P1_U2692 = ~new_P1_U7435 | ~new_P1_U7434;
  assign new_P1_U2693 = ~new_P1_U7437 | ~new_P1_U7436;
  assign new_P1_U2694 = ~new_P1_U7439 | ~new_P1_U7438;
  assign new_P1_U2695 = ~new_P1_U7441 | ~new_P1_U7440;
  assign new_P1_U2696 = ~new_P1_U7443 | ~new_P1_U7442;
  assign new_P1_U2697 = ~new_P1_U7445 | ~new_P1_U7444;
  assign new_P1_U2698 = ~new_P1_U7447 | ~new_P1_U7446;
  assign new_P1_U2699 = ~new_P1_U7449 | ~new_P1_U7448;
  assign new_P1_U2700 = ~new_P1_U7451 | ~new_P1_U7450;
  assign new_P1_U2701 = ~new_P1_U7393 | ~new_P1_U7392;
  assign new_P1_U2702 = ~new_P1_U7395 | ~new_P1_U7394;
  assign new_P1_U2703 = ~new_P1_U7397 | ~new_P1_U7396;
  assign new_P1_U2704 = ~new_P1_U7399 | ~new_P1_U7398;
  assign new_P1_U2705 = ~new_P1_U7401 | ~new_P1_U7400;
  assign new_P1_U2706 = ~new_P1_U7403 | ~new_P1_U7402;
  assign new_P1_U2707 = ~new_P1_U7409 | ~new_P1_U7408;
  assign new_P1_U2708 = ~new_P1_U7431 | ~new_P1_U7430;
  assign new_P1_U2709 = ~new_P1_U7453 | ~new_P1_U7452;
  assign new_P1_U2710 = ~new_P1_U7455 | ~new_P1_U7454;
  assign new_P1_U2711 = ~new_P1_U7377 | ~new_P1_U7376;
  assign new_P1_U2712 = ~new_P1_U7379 | ~new_P1_U7378;
  assign new_P1_U2713 = ~new_P1_U4165 | ~new_P1_U4239;
  assign new_P1_U2714 = ~new_P1_U3434 | ~new_P1_U4166 | ~new_P1_U7386 | ~new_P1_U7385;
  assign new_P1_U2715 = ~new_P1_U4239 | ~new_P1_U4167;
  assign new_P1_U2716 = ~new_P1_U7365 | ~new_P1_U7364;
  assign new_P1_U2717 = ~new_P1_U7367 | ~new_P1_U7366;
  assign new_P1_U2718 = ~new_P1_U4161 | ~new_P1_U7368;
  assign new_P1_U2719 = ~new_P1_U4162 | ~new_P1_U7370;
  assign new_P1_U2720 = ~new_P1_U4163 | ~new_P1_U7372;
  assign new_P1_U2721 = ~new_P1_U4164 | ~new_P1_U7374;
  assign new_P1_U2722 = ~new_P1_U4159 | ~new_P1_U4192;
  assign new_P1_U2723 = new_P1_U7236 & new_P1_U7083;
  assign new_P1_U2724 = new_P1_U7253 & new_P1_U7083;
  assign new_P1_U2725 = new_P1_U7270 & new_P1_U7083;
  assign new_P1_U2726 = new_P1_U7620 & new_P1_U7083;
  assign new_P1_U2727 = new_P1_U7302 & new_P1_U7083;
  assign new_P1_U2728 = new_P1_U7319 & new_P1_U7083;
  assign new_P1_U2729 = new_P1_U7336 & new_P1_U7083;
  assign new_P1_U2730 = new_P1_U7353 & new_P1_U7083;
  assign new_P1_U2731 = ~new_P1_U2606 | ~new_P1_U7354;
  assign new_P1_U2732 = new_P1_U7083 & new_P1_U7082;
  assign new_P1_U2733 = new_P1_U7114 & new_P1_U7083;
  assign new_P1_U2734 = new_P1_U7131 & new_P1_U7083;
  assign new_P1_U2735 = new_P1_U7618 & new_P1_U7083;
  assign new_P1_U2736 = new_P1_U7163 & new_P1_U7083;
  assign new_P1_U2737 = new_P1_U7180 & new_P1_U7083;
  assign new_P1_U2738 = new_P1_U7197 & new_P1_U7083;
  assign new_P1_U2739 = new_P1_U7214 & new_P1_U7083;
  assign new_P1_U2740 = P1_INSTQUEUERD_ADDR_REG_4_ & new_P1_U7063;
  assign new_P1_U2741 = ~new_P1_U4078 | ~new_P1_U7096;
  assign new_P1_U2742 = new_P1_U7492 & new_P1_U7491;
  assign new_P1_U2743 = new_P1_U7506 & new_P1_U7470;
  assign new_P1_U2744 = new_P1_U7479 & new_P1_U7478;
  assign new_P1_U2745 = ~new_P1_U7048 | ~new_P1_U7047;
  assign new_P1_U2746 = ~new_P1_U7050 | ~new_P1_U7049;
  assign new_P1_U2747 = ~new_P1_U7052 | ~new_P1_U7051;
  assign new_P1_U2748 = ~new_P1_U7616 | ~new_P1_U7053;
  assign new_P1_U2749 = ~new_P1_U7055 | ~new_P1_U7054;
  assign new_P1_U2750 = ~new_P1_U7057 | ~new_P1_U7056;
  assign new_P1_U2751 = ~new_P1_U4061 | ~new_P1_U7058;
  assign new_P1_U2752 = ~new_P1_U7061 | ~new_P1_U4062 | ~new_P1_U7060;
  assign new_P1_U2753 = new_P1_U6957 & new_P1_U6909;
  assign new_P1_U2754 = new_P1_U6974 & new_P1_U6909;
  assign new_P1_U2755 = new_P1_U6991 & new_P1_U6909;
  assign new_P1_U2756 = new_P1_U7615 & new_P1_U6909;
  assign new_P1_U2757 = new_P1_U7023 & new_P1_U6909;
  assign new_P1_U2758 = new_P1_U7040 & new_P1_U6909;
  assign new_P1_U2759 = new_P1_U6909 & new_P1_U6908;
  assign new_P1_U2760 = new_P1_U6926 & new_P1_U6909;
  assign new_P1_U2761 = ~new_P1_U6928 | ~new_P1_U6927;
  assign new_P1_U2762 = ~new_P1_U6930 | ~new_P1_U6929;
  assign new_P1_U2763 = ~new_P1_U6932 | ~new_P1_U6931;
  assign new_P1_U2764 = ~new_P1_U6934 | ~new_P1_U6933;
  assign new_P1_U2765 = ~new_P1_U6937 | ~new_P1_U6936 | ~new_P1_U6935;
  assign new_P1_U2766 = ~new_P1_U6940 | ~new_P1_U6939 | ~new_P1_U6938;
  assign new_P1_U2767 = ~new_P1_U7042 | ~new_P1_U7043 | ~new_P1_U7041;
  assign new_P1_U2768 = ~new_P1_U7045 | ~new_P1_U7046 | ~new_P1_U7044;
  assign new_P1_U2769 = new_P1_R2144_U145 & new_P1_U4159;
  assign new_P1_U2770 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2771 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2772 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2773 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2774 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2775 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2776 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2777 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2778 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2779 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2780 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2781 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2782 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2783 = new_P1_U4159 & new_P1_R2144_U145;
  assign new_P1_U2784 = new_P1_U4159 & new_P1_R2144_U11;
  assign new_P1_U2785 = new_P1_U4159 & new_P1_R2144_U37;
  assign new_P1_U2786 = new_P1_U4159 & new_P1_R2144_U38;
  assign new_P1_U2787 = new_P1_U4159 & new_P1_R2144_U39;
  assign new_P1_U2788 = new_P1_U4159 & new_P1_R2144_U40;
  assign new_P1_U2789 = new_P1_U4159 & new_P1_R2144_U41;
  assign new_P1_U2790 = new_P1_U4159 & new_P1_R2144_U42;
  assign new_P1_U2791 = new_P1_U4159 & new_P1_R2144_U30;
  assign new_P1_U2792 = ~new_P1_U6872 | ~new_P1_U6871;
  assign new_P1_U2793 = ~new_P1_U6874 | ~new_P1_U6873;
  assign new_P1_U2794 = ~new_P1_U6876 | ~new_P1_U6875;
  assign new_P1_U2795 = ~new_P1_U6878 | ~new_P1_U6877;
  assign new_P1_U2796 = ~new_P1_U6880 | ~new_P1_U6879;
  assign new_P1_U2797 = ~new_P1_U6882 | ~new_P1_U6881;
  assign new_P1_U2798 = ~new_P1_U6883 | ~new_P1_U6884 | ~new_P1_U6885;
  assign new_P1_U2799 = ~new_P1_U6886 | ~new_P1_U4028 | ~new_P1_U6887;
  assign new_P1_U2800 = ~new_P1_U6889 | ~new_P1_U6890 | ~new_P1_U6891;
  assign n7283 = ~new_P1_U7498 | ~new_P1_U6617 | ~new_P1_U3432;
  assign n7274 = ~new_P1_U7650 | ~new_P1_U6613;
  assign n7269 = ~new_P1_U6612 | ~new_P1_U6611;
  assign n7259 = ~new_P1_U4243 | ~new_P1_U7769 | ~new_P1_U7768;
  assign n7249 = ~new_P1_U4243 | ~new_P1_U7765 | ~new_P1_U7764;
  assign n7239 = ~new_P1_U6601 | ~new_P1_U4248;
  assign n7224 = ~new_P1_U4240 | ~new_P1_U7757 | ~new_P1_U7756;
  assign n7214 = ~new_P1_U4240 | ~new_P1_U7747 | ~new_P1_U7746;
  assign n7209 = ~new_P1_U6595 | ~new_P1_U6591 | ~new_P1_U3949 | ~new_P1_U6593 | ~new_P1_U3948;
  assign n7204 = ~new_P1_U6588 | ~new_P1_U6584 | ~new_P1_U3947 | ~new_P1_U6586 | ~new_P1_U3946;
  assign n7199 = ~new_P1_U6581 | ~new_P1_U6577 | ~new_P1_U3945 | ~new_P1_U6579 | ~new_P1_U3944;
  assign n7194 = ~new_P1_U6574 | ~new_P1_U6570 | ~new_P1_U3943 | ~new_P1_U6572 | ~new_P1_U3942;
  assign n7189 = ~new_P1_U6567 | ~new_P1_U6563 | ~new_P1_U3941 | ~new_P1_U6565 | ~new_P1_U3940;
  assign n7184 = ~new_P1_U6560 | ~new_P1_U6556 | ~new_P1_U3939 | ~new_P1_U6558 | ~new_P1_U3938;
  assign n7179 = ~new_P1_U6553 | ~new_P1_U6549 | ~new_P1_U3937 | ~new_P1_U6551 | ~new_P1_U3936;
  assign n7174 = ~new_P1_U6546 | ~new_P1_U6542 | ~new_P1_U3935 | ~new_P1_U6544 | ~new_P1_U3934;
  assign n7169 = ~new_P1_U6539 | ~new_P1_U6535 | ~new_P1_U3933 | ~new_P1_U6537 | ~new_P1_U3932;
  assign n7164 = ~new_P1_U6532 | ~new_P1_U6528 | ~new_P1_U3931 | ~new_P1_U6530 | ~new_P1_U3930;
  assign n7159 = ~new_P1_U6525 | ~new_P1_U6521 | ~new_P1_U3929 | ~new_P1_U6523 | ~new_P1_U3928;
  assign n7154 = ~new_P1_U6518 | ~new_P1_U6514 | ~new_P1_U3927 | ~new_P1_U6516 | ~new_P1_U3926;
  assign n7149 = ~new_P1_U6511 | ~new_P1_U6507 | ~new_P1_U3925 | ~new_P1_U3924 | ~new_P1_U6509;
  assign n7144 = ~new_P1_U6504 | ~new_P1_U6500 | ~new_P1_U3923 | ~new_P1_U3922 | ~new_P1_U6502;
  assign n7139 = ~new_P1_U6497 | ~new_P1_U6493 | ~new_P1_U3921 | ~new_P1_U3920 | ~new_P1_U6495;
  assign n7134 = ~new_P1_U6490 | ~new_P1_U3918 | ~new_P1_U3919 | ~new_P1_U6488 | ~new_P1_U6487;
  assign n7129 = ~new_P1_U6483 | ~new_P1_U3916 | ~new_P1_U3917 | ~new_P1_U6481 | ~new_P1_U6480;
  assign n7124 = ~new_P1_U6476 | ~new_P1_U6473 | ~new_P1_U3914 | ~new_P1_U3915 | ~new_P1_U6474;
  assign n7119 = ~new_P1_U6469 | ~new_P1_U6466 | ~new_P1_U3912 | ~new_P1_U3913 | ~new_P1_U6467;
  assign n7114 = ~new_P1_U6462 | ~new_P1_U6459 | ~new_P1_U3910 | ~new_P1_U3911 | ~new_P1_U6460;
  assign n7109 = ~new_P1_U6455 | ~new_P1_U6452 | ~new_P1_U3908 | ~new_P1_U3909 | ~new_P1_U6453;
  assign n7104 = ~new_P1_U6448 | ~new_P1_U6445 | ~new_P1_U3906 | ~new_P1_U3907 | ~new_P1_U6446;
  assign n7099 = ~new_P1_U6441 | ~new_P1_U6438 | ~new_P1_U3904 | ~new_P1_U3905 | ~new_P1_U6439;
  assign n7094 = ~new_P1_U6434 | ~new_P1_U6431 | ~new_P1_U3902 | ~new_P1_U3903 | ~new_P1_U6432;
  assign n7089 = ~new_P1_U6427 | ~new_P1_U6424 | ~new_P1_U3900 | ~new_P1_U3901 | ~new_P1_U6425;
  assign n7084 = ~new_P1_U6420 | ~new_P1_U6417 | ~new_P1_U3898 | ~new_P1_U3899 | ~new_P1_U6418;
  assign n7079 = ~new_P1_U3897 | ~new_P1_U6410 | ~new_P1_U3896 | ~new_P1_U6409;
  assign n7074 = ~new_P1_U6402 | ~new_P1_U6403 | ~new_P1_U3895 | ~new_P1_U3894 | ~new_P1_U6401;
  assign n7069 = ~new_P1_U3893 | ~new_P1_U6394 | ~new_P1_U6393 | ~new_P1_U6392;
  assign n7064 = ~new_P1_U3892 | ~new_P1_U6386 | ~new_P1_U6385 | ~new_P1_U6384;
  assign n7059 = ~new_P1_U3891 | ~new_P1_U6378 | ~new_P1_U6377 | ~new_P1_U6376;
  assign n7054 = ~new_P1_U3890 | ~new_P1_U6370 | ~new_P1_U6369 | ~new_P1_U6368;
  assign n7049 = ~new_P1_U6359 | ~new_P1_U6358;
  assign n7044 = ~new_P1_U6355 | ~new_P1_U6356 | ~new_P1_U6357;
  assign n7039 = ~new_P1_U6352 | ~new_P1_U6353 | ~new_P1_U6354;
  assign n7034 = ~new_P1_U6349 | ~new_P1_U6350 | ~new_P1_U6351;
  assign n7029 = ~new_P1_U6346 | ~new_P1_U6347 | ~new_P1_U6348;
  assign n7024 = ~new_P1_U6343 | ~new_P1_U6344 | ~new_P1_U6345;
  assign n7019 = ~new_P1_U6340 | ~new_P1_U6341 | ~new_P1_U6342;
  assign n7014 = ~new_P1_U6337 | ~new_P1_U6338 | ~new_P1_U6339;
  assign n7009 = ~new_P1_U6334 | ~new_P1_U6335 | ~new_P1_U6336;
  assign n7004 = ~new_P1_U6331 | ~new_P1_U6332 | ~new_P1_U6333;
  assign n6999 = ~new_P1_U6328 | ~new_P1_U6329 | ~new_P1_U6330;
  assign n6994 = ~new_P1_U6325 | ~new_P1_U6326 | ~new_P1_U6327;
  assign n6989 = ~new_P1_U6322 | ~new_P1_U6323 | ~new_P1_U6324;
  assign n6984 = ~new_P1_U6319 | ~new_P1_U6320 | ~new_P1_U6321;
  assign n6979 = ~new_P1_U6316 | ~new_P1_U6317 | ~new_P1_U6318;
  assign n6974 = ~new_P1_U6313 | ~new_P1_U6314 | ~new_P1_U6315;
  assign n6969 = ~new_P1_U6310 | ~new_P1_U6311 | ~new_P1_U6312;
  assign n6964 = ~new_P1_U6307 | ~new_P1_U6308 | ~new_P1_U6309;
  assign n6959 = ~new_P1_U6304 | ~new_P1_U6305 | ~new_P1_U6306;
  assign n6954 = ~new_P1_U6301 | ~new_P1_U6302 | ~new_P1_U6303;
  assign n6949 = ~new_P1_U6298 | ~new_P1_U6299 | ~new_P1_U6300;
  assign n6944 = ~new_P1_U6295 | ~new_P1_U6296 | ~new_P1_U6297;
  assign n6939 = ~new_P1_U6292 | ~new_P1_U6293 | ~new_P1_U6294;
  assign n6934 = ~new_P1_U6289 | ~new_P1_U6290 | ~new_P1_U6291;
  assign n6929 = ~new_P1_U6286 | ~new_P1_U6287 | ~new_P1_U6288;
  assign n6924 = ~new_P1_U6283 | ~new_P1_U6284 | ~new_P1_U6285;
  assign n6919 = ~new_P1_U6280 | ~new_P1_U6281 | ~new_P1_U6282;
  assign n6914 = ~new_P1_U6277 | ~new_P1_U6278 | ~new_P1_U6279;
  assign n6909 = ~new_P1_U6274 | ~new_P1_U6275 | ~new_P1_U6276;
  assign n6904 = ~new_P1_U6271 | ~new_P1_U6272 | ~new_P1_U6273;
  assign n6899 = ~new_P1_U6268 | ~new_P1_U6269 | ~new_P1_U6270;
  assign n6894 = ~new_P1_U6267 | ~new_P1_U6266 | ~new_P1_U6265;
  assign n6889 = ~new_P1_U4176 | ~new_P1_U6262;
  assign n6884 = ~new_P1_U6260 | ~new_P1_U6261 | ~new_P1_U6259 | ~new_P1_U6258;
  assign n6879 = ~new_P1_U6256 | ~new_P1_U6257 | ~new_P1_U6255 | ~new_P1_U6254;
  assign n6874 = ~new_P1_U6252 | ~new_P1_U6253 | ~new_P1_U6251 | ~new_P1_U6250;
  assign n6869 = ~new_P1_U6248 | ~new_P1_U6249 | ~new_P1_U6247 | ~new_P1_U6246;
  assign n6864 = ~new_P1_U6244 | ~new_P1_U6245 | ~new_P1_U6243 | ~new_P1_U6242;
  assign n6859 = ~new_P1_U6240 | ~new_P1_U6241 | ~new_P1_U6239 | ~new_P1_U6238;
  assign n6854 = ~new_P1_U6236 | ~new_P1_U6237 | ~new_P1_U6235 | ~new_P1_U6234;
  assign n6849 = ~new_P1_U6232 | ~new_P1_U6233 | ~new_P1_U6231 | ~new_P1_U6230;
  assign n6844 = ~new_P1_U6228 | ~new_P1_U6229 | ~new_P1_U6227 | ~new_P1_U6226;
  assign n6839 = ~new_P1_U6224 | ~new_P1_U6225 | ~new_P1_U6223 | ~new_P1_U6222;
  assign n6834 = ~new_P1_U6220 | ~new_P1_U6221 | ~new_P1_U6219 | ~new_P1_U6218;
  assign n6829 = ~new_P1_U6216 | ~new_P1_U6217 | ~new_P1_U6215 | ~new_P1_U6214;
  assign n6824 = ~new_P1_U6212 | ~new_P1_U6213 | ~new_P1_U6211 | ~new_P1_U6210;
  assign n6819 = ~new_P1_U6208 | ~new_P1_U6209 | ~new_P1_U6207 | ~new_P1_U6206;
  assign n6814 = ~new_P1_U6204 | ~new_P1_U6205 | ~new_P1_U6203 | ~new_P1_U6202;
  assign n6809 = ~new_P1_U6200 | ~new_P1_U6201 | ~new_P1_U6199;
  assign n6804 = ~new_P1_U6197 | ~new_P1_U6198 | ~new_P1_U6196;
  assign n6799 = ~new_P1_U6194 | ~new_P1_U6195 | ~new_P1_U6193;
  assign n6794 = ~new_P1_U6191 | ~new_P1_U6192 | ~new_P1_U6190;
  assign n6789 = ~new_P1_U6188 | ~new_P1_U6189 | ~new_P1_U6187;
  assign n6784 = ~new_P1_U6185 | ~new_P1_U6186 | ~new_P1_U6184;
  assign n6779 = ~new_P1_U6182 | ~new_P1_U6183 | ~new_P1_U6181;
  assign n6774 = ~new_P1_U6179 | ~new_P1_U6180 | ~new_P1_U6178;
  assign n6769 = ~new_P1_U6176 | ~new_P1_U6177 | ~new_P1_U6175;
  assign n6764 = ~new_P1_U6173 | ~new_P1_U6174 | ~new_P1_U6172;
  assign n6759 = ~new_P1_U6170 | ~new_P1_U6171 | ~new_P1_U6169;
  assign n6754 = ~new_P1_U6167 | ~new_P1_U6168 | ~new_P1_U6166;
  assign n6749 = ~new_P1_U6164 | ~new_P1_U6165 | ~new_P1_U6163;
  assign n6744 = ~new_P1_U6161 | ~new_P1_U6162 | ~new_P1_U6160;
  assign n6739 = ~new_P1_U6159 | ~new_P1_U6158 | ~new_P1_U6157;
  assign n6734 = ~new_P1_U6156 | ~new_P1_U6155 | ~new_P1_U6154;
  assign n6729 = P1_DATAO_REG_31_ & new_P1_U6055;
  assign n6724 = ~new_P1_U3882 | ~new_P1_U6146;
  assign n6719 = ~new_P1_U3881 | ~new_P1_U6143;
  assign n6714 = ~new_P1_U3880 | ~new_P1_U6140;
  assign n6709 = ~new_P1_U3879 | ~new_P1_U6137;
  assign n6704 = ~new_P1_U3878 | ~new_P1_U6134;
  assign n6699 = ~new_P1_U3877 | ~new_P1_U6131;
  assign n6694 = ~new_P1_U3876 | ~new_P1_U6128;
  assign n6689 = ~new_P1_U3875 | ~new_P1_U6125;
  assign n6684 = ~new_P1_U3874 | ~new_P1_U6122;
  assign n6679 = ~new_P1_U3873 | ~new_P1_U6119;
  assign n6674 = ~new_P1_U3872 | ~new_P1_U6116;
  assign n6669 = ~new_P1_U3871 | ~new_P1_U6113;
  assign n6664 = ~new_P1_U3870 | ~new_P1_U6110;
  assign n6659 = ~new_P1_U3869 | ~new_P1_U6107;
  assign n6654 = ~new_P1_U3868 | ~new_P1_U6104;
  assign n6649 = ~new_P1_U6103 | ~new_P1_U6102 | ~new_P1_U6101;
  assign n6644 = ~new_P1_U6100 | ~new_P1_U6099 | ~new_P1_U6098;
  assign n6639 = ~new_P1_U6097 | ~new_P1_U6096 | ~new_P1_U6095;
  assign n6634 = ~new_P1_U6094 | ~new_P1_U6093 | ~new_P1_U6092;
  assign n6629 = ~new_P1_U6091 | ~new_P1_U6090 | ~new_P1_U6089;
  assign n6624 = ~new_P1_U6088 | ~new_P1_U6087 | ~new_P1_U6086;
  assign n6619 = ~new_P1_U6085 | ~new_P1_U6084 | ~new_P1_U6083;
  assign n6614 = ~new_P1_U6082 | ~new_P1_U6081 | ~new_P1_U6080;
  assign n6609 = ~new_P1_U6079 | ~new_P1_U6078 | ~new_P1_U6077;
  assign n6604 = ~new_P1_U6076 | ~new_P1_U6075 | ~new_P1_U6074;
  assign n6599 = ~new_P1_U6073 | ~new_P1_U6072 | ~new_P1_U6071;
  assign n6594 = ~new_P1_U6070 | ~new_P1_U6069 | ~new_P1_U6068;
  assign n6589 = ~new_P1_U6067 | ~new_P1_U6066 | ~new_P1_U6065;
  assign n6584 = ~new_P1_U6064 | ~new_P1_U6063 | ~new_P1_U6062;
  assign n6579 = ~new_P1_U6061 | ~new_P1_U6060 | ~new_P1_U6059;
  assign n6574 = ~new_P1_U6058 | ~new_P1_U6057 | ~new_P1_U6056;
  assign n6569 = ~new_P1_U7540 | ~new_P1_U7542;
  assign n6564 = ~new_P1_U7539 | ~new_P1_U7544;
  assign n6559 = ~new_P1_U7538 | ~new_P1_U7546;
  assign n6554 = ~new_P1_U7537 | ~new_P1_U7548;
  assign n6549 = ~new_P1_U7536 | ~new_P1_U7550;
  assign n6544 = ~new_P1_U7535 | ~new_P1_U7552;
  assign n6539 = ~new_P1_U7534 | ~new_P1_U7554;
  assign n6534 = ~new_P1_U7533 | ~new_P1_U7556;
  assign n6529 = ~new_P1_U7532 | ~new_P1_U7558;
  assign n6524 = ~new_P1_U7531 | ~new_P1_U7560;
  assign n6519 = ~new_P1_U7530 | ~new_P1_U7562;
  assign n6514 = ~new_P1_U7529 | ~new_P1_U7564;
  assign n6509 = ~new_P1_U7528 | ~new_P1_U7566;
  assign n6504 = ~new_P1_U7527 | ~new_P1_U7568;
  assign n6499 = ~new_P1_U7526 | ~new_P1_U7570;
  assign n6494 = ~new_P1_U7525 | ~new_P1_U7572;
  assign n6489 = ~new_P1_U7524 | ~new_P1_U7574;
  assign n6484 = ~new_P1_U7523 | ~new_P1_U7576;
  assign n6479 = ~new_P1_U7522 | ~new_P1_U7578;
  assign n6474 = ~new_P1_U7521 | ~new_P1_U7580;
  assign n6469 = ~new_P1_U7520 | ~new_P1_U7582;
  assign n6464 = ~new_P1_U7519 | ~new_P1_U7584;
  assign n6459 = ~new_P1_U7518 | ~new_P1_U7586;
  assign n6454 = ~new_P1_U7517 | ~new_P1_U7588;
  assign n6449 = ~new_P1_U7516 | ~new_P1_U7590;
  assign n6444 = ~new_P1_U7515 | ~new_P1_U7592;
  assign n6439 = ~new_P1_U7514 | ~new_P1_U7594;
  assign n6434 = ~new_P1_U7513 | ~new_P1_U7596;
  assign n6429 = ~new_P1_U7512 | ~new_P1_U7598;
  assign n6424 = ~new_P1_U7511 | ~new_P1_U7600;
  assign n6419 = ~new_P1_U7510 | ~new_P1_U7602;
  assign n6414 = ~new_P1_U5957 | ~new_P1_U5955 | ~new_P1_U5958 | ~new_P1_U5956 | ~new_P1_U5954;
  assign n6409 = ~new_P1_U5952 | ~new_P1_U5950 | ~new_P1_U5953 | ~new_P1_U5951 | ~new_P1_U5949;
  assign n6404 = ~new_P1_U5947 | ~new_P1_U5945 | ~new_P1_U5948 | ~new_P1_U5946 | ~new_P1_U5944;
  assign n6399 = ~new_P1_U5942 | ~new_P1_U5940 | ~new_P1_U5943 | ~new_P1_U5941 | ~new_P1_U5939;
  assign n6394 = ~new_P1_U5937 | ~new_P1_U5935 | ~new_P1_U5938 | ~new_P1_U5936 | ~new_P1_U5934;
  assign n6389 = ~new_P1_U5932 | ~new_P1_U5930 | ~new_P1_U5933 | ~new_P1_U5931 | ~new_P1_U5929;
  assign n6384 = ~new_P1_U5927 | ~new_P1_U5925 | ~new_P1_U5928 | ~new_P1_U5926 | ~new_P1_U5924;
  assign n6379 = ~new_P1_U5922 | ~new_P1_U5920 | ~new_P1_U5923 | ~new_P1_U5921 | ~new_P1_U5919;
  assign n6374 = ~new_P1_U5917 | ~new_P1_U5915 | ~new_P1_U5918 | ~new_P1_U5916 | ~new_P1_U5914;
  assign n6369 = ~new_P1_U5912 | ~new_P1_U5910 | ~new_P1_U5913 | ~new_P1_U5911 | ~new_P1_U5909;
  assign n6364 = ~new_P1_U5907 | ~new_P1_U5905 | ~new_P1_U5908 | ~new_P1_U5906 | ~new_P1_U5904;
  assign n6359 = ~new_P1_U5902 | ~new_P1_U5900 | ~new_P1_U5903 | ~new_P1_U5901 | ~new_P1_U5899;
  assign n6354 = ~new_P1_U5897 | ~new_P1_U5895 | ~new_P1_U5898 | ~new_P1_U5896 | ~new_P1_U5894;
  assign n6349 = ~new_P1_U5892 | ~new_P1_U5890 | ~new_P1_U5893 | ~new_P1_U5891 | ~new_P1_U5889;
  assign n6344 = ~new_P1_U5887 | ~new_P1_U5885 | ~new_P1_U5888 | ~new_P1_U5886 | ~new_P1_U5884;
  assign n6339 = ~new_P1_U5882 | ~new_P1_U5880 | ~new_P1_U5883 | ~new_P1_U5881 | ~new_P1_U5879;
  assign n6334 = ~new_P1_U5877 | ~new_P1_U5875 | ~new_P1_U5878 | ~new_P1_U5876 | ~new_P1_U5874;
  assign n6329 = ~new_P1_U5872 | ~new_P1_U5870 | ~new_P1_U5873 | ~new_P1_U5871 | ~new_P1_U5869;
  assign n6324 = ~new_P1_U5867 | ~new_P1_U5865 | ~new_P1_U5868 | ~new_P1_U5866 | ~new_P1_U5864;
  assign n6319 = ~new_P1_U5862 | ~new_P1_U5860 | ~new_P1_U5863 | ~new_P1_U5861 | ~new_P1_U5859;
  assign n6314 = ~new_P1_U5857 | ~new_P1_U5855 | ~new_P1_U5858 | ~new_P1_U5856 | ~new_P1_U5854;
  assign n6309 = ~new_P1_U5852 | ~new_P1_U5850 | ~new_P1_U5853 | ~new_P1_U5851 | ~new_P1_U5849;
  assign n6304 = ~new_P1_U5847 | ~new_P1_U5845 | ~new_P1_U5848 | ~new_P1_U5846 | ~new_P1_U5844;
  assign n6299 = ~new_P1_U5842 | ~new_P1_U5840 | ~new_P1_U5843 | ~new_P1_U5841 | ~new_P1_U5839;
  assign n6294 = ~new_P1_U5837 | ~new_P1_U5838 | ~new_P1_U5835 | ~new_P1_U5836 | ~new_P1_U5834;
  assign n6289 = ~new_P1_U5832 | ~new_P1_U5833 | ~new_P1_U5830 | ~new_P1_U5831 | ~new_P1_U5829;
  assign n6284 = ~new_P1_U5827 | ~new_P1_U5828 | ~new_P1_U5825 | ~new_P1_U5826 | ~new_P1_U5824;
  assign n6279 = ~new_P1_U5822 | ~new_P1_U5823 | ~new_P1_U5820 | ~new_P1_U5821 | ~new_P1_U5819;
  assign n6274 = ~new_P1_U5817 | ~new_P1_U5818 | ~new_P1_U5815 | ~new_P1_U5816 | ~new_P1_U5814;
  assign n6269 = ~new_P1_U5812 | ~new_P1_U5813 | ~new_P1_U5810 | ~new_P1_U5811 | ~new_P1_U5809;
  assign n6264 = ~new_P1_U5807 | ~new_P1_U5808 | ~new_P1_U5806 | ~new_P1_U5805 | ~new_P1_U5804;
  assign n6259 = ~new_P1_U5802 | ~new_P1_U5803 | ~new_P1_U5801 | ~new_P1_U5800 | ~new_P1_U5799;
  assign n6254 = ~new_P1_U5789 | ~new_P1_U5787 | ~new_P1_U3861 | ~new_P1_U3859;
  assign n6249 = ~new_P1_U5782 | ~new_P1_U5780 | ~new_P1_U3858 | ~new_P1_U3856;
  assign n6244 = ~new_P1_U5775 | ~new_P1_U5773 | ~new_P1_U3855 | ~new_P1_U3853;
  assign n6239 = ~new_P1_U5768 | ~new_P1_U5766 | ~new_P1_U3852 | ~new_P1_U3850;
  assign n6234 = ~new_P1_U5761 | ~new_P1_U5759 | ~new_P1_U3849 | ~new_P1_U3847;
  assign n6229 = ~new_P1_U5754 | ~new_P1_U5752 | ~new_P1_U3846 | ~new_P1_U3844;
  assign n6224 = ~new_P1_U5747 | ~new_P1_U5745 | ~new_P1_U3843 | ~new_P1_U3841;
  assign n6219 = ~new_P1_U5740 | ~new_P1_U5738 | ~new_P1_U3840 | ~new_P1_U3838;
  assign n6214 = ~new_P1_U5733 | ~new_P1_U5731 | ~new_P1_U3837 | ~new_P1_U3835;
  assign n6209 = ~new_P1_U5726 | ~new_P1_U5724 | ~new_P1_U3834 | ~new_P1_U3832;
  assign n6204 = ~new_P1_U5719 | ~new_P1_U5717 | ~new_P1_U3831 | ~new_P1_U3829;
  assign n6199 = ~new_P1_U5712 | ~new_P1_U5710 | ~new_P1_U3828 | ~new_P1_U3826;
  assign n6194 = ~new_P1_U5705 | ~new_P1_U5703 | ~new_P1_U3825 | ~new_P1_U3823;
  assign n6189 = ~new_P1_U5698 | ~new_P1_U5696 | ~new_P1_U3822 | ~new_P1_U3820;
  assign n6184 = ~new_P1_U5691 | ~new_P1_U5689 | ~new_P1_U3819 | ~new_P1_U3817;
  assign n6179 = ~new_P1_U5684 | ~new_P1_U5682 | ~new_P1_U3816 | ~new_P1_U3814;
  assign n6174 = ~new_P1_U5677 | ~new_P1_U5675 | ~new_P1_U3813 | ~new_P1_U3811;
  assign n6169 = ~new_P1_U5670 | ~new_P1_U5668 | ~new_P1_U3810 | ~new_P1_U3808;
  assign n6164 = ~new_P1_U5663 | ~new_P1_U5661 | ~new_P1_U3807 | ~new_P1_U3805;
  assign n6159 = ~new_P1_U5656 | ~new_P1_U3802 | ~new_P1_U3804;
  assign n6154 = ~new_P1_U5649 | ~new_P1_U3799 | ~new_P1_U3801;
  assign n6149 = ~new_P1_U5642 | ~new_P1_U3796 | ~new_P1_U3798;
  assign n6144 = ~new_P1_U5635 | ~new_P1_U3793 | ~new_P1_U3795;
  assign n6139 = ~new_P1_U5628 | ~new_P1_U3790 | ~new_P1_U3792;
  assign n6134 = ~new_P1_U5621 | ~new_P1_U3787 | ~new_P1_U3789;
  assign n6129 = ~new_P1_U5614 | ~new_P1_U3784 | ~new_P1_U3786;
  assign n6124 = ~new_P1_U5607 | ~new_P1_U3781 | ~new_P1_U3783;
  assign n6119 = ~new_P1_U5600 | ~new_P1_U3778 | ~new_P1_U3780;
  assign n6114 = ~new_P1_U3775 | ~new_P1_U3776;
  assign n6109 = ~new_P1_U3774 | ~new_P1_U3772 | ~new_P1_U3771;
  assign n6104 = ~new_P1_U3770 | ~new_P1_U3768 | ~new_P1_U3767;
  assign n6099 = ~new_P1_U3766 | ~new_P1_U3764 | ~new_P1_U3763;
  assign n6074 = P1_INSTQUEUEWR_ADDR_REG_4_ & new_P1_U5537;
  assign n6044 = ~new_P1_U3730 | ~new_P1_U5460 | ~new_P1_U5459;
  assign n6039 = ~new_P1_U3729 | ~new_P1_U5455 | ~new_P1_U5454;
  assign n6034 = ~new_P1_U3728 | ~new_P1_U5450 | ~new_P1_U5449;
  assign n6029 = ~new_P1_U3727 | ~new_P1_U5445 | ~new_P1_U5444;
  assign n6024 = ~new_P1_U3726 | ~new_P1_U7612 | ~new_P1_U5440;
  assign n6019 = ~new_P1_U3725 | ~new_P1_U5436 | ~new_P1_U5435;
  assign n6014 = ~new_P1_U3724 | ~new_P1_U5431 | ~new_P1_U5430;
  assign n6009 = ~new_P1_U3723 | ~new_P1_U5426 | ~new_P1_U5425;
  assign n6004 = ~new_P1_U3721 | ~new_P1_U5404 | ~new_P1_U5403;
  assign n5999 = ~new_P1_U3720 | ~new_P1_U5399 | ~new_P1_U5398;
  assign n5994 = ~new_P1_U3719 | ~new_P1_U5394 | ~new_P1_U5393;
  assign n5989 = ~new_P1_U3718 | ~new_P1_U5389 | ~new_P1_U5388;
  assign n5984 = ~new_P1_U3717 | ~new_P1_U5384 | ~new_P1_U5383;
  assign n5979 = ~new_P1_U3716 | ~new_P1_U5379 | ~new_P1_U5378;
  assign n5974 = ~new_P1_U3715 | ~new_P1_U5374 | ~new_P1_U5373;
  assign n5969 = ~new_P1_U3714 | ~new_P1_U5369 | ~new_P1_U5368;
  assign n5964 = ~new_P1_U3712 | ~new_P1_U5346 | ~new_P1_U5345;
  assign n5959 = ~new_P1_U3711 | ~new_P1_U5341 | ~new_P1_U5340;
  assign n5954 = ~new_P1_U3710 | ~new_P1_U5336 | ~new_P1_U5335;
  assign n5949 = ~new_P1_U3709 | ~new_P1_U5331 | ~new_P1_U5330;
  assign n5944 = ~new_P1_U3708 | ~new_P1_U5326 | ~new_P1_U5325;
  assign n5939 = ~new_P1_U3707 | ~new_P1_U5321 | ~new_P1_U5320;
  assign n5934 = ~new_P1_U3706 | ~new_P1_U5316 | ~new_P1_U5315;
  assign n5929 = ~new_P1_U3705 | ~new_P1_U5311 | ~new_P1_U5310;
  assign n5924 = ~new_P1_U3703 | ~new_P1_U5289 | ~new_P1_U5288;
  assign n5919 = ~new_P1_U3702 | ~new_P1_U5284 | ~new_P1_U5283;
  assign n5914 = ~new_P1_U3701 | ~new_P1_U5279 | ~new_P1_U5278;
  assign n5909 = ~new_P1_U3700 | ~new_P1_U5274 | ~new_P1_U5273;
  assign n5904 = ~new_P1_U3699 | ~new_P1_U5269 | ~new_P1_U5268;
  assign n5899 = ~new_P1_U3698 | ~new_P1_U5264 | ~new_P1_U5263;
  assign n5894 = ~new_P1_U3697 | ~new_P1_U5259 | ~new_P1_U5258;
  assign n5889 = ~new_P1_U3696 | ~new_P1_U5254 | ~new_P1_U5253;
  assign n5884 = ~new_P1_U3694 | ~new_P1_U5231 | ~new_P1_U5230;
  assign n5879 = ~new_P1_U3693 | ~new_P1_U5226 | ~new_P1_U5225;
  assign n5874 = ~new_P1_U3692 | ~new_P1_U5221 | ~new_P1_U5220;
  assign n5869 = ~new_P1_U3691 | ~new_P1_U5216 | ~new_P1_U5215;
  assign n5864 = ~new_P1_U3690 | ~new_P1_U5211 | ~new_P1_U5210;
  assign n5859 = ~new_P1_U3689 | ~new_P1_U5206 | ~new_P1_U5205;
  assign n5854 = ~new_P1_U3688 | ~new_P1_U5201 | ~new_P1_U5200;
  assign n5849 = ~new_P1_U3687 | ~new_P1_U5196 | ~new_P1_U5195;
  assign n5844 = ~new_P1_U3685 | ~new_P1_U5174 | ~new_P1_U5173;
  assign n5839 = ~new_P1_U3684 | ~new_P1_U5169 | ~new_P1_U5168;
  assign n5834 = ~new_P1_U3683 | ~new_P1_U5164 | ~new_P1_U5163;
  assign n5829 = ~new_P1_U3682 | ~new_P1_U5159 | ~new_P1_U5158;
  assign n5824 = ~new_P1_U3681 | ~new_P1_U5154 | ~new_P1_U5153;
  assign n5819 = ~new_P1_U3680 | ~new_P1_U5149 | ~new_P1_U5148;
  assign n5814 = ~new_P1_U3679 | ~new_P1_U5144 | ~new_P1_U5143;
  assign n5809 = ~new_P1_U3678 | ~new_P1_U5139 | ~new_P1_U5138;
  assign n5804 = ~new_P1_U3676 | ~new_P1_U5116 | ~new_P1_U5115;
  assign n5799 = ~new_P1_U3675 | ~new_P1_U5111 | ~new_P1_U5110;
  assign n5794 = ~new_P1_U3674 | ~new_P1_U5106 | ~new_P1_U5105;
  assign n5789 = ~new_P1_U3673 | ~new_P1_U5101 | ~new_P1_U5100;
  assign n5784 = ~new_P1_U3672 | ~new_P1_U5096 | ~new_P1_U5095;
  assign n5779 = ~new_P1_U3671 | ~new_P1_U5091 | ~new_P1_U5090;
  assign n5774 = ~new_P1_U3670 | ~new_P1_U5086 | ~new_P1_U5085;
  assign n5769 = ~new_P1_U3669 | ~new_P1_U5081 | ~new_P1_U5080;
  assign n5764 = ~new_P1_U3667 | ~new_P1_U5059 | ~new_P1_U5058;
  assign n5759 = ~new_P1_U3666 | ~new_P1_U5054 | ~new_P1_U5053;
  assign n5754 = ~new_P1_U3665 | ~new_P1_U5049 | ~new_P1_U5048;
  assign n5749 = ~new_P1_U3664 | ~new_P1_U5044 | ~new_P1_U5043;
  assign n5744 = ~new_P1_U3663 | ~new_P1_U5039 | ~new_P1_U5038;
  assign n5739 = ~new_P1_U3662 | ~new_P1_U5034 | ~new_P1_U5033;
  assign n5734 = ~new_P1_U3661 | ~new_P1_U5029 | ~new_P1_U5028;
  assign n5729 = ~new_P1_U3660 | ~new_P1_U5024 | ~new_P1_U5023;
  assign n5724 = ~new_P1_U3658 | ~new_P1_U5003 | ~new_P1_U5002;
  assign n5719 = ~new_P1_U3657 | ~new_P1_U4998 | ~new_P1_U4997;
  assign n5714 = ~new_P1_U3656 | ~new_P1_U4993 | ~new_P1_U4992;
  assign n5709 = ~new_P1_U3655 | ~new_P1_U4988 | ~new_P1_U4987;
  assign n5704 = ~new_P1_U3654 | ~new_P1_U4983 | ~new_P1_U4982;
  assign n5699 = ~new_P1_U3653 | ~new_P1_U4978 | ~new_P1_U4977;
  assign n5694 = ~new_P1_U3652 | ~new_P1_U4973 | ~new_P1_U4972;
  assign n5689 = ~new_P1_U3651 | ~new_P1_U4968 | ~new_P1_U4967;
  assign n5684 = ~new_P1_U3649 | ~new_P1_U4946 | ~new_P1_U4945;
  assign n5679 = ~new_P1_U3648 | ~new_P1_U4941 | ~new_P1_U4940;
  assign n5674 = ~new_P1_U3647 | ~new_P1_U4936 | ~new_P1_U4935;
  assign n5669 = ~new_P1_U3646 | ~new_P1_U4931 | ~new_P1_U4930;
  assign n5664 = ~new_P1_U3645 | ~new_P1_U4926 | ~new_P1_U4925;
  assign n5659 = ~new_P1_U3644 | ~new_P1_U4921 | ~new_P1_U4920;
  assign n5654 = ~new_P1_U3643 | ~new_P1_U4916 | ~new_P1_U4915;
  assign n5649 = ~new_P1_U3642 | ~new_P1_U4911 | ~new_P1_U4910;
  assign n5644 = ~new_P1_U3640 | ~new_P1_U4888 | ~new_P1_U4887;
  assign n5639 = ~new_P1_U3639 | ~new_P1_U4883 | ~new_P1_U4882;
  assign n5634 = ~new_P1_U3638 | ~new_P1_U4878 | ~new_P1_U4877;
  assign n5629 = ~new_P1_U3637 | ~new_P1_U4873 | ~new_P1_U4872;
  assign n5624 = ~new_P1_U3636 | ~new_P1_U4868 | ~new_P1_U4867;
  assign n5619 = ~new_P1_U3635 | ~new_P1_U4863 | ~new_P1_U4862;
  assign n5614 = ~new_P1_U3634 | ~new_P1_U4858 | ~new_P1_U4857;
  assign n5609 = ~new_P1_U3633 | ~new_P1_U4853 | ~new_P1_U4852;
  assign n5604 = ~new_P1_U3631 | ~new_P1_U4831 | ~new_P1_U4830;
  assign n5599 = ~new_P1_U3630 | ~new_P1_U4826 | ~new_P1_U4825;
  assign n5594 = ~new_P1_U3629 | ~new_P1_U4821 | ~new_P1_U4820;
  assign n5589 = ~new_P1_U3628 | ~new_P1_U4816 | ~new_P1_U4815;
  assign n5584 = ~new_P1_U3627 | ~new_P1_U4811 | ~new_P1_U4810;
  assign n5579 = ~new_P1_U3626 | ~new_P1_U4806 | ~new_P1_U4805;
  assign n5574 = ~new_P1_U3625 | ~new_P1_U4801 | ~new_P1_U4800;
  assign n5569 = ~new_P1_U3624 | ~new_P1_U4796 | ~new_P1_U4795;
  assign n5564 = ~new_P1_U3622 | ~new_P1_U4773 | ~new_P1_U4772;
  assign n5559 = ~new_P1_U3621 | ~new_P1_U4768 | ~new_P1_U4767;
  assign n5554 = ~new_P1_U3620 | ~new_P1_U4763 | ~new_P1_U4762;
  assign n5549 = ~new_P1_U3619 | ~new_P1_U4758 | ~new_P1_U4757;
  assign n5544 = ~new_P1_U3618 | ~new_P1_U4753 | ~new_P1_U4752;
  assign n5539 = ~new_P1_U3617 | ~new_P1_U4748 | ~new_P1_U4747;
  assign n5534 = ~new_P1_U3616 | ~new_P1_U4743 | ~new_P1_U4742;
  assign n5529 = ~new_P1_U3615 | ~new_P1_U4738 | ~new_P1_U4737;
  assign n5524 = ~new_P1_U3613 | ~new_P1_U4716 | ~new_P1_U4715;
  assign n5519 = ~new_P1_U3612 | ~new_P1_U4711 | ~new_P1_U4710;
  assign n5514 = ~new_P1_U3611 | ~new_P1_U4706 | ~new_P1_U4705;
  assign n5509 = ~new_P1_U3610 | ~new_P1_U4701 | ~new_P1_U4700;
  assign n5504 = ~new_P1_U3609 | ~new_P1_U4696 | ~new_P1_U4695;
  assign n5499 = ~new_P1_U3608 | ~new_P1_U4691 | ~new_P1_U4690;
  assign n5494 = ~new_P1_U3607 | ~new_P1_U4686 | ~new_P1_U4685;
  assign n5489 = ~new_P1_U3606 | ~new_P1_U4681 | ~new_P1_U4680;
  assign n5484 = ~new_P1_U3604 | ~new_P1_U4657 | ~new_P1_U4656;
  assign n5479 = ~new_P1_U3603 | ~new_P1_U4652 | ~new_P1_U4651;
  assign n5474 = ~new_P1_U3602 | ~new_P1_U4647 | ~new_P1_U4646;
  assign n5469 = ~new_P1_U3601 | ~new_P1_U4642 | ~new_P1_U4641;
  assign n5464 = ~new_P1_U3600 | ~new_P1_U4637 | ~new_P1_U4636;
  assign n5459 = ~new_P1_U3599 | ~new_P1_U4632 | ~new_P1_U4631;
  assign n5454 = ~new_P1_U3598 | ~new_P1_U4627 | ~new_P1_U4626;
  assign n5449 = ~new_P1_U3597 | ~new_P1_U4622 | ~new_P1_U4621;
  assign n5444 = ~new_P1_U3595 | ~new_P1_U4599 | ~new_P1_U4598;
  assign n5439 = ~new_P1_U3594 | ~new_P1_U4594 | ~new_P1_U4593;
  assign n5434 = ~new_P1_U3593 | ~new_P1_U4589 | ~new_P1_U4588;
  assign n5429 = ~new_P1_U3592 | ~new_P1_U4584 | ~new_P1_U4583;
  assign n5424 = ~new_P1_U3591 | ~new_P1_U4579 | ~new_P1_U4578;
  assign n5419 = ~new_P1_U3590 | ~new_P1_U4574 | ~new_P1_U4573;
  assign n5414 = ~new_P1_U3589 | ~new_P1_U4569 | ~new_P1_U4568;
  assign n5409 = ~new_P1_U3588 | ~new_P1_U4564 | ~new_P1_U4563;
  assign n5404 = ~new_P1_U3586 | ~new_P1_U7690 | ~new_P1_U7689;
  assign n5399 = ~new_P1_U4244 | ~new_P1_U4518 | ~new_P1_U4520 | ~new_P1_U4519;
  assign n5394 = ~new_P1_U3582 | ~new_P1_U4516;
  assign n5384 = P1_DATAWIDTH_REG_31_ & new_P1_U7650;
  assign n5379 = P1_DATAWIDTH_REG_30_ & new_P1_U7650;
  assign n5374 = P1_DATAWIDTH_REG_29_ & new_P1_U7650;
  assign n5369 = P1_DATAWIDTH_REG_28_ & new_P1_U7650;
  assign n5364 = P1_DATAWIDTH_REG_27_ & new_P1_U7650;
  assign n5359 = P1_DATAWIDTH_REG_26_ & new_P1_U7650;
  assign n5354 = P1_DATAWIDTH_REG_25_ & new_P1_U7650;
  assign n5349 = P1_DATAWIDTH_REG_24_ & new_P1_U7650;
  assign n5344 = P1_DATAWIDTH_REG_23_ & new_P1_U7650;
  assign n5339 = P1_DATAWIDTH_REG_22_ & new_P1_U7650;
  assign n5334 = P1_DATAWIDTH_REG_21_ & new_P1_U7650;
  assign n5329 = P1_DATAWIDTH_REG_20_ & new_P1_U7650;
  assign n5324 = P1_DATAWIDTH_REG_19_ & new_P1_U7650;
  assign n5319 = P1_DATAWIDTH_REG_18_ & new_P1_U7650;
  assign n5314 = P1_DATAWIDTH_REG_17_ & new_P1_U7650;
  assign n5309 = P1_DATAWIDTH_REG_16_ & new_P1_U7650;
  assign n5304 = P1_DATAWIDTH_REG_15_ & new_P1_U7650;
  assign n5299 = P1_DATAWIDTH_REG_14_ & new_P1_U7650;
  assign n5294 = P1_DATAWIDTH_REG_13_ & new_P1_U7650;
  assign n5289 = P1_DATAWIDTH_REG_12_ & new_P1_U7650;
  assign n5284 = P1_DATAWIDTH_REG_11_ & new_P1_U7650;
  assign n5279 = P1_DATAWIDTH_REG_10_ & new_P1_U7650;
  assign n5274 = P1_DATAWIDTH_REG_9_ & new_P1_U7650;
  assign n5269 = P1_DATAWIDTH_REG_8_ & new_P1_U7650;
  assign n5264 = P1_DATAWIDTH_REG_7_ & new_P1_U7650;
  assign n5259 = P1_DATAWIDTH_REG_6_ & new_P1_U7650;
  assign n5254 = P1_DATAWIDTH_REG_5_ & new_P1_U7650;
  assign n5249 = P1_DATAWIDTH_REG_4_ & new_P1_U7650;
  assign n5244 = P1_DATAWIDTH_REG_3_ & new_P1_U7650;
  assign n5239 = P1_DATAWIDTH_REG_2_ & new_P1_U7650;
  assign n5224 = ~new_P1_U4375 | ~new_P1_U7647 | ~new_P1_U7646;
  assign n5219 = ~new_P1_U3495 | ~new_P1_U7645 | ~new_P1_U7644;
  assign n5214 = ~new_P1_U3494 | ~new_P1_U4369;
  assign n5210 = ~new_P1_U4356 | ~new_P1_U4355 | ~new_P1_U4354;
  assign n5206 = ~new_P1_U4353 | ~new_P1_U4352 | ~new_P1_U4351;
  assign n5202 = ~new_P1_U4350 | ~new_P1_U4349 | ~new_P1_U4348;
  assign n5198 = ~new_P1_U4347 | ~new_P1_U4346 | ~new_P1_U4345;
  assign n5194 = ~new_P1_U4344 | ~new_P1_U4343 | ~new_P1_U4342;
  assign n5190 = ~new_P1_U4341 | ~new_P1_U4340 | ~new_P1_U4339;
  assign n5186 = ~new_P1_U4338 | ~new_P1_U4337 | ~new_P1_U4336;
  assign n5182 = ~new_P1_U4335 | ~new_P1_U4334 | ~new_P1_U4333;
  assign n5178 = ~new_P1_U4332 | ~new_P1_U4331 | ~new_P1_U4330;
  assign n5174 = ~new_P1_U4329 | ~new_P1_U4328 | ~new_P1_U4327;
  assign n5170 = ~new_P1_U4326 | ~new_P1_U4325 | ~new_P1_U4324;
  assign n5166 = ~new_P1_U4323 | ~new_P1_U4322 | ~new_P1_U4321;
  assign n5162 = ~new_P1_U4320 | ~new_P1_U4319 | ~new_P1_U4318;
  assign n5158 = ~new_P1_U4317 | ~new_P1_U4316 | ~new_P1_U4315;
  assign n5154 = ~new_P1_U4314 | ~new_P1_U4313 | ~new_P1_U4312;
  assign n5150 = ~new_P1_U4311 | ~new_P1_U4310 | ~new_P1_U4309;
  assign n5146 = ~new_P1_U4308 | ~new_P1_U4307 | ~new_P1_U4306;
  assign n5142 = ~new_P1_U4305 | ~new_P1_U4304 | ~new_P1_U4303;
  assign n5138 = ~new_P1_U4302 | ~new_P1_U4301 | ~new_P1_U4300;
  assign n5134 = ~new_P1_U4299 | ~new_P1_U4298 | ~new_P1_U4297;
  assign n5130 = ~new_P1_U4296 | ~new_P1_U4295 | ~new_P1_U4294;
  assign n5126 = ~new_P1_U4293 | ~new_P1_U4292 | ~new_P1_U4291;
  assign n5122 = ~new_P1_U4290 | ~new_P1_U4289 | ~new_P1_U4288;
  assign n5118 = ~new_P1_U4287 | ~new_P1_U4286 | ~new_P1_U4285;
  assign n5114 = ~new_P1_U4284 | ~new_P1_U4283 | ~new_P1_U4282;
  assign n5110 = ~new_P1_U4281 | ~new_P1_U4280 | ~new_P1_U4279;
  assign n5106 = ~new_P1_U4278 | ~new_P1_U4277 | ~new_P1_U4276;
  assign n5102 = ~new_P1_U4275 | ~new_P1_U4274 | ~new_P1_U4273;
  assign n5098 = ~new_P1_U4272 | ~new_P1_U4271 | ~new_P1_U4270;
  assign n5094 = ~new_P1_U4269 | ~new_P1_U4268 | ~new_P1_U4267;
  assign new_P1_U3227 = ~new_P1_U3998 | ~new_P1_U3999 | ~new_P1_U4001 | ~new_P1_U4000;
  assign new_P1_U3228 = ~new_P1_U3994 | ~new_P1_U3995 | ~new_P1_U3997 | ~new_P1_U3996;
  assign new_P1_U3229 = ~new_P1_U3990 | ~new_P1_U3991 | ~new_P1_U3993 | ~new_P1_U3992;
  assign new_P1_U3230 = ~new_P1_U3986 | ~new_P1_U3987 | ~new_P1_U3989 | ~new_P1_U3988;
  assign new_P1_U3231 = ~new_P1_U3982 | ~new_P1_U3983 | ~new_P1_U3985 | ~new_P1_U3984;
  assign new_P1_U3232 = ~new_P1_U3978 | ~new_P1_U3979 | ~new_P1_U3981 | ~new_P1_U3980;
  assign new_P1_U3233 = ~new_P1_U3974 | ~new_P1_U3975 | ~new_P1_U3977 | ~new_P1_U3976;
  assign new_P1_U3234 = ~new_P1_U3970 | ~new_P1_U3971 | ~new_P1_U3973 | ~new_P1_U3972;
  assign new_P1_U3235 = ~new_P1_U3329 | ~new_P1_U3323;
  assign new_P1_U3236 = ~new_P1_U2432 | ~new_P1_U3235;
  assign new_P1_U3237 = ~new_P1_U2432 | ~new_P1_U4543;
  assign new_P1_U3238 = ~new_P1_U2434 | ~new_P1_U3235;
  assign new_P1_U3239 = ~new_P1_U2434 | ~new_P1_U4543;
  assign new_P1_U3240 = ~new_P1_U2433 | ~new_P1_U3235;
  assign new_P1_U3241 = ~new_P1_U2433 | ~new_P1_U4543;
  assign new_P1_U3242 = ~new_P1_U2435 | ~new_P1_U3235;
  assign new_P1_U3243 = ~new_P1_U2435 | ~new_P1_U4543;
  assign new_P1_U3244 = ~new_P1_U5463 | ~new_P1_U3391 | ~new_P1_U3394;
  assign new_P1_U3245 = ~new_P1_U7086 | ~new_P1_U5464;
  assign new_P1_U3246 = ~new_P1_U4156 | ~new_P1_U4158 | ~new_P1_U7792 | ~new_P1_U7791;
  assign new_P1_U3247 = ~P1_REQUESTPENDING_REG;
  assign new_P1_U3248 = ~P1_STATE_REG_1_;
  assign new_P1_U3249 = ~P1_STATE_REG_1_ | ~new_P1_U3258;
  assign new_P1_U3250 = ~new_P1_U4221 | ~new_P1_U3251;
  assign new_P1_U3251 = ~P1_STATE_REG_2_;
  assign new_P1_U3252 = ~P1_STATE_REG_2_ | ~new_P1_U4221;
  assign new_P1_U3253 = ~P1_REIP_REG_1_;
  assign new_P1_U3254 = ~P1_STATE_REG_1_ | ~new_P1_U3251;
  assign new_P1_U3255 = P1_STATE_REG_1_ | P1_STATE_REG_2_;
  assign new_P1_U3256 = ~HOLD;
  assign new_P1_U3257 = ~new_U210;
  assign new_P1_U3258 = ~P1_STATE_REG_0_;
  assign new_P1_U3259 = ~P1_STATE_REG_0_ | ~new_P1_U3260;
  assign new_P1_U3260 = ~P1_REQUESTPENDING_REG | ~new_P1_U3256;
  assign new_P1_U3261 = HOLD | P1_REQUESTPENDING_REG;
  assign new_P1_U3262 = ~P1_STATE2_REG_1_;
  assign new_P1_U3263 = ~P1_STATE2_REG_2_;
  assign new_P1_U3264 = ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3265 = ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3266 = ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3267 = ~new_P1_U3270 | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3268 = P1_INSTQUEUERD_ADDR_REG_2_ | P1_INSTQUEUERD_ADDR_REG_0_ | P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3269 = P1_INSTQUEUERD_ADDR_REG_1_ | P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3270 = ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3271 = ~new_P1_U3564 | ~new_P1_U3565 | ~new_P1_U3567 | ~new_P1_U3566;
  assign new_P1_U3272 = ~new_P1_U4496 | ~new_P1_U3258;
  assign new_P1_U3273 = ~new_P1_R2167_U17;
  assign new_P1_U3274 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3270;
  assign new_P1_U3275 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3276 = ~new_P1_U3516 | ~new_P1_U3517 | ~new_P1_U3519 | ~new_P1_U3518;
  assign new_P1_U3277 = ~new_P1_U3536 | ~new_P1_U3537 | ~new_P1_U3538 | ~new_P1_U3539 | ~new_P1_U4170;
  assign new_P1_U3278 = ~new_P1_U3554 | ~new_P1_U3555 | ~new_P1_U3557 | ~new_P1_U3556;
  assign new_P1_U3279 = ~new_P1_U3559 | ~new_P1_U3558;
  assign new_P1_U3280 = P1_STATEBS16_REG | new_U210;
  assign new_P1_U3281 = ~new_P1_R2167_U17 | ~new_P1_U4497;
  assign new_P1_U3282 = ~new_P1_U4477 | ~new_P1_U3284;
  assign new_P1_U3283 = ~new_P1_U3508 | ~new_P1_U3509 | ~new_P1_U3511 | ~new_P1_U3510;
  assign new_P1_U3284 = ~new_P1_U3560 | ~new_P1_U3561 | ~new_P1_U3563 | ~new_P1_U3562;
  assign new_P1_U3285 = ~new_P1_U2473 | ~new_P1_U4501;
  assign new_P1_U3286 = ~new_P1_U2389 | ~new_P1_U3283;
  assign new_P1_U3287 = ~new_P1_U4494 | ~new_P1_U4477;
  assign new_P1_U3288 = ~new_P1_U4249 | ~new_P1_U2447;
  assign new_P1_U3289 = ~new_P1_U3278 | ~new_P1_U4173 | ~new_P1_U4460 | ~new_P1_U3391;
  assign new_P1_U3290 = ~new_P1_U3271 | ~new_P1_U3283;
  assign new_P1_U3291 = ~new_P1_U4190 | ~new_P1_U3284;
  assign new_P1_U3292 = ~new_P1_U4256 | ~new_P1_U2431;
  assign new_P1_U3293 = ~new_P1_LT_563_U6 | ~new_P1_U4225 | ~new_P1_U7626 | ~new_P1_U4178 | ~new_P1_U4509;
  assign new_P1_U3294 = ~P1_STATE2_REG_0_;
  assign new_P1_U3295 = ~P1_STATE2_REG_0_ | ~new_P1_U7604;
  assign new_P1_U3296 = ~P1_STATE2_REG_3_;
  assign new_P1_U3297 = ~P1_STATE2_REG_2_ | ~new_P1_U3262;
  assign new_P1_U3298 = P1_STATE2_REG_2_ | P1_STATE2_REG_1_;
  assign new_P1_U3299 = ~P1_STATE2_REG_3_ | ~new_P1_R2167_U17;
  assign new_P1_U3300 = ~new_P1_U4547 | ~new_P1_U3294;
  assign new_P1_U3301 = ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P1_U3302 = ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P1_U3303 = ~P1_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P1_U3304 = ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P1_U3305 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P1_U3306 = ~new_P1_U4533 | ~new_P1_U2478;
  assign new_P1_U3307 = P1_STATE2_REG_2_ | P1_STATE2_REG_3_;
  assign new_P1_U3308 = ~P1_STATEBS16_REG;
  assign new_P1_U3309 = ~new_P1_R2144_U43;
  assign new_P1_U3310 = ~new_P1_R2144_U50;
  assign new_P1_U3311 = ~new_P1_R2144_U49;
  assign new_P1_U3312 = ~new_P1_R2144_U8;
  assign new_P1_U3313 = ~new_P1_R2144_U50 | ~new_P1_R2144_U43;
  assign new_P1_U3314 = ~new_P1_U3332 | ~new_P1_U3309;
  assign new_P1_U3315 = ~new_P1_U4527 | ~new_P1_U2475;
  assign new_P1_U3316 = ~new_P1_R2182_U25;
  assign new_P1_U3317 = ~new_P1_R2182_U42;
  assign new_P1_U3318 = ~new_P1_R2182_U34;
  assign new_P1_U3319 = ~new_P1_R2182_U33;
  assign new_P1_U3320 = ~new_P1_U4209 | ~new_P1_U3308;
  assign new_P1_U3321 = ~new_P1_U3306 | ~new_P1_U4535;
  assign new_P1_U3322 = ~new_P1_U3306 | ~new_P1_U4544;
  assign new_P1_U3323 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_U3301;
  assign new_P1_U3324 = ~new_P1_U4542 | ~new_P1_U2478;
  assign new_P1_U3325 = ~new_P1_R2144_U50 | ~new_P1_U3309;
  assign new_P1_U3326 = ~new_P1_R2144_U43 | ~new_P1_U3332;
  assign new_P1_U3327 = ~new_P1_U4600 | ~new_P1_U2475;
  assign new_P1_U3328 = ~new_P1_U3324 | ~new_P1_U4603;
  assign new_P1_U3329 = ~P1_INSTQUEUEWR_ADDR_REG_0_ | ~new_P1_U3302;
  assign new_P1_U3330 = ~new_P1_U4541 | ~new_P1_U2478;
  assign new_P1_U3331 = ~new_P1_R2144_U43 | ~new_P1_U3310;
  assign new_P1_U3332 = ~new_P1_U3325 | ~new_P1_U3331;
  assign new_P1_U3333 = ~new_P1_U4526 | ~new_P1_U3309;
  assign new_P1_U3334 = ~new_P1_U4658 | ~new_P1_U2475;
  assign new_P1_U3335 = ~new_P1_U3330 | ~new_P1_U4661;
  assign new_P1_U3336 = ~new_P1_U3330 | ~new_P1_U4663;
  assign new_P1_U3337 = ~new_P1_U2488 | ~new_P1_U2478;
  assign new_P1_U3338 = ~new_P1_U2485 | ~new_P1_U2475;
  assign new_P1_U3339 = ~new_P1_U3337 | ~new_P1_U4719;
  assign new_P1_U3340 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_U3304;
  assign new_P1_U3341 = ~new_P1_U4538 | ~new_P1_U4533;
  assign new_P1_U3342 = ~new_P1_R2144_U8 | ~new_P1_U3311;
  assign new_P1_U3343 = ~new_P1_U2490 | ~new_P1_U4527;
  assign new_P1_U3344 = ~new_P1_U3341 | ~new_P1_U4776;
  assign new_P1_U3345 = ~new_P1_U3341 | ~new_P1_U4778;
  assign new_P1_U3346 = ~new_P1_U4538 | ~new_P1_U4542;
  assign new_P1_U3347 = ~new_P1_U2490 | ~new_P1_U4600;
  assign new_P1_U3348 = ~new_P1_U3346 | ~new_P1_U4834;
  assign new_P1_U3349 = ~new_P1_U4538 | ~new_P1_U4541;
  assign new_P1_U3350 = ~new_P1_U2490 | ~new_P1_U4658;
  assign new_P1_U3351 = ~new_P1_U3349 | ~new_P1_U4891;
  assign new_P1_U3352 = ~new_P1_U3349 | ~new_P1_U4893;
  assign new_P1_U3353 = ~new_P1_U4538 | ~new_P1_U2488;
  assign new_P1_U3354 = ~new_P1_U2490 | ~new_P1_U2485;
  assign new_P1_U3355 = ~new_P1_U3353 | ~new_P1_U4949;
  assign new_P1_U3356 = ~new_P1_U2479 | ~new_P1_U4533;
  assign new_P1_U3357 = ~new_P1_U2474 | ~new_P1_U4528;
  assign new_P1_U3358 = ~new_P1_U3357 | ~new_P1_U3342 | ~new_P1_U4530;
  assign new_P1_U3359 = ~new_P1_U2499 | ~new_P1_U4527;
  assign new_P1_U3360 = ~new_P1_U3356 | ~new_P1_U3340 | ~new_P1_U4539;
  assign new_P1_U3361 = ~new_P1_U3356 | ~new_P1_U5005;
  assign new_P1_U3362 = ~new_P1_U3356 | ~new_P1_U5007;
  assign new_P1_U3363 = ~new_P1_U4542 | ~new_P1_U2479;
  assign new_P1_U3364 = ~new_P1_U2499 | ~new_P1_U4600;
  assign new_P1_U3365 = ~new_P1_U3363 | ~new_P1_U5062;
  assign new_P1_U3366 = ~new_P1_U4541 | ~new_P1_U2479;
  assign new_P1_U3367 = ~new_P1_U2499 | ~new_P1_U4658;
  assign new_P1_U3368 = ~new_P1_U3366 | ~new_P1_U5119;
  assign new_P1_U3369 = ~new_P1_U3366 | ~new_P1_U5121;
  assign new_P1_U3370 = ~new_P1_U2488 | ~new_P1_U2479;
  assign new_P1_U3371 = ~new_P1_U2499 | ~new_P1_U2485;
  assign new_P1_U3372 = ~new_P1_U3370 | ~new_P1_U5177;
  assign new_P1_U3373 = ~new_P1_U2510 | ~new_P1_U4533;
  assign new_P1_U3374 = ~new_P1_U2507 | ~new_P1_U4527;
  assign new_P1_U3375 = ~new_P1_U3373 | ~new_P1_U5234;
  assign new_P1_U3376 = ~new_P1_U3373 | ~new_P1_U5236;
  assign new_P1_U3377 = ~new_P1_U2510 | ~new_P1_U4542;
  assign new_P1_U3378 = ~new_P1_U2507 | ~new_P1_U4600;
  assign new_P1_U3379 = ~new_P1_U3377 | ~new_P1_U5292;
  assign new_P1_U3380 = ~new_P1_U2510 | ~new_P1_U4541;
  assign new_P1_U3381 = ~new_P1_U2507 | ~new_P1_U4658;
  assign new_P1_U3382 = ~new_P1_U3380 | ~new_P1_U5349;
  assign new_P1_U3383 = ~new_P1_U3380 | ~new_P1_U5351;
  assign new_P1_U3384 = ~new_P1_U2510 | ~new_P1_U2488;
  assign new_P1_U3385 = ~new_P1_U2507 | ~new_P1_U2485;
  assign new_P1_U3386 = ~new_P1_U3384 | ~new_P1_U5407;
  assign new_P1_U3387 = ~P1_FLUSH_REG;
  assign new_P1_U3388 = ~new_P1_GTE_485_U6;
  assign new_P1_U3389 = ~new_P1_U3284 | ~new_P1_U3278;
  assign new_P1_U3390 = ~new_P1_U3284 | ~new_P1_U3271;
  assign new_P1_U3391 = ~new_P1_U3512 | ~new_P1_U3513 | ~new_P1_U3515 | ~new_P1_U3514;
  assign new_P1_U3392 = ~new_P1_U7628 | ~new_P1_U5490 | ~new_P1_U5489;
  assign new_P1_U3393 = ~new_P1_U4399 | ~new_P1_U3284;
  assign new_P1_U3394 = ~new_P1_U2605 | ~new_P1_U3277;
  assign new_P1_U3395 = ~new_P1_U4494 | ~new_P1_U4399 | ~new_P1_U7494;
  assign new_P1_U3396 = ~new_P1_U3741 | ~new_P1_U4247;
  assign new_P1_U3397 = ~new_P1_U4399 | ~new_P1_U4494 | ~new_P1_U2605 | ~new_P1_U7494 | ~new_P1_U4477;
  assign new_P1_U3398 = ~new_P1_U4400 | ~new_P1_U4449 | ~new_P1_U4171 | ~new_P1_U2605 | ~new_P1_U4460;
  assign new_P1_U3399 = ~new_P1_U4234 | ~new_P1_U4199 | ~new_P1_U4477;
  assign new_P1_U3400 = ~new_P1_U2449 | ~new_P1_U2447;
  assign new_P1_U3401 = ~new_P1_U3444 | ~new_P1_U5510;
  assign new_P1_U3402 = ~new_P1_U3269 | ~new_P1_U3275;
  assign new_P1_U3403 = ~new_P1_LT_589_U6;
  assign new_P1_U3404 = ~new_P1_U5536 | ~new_P1_U4242 | ~new_P1_U3300;
  assign new_P1_U3405 = ~new_P1_U3284 | ~P1_STATE2_REG_0_ | ~new_P1_U3278;
  assign new_P1_U3406 = ~new_P1_U3271 | ~new_P1_U3273;
  assign new_P1_U3407 = ~new_P1_U3277 | ~new_P1_U3391;
  assign new_P1_U3408 = ~new_P1_U2427 | ~new_P1_U3294;
  assign new_P1_U3409 = ~new_P1_U4460 | ~new_P1_U3391;
  assign new_P1_U3410 = ~new_P1_U4253 | ~new_P1_U3278;
  assign new_P1_U3411 = ~new_P1_U4190 | ~new_P1_U2452;
  assign new_P1_U3412 = ~P1_STATE2_REG_2_ | ~new_P1_U3271;
  assign new_P1_U3413 = ~P1_REIP_REG_0_;
  assign new_P1_U3414 = ~new_P1_U3756 | ~new_P1_U5562;
  assign new_P1_U3415 = ~new_P1_U4400 | ~new_P1_U4173;
  assign new_P1_U3416 = ~new_P1_U3863 | ~new_P1_U4248;
  assign new_P1_U3417 = ~new_P1_U6054 | ~new_P1_U6053;
  assign new_P1_U3418 = ~P1_STATE2_REG_0_ | ~new_P1_U4494;
  assign new_P1_U3419 = ~new_P1_U4399 | ~new_P1_U7494;
  assign new_P1_U3420 = ~new_P1_U4206 | ~new_P1_U4477;
  assign new_P1_U3421 = ~new_P1_U4194 | ~new_P1_U2431;
  assign new_P1_U3422 = ~new_P1_U4210 | ~P1_STATE2_REG_0_;
  assign new_P1_U3423 = ~new_P1_U4503 | ~new_P1_U3391;
  assign new_P1_U3424 = ~new_P1_U4235 | ~new_P1_U6153;
  assign new_P1_U3425 = ~P1_STATE2_REG_0_ | ~new_P1_U4216;
  assign new_P1_U3426 = ~new_P1_U4235 | ~new_P1_U6264;
  assign new_P1_U3427 = ~new_P1_U2452 | ~new_P1_U3886 | ~P1_STATE2_REG_0_ | ~new_P1_U4249;
  assign new_P1_U3428 = ~new_P1_U3866 | ~new_P1_U2447;
  assign new_P1_U3429 = ~P1_EBX_REG_31_;
  assign new_P1_U3430 = ~new_P1_R2337_U69;
  assign new_P1_U3431 = ~new_P1_U4228 | ~new_P1_U3887;
  assign new_P1_U3432 = ~new_P1_U4209 | ~new_P1_U3262;
  assign new_P1_U3433 = ~new_P1_U3952 | ~new_P1_U3955 | ~new_P1_U3962 | ~new_P1_U3958;
  assign new_P1_U3434 = ~new_P1_U4206 | ~new_P1_U3271;
  assign new_P1_U3435 = ~P1_CODEFETCH_REG;
  assign new_P1_U3436 = ~P1_READREQUEST_REG;
  assign new_P1_U3437 = ~new_P1_U2447 | ~new_P1_U4498;
  assign new_P1_U3438 = ~new_P1_U3267 | ~new_P1_U5482;
  assign new_P1_U3439 = ~new_P1_U4449 | ~P1_STATE2_REG_2_;
  assign new_P1_U3440 = ~P1_STATEBS16_REG | ~new_P1_U3263;
  assign new_P1_U3441 = ~new_P1_U3234;
  assign new_P1_U3442 = ~new_P1_U5479 | ~new_P1_U5478;
  assign new_P1_U3443 = ~new_P1_U2450 | ~new_P1_U3441;
  assign new_P1_U3444 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3264;
  assign new_P1_U3445 = ~new_P1_U3274 | ~new_P1_U7064;
  assign new_P1_U3446 = ~new_P1_U4197 | ~new_P1_U4234;
  assign new_P1_U3447 = ~new_P1_U4250 | ~new_P1_U4231 | ~new_P1_U4400;
  assign new_P1_U3448 = ~new_P1_U4250 | ~new_P1_U4231 | ~new_P1_U3278;
  assign new_P1_U3449 = ~new_P1_U4477 | ~new_P1_U4496;
  assign new_P1_U3450 = ~new_P1_U4077 | ~new_P1_U4075 | ~new_P1_U4074 | ~new_P1_U7093;
  assign new_P1_U3451 = ~new_P1_U4254 | ~new_P1_U4266;
  assign new_P1_U3452 = ~new_P1_U4183 | ~new_P1_U3268;
  assign new_P1_U3453 = ~P1_STATE2_REG_0_ | ~new_P1_U2605;
  assign new_P1_U3454 = ~new_P1_U7692 | ~new_P1_U7691;
  assign new_P1_U3455 = ~new_P1_U7695 | ~new_P1_U7694;
  assign new_P1_U3456 = ~new_P1_U7719 | ~new_P1_U7718;
  assign new_P1_U3457 = ~new_P1_U7789 | ~new_P1_U7788;
  assign n5074 = ~new_P1_U7634 | ~new_P1_U7633;
  assign n5079 = ~new_P1_U7636 | ~new_P1_U7635;
  assign n5084 = ~new_P1_U7638 | ~new_P1_U7637;
  assign n5089 = ~new_P1_U7640 | ~new_P1_U7639;
  assign new_P1_U3462 = ~new_P1_U7649 | ~new_P1_U7648;
  assign new_P1_U3463 = new_P1_U3255 & new_P1_U4179;
  assign n5229 = ~new_P1_U7652 | ~new_P1_U7651;
  assign n5234 = ~new_P1_U7654 | ~new_P1_U7653;
  assign n5389 = ~new_P1_U7686 | ~new_P1_U7685;
  assign new_P1_U3467 = new_P1_R2182_U24 & new_P1_U2427 & new_P1_U4215;
  assign n6049 = ~new_P1_U7702 | ~new_P1_U7701;
  assign n6054 = ~new_P1_U7709 | ~new_P1_U7708;
  assign new_P1_U3470 = ~new_P1_U7711 | ~new_P1_U7710;
  assign new_P1_U3471 = ~new_P1_U7714 | ~new_P1_U7713;
  assign n6059 = ~new_P1_U7722 | ~new_P1_U7721;
  assign n6064 = ~new_P1_U7724 | ~new_P1_U7723;
  assign n6069 = ~new_P1_U7728 | ~new_P1_U7727;
  assign n6079 = ~new_P1_U7730 | ~new_P1_U7729;
  assign n6084 = ~new_P1_U7735 | ~new_P1_U7734;
  assign n6089 = ~new_P1_U7737 | ~new_P1_U7736;
  assign n6094 = ~new_P1_U7739 | ~new_P1_U7738;
  assign new_P1_U3479 = new_P1_R2358_U22 & new_P1_U4449;
  assign new_P1_U3480 = ~P1_DATAWIDTH_REG_1_ & ~P1_REIP_REG_1_;
  assign n7219 = ~new_P1_U7755 | ~new_P1_U7754;
  assign n7229 = ~new_P1_U7759 | ~new_P1_U7758;
  assign n7234 = ~new_P1_U7761 | ~new_P1_U7760;
  assign n7244 = ~new_P1_U7763 | ~new_P1_U7762;
  assign n7254 = ~new_P1_U7767 | ~new_P1_U7766;
  assign n7264 = ~new_P1_U7771 | ~new_P1_U7770;
  assign n7278 = ~new_P1_U7773 | ~new_P1_U7772;
  assign new_P1_U3488 = new_P1_R2182_U24 & new_P1_U4215;
  assign new_P1_U3489 = ~new_P1_U7775 | ~new_P1_U7774;
  assign new_P1_U3490 = ~new_P1_U7777 | ~new_P1_U7776;
  assign new_P1_U3491 = ~new_P1_U7779 | ~new_P1_U7778;
  assign new_P1_U3492 = ~new_P1_U7781 | ~new_P1_U7780;
  assign new_P1_U3493 = ~new_P1_U7783 | ~new_P1_U7782;
  assign new_P1_U3494 = new_P1_U4368 & new_P1_U3252;
  assign new_P1_U3495 = new_P1_U4370 & new_P1_U3250;
  assign new_P1_U3496 = P1_REQUESTPENDING_REG & P1_STATE_REG_0_;
  assign new_P1_U3497 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3498 = P1_INSTQUEUERD_ADDR_REG_0_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3499 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3500 = P1_INSTQUEUERD_ADDR_REG_0_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3501 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3502 = P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3503 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3504 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3505 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3506 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3507 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3508 = new_P1_U4383 & new_P1_U4384 & new_P1_U4386 & new_P1_U4385;
  assign new_P1_U3509 = new_P1_U4387 & new_P1_U4388 & new_P1_U4390 & new_P1_U4389;
  assign new_P1_U3510 = new_P1_U4391 & new_P1_U4392 & new_P1_U4394 & new_P1_U4393;
  assign new_P1_U3511 = new_P1_U4395 & new_P1_U4396 & new_P1_U4398 & new_P1_U4397;
  assign new_P1_U3512 = new_P1_U4433 & new_P1_U4434 & new_P1_U4436 & new_P1_U4435;
  assign new_P1_U3513 = new_P1_U4437 & new_P1_U4438 & new_P1_U4440 & new_P1_U4439;
  assign new_P1_U3514 = new_P1_U4441 & new_P1_U4442 & new_P1_U4444 & new_P1_U4443;
  assign new_P1_U3515 = new_P1_U4445 & new_P1_U4446 & new_P1_U4448 & new_P1_U4447;
  assign new_P1_U3516 = new_P1_U4416 & new_P1_U4417 & new_P1_U4419 & new_P1_U4418;
  assign new_P1_U3517 = new_P1_U4420 & new_P1_U4421 & new_P1_U4423 & new_P1_U4422;
  assign new_P1_U3518 = new_P1_U4424 & new_P1_U4425 & new_P1_U4427 & new_P1_U4426;
  assign new_P1_U3519 = new_P1_U4428 & new_P1_U4429 & new_P1_U4431 & new_P1_U4430;
  assign new_P1_U3520 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3521 = P1_INSTQUEUE_REG_5__5_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3522 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3523 = P1_INSTQUEUE_REG_6__5_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3524 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUE_REG_8__5_;
  assign new_P1_U3525 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3526 = P1_INSTQUEUE_REG_10__5_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3527 = P1_INSTQUEUE_REG_12__5_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3528 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3529 = P1_INSTQUEUE_REG_9__5_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3530 = new_P1_U4401 & new_P1_U4402 & new_P1_U4404 & new_P1_U4403;
  assign new_P1_U3531 = new_P1_U4405 & new_P1_U4406 & new_P1_U4408 & new_P1_U4407;
  assign new_P1_U3532 = new_P1_U4409 & new_P1_U4410 & new_P1_U4412 & new_P1_U4411;
  assign new_P1_U3533 = new_P1_U4414 & new_P1_U4413;
  assign new_P1_U3534 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3535 = P1_INSTQUEUE_REG_3__6_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3536 = new_P1_U4450 & new_P1_U4451 & new_P1_U4453 & new_P1_U4452;
  assign new_P1_U3537 = new_P1_U4456 & new_P1_U4455 & new_P1_U4454;
  assign new_P1_U3538 = new_P1_U4459 & new_P1_U4458 & new_P1_U4457;
  assign new_P1_U3539 = new_P1_U7675 & new_P1_U7676 & new_P1_U7678 & new_P1_U7677;
  assign new_P1_U3540 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3541 = P1_INSTQUEUE_REG_1__4_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U3542 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3543 = P1_INSTQUEUE_REG_4__4_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3544 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U3545 = P1_INSTQUEUE_REG_12__4_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3546 = P1_INSTQUEUERD_ADDR_REG_0_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3547 = P1_INSTQUEUE_REG_13__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3548 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3549 = P1_INSTQUEUE_REG_6__4_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3550 = P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3551 = P1_INSTQUEUE_REG_14__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3552 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U3553 = P1_INSTQUEUE_REG_9__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U3554 = new_P1_U7655 & new_P1_U7656 & new_P1_U7658 & new_P1_U7657;
  assign new_P1_U3555 = new_P1_U7659 & new_P1_U7660 & new_P1_U7662 & new_P1_U7661;
  assign new_P1_U3556 = new_P1_U7663 & new_P1_U7664 & new_P1_U7666 & new_P1_U7665;
  assign new_P1_U3557 = new_P1_U7667 & new_P1_U7668 & new_P1_U7670 & new_P1_U7669;
  assign new_P1_U3558 = new_P1_U7494 & new_P1_U3391 & new_P1_U3283;
  assign new_P1_U3559 = new_P1_U4400 & new_P1_U4460 & new_P1_U2605;
  assign new_P1_U3560 = new_P1_U4478 & new_P1_U4479 & new_P1_U4481 & new_P1_U4480;
  assign new_P1_U3561 = new_P1_U4482 & new_P1_U4483 & new_P1_U4485 & new_P1_U4484;
  assign new_P1_U3562 = new_P1_U4486 & new_P1_U4487 & new_P1_U4489 & new_P1_U4488;
  assign new_P1_U3563 = new_P1_U4490 & new_P1_U4491 & new_P1_U4493 & new_P1_U4492;
  assign new_P1_U3564 = new_P1_U4461 & new_P1_U4462 & new_P1_U4464 & new_P1_U4463;
  assign new_P1_U3565 = new_P1_U4465 & new_P1_U4466 & new_P1_U4468 & new_P1_U4467;
  assign new_P1_U3566 = new_P1_U4469 & new_P1_U4470 & new_P1_U4472 & new_P1_U4471;
  assign new_P1_U3567 = new_P1_U4473 & new_P1_U4474 & new_P1_U4476 & new_P1_U4475;
  assign new_P1_U3568 = new_P1_U4377 & new_P1_U4208;
  assign new_P1_U3569 = new_P1_U4416 & new_P1_U4417 & new_P1_U4419 & new_P1_U4418;
  assign new_P1_U3570 = new_P1_U4420 & new_P1_U4421 & new_P1_U4423 & new_P1_U4422;
  assign new_P1_U3571 = new_P1_U4424 & new_P1_U4425 & new_P1_U4427 & new_P1_U4426;
  assign new_P1_U3572 = new_P1_U4428 & new_P1_U4429 & new_P1_U4431 & new_P1_U4430;
  assign new_P1_U3573 = new_P1_U4401 & new_P1_U4402 & new_P1_U4404 & new_P1_U4403;
  assign new_P1_U3574 = new_P1_U4405 & new_P1_U4406 & new_P1_U4408 & new_P1_U4407;
  assign new_P1_U3575 = new_P1_U4409 & new_P1_U4410 & new_P1_U4412 & new_P1_U4411;
  assign new_P1_U3576 = new_P1_U4414 & new_P1_U4413;
  assign new_P1_U3577 = new_P1_U4399 & new_P1_U4171;
  assign new_P1_U3578 = new_P1_U4249 & new_P1_U3283;
  assign new_P1_U3579 = new_P1_U7494 & new_P1_U4400 & new_P1_U3284 & new_P1_U3283;
  assign new_P1_U3580 = new_P1_U4217 & new_P1_U3400;
  assign new_P1_U3581 = P1_STATE2_REG_2_ & new_P1_U7603;
  assign new_P1_U3582 = new_P1_U4515 & new_P1_U3297;
  assign new_P1_U3583 = new_P1_U2427 & new_P1_U3257;
  assign new_P1_U3584 = P1_STATE2_REG_3_ & P1_STATE2_REG_0_;
  assign new_P1_U3585 = new_P1_U4246 & new_P1_U4241;
  assign new_P1_U3586 = new_P1_U3585 & new_P1_U4523;
  assign new_P1_U3587 = new_P1_U4224 & new_P1_U4552 & new_P1_U4553;
  assign new_P1_U3588 = new_P1_U4562 & new_P1_U4561 & new_P1_U4560;
  assign new_P1_U3589 = new_P1_U4567 & new_P1_U4566 & new_P1_U4565;
  assign new_P1_U3590 = new_P1_U4572 & new_P1_U4571 & new_P1_U4570;
  assign new_P1_U3591 = new_P1_U4577 & new_P1_U4576 & new_P1_U4575;
  assign new_P1_U3592 = new_P1_U4582 & new_P1_U4581 & new_P1_U4580;
  assign new_P1_U3593 = new_P1_U4587 & new_P1_U4586 & new_P1_U4585;
  assign new_P1_U3594 = new_P1_U4592 & new_P1_U4591 & new_P1_U4590;
  assign new_P1_U3595 = new_P1_U4597 & new_P1_U4596 & new_P1_U4595;
  assign new_P1_U3596 = new_P1_U4224 & new_P1_U4610 & new_P1_U4611;
  assign new_P1_U3597 = new_P1_U4620 & new_P1_U4619 & new_P1_U4618;
  assign new_P1_U3598 = new_P1_U4625 & new_P1_U4624 & new_P1_U4623;
  assign new_P1_U3599 = new_P1_U4630 & new_P1_U4629 & new_P1_U4628;
  assign new_P1_U3600 = new_P1_U4635 & new_P1_U4634 & new_P1_U4633;
  assign new_P1_U3601 = new_P1_U4640 & new_P1_U4639 & new_P1_U4638;
  assign new_P1_U3602 = new_P1_U4645 & new_P1_U4644 & new_P1_U4643;
  assign new_P1_U3603 = new_P1_U4650 & new_P1_U4649 & new_P1_U4648;
  assign new_P1_U3604 = new_P1_U4655 & new_P1_U4654 & new_P1_U4653;
  assign new_P1_U3605 = new_P1_U4224 & new_P1_U4669 & new_P1_U4670;
  assign new_P1_U3606 = new_P1_U4679 & new_P1_U4678 & new_P1_U4677;
  assign new_P1_U3607 = new_P1_U4684 & new_P1_U4683 & new_P1_U4682;
  assign new_P1_U3608 = new_P1_U4689 & new_P1_U4688 & new_P1_U4687;
  assign new_P1_U3609 = new_P1_U4694 & new_P1_U4693 & new_P1_U4692;
  assign new_P1_U3610 = new_P1_U4699 & new_P1_U4698 & new_P1_U4697;
  assign new_P1_U3611 = new_P1_U4704 & new_P1_U4703 & new_P1_U4702;
  assign new_P1_U3612 = new_P1_U4709 & new_P1_U4708 & new_P1_U4707;
  assign new_P1_U3613 = new_P1_U4714 & new_P1_U4713 & new_P1_U4712;
  assign new_P1_U3614 = new_P1_U4224 & new_P1_U4726 & new_P1_U4727;
  assign new_P1_U3615 = new_P1_U4736 & new_P1_U4735 & new_P1_U4734;
  assign new_P1_U3616 = new_P1_U4741 & new_P1_U4740 & new_P1_U4739;
  assign new_P1_U3617 = new_P1_U4746 & new_P1_U4745 & new_P1_U4744;
  assign new_P1_U3618 = new_P1_U4751 & new_P1_U4750 & new_P1_U4749;
  assign new_P1_U3619 = new_P1_U4756 & new_P1_U4755 & new_P1_U4754;
  assign new_P1_U3620 = new_P1_U4761 & new_P1_U4760 & new_P1_U4759;
  assign new_P1_U3621 = new_P1_U4766 & new_P1_U4765 & new_P1_U4764;
  assign new_P1_U3622 = new_P1_U4771 & new_P1_U4770 & new_P1_U4769;
  assign new_P1_U3623 = new_P1_U4224 & new_P1_U4784 & new_P1_U4785;
  assign new_P1_U3624 = new_P1_U4794 & new_P1_U4793 & new_P1_U4792;
  assign new_P1_U3625 = new_P1_U4799 & new_P1_U4798 & new_P1_U4797;
  assign new_P1_U3626 = new_P1_U4804 & new_P1_U4803 & new_P1_U4802;
  assign new_P1_U3627 = new_P1_U4809 & new_P1_U4808 & new_P1_U4807;
  assign new_P1_U3628 = new_P1_U4814 & new_P1_U4813 & new_P1_U4812;
  assign new_P1_U3629 = new_P1_U4819 & new_P1_U4818 & new_P1_U4817;
  assign new_P1_U3630 = new_P1_U4824 & new_P1_U4823 & new_P1_U4822;
  assign new_P1_U3631 = new_P1_U4829 & new_P1_U4828 & new_P1_U4827;
  assign new_P1_U3632 = new_P1_U4224 & new_P1_U4841 & new_P1_U4842;
  assign new_P1_U3633 = new_P1_U4851 & new_P1_U4850 & new_P1_U4849;
  assign new_P1_U3634 = new_P1_U4856 & new_P1_U4855 & new_P1_U4854;
  assign new_P1_U3635 = new_P1_U4861 & new_P1_U4860 & new_P1_U4859;
  assign new_P1_U3636 = new_P1_U4866 & new_P1_U4865 & new_P1_U4864;
  assign new_P1_U3637 = new_P1_U4871 & new_P1_U4870 & new_P1_U4869;
  assign new_P1_U3638 = new_P1_U4876 & new_P1_U4875 & new_P1_U4874;
  assign new_P1_U3639 = new_P1_U4881 & new_P1_U4880 & new_P1_U4879;
  assign new_P1_U3640 = new_P1_U4886 & new_P1_U4885 & new_P1_U4884;
  assign new_P1_U3641 = new_P1_U4224 & new_P1_U4899 & new_P1_U4900;
  assign new_P1_U3642 = new_P1_U4909 & new_P1_U4908 & new_P1_U4907;
  assign new_P1_U3643 = new_P1_U4914 & new_P1_U4913 & new_P1_U4912;
  assign new_P1_U3644 = new_P1_U4919 & new_P1_U4918 & new_P1_U4917;
  assign new_P1_U3645 = new_P1_U4924 & new_P1_U4923 & new_P1_U4922;
  assign new_P1_U3646 = new_P1_U4929 & new_P1_U4928 & new_P1_U4927;
  assign new_P1_U3647 = new_P1_U4934 & new_P1_U4933 & new_P1_U4932;
  assign new_P1_U3648 = new_P1_U4939 & new_P1_U4938 & new_P1_U4937;
  assign new_P1_U3649 = new_P1_U4944 & new_P1_U4943 & new_P1_U4942;
  assign new_P1_U3650 = new_P1_U4224 & new_P1_U4956 & new_P1_U4957;
  assign new_P1_U3651 = new_P1_U4966 & new_P1_U4965 & new_P1_U4964;
  assign new_P1_U3652 = new_P1_U4971 & new_P1_U4970 & new_P1_U4969;
  assign new_P1_U3653 = new_P1_U4976 & new_P1_U4975 & new_P1_U4974;
  assign new_P1_U3654 = new_P1_U4981 & new_P1_U4980 & new_P1_U4979;
  assign new_P1_U3655 = new_P1_U4986 & new_P1_U4985 & new_P1_U4984;
  assign new_P1_U3656 = new_P1_U4991 & new_P1_U4990 & new_P1_U4989;
  assign new_P1_U3657 = new_P1_U4996 & new_P1_U4995 & new_P1_U4994;
  assign new_P1_U3658 = new_P1_U5001 & new_P1_U5000 & new_P1_U4999;
  assign new_P1_U3659 = new_P1_U4224 & new_P1_U5012 & new_P1_U5013;
  assign new_P1_U3660 = new_P1_U5022 & new_P1_U5021 & new_P1_U5020;
  assign new_P1_U3661 = new_P1_U5027 & new_P1_U5026 & new_P1_U5025;
  assign new_P1_U3662 = new_P1_U5032 & new_P1_U5031 & new_P1_U5030;
  assign new_P1_U3663 = new_P1_U5037 & new_P1_U5036 & new_P1_U5035;
  assign new_P1_U3664 = new_P1_U5042 & new_P1_U5041 & new_P1_U5040;
  assign new_P1_U3665 = new_P1_U5047 & new_P1_U5046 & new_P1_U5045;
  assign new_P1_U3666 = new_P1_U5052 & new_P1_U5051 & new_P1_U5050;
  assign new_P1_U3667 = new_P1_U5057 & new_P1_U5056 & new_P1_U5055;
  assign new_P1_U3668 = new_P1_U4224 & new_P1_U5069 & new_P1_U5070;
  assign new_P1_U3669 = new_P1_U5079 & new_P1_U5078 & new_P1_U5077;
  assign new_P1_U3670 = new_P1_U5084 & new_P1_U5083 & new_P1_U5082;
  assign new_P1_U3671 = new_P1_U5089 & new_P1_U5088 & new_P1_U5087;
  assign new_P1_U3672 = new_P1_U5094 & new_P1_U5093 & new_P1_U5092;
  assign new_P1_U3673 = new_P1_U5099 & new_P1_U5098 & new_P1_U5097;
  assign new_P1_U3674 = new_P1_U5104 & new_P1_U5103 & new_P1_U5102;
  assign new_P1_U3675 = new_P1_U5109 & new_P1_U5108 & new_P1_U5107;
  assign new_P1_U3676 = new_P1_U5114 & new_P1_U5113 & new_P1_U5112;
  assign new_P1_U3677 = new_P1_U4224 & new_P1_U5127 & new_P1_U5128;
  assign new_P1_U3678 = new_P1_U5137 & new_P1_U5136 & new_P1_U5135;
  assign new_P1_U3679 = new_P1_U5142 & new_P1_U5141 & new_P1_U5140;
  assign new_P1_U3680 = new_P1_U5147 & new_P1_U5146 & new_P1_U5145;
  assign new_P1_U3681 = new_P1_U5152 & new_P1_U5151 & new_P1_U5150;
  assign new_P1_U3682 = new_P1_U5157 & new_P1_U5156 & new_P1_U5155;
  assign new_P1_U3683 = new_P1_U5162 & new_P1_U5161 & new_P1_U5160;
  assign new_P1_U3684 = new_P1_U5167 & new_P1_U5166 & new_P1_U5165;
  assign new_P1_U3685 = new_P1_U5172 & new_P1_U5171 & new_P1_U5170;
  assign new_P1_U3686 = new_P1_U4224 & new_P1_U5184 & new_P1_U5185;
  assign new_P1_U3687 = new_P1_U5194 & new_P1_U5193 & new_P1_U5192;
  assign new_P1_U3688 = new_P1_U5199 & new_P1_U5198 & new_P1_U5197;
  assign new_P1_U3689 = new_P1_U5204 & new_P1_U5203 & new_P1_U5202;
  assign new_P1_U3690 = new_P1_U5209 & new_P1_U5208 & new_P1_U5207;
  assign new_P1_U3691 = new_P1_U5214 & new_P1_U5213 & new_P1_U5212;
  assign new_P1_U3692 = new_P1_U5219 & new_P1_U5218 & new_P1_U5217;
  assign new_P1_U3693 = new_P1_U5224 & new_P1_U5223 & new_P1_U5222;
  assign new_P1_U3694 = new_P1_U5229 & new_P1_U5228 & new_P1_U5227;
  assign new_P1_U3695 = new_P1_U4224 & new_P1_U5242 & new_P1_U5243;
  assign new_P1_U3696 = new_P1_U5252 & new_P1_U5251 & new_P1_U5250;
  assign new_P1_U3697 = new_P1_U5257 & new_P1_U5256 & new_P1_U5255;
  assign new_P1_U3698 = new_P1_U5262 & new_P1_U5261 & new_P1_U5260;
  assign new_P1_U3699 = new_P1_U5267 & new_P1_U5266 & new_P1_U5265;
  assign new_P1_U3700 = new_P1_U5272 & new_P1_U5271 & new_P1_U5270;
  assign new_P1_U3701 = new_P1_U5277 & new_P1_U5276 & new_P1_U5275;
  assign new_P1_U3702 = new_P1_U5282 & new_P1_U5281 & new_P1_U5280;
  assign new_P1_U3703 = new_P1_U5287 & new_P1_U5286 & new_P1_U5285;
  assign new_P1_U3704 = new_P1_U4224 & new_P1_U5299 & new_P1_U5300;
  assign new_P1_U3705 = new_P1_U5309 & new_P1_U5308 & new_P1_U5307;
  assign new_P1_U3706 = new_P1_U5314 & new_P1_U5313 & new_P1_U5312;
  assign new_P1_U3707 = new_P1_U5319 & new_P1_U5318 & new_P1_U5317;
  assign new_P1_U3708 = new_P1_U5324 & new_P1_U5323 & new_P1_U5322;
  assign new_P1_U3709 = new_P1_U5329 & new_P1_U5328 & new_P1_U5327;
  assign new_P1_U3710 = new_P1_U5334 & new_P1_U5333 & new_P1_U5332;
  assign new_P1_U3711 = new_P1_U5339 & new_P1_U5338 & new_P1_U5337;
  assign new_P1_U3712 = new_P1_U5344 & new_P1_U5343 & new_P1_U5342;
  assign new_P1_U3713 = new_P1_U4224 & new_P1_U5357 & new_P1_U5358;
  assign new_P1_U3714 = new_P1_U5367 & new_P1_U5366 & new_P1_U5365;
  assign new_P1_U3715 = new_P1_U5372 & new_P1_U5371 & new_P1_U5370;
  assign new_P1_U3716 = new_P1_U5377 & new_P1_U5376 & new_P1_U5375;
  assign new_P1_U3717 = new_P1_U5382 & new_P1_U5381 & new_P1_U5380;
  assign new_P1_U3718 = new_P1_U5387 & new_P1_U5386 & new_P1_U5385;
  assign new_P1_U3719 = new_P1_U5392 & new_P1_U5391 & new_P1_U5390;
  assign new_P1_U3720 = new_P1_U5397 & new_P1_U5396 & new_P1_U5395;
  assign new_P1_U3721 = new_P1_U5402 & new_P1_U5401 & new_P1_U5400;
  assign new_P1_U3722 = new_P1_U4224 & new_P1_U5414 & new_P1_U5415;
  assign new_P1_U3723 = new_P1_U5424 & new_P1_U5423 & new_P1_U5422;
  assign new_P1_U3724 = new_P1_U5429 & new_P1_U5428 & new_P1_U5427;
  assign new_P1_U3725 = new_P1_U5434 & new_P1_U5433 & new_P1_U5432;
  assign new_P1_U3726 = new_P1_U5439 & new_P1_U5438 & new_P1_U5437;
  assign new_P1_U3727 = new_P1_U5443 & new_P1_U5442 & new_P1_U5441;
  assign new_P1_U3728 = new_P1_U5448 & new_P1_U5447 & new_P1_U5446;
  assign new_P1_U3729 = new_P1_U5453 & new_P1_U5452 & new_P1_U5451;
  assign new_P1_U3730 = new_P1_U5458 & new_P1_U5457 & new_P1_U5456;
  assign new_P1_U3731 = P1_FLUSH_REG & P1_STATE2_REG_0_;
  assign new_P1_U3732 = new_P1_U4494 & new_P1_U4399;
  assign new_P1_U3733 = new_P1_U4497 & new_P1_U3257;
  assign new_P1_U3734 = new_P1_U4210 & new_P1_U3257;
  assign new_P1_U3735 = new_P1_U7496 & new_P1_U4217;
  assign new_P1_U3736 = new_P1_U5471 & new_P1_U5472;
  assign new_P1_U3737 = new_P1_U3736 & new_P1_U5470;
  assign new_P1_U3738 = new_P1_U3737 & new_P1_U2518;
  assign new_P1_U3739 = new_P1_U5475 & new_P1_U4242;
  assign new_P1_U3740 = new_P1_U5486 & new_P1_U5485;
  assign new_P1_U3741 = new_P1_U4449 & new_P1_U4400;
  assign new_P1_U3742 = new_P1_U5496 & new_P1_U3393;
  assign new_P1_U3743 = new_P1_U5498 & new_P1_U5497;
  assign new_P1_U3744 = new_P1_U3743 & new_P1_U3742 & new_P1_U5500 & new_P1_U7627;
  assign new_P1_U3745 = new_P1_U4263 & new_P1_U3397;
  assign new_P1_U3746 = new_P1_U3279 & new_P1_U2520 & new_P1_U3745 & new_P1_U3411 & new_P1_U3288;
  assign new_P1_U3747 = new_P1_U3748 & new_P1_U5502;
  assign new_P1_U3748 = new_P1_U5505 & new_P1_U5504;
  assign new_P1_U3749 = new_P1_U5513 & new_P1_U7717 & new_P1_U7716;
  assign new_P1_U3750 = new_P1_U5524 & new_P1_U5522;
  assign new_P1_U3751 = new_P1_U5543 & new_P1_U5544;
  assign new_P1_U3752 = new_P1_U5547 & new_P1_U5548;
  assign new_P1_U3753 = new_P1_U5552 & new_P1_U5553;
  assign new_P1_U3754 = new_P1_U5558 & new_P1_U3257;
  assign new_P1_U3755 = new_P1_U3284 & new_P1_U3407;
  assign new_P1_U3756 = new_P1_U5563 & new_P1_U5561;
  assign new_P1_U3757 = new_P1_U5567 & new_P1_U3398 & new_P1_U3399;
  assign new_P1_U3758 = new_P1_U3757 & new_P1_U2520 & new_P1_U5568;
  assign new_P1_U3759 = new_P1_U4186 & new_P1_U3284;
  assign new_P1_U3760 = new_P1_U3448 & new_P1_U3288 & new_P1_U4217;
  assign new_P1_U3761 = new_P1_U5566 & new_P1_U7507;
  assign new_P1_U3762 = new_P1_U7508 & P1_STATE2_REG_2_;
  assign new_P1_U3763 = new_P1_U5571 & new_P1_U5570;
  assign new_P1_U3764 = new_P1_U5573 & new_P1_U5572;
  assign new_P1_U3765 = new_P1_U5575 & new_P1_U5576;
  assign new_P1_U3766 = new_P1_U3765 & new_P1_U5574;
  assign new_P1_U3767 = new_P1_U5578 & new_P1_U5577;
  assign new_P1_U3768 = new_P1_U5580 & new_P1_U5579;
  assign new_P1_U3769 = new_P1_U5582 & new_P1_U5583;
  assign new_P1_U3770 = new_P1_U3769 & new_P1_U5581;
  assign new_P1_U3771 = new_P1_U5585 & new_P1_U5584;
  assign new_P1_U3772 = new_P1_U5587 & new_P1_U5586;
  assign new_P1_U3773 = new_P1_U5589 & new_P1_U5590;
  assign new_P1_U3774 = new_P1_U3773 & new_P1_U5588;
  assign new_P1_U3775 = new_P1_U5594 & new_P1_U5592 & new_P1_U5591;
  assign new_P1_U3776 = new_P1_U5593 & new_P1_U3777 & new_P1_U5595;
  assign new_P1_U3777 = new_P1_U5596 & new_P1_U5597;
  assign new_P1_U3778 = new_P1_U5601 & new_P1_U5599 & new_P1_U5598;
  assign new_P1_U3779 = new_P1_U5603 & new_P1_U5604;
  assign new_P1_U3780 = new_P1_U3779 & new_P1_U5602;
  assign new_P1_U3781 = new_P1_U5608 & new_P1_U5606 & new_P1_U5605;
  assign new_P1_U3782 = new_P1_U5610 & new_P1_U5611;
  assign new_P1_U3783 = new_P1_U3782 & new_P1_U5609;
  assign new_P1_U3784 = new_P1_U5615 & new_P1_U5613 & new_P1_U5612;
  assign new_P1_U3785 = new_P1_U5617 & new_P1_U5618;
  assign new_P1_U3786 = new_P1_U3785 & new_P1_U5616;
  assign new_P1_U3787 = new_P1_U5622 & new_P1_U5620 & new_P1_U5619;
  assign new_P1_U3788 = new_P1_U5624 & new_P1_U5625;
  assign new_P1_U3789 = new_P1_U3788 & new_P1_U5623;
  assign new_P1_U3790 = new_P1_U5629 & new_P1_U5627 & new_P1_U5626;
  assign new_P1_U3791 = new_P1_U5631 & new_P1_U5632;
  assign new_P1_U3792 = new_P1_U3791 & new_P1_U5630;
  assign new_P1_U3793 = new_P1_U5636 & new_P1_U5634 & new_P1_U5633;
  assign new_P1_U3794 = new_P1_U5638 & new_P1_U5639;
  assign new_P1_U3795 = new_P1_U3794 & new_P1_U5637;
  assign new_P1_U3796 = new_P1_U5643 & new_P1_U5641 & new_P1_U5640;
  assign new_P1_U3797 = new_P1_U5645 & new_P1_U5646;
  assign new_P1_U3798 = new_P1_U3797 & new_P1_U5644;
  assign new_P1_U3799 = new_P1_U5650 & new_P1_U5648 & new_P1_U5647;
  assign new_P1_U3800 = new_P1_U5652 & new_P1_U5653;
  assign new_P1_U3801 = new_P1_U3800 & new_P1_U5651;
  assign new_P1_U3802 = new_P1_U5657 & new_P1_U5655 & new_P1_U5654;
  assign new_P1_U3803 = new_P1_U5659 & new_P1_U5660;
  assign new_P1_U3804 = new_P1_U3803 & new_P1_U5658;
  assign new_P1_U3805 = new_P1_U5662 & new_P1_U5664;
  assign new_P1_U3806 = new_P1_U5666 & new_P1_U5667;
  assign new_P1_U3807 = new_P1_U3806 & new_P1_U5665;
  assign new_P1_U3808 = new_P1_U5669 & new_P1_U5671;
  assign new_P1_U3809 = new_P1_U5673 & new_P1_U5674;
  assign new_P1_U3810 = new_P1_U3809 & new_P1_U5672;
  assign new_P1_U3811 = new_P1_U5676 & new_P1_U5678;
  assign new_P1_U3812 = new_P1_U5680 & new_P1_U5681;
  assign new_P1_U3813 = new_P1_U3812 & new_P1_U5679;
  assign new_P1_U3814 = new_P1_U5683 & new_P1_U5685;
  assign new_P1_U3815 = new_P1_U5687 & new_P1_U5688;
  assign new_P1_U3816 = new_P1_U3815 & new_P1_U5686;
  assign new_P1_U3817 = new_P1_U5690 & new_P1_U5692;
  assign new_P1_U3818 = new_P1_U5694 & new_P1_U5695;
  assign new_P1_U3819 = new_P1_U3818 & new_P1_U5693;
  assign new_P1_U3820 = new_P1_U5697 & new_P1_U5699;
  assign new_P1_U3821 = new_P1_U5701 & new_P1_U5702;
  assign new_P1_U3822 = new_P1_U3821 & new_P1_U5700;
  assign new_P1_U3823 = new_P1_U5704 & new_P1_U5706;
  assign new_P1_U3824 = new_P1_U5708 & new_P1_U5709;
  assign new_P1_U3825 = new_P1_U3824 & new_P1_U5707;
  assign new_P1_U3826 = new_P1_U5711 & new_P1_U5713;
  assign new_P1_U3827 = new_P1_U5715 & new_P1_U5716;
  assign new_P1_U3828 = new_P1_U3827 & new_P1_U5714;
  assign new_P1_U3829 = new_P1_U5718 & new_P1_U5720;
  assign new_P1_U3830 = new_P1_U5722 & new_P1_U5723;
  assign new_P1_U3831 = new_P1_U3830 & new_P1_U5721;
  assign new_P1_U3832 = new_P1_U5725 & new_P1_U5727;
  assign new_P1_U3833 = new_P1_U5729 & new_P1_U5730;
  assign new_P1_U3834 = new_P1_U3833 & new_P1_U5728;
  assign new_P1_U3835 = new_P1_U5732 & new_P1_U5734;
  assign new_P1_U3836 = new_P1_U5736 & new_P1_U5737;
  assign new_P1_U3837 = new_P1_U3836 & new_P1_U5735;
  assign new_P1_U3838 = new_P1_U5739 & new_P1_U5741;
  assign new_P1_U3839 = new_P1_U5743 & new_P1_U5744;
  assign new_P1_U3840 = new_P1_U3839 & new_P1_U5742;
  assign new_P1_U3841 = new_P1_U5746 & new_P1_U5748;
  assign new_P1_U3842 = new_P1_U5750 & new_P1_U5751;
  assign new_P1_U3843 = new_P1_U3842 & new_P1_U5749;
  assign new_P1_U3844 = new_P1_U5753 & new_P1_U5755;
  assign new_P1_U3845 = new_P1_U5757 & new_P1_U5758;
  assign new_P1_U3846 = new_P1_U3845 & new_P1_U5756;
  assign new_P1_U3847 = new_P1_U5760 & new_P1_U5762;
  assign new_P1_U3848 = new_P1_U5764 & new_P1_U5765;
  assign new_P1_U3849 = new_P1_U3848 & new_P1_U5763;
  assign new_P1_U3850 = new_P1_U5767 & new_P1_U5769;
  assign new_P1_U3851 = new_P1_U5771 & new_P1_U5772;
  assign new_P1_U3852 = new_P1_U3851 & new_P1_U5770;
  assign new_P1_U3853 = new_P1_U5774 & new_P1_U5776;
  assign new_P1_U3854 = new_P1_U5778 & new_P1_U5779;
  assign new_P1_U3855 = new_P1_U3854 & new_P1_U5777;
  assign new_P1_U3856 = new_P1_U5781 & new_P1_U5783;
  assign new_P1_U3857 = new_P1_U5785 & new_P1_U5786;
  assign new_P1_U3858 = new_P1_U3857 & new_P1_U5784;
  assign new_P1_U3859 = new_P1_U5788 & new_P1_U5790;
  assign new_P1_U3860 = new_P1_U5792 & new_P1_U5793;
  assign new_P1_U3861 = new_P1_U3860 & new_P1_U5791;
  assign new_P1_U3862 = new_P1_U7494 & new_P1_U3283 & new_P1_U3262;
  assign new_P1_U3863 = new_P1_U5794 & new_P1_U3408;
  assign new_P1_U3864 = P1_STATE2_REG_1_ & P1_STATEBS16_REG;
  assign new_P1_U3865 = new_P1_U2368 & new_P1_U3284;
  assign new_P1_U3866 = new_P1_U2449 & P1_STATE2_REG_0_;
  assign new_P1_U3867 = new_P1_U4208 & new_P1_U2368;
  assign new_P1_U3868 = new_P1_U6105 & new_P1_U6106;
  assign new_P1_U3869 = new_P1_U6108 & new_P1_U6109;
  assign new_P1_U3870 = new_P1_U6111 & new_P1_U6112;
  assign new_P1_U3871 = new_P1_U6114 & new_P1_U6115;
  assign new_P1_U3872 = new_P1_U6117 & new_P1_U6118;
  assign new_P1_U3873 = new_P1_U6120 & new_P1_U6121;
  assign new_P1_U3874 = new_P1_U6123 & new_P1_U6124;
  assign new_P1_U3875 = new_P1_U6126 & new_P1_U6127;
  assign new_P1_U3876 = new_P1_U6129 & new_P1_U6130;
  assign new_P1_U3877 = new_P1_U6132 & new_P1_U6133;
  assign new_P1_U3878 = new_P1_U6135 & new_P1_U6136;
  assign new_P1_U3879 = new_P1_U6138 & new_P1_U6139;
  assign new_P1_U3880 = new_P1_U6141 & new_P1_U6142;
  assign new_P1_U3881 = new_P1_U6144 & new_P1_U6145;
  assign new_P1_U3882 = new_P1_U6147 & new_P1_U6148;
  assign new_P1_U3883 = new_P1_U6151 & new_P1_U6150;
  assign new_P1_U3884 = new_P1_U2605 & new_P1_U3391;
  assign new_P1_U3885 = new_P1_U7494 & P1_STATE2_REG_0_ & new_P1_U3271;
  assign new_P1_U3886 = new_P1_U4399 & new_P1_U4171;
  assign new_P1_U3887 = new_P1_U6362 & new_P1_U4241 & new_P1_U4244;
  assign new_P1_U3888 = ~new_U210 & ~P1_STATEBS16_REG;
  assign new_P1_U3889 = new_P1_U4494 & new_P1_U4186;
  assign new_P1_U3890 = new_P1_U6371 & new_P1_U6374 & new_P1_U6375 & new_P1_U6373 & new_P1_U6372;
  assign new_P1_U3891 = new_P1_U6379 & new_P1_U6382 & new_P1_U6383 & new_P1_U6381 & new_P1_U6380;
  assign new_P1_U3892 = new_P1_U6387 & new_P1_U6390 & new_P1_U6391 & new_P1_U6389 & new_P1_U6388;
  assign new_P1_U3893 = new_P1_U6395 & new_P1_U6398 & new_P1_U6399 & new_P1_U6397 & new_P1_U6396;
  assign new_P1_U3894 = new_P1_U6400 & new_P1_U4227;
  assign new_P1_U3895 = new_P1_U6406 & new_P1_U6407 & new_P1_U6405 & new_P1_U6404;
  assign new_P1_U3896 = new_P1_U6408 & new_P1_U4227;
  assign new_P1_U3897 = new_P1_U6411 & new_P1_U6414 & new_P1_U6415 & new_P1_U6413 & new_P1_U6412;
  assign new_P1_U3898 = new_P1_U6416 & new_P1_U4227;
  assign new_P1_U3899 = new_P1_U6421 & new_P1_U6422 & new_P1_U6419;
  assign new_P1_U3900 = new_P1_U6423 & new_P1_U4227;
  assign new_P1_U3901 = new_P1_U6428 & new_P1_U6429 & new_P1_U6426;
  assign new_P1_U3902 = new_P1_U6430 & new_P1_U4227;
  assign new_P1_U3903 = new_P1_U6435 & new_P1_U6436 & new_P1_U6433;
  assign new_P1_U3904 = new_P1_U6437 & new_P1_U4227;
  assign new_P1_U3905 = new_P1_U6442 & new_P1_U6443 & new_P1_U6440;
  assign new_P1_U3906 = new_P1_U6444 & new_P1_U4227;
  assign new_P1_U3907 = new_P1_U6449 & new_P1_U6450 & new_P1_U6447;
  assign new_P1_U3908 = new_P1_U6451 & new_P1_U4227;
  assign new_P1_U3909 = new_P1_U6456 & new_P1_U6457 & new_P1_U6454;
  assign new_P1_U3910 = new_P1_U6458 & new_P1_U4227;
  assign new_P1_U3911 = new_P1_U6463 & new_P1_U6464 & new_P1_U6461;
  assign new_P1_U3912 = new_P1_U6465 & new_P1_U4227;
  assign new_P1_U3913 = new_P1_U6470 & new_P1_U6471 & new_P1_U6468;
  assign new_P1_U3914 = new_P1_U6472 & new_P1_U4227;
  assign new_P1_U3915 = new_P1_U6477 & new_P1_U6478 & new_P1_U6475;
  assign new_P1_U3916 = new_P1_U6479 & new_P1_U4227;
  assign new_P1_U3917 = new_P1_U6484 & new_P1_U6485 & new_P1_U6482;
  assign new_P1_U3918 = new_P1_U6486 & new_P1_U4227;
  assign new_P1_U3919 = new_P1_U6491 & new_P1_U6492 & new_P1_U6489;
  assign new_P1_U3920 = new_P1_U4227 & new_P1_U6494;
  assign new_P1_U3921 = new_P1_U6498 & new_P1_U6499 & new_P1_U6496;
  assign new_P1_U3922 = new_P1_U4227 & new_P1_U6501;
  assign new_P1_U3923 = new_P1_U6505 & new_P1_U6506 & new_P1_U6503;
  assign new_P1_U3924 = new_P1_U4227 & new_P1_U6508;
  assign new_P1_U3925 = new_P1_U6512 & new_P1_U6513 & new_P1_U6510;
  assign new_P1_U3926 = new_P1_U6517 & new_P1_U6515;
  assign new_P1_U3927 = new_P1_U6519 & new_P1_U6520;
  assign new_P1_U3928 = new_P1_U6524 & new_P1_U6522;
  assign new_P1_U3929 = new_P1_U6526 & new_P1_U6527;
  assign new_P1_U3930 = new_P1_U6531 & new_P1_U6529;
  assign new_P1_U3931 = new_P1_U6533 & new_P1_U6534;
  assign new_P1_U3932 = new_P1_U6538 & new_P1_U6536;
  assign new_P1_U3933 = new_P1_U6540 & new_P1_U6541;
  assign new_P1_U3934 = new_P1_U6545 & new_P1_U6543;
  assign new_P1_U3935 = new_P1_U6547 & new_P1_U6548;
  assign new_P1_U3936 = new_P1_U6552 & new_P1_U6550;
  assign new_P1_U3937 = new_P1_U6554 & new_P1_U6555;
  assign new_P1_U3938 = new_P1_U6559 & new_P1_U6557;
  assign new_P1_U3939 = new_P1_U6561 & new_P1_U6562;
  assign new_P1_U3940 = new_P1_U6566 & new_P1_U6564;
  assign new_P1_U3941 = new_P1_U6568 & new_P1_U6569;
  assign new_P1_U3942 = new_P1_U6573 & new_P1_U6571;
  assign new_P1_U3943 = new_P1_U6575 & new_P1_U6576;
  assign new_P1_U3944 = new_P1_U6580 & new_P1_U6578;
  assign new_P1_U3945 = new_P1_U6582 & new_P1_U6583;
  assign new_P1_U3946 = new_P1_U6587 & new_P1_U6585;
  assign new_P1_U3947 = new_P1_U6589 & new_P1_U6590;
  assign new_P1_U3948 = new_P1_U6594 & new_P1_U6592;
  assign new_P1_U3949 = new_P1_U6596 & new_P1_U6597;
  assign new_P1_U3950 = ~P1_DATAWIDTH_REG_5_ & ~P1_DATAWIDTH_REG_4_ & ~P1_DATAWIDTH_REG_2_ & ~P1_DATAWIDTH_REG_3_;
  assign new_P1_U3951 = ~P1_DATAWIDTH_REG_9_ & ~P1_DATAWIDTH_REG_8_ & ~P1_DATAWIDTH_REG_6_ & ~P1_DATAWIDTH_REG_7_;
  assign new_P1_U3952 = new_P1_U3951 & new_P1_U3950;
  assign new_P1_U3953 = ~P1_DATAWIDTH_REG_13_ & ~P1_DATAWIDTH_REG_12_ & ~P1_DATAWIDTH_REG_10_ & ~P1_DATAWIDTH_REG_11_;
  assign new_P1_U3954 = ~P1_DATAWIDTH_REG_17_ & ~P1_DATAWIDTH_REG_16_ & ~P1_DATAWIDTH_REG_14_ & ~P1_DATAWIDTH_REG_15_;
  assign new_P1_U3955 = new_P1_U3954 & new_P1_U3953;
  assign new_P1_U3956 = ~P1_DATAWIDTH_REG_21_ & ~P1_DATAWIDTH_REG_20_ & ~P1_DATAWIDTH_REG_18_ & ~P1_DATAWIDTH_REG_19_;
  assign new_P1_U3957 = ~P1_DATAWIDTH_REG_25_ & ~P1_DATAWIDTH_REG_24_ & ~P1_DATAWIDTH_REG_22_ & ~P1_DATAWIDTH_REG_23_;
  assign new_P1_U3958 = new_P1_U3957 & new_P1_U3956;
  assign new_P1_U3959 = ~P1_DATAWIDTH_REG_26_ & ~P1_DATAWIDTH_REG_27_;
  assign new_P1_U3960 = ~P1_DATAWIDTH_REG_28_ & ~P1_DATAWIDTH_REG_29_;
  assign new_P1_U3961 = ~P1_DATAWIDTH_REG_30_ & ~P1_DATAWIDTH_REG_31_;
  assign new_P1_U3962 = new_P1_U3959 & new_P1_U3960 & new_P1_U3961 & new_P1_U6598;
  assign new_P1_U3963 = ~P1_DATAWIDTH_REG_1_ & ~P1_REIP_REG_0_ & ~P1_DATAWIDTH_REG_0_;
  assign new_P1_U3964 = P1_STATE2_REG_2_ & new_P1_U3257;
  assign new_P1_U3965 = new_P1_U6608 & new_P1_U3298;
  assign new_P1_U3966 = ~new_U210 & ~P1_STATE2_REG_0_;
  assign new_P1_U3967 = new_P1_U6602 & new_P1_U3307 & new_P1_U3408;
  assign new_P1_U3968 = P1_STATE2_REG_2_ & new_P1_U3287;
  assign new_P1_U3969 = new_P1_U4235 & new_P1_U4206;
  assign new_P1_U3970 = new_P1_U6618 & new_P1_U6619 & new_P1_U6621 & new_P1_U6620;
  assign new_P1_U3971 = new_P1_U6622 & new_P1_U6623 & new_P1_U6625 & new_P1_U6624;
  assign new_P1_U3972 = new_P1_U6626 & new_P1_U6627 & new_P1_U6629 & new_P1_U6628;
  assign new_P1_U3973 = new_P1_U6630 & new_P1_U6631 & new_P1_U6633 & new_P1_U6632;
  assign new_P1_U3974 = new_P1_U6634 & new_P1_U6635 & new_P1_U6637 & new_P1_U6636;
  assign new_P1_U3975 = new_P1_U6638 & new_P1_U6639 & new_P1_U6641 & new_P1_U6640;
  assign new_P1_U3976 = new_P1_U6642 & new_P1_U6643 & new_P1_U6645 & new_P1_U6644;
  assign new_P1_U3977 = new_P1_U6646 & new_P1_U6647 & new_P1_U6649 & new_P1_U6648;
  assign new_P1_U3978 = new_P1_U6650 & new_P1_U6651 & new_P1_U6653 & new_P1_U6652;
  assign new_P1_U3979 = new_P1_U6654 & new_P1_U6655 & new_P1_U6657 & new_P1_U6656;
  assign new_P1_U3980 = new_P1_U6658 & new_P1_U6659 & new_P1_U6661 & new_P1_U6660;
  assign new_P1_U3981 = new_P1_U6662 & new_P1_U6663 & new_P1_U6665 & new_P1_U6664;
  assign new_P1_U3982 = new_P1_U6666 & new_P1_U6667 & new_P1_U6669 & new_P1_U6668;
  assign new_P1_U3983 = new_P1_U6670 & new_P1_U6671 & new_P1_U6673 & new_P1_U6672;
  assign new_P1_U3984 = new_P1_U6674 & new_P1_U6675 & new_P1_U6677 & new_P1_U6676;
  assign new_P1_U3985 = new_P1_U6678 & new_P1_U6679 & new_P1_U7613 & new_P1_U6680;
  assign new_P1_U3986 = new_P1_U6681 & new_P1_U6682 & new_P1_U6684 & new_P1_U6683;
  assign new_P1_U3987 = new_P1_U6685 & new_P1_U6686 & new_P1_U6688 & new_P1_U6687;
  assign new_P1_U3988 = new_P1_U6689 & new_P1_U6690 & new_P1_U6692 & new_P1_U6691;
  assign new_P1_U3989 = new_P1_U6693 & new_P1_U6694 & new_P1_U6696 & new_P1_U6695;
  assign new_P1_U3990 = new_P1_U6697 & new_P1_U6698 & new_P1_U6700 & new_P1_U6699;
  assign new_P1_U3991 = new_P1_U6701 & new_P1_U6702 & new_P1_U6704 & new_P1_U6703;
  assign new_P1_U3992 = new_P1_U6705 & new_P1_U6706 & new_P1_U6708 & new_P1_U6707;
  assign new_P1_U3993 = new_P1_U6709 & new_P1_U6710 & new_P1_U6712 & new_P1_U6711;
  assign new_P1_U3994 = new_P1_U6713 & new_P1_U6714 & new_P1_U6716 & new_P1_U6715;
  assign new_P1_U3995 = new_P1_U6717 & new_P1_U6718 & new_P1_U6720 & new_P1_U6719;
  assign new_P1_U3996 = new_P1_U6721 & new_P1_U6722 & new_P1_U6724 & new_P1_U6723;
  assign new_P1_U3997 = new_P1_U6725 & new_P1_U6726 & new_P1_U6728 & new_P1_U6727;
  assign new_P1_U3998 = new_P1_U6729 & new_P1_U6730 & new_P1_U6732 & new_P1_U6731;
  assign new_P1_U3999 = new_P1_U6733 & new_P1_U6734 & new_P1_U6736 & new_P1_U6735;
  assign new_P1_U4000 = new_P1_U6737 & new_P1_U6738 & new_P1_U6740 & new_P1_U6739;
  assign new_P1_U4001 = new_P1_U6741 & new_P1_U6742 & new_P1_U6744 & new_P1_U6743;
  assign new_P1_U4002 = new_P1_U6749 & new_P1_U6748;
  assign new_P1_U4003 = new_P1_U6752 & new_P1_U6751;
  assign new_P1_U4004 = new_P1_U6755 & new_P1_U6754;
  assign new_P1_U4005 = new_P1_U6758 & new_P1_U6757;
  assign new_P1_U4006 = new_P1_U6760 & new_P1_U4007;
  assign new_P1_U4007 = new_P1_U6762 & new_P1_U6761;
  assign new_P1_U4008 = new_P1_U6764 & new_P1_U6765;
  assign new_P1_U4009 = new_P1_U6774 & new_P1_U6772 & new_P1_U6773;
  assign new_P1_U4010 = new_P1_U6776 & new_P1_U6777;
  assign new_P1_U4011 = new_P1_U6783 & new_P1_U6781 & new_P1_U6782;
  assign new_P1_U4012 = new_P1_U6787 & new_P1_U6785 & new_P1_U6786;
  assign new_P1_U4013 = new_P1_U6791 & new_P1_U6789 & new_P1_U6790;
  assign new_P1_U4014 = new_P1_U6795 & new_P1_U6793 & new_P1_U6794;
  assign new_P1_U4015 = new_P1_U6799 & new_P1_U6797 & new_P1_U6798;
  assign new_P1_U4016 = new_P1_U6803 & new_P1_U6801 & new_P1_U6802;
  assign new_P1_U4017 = new_P1_U6807 & new_P1_U6805 & new_P1_U6806;
  assign new_P1_U4018 = new_P1_U6811 & new_P1_U6809 & new_P1_U6810;
  assign new_P1_U4019 = new_P1_U6815 & new_P1_U6813 & new_P1_U6814;
  assign new_P1_U4020 = new_P1_U6819 & new_P1_U6817 & new_P1_U6818;
  assign new_P1_U4021 = new_P1_U6821 & new_P1_U6822;
  assign new_P1_U4022 = new_P1_U6828 & new_P1_U6826 & new_P1_U6827;
  assign new_P1_U4023 = new_P1_U6832 & new_P1_U6830 & new_P1_U6831;
  assign new_P1_U4024 = new_P1_U6836 & new_P1_U6834 & new_P1_U6835;
  assign new_P1_U4025 = new_P1_U6840 & new_P1_U6838 & new_P1_U6839;
  assign new_P1_U4026 = new_P1_U6858 & new_P1_U6857;
  assign new_P1_U4027 = new_P1_U6860 & new_P1_U6861;
  assign new_P1_U4028 = new_P1_U3283 & new_P1_U7494 & new_P1_U6888;
  assign new_P1_U4029 = new_P1_U6892 & new_P1_U6893 & new_P1_U6895 & new_P1_U6894;
  assign new_P1_U4030 = new_P1_U6896 & new_P1_U6897 & new_P1_U6899 & new_P1_U6898;
  assign new_P1_U4031 = new_P1_U6900 & new_P1_U6901 & new_P1_U6903 & new_P1_U6902;
  assign new_P1_U4032 = new_P1_U6904 & new_P1_U6905 & new_P1_U6907 & new_P1_U6906;
  assign new_P1_U4033 = new_P1_U6910 & new_P1_U6911 & new_P1_U6913 & new_P1_U6912;
  assign new_P1_U4034 = new_P1_U6914 & new_P1_U6915 & new_P1_U6917 & new_P1_U6916;
  assign new_P1_U4035 = new_P1_U6918 & new_P1_U6919 & new_P1_U6921 & new_P1_U6920;
  assign new_P1_U4036 = new_P1_U6922 & new_P1_U6923 & new_P1_U6925 & new_P1_U6924;
  assign new_P1_U4037 = new_P1_U6941 & new_P1_U6942 & new_P1_U6944 & new_P1_U6943;
  assign new_P1_U4038 = new_P1_U6945 & new_P1_U6946 & new_P1_U6948 & new_P1_U6947;
  assign new_P1_U4039 = new_P1_U6949 & new_P1_U6950 & new_P1_U6952 & new_P1_U6951;
  assign new_P1_U4040 = new_P1_U6953 & new_P1_U6954 & new_P1_U6956 & new_P1_U6955;
  assign new_P1_U4041 = new_P1_U6958 & new_P1_U6959 & new_P1_U6961 & new_P1_U6960;
  assign new_P1_U4042 = new_P1_U6962 & new_P1_U6963 & new_P1_U6965 & new_P1_U6964;
  assign new_P1_U4043 = new_P1_U6966 & new_P1_U6967 & new_P1_U6969 & new_P1_U6968;
  assign new_P1_U4044 = new_P1_U6970 & new_P1_U6971 & new_P1_U6973 & new_P1_U6972;
  assign new_P1_U4045 = new_P1_U6975 & new_P1_U6976 & new_P1_U6978 & new_P1_U6977;
  assign new_P1_U4046 = new_P1_U6979 & new_P1_U6980 & new_P1_U6982 & new_P1_U6981;
  assign new_P1_U4047 = new_P1_U6983 & new_P1_U6984 & new_P1_U6986 & new_P1_U6985;
  assign new_P1_U4048 = new_P1_U6987 & new_P1_U6988 & new_P1_U6990 & new_P1_U6989;
  assign new_P1_U4049 = new_P1_U6992 & new_P1_U6993 & new_P1_U6995 & new_P1_U6994;
  assign new_P1_U4050 = new_P1_U6996 & new_P1_U6997 & new_P1_U6999 & new_P1_U6998;
  assign new_P1_U4051 = new_P1_U7000 & new_P1_U7001 & new_P1_U7003 & new_P1_U7002;
  assign new_P1_U4052 = new_P1_U7004 & new_P1_U7005 & new_P1_U7614 & new_P1_U7006;
  assign new_P1_U4053 = new_P1_U7007 & new_P1_U7008 & new_P1_U7010 & new_P1_U7009;
  assign new_P1_U4054 = new_P1_U7011 & new_P1_U7012 & new_P1_U7014 & new_P1_U7013;
  assign new_P1_U4055 = new_P1_U7015 & new_P1_U7016 & new_P1_U7018 & new_P1_U7017;
  assign new_P1_U4056 = new_P1_U7019 & new_P1_U7020 & new_P1_U7022 & new_P1_U7021;
  assign new_P1_U4057 = new_P1_U7024 & new_P1_U7025 & new_P1_U7027 & new_P1_U7026;
  assign new_P1_U4058 = new_P1_U7028 & new_P1_U7029 & new_P1_U7031 & new_P1_U7030;
  assign new_P1_U4059 = new_P1_U7032 & new_P1_U7033 & new_P1_U7035 & new_P1_U7034;
  assign new_P1_U4060 = new_P1_U7036 & new_P1_U7037 & new_P1_U7039 & new_P1_U7038;
  assign new_P1_U4061 = new_P1_U7059 & new_P1_U3443;
  assign new_P1_U4062 = P1_STATE2_REG_0_ & new_P1_U7062;
  assign new_P1_U4063 = new_P1_U7066 & new_P1_U7067 & new_P1_U7069 & new_P1_U7068;
  assign new_P1_U4064 = new_P1_U7070 & new_P1_U7071 & new_P1_U7073 & new_P1_U7072;
  assign new_P1_U4065 = new_P1_U7074 & new_P1_U7075 & new_P1_U7077 & new_P1_U7076;
  assign new_P1_U4066 = new_P1_U7078 & new_P1_U7079 & new_P1_U7081 & new_P1_U7080;
  assign new_P1_U4067 = new_P1_U4256 & P1_STATE2_REG_0_;
  assign new_P1_U4068 = new_P1_U4401 & new_P1_U4403 & new_P1_U4405 & new_P1_U4404;
  assign new_P1_U4069 = new_P1_U4408 & new_P1_U4407 & new_P1_U4406;
  assign new_P1_U4070 = new_P1_U4409 & new_P1_U4410 & new_P1_U4412 & new_P1_U4411;
  assign new_P1_U4071 = new_P1_U4414 & new_P1_U4413;
  assign new_P1_U4072 = new_P1_U4400 & new_P1_U3391;
  assign new_P1_U4073 = P1_STATE2_REG_0_ & new_P1_U3284;
  assign new_P1_U4074 = new_P1_U7090 & new_P1_U7089;
  assign new_P1_U4075 = new_P1_U7473 & new_P1_U7472 & new_P1_U3434;
  assign new_P1_U4076 = new_P1_U7474 & new_P1_U7475 & new_P1_U7476;
  assign new_P1_U4077 = new_P1_U4076 & new_P1_U2606 & new_P1_U7477;
  assign new_P1_U4078 = new_P1_U7097 & new_P1_U7095;
  assign new_P1_U4079 = new_P1_U7098 & new_P1_U7099 & new_P1_U7101 & new_P1_U7100;
  assign new_P1_U4080 = new_P1_U7102 & new_P1_U7103 & new_P1_U7105 & new_P1_U7104;
  assign new_P1_U4081 = new_P1_U7106 & new_P1_U7107 & new_P1_U7109 & new_P1_U7108;
  assign new_P1_U4082 = new_P1_U7110 & new_P1_U7111 & new_P1_U7113 & new_P1_U7112;
  assign new_P1_U4083 = new_P1_U7115 & new_P1_U7116 & new_P1_U7118 & new_P1_U7117;
  assign new_P1_U4084 = new_P1_U7119 & new_P1_U7120 & new_P1_U7122 & new_P1_U7121;
  assign new_P1_U4085 = new_P1_U7123 & new_P1_U7124 & new_P1_U7126 & new_P1_U7125;
  assign new_P1_U4086 = new_P1_U7127 & new_P1_U7128 & new_P1_U7130 & new_P1_U7129;
  assign new_P1_U4087 = new_P1_U7132 & new_P1_U7133 & new_P1_U7135 & new_P1_U7134;
  assign new_P1_U4088 = new_P1_U7136 & new_P1_U7137 & new_P1_U7139 & new_P1_U7138;
  assign new_P1_U4089 = new_P1_U7140 & new_P1_U7141 & new_P1_U7143 & new_P1_U7142;
  assign new_P1_U4090 = new_P1_U7145 & new_P1_U7144;
  assign new_P1_U4091 = new_P1_U4090 & new_P1_U7617 & new_P1_U7146;
  assign new_P1_U4092 = new_P1_U7147 & new_P1_U7148 & new_P1_U7150 & new_P1_U7149;
  assign new_P1_U4093 = new_P1_U7151 & new_P1_U7152 & new_P1_U7154 & new_P1_U7153;
  assign new_P1_U4094 = new_P1_U7155 & new_P1_U7156 & new_P1_U7158 & new_P1_U7157;
  assign new_P1_U4095 = new_P1_U7159 & new_P1_U7160 & new_P1_U7162 & new_P1_U7161;
  assign new_P1_U4096 = new_P1_U7164 & new_P1_U7165 & new_P1_U7167 & new_P1_U7166;
  assign new_P1_U4097 = new_P1_U7168 & new_P1_U7169 & new_P1_U7171 & new_P1_U7170;
  assign new_P1_U4098 = new_P1_U7172 & new_P1_U7173 & new_P1_U7175 & new_P1_U7174;
  assign new_P1_U4099 = new_P1_U7176 & new_P1_U7177 & new_P1_U7179 & new_P1_U7178;
  assign new_P1_U4100 = new_P1_U7181 & new_P1_U7182 & new_P1_U7184 & new_P1_U7183;
  assign new_P1_U4101 = new_P1_U7185 & new_P1_U7186 & new_P1_U7188 & new_P1_U7187;
  assign new_P1_U4102 = new_P1_U7189 & new_P1_U7190 & new_P1_U7192 & new_P1_U7191;
  assign new_P1_U4103 = new_P1_U7193 & new_P1_U7194 & new_P1_U7196 & new_P1_U7195;
  assign new_P1_U4104 = new_P1_U7198 & new_P1_U7199 & new_P1_U7201 & new_P1_U7200;
  assign new_P1_U4105 = new_P1_U7202 & new_P1_U7203 & new_P1_U7205 & new_P1_U7204;
  assign new_P1_U4106 = new_P1_U7206 & new_P1_U7207 & new_P1_U7209 & new_P1_U7208;
  assign new_P1_U4107 = new_P1_U7210 & new_P1_U7211 & new_P1_U7213 & new_P1_U7212;
  assign new_P1_U4108 = new_P1_U7215 & new_P1_U3264;
  assign new_P1_U4109 = new_P1_U7216 & new_P1_U7215;
  assign new_P1_U4110 = new_P1_U7217 & new_P1_U3265;
  assign new_P1_U4111 = new_P1_U7089 & new_P1_U3427;
  assign new_P1_U4112 = new_P1_U7218 & new_P1_U7217;
  assign new_P1_U4113 = new_P1_U7473 & new_P1_U4112 & new_P1_U7472;
  assign new_P1_U4114 = new_P1_U4113 & new_P1_U4111 & new_P1_U7090 & new_P1_U3434;
  assign new_P1_U4115 = new_P1_U7474 & new_P1_U7476 & new_P1_U7486 & new_P1_U7480;
  assign new_P1_U4116 = new_P1_U7487 & new_P1_U7488 & new_P1_U7505 & new_P1_U7489;
  assign new_P1_U4117 = new_P1_U7090 & new_P1_U7089;
  assign new_P1_U4118 = new_P1_U7473 & new_P1_U7472 & new_P1_U3434;
  assign new_P1_U4119 = new_P1_U7474 & new_P1_U7475 & new_P1_U7476;
  assign new_P1_U4120 = new_P1_U4119 & new_P1_U2606 & new_P1_U2608 & new_P1_U7477;
  assign new_P1_U4121 = new_P1_U7220 & new_P1_U7221 & new_P1_U7223 & new_P1_U7222;
  assign new_P1_U4122 = new_P1_U7224 & new_P1_U7225 & new_P1_U7227 & new_P1_U7226;
  assign new_P1_U4123 = new_P1_U7228 & new_P1_U7229 & new_P1_U7231 & new_P1_U7230;
  assign new_P1_U4124 = new_P1_U7232 & new_P1_U7233 & new_P1_U7235 & new_P1_U7234;
  assign new_P1_U4125 = new_P1_U7237 & new_P1_U7238 & new_P1_U7240 & new_P1_U7239;
  assign new_P1_U4126 = new_P1_U7241 & new_P1_U7242 & new_P1_U7244 & new_P1_U7243;
  assign new_P1_U4127 = new_P1_U7245 & new_P1_U7246 & new_P1_U7248 & new_P1_U7247;
  assign new_P1_U4128 = new_P1_U7249 & new_P1_U7250 & new_P1_U7252 & new_P1_U7251;
  assign new_P1_U4129 = new_P1_U7254 & new_P1_U7255 & new_P1_U7257 & new_P1_U7256;
  assign new_P1_U4130 = new_P1_U7258 & new_P1_U7259 & new_P1_U7261 & new_P1_U7260;
  assign new_P1_U4131 = new_P1_U7262 & new_P1_U7263 & new_P1_U7265 & new_P1_U7264;
  assign new_P1_U4132 = new_P1_U7266 & new_P1_U7267 & new_P1_U7269 & new_P1_U7268;
  assign new_P1_U4133 = new_P1_U7271 & new_P1_U7272 & new_P1_U7274 & new_P1_U7273;
  assign new_P1_U4134 = new_P1_U7275 & new_P1_U7276 & new_P1_U7278 & new_P1_U7277;
  assign new_P1_U4135 = new_P1_U7279 & new_P1_U7280 & new_P1_U7282 & new_P1_U7281;
  assign new_P1_U4136 = new_P1_U7283 & new_P1_U7284 & new_P1_U7619 & new_P1_U7285;
  assign new_P1_U4137 = new_P1_U7286 & new_P1_U7287 & new_P1_U7289 & new_P1_U7288;
  assign new_P1_U4138 = new_P1_U7290 & new_P1_U7291 & new_P1_U7293 & new_P1_U7292;
  assign new_P1_U4139 = new_P1_U7294 & new_P1_U7295 & new_P1_U7297 & new_P1_U7296;
  assign new_P1_U4140 = new_P1_U7298 & new_P1_U7299 & new_P1_U7301 & new_P1_U7300;
  assign new_P1_U4141 = new_P1_U7303 & new_P1_U7304 & new_P1_U7306 & new_P1_U7305;
  assign new_P1_U4142 = new_P1_U7307 & new_P1_U7308 & new_P1_U7310 & new_P1_U7309;
  assign new_P1_U4143 = new_P1_U7311 & new_P1_U7312 & new_P1_U7314 & new_P1_U7313;
  assign new_P1_U4144 = new_P1_U7315 & new_P1_U7316 & new_P1_U7318 & new_P1_U7317;
  assign new_P1_U4145 = new_P1_U7320 & new_P1_U7321 & new_P1_U7323 & new_P1_U7322;
  assign new_P1_U4146 = new_P1_U7324 & new_P1_U7325 & new_P1_U7327 & new_P1_U7326;
  assign new_P1_U4147 = new_P1_U7328 & new_P1_U7329 & new_P1_U7331 & new_P1_U7330;
  assign new_P1_U4148 = new_P1_U7332 & new_P1_U7333 & new_P1_U7335 & new_P1_U7334;
  assign new_P1_U4149 = new_P1_U7337 & new_P1_U7338 & new_P1_U7340 & new_P1_U7339;
  assign new_P1_U4150 = new_P1_U7341 & new_P1_U7342 & new_P1_U7344 & new_P1_U7343;
  assign new_P1_U4151 = new_P1_U7345 & new_P1_U7346 & new_P1_U7348 & new_P1_U7347;
  assign new_P1_U4152 = new_P1_U7349 & new_P1_U7350 & new_P1_U7352 & new_P1_U7351;
  assign new_P1_U4153 = new_P1_U3284 & new_P1_U3419;
  assign new_P1_U4154 = new_P1_U3283 & new_P1_U3391;
  assign new_P1_U4155 = new_P1_U4263 & new_P1_U7357 & new_P1_U7358;
  assign new_P1_U4156 = new_P1_U4155 & new_P1_U7359;
  assign new_P1_U4157 = P1_STATE2_REG_0_ & new_P1_U2427;
  assign new_P1_U4158 = new_P1_U4157 & new_P1_U7360;
  assign new_P1_U4159 = new_P1_U3271 & new_P1_U4173;
  assign new_P1_U4160 = P1_STATE2_REG_0_ & new_P1_U4173;
  assign new_P1_U4161 = new_P1_U7369 & P1_STATE2_REG_0_;
  assign new_P1_U4162 = new_P1_U7371 & new_P1_U2603;
  assign new_P1_U4163 = new_P1_U7373 & P1_STATE2_REG_0_;
  assign new_P1_U4164 = new_P1_U7375 & new_P1_U2603;
  assign new_P1_U4165 = new_P1_U7382 & new_P1_U7383;
  assign new_P1_U4166 = new_P1_U3453 & new_P1_U7384;
  assign new_P1_U4167 = new_P1_U7387 & new_P1_U7389 & new_P1_U7388;
  assign new_P1_U4168 = new_P1_U7462 & new_P1_U7461;
  assign new_P1_U4169 = new_P1_U7465 & new_P1_U7464;
  assign new_P1_U4170 = new_P1_U7674 & new_P1_U7673;
  assign new_P1_U4171 = ~new_P1_U3569 | ~new_P1_U3570 | ~new_P1_U3572 | ~new_P1_U3571;
  assign new_P1_U4172 = ~new_P1_U3739 | ~new_P1_U5474;
  assign new_P1_U4173 = ~new_P1_U3573 | ~new_P1_U3574 | ~new_P1_U3575 | ~new_P1_U3576 | ~new_P1_U2607;
  assign new_P1_U4174 = ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_U4175 = new_P1_U7726 & new_P1_U7725;
  assign new_P1_U4176 = new_P1_U7745 & new_P1_U7744;
  assign new_P1_U4177 = ~new_P1_U2368 | ~new_P1_U3285;
  assign new_P1_U4178 = ~new_P1_U4508 | ~new_P1_U3391;
  assign new_P1_U4179 = ~BS16;
  assign new_P1_U4180 = ~new_P1_U3967 | ~new_P1_U4228;
  assign new_P1_U4181 = ~new_P1_U4228 | ~new_P1_U3432;
  assign new_P1_U4182 = ~new_P1_U3738 | ~new_P1_U7698 | ~new_P1_U7697;
  assign new_P1_U4183 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3269;
  assign new_P1_U4184 = ~new_P1_U3452;
  assign new_P1_U4185 = ~HOLD | ~new_P1_U3257;
  assign new_P1_U4186 = ~new_P1_U3412;
  assign new_P1_U4187 = ~new_P1_U3440;
  assign new_P1_U4188 = ~new_P1_U3439;
  assign new_P1_U4189 = ~new_P1_U3393;
  assign new_P1_U4190 = ~new_P1_U3290;
  assign new_P1_U4191 = ~new_P1_U3449;
  assign new_P1_U4192 = ~new_P1_U3405;
  assign new_P1_U4193 = ~new_P1_U3434;
  assign new_P1_U4194 = ~new_P1_U3420;
  assign new_P1_U4195 = ~new_P1_U4265 | ~new_P1_U3271;
  assign new_P1_U4196 = ~new_P1_U4460 | ~new_P1_U2605;
  assign new_P1_U4197 = ~new_P1_U3396;
  assign new_P1_U4198 = ~new_P1_U3425;
  assign new_P1_U4199 = ~new_P1_U3289;
  assign new_P1_U4200 = ~new_P1_U3421;
  assign new_P1_U4201 = ~new_P1_U3422;
  assign new_P1_U4202 = ~new_P1_U3428;
  assign new_P1_U4203 = ~new_P1_U3408;
  assign new_P1_U4204 = ~new_P1_U3427;
  assign new_P1_U4205 = ~new_P1_U4197 | ~new_P1_U3885 | ~new_P1_U4189;
  assign new_P1_U4206 = ~new_P1_U3418;
  assign new_P1_U4207 = ~new_P1_U3443;
  assign new_P1_U4208 = ~new_P1_U3282;
  assign new_P1_U4209 = ~new_P1_U3307;
  assign new_P1_U4210 = ~new_P1_U3390;
  assign new_P1_U4211 = ~new_P1_U3446;
  assign new_P1_U4212 = ~new_P1_U3447;
  assign new_P1_U4213 = ~new_P1_U3448;
  assign new_P1_U4214 = ~new_P1_U3400;
  assign new_P1_U4215 = ~new_P1_U3288;
  assign new_P1_U4216 = ~new_P1_U3292;
  assign new_P1_U4217 = ~new_P1_U3578 | ~new_P1_U2431;
  assign new_P1_U4218 = ~new_P1_U3399;
  assign new_P1_U4219 = ~new_P1_U4449 | ~new_P1_U3271;
  assign new_P1_U4220 = ~new_P1_U3433;
  assign new_P1_U4221 = ~new_P1_U3249;
  assign new_P1_U4222 = ~new_P1_U3426;
  assign new_P1_U4223 = ~new_P1_U3424;
  assign new_P1_U4224 = ~new_P1_U3300;
  assign new_P1_U4225 = ~new_P1_LT_563_1260_U6;
  assign new_P1_U4226 = ~new_P1_U3320;
  assign new_P1_U4227 = ~new_P1_U4255 | ~new_P1_U3431;
  assign new_P1_U4228 = ~new_P1_U4235 | ~new_P1_U7500;
  assign new_P1_U4229 = ~new_P1_U2362 | ~new_P1_U3272;
  assign new_P1_U4230 = ~new_P1_U2363 | ~new_P1_U4377;
  assign new_P1_U4231 = ~new_P1_U3407;
  assign new_P1_U4232 = ~new_P1_U3252;
  assign new_P1_U4233 = ~new_P1_U3250;
  assign new_P1_U4234 = ~new_P1_U3395;
  assign new_P1_U4235 = ~new_P1_U3297;
  assign new_P1_U4236 = ~new_P1_U3398;
  assign new_P1_U4237 = ~new_P1_U4178;
  assign new_P1_U4238 = ~new_P1_U3357;
  assign new_P1_U4239 = ~new_P1_U4477 | ~new_P1_U7381;
  assign new_P1_U4240 = ~new_P1_U3963 | ~new_P1_U4220;
  assign new_P1_U4241 = ~new_P1_U3584 | ~new_P1_U4261;
  assign new_P1_U4242 = ~new_P1_U3731 | ~new_P1_U2428;
  assign new_P1_U4243 = ~new_P1_U4364 | ~new_P1_U3258;
  assign new_P1_U4244 = ~new_P1_U2352 | ~P1_STATE2_REG_1_ | ~new_P1_U3294;
  assign new_P1_U4245 = ~new_P1_U2428 | ~new_P1_U3403;
  assign new_P1_U4246 = ~new_U210 | ~P1_STATE2_REG_0_ | ~new_P1_U3263;
  assign new_P1_U4247 = ~new_P1_U3394;
  assign new_P1_U4248 = ~new_P1_U2448 | ~new_P1_U3862 | ~new_P1_U2451 | ~new_P1_U2353;
  assign new_P1_U4249 = ~new_P1_U3287;
  assign new_P1_U4250 = ~new_P1_U3397;
  assign new_P1_U4251 = ~new_P1_U3415;
  assign new_P1_U4252 = ~new_P1_U3299;
  assign new_P1_U4253 = ~new_P1_U3409;
  assign new_P1_U4254 = ~new_P1_U3419;
  assign new_P1_U4255 = ~new_P1_U3432;
  assign new_P1_U4256 = ~new_P1_U3291;
  assign new_P1_U4257 = ~new_P1_U3389;
  assign new_P1_U4258 = ~new_P1_U3254;
  assign new_P1_U4259 = ~new_P1_U3281;
  assign new_P1_U4260 = ~new_P1_U3406;
  assign new_P1_U4261 = ~new_P1_U3298;
  assign new_P1_U4262 = ~new_P1_U3286;
  assign new_P1_U4263 = ~new_P1_U4236 | ~new_P1_U4399;
  assign new_P1_U4264 = ~new_P1_U3411;
  assign new_P1_U4265 = ~new_P1_U3453;
  assign new_P1_U4266 = ~new_P1_U3410;
  assign new_P1_U4267 = ~P1_REIP_REG_31_ | ~new_P1_U4233;
  assign new_P1_U4268 = ~P1_REIP_REG_30_ | ~new_P1_U4232;
  assign new_P1_U4269 = ~P1_ADDRESS_REG_29_ | ~new_P1_U3249;
  assign new_P1_U4270 = ~P1_REIP_REG_30_ | ~new_P1_U4233;
  assign new_P1_U4271 = ~P1_REIP_REG_29_ | ~new_P1_U4232;
  assign new_P1_U4272 = ~P1_ADDRESS_REG_28_ | ~new_P1_U3249;
  assign new_P1_U4273 = ~P1_REIP_REG_29_ | ~new_P1_U4233;
  assign new_P1_U4274 = ~P1_REIP_REG_28_ | ~new_P1_U4232;
  assign new_P1_U4275 = ~P1_ADDRESS_REG_27_ | ~new_P1_U3249;
  assign new_P1_U4276 = ~P1_REIP_REG_28_ | ~new_P1_U4233;
  assign new_P1_U4277 = ~P1_REIP_REG_27_ | ~new_P1_U4232;
  assign new_P1_U4278 = ~P1_ADDRESS_REG_26_ | ~new_P1_U3249;
  assign new_P1_U4279 = ~P1_REIP_REG_27_ | ~new_P1_U4233;
  assign new_P1_U4280 = ~P1_REIP_REG_26_ | ~new_P1_U4232;
  assign new_P1_U4281 = ~P1_ADDRESS_REG_25_ | ~new_P1_U3249;
  assign new_P1_U4282 = ~P1_REIP_REG_26_ | ~new_P1_U4233;
  assign new_P1_U4283 = ~P1_REIP_REG_25_ | ~new_P1_U4232;
  assign new_P1_U4284 = ~P1_ADDRESS_REG_24_ | ~new_P1_U3249;
  assign new_P1_U4285 = ~P1_REIP_REG_25_ | ~new_P1_U4233;
  assign new_P1_U4286 = ~P1_REIP_REG_24_ | ~new_P1_U4232;
  assign new_P1_U4287 = ~P1_ADDRESS_REG_23_ | ~new_P1_U3249;
  assign new_P1_U4288 = ~P1_REIP_REG_24_ | ~new_P1_U4233;
  assign new_P1_U4289 = ~P1_REIP_REG_23_ | ~new_P1_U4232;
  assign new_P1_U4290 = ~P1_ADDRESS_REG_22_ | ~new_P1_U3249;
  assign new_P1_U4291 = ~P1_REIP_REG_23_ | ~new_P1_U4233;
  assign new_P1_U4292 = ~P1_REIP_REG_22_ | ~new_P1_U4232;
  assign new_P1_U4293 = ~P1_ADDRESS_REG_21_ | ~new_P1_U3249;
  assign new_P1_U4294 = ~P1_REIP_REG_22_ | ~new_P1_U4233;
  assign new_P1_U4295 = ~P1_REIP_REG_21_ | ~new_P1_U4232;
  assign new_P1_U4296 = ~P1_ADDRESS_REG_20_ | ~new_P1_U3249;
  assign new_P1_U4297 = ~P1_REIP_REG_21_ | ~new_P1_U4233;
  assign new_P1_U4298 = ~P1_REIP_REG_20_ | ~new_P1_U4232;
  assign new_P1_U4299 = ~P1_ADDRESS_REG_19_ | ~new_P1_U3249;
  assign new_P1_U4300 = ~P1_REIP_REG_20_ | ~new_P1_U4233;
  assign new_P1_U4301 = ~P1_REIP_REG_19_ | ~new_P1_U4232;
  assign new_P1_U4302 = ~P1_ADDRESS_REG_18_ | ~new_P1_U3249;
  assign new_P1_U4303 = ~P1_REIP_REG_19_ | ~new_P1_U4233;
  assign new_P1_U4304 = ~P1_REIP_REG_18_ | ~new_P1_U4232;
  assign new_P1_U4305 = ~P1_ADDRESS_REG_17_ | ~new_P1_U3249;
  assign new_P1_U4306 = ~P1_REIP_REG_18_ | ~new_P1_U4233;
  assign new_P1_U4307 = ~P1_REIP_REG_17_ | ~new_P1_U4232;
  assign new_P1_U4308 = ~P1_ADDRESS_REG_16_ | ~new_P1_U3249;
  assign new_P1_U4309 = ~P1_REIP_REG_17_ | ~new_P1_U4233;
  assign new_P1_U4310 = ~P1_REIP_REG_16_ | ~new_P1_U4232;
  assign new_P1_U4311 = ~P1_ADDRESS_REG_15_ | ~new_P1_U3249;
  assign new_P1_U4312 = ~P1_REIP_REG_16_ | ~new_P1_U4233;
  assign new_P1_U4313 = ~P1_REIP_REG_15_ | ~new_P1_U4232;
  assign new_P1_U4314 = ~P1_ADDRESS_REG_14_ | ~new_P1_U3249;
  assign new_P1_U4315 = ~P1_REIP_REG_15_ | ~new_P1_U4233;
  assign new_P1_U4316 = ~P1_REIP_REG_14_ | ~new_P1_U4232;
  assign new_P1_U4317 = ~P1_ADDRESS_REG_13_ | ~new_P1_U3249;
  assign new_P1_U4318 = ~P1_REIP_REG_14_ | ~new_P1_U4233;
  assign new_P1_U4319 = ~P1_REIP_REG_13_ | ~new_P1_U4232;
  assign new_P1_U4320 = ~P1_ADDRESS_REG_12_ | ~new_P1_U3249;
  assign new_P1_U4321 = ~P1_REIP_REG_13_ | ~new_P1_U4233;
  assign new_P1_U4322 = ~P1_REIP_REG_12_ | ~new_P1_U4232;
  assign new_P1_U4323 = ~P1_ADDRESS_REG_11_ | ~new_P1_U3249;
  assign new_P1_U4324 = ~P1_REIP_REG_12_ | ~new_P1_U4233;
  assign new_P1_U4325 = ~P1_REIP_REG_11_ | ~new_P1_U4232;
  assign new_P1_U4326 = ~P1_ADDRESS_REG_10_ | ~new_P1_U3249;
  assign new_P1_U4327 = ~P1_REIP_REG_11_ | ~new_P1_U4233;
  assign new_P1_U4328 = ~P1_REIP_REG_10_ | ~new_P1_U4232;
  assign new_P1_U4329 = ~P1_ADDRESS_REG_9_ | ~new_P1_U3249;
  assign new_P1_U4330 = ~P1_REIP_REG_10_ | ~new_P1_U4233;
  assign new_P1_U4331 = ~P1_REIP_REG_9_ | ~new_P1_U4232;
  assign new_P1_U4332 = ~P1_ADDRESS_REG_8_ | ~new_P1_U3249;
  assign new_P1_U4333 = ~P1_REIP_REG_9_ | ~new_P1_U4233;
  assign new_P1_U4334 = ~P1_REIP_REG_8_ | ~new_P1_U4232;
  assign new_P1_U4335 = ~P1_ADDRESS_REG_7_ | ~new_P1_U3249;
  assign new_P1_U4336 = ~P1_REIP_REG_8_ | ~new_P1_U4233;
  assign new_P1_U4337 = ~P1_REIP_REG_7_ | ~new_P1_U4232;
  assign new_P1_U4338 = ~P1_ADDRESS_REG_6_ | ~new_P1_U3249;
  assign new_P1_U4339 = ~P1_REIP_REG_7_ | ~new_P1_U4233;
  assign new_P1_U4340 = ~P1_REIP_REG_6_ | ~new_P1_U4232;
  assign new_P1_U4341 = ~P1_ADDRESS_REG_5_ | ~new_P1_U3249;
  assign new_P1_U4342 = ~P1_REIP_REG_6_ | ~new_P1_U4233;
  assign new_P1_U4343 = ~P1_REIP_REG_5_ | ~new_P1_U4232;
  assign new_P1_U4344 = ~P1_ADDRESS_REG_4_ | ~new_P1_U3249;
  assign new_P1_U4345 = ~P1_REIP_REG_5_ | ~new_P1_U4233;
  assign new_P1_U4346 = ~P1_REIP_REG_4_ | ~new_P1_U4232;
  assign new_P1_U4347 = ~P1_ADDRESS_REG_3_ | ~new_P1_U3249;
  assign new_P1_U4348 = ~P1_REIP_REG_4_ | ~new_P1_U4233;
  assign new_P1_U4349 = ~P1_REIP_REG_3_ | ~new_P1_U4232;
  assign new_P1_U4350 = ~P1_ADDRESS_REG_2_ | ~new_P1_U3249;
  assign new_P1_U4351 = ~P1_REIP_REG_3_ | ~new_P1_U4233;
  assign new_P1_U4352 = ~P1_REIP_REG_2_ | ~new_P1_U4232;
  assign new_P1_U4353 = ~P1_ADDRESS_REG_1_ | ~new_P1_U3249;
  assign new_P1_U4354 = ~P1_REIP_REG_2_ | ~new_P1_U4233;
  assign new_P1_U4355 = ~P1_REIP_REG_1_ | ~new_P1_U4232;
  assign new_P1_U4356 = ~P1_ADDRESS_REG_0_ | ~new_P1_U3249;
  assign new_P1_U4357 = ~new_P1_U3260;
  assign new_P1_U4358 = ~new_P1_U4357 | ~new_P1_U3257;
  assign new_P1_U4359 = ~NA | ~new_P1_U4258;
  assign new_P1_U4360 = ~new_P1_U3261;
  assign new_P1_U4361 = ~new_P1_U4360 | ~new_P1_U3257;
  assign new_P1_U4362 = P1_STATE_REG_0_ | NA;
  assign new_P1_U4363 = ~new_P1_U7623 | ~new_P1_U7622 | ~new_P1_U4362;
  assign new_P1_U4364 = ~new_P1_U3255;
  assign new_P1_U4365 = ~new_P1_U4364 | ~HOLD | ~new_P1_U3247;
  assign new_P1_U4366 = ~new_U210 | ~P1_STATE_REG_1_ | ~new_P1_U3261;
  assign new_P1_U4367 = ~new_P1_U4366 | ~new_P1_U4365;
  assign new_P1_U4368 = ~new_P1_U4367 | ~P1_STATE_REG_0_ | ~new_P1_U4359;
  assign new_P1_U4369 = ~P1_STATE_REG_2_ | ~new_P1_U4363;
  assign new_P1_U4370 = ~new_U210 | ~new_P1_U4221;
  assign new_P1_U4371 = ~new_P1_U3496 | ~new_P1_U7625;
  assign new_P1_U4372 = ~P1_STATE_REG_2_ | ~new_P1_U3260;
  assign new_P1_U4373 = ~NA | ~new_P1_U3258;
  assign new_P1_U4374 = ~new_P1_U4373 | ~new_P1_U4372;
  assign new_P1_U4375 = ~new_P1_U4374 | ~new_P1_U3248;
  assign new_P1_U4376 = ~new_P1_U4179 | ~new_P1_U3255;
  assign new_P1_U4377 = ~new_P1_U3280;
  assign new_P1_U4378 = ~new_P1_U3269;
  assign new_P1_U4379 = ~new_P1_U3444;
  assign new_P1_U4380 = ~new_P1_U3268;
  assign new_P1_U4381 = ~new_P1_U3274;
  assign new_P1_U4382 = ~new_P1_U3267;
  assign new_P1_U4383 = ~P1_INSTQUEUE_REG_7__3_ | ~new_P1_U4382;
  assign new_P1_U4384 = ~P1_INSTQUEUE_REG_0__3_ | ~new_P1_U2472;
  assign new_P1_U4385 = ~P1_INSTQUEUE_REG_1__3_ | ~new_P1_U2471;
  assign new_P1_U4386 = ~P1_INSTQUEUE_REG_2__3_ | ~new_P1_U2470;
  assign new_P1_U4387 = ~P1_INSTQUEUE_REG_3__3_ | ~new_P1_U2468;
  assign new_P1_U4388 = ~P1_INSTQUEUE_REG_4__3_ | ~new_P1_U2467;
  assign new_P1_U4389 = ~P1_INSTQUEUE_REG_5__3_ | ~new_P1_U2466;
  assign new_P1_U4390 = ~P1_INSTQUEUE_REG_6__3_ | ~new_P1_U2465;
  assign new_P1_U4391 = ~P1_INSTQUEUE_REG_8__3_ | ~new_P1_U2464;
  assign new_P1_U4392 = ~P1_INSTQUEUE_REG_9__3_ | ~new_P1_U2463;
  assign new_P1_U4393 = ~P1_INSTQUEUE_REG_10__3_ | ~new_P1_U2461;
  assign new_P1_U4394 = ~P1_INSTQUEUE_REG_11__3_ | ~new_P1_U2459;
  assign new_P1_U4395 = ~P1_INSTQUEUE_REG_12__3_ | ~new_P1_U2458;
  assign new_P1_U4396 = ~P1_INSTQUEUE_REG_13__3_ | ~new_P1_U2457;
  assign new_P1_U4397 = ~P1_INSTQUEUE_REG_14__3_ | ~new_P1_U2455;
  assign new_P1_U4398 = ~P1_INSTQUEUE_REG_15__3_ | ~new_P1_U2453;
  assign new_P1_U4399 = ~new_P1_U3283;
  assign new_P1_U4400 = ~new_P1_U3278;
  assign new_P1_U4401 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUE_REG_7__5_ | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3270;
  assign new_P1_U4402 = ~new_P1_U4380 | ~P1_INSTQUEUE_REG_0__5_ | ~new_P1_U3270;
  assign new_P1_U4403 = ~new_P1_U3265 | ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUE_REG_1__5_ | ~new_P1_U2469;
  assign new_P1_U4404 = ~new_P1_U3266 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_2__5_ | ~new_P1_U2469;
  assign new_P1_U4405 = ~new_P1_U3270 | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~P1_INSTQUEUE_REG_4__5_ | ~new_P1_U4378;
  assign new_P1_U4406 = ~new_P1_U3521 | ~new_P1_U3520 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U4407 = ~new_P1_U3523 | ~new_P1_U3522 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U4408 = ~new_P1_U3524 | ~new_P1_U4380;
  assign new_P1_U4409 = ~new_P1_U3526 | ~new_P1_U3525 | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U4410 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~P1_INSTQUEUE_REG_11__5_ | ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3264;
  assign new_P1_U4411 = ~new_P1_U3527 | ~new_P1_U4378 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U4412 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~P1_INSTQUEUE_REG_13__5_ | ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3265;
  assign new_P1_U4413 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~P1_INSTQUEUE_REG_14__5_ | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3266;
  assign new_P1_U4414 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~P1_INSTQUEUE_REG_15__5_ | ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U4415 = ~new_P1_U4173;
  assign new_P1_U4416 = ~P1_INSTQUEUE_REG_7__2_ | ~new_P1_U4382;
  assign new_P1_U4417 = ~P1_INSTQUEUE_REG_0__2_ | ~new_P1_U2472;
  assign new_P1_U4418 = ~P1_INSTQUEUE_REG_1__2_ | ~new_P1_U2471;
  assign new_P1_U4419 = ~P1_INSTQUEUE_REG_2__2_ | ~new_P1_U2470;
  assign new_P1_U4420 = ~P1_INSTQUEUE_REG_3__2_ | ~new_P1_U2468;
  assign new_P1_U4421 = ~P1_INSTQUEUE_REG_4__2_ | ~new_P1_U2467;
  assign new_P1_U4422 = ~P1_INSTQUEUE_REG_5__2_ | ~new_P1_U2466;
  assign new_P1_U4423 = ~P1_INSTQUEUE_REG_6__2_ | ~new_P1_U2465;
  assign new_P1_U4424 = ~P1_INSTQUEUE_REG_8__2_ | ~new_P1_U2464;
  assign new_P1_U4425 = ~P1_INSTQUEUE_REG_9__2_ | ~new_P1_U2463;
  assign new_P1_U4426 = ~P1_INSTQUEUE_REG_10__2_ | ~new_P1_U2461;
  assign new_P1_U4427 = ~P1_INSTQUEUE_REG_11__2_ | ~new_P1_U2459;
  assign new_P1_U4428 = ~P1_INSTQUEUE_REG_12__2_ | ~new_P1_U2458;
  assign new_P1_U4429 = ~P1_INSTQUEUE_REG_13__2_ | ~new_P1_U2457;
  assign new_P1_U4430 = ~P1_INSTQUEUE_REG_14__2_ | ~new_P1_U2455;
  assign new_P1_U4431 = ~P1_INSTQUEUE_REG_15__2_ | ~new_P1_U2453;
  assign new_P1_U4432 = ~new_P1_U4171;
  assign new_P1_U4433 = ~P1_INSTQUEUE_REG_7__7_ | ~new_P1_U4382;
  assign new_P1_U4434 = ~P1_INSTQUEUE_REG_0__7_ | ~new_P1_U2472;
  assign new_P1_U4435 = ~P1_INSTQUEUE_REG_1__7_ | ~new_P1_U2471;
  assign new_P1_U4436 = ~P1_INSTQUEUE_REG_2__7_ | ~new_P1_U2470;
  assign new_P1_U4437 = ~P1_INSTQUEUE_REG_3__7_ | ~new_P1_U2468;
  assign new_P1_U4438 = ~P1_INSTQUEUE_REG_4__7_ | ~new_P1_U2467;
  assign new_P1_U4439 = ~P1_INSTQUEUE_REG_5__7_ | ~new_P1_U2466;
  assign new_P1_U4440 = ~P1_INSTQUEUE_REG_6__7_ | ~new_P1_U2465;
  assign new_P1_U4441 = ~P1_INSTQUEUE_REG_8__7_ | ~new_P1_U2464;
  assign new_P1_U4442 = ~P1_INSTQUEUE_REG_9__7_ | ~new_P1_U2463;
  assign new_P1_U4443 = ~P1_INSTQUEUE_REG_10__7_ | ~new_P1_U2461;
  assign new_P1_U4444 = ~P1_INSTQUEUE_REG_11__7_ | ~new_P1_U2459;
  assign new_P1_U4445 = ~P1_INSTQUEUE_REG_12__7_ | ~new_P1_U2458;
  assign new_P1_U4446 = ~P1_INSTQUEUE_REG_13__7_ | ~new_P1_U2457;
  assign new_P1_U4447 = ~P1_INSTQUEUE_REG_14__7_ | ~new_P1_U2455;
  assign new_P1_U4448 = ~P1_INSTQUEUE_REG_15__7_ | ~new_P1_U2453;
  assign new_P1_U4449 = ~new_P1_U3391;
  assign new_P1_U4450 = ~P1_INSTQUEUE_REG_7__6_ | ~new_P1_U3498 | ~new_P1_U4381;
  assign new_P1_U4451 = ~new_P1_U2456 | ~P1_INSTQUEUE_REG_1__6_ | ~new_P1_U2469;
  assign new_P1_U4452 = ~new_P1_U2454 | ~P1_INSTQUEUE_REG_2__6_ | ~new_P1_U2469;
  assign new_P1_U4453 = ~new_P1_U4381 | ~P1_INSTQUEUE_REG_4__6_ | ~new_P1_U4378;
  assign new_P1_U4454 = ~P1_INSTQUEUE_REG_5__6_ | ~new_P1_U2456 | ~new_P1_U4381;
  assign new_P1_U4455 = ~P1_INSTQUEUE_REG_6__6_ | ~new_P1_U2454 | ~new_P1_U4381;
  assign new_P1_U4456 = ~new_P1_U3507 | ~P1_INSTQUEUE_REG_12__6_ | ~new_P1_U4378;
  assign new_P1_U4457 = ~P1_INSTQUEUE_REG_13__6_ | ~new_P1_U3507 | ~new_P1_U2456;
  assign new_P1_U4458 = ~P1_INSTQUEUE_REG_14__6_ | ~new_P1_U3507 | ~new_P1_U2454;
  assign new_P1_U4459 = ~P1_INSTQUEUE_REG_15__6_ | ~new_P1_U3507 | ~new_P1_U3498;
  assign new_P1_U4460 = ~new_P1_U3277;
  assign new_P1_U4461 = ~P1_INSTQUEUE_REG_7__1_ | ~new_P1_U4382;
  assign new_P1_U4462 = ~P1_INSTQUEUE_REG_0__1_ | ~new_P1_U2472;
  assign new_P1_U4463 = ~P1_INSTQUEUE_REG_1__1_ | ~new_P1_U2471;
  assign new_P1_U4464 = ~P1_INSTQUEUE_REG_2__1_ | ~new_P1_U2470;
  assign new_P1_U4465 = ~P1_INSTQUEUE_REG_3__1_ | ~new_P1_U2468;
  assign new_P1_U4466 = ~P1_INSTQUEUE_REG_4__1_ | ~new_P1_U2467;
  assign new_P1_U4467 = ~P1_INSTQUEUE_REG_5__1_ | ~new_P1_U2466;
  assign new_P1_U4468 = ~P1_INSTQUEUE_REG_6__1_ | ~new_P1_U2465;
  assign new_P1_U4469 = ~P1_INSTQUEUE_REG_8__1_ | ~new_P1_U2464;
  assign new_P1_U4470 = ~P1_INSTQUEUE_REG_9__1_ | ~new_P1_U2463;
  assign new_P1_U4471 = ~P1_INSTQUEUE_REG_10__1_ | ~new_P1_U2461;
  assign new_P1_U4472 = ~P1_INSTQUEUE_REG_11__1_ | ~new_P1_U2459;
  assign new_P1_U4473 = ~P1_INSTQUEUE_REG_12__1_ | ~new_P1_U2458;
  assign new_P1_U4474 = ~P1_INSTQUEUE_REG_13__1_ | ~new_P1_U2457;
  assign new_P1_U4475 = ~P1_INSTQUEUE_REG_14__1_ | ~new_P1_U2455;
  assign new_P1_U4476 = ~P1_INSTQUEUE_REG_15__1_ | ~new_P1_U2453;
  assign new_P1_U4477 = ~new_P1_U3271;
  assign new_P1_U4478 = ~P1_INSTQUEUE_REG_7__0_ | ~new_P1_U4382;
  assign new_P1_U4479 = ~P1_INSTQUEUE_REG_0__0_ | ~new_P1_U2472;
  assign new_P1_U4480 = ~P1_INSTQUEUE_REG_1__0_ | ~new_P1_U2471;
  assign new_P1_U4481 = ~P1_INSTQUEUE_REG_2__0_ | ~new_P1_U2470;
  assign new_P1_U4482 = ~P1_INSTQUEUE_REG_3__0_ | ~new_P1_U2468;
  assign new_P1_U4483 = ~P1_INSTQUEUE_REG_4__0_ | ~new_P1_U2467;
  assign new_P1_U4484 = ~P1_INSTQUEUE_REG_5__0_ | ~new_P1_U2466;
  assign new_P1_U4485 = ~P1_INSTQUEUE_REG_6__0_ | ~new_P1_U2465;
  assign new_P1_U4486 = ~P1_INSTQUEUE_REG_8__0_ | ~new_P1_U2464;
  assign new_P1_U4487 = ~P1_INSTQUEUE_REG_9__0_ | ~new_P1_U2463;
  assign new_P1_U4488 = ~P1_INSTQUEUE_REG_10__0_ | ~new_P1_U2461;
  assign new_P1_U4489 = ~P1_INSTQUEUE_REG_11__0_ | ~new_P1_U2459;
  assign new_P1_U4490 = ~P1_INSTQUEUE_REG_12__0_ | ~new_P1_U2458;
  assign new_P1_U4491 = ~P1_INSTQUEUE_REG_13__0_ | ~new_P1_U2457;
  assign new_P1_U4492 = ~P1_INSTQUEUE_REG_14__0_ | ~new_P1_U2455;
  assign new_P1_U4493 = ~P1_INSTQUEUE_REG_15__0_ | ~new_P1_U2453;
  assign new_P1_U4494 = ~new_P1_U3284;
  assign new_P1_U4495 = ~P1_STATE_REG_2_ | ~new_P1_U3248;
  assign new_P1_U4496 = ~new_P1_U3254 | ~new_P1_U4495;
  assign new_P1_U4497 = ~new_P1_U3272;
  assign new_P1_U4498 = ~new_P1_U4477 | ~new_P1_U3388;
  assign new_P1_U4499 = ~new_P1_U3437;
  assign new_P1_U4500 = ~new_P1_U3287 | ~new_P1_U3272 | ~new_P1_U3390;
  assign new_P1_U4501 = ~new_P1_U4500 | ~new_P1_U3257;
  assign new_P1_U4502 = ~new_P1_U3285;
  assign new_P1_U4503 = ~new_P1_U4460 | ~new_P1_U4173;
  assign new_P1_U4504 = ~new_P1_U4196 | ~new_P1_U3286;
  assign new_P1_U4505 = ~new_P1_U4504 | ~new_P1_U3579;
  assign new_P1_U4506 = ~new_P1_U3580 | ~new_P1_U4505;
  assign new_P1_U4507 = ~new_P1_U4215 | ~new_P1_U3388;
  assign new_P1_U4508 = ~new_P1_U4507 | ~new_P1_U7682 | ~new_P1_U7681;
  assign new_P1_U4509 = ~new_P1_U2448 | ~new_P1_U4262;
  assign new_P1_U4510 = P1_MORE_REG | P1_FLUSH_REG;
  assign new_P1_U4511 = ~new_P1_U3293;
  assign new_P1_U4512 = ~new_P1_U4511 | ~new_P1_U3262;
  assign new_P1_U4513 = ~P1_STATE2_REG_1_ | ~new_U210;
  assign new_P1_U4514 = ~new_P1_U3295;
  assign new_P1_U4515 = ~P1_STATE2_REG_1_ | ~new_P1_U7688 | ~new_P1_U7687;
  assign new_P1_U4516 = ~P1_STATE2_REG_2_ | ~new_P1_U3295;
  assign new_P1_U4517 = ~new_P1_U7604 | ~new_P1_U4246;
  assign new_P1_U4518 = ~new_P1_U3583 | ~new_P1_U4514;
  assign new_P1_U4519 = ~P1_STATE2_REG_1_ | ~new_P1_U4517;
  assign new_P1_U4520 = ~new_P1_U2368 | ~new_P1_U7604;
  assign new_P1_U4521 = ~new_P1_U4252 | ~new_P1_U4261;
  assign new_P1_U4522 = ~new_P1_U7604 | ~new_P1_U4245;
  assign new_P1_U4523 = ~new_P1_U2368 | ~new_P1_U3293;
  assign new_P1_U4524 = ~new_P1_U3325;
  assign new_P1_U4525 = ~new_P1_U3331;
  assign new_P1_U4526 = ~new_P1_U3332;
  assign new_P1_U4527 = ~new_P1_U3314;
  assign new_P1_U4528 = ~new_P1_U3313;
  assign new_P1_U4529 = ~new_P1_U3342;
  assign new_P1_U4530 = ~new_P1_R2144_U8 | ~new_P1_U3313;
  assign new_P1_U4531 = ~new_P1_U3358;
  assign new_P1_U4532 = ~new_P1_U3315;
  assign new_P1_U4533 = ~new_P1_U3305;
  assign new_P1_U4534 = ~new_P1_U3306;
  assign new_P1_U4535 = ~new_P1_U2438 | ~new_P1_U2442;
  assign new_P1_U4536 = ~new_P1_U3321;
  assign new_P1_U4537 = ~new_P1_U3356;
  assign new_P1_U4538 = ~new_P1_U3340;
  assign new_P1_U4539 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_U3305;
  assign new_P1_U4540 = ~new_P1_U3360;
  assign new_P1_U4541 = ~new_P1_U3329;
  assign new_P1_U4542 = ~new_P1_U3323;
  assign new_P1_U4543 = ~new_P1_U3235;
  assign new_P1_U4544 = ~new_P1_U2432 | ~new_P1_U2436;
  assign new_P1_U4545 = ~new_P1_U3322;
  assign new_P1_U4546 = ~P1_STATE2_REG_1_ | ~new_P1_U3263;
  assign new_P1_U4547 = ~new_P1_U3299 | ~new_P1_U4546 | ~new_P1_U3297;
  assign new_P1_U4548 = ~new_P1_U4528 | ~new_P1_U2476;
  assign new_P1_U4549 = ~new_P1_U2480 | ~new_P1_U2358;
  assign new_P1_U4550 = ~new_P1_U3320 | ~new_P1_U4549;
  assign new_P1_U4551 = ~new_P1_U4536 | ~new_P1_U4550;
  assign new_P1_U4552 = ~P1_STATE2_REG_3_ | ~new_P1_U3306;
  assign new_P1_U4553 = ~new_P1_U4545 | ~P1_STATE2_REG_2_;
  assign new_P1_U4554 = ~new_P1_U4551 | ~new_P1_U3587;
  assign new_P1_U4555 = ~new_P1_U2480 | ~new_P1_U2388;
  assign new_P1_U4556 = ~new_P1_U3320 | ~new_P1_U4555;
  assign new_P1_U4557 = ~new_P1_U4556 | ~new_P1_U3321;
  assign new_P1_U4558 = ~P1_STATE2_REG_2_ | ~new_P1_U3322;
  assign new_P1_U4559 = ~new_P1_U4558 | ~new_P1_U4557;
  assign new_P1_U4560 = ~new_P1_U2415 | ~new_P1_U4534;
  assign new_P1_U4561 = ~new_P1_U2413 | ~new_P1_U2477;
  assign new_P1_U4562 = ~new_P1_U2412 | ~new_P1_U4532;
  assign new_P1_U4563 = ~new_P1_U2397 | ~new_P1_U4559;
  assign new_P1_U4564 = ~P1_INSTQUEUE_REG_15__7_ | ~new_P1_U4554;
  assign new_P1_U4565 = ~new_P1_U2416 | ~new_P1_U4534;
  assign new_P1_U4566 = ~new_P1_U2411 | ~new_P1_U2477;
  assign new_P1_U4567 = ~new_P1_U2410 | ~new_P1_U4532;
  assign new_P1_U4568 = ~new_P1_U2396 | ~new_P1_U4559;
  assign new_P1_U4569 = ~P1_INSTQUEUE_REG_15__6_ | ~new_P1_U4554;
  assign new_P1_U4570 = ~new_P1_U2420 | ~new_P1_U4534;
  assign new_P1_U4571 = ~new_P1_U2409 | ~new_P1_U2477;
  assign new_P1_U4572 = ~new_P1_U2408 | ~new_P1_U4532;
  assign new_P1_U4573 = ~new_P1_U2395 | ~new_P1_U4559;
  assign new_P1_U4574 = ~P1_INSTQUEUE_REG_15__5_ | ~new_P1_U4554;
  assign new_P1_U4575 = ~new_P1_U2419 | ~new_P1_U4534;
  assign new_P1_U4576 = ~new_P1_U2407 | ~new_P1_U2477;
  assign new_P1_U4577 = ~new_P1_U2406 | ~new_P1_U4532;
  assign new_P1_U4578 = ~new_P1_U2394 | ~new_P1_U4559;
  assign new_P1_U4579 = ~P1_INSTQUEUE_REG_15__4_ | ~new_P1_U4554;
  assign new_P1_U4580 = ~new_P1_U2418 | ~new_P1_U4534;
  assign new_P1_U4581 = ~new_P1_U2405 | ~new_P1_U2477;
  assign new_P1_U4582 = ~new_P1_U2404 | ~new_P1_U4532;
  assign new_P1_U4583 = ~new_P1_U2393 | ~new_P1_U4559;
  assign new_P1_U4584 = ~P1_INSTQUEUE_REG_15__3_ | ~new_P1_U4554;
  assign new_P1_U4585 = ~new_P1_U2421 | ~new_P1_U4534;
  assign new_P1_U4586 = ~new_P1_U2403 | ~new_P1_U2477;
  assign new_P1_U4587 = ~new_P1_U2402 | ~new_P1_U4532;
  assign new_P1_U4588 = ~new_P1_U2392 | ~new_P1_U4559;
  assign new_P1_U4589 = ~P1_INSTQUEUE_REG_15__2_ | ~new_P1_U4554;
  assign new_P1_U4590 = ~new_P1_U2414 | ~new_P1_U4534;
  assign new_P1_U4591 = ~new_P1_U2401 | ~new_P1_U2477;
  assign new_P1_U4592 = ~new_P1_U2400 | ~new_P1_U4532;
  assign new_P1_U4593 = ~new_P1_U2391 | ~new_P1_U4559;
  assign new_P1_U4594 = ~P1_INSTQUEUE_REG_15__1_ | ~new_P1_U4554;
  assign new_P1_U4595 = ~new_P1_U2417 | ~new_P1_U4534;
  assign new_P1_U4596 = ~new_P1_U2399 | ~new_P1_U2477;
  assign new_P1_U4597 = ~new_P1_U2398 | ~new_P1_U4532;
  assign new_P1_U4598 = ~new_P1_U2390 | ~new_P1_U4559;
  assign new_P1_U4599 = ~P1_INSTQUEUE_REG_15__0_ | ~new_P1_U4554;
  assign new_P1_U4600 = ~new_P1_U3326;
  assign new_P1_U4601 = ~new_P1_U3327;
  assign new_P1_U4602 = ~new_P1_U3324;
  assign new_P1_U4603 = ~new_P1_U2443 | ~new_P1_U2438;
  assign new_P1_U4604 = ~new_P1_U3328;
  assign new_P1_U4605 = ~new_P1_U3236;
  assign new_P1_U4606 = ~new_P1_U4524 | ~new_P1_U2476;
  assign new_P1_U4607 = ~new_P1_U2482 | ~new_P1_U2358;
  assign new_P1_U4608 = ~new_P1_U3320 | ~new_P1_U4607;
  assign new_P1_U4609 = ~new_P1_U4604 | ~new_P1_U4608;
  assign new_P1_U4610 = ~P1_STATE2_REG_3_ | ~new_P1_U3324;
  assign new_P1_U4611 = ~P1_STATE2_REG_2_ | ~new_P1_U3236;
  assign new_P1_U4612 = ~new_P1_U4609 | ~new_P1_U3596;
  assign new_P1_U4613 = ~new_P1_U2482 | ~new_P1_U2388;
  assign new_P1_U4614 = ~new_P1_U3320 | ~new_P1_U4613;
  assign new_P1_U4615 = ~new_P1_U4614 | ~new_P1_U3328;
  assign new_P1_U4616 = ~P1_STATE2_REG_2_ | ~new_P1_U4605;
  assign new_P1_U4617 = ~new_P1_U4616 | ~new_P1_U4615;
  assign new_P1_U4618 = ~new_P1_U4602 | ~new_P1_U2415;
  assign new_P1_U4619 = ~new_P1_U2481 | ~new_P1_U2413;
  assign new_P1_U4620 = ~new_P1_U4601 | ~new_P1_U2412;
  assign new_P1_U4621 = ~new_P1_U2397 | ~new_P1_U4617;
  assign new_P1_U4622 = ~P1_INSTQUEUE_REG_14__7_ | ~new_P1_U4612;
  assign new_P1_U4623 = ~new_P1_U4602 | ~new_P1_U2416;
  assign new_P1_U4624 = ~new_P1_U2481 | ~new_P1_U2411;
  assign new_P1_U4625 = ~new_P1_U4601 | ~new_P1_U2410;
  assign new_P1_U4626 = ~new_P1_U2396 | ~new_P1_U4617;
  assign new_P1_U4627 = ~P1_INSTQUEUE_REG_14__6_ | ~new_P1_U4612;
  assign new_P1_U4628 = ~new_P1_U4602 | ~new_P1_U2420;
  assign new_P1_U4629 = ~new_P1_U2481 | ~new_P1_U2409;
  assign new_P1_U4630 = ~new_P1_U4601 | ~new_P1_U2408;
  assign new_P1_U4631 = ~new_P1_U2395 | ~new_P1_U4617;
  assign new_P1_U4632 = ~P1_INSTQUEUE_REG_14__5_ | ~new_P1_U4612;
  assign new_P1_U4633 = ~new_P1_U4602 | ~new_P1_U2419;
  assign new_P1_U4634 = ~new_P1_U2481 | ~new_P1_U2407;
  assign new_P1_U4635 = ~new_P1_U4601 | ~new_P1_U2406;
  assign new_P1_U4636 = ~new_P1_U2394 | ~new_P1_U4617;
  assign new_P1_U4637 = ~P1_INSTQUEUE_REG_14__4_ | ~new_P1_U4612;
  assign new_P1_U4638 = ~new_P1_U4602 | ~new_P1_U2418;
  assign new_P1_U4639 = ~new_P1_U2481 | ~new_P1_U2405;
  assign new_P1_U4640 = ~new_P1_U4601 | ~new_P1_U2404;
  assign new_P1_U4641 = ~new_P1_U2393 | ~new_P1_U4617;
  assign new_P1_U4642 = ~P1_INSTQUEUE_REG_14__3_ | ~new_P1_U4612;
  assign new_P1_U4643 = ~new_P1_U4602 | ~new_P1_U2421;
  assign new_P1_U4644 = ~new_P1_U2481 | ~new_P1_U2403;
  assign new_P1_U4645 = ~new_P1_U4601 | ~new_P1_U2402;
  assign new_P1_U4646 = ~new_P1_U2392 | ~new_P1_U4617;
  assign new_P1_U4647 = ~P1_INSTQUEUE_REG_14__2_ | ~new_P1_U4612;
  assign new_P1_U4648 = ~new_P1_U4602 | ~new_P1_U2414;
  assign new_P1_U4649 = ~new_P1_U2481 | ~new_P1_U2401;
  assign new_P1_U4650 = ~new_P1_U4601 | ~new_P1_U2400;
  assign new_P1_U4651 = ~new_P1_U2391 | ~new_P1_U4617;
  assign new_P1_U4652 = ~P1_INSTQUEUE_REG_14__1_ | ~new_P1_U4612;
  assign new_P1_U4653 = ~new_P1_U4602 | ~new_P1_U2417;
  assign new_P1_U4654 = ~new_P1_U2481 | ~new_P1_U2399;
  assign new_P1_U4655 = ~new_P1_U4601 | ~new_P1_U2398;
  assign new_P1_U4656 = ~new_P1_U2390 | ~new_P1_U4617;
  assign new_P1_U4657 = ~P1_INSTQUEUE_REG_14__0_ | ~new_P1_U4612;
  assign new_P1_U4658 = ~new_P1_U3333;
  assign new_P1_U4659 = ~new_P1_U3334;
  assign new_P1_U4660 = ~new_P1_U3330;
  assign new_P1_U4661 = ~new_P1_U2444 | ~new_P1_U2438;
  assign new_P1_U4662 = ~new_P1_U3335;
  assign new_P1_U4663 = ~new_P1_U2437 | ~new_P1_U2432;
  assign new_P1_U4664 = ~new_P1_U3336;
  assign new_P1_U4665 = ~new_P1_U4525 | ~new_P1_U2476;
  assign new_P1_U4666 = ~new_P1_U2484 | ~new_P1_U2358;
  assign new_P1_U4667 = ~new_P1_U3320 | ~new_P1_U4666;
  assign new_P1_U4668 = ~new_P1_U4662 | ~new_P1_U4667;
  assign new_P1_U4669 = ~P1_STATE2_REG_3_ | ~new_P1_U3330;
  assign new_P1_U4670 = ~new_P1_U4664 | ~P1_STATE2_REG_2_;
  assign new_P1_U4671 = ~new_P1_U4668 | ~new_P1_U3605;
  assign new_P1_U4672 = ~new_P1_U2484 | ~new_P1_U2388;
  assign new_P1_U4673 = ~new_P1_U3320 | ~new_P1_U4672;
  assign new_P1_U4674 = ~new_P1_U4673 | ~new_P1_U3335;
  assign new_P1_U4675 = ~P1_STATE2_REG_2_ | ~new_P1_U3336;
  assign new_P1_U4676 = ~new_P1_U4675 | ~new_P1_U4674;
  assign new_P1_U4677 = ~new_P1_U4660 | ~new_P1_U2415;
  assign new_P1_U4678 = ~new_P1_U2483 | ~new_P1_U2413;
  assign new_P1_U4679 = ~new_P1_U4659 | ~new_P1_U2412;
  assign new_P1_U4680 = ~new_P1_U2397 | ~new_P1_U4676;
  assign new_P1_U4681 = ~P1_INSTQUEUE_REG_13__7_ | ~new_P1_U4671;
  assign new_P1_U4682 = ~new_P1_U4660 | ~new_P1_U2416;
  assign new_P1_U4683 = ~new_P1_U2483 | ~new_P1_U2411;
  assign new_P1_U4684 = ~new_P1_U4659 | ~new_P1_U2410;
  assign new_P1_U4685 = ~new_P1_U2396 | ~new_P1_U4676;
  assign new_P1_U4686 = ~P1_INSTQUEUE_REG_13__6_ | ~new_P1_U4671;
  assign new_P1_U4687 = ~new_P1_U4660 | ~new_P1_U2420;
  assign new_P1_U4688 = ~new_P1_U2483 | ~new_P1_U2409;
  assign new_P1_U4689 = ~new_P1_U4659 | ~new_P1_U2408;
  assign new_P1_U4690 = ~new_P1_U2395 | ~new_P1_U4676;
  assign new_P1_U4691 = ~P1_INSTQUEUE_REG_13__5_ | ~new_P1_U4671;
  assign new_P1_U4692 = ~new_P1_U4660 | ~new_P1_U2419;
  assign new_P1_U4693 = ~new_P1_U2483 | ~new_P1_U2407;
  assign new_P1_U4694 = ~new_P1_U4659 | ~new_P1_U2406;
  assign new_P1_U4695 = ~new_P1_U2394 | ~new_P1_U4676;
  assign new_P1_U4696 = ~P1_INSTQUEUE_REG_13__4_ | ~new_P1_U4671;
  assign new_P1_U4697 = ~new_P1_U4660 | ~new_P1_U2418;
  assign new_P1_U4698 = ~new_P1_U2483 | ~new_P1_U2405;
  assign new_P1_U4699 = ~new_P1_U4659 | ~new_P1_U2404;
  assign new_P1_U4700 = ~new_P1_U2393 | ~new_P1_U4676;
  assign new_P1_U4701 = ~P1_INSTQUEUE_REG_13__3_ | ~new_P1_U4671;
  assign new_P1_U4702 = ~new_P1_U4660 | ~new_P1_U2421;
  assign new_P1_U4703 = ~new_P1_U2483 | ~new_P1_U2403;
  assign new_P1_U4704 = ~new_P1_U4659 | ~new_P1_U2402;
  assign new_P1_U4705 = ~new_P1_U2392 | ~new_P1_U4676;
  assign new_P1_U4706 = ~P1_INSTQUEUE_REG_13__2_ | ~new_P1_U4671;
  assign new_P1_U4707 = ~new_P1_U4660 | ~new_P1_U2414;
  assign new_P1_U4708 = ~new_P1_U2483 | ~new_P1_U2401;
  assign new_P1_U4709 = ~new_P1_U4659 | ~new_P1_U2400;
  assign new_P1_U4710 = ~new_P1_U2391 | ~new_P1_U4676;
  assign new_P1_U4711 = ~P1_INSTQUEUE_REG_13__1_ | ~new_P1_U4671;
  assign new_P1_U4712 = ~new_P1_U4660 | ~new_P1_U2417;
  assign new_P1_U4713 = ~new_P1_U2483 | ~new_P1_U2399;
  assign new_P1_U4714 = ~new_P1_U4659 | ~new_P1_U2398;
  assign new_P1_U4715 = ~new_P1_U2390 | ~new_P1_U4676;
  assign new_P1_U4716 = ~P1_INSTQUEUE_REG_13__0_ | ~new_P1_U4671;
  assign new_P1_U4717 = ~new_P1_U3338;
  assign new_P1_U4718 = ~new_P1_U3337;
  assign new_P1_U4719 = ~new_P1_U2445 | ~new_P1_U2438;
  assign new_P1_U4720 = ~new_P1_U3339;
  assign new_P1_U4721 = ~new_P1_U3237;
  assign new_P1_U4722 = ~new_P1_U2486 | ~new_P1_U2476;
  assign new_P1_U4723 = ~new_P1_U2489 | ~new_P1_U2358;
  assign new_P1_U4724 = ~new_P1_U3320 | ~new_P1_U4723;
  assign new_P1_U4725 = ~new_P1_U4720 | ~new_P1_U4724;
  assign new_P1_U4726 = ~P1_STATE2_REG_3_ | ~new_P1_U3337;
  assign new_P1_U4727 = ~P1_STATE2_REG_2_ | ~new_P1_U3237;
  assign new_P1_U4728 = ~new_P1_U4725 | ~new_P1_U3614;
  assign new_P1_U4729 = ~new_P1_U2489 | ~new_P1_U2388;
  assign new_P1_U4730 = ~new_P1_U3320 | ~new_P1_U4729;
  assign new_P1_U4731 = ~new_P1_U4730 | ~new_P1_U3339;
  assign new_P1_U4732 = ~P1_STATE2_REG_2_ | ~new_P1_U4721;
  assign new_P1_U4733 = ~new_P1_U4732 | ~new_P1_U4731;
  assign new_P1_U4734 = ~new_P1_U4718 | ~new_P1_U2415;
  assign new_P1_U4735 = ~new_P1_U2487 | ~new_P1_U2413;
  assign new_P1_U4736 = ~new_P1_U4717 | ~new_P1_U2412;
  assign new_P1_U4737 = ~new_P1_U2397 | ~new_P1_U4733;
  assign new_P1_U4738 = ~P1_INSTQUEUE_REG_12__7_ | ~new_P1_U4728;
  assign new_P1_U4739 = ~new_P1_U4718 | ~new_P1_U2416;
  assign new_P1_U4740 = ~new_P1_U2487 | ~new_P1_U2411;
  assign new_P1_U4741 = ~new_P1_U4717 | ~new_P1_U2410;
  assign new_P1_U4742 = ~new_P1_U2396 | ~new_P1_U4733;
  assign new_P1_U4743 = ~P1_INSTQUEUE_REG_12__6_ | ~new_P1_U4728;
  assign new_P1_U4744 = ~new_P1_U4718 | ~new_P1_U2420;
  assign new_P1_U4745 = ~new_P1_U2487 | ~new_P1_U2409;
  assign new_P1_U4746 = ~new_P1_U4717 | ~new_P1_U2408;
  assign new_P1_U4747 = ~new_P1_U2395 | ~new_P1_U4733;
  assign new_P1_U4748 = ~P1_INSTQUEUE_REG_12__5_ | ~new_P1_U4728;
  assign new_P1_U4749 = ~new_P1_U4718 | ~new_P1_U2419;
  assign new_P1_U4750 = ~new_P1_U2487 | ~new_P1_U2407;
  assign new_P1_U4751 = ~new_P1_U4717 | ~new_P1_U2406;
  assign new_P1_U4752 = ~new_P1_U2394 | ~new_P1_U4733;
  assign new_P1_U4753 = ~P1_INSTQUEUE_REG_12__4_ | ~new_P1_U4728;
  assign new_P1_U4754 = ~new_P1_U4718 | ~new_P1_U2418;
  assign new_P1_U4755 = ~new_P1_U2487 | ~new_P1_U2405;
  assign new_P1_U4756 = ~new_P1_U4717 | ~new_P1_U2404;
  assign new_P1_U4757 = ~new_P1_U2393 | ~new_P1_U4733;
  assign new_P1_U4758 = ~P1_INSTQUEUE_REG_12__3_ | ~new_P1_U4728;
  assign new_P1_U4759 = ~new_P1_U4718 | ~new_P1_U2421;
  assign new_P1_U4760 = ~new_P1_U2487 | ~new_P1_U2403;
  assign new_P1_U4761 = ~new_P1_U4717 | ~new_P1_U2402;
  assign new_P1_U4762 = ~new_P1_U2392 | ~new_P1_U4733;
  assign new_P1_U4763 = ~P1_INSTQUEUE_REG_12__2_ | ~new_P1_U4728;
  assign new_P1_U4764 = ~new_P1_U4718 | ~new_P1_U2414;
  assign new_P1_U4765 = ~new_P1_U2487 | ~new_P1_U2401;
  assign new_P1_U4766 = ~new_P1_U4717 | ~new_P1_U2400;
  assign new_P1_U4767 = ~new_P1_U2391 | ~new_P1_U4733;
  assign new_P1_U4768 = ~P1_INSTQUEUE_REG_12__1_ | ~new_P1_U4728;
  assign new_P1_U4769 = ~new_P1_U4718 | ~new_P1_U2417;
  assign new_P1_U4770 = ~new_P1_U2487 | ~new_P1_U2399;
  assign new_P1_U4771 = ~new_P1_U4717 | ~new_P1_U2398;
  assign new_P1_U4772 = ~new_P1_U2390 | ~new_P1_U4733;
  assign new_P1_U4773 = ~P1_INSTQUEUE_REG_12__0_ | ~new_P1_U4728;
  assign new_P1_U4774 = ~new_P1_U3343;
  assign new_P1_U4775 = ~new_P1_U3341;
  assign new_P1_U4776 = ~new_P1_U2440 | ~new_P1_U2442;
  assign new_P1_U4777 = ~new_P1_U3344;
  assign new_P1_U4778 = ~new_P1_U2434 | ~new_P1_U2436;
  assign new_P1_U4779 = ~new_P1_U3345;
  assign new_P1_U4780 = ~new_P1_U4529 | ~new_P1_U4528;
  assign new_P1_U4781 = ~new_P1_U2492 | ~new_P1_U2358;
  assign new_P1_U4782 = ~new_P1_U3320 | ~new_P1_U4781;
  assign new_P1_U4783 = ~new_P1_U4777 | ~new_P1_U4782;
  assign new_P1_U4784 = ~P1_STATE2_REG_3_ | ~new_P1_U3341;
  assign new_P1_U4785 = ~new_P1_U4779 | ~P1_STATE2_REG_2_;
  assign new_P1_U4786 = ~new_P1_U4783 | ~new_P1_U3623;
  assign new_P1_U4787 = ~new_P1_U2492 | ~new_P1_U2388;
  assign new_P1_U4788 = ~new_P1_U3320 | ~new_P1_U4787;
  assign new_P1_U4789 = ~new_P1_U4788 | ~new_P1_U3344;
  assign new_P1_U4790 = ~P1_STATE2_REG_2_ | ~new_P1_U3345;
  assign new_P1_U4791 = ~new_P1_U4790 | ~new_P1_U4789;
  assign new_P1_U4792 = ~new_P1_U4775 | ~new_P1_U2415;
  assign new_P1_U4793 = ~new_P1_U2491 | ~new_P1_U2413;
  assign new_P1_U4794 = ~new_P1_U4774 | ~new_P1_U2412;
  assign new_P1_U4795 = ~new_P1_U2397 | ~new_P1_U4791;
  assign new_P1_U4796 = ~P1_INSTQUEUE_REG_11__7_ | ~new_P1_U4786;
  assign new_P1_U4797 = ~new_P1_U4775 | ~new_P1_U2416;
  assign new_P1_U4798 = ~new_P1_U2491 | ~new_P1_U2411;
  assign new_P1_U4799 = ~new_P1_U4774 | ~new_P1_U2410;
  assign new_P1_U4800 = ~new_P1_U2396 | ~new_P1_U4791;
  assign new_P1_U4801 = ~P1_INSTQUEUE_REG_11__6_ | ~new_P1_U4786;
  assign new_P1_U4802 = ~new_P1_U4775 | ~new_P1_U2420;
  assign new_P1_U4803 = ~new_P1_U2491 | ~new_P1_U2409;
  assign new_P1_U4804 = ~new_P1_U4774 | ~new_P1_U2408;
  assign new_P1_U4805 = ~new_P1_U2395 | ~new_P1_U4791;
  assign new_P1_U4806 = ~P1_INSTQUEUE_REG_11__5_ | ~new_P1_U4786;
  assign new_P1_U4807 = ~new_P1_U4775 | ~new_P1_U2419;
  assign new_P1_U4808 = ~new_P1_U2491 | ~new_P1_U2407;
  assign new_P1_U4809 = ~new_P1_U4774 | ~new_P1_U2406;
  assign new_P1_U4810 = ~new_P1_U2394 | ~new_P1_U4791;
  assign new_P1_U4811 = ~P1_INSTQUEUE_REG_11__4_ | ~new_P1_U4786;
  assign new_P1_U4812 = ~new_P1_U4775 | ~new_P1_U2418;
  assign new_P1_U4813 = ~new_P1_U2491 | ~new_P1_U2405;
  assign new_P1_U4814 = ~new_P1_U4774 | ~new_P1_U2404;
  assign new_P1_U4815 = ~new_P1_U2393 | ~new_P1_U4791;
  assign new_P1_U4816 = ~P1_INSTQUEUE_REG_11__3_ | ~new_P1_U4786;
  assign new_P1_U4817 = ~new_P1_U4775 | ~new_P1_U2421;
  assign new_P1_U4818 = ~new_P1_U2491 | ~new_P1_U2403;
  assign new_P1_U4819 = ~new_P1_U4774 | ~new_P1_U2402;
  assign new_P1_U4820 = ~new_P1_U2392 | ~new_P1_U4791;
  assign new_P1_U4821 = ~P1_INSTQUEUE_REG_11__2_ | ~new_P1_U4786;
  assign new_P1_U4822 = ~new_P1_U4775 | ~new_P1_U2414;
  assign new_P1_U4823 = ~new_P1_U2491 | ~new_P1_U2401;
  assign new_P1_U4824 = ~new_P1_U4774 | ~new_P1_U2400;
  assign new_P1_U4825 = ~new_P1_U2391 | ~new_P1_U4791;
  assign new_P1_U4826 = ~P1_INSTQUEUE_REG_11__1_ | ~new_P1_U4786;
  assign new_P1_U4827 = ~new_P1_U4775 | ~new_P1_U2417;
  assign new_P1_U4828 = ~new_P1_U2491 | ~new_P1_U2399;
  assign new_P1_U4829 = ~new_P1_U4774 | ~new_P1_U2398;
  assign new_P1_U4830 = ~new_P1_U2390 | ~new_P1_U4791;
  assign new_P1_U4831 = ~P1_INSTQUEUE_REG_11__0_ | ~new_P1_U4786;
  assign new_P1_U4832 = ~new_P1_U3347;
  assign new_P1_U4833 = ~new_P1_U3346;
  assign new_P1_U4834 = ~new_P1_U2440 | ~new_P1_U2443;
  assign new_P1_U4835 = ~new_P1_U3348;
  assign new_P1_U4836 = ~new_P1_U3238;
  assign new_P1_U4837 = ~new_P1_U4529 | ~new_P1_U4524;
  assign new_P1_U4838 = ~new_P1_U2494 | ~new_P1_U2358;
  assign new_P1_U4839 = ~new_P1_U3320 | ~new_P1_U4838;
  assign new_P1_U4840 = ~new_P1_U4835 | ~new_P1_U4839;
  assign new_P1_U4841 = ~P1_STATE2_REG_3_ | ~new_P1_U3346;
  assign new_P1_U4842 = ~P1_STATE2_REG_2_ | ~new_P1_U3238;
  assign new_P1_U4843 = ~new_P1_U4840 | ~new_P1_U3632;
  assign new_P1_U4844 = ~new_P1_U2494 | ~new_P1_U2388;
  assign new_P1_U4845 = ~new_P1_U3320 | ~new_P1_U4844;
  assign new_P1_U4846 = ~new_P1_U4845 | ~new_P1_U3348;
  assign new_P1_U4847 = ~P1_STATE2_REG_2_ | ~new_P1_U4836;
  assign new_P1_U4848 = ~new_P1_U4847 | ~new_P1_U4846;
  assign new_P1_U4849 = ~new_P1_U4833 | ~new_P1_U2415;
  assign new_P1_U4850 = ~new_P1_U2493 | ~new_P1_U2413;
  assign new_P1_U4851 = ~new_P1_U4832 | ~new_P1_U2412;
  assign new_P1_U4852 = ~new_P1_U2397 | ~new_P1_U4848;
  assign new_P1_U4853 = ~P1_INSTQUEUE_REG_10__7_ | ~new_P1_U4843;
  assign new_P1_U4854 = ~new_P1_U4833 | ~new_P1_U2416;
  assign new_P1_U4855 = ~new_P1_U2493 | ~new_P1_U2411;
  assign new_P1_U4856 = ~new_P1_U4832 | ~new_P1_U2410;
  assign new_P1_U4857 = ~new_P1_U2396 | ~new_P1_U4848;
  assign new_P1_U4858 = ~P1_INSTQUEUE_REG_10__6_ | ~new_P1_U4843;
  assign new_P1_U4859 = ~new_P1_U4833 | ~new_P1_U2420;
  assign new_P1_U4860 = ~new_P1_U2493 | ~new_P1_U2409;
  assign new_P1_U4861 = ~new_P1_U4832 | ~new_P1_U2408;
  assign new_P1_U4862 = ~new_P1_U2395 | ~new_P1_U4848;
  assign new_P1_U4863 = ~P1_INSTQUEUE_REG_10__5_ | ~new_P1_U4843;
  assign new_P1_U4864 = ~new_P1_U4833 | ~new_P1_U2419;
  assign new_P1_U4865 = ~new_P1_U2493 | ~new_P1_U2407;
  assign new_P1_U4866 = ~new_P1_U4832 | ~new_P1_U2406;
  assign new_P1_U4867 = ~new_P1_U2394 | ~new_P1_U4848;
  assign new_P1_U4868 = ~P1_INSTQUEUE_REG_10__4_ | ~new_P1_U4843;
  assign new_P1_U4869 = ~new_P1_U4833 | ~new_P1_U2418;
  assign new_P1_U4870 = ~new_P1_U2493 | ~new_P1_U2405;
  assign new_P1_U4871 = ~new_P1_U4832 | ~new_P1_U2404;
  assign new_P1_U4872 = ~new_P1_U2393 | ~new_P1_U4848;
  assign new_P1_U4873 = ~P1_INSTQUEUE_REG_10__3_ | ~new_P1_U4843;
  assign new_P1_U4874 = ~new_P1_U4833 | ~new_P1_U2421;
  assign new_P1_U4875 = ~new_P1_U2493 | ~new_P1_U2403;
  assign new_P1_U4876 = ~new_P1_U4832 | ~new_P1_U2402;
  assign new_P1_U4877 = ~new_P1_U2392 | ~new_P1_U4848;
  assign new_P1_U4878 = ~P1_INSTQUEUE_REG_10__2_ | ~new_P1_U4843;
  assign new_P1_U4879 = ~new_P1_U4833 | ~new_P1_U2414;
  assign new_P1_U4880 = ~new_P1_U2493 | ~new_P1_U2401;
  assign new_P1_U4881 = ~new_P1_U4832 | ~new_P1_U2400;
  assign new_P1_U4882 = ~new_P1_U2391 | ~new_P1_U4848;
  assign new_P1_U4883 = ~P1_INSTQUEUE_REG_10__1_ | ~new_P1_U4843;
  assign new_P1_U4884 = ~new_P1_U4833 | ~new_P1_U2417;
  assign new_P1_U4885 = ~new_P1_U2493 | ~new_P1_U2399;
  assign new_P1_U4886 = ~new_P1_U4832 | ~new_P1_U2398;
  assign new_P1_U4887 = ~new_P1_U2390 | ~new_P1_U4848;
  assign new_P1_U4888 = ~P1_INSTQUEUE_REG_10__0_ | ~new_P1_U4843;
  assign new_P1_U4889 = ~new_P1_U3350;
  assign new_P1_U4890 = ~new_P1_U3349;
  assign new_P1_U4891 = ~new_P1_U2440 | ~new_P1_U2444;
  assign new_P1_U4892 = ~new_P1_U3351;
  assign new_P1_U4893 = ~new_P1_U2434 | ~new_P1_U2437;
  assign new_P1_U4894 = ~new_P1_U3352;
  assign new_P1_U4895 = ~new_P1_U4529 | ~new_P1_U4525;
  assign new_P1_U4896 = ~new_P1_U2496 | ~new_P1_U2358;
  assign new_P1_U4897 = ~new_P1_U3320 | ~new_P1_U4896;
  assign new_P1_U4898 = ~new_P1_U4892 | ~new_P1_U4897;
  assign new_P1_U4899 = ~P1_STATE2_REG_3_ | ~new_P1_U3349;
  assign new_P1_U4900 = ~new_P1_U4894 | ~P1_STATE2_REG_2_;
  assign new_P1_U4901 = ~new_P1_U4898 | ~new_P1_U3641;
  assign new_P1_U4902 = ~new_P1_U2496 | ~new_P1_U2388;
  assign new_P1_U4903 = ~new_P1_U3320 | ~new_P1_U4902;
  assign new_P1_U4904 = ~new_P1_U4903 | ~new_P1_U3351;
  assign new_P1_U4905 = ~P1_STATE2_REG_2_ | ~new_P1_U3352;
  assign new_P1_U4906 = ~new_P1_U4905 | ~new_P1_U4904;
  assign new_P1_U4907 = ~new_P1_U4890 | ~new_P1_U2415;
  assign new_P1_U4908 = ~new_P1_U2495 | ~new_P1_U2413;
  assign new_P1_U4909 = ~new_P1_U4889 | ~new_P1_U2412;
  assign new_P1_U4910 = ~new_P1_U2397 | ~new_P1_U4906;
  assign new_P1_U4911 = ~P1_INSTQUEUE_REG_9__7_ | ~new_P1_U4901;
  assign new_P1_U4912 = ~new_P1_U4890 | ~new_P1_U2416;
  assign new_P1_U4913 = ~new_P1_U2495 | ~new_P1_U2411;
  assign new_P1_U4914 = ~new_P1_U4889 | ~new_P1_U2410;
  assign new_P1_U4915 = ~new_P1_U2396 | ~new_P1_U4906;
  assign new_P1_U4916 = ~P1_INSTQUEUE_REG_9__6_ | ~new_P1_U4901;
  assign new_P1_U4917 = ~new_P1_U4890 | ~new_P1_U2420;
  assign new_P1_U4918 = ~new_P1_U2495 | ~new_P1_U2409;
  assign new_P1_U4919 = ~new_P1_U4889 | ~new_P1_U2408;
  assign new_P1_U4920 = ~new_P1_U2395 | ~new_P1_U4906;
  assign new_P1_U4921 = ~P1_INSTQUEUE_REG_9__5_ | ~new_P1_U4901;
  assign new_P1_U4922 = ~new_P1_U4890 | ~new_P1_U2419;
  assign new_P1_U4923 = ~new_P1_U2495 | ~new_P1_U2407;
  assign new_P1_U4924 = ~new_P1_U4889 | ~new_P1_U2406;
  assign new_P1_U4925 = ~new_P1_U2394 | ~new_P1_U4906;
  assign new_P1_U4926 = ~P1_INSTQUEUE_REG_9__4_ | ~new_P1_U4901;
  assign new_P1_U4927 = ~new_P1_U4890 | ~new_P1_U2418;
  assign new_P1_U4928 = ~new_P1_U2495 | ~new_P1_U2405;
  assign new_P1_U4929 = ~new_P1_U4889 | ~new_P1_U2404;
  assign new_P1_U4930 = ~new_P1_U2393 | ~new_P1_U4906;
  assign new_P1_U4931 = ~P1_INSTQUEUE_REG_9__3_ | ~new_P1_U4901;
  assign new_P1_U4932 = ~new_P1_U4890 | ~new_P1_U2421;
  assign new_P1_U4933 = ~new_P1_U2495 | ~new_P1_U2403;
  assign new_P1_U4934 = ~new_P1_U4889 | ~new_P1_U2402;
  assign new_P1_U4935 = ~new_P1_U2392 | ~new_P1_U4906;
  assign new_P1_U4936 = ~P1_INSTQUEUE_REG_9__2_ | ~new_P1_U4901;
  assign new_P1_U4937 = ~new_P1_U4890 | ~new_P1_U2414;
  assign new_P1_U4938 = ~new_P1_U2495 | ~new_P1_U2401;
  assign new_P1_U4939 = ~new_P1_U4889 | ~new_P1_U2400;
  assign new_P1_U4940 = ~new_P1_U2391 | ~new_P1_U4906;
  assign new_P1_U4941 = ~P1_INSTQUEUE_REG_9__1_ | ~new_P1_U4901;
  assign new_P1_U4942 = ~new_P1_U4890 | ~new_P1_U2417;
  assign new_P1_U4943 = ~new_P1_U2495 | ~new_P1_U2399;
  assign new_P1_U4944 = ~new_P1_U4889 | ~new_P1_U2398;
  assign new_P1_U4945 = ~new_P1_U2390 | ~new_P1_U4906;
  assign new_P1_U4946 = ~P1_INSTQUEUE_REG_9__0_ | ~new_P1_U4901;
  assign new_P1_U4947 = ~new_P1_U3354;
  assign new_P1_U4948 = ~new_P1_U3353;
  assign new_P1_U4949 = ~new_P1_U2440 | ~new_P1_U2445;
  assign new_P1_U4950 = ~new_P1_U3355;
  assign new_P1_U4951 = ~new_P1_U3239;
  assign new_P1_U4952 = ~new_P1_U4529 | ~new_P1_U2486;
  assign new_P1_U4953 = ~new_P1_U2498 | ~new_P1_U2358;
  assign new_P1_U4954 = ~new_P1_U3320 | ~new_P1_U4953;
  assign new_P1_U4955 = ~new_P1_U4950 | ~new_P1_U4954;
  assign new_P1_U4956 = ~P1_STATE2_REG_3_ | ~new_P1_U3353;
  assign new_P1_U4957 = ~P1_STATE2_REG_2_ | ~new_P1_U3239;
  assign new_P1_U4958 = ~new_P1_U4955 | ~new_P1_U3650;
  assign new_P1_U4959 = ~new_P1_U2498 | ~new_P1_U2388;
  assign new_P1_U4960 = ~new_P1_U3320 | ~new_P1_U4959;
  assign new_P1_U4961 = ~new_P1_U4960 | ~new_P1_U3355;
  assign new_P1_U4962 = ~P1_STATE2_REG_2_ | ~new_P1_U4951;
  assign new_P1_U4963 = ~new_P1_U4962 | ~new_P1_U4961;
  assign new_P1_U4964 = ~new_P1_U4948 | ~new_P1_U2415;
  assign new_P1_U4965 = ~new_P1_U2497 | ~new_P1_U2413;
  assign new_P1_U4966 = ~new_P1_U4947 | ~new_P1_U2412;
  assign new_P1_U4967 = ~new_P1_U2397 | ~new_P1_U4963;
  assign new_P1_U4968 = ~P1_INSTQUEUE_REG_8__7_ | ~new_P1_U4958;
  assign new_P1_U4969 = ~new_P1_U4948 | ~new_P1_U2416;
  assign new_P1_U4970 = ~new_P1_U2497 | ~new_P1_U2411;
  assign new_P1_U4971 = ~new_P1_U4947 | ~new_P1_U2410;
  assign new_P1_U4972 = ~new_P1_U2396 | ~new_P1_U4963;
  assign new_P1_U4973 = ~P1_INSTQUEUE_REG_8__6_ | ~new_P1_U4958;
  assign new_P1_U4974 = ~new_P1_U4948 | ~new_P1_U2420;
  assign new_P1_U4975 = ~new_P1_U2497 | ~new_P1_U2409;
  assign new_P1_U4976 = ~new_P1_U4947 | ~new_P1_U2408;
  assign new_P1_U4977 = ~new_P1_U2395 | ~new_P1_U4963;
  assign new_P1_U4978 = ~P1_INSTQUEUE_REG_8__5_ | ~new_P1_U4958;
  assign new_P1_U4979 = ~new_P1_U4948 | ~new_P1_U2419;
  assign new_P1_U4980 = ~new_P1_U2497 | ~new_P1_U2407;
  assign new_P1_U4981 = ~new_P1_U4947 | ~new_P1_U2406;
  assign new_P1_U4982 = ~new_P1_U2394 | ~new_P1_U4963;
  assign new_P1_U4983 = ~P1_INSTQUEUE_REG_8__4_ | ~new_P1_U4958;
  assign new_P1_U4984 = ~new_P1_U4948 | ~new_P1_U2418;
  assign new_P1_U4985 = ~new_P1_U2497 | ~new_P1_U2405;
  assign new_P1_U4986 = ~new_P1_U4947 | ~new_P1_U2404;
  assign new_P1_U4987 = ~new_P1_U2393 | ~new_P1_U4963;
  assign new_P1_U4988 = ~P1_INSTQUEUE_REG_8__3_ | ~new_P1_U4958;
  assign new_P1_U4989 = ~new_P1_U4948 | ~new_P1_U2421;
  assign new_P1_U4990 = ~new_P1_U2497 | ~new_P1_U2403;
  assign new_P1_U4991 = ~new_P1_U4947 | ~new_P1_U2402;
  assign new_P1_U4992 = ~new_P1_U2392 | ~new_P1_U4963;
  assign new_P1_U4993 = ~P1_INSTQUEUE_REG_8__2_ | ~new_P1_U4958;
  assign new_P1_U4994 = ~new_P1_U4948 | ~new_P1_U2414;
  assign new_P1_U4995 = ~new_P1_U2497 | ~new_P1_U2401;
  assign new_P1_U4996 = ~new_P1_U4947 | ~new_P1_U2400;
  assign new_P1_U4997 = ~new_P1_U2391 | ~new_P1_U4963;
  assign new_P1_U4998 = ~P1_INSTQUEUE_REG_8__1_ | ~new_P1_U4958;
  assign new_P1_U4999 = ~new_P1_U4948 | ~new_P1_U2417;
  assign new_P1_U5000 = ~new_P1_U2497 | ~new_P1_U2399;
  assign new_P1_U5001 = ~new_P1_U4947 | ~new_P1_U2398;
  assign new_P1_U5002 = ~new_P1_U2390 | ~new_P1_U4963;
  assign new_P1_U5003 = ~P1_INSTQUEUE_REG_8__0_ | ~new_P1_U4958;
  assign new_P1_U5004 = ~new_P1_U3359;
  assign new_P1_U5005 = ~new_P1_U2439 | ~new_P1_U2442;
  assign new_P1_U5006 = ~new_P1_U3361;
  assign new_P1_U5007 = ~new_P1_U2433 | ~new_P1_U2436;
  assign new_P1_U5008 = ~new_P1_U3362;
  assign new_P1_U5009 = ~new_P1_U2500 | ~new_P1_U2358;
  assign new_P1_U5010 = ~new_P1_U3320 | ~new_P1_U5009;
  assign new_P1_U5011 = ~new_P1_U5006 | ~new_P1_U5010;
  assign new_P1_U5012 = ~P1_STATE2_REG_3_ | ~new_P1_U3356;
  assign new_P1_U5013 = ~new_P1_U5008 | ~P1_STATE2_REG_2_;
  assign new_P1_U5014 = ~new_P1_U5011 | ~new_P1_U3659;
  assign new_P1_U5015 = ~new_P1_U2500 | ~new_P1_U2388;
  assign new_P1_U5016 = ~new_P1_U3320 | ~new_P1_U5015;
  assign new_P1_U5017 = ~new_P1_U5016 | ~new_P1_U3361;
  assign new_P1_U5018 = ~P1_STATE2_REG_2_ | ~new_P1_U3362;
  assign new_P1_U5019 = ~new_P1_U5018 | ~new_P1_U5017;
  assign new_P1_U5020 = ~new_P1_U4537 | ~new_P1_U2415;
  assign new_P1_U5021 = ~new_P1_U4238 | ~new_P1_U2413;
  assign new_P1_U5022 = ~new_P1_U5004 | ~new_P1_U2412;
  assign new_P1_U5023 = ~new_P1_U2397 | ~new_P1_U5019;
  assign new_P1_U5024 = ~P1_INSTQUEUE_REG_7__7_ | ~new_P1_U5014;
  assign new_P1_U5025 = ~new_P1_U4537 | ~new_P1_U2416;
  assign new_P1_U5026 = ~new_P1_U4238 | ~new_P1_U2411;
  assign new_P1_U5027 = ~new_P1_U5004 | ~new_P1_U2410;
  assign new_P1_U5028 = ~new_P1_U2396 | ~new_P1_U5019;
  assign new_P1_U5029 = ~P1_INSTQUEUE_REG_7__6_ | ~new_P1_U5014;
  assign new_P1_U5030 = ~new_P1_U4537 | ~new_P1_U2420;
  assign new_P1_U5031 = ~new_P1_U4238 | ~new_P1_U2409;
  assign new_P1_U5032 = ~new_P1_U5004 | ~new_P1_U2408;
  assign new_P1_U5033 = ~new_P1_U2395 | ~new_P1_U5019;
  assign new_P1_U5034 = ~P1_INSTQUEUE_REG_7__5_ | ~new_P1_U5014;
  assign new_P1_U5035 = ~new_P1_U4537 | ~new_P1_U2419;
  assign new_P1_U5036 = ~new_P1_U4238 | ~new_P1_U2407;
  assign new_P1_U5037 = ~new_P1_U5004 | ~new_P1_U2406;
  assign new_P1_U5038 = ~new_P1_U2394 | ~new_P1_U5019;
  assign new_P1_U5039 = ~P1_INSTQUEUE_REG_7__4_ | ~new_P1_U5014;
  assign new_P1_U5040 = ~new_P1_U4537 | ~new_P1_U2418;
  assign new_P1_U5041 = ~new_P1_U4238 | ~new_P1_U2405;
  assign new_P1_U5042 = ~new_P1_U5004 | ~new_P1_U2404;
  assign new_P1_U5043 = ~new_P1_U2393 | ~new_P1_U5019;
  assign new_P1_U5044 = ~P1_INSTQUEUE_REG_7__3_ | ~new_P1_U5014;
  assign new_P1_U5045 = ~new_P1_U4537 | ~new_P1_U2421;
  assign new_P1_U5046 = ~new_P1_U4238 | ~new_P1_U2403;
  assign new_P1_U5047 = ~new_P1_U5004 | ~new_P1_U2402;
  assign new_P1_U5048 = ~new_P1_U2392 | ~new_P1_U5019;
  assign new_P1_U5049 = ~P1_INSTQUEUE_REG_7__2_ | ~new_P1_U5014;
  assign new_P1_U5050 = ~new_P1_U4537 | ~new_P1_U2414;
  assign new_P1_U5051 = ~new_P1_U4238 | ~new_P1_U2401;
  assign new_P1_U5052 = ~new_P1_U5004 | ~new_P1_U2400;
  assign new_P1_U5053 = ~new_P1_U2391 | ~new_P1_U5019;
  assign new_P1_U5054 = ~P1_INSTQUEUE_REG_7__1_ | ~new_P1_U5014;
  assign new_P1_U5055 = ~new_P1_U4537 | ~new_P1_U2417;
  assign new_P1_U5056 = ~new_P1_U4238 | ~new_P1_U2399;
  assign new_P1_U5057 = ~new_P1_U5004 | ~new_P1_U2398;
  assign new_P1_U5058 = ~new_P1_U2390 | ~new_P1_U5019;
  assign new_P1_U5059 = ~P1_INSTQUEUE_REG_7__0_ | ~new_P1_U5014;
  assign new_P1_U5060 = ~new_P1_U3364;
  assign new_P1_U5061 = ~new_P1_U3363;
  assign new_P1_U5062 = ~new_P1_U2439 | ~new_P1_U2443;
  assign new_P1_U5063 = ~new_P1_U3365;
  assign new_P1_U5064 = ~new_P1_U3240;
  assign new_P1_U5065 = ~new_P1_U4524 | ~new_P1_U2474;
  assign new_P1_U5066 = ~new_P1_U2502 | ~new_P1_U2358;
  assign new_P1_U5067 = ~new_P1_U3320 | ~new_P1_U5066;
  assign new_P1_U5068 = ~new_P1_U5063 | ~new_P1_U5067;
  assign new_P1_U5069 = ~P1_STATE2_REG_3_ | ~new_P1_U3363;
  assign new_P1_U5070 = ~P1_STATE2_REG_2_ | ~new_P1_U3240;
  assign new_P1_U5071 = ~new_P1_U5068 | ~new_P1_U3668;
  assign new_P1_U5072 = ~new_P1_U2502 | ~new_P1_U2388;
  assign new_P1_U5073 = ~new_P1_U3320 | ~new_P1_U5072;
  assign new_P1_U5074 = ~new_P1_U5073 | ~new_P1_U3365;
  assign new_P1_U5075 = ~P1_STATE2_REG_2_ | ~new_P1_U5064;
  assign new_P1_U5076 = ~new_P1_U5075 | ~new_P1_U5074;
  assign new_P1_U5077 = ~new_P1_U5061 | ~new_P1_U2415;
  assign new_P1_U5078 = ~new_P1_U2501 | ~new_P1_U2413;
  assign new_P1_U5079 = ~new_P1_U5060 | ~new_P1_U2412;
  assign new_P1_U5080 = ~new_P1_U2397 | ~new_P1_U5076;
  assign new_P1_U5081 = ~P1_INSTQUEUE_REG_6__7_ | ~new_P1_U5071;
  assign new_P1_U5082 = ~new_P1_U5061 | ~new_P1_U2416;
  assign new_P1_U5083 = ~new_P1_U2501 | ~new_P1_U2411;
  assign new_P1_U5084 = ~new_P1_U5060 | ~new_P1_U2410;
  assign new_P1_U5085 = ~new_P1_U2396 | ~new_P1_U5076;
  assign new_P1_U5086 = ~P1_INSTQUEUE_REG_6__6_ | ~new_P1_U5071;
  assign new_P1_U5087 = ~new_P1_U5061 | ~new_P1_U2420;
  assign new_P1_U5088 = ~new_P1_U2501 | ~new_P1_U2409;
  assign new_P1_U5089 = ~new_P1_U5060 | ~new_P1_U2408;
  assign new_P1_U5090 = ~new_P1_U2395 | ~new_P1_U5076;
  assign new_P1_U5091 = ~P1_INSTQUEUE_REG_6__5_ | ~new_P1_U5071;
  assign new_P1_U5092 = ~new_P1_U5061 | ~new_P1_U2419;
  assign new_P1_U5093 = ~new_P1_U2501 | ~new_P1_U2407;
  assign new_P1_U5094 = ~new_P1_U5060 | ~new_P1_U2406;
  assign new_P1_U5095 = ~new_P1_U2394 | ~new_P1_U5076;
  assign new_P1_U5096 = ~P1_INSTQUEUE_REG_6__4_ | ~new_P1_U5071;
  assign new_P1_U5097 = ~new_P1_U5061 | ~new_P1_U2418;
  assign new_P1_U5098 = ~new_P1_U2501 | ~new_P1_U2405;
  assign new_P1_U5099 = ~new_P1_U5060 | ~new_P1_U2404;
  assign new_P1_U5100 = ~new_P1_U2393 | ~new_P1_U5076;
  assign new_P1_U5101 = ~P1_INSTQUEUE_REG_6__3_ | ~new_P1_U5071;
  assign new_P1_U5102 = ~new_P1_U5061 | ~new_P1_U2421;
  assign new_P1_U5103 = ~new_P1_U2501 | ~new_P1_U2403;
  assign new_P1_U5104 = ~new_P1_U5060 | ~new_P1_U2402;
  assign new_P1_U5105 = ~new_P1_U2392 | ~new_P1_U5076;
  assign new_P1_U5106 = ~P1_INSTQUEUE_REG_6__2_ | ~new_P1_U5071;
  assign new_P1_U5107 = ~new_P1_U5061 | ~new_P1_U2414;
  assign new_P1_U5108 = ~new_P1_U2501 | ~new_P1_U2401;
  assign new_P1_U5109 = ~new_P1_U5060 | ~new_P1_U2400;
  assign new_P1_U5110 = ~new_P1_U2391 | ~new_P1_U5076;
  assign new_P1_U5111 = ~P1_INSTQUEUE_REG_6__1_ | ~new_P1_U5071;
  assign new_P1_U5112 = ~new_P1_U5061 | ~new_P1_U2417;
  assign new_P1_U5113 = ~new_P1_U2501 | ~new_P1_U2399;
  assign new_P1_U5114 = ~new_P1_U5060 | ~new_P1_U2398;
  assign new_P1_U5115 = ~new_P1_U2390 | ~new_P1_U5076;
  assign new_P1_U5116 = ~P1_INSTQUEUE_REG_6__0_ | ~new_P1_U5071;
  assign new_P1_U5117 = ~new_P1_U3367;
  assign new_P1_U5118 = ~new_P1_U3366;
  assign new_P1_U5119 = ~new_P1_U2439 | ~new_P1_U2444;
  assign new_P1_U5120 = ~new_P1_U3368;
  assign new_P1_U5121 = ~new_P1_U2433 | ~new_P1_U2437;
  assign new_P1_U5122 = ~new_P1_U3369;
  assign new_P1_U5123 = ~new_P1_U4525 | ~new_P1_U2474;
  assign new_P1_U5124 = ~new_P1_U2504 | ~new_P1_U2358;
  assign new_P1_U5125 = ~new_P1_U3320 | ~new_P1_U5124;
  assign new_P1_U5126 = ~new_P1_U5120 | ~new_P1_U5125;
  assign new_P1_U5127 = ~P1_STATE2_REG_3_ | ~new_P1_U3366;
  assign new_P1_U5128 = ~new_P1_U5122 | ~P1_STATE2_REG_2_;
  assign new_P1_U5129 = ~new_P1_U5126 | ~new_P1_U3677;
  assign new_P1_U5130 = ~new_P1_U2504 | ~new_P1_U2388;
  assign new_P1_U5131 = ~new_P1_U3320 | ~new_P1_U5130;
  assign new_P1_U5132 = ~new_P1_U5131 | ~new_P1_U3368;
  assign new_P1_U5133 = ~P1_STATE2_REG_2_ | ~new_P1_U3369;
  assign new_P1_U5134 = ~new_P1_U5133 | ~new_P1_U5132;
  assign new_P1_U5135 = ~new_P1_U5118 | ~new_P1_U2415;
  assign new_P1_U5136 = ~new_P1_U2503 | ~new_P1_U2413;
  assign new_P1_U5137 = ~new_P1_U5117 | ~new_P1_U2412;
  assign new_P1_U5138 = ~new_P1_U2397 | ~new_P1_U5134;
  assign new_P1_U5139 = ~P1_INSTQUEUE_REG_5__7_ | ~new_P1_U5129;
  assign new_P1_U5140 = ~new_P1_U5118 | ~new_P1_U2416;
  assign new_P1_U5141 = ~new_P1_U2503 | ~new_P1_U2411;
  assign new_P1_U5142 = ~new_P1_U5117 | ~new_P1_U2410;
  assign new_P1_U5143 = ~new_P1_U2396 | ~new_P1_U5134;
  assign new_P1_U5144 = ~P1_INSTQUEUE_REG_5__6_ | ~new_P1_U5129;
  assign new_P1_U5145 = ~new_P1_U5118 | ~new_P1_U2420;
  assign new_P1_U5146 = ~new_P1_U2503 | ~new_P1_U2409;
  assign new_P1_U5147 = ~new_P1_U5117 | ~new_P1_U2408;
  assign new_P1_U5148 = ~new_P1_U2395 | ~new_P1_U5134;
  assign new_P1_U5149 = ~P1_INSTQUEUE_REG_5__5_ | ~new_P1_U5129;
  assign new_P1_U5150 = ~new_P1_U5118 | ~new_P1_U2419;
  assign new_P1_U5151 = ~new_P1_U2503 | ~new_P1_U2407;
  assign new_P1_U5152 = ~new_P1_U5117 | ~new_P1_U2406;
  assign new_P1_U5153 = ~new_P1_U2394 | ~new_P1_U5134;
  assign new_P1_U5154 = ~P1_INSTQUEUE_REG_5__4_ | ~new_P1_U5129;
  assign new_P1_U5155 = ~new_P1_U5118 | ~new_P1_U2418;
  assign new_P1_U5156 = ~new_P1_U2503 | ~new_P1_U2405;
  assign new_P1_U5157 = ~new_P1_U5117 | ~new_P1_U2404;
  assign new_P1_U5158 = ~new_P1_U2393 | ~new_P1_U5134;
  assign new_P1_U5159 = ~P1_INSTQUEUE_REG_5__3_ | ~new_P1_U5129;
  assign new_P1_U5160 = ~new_P1_U5118 | ~new_P1_U2421;
  assign new_P1_U5161 = ~new_P1_U2503 | ~new_P1_U2403;
  assign new_P1_U5162 = ~new_P1_U5117 | ~new_P1_U2402;
  assign new_P1_U5163 = ~new_P1_U2392 | ~new_P1_U5134;
  assign new_P1_U5164 = ~P1_INSTQUEUE_REG_5__2_ | ~new_P1_U5129;
  assign new_P1_U5165 = ~new_P1_U5118 | ~new_P1_U2414;
  assign new_P1_U5166 = ~new_P1_U2503 | ~new_P1_U2401;
  assign new_P1_U5167 = ~new_P1_U5117 | ~new_P1_U2400;
  assign new_P1_U5168 = ~new_P1_U2391 | ~new_P1_U5134;
  assign new_P1_U5169 = ~P1_INSTQUEUE_REG_5__1_ | ~new_P1_U5129;
  assign new_P1_U5170 = ~new_P1_U5118 | ~new_P1_U2417;
  assign new_P1_U5171 = ~new_P1_U2503 | ~new_P1_U2399;
  assign new_P1_U5172 = ~new_P1_U5117 | ~new_P1_U2398;
  assign new_P1_U5173 = ~new_P1_U2390 | ~new_P1_U5134;
  assign new_P1_U5174 = ~P1_INSTQUEUE_REG_5__0_ | ~new_P1_U5129;
  assign new_P1_U5175 = ~new_P1_U3371;
  assign new_P1_U5176 = ~new_P1_U3370;
  assign new_P1_U5177 = ~new_P1_U2439 | ~new_P1_U2445;
  assign new_P1_U5178 = ~new_P1_U3372;
  assign new_P1_U5179 = ~new_P1_U3241;
  assign new_P1_U5180 = ~new_P1_U2486 | ~new_P1_U2474;
  assign new_P1_U5181 = ~new_P1_U2506 | ~new_P1_U2358;
  assign new_P1_U5182 = ~new_P1_U3320 | ~new_P1_U5181;
  assign new_P1_U5183 = ~new_P1_U5178 | ~new_P1_U5182;
  assign new_P1_U5184 = ~P1_STATE2_REG_3_ | ~new_P1_U3370;
  assign new_P1_U5185 = ~P1_STATE2_REG_2_ | ~new_P1_U3241;
  assign new_P1_U5186 = ~new_P1_U5183 | ~new_P1_U3686;
  assign new_P1_U5187 = ~new_P1_U2506 | ~new_P1_U2388;
  assign new_P1_U5188 = ~new_P1_U3320 | ~new_P1_U5187;
  assign new_P1_U5189 = ~new_P1_U5188 | ~new_P1_U3372;
  assign new_P1_U5190 = ~P1_STATE2_REG_2_ | ~new_P1_U5179;
  assign new_P1_U5191 = ~new_P1_U5190 | ~new_P1_U5189;
  assign new_P1_U5192 = ~new_P1_U5176 | ~new_P1_U2415;
  assign new_P1_U5193 = ~new_P1_U2505 | ~new_P1_U2413;
  assign new_P1_U5194 = ~new_P1_U5175 | ~new_P1_U2412;
  assign new_P1_U5195 = ~new_P1_U2397 | ~new_P1_U5191;
  assign new_P1_U5196 = ~P1_INSTQUEUE_REG_4__7_ | ~new_P1_U5186;
  assign new_P1_U5197 = ~new_P1_U5176 | ~new_P1_U2416;
  assign new_P1_U5198 = ~new_P1_U2505 | ~new_P1_U2411;
  assign new_P1_U5199 = ~new_P1_U5175 | ~new_P1_U2410;
  assign new_P1_U5200 = ~new_P1_U2396 | ~new_P1_U5191;
  assign new_P1_U5201 = ~P1_INSTQUEUE_REG_4__6_ | ~new_P1_U5186;
  assign new_P1_U5202 = ~new_P1_U5176 | ~new_P1_U2420;
  assign new_P1_U5203 = ~new_P1_U2505 | ~new_P1_U2409;
  assign new_P1_U5204 = ~new_P1_U5175 | ~new_P1_U2408;
  assign new_P1_U5205 = ~new_P1_U2395 | ~new_P1_U5191;
  assign new_P1_U5206 = ~P1_INSTQUEUE_REG_4__5_ | ~new_P1_U5186;
  assign new_P1_U5207 = ~new_P1_U5176 | ~new_P1_U2419;
  assign new_P1_U5208 = ~new_P1_U2505 | ~new_P1_U2407;
  assign new_P1_U5209 = ~new_P1_U5175 | ~new_P1_U2406;
  assign new_P1_U5210 = ~new_P1_U2394 | ~new_P1_U5191;
  assign new_P1_U5211 = ~P1_INSTQUEUE_REG_4__4_ | ~new_P1_U5186;
  assign new_P1_U5212 = ~new_P1_U5176 | ~new_P1_U2418;
  assign new_P1_U5213 = ~new_P1_U2505 | ~new_P1_U2405;
  assign new_P1_U5214 = ~new_P1_U5175 | ~new_P1_U2404;
  assign new_P1_U5215 = ~new_P1_U2393 | ~new_P1_U5191;
  assign new_P1_U5216 = ~P1_INSTQUEUE_REG_4__3_ | ~new_P1_U5186;
  assign new_P1_U5217 = ~new_P1_U5176 | ~new_P1_U2421;
  assign new_P1_U5218 = ~new_P1_U2505 | ~new_P1_U2403;
  assign new_P1_U5219 = ~new_P1_U5175 | ~new_P1_U2402;
  assign new_P1_U5220 = ~new_P1_U2392 | ~new_P1_U5191;
  assign new_P1_U5221 = ~P1_INSTQUEUE_REG_4__2_ | ~new_P1_U5186;
  assign new_P1_U5222 = ~new_P1_U5176 | ~new_P1_U2414;
  assign new_P1_U5223 = ~new_P1_U2505 | ~new_P1_U2401;
  assign new_P1_U5224 = ~new_P1_U5175 | ~new_P1_U2400;
  assign new_P1_U5225 = ~new_P1_U2391 | ~new_P1_U5191;
  assign new_P1_U5226 = ~P1_INSTQUEUE_REG_4__1_ | ~new_P1_U5186;
  assign new_P1_U5227 = ~new_P1_U5176 | ~new_P1_U2417;
  assign new_P1_U5228 = ~new_P1_U2505 | ~new_P1_U2399;
  assign new_P1_U5229 = ~new_P1_U5175 | ~new_P1_U2398;
  assign new_P1_U5230 = ~new_P1_U2390 | ~new_P1_U5191;
  assign new_P1_U5231 = ~P1_INSTQUEUE_REG_4__0_ | ~new_P1_U5186;
  assign new_P1_U5232 = ~new_P1_U3374;
  assign new_P1_U5233 = ~new_P1_U3373;
  assign new_P1_U5234 = ~new_P1_U2441 | ~new_P1_U2442;
  assign new_P1_U5235 = ~new_P1_U3375;
  assign new_P1_U5236 = ~new_P1_U2435 | ~new_P1_U2436;
  assign new_P1_U5237 = ~new_P1_U3376;
  assign new_P1_U5238 = ~new_P1_U2508 | ~new_P1_U4528;
  assign new_P1_U5239 = ~new_P1_U2511 | ~new_P1_U2358;
  assign new_P1_U5240 = ~new_P1_U3320 | ~new_P1_U5239;
  assign new_P1_U5241 = ~new_P1_U5235 | ~new_P1_U5240;
  assign new_P1_U5242 = ~P1_STATE2_REG_3_ | ~new_P1_U3373;
  assign new_P1_U5243 = ~new_P1_U5237 | ~P1_STATE2_REG_2_;
  assign new_P1_U5244 = ~new_P1_U5241 | ~new_P1_U3695;
  assign new_P1_U5245 = ~new_P1_U2511 | ~new_P1_U2388;
  assign new_P1_U5246 = ~new_P1_U3320 | ~new_P1_U5245;
  assign new_P1_U5247 = ~new_P1_U5246 | ~new_P1_U3375;
  assign new_P1_U5248 = ~P1_STATE2_REG_2_ | ~new_P1_U3376;
  assign new_P1_U5249 = ~new_P1_U5248 | ~new_P1_U5247;
  assign new_P1_U5250 = ~new_P1_U5233 | ~new_P1_U2415;
  assign new_P1_U5251 = ~new_P1_U2509 | ~new_P1_U2413;
  assign new_P1_U5252 = ~new_P1_U5232 | ~new_P1_U2412;
  assign new_P1_U5253 = ~new_P1_U2397 | ~new_P1_U5249;
  assign new_P1_U5254 = ~P1_INSTQUEUE_REG_3__7_ | ~new_P1_U5244;
  assign new_P1_U5255 = ~new_P1_U5233 | ~new_P1_U2416;
  assign new_P1_U5256 = ~new_P1_U2509 | ~new_P1_U2411;
  assign new_P1_U5257 = ~new_P1_U5232 | ~new_P1_U2410;
  assign new_P1_U5258 = ~new_P1_U2396 | ~new_P1_U5249;
  assign new_P1_U5259 = ~P1_INSTQUEUE_REG_3__6_ | ~new_P1_U5244;
  assign new_P1_U5260 = ~new_P1_U5233 | ~new_P1_U2420;
  assign new_P1_U5261 = ~new_P1_U2509 | ~new_P1_U2409;
  assign new_P1_U5262 = ~new_P1_U5232 | ~new_P1_U2408;
  assign new_P1_U5263 = ~new_P1_U2395 | ~new_P1_U5249;
  assign new_P1_U5264 = ~P1_INSTQUEUE_REG_3__5_ | ~new_P1_U5244;
  assign new_P1_U5265 = ~new_P1_U5233 | ~new_P1_U2419;
  assign new_P1_U5266 = ~new_P1_U2509 | ~new_P1_U2407;
  assign new_P1_U5267 = ~new_P1_U5232 | ~new_P1_U2406;
  assign new_P1_U5268 = ~new_P1_U2394 | ~new_P1_U5249;
  assign new_P1_U5269 = ~P1_INSTQUEUE_REG_3__4_ | ~new_P1_U5244;
  assign new_P1_U5270 = ~new_P1_U5233 | ~new_P1_U2418;
  assign new_P1_U5271 = ~new_P1_U2509 | ~new_P1_U2405;
  assign new_P1_U5272 = ~new_P1_U5232 | ~new_P1_U2404;
  assign new_P1_U5273 = ~new_P1_U2393 | ~new_P1_U5249;
  assign new_P1_U5274 = ~P1_INSTQUEUE_REG_3__3_ | ~new_P1_U5244;
  assign new_P1_U5275 = ~new_P1_U5233 | ~new_P1_U2421;
  assign new_P1_U5276 = ~new_P1_U2509 | ~new_P1_U2403;
  assign new_P1_U5277 = ~new_P1_U5232 | ~new_P1_U2402;
  assign new_P1_U5278 = ~new_P1_U2392 | ~new_P1_U5249;
  assign new_P1_U5279 = ~P1_INSTQUEUE_REG_3__2_ | ~new_P1_U5244;
  assign new_P1_U5280 = ~new_P1_U5233 | ~new_P1_U2414;
  assign new_P1_U5281 = ~new_P1_U2509 | ~new_P1_U2401;
  assign new_P1_U5282 = ~new_P1_U5232 | ~new_P1_U2400;
  assign new_P1_U5283 = ~new_P1_U2391 | ~new_P1_U5249;
  assign new_P1_U5284 = ~P1_INSTQUEUE_REG_3__1_ | ~new_P1_U5244;
  assign new_P1_U5285 = ~new_P1_U5233 | ~new_P1_U2417;
  assign new_P1_U5286 = ~new_P1_U2509 | ~new_P1_U2399;
  assign new_P1_U5287 = ~new_P1_U5232 | ~new_P1_U2398;
  assign new_P1_U5288 = ~new_P1_U2390 | ~new_P1_U5249;
  assign new_P1_U5289 = ~P1_INSTQUEUE_REG_3__0_ | ~new_P1_U5244;
  assign new_P1_U5290 = ~new_P1_U3378;
  assign new_P1_U5291 = ~new_P1_U3377;
  assign new_P1_U5292 = ~new_P1_U2441 | ~new_P1_U2443;
  assign new_P1_U5293 = ~new_P1_U3379;
  assign new_P1_U5294 = ~new_P1_U3242;
  assign new_P1_U5295 = ~new_P1_U2508 | ~new_P1_U4524;
  assign new_P1_U5296 = ~new_P1_U2513 | ~new_P1_U2358;
  assign new_P1_U5297 = ~new_P1_U3320 | ~new_P1_U5296;
  assign new_P1_U5298 = ~new_P1_U5293 | ~new_P1_U5297;
  assign new_P1_U5299 = ~P1_STATE2_REG_3_ | ~new_P1_U3377;
  assign new_P1_U5300 = ~P1_STATE2_REG_2_ | ~new_P1_U3242;
  assign new_P1_U5301 = ~new_P1_U5298 | ~new_P1_U3704;
  assign new_P1_U5302 = ~new_P1_U2513 | ~new_P1_U2388;
  assign new_P1_U5303 = ~new_P1_U3320 | ~new_P1_U5302;
  assign new_P1_U5304 = ~new_P1_U5303 | ~new_P1_U3379;
  assign new_P1_U5305 = ~P1_STATE2_REG_2_ | ~new_P1_U5294;
  assign new_P1_U5306 = ~new_P1_U5305 | ~new_P1_U5304;
  assign new_P1_U5307 = ~new_P1_U5291 | ~new_P1_U2415;
  assign new_P1_U5308 = ~new_P1_U2512 | ~new_P1_U2413;
  assign new_P1_U5309 = ~new_P1_U5290 | ~new_P1_U2412;
  assign new_P1_U5310 = ~new_P1_U2397 | ~new_P1_U5306;
  assign new_P1_U5311 = ~P1_INSTQUEUE_REG_2__7_ | ~new_P1_U5301;
  assign new_P1_U5312 = ~new_P1_U5291 | ~new_P1_U2416;
  assign new_P1_U5313 = ~new_P1_U2512 | ~new_P1_U2411;
  assign new_P1_U5314 = ~new_P1_U5290 | ~new_P1_U2410;
  assign new_P1_U5315 = ~new_P1_U2396 | ~new_P1_U5306;
  assign new_P1_U5316 = ~P1_INSTQUEUE_REG_2__6_ | ~new_P1_U5301;
  assign new_P1_U5317 = ~new_P1_U5291 | ~new_P1_U2420;
  assign new_P1_U5318 = ~new_P1_U2512 | ~new_P1_U2409;
  assign new_P1_U5319 = ~new_P1_U5290 | ~new_P1_U2408;
  assign new_P1_U5320 = ~new_P1_U2395 | ~new_P1_U5306;
  assign new_P1_U5321 = ~P1_INSTQUEUE_REG_2__5_ | ~new_P1_U5301;
  assign new_P1_U5322 = ~new_P1_U5291 | ~new_P1_U2419;
  assign new_P1_U5323 = ~new_P1_U2512 | ~new_P1_U2407;
  assign new_P1_U5324 = ~new_P1_U5290 | ~new_P1_U2406;
  assign new_P1_U5325 = ~new_P1_U2394 | ~new_P1_U5306;
  assign new_P1_U5326 = ~P1_INSTQUEUE_REG_2__4_ | ~new_P1_U5301;
  assign new_P1_U5327 = ~new_P1_U5291 | ~new_P1_U2418;
  assign new_P1_U5328 = ~new_P1_U2512 | ~new_P1_U2405;
  assign new_P1_U5329 = ~new_P1_U5290 | ~new_P1_U2404;
  assign new_P1_U5330 = ~new_P1_U2393 | ~new_P1_U5306;
  assign new_P1_U5331 = ~P1_INSTQUEUE_REG_2__3_ | ~new_P1_U5301;
  assign new_P1_U5332 = ~new_P1_U5291 | ~new_P1_U2421;
  assign new_P1_U5333 = ~new_P1_U2512 | ~new_P1_U2403;
  assign new_P1_U5334 = ~new_P1_U5290 | ~new_P1_U2402;
  assign new_P1_U5335 = ~new_P1_U2392 | ~new_P1_U5306;
  assign new_P1_U5336 = ~P1_INSTQUEUE_REG_2__2_ | ~new_P1_U5301;
  assign new_P1_U5337 = ~new_P1_U5291 | ~new_P1_U2414;
  assign new_P1_U5338 = ~new_P1_U2512 | ~new_P1_U2401;
  assign new_P1_U5339 = ~new_P1_U5290 | ~new_P1_U2400;
  assign new_P1_U5340 = ~new_P1_U2391 | ~new_P1_U5306;
  assign new_P1_U5341 = ~P1_INSTQUEUE_REG_2__1_ | ~new_P1_U5301;
  assign new_P1_U5342 = ~new_P1_U5291 | ~new_P1_U2417;
  assign new_P1_U5343 = ~new_P1_U2512 | ~new_P1_U2399;
  assign new_P1_U5344 = ~new_P1_U5290 | ~new_P1_U2398;
  assign new_P1_U5345 = ~new_P1_U2390 | ~new_P1_U5306;
  assign new_P1_U5346 = ~P1_INSTQUEUE_REG_2__0_ | ~new_P1_U5301;
  assign new_P1_U5347 = ~new_P1_U3381;
  assign new_P1_U5348 = ~new_P1_U3380;
  assign new_P1_U5349 = ~new_P1_U2441 | ~new_P1_U2444;
  assign new_P1_U5350 = ~new_P1_U3382;
  assign new_P1_U5351 = ~new_P1_U2435 | ~new_P1_U2437;
  assign new_P1_U5352 = ~new_P1_U3383;
  assign new_P1_U5353 = ~new_P1_U2508 | ~new_P1_U4525;
  assign new_P1_U5354 = ~new_P1_U2515 | ~new_P1_U2358;
  assign new_P1_U5355 = ~new_P1_U3320 | ~new_P1_U5354;
  assign new_P1_U5356 = ~new_P1_U5350 | ~new_P1_U5355;
  assign new_P1_U5357 = ~P1_STATE2_REG_3_ | ~new_P1_U3380;
  assign new_P1_U5358 = ~new_P1_U5352 | ~P1_STATE2_REG_2_;
  assign new_P1_U5359 = ~new_P1_U5356 | ~new_P1_U3713;
  assign new_P1_U5360 = ~new_P1_U2515 | ~new_P1_U2388;
  assign new_P1_U5361 = ~new_P1_U3320 | ~new_P1_U5360;
  assign new_P1_U5362 = ~new_P1_U5361 | ~new_P1_U3382;
  assign new_P1_U5363 = ~P1_STATE2_REG_2_ | ~new_P1_U3383;
  assign new_P1_U5364 = ~new_P1_U5363 | ~new_P1_U5362;
  assign new_P1_U5365 = ~new_P1_U5348 | ~new_P1_U2415;
  assign new_P1_U5366 = ~new_P1_U2514 | ~new_P1_U2413;
  assign new_P1_U5367 = ~new_P1_U5347 | ~new_P1_U2412;
  assign new_P1_U5368 = ~new_P1_U2397 | ~new_P1_U5364;
  assign new_P1_U5369 = ~P1_INSTQUEUE_REG_1__7_ | ~new_P1_U5359;
  assign new_P1_U5370 = ~new_P1_U5348 | ~new_P1_U2416;
  assign new_P1_U5371 = ~new_P1_U2514 | ~new_P1_U2411;
  assign new_P1_U5372 = ~new_P1_U5347 | ~new_P1_U2410;
  assign new_P1_U5373 = ~new_P1_U2396 | ~new_P1_U5364;
  assign new_P1_U5374 = ~P1_INSTQUEUE_REG_1__6_ | ~new_P1_U5359;
  assign new_P1_U5375 = ~new_P1_U5348 | ~new_P1_U2420;
  assign new_P1_U5376 = ~new_P1_U2514 | ~new_P1_U2409;
  assign new_P1_U5377 = ~new_P1_U5347 | ~new_P1_U2408;
  assign new_P1_U5378 = ~new_P1_U2395 | ~new_P1_U5364;
  assign new_P1_U5379 = ~P1_INSTQUEUE_REG_1__5_ | ~new_P1_U5359;
  assign new_P1_U5380 = ~new_P1_U5348 | ~new_P1_U2419;
  assign new_P1_U5381 = ~new_P1_U2514 | ~new_P1_U2407;
  assign new_P1_U5382 = ~new_P1_U5347 | ~new_P1_U2406;
  assign new_P1_U5383 = ~new_P1_U2394 | ~new_P1_U5364;
  assign new_P1_U5384 = ~P1_INSTQUEUE_REG_1__4_ | ~new_P1_U5359;
  assign new_P1_U5385 = ~new_P1_U5348 | ~new_P1_U2418;
  assign new_P1_U5386 = ~new_P1_U2514 | ~new_P1_U2405;
  assign new_P1_U5387 = ~new_P1_U5347 | ~new_P1_U2404;
  assign new_P1_U5388 = ~new_P1_U2393 | ~new_P1_U5364;
  assign new_P1_U5389 = ~P1_INSTQUEUE_REG_1__3_ | ~new_P1_U5359;
  assign new_P1_U5390 = ~new_P1_U5348 | ~new_P1_U2421;
  assign new_P1_U5391 = ~new_P1_U2514 | ~new_P1_U2403;
  assign new_P1_U5392 = ~new_P1_U5347 | ~new_P1_U2402;
  assign new_P1_U5393 = ~new_P1_U2392 | ~new_P1_U5364;
  assign new_P1_U5394 = ~P1_INSTQUEUE_REG_1__2_ | ~new_P1_U5359;
  assign new_P1_U5395 = ~new_P1_U5348 | ~new_P1_U2414;
  assign new_P1_U5396 = ~new_P1_U2514 | ~new_P1_U2401;
  assign new_P1_U5397 = ~new_P1_U5347 | ~new_P1_U2400;
  assign new_P1_U5398 = ~new_P1_U2391 | ~new_P1_U5364;
  assign new_P1_U5399 = ~P1_INSTQUEUE_REG_1__1_ | ~new_P1_U5359;
  assign new_P1_U5400 = ~new_P1_U5348 | ~new_P1_U2417;
  assign new_P1_U5401 = ~new_P1_U2514 | ~new_P1_U2399;
  assign new_P1_U5402 = ~new_P1_U5347 | ~new_P1_U2398;
  assign new_P1_U5403 = ~new_P1_U2390 | ~new_P1_U5364;
  assign new_P1_U5404 = ~P1_INSTQUEUE_REG_1__0_ | ~new_P1_U5359;
  assign new_P1_U5405 = ~new_P1_U3385;
  assign new_P1_U5406 = ~new_P1_U3384;
  assign new_P1_U5407 = ~new_P1_U2441 | ~new_P1_U2445;
  assign new_P1_U5408 = ~new_P1_U3386;
  assign new_P1_U5409 = ~new_P1_U3243;
  assign new_P1_U5410 = ~new_P1_U2508 | ~new_P1_U2486;
  assign new_P1_U5411 = ~new_P1_U2517 | ~new_P1_U2358;
  assign new_P1_U5412 = ~new_P1_U3320 | ~new_P1_U5411;
  assign new_P1_U5413 = ~new_P1_U5408 | ~new_P1_U5412;
  assign new_P1_U5414 = ~P1_STATE2_REG_3_ | ~new_P1_U3384;
  assign new_P1_U5415 = ~P1_STATE2_REG_2_ | ~new_P1_U3243;
  assign new_P1_U5416 = ~new_P1_U5413 | ~new_P1_U3722;
  assign new_P1_U5417 = ~new_P1_U2517 | ~new_P1_U2388;
  assign new_P1_U5418 = ~new_P1_U3320 | ~new_P1_U5417;
  assign new_P1_U5419 = ~new_P1_U5418 | ~new_P1_U3386;
  assign new_P1_U5420 = ~P1_STATE2_REG_2_ | ~new_P1_U5409;
  assign new_P1_U5421 = ~new_P1_U5420 | ~new_P1_U5419;
  assign new_P1_U5422 = ~new_P1_U5406 | ~new_P1_U2415;
  assign new_P1_U5423 = ~new_P1_U2516 | ~new_P1_U2413;
  assign new_P1_U5424 = ~new_P1_U5405 | ~new_P1_U2412;
  assign new_P1_U5425 = ~new_P1_U2397 | ~new_P1_U5421;
  assign new_P1_U5426 = ~P1_INSTQUEUE_REG_0__7_ | ~new_P1_U5416;
  assign new_P1_U5427 = ~new_P1_U5406 | ~new_P1_U2416;
  assign new_P1_U5428 = ~new_P1_U2516 | ~new_P1_U2411;
  assign new_P1_U5429 = ~new_P1_U5405 | ~new_P1_U2410;
  assign new_P1_U5430 = ~new_P1_U2396 | ~new_P1_U5421;
  assign new_P1_U5431 = ~P1_INSTQUEUE_REG_0__6_ | ~new_P1_U5416;
  assign new_P1_U5432 = ~new_P1_U5406 | ~new_P1_U2420;
  assign new_P1_U5433 = ~new_P1_U2516 | ~new_P1_U2409;
  assign new_P1_U5434 = ~new_P1_U5405 | ~new_P1_U2408;
  assign new_P1_U5435 = ~new_P1_U2395 | ~new_P1_U5421;
  assign new_P1_U5436 = ~P1_INSTQUEUE_REG_0__5_ | ~new_P1_U5416;
  assign new_P1_U5437 = ~new_P1_U5406 | ~new_P1_U2419;
  assign new_P1_U5438 = ~new_P1_U2516 | ~new_P1_U2407;
  assign new_P1_U5439 = ~new_P1_U5405 | ~new_P1_U2406;
  assign new_P1_U5440 = ~new_P1_U2394 | ~new_P1_U5421;
  assign new_P1_U5441 = ~new_P1_U5406 | ~new_P1_U2418;
  assign new_P1_U5442 = ~new_P1_U2516 | ~new_P1_U2405;
  assign new_P1_U5443 = ~new_P1_U5405 | ~new_P1_U2404;
  assign new_P1_U5444 = ~new_P1_U2393 | ~new_P1_U5421;
  assign new_P1_U5445 = ~P1_INSTQUEUE_REG_0__3_ | ~new_P1_U5416;
  assign new_P1_U5446 = ~new_P1_U5406 | ~new_P1_U2421;
  assign new_P1_U5447 = ~new_P1_U2516 | ~new_P1_U2403;
  assign new_P1_U5448 = ~new_P1_U5405 | ~new_P1_U2402;
  assign new_P1_U5449 = ~new_P1_U2392 | ~new_P1_U5421;
  assign new_P1_U5450 = ~P1_INSTQUEUE_REG_0__2_ | ~new_P1_U5416;
  assign new_P1_U5451 = ~new_P1_U5406 | ~new_P1_U2414;
  assign new_P1_U5452 = ~new_P1_U2516 | ~new_P1_U2401;
  assign new_P1_U5453 = ~new_P1_U5405 | ~new_P1_U2400;
  assign new_P1_U5454 = ~new_P1_U2391 | ~new_P1_U5421;
  assign new_P1_U5455 = ~P1_INSTQUEUE_REG_0__1_ | ~new_P1_U5416;
  assign new_P1_U5456 = ~new_P1_U5406 | ~new_P1_U2417;
  assign new_P1_U5457 = ~new_P1_U2516 | ~new_P1_U2399;
  assign new_P1_U5458 = ~new_P1_U5405 | ~new_P1_U2398;
  assign new_P1_U5459 = ~new_P1_U2390 | ~new_P1_U5421;
  assign new_P1_U5460 = ~P1_INSTQUEUE_REG_0__0_ | ~new_P1_U5416;
  assign new_P1_U5461 = ~new_P1_U3423;
  assign new_P1_U5462 = ~new_P1_U4503 | ~new_P1_U3391 | ~new_P1_U3394;
  assign new_P1_U5463 = ~new_P1_U4460 | ~new_P1_U4400 | ~new_P1_U4173;
  assign new_P1_U5464 = ~new_P1_U3244;
  assign new_P1_U5465 = ~new_P1_U4494 | ~new_P1_U3289;
  assign new_P1_U5466 = ~new_P1_U5464 | ~new_P1_U5465 | ~new_P1_U3283;
  assign new_P1_U5467 = ~new_P1_U3732 | ~new_P1_U2452;
  assign new_P1_U5468 = ~new_P1_U4208 | ~new_P1_U5462;
  assign new_P1_U5469 = ~new_P1_U3733 | ~new_P1_U7609;
  assign new_P1_U5470 = ~new_P1_GTE_485_U6 | ~new_P1_U4215 | ~new_P1_U3257;
  assign new_P1_U5471 = ~new_P1_U2449 | ~new_P1_U7494;
  assign new_P1_U5472 = ~new_P1_U4257 | ~new_P1_U4503;
  assign new_P1_U5473 = ~new_P1_U4182;
  assign new_P1_U5474 = ~new_P1_U2368 | ~new_P1_U4182;
  assign new_P1_U5475 = ~P1_STATE2_REG_3_ | ~new_P1_U3294;
  assign new_P1_U5476 = ~new_P1_U4172;
  assign new_P1_U5477 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U5478 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U5477;
  assign new_P1_U5479 = ~new_P1_U4381 | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U5480 = ~new_P1_U3442;
  assign new_P1_U5481 = ~new_P1_U3498 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U5482 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U5481;
  assign new_P1_U5483 = ~new_P1_U3438;
  assign new_P1_U5484 = ~new_P1_U3275 | ~new_P1_U3264;
  assign new_P1_U5485 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U5484;
  assign new_P1_U5486 = ~new_P1_U2469 | ~new_P1_U3275;
  assign new_P1_U5487 = ~new_P1_U4494 | ~new_P1_U3290;
  assign new_P1_U5488 = ~new_P1_U4400 | ~new_P1_U2605;
  assign new_P1_U5489 = ~new_P1_U7494 | ~new_P1_U7704 | ~new_P1_U7703;
  assign new_P1_U5490 = ~new_P1_U4449 | ~new_P1_U5488;
  assign new_P1_U5491 = ~new_P1_U3409 | ~new_P1_U4400 | ~new_P1_U3394;
  assign new_P1_U5492 = ~new_P1_U5491 | ~new_P1_U4171;
  assign new_P1_U5493 = ~new_P1_U7629 | ~new_P1_U5492;
  assign new_P1_U5494 = ~new_P1_U4460 | ~new_P1_U4171;
  assign new_P1_U5495 = ~new_P1_U3395 | ~new_P1_U5494;
  assign new_P1_U5496 = ~new_P1_U4208 | ~new_P1_U5462;
  assign new_P1_U5497 = ~new_P1_U4257 | ~new_P1_U4503;
  assign new_P1_U5498 = ~new_P1_U5495 | ~new_P1_U3271;
  assign new_P1_U5499 = ~new_P1_U4494 | ~new_P1_U7707;
  assign new_P1_U5500 = ~new_P1_U4190 | ~new_P1_U3244;
  assign new_P1_U5501 = ~new_P1_U3292 | ~new_P1_U4217;
  assign new_P1_U5502 = ~new_P1_U3740 | ~new_P1_U5501;
  assign new_P1_U5503 = ~new_P1_R2182_U25 | ~new_P1_U7509;
  assign new_P1_U5504 = ~new_P1_U4218 | ~new_P1_U3438;
  assign new_P1_U5505 = ~new_P1_U4214 | ~new_P1_U3442;
  assign new_P1_U5506 = ~new_P1_U5503 | ~new_P1_U3747;
  assign new_P1_U5507 = ~new_P1_U4252 | ~new_P1_U3438;
  assign new_P1_U5508 = ~new_P1_U2427 | ~new_P1_U5506;
  assign new_P1_U5509 = ~new_P1_U5508 | ~new_P1_U5507;
  assign new_P1_U5510 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3275;
  assign new_P1_U5511 = ~new_P1_U3401;
  assign new_P1_U5512 = ~new_P1_R2182_U42 | ~new_P1_U7509;
  assign new_P1_U5513 = ~new_P1_U4214 | ~new_P1_U3456;
  assign new_P1_U5514 = ~new_P1_U3749 | ~new_P1_U5512;
  assign new_P1_U5515 = ~new_P1_U2446 | ~new_P1_U3470;
  assign new_P1_U5516 = ~new_P1_U4252 | ~new_P1_U3401;
  assign new_P1_U5517 = ~new_P1_U2427 | ~new_P1_U5514;
  assign new_P1_U5518 = ~new_P1_U5516 | ~new_P1_U5517 | ~new_P1_U5515;
  assign new_P1_U5519 = ~new_P1_U3402;
  assign new_P1_U5520 = ~new_P1_U2431 | ~new_P1_U4249;
  assign new_P1_U5521 = ~new_P1_U3292 | ~new_P1_U5520;
  assign new_P1_U5522 = ~new_P1_U5519 | ~new_P1_U5521;
  assign new_P1_U5523 = ~new_P1_R2182_U33 | ~new_P1_U7509;
  assign new_P1_U5524 = ~new_P1_U4214 | ~new_P1_U3265;
  assign new_P1_U5525 = ~new_P1_U3750 | ~new_P1_U5523;
  assign new_P1_U5526 = ~new_P1_U7712 | ~new_P1_U2446;
  assign new_P1_U5527 = ~new_P1_U5519 | ~new_P1_U4252;
  assign new_P1_U5528 = ~new_P1_U2427 | ~new_P1_U5525;
  assign new_P1_U5529 = ~new_P1_U5527 | ~new_P1_U5528 | ~new_P1_U5526;
  assign new_P1_U5530 = ~new_P1_R2182_U34 | ~new_P1_U7509;
  assign new_P1_U5531 = ~new_P1_U4175 | ~new_P1_U5530;
  assign new_P1_U5532 = ~new_P1_U4252 | ~new_P1_U3266;
  assign new_P1_U5533 = ~new_P1_U2427 | ~new_P1_U5531;
  assign new_P1_U5534 = ~new_P1_U7715 | ~P1_STATE2_REG_1_;
  assign new_P1_U5535 = ~new_P1_U5532 | ~new_P1_U5533 | ~new_P1_U5534;
  assign new_P1_U5536 = ~new_P1_LT_589_U6 | ~new_P1_U2428 | ~P1_STATE2_REG_0_;
  assign new_P1_U5537 = ~new_P1_U3404;
  assign new_P1_U5538 = ~P1_STATE2_REG_1_ | ~new_P1_U3296;
  assign new_P1_U5539 = ~new_P1_U4527 | ~new_P1_U3454;
  assign new_P1_U5540 = ~new_P1_U3358 | ~new_P1_U5539;
  assign new_P1_U5541 = ~new_P1_U3359 | ~new_P1_U5540;
  assign new_P1_U5542 = ~new_P1_U2388 | ~new_P1_U5541;
  assign new_P1_U5543 = ~new_P1_R2182_U25 | ~new_P1_U5538;
  assign new_P1_U5544 = ~new_P1_U4226 | ~new_P1_R2144_U8;
  assign new_P1_U5545 = ~new_P1_U3751 | ~new_P1_U5542;
  assign new_P1_U5546 = ~new_P1_U2388 | ~new_P1_U7733;
  assign new_P1_U5547 = ~new_P1_R2182_U42 | ~new_P1_U5538;
  assign new_P1_U5548 = ~new_P1_U4226 | ~new_P1_R2144_U49;
  assign new_P1_U5549 = ~new_P1_U3752 | ~new_P1_U5546;
  assign new_P1_U5550 = ~new_P1_U3326 | ~new_P1_U3333;
  assign new_P1_U5551 = ~new_P1_U2388 | ~new_P1_U5550;
  assign new_P1_U5552 = ~new_P1_R2182_U33 | ~new_P1_U5538;
  assign new_P1_U5553 = ~new_P1_U4226 | ~new_P1_R2144_U50;
  assign new_P1_U5554 = ~new_P1_U3753 | ~new_P1_U5551;
  assign new_P1_U5555 = ~new_P1_R2182_U34 | ~new_P1_U5538;
  assign new_P1_U5556 = ~new_P1_R2144_U43 | ~new_P1_U4209;
  assign new_P1_U5557 = ~new_P1_U4245 | ~new_P1_U5555 | ~new_P1_U5556;
  assign new_P1_U5558 = ~new_P1_U4477 | ~new_P1_U3272;
  assign new_P1_U5559 = ~new_P1_U4260 | ~new_P1_U2431;
  assign new_P1_U5560 = ~new_P1_U7742 | ~new_P1_U7743 | ~new_P1_U2518 | ~new_P1_U5559;
  assign new_P1_U5561 = ~new_P1_U4192 | ~new_P1_U4235 | ~new_P1_U4503;
  assign new_P1_U5562 = ~new_P1_U2368 | ~new_P1_U5560;
  assign new_P1_U5563 = ~new_P1_U4203 | ~new_P1_U3263;
  assign new_P1_U5564 = ~new_P1_U3414;
  assign new_P1_U5565 = ~new_P1_U4262 | ~new_P1_U4208;
  assign new_P1_U5566 = ~new_P1_U4256 | ~new_P1_U2389;
  assign new_P1_U5567 = ~new_P1_U4266 | ~new_P1_U4250;
  assign new_P1_U5568 = ~new_P1_U4264 | ~new_P1_U4494;
  assign new_P1_U5569 = ~new_P1_U3758 | ~new_P1_U2519;
  assign new_P1_U5570 = ~new_P1_R2099_U86 | ~new_P1_U2380;
  assign new_P1_U5571 = ~new_P1_R2027_U5 | ~new_P1_U2378;
  assign new_P1_U5572 = ~new_P1_R2278_U99 | ~new_P1_U2377;
  assign new_P1_U5573 = ~new_P1_ADD_405_U4 | ~new_P1_U2375;
  assign new_P1_U5574 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_U2374;
  assign new_P1_U5575 = ~P1_REIP_REG_0_ | ~new_P1_U2370;
  assign new_P1_U5576 = ~new_P1_U5564 | ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_U5577 = ~new_P1_R2099_U87 | ~new_P1_U2380;
  assign new_P1_U5578 = ~new_P1_R2027_U71 | ~new_P1_U2378;
  assign new_P1_U5579 = ~new_P1_R2278_U19 | ~new_P1_U2377;
  assign new_P1_U5580 = ~new_P1_ADD_405_U85 | ~new_P1_U2375;
  assign new_P1_U5581 = ~new_P1_ADD_515_U4 | ~new_P1_U2374;
  assign new_P1_U5582 = ~new_P1_U2370 | ~P1_REIP_REG_1_;
  assign new_P1_U5583 = ~new_P1_U5564 | ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_U5584 = ~new_P1_R2099_U138 | ~new_P1_U2380;
  assign new_P1_U5585 = ~new_P1_R2027_U60 | ~new_P1_U2378;
  assign new_P1_U5586 = ~new_P1_R2278_U107 | ~new_P1_U2377;
  assign new_P1_U5587 = ~new_P1_ADD_405_U5 | ~new_P1_U2375;
  assign new_P1_U5588 = ~new_P1_ADD_515_U67 | ~new_P1_U2374;
  assign new_P1_U5589 = ~new_P1_U2370 | ~P1_REIP_REG_2_;
  assign new_P1_U5590 = ~P1_INSTADDRPOINTER_REG_2_ | ~new_P1_U5564;
  assign new_P1_U5591 = ~new_P1_R2099_U42 | ~new_P1_U2380;
  assign new_P1_U5592 = ~new_P1_R2027_U57 | ~new_P1_U2378;
  assign new_P1_U5593 = ~new_P1_R2278_U105 | ~new_P1_U2377;
  assign new_P1_U5594 = ~new_P1_ADD_405_U95 | ~new_P1_U2375;
  assign new_P1_U5595 = ~new_P1_ADD_515_U85 | ~new_P1_U2374;
  assign new_P1_U5596 = ~new_P1_U2370 | ~P1_REIP_REG_3_;
  assign new_P1_U5597 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_U5564;
  assign new_P1_U5598 = ~new_P1_R2099_U41 | ~new_P1_U2380;
  assign new_P1_U5599 = ~new_P1_R2027_U56 | ~new_P1_U2378;
  assign new_P1_U5600 = ~new_P1_R2278_U104 | ~new_P1_U2377;
  assign new_P1_U5601 = ~new_P1_ADD_405_U76 | ~new_P1_U2375;
  assign new_P1_U5602 = ~new_P1_ADD_515_U76 | ~new_P1_U2374;
  assign new_P1_U5603 = ~new_P1_U2370 | ~P1_REIP_REG_4_;
  assign new_P1_U5604 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_U5564;
  assign new_P1_U5605 = ~new_P1_R2099_U40 | ~new_P1_U2380;
  assign new_P1_U5606 = ~new_P1_R2027_U55 | ~new_P1_U2378;
  assign new_P1_U5607 = ~new_P1_R2278_U17 | ~new_P1_U2377;
  assign new_P1_U5608 = ~new_P1_ADD_405_U79 | ~new_P1_U2375;
  assign new_P1_U5609 = ~new_P1_ADD_515_U79 | ~new_P1_U2374;
  assign new_P1_U5610 = ~new_P1_U2370 | ~P1_REIP_REG_5_;
  assign new_P1_U5611 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_U5564;
  assign new_P1_U5612 = ~new_P1_R2099_U39 | ~new_P1_U2380;
  assign new_P1_U5613 = ~new_P1_R2027_U54 | ~new_P1_U2378;
  assign new_P1_U5614 = ~new_P1_R2278_U103 | ~new_P1_U2377;
  assign new_P1_U5615 = ~new_P1_ADD_405_U63 | ~new_P1_U2375;
  assign new_P1_U5616 = ~new_P1_ADD_515_U62 | ~new_P1_U2374;
  assign new_P1_U5617 = ~new_P1_U2370 | ~P1_REIP_REG_6_;
  assign new_P1_U5618 = ~P1_INSTADDRPOINTER_REG_6_ | ~new_P1_U5564;
  assign new_P1_U5619 = ~new_P1_R2099_U38 | ~new_P1_U2380;
  assign new_P1_U5620 = ~new_P1_R2027_U53 | ~new_P1_U2378;
  assign new_P1_U5621 = ~new_P1_R2278_U18 | ~new_P1_U2377;
  assign new_P1_U5622 = ~new_P1_ADD_405_U89 | ~new_P1_U2375;
  assign new_P1_U5623 = ~new_P1_ADD_515_U89 | ~new_P1_U2374;
  assign new_P1_U5624 = ~new_P1_U2370 | ~P1_REIP_REG_7_;
  assign new_P1_U5625 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_U5564;
  assign new_P1_U5626 = ~new_P1_R2099_U37 | ~new_P1_U2380;
  assign new_P1_U5627 = ~new_P1_R2027_U52 | ~new_P1_U2378;
  assign new_P1_U5628 = ~new_P1_R2278_U102 | ~new_P1_U2377;
  assign new_P1_U5629 = ~new_P1_ADD_405_U80 | ~new_P1_U2375;
  assign new_P1_U5630 = ~new_P1_ADD_515_U80 | ~new_P1_U2374;
  assign new_P1_U5631 = ~new_P1_U2370 | ~P1_REIP_REG_8_;
  assign new_P1_U5632 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_U5564;
  assign new_P1_U5633 = ~new_P1_R2099_U36 | ~new_P1_U2380;
  assign new_P1_U5634 = ~new_P1_R2027_U51 | ~new_P1_U2378;
  assign new_P1_U5635 = ~new_P1_R2278_U101 | ~new_P1_U2377;
  assign new_P1_U5636 = ~new_P1_ADD_405_U70 | ~new_P1_U2375;
  assign new_P1_U5637 = ~new_P1_ADD_515_U70 | ~new_P1_U2374;
  assign new_P1_U5638 = ~new_P1_U2370 | ~P1_REIP_REG_9_;
  assign new_P1_U5639 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_U5564;
  assign new_P1_U5640 = ~new_P1_R2099_U85 | ~new_P1_U2380;
  assign new_P1_U5641 = ~new_P1_R2027_U81 | ~new_P1_U2378;
  assign new_P1_U5642 = ~new_P1_R2278_U126 | ~new_P1_U2377;
  assign new_P1_U5643 = ~new_P1_ADD_405_U83 | ~new_P1_U2375;
  assign new_P1_U5644 = ~new_P1_ADD_515_U83 | ~new_P1_U2374;
  assign new_P1_U5645 = ~new_P1_U2370 | ~P1_REIP_REG_10_;
  assign new_P1_U5646 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_U5564;
  assign new_P1_U5647 = ~new_P1_R2099_U84 | ~new_P1_U2380;
  assign new_P1_U5648 = ~new_P1_R2027_U80 | ~new_P1_U2378;
  assign new_P1_U5649 = ~new_P1_R2278_U15 | ~new_P1_U2377;
  assign new_P1_U5650 = ~new_P1_ADD_405_U73 | ~new_P1_U2375;
  assign new_P1_U5651 = ~new_P1_ADD_515_U73 | ~new_P1_U2374;
  assign new_P1_U5652 = ~new_P1_U2370 | ~P1_REIP_REG_11_;
  assign new_P1_U5653 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_U5564;
  assign new_P1_U5654 = ~new_P1_R2099_U83 | ~new_P1_U2380;
  assign new_P1_U5655 = ~new_P1_R2027_U79 | ~new_P1_U2378;
  assign new_P1_U5656 = ~new_P1_R2278_U125 | ~new_P1_U2377;
  assign new_P1_U5657 = ~new_P1_ADD_405_U88 | ~new_P1_U2375;
  assign new_P1_U5658 = ~new_P1_ADD_515_U88 | ~new_P1_U2374;
  assign new_P1_U5659 = ~new_P1_U2370 | ~P1_REIP_REG_12_;
  assign new_P1_U5660 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_U5564;
  assign new_P1_U5661 = ~new_P1_R2099_U82 | ~new_P1_U2380;
  assign new_P1_U5662 = ~new_P1_R2027_U78 | ~new_P1_U2378;
  assign new_P1_U5663 = ~new_P1_R2278_U123 | ~new_P1_U2377;
  assign new_P1_U5664 = ~new_P1_ADD_405_U69 | ~new_P1_U2375;
  assign new_P1_U5665 = ~new_P1_ADD_515_U69 | ~new_P1_U2374;
  assign new_P1_U5666 = ~new_P1_U2370 | ~P1_REIP_REG_13_;
  assign new_P1_U5667 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_U5564;
  assign new_P1_U5668 = ~new_P1_R2099_U81 | ~new_P1_U2380;
  assign new_P1_U5669 = ~new_P1_R2027_U77 | ~new_P1_U2378;
  assign new_P1_U5670 = ~new_P1_R2278_U122 | ~new_P1_U2377;
  assign new_P1_U5671 = ~new_P1_ADD_405_U78 | ~new_P1_U2375;
  assign new_P1_U5672 = ~new_P1_ADD_515_U78 | ~new_P1_U2374;
  assign new_P1_U5673 = ~new_P1_U2370 | ~P1_REIP_REG_14_;
  assign new_P1_U5674 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_U5564;
  assign new_P1_U5675 = ~new_P1_R2099_U80 | ~new_P1_U2380;
  assign new_P1_U5676 = ~new_P1_R2027_U76 | ~new_P1_U2378;
  assign new_P1_U5677 = ~new_P1_R2278_U20 | ~new_P1_U2377;
  assign new_P1_U5678 = ~new_P1_ADD_405_U75 | ~new_P1_U2375;
  assign new_P1_U5679 = ~new_P1_ADD_515_U75 | ~new_P1_U2374;
  assign new_P1_U5680 = ~new_P1_U2370 | ~P1_REIP_REG_15_;
  assign new_P1_U5681 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_U5564;
  assign new_P1_U5682 = ~new_P1_R2099_U79 | ~new_P1_U2380;
  assign new_P1_U5683 = ~new_P1_R2027_U75 | ~new_P1_U2378;
  assign new_P1_U5684 = ~new_P1_R2278_U121 | ~new_P1_U2377;
  assign new_P1_U5685 = ~new_P1_ADD_405_U91 | ~new_P1_U2375;
  assign new_P1_U5686 = ~new_P1_ADD_515_U91 | ~new_P1_U2374;
  assign new_P1_U5687 = ~new_P1_U2370 | ~P1_REIP_REG_16_;
  assign new_P1_U5688 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_U5564;
  assign new_P1_U5689 = ~new_P1_R2099_U78 | ~new_P1_U2380;
  assign new_P1_U5690 = ~new_P1_R2027_U74 | ~new_P1_U2378;
  assign new_P1_U5691 = ~new_P1_R2278_U120 | ~new_P1_U2377;
  assign new_P1_U5692 = ~new_P1_ADD_405_U67 | ~new_P1_U2375;
  assign new_P1_U5693 = ~new_P1_ADD_515_U66 | ~new_P1_U2374;
  assign new_P1_U5694 = ~new_P1_U2370 | ~P1_REIP_REG_17_;
  assign new_P1_U5695 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_U5564;
  assign new_P1_U5696 = ~new_P1_R2099_U77 | ~new_P1_U2380;
  assign new_P1_U5697 = ~new_P1_R2027_U73 | ~new_P1_U2378;
  assign new_P1_U5698 = ~new_P1_R2278_U119 | ~new_P1_U2377;
  assign new_P1_U5699 = ~new_P1_ADD_405_U72 | ~new_P1_U2375;
  assign new_P1_U5700 = ~new_P1_ADD_515_U72 | ~new_P1_U2374;
  assign new_P1_U5701 = ~new_P1_U2370 | ~P1_REIP_REG_18_;
  assign new_P1_U5702 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_U5564;
  assign new_P1_U5703 = ~new_P1_R2099_U76 | ~new_P1_U2380;
  assign new_P1_U5704 = ~new_P1_R2027_U72 | ~new_P1_U2378;
  assign new_P1_U5705 = ~new_P1_R2278_U118 | ~new_P1_U2377;
  assign new_P1_U5706 = ~new_P1_ADD_405_U82 | ~new_P1_U2375;
  assign new_P1_U5707 = ~new_P1_ADD_515_U82 | ~new_P1_U2374;
  assign new_P1_U5708 = ~new_P1_U2370 | ~P1_REIP_REG_19_;
  assign new_P1_U5709 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_U5564;
  assign new_P1_U5710 = ~new_P1_R2099_U75 | ~new_P1_U2380;
  assign new_P1_U5711 = ~new_P1_R2027_U70 | ~new_P1_U2378;
  assign new_P1_U5712 = ~new_P1_R2278_U117 | ~new_P1_U2377;
  assign new_P1_U5713 = ~new_P1_ADD_405_U68 | ~new_P1_U2375;
  assign new_P1_U5714 = ~new_P1_ADD_515_U68 | ~new_P1_U2374;
  assign new_P1_U5715 = ~new_P1_U2370 | ~P1_REIP_REG_20_;
  assign new_P1_U5716 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_U5564;
  assign new_P1_U5717 = ~new_P1_R2099_U74 | ~new_P1_U2380;
  assign new_P1_U5718 = ~new_P1_R2027_U69 | ~new_P1_U2378;
  assign new_P1_U5719 = ~new_P1_R2278_U116 | ~new_P1_U2377;
  assign new_P1_U5720 = ~new_P1_ADD_405_U87 | ~new_P1_U2375;
  assign new_P1_U5721 = ~new_P1_ADD_515_U87 | ~new_P1_U2374;
  assign new_P1_U5722 = ~new_P1_U2370 | ~P1_REIP_REG_21_;
  assign new_P1_U5723 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_U5564;
  assign new_P1_U5724 = ~new_P1_R2099_U73 | ~new_P1_U2380;
  assign new_P1_U5725 = ~new_P1_R2027_U68 | ~new_P1_U2378;
  assign new_P1_U5726 = ~new_P1_R2278_U115 | ~new_P1_U2377;
  assign new_P1_U5727 = ~new_P1_ADD_405_U71 | ~new_P1_U2375;
  assign new_P1_U5728 = ~new_P1_ADD_515_U71 | ~new_P1_U2374;
  assign new_P1_U5729 = ~new_P1_U2370 | ~P1_REIP_REG_22_;
  assign new_P1_U5730 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_U5564;
  assign new_P1_U5731 = ~new_P1_R2099_U72 | ~new_P1_U2380;
  assign new_P1_U5732 = ~new_P1_R2027_U67 | ~new_P1_U2378;
  assign new_P1_U5733 = ~new_P1_R2278_U114 | ~new_P1_U2377;
  assign new_P1_U5734 = ~new_P1_ADD_405_U81 | ~new_P1_U2375;
  assign new_P1_U5735 = ~new_P1_ADD_515_U81 | ~new_P1_U2374;
  assign new_P1_U5736 = ~new_P1_U2370 | ~P1_REIP_REG_23_;
  assign new_P1_U5737 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_U5564;
  assign new_P1_U5738 = ~new_P1_R2099_U71 | ~new_P1_U2380;
  assign new_P1_U5739 = ~new_P1_R2027_U66 | ~new_P1_U2378;
  assign new_P1_U5740 = ~new_P1_R2278_U113 | ~new_P1_U2377;
  assign new_P1_U5741 = ~new_P1_ADD_405_U66 | ~new_P1_U2375;
  assign new_P1_U5742 = ~new_P1_ADD_515_U65 | ~new_P1_U2374;
  assign new_P1_U5743 = ~new_P1_U2370 | ~P1_REIP_REG_24_;
  assign new_P1_U5744 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_U5564;
  assign new_P1_U5745 = ~new_P1_R2099_U70 | ~new_P1_U2380;
  assign new_P1_U5746 = ~new_P1_R2027_U65 | ~new_P1_U2378;
  assign new_P1_U5747 = ~new_P1_R2278_U112 | ~new_P1_U2377;
  assign new_P1_U5748 = ~new_P1_ADD_405_U90 | ~new_P1_U2375;
  assign new_P1_U5749 = ~new_P1_ADD_515_U90 | ~new_P1_U2374;
  assign new_P1_U5750 = ~new_P1_U2370 | ~P1_REIP_REG_25_;
  assign new_P1_U5751 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_U5564;
  assign new_P1_U5752 = ~new_P1_R2099_U69 | ~new_P1_U2380;
  assign new_P1_U5753 = ~new_P1_R2027_U64 | ~new_P1_U2378;
  assign new_P1_U5754 = ~new_P1_R2278_U111 | ~new_P1_U2377;
  assign new_P1_U5755 = ~new_P1_ADD_405_U74 | ~new_P1_U2375;
  assign new_P1_U5756 = ~new_P1_ADD_515_U74 | ~new_P1_U2374;
  assign new_P1_U5757 = ~new_P1_U2370 | ~P1_REIP_REG_26_;
  assign new_P1_U5758 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_U5564;
  assign new_P1_U5759 = ~new_P1_R2099_U68 | ~new_P1_U2380;
  assign new_P1_U5760 = ~new_P1_R2027_U63 | ~new_P1_U2378;
  assign new_P1_U5761 = ~new_P1_R2278_U110 | ~new_P1_U2377;
  assign new_P1_U5762 = ~new_P1_ADD_405_U77 | ~new_P1_U2375;
  assign new_P1_U5763 = ~new_P1_ADD_515_U77 | ~new_P1_U2374;
  assign new_P1_U5764 = ~new_P1_U2370 | ~P1_REIP_REG_27_;
  assign new_P1_U5765 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_U5564;
  assign new_P1_U5766 = ~new_P1_R2099_U67 | ~new_P1_U2380;
  assign new_P1_U5767 = ~new_P1_R2027_U62 | ~new_P1_U2378;
  assign new_P1_U5768 = ~new_P1_R2278_U109 | ~new_P1_U2377;
  assign new_P1_U5769 = ~new_P1_ADD_405_U86 | ~new_P1_U2375;
  assign new_P1_U5770 = ~new_P1_ADD_515_U86 | ~new_P1_U2374;
  assign new_P1_U5771 = ~new_P1_U2370 | ~P1_REIP_REG_28_;
  assign new_P1_U5772 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_U5564;
  assign new_P1_U5773 = ~new_P1_R2099_U66 | ~new_P1_U2380;
  assign new_P1_U5774 = ~new_P1_R2027_U61 | ~new_P1_U2378;
  assign new_P1_U5775 = ~new_P1_R2278_U108 | ~new_P1_U2377;
  assign new_P1_U5776 = ~new_P1_ADD_405_U65 | ~new_P1_U2375;
  assign new_P1_U5777 = ~new_P1_ADD_515_U64 | ~new_P1_U2374;
  assign new_P1_U5778 = ~new_P1_U2370 | ~P1_REIP_REG_29_;
  assign new_P1_U5779 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_U5564;
  assign new_P1_U5780 = ~new_P1_R2099_U65 | ~new_P1_U2380;
  assign new_P1_U5781 = ~new_P1_R2027_U59 | ~new_P1_U2378;
  assign new_P1_U5782 = ~new_P1_R2278_U106 | ~new_P1_U2377;
  assign new_P1_U5783 = ~new_P1_ADD_405_U64 | ~new_P1_U2375;
  assign new_P1_U5784 = ~new_P1_ADD_515_U63 | ~new_P1_U2374;
  assign new_P1_U5785 = ~new_P1_U2370 | ~P1_REIP_REG_30_;
  assign new_P1_U5786 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_U5564;
  assign new_P1_U5787 = ~new_P1_R2099_U64 | ~new_P1_U2380;
  assign new_P1_U5788 = ~new_P1_R2027_U58 | ~new_P1_U2378;
  assign new_P1_U5789 = ~new_P1_R2278_U16 | ~new_P1_U2377;
  assign new_P1_U5790 = ~new_P1_ADD_405_U84 | ~new_P1_U2375;
  assign new_P1_U5791 = ~new_P1_ADD_515_U84 | ~new_P1_U2374;
  assign new_P1_U5792 = ~new_P1_U2370 | ~P1_REIP_REG_31_;
  assign new_P1_U5793 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_U5564;
  assign new_P1_U5794 = ~new_P1_U4209 | ~new_P1_U3294;
  assign new_P1_U5795 = ~new_P1_U3416;
  assign new_P1_U5796 = ~P1_STATE2_REG_2_ | ~new_P1_U3294;
  assign new_P1_U5797 = ~P1_STATE2_REG_1_ | ~new_P1_U3308;
  assign new_P1_U5798 = ~new_P1_U5797 | ~new_P1_U5796;
  assign new_P1_U5799 = ~P1_PHYADDRPOINTER_REG_0_ | ~new_P1_U2376;
  assign new_P1_U5800 = ~new_P1_U2372 | ~new_P1_R2278_U99;
  assign new_P1_U5801 = ~new_P1_U2365 | ~P1_REIP_REG_0_;
  assign new_P1_U5802 = ~new_P1_R2358_U76 | ~new_P1_U2364;
  assign new_P1_U5803 = ~P1_PHYADDRPOINTER_REG_0_ | ~new_P1_U5795;
  assign new_P1_U5804 = ~new_P1_R2337_U4 | ~new_P1_U2376;
  assign new_P1_U5805 = ~new_P1_U2372 | ~new_P1_R2278_U19;
  assign new_P1_U5806 = ~new_P1_U2365 | ~P1_REIP_REG_1_;
  assign new_P1_U5807 = ~new_P1_R2358_U107 | ~new_P1_U2364;
  assign new_P1_U5808 = ~P1_PHYADDRPOINTER_REG_1_ | ~new_P1_U5795;
  assign new_P1_U5809 = ~new_P1_R2337_U71 | ~new_P1_U2376;
  assign new_P1_U5810 = ~new_P1_U2372 | ~new_P1_R2278_U107;
  assign new_P1_U5811 = ~new_P1_U2365 | ~P1_REIP_REG_2_;
  assign new_P1_U5812 = ~new_P1_R2358_U18 | ~new_P1_U2364;
  assign new_P1_U5813 = ~P1_PHYADDRPOINTER_REG_2_ | ~new_P1_U5795;
  assign new_P1_U5814 = ~new_P1_R2337_U68 | ~new_P1_U2376;
  assign new_P1_U5815 = ~new_P1_U2372 | ~new_P1_R2278_U105;
  assign new_P1_U5816 = ~new_P1_U2365 | ~P1_REIP_REG_3_;
  assign new_P1_U5817 = ~new_P1_R2358_U19 | ~new_P1_U2364;
  assign new_P1_U5818 = ~P1_PHYADDRPOINTER_REG_3_ | ~new_P1_U5795;
  assign new_P1_U5819 = ~new_P1_R2337_U67 | ~new_P1_U2376;
  assign new_P1_U5820 = ~new_P1_U2372 | ~new_P1_R2278_U104;
  assign new_P1_U5821 = ~new_P1_U2365 | ~P1_REIP_REG_4_;
  assign new_P1_U5822 = ~new_P1_R2358_U84 | ~new_P1_U2364;
  assign new_P1_U5823 = ~P1_PHYADDRPOINTER_REG_4_ | ~new_P1_U5795;
  assign new_P1_U5824 = ~new_P1_R2337_U66 | ~new_P1_U2376;
  assign new_P1_U5825 = ~new_P1_U2372 | ~new_P1_R2278_U17;
  assign new_P1_U5826 = ~new_P1_U2365 | ~P1_REIP_REG_5_;
  assign new_P1_U5827 = ~new_P1_R2358_U82 | ~new_P1_U2364;
  assign new_P1_U5828 = ~P1_PHYADDRPOINTER_REG_5_ | ~new_P1_U5795;
  assign new_P1_U5829 = ~new_P1_R2337_U65 | ~new_P1_U2376;
  assign new_P1_U5830 = ~new_P1_U2372 | ~new_P1_R2278_U103;
  assign new_P1_U5831 = ~new_P1_U2365 | ~P1_REIP_REG_6_;
  assign new_P1_U5832 = ~new_P1_R2358_U20 | ~new_P1_U2364;
  assign new_P1_U5833 = ~P1_PHYADDRPOINTER_REG_6_ | ~new_P1_U5795;
  assign new_P1_U5834 = ~new_P1_R2337_U64 | ~new_P1_U2376;
  assign new_P1_U5835 = ~new_P1_U2372 | ~new_P1_R2278_U18;
  assign new_P1_U5836 = ~new_P1_U2365 | ~P1_REIP_REG_7_;
  assign new_P1_U5837 = ~new_P1_R2358_U21 | ~new_P1_U2364;
  assign new_P1_U5838 = ~P1_PHYADDRPOINTER_REG_7_ | ~new_P1_U5795;
  assign new_P1_U5839 = ~new_P1_R2337_U63 | ~new_P1_U2376;
  assign new_P1_U5840 = ~new_P1_U2372 | ~new_P1_R2278_U102;
  assign new_P1_U5841 = ~new_P1_U2365 | ~P1_REIP_REG_8_;
  assign new_P1_U5842 = ~new_P1_R2358_U80 | ~new_P1_U2364;
  assign new_P1_U5843 = ~P1_PHYADDRPOINTER_REG_8_ | ~new_P1_U5795;
  assign new_P1_U5844 = ~new_P1_R2337_U62 | ~new_P1_U2376;
  assign new_P1_U5845 = ~new_P1_U2372 | ~new_P1_R2278_U101;
  assign new_P1_U5846 = ~new_P1_U2365 | ~P1_REIP_REG_9_;
  assign new_P1_U5847 = ~new_P1_R2358_U78 | ~new_P1_U2364;
  assign new_P1_U5848 = ~P1_PHYADDRPOINTER_REG_9_ | ~new_P1_U5795;
  assign new_P1_U5849 = ~new_P1_R2337_U91 | ~new_P1_U2376;
  assign new_P1_U5850 = ~new_P1_U2372 | ~new_P1_R2278_U126;
  assign new_P1_U5851 = ~new_P1_U2365 | ~P1_REIP_REG_10_;
  assign new_P1_U5852 = ~new_P1_R2358_U14 | ~new_P1_U2364;
  assign new_P1_U5853 = ~P1_PHYADDRPOINTER_REG_10_ | ~new_P1_U5795;
  assign new_P1_U5854 = ~new_P1_R2337_U90 | ~new_P1_U2376;
  assign new_P1_U5855 = ~new_P1_U2372 | ~new_P1_R2278_U15;
  assign new_P1_U5856 = ~new_P1_U2365 | ~P1_REIP_REG_11_;
  assign new_P1_U5857 = ~new_P1_R2358_U15 | ~new_P1_U2364;
  assign new_P1_U5858 = ~P1_PHYADDRPOINTER_REG_11_ | ~new_P1_U5795;
  assign new_P1_U5859 = ~new_P1_R2337_U89 | ~new_P1_U2376;
  assign new_P1_U5860 = ~new_P1_U2372 | ~new_P1_R2278_U125;
  assign new_P1_U5861 = ~new_P1_U2365 | ~P1_REIP_REG_12_;
  assign new_P1_U5862 = ~new_P1_R2358_U119 | ~new_P1_U2364;
  assign new_P1_U5863 = ~P1_PHYADDRPOINTER_REG_12_ | ~new_P1_U5795;
  assign new_P1_U5864 = ~new_P1_R2337_U88 | ~new_P1_U2376;
  assign new_P1_U5865 = ~new_P1_U2372 | ~new_P1_R2278_U123;
  assign new_P1_U5866 = ~new_P1_U2365 | ~P1_REIP_REG_13_;
  assign new_P1_U5867 = ~new_P1_R2358_U117 | ~new_P1_U2364;
  assign new_P1_U5868 = ~P1_PHYADDRPOINTER_REG_13_ | ~new_P1_U5795;
  assign new_P1_U5869 = ~new_P1_R2337_U87 | ~new_P1_U2376;
  assign new_P1_U5870 = ~new_P1_U2372 | ~new_P1_R2278_U122;
  assign new_P1_U5871 = ~new_P1_U2365 | ~P1_REIP_REG_14_;
  assign new_P1_U5872 = ~new_P1_R2358_U16 | ~new_P1_U2364;
  assign new_P1_U5873 = ~P1_PHYADDRPOINTER_REG_14_ | ~new_P1_U5795;
  assign new_P1_U5874 = ~new_P1_R2337_U86 | ~new_P1_U2376;
  assign new_P1_U5875 = ~new_P1_U2372 | ~new_P1_R2278_U20;
  assign new_P1_U5876 = ~new_P1_U2365 | ~P1_REIP_REG_15_;
  assign new_P1_U5877 = ~new_P1_R2358_U17 | ~new_P1_U2364;
  assign new_P1_U5878 = ~P1_PHYADDRPOINTER_REG_15_ | ~new_P1_U5795;
  assign new_P1_U5879 = ~new_P1_R2337_U85 | ~new_P1_U2376;
  assign new_P1_U5880 = ~new_P1_U2372 | ~new_P1_R2278_U121;
  assign new_P1_U5881 = ~new_P1_U2365 | ~P1_REIP_REG_16_;
  assign new_P1_U5882 = ~new_P1_R2358_U115 | ~new_P1_U2364;
  assign new_P1_U5883 = ~P1_PHYADDRPOINTER_REG_16_ | ~new_P1_U5795;
  assign new_P1_U5884 = ~new_P1_R2337_U84 | ~new_P1_U2376;
  assign new_P1_U5885 = ~new_P1_U2372 | ~new_P1_R2278_U120;
  assign new_P1_U5886 = ~new_P1_U2365 | ~P1_REIP_REG_17_;
  assign new_P1_U5887 = ~new_P1_R2358_U113 | ~new_P1_U2364;
  assign new_P1_U5888 = ~P1_PHYADDRPOINTER_REG_17_ | ~new_P1_U5795;
  assign new_P1_U5889 = ~new_P1_R2337_U83 | ~new_P1_U2376;
  assign new_P1_U5890 = ~new_P1_U2372 | ~new_P1_R2278_U119;
  assign new_P1_U5891 = ~new_P1_U2365 | ~P1_REIP_REG_18_;
  assign new_P1_U5892 = ~new_P1_R2358_U111 | ~new_P1_U2364;
  assign new_P1_U5893 = ~P1_PHYADDRPOINTER_REG_18_ | ~new_P1_U5795;
  assign new_P1_U5894 = ~new_P1_R2337_U82 | ~new_P1_U2376;
  assign new_P1_U5895 = ~new_P1_U2372 | ~new_P1_R2278_U118;
  assign new_P1_U5896 = ~new_P1_U2365 | ~P1_REIP_REG_19_;
  assign new_P1_U5897 = ~new_P1_R2358_U109 | ~new_P1_U2364;
  assign new_P1_U5898 = ~P1_PHYADDRPOINTER_REG_19_ | ~new_P1_U5795;
  assign new_P1_U5899 = ~new_P1_R2337_U81 | ~new_P1_U2376;
  assign new_P1_U5900 = ~new_P1_U2372 | ~new_P1_R2278_U117;
  assign new_P1_U5901 = ~new_P1_U2365 | ~P1_REIP_REG_20_;
  assign new_P1_U5902 = ~new_P1_R2358_U105 | ~new_P1_U2364;
  assign new_P1_U5903 = ~P1_PHYADDRPOINTER_REG_20_ | ~new_P1_U5795;
  assign new_P1_U5904 = ~new_P1_R2337_U80 | ~new_P1_U2376;
  assign new_P1_U5905 = ~new_P1_U2372 | ~new_P1_R2278_U116;
  assign new_P1_U5906 = ~new_P1_U2365 | ~P1_REIP_REG_21_;
  assign new_P1_U5907 = ~new_P1_R2358_U103 | ~new_P1_U2364;
  assign new_P1_U5908 = ~P1_PHYADDRPOINTER_REG_21_ | ~new_P1_U5795;
  assign new_P1_U5909 = ~new_P1_R2337_U79 | ~new_P1_U2376;
  assign new_P1_U5910 = ~new_P1_U2372 | ~new_P1_R2278_U115;
  assign new_P1_U5911 = ~new_P1_U2365 | ~P1_REIP_REG_22_;
  assign new_P1_U5912 = ~new_P1_R2358_U101 | ~new_P1_U2364;
  assign new_P1_U5913 = ~P1_PHYADDRPOINTER_REG_22_ | ~new_P1_U5795;
  assign new_P1_U5914 = ~new_P1_R2337_U78 | ~new_P1_U2376;
  assign new_P1_U5915 = ~new_P1_U2372 | ~new_P1_R2278_U114;
  assign new_P1_U5916 = ~new_P1_U2365 | ~P1_REIP_REG_23_;
  assign new_P1_U5917 = ~new_P1_R2358_U99 | ~new_P1_U2364;
  assign new_P1_U5918 = ~P1_PHYADDRPOINTER_REG_23_ | ~new_P1_U5795;
  assign new_P1_U5919 = ~new_P1_R2337_U77 | ~new_P1_U2376;
  assign new_P1_U5920 = ~new_P1_U2372 | ~new_P1_R2278_U113;
  assign new_P1_U5921 = ~new_P1_U2365 | ~P1_REIP_REG_24_;
  assign new_P1_U5922 = ~new_P1_R2358_U97 | ~new_P1_U2364;
  assign new_P1_U5923 = ~P1_PHYADDRPOINTER_REG_24_ | ~new_P1_U5795;
  assign new_P1_U5924 = ~new_P1_R2337_U76 | ~new_P1_U2376;
  assign new_P1_U5925 = ~new_P1_U2372 | ~new_P1_R2278_U112;
  assign new_P1_U5926 = ~new_P1_U2365 | ~P1_REIP_REG_25_;
  assign new_P1_U5927 = ~new_P1_R2358_U95 | ~new_P1_U2364;
  assign new_P1_U5928 = ~P1_PHYADDRPOINTER_REG_25_ | ~new_P1_U5795;
  assign new_P1_U5929 = ~new_P1_R2337_U75 | ~new_P1_U2376;
  assign new_P1_U5930 = ~new_P1_U2372 | ~new_P1_R2278_U111;
  assign new_P1_U5931 = ~new_P1_U2365 | ~P1_REIP_REG_26_;
  assign new_P1_U5932 = ~new_P1_R2358_U93 | ~new_P1_U2364;
  assign new_P1_U5933 = ~P1_PHYADDRPOINTER_REG_26_ | ~new_P1_U5795;
  assign new_P1_U5934 = ~new_P1_R2337_U74 | ~new_P1_U2376;
  assign new_P1_U5935 = ~new_P1_U2372 | ~new_P1_R2278_U110;
  assign new_P1_U5936 = ~new_P1_U2365 | ~P1_REIP_REG_27_;
  assign new_P1_U5937 = ~new_P1_R2358_U91 | ~new_P1_U2364;
  assign new_P1_U5938 = ~P1_PHYADDRPOINTER_REG_27_ | ~new_P1_U5795;
  assign new_P1_U5939 = ~new_P1_R2337_U73 | ~new_P1_U2376;
  assign new_P1_U5940 = ~new_P1_U2372 | ~new_P1_R2278_U109;
  assign new_P1_U5941 = ~new_P1_U2365 | ~P1_REIP_REG_28_;
  assign new_P1_U5942 = ~new_P1_R2358_U89 | ~new_P1_U2364;
  assign new_P1_U5943 = ~P1_PHYADDRPOINTER_REG_28_ | ~new_P1_U5795;
  assign new_P1_U5944 = ~new_P1_R2337_U72 | ~new_P1_U2376;
  assign new_P1_U5945 = ~new_P1_U2372 | ~new_P1_R2278_U108;
  assign new_P1_U5946 = ~new_P1_U2365 | ~P1_REIP_REG_29_;
  assign new_P1_U5947 = ~new_P1_R2358_U87 | ~new_P1_U2364;
  assign new_P1_U5948 = ~P1_PHYADDRPOINTER_REG_29_ | ~new_P1_U5795;
  assign new_P1_U5949 = ~new_P1_R2337_U70 | ~new_P1_U2376;
  assign new_P1_U5950 = ~new_P1_U2372 | ~new_P1_R2278_U106;
  assign new_P1_U5951 = ~new_P1_U2365 | ~P1_REIP_REG_30_;
  assign new_P1_U5952 = ~new_P1_R2358_U85 | ~new_P1_U2364;
  assign new_P1_U5953 = ~P1_PHYADDRPOINTER_REG_30_ | ~new_P1_U5795;
  assign new_P1_U5954 = ~new_P1_R2337_U69 | ~new_P1_U2376;
  assign new_P1_U5955 = ~new_P1_U2372 | ~new_P1_R2278_U16;
  assign new_P1_U5956 = ~new_P1_U2365 | ~P1_REIP_REG_31_;
  assign new_P1_U5957 = ~new_P1_R2358_U22 | ~new_P1_U2364;
  assign new_P1_U5958 = ~P1_PHYADDRPOINTER_REG_31_ | ~new_P1_U5795;
  assign new_P1_U5959 = ~new_U210 | ~new_P1_U3282;
  assign new_P1_U5960 = ~P1_EAX_REG_15_ | ~new_P1_U2382;
  assign new_P1_U5961 = ~new_U340 | ~new_P1_U2381;
  assign new_P1_U5962 = ~new_P1_U5961 | ~new_P1_U5960;
  assign new_P1_U5963 = ~P1_EAX_REG_14_ | ~new_P1_U2382;
  assign new_P1_U5964 = ~new_U341 | ~new_P1_U2381;
  assign new_P1_U5965 = ~new_P1_U5964 | ~new_P1_U5963;
  assign new_P1_U5966 = ~P1_EAX_REG_13_ | ~new_P1_U2382;
  assign new_P1_U5967 = ~new_U342 | ~new_P1_U2381;
  assign new_P1_U5968 = ~new_P1_U5967 | ~new_P1_U5966;
  assign new_P1_U5969 = ~P1_EAX_REG_12_ | ~new_P1_U2382;
  assign new_P1_U5970 = ~new_U343 | ~new_P1_U2381;
  assign new_P1_U5971 = ~new_P1_U5970 | ~new_P1_U5969;
  assign new_P1_U5972 = ~P1_EAX_REG_11_ | ~new_P1_U2382;
  assign new_P1_U5973 = ~new_U344 | ~new_P1_U2381;
  assign new_P1_U5974 = ~new_P1_U5973 | ~new_P1_U5972;
  assign new_P1_U5975 = ~P1_EAX_REG_10_ | ~new_P1_U2382;
  assign new_P1_U5976 = ~new_U345 | ~new_P1_U2381;
  assign new_P1_U5977 = ~new_P1_U5976 | ~new_P1_U5975;
  assign new_P1_U5978 = ~P1_EAX_REG_9_ | ~new_P1_U2382;
  assign new_P1_U5979 = ~new_U315 | ~new_P1_U2381;
  assign new_P1_U5980 = ~new_P1_U5979 | ~new_P1_U5978;
  assign new_P1_U5981 = ~P1_EAX_REG_8_ | ~new_P1_U2382;
  assign new_P1_U5982 = ~new_U316 | ~new_P1_U2381;
  assign new_P1_U5983 = ~new_P1_U5982 | ~new_P1_U5981;
  assign new_P1_U5984 = ~P1_EAX_REG_7_ | ~new_P1_U2382;
  assign new_P1_U5985 = ~new_P1_U2381 | ~new_U317;
  assign new_P1_U5986 = ~new_P1_U5985 | ~new_P1_U5984;
  assign new_P1_U5987 = ~P1_EAX_REG_6_ | ~new_P1_U2382;
  assign new_P1_U5988 = ~new_P1_U2381 | ~new_U318;
  assign new_P1_U5989 = ~new_P1_U5988 | ~new_P1_U5987;
  assign new_P1_U5990 = ~P1_EAX_REG_5_ | ~new_P1_U2382;
  assign new_P1_U5991 = ~new_P1_U2381 | ~new_U319;
  assign new_P1_U5992 = ~new_P1_U5991 | ~new_P1_U5990;
  assign new_P1_U5993 = ~P1_EAX_REG_4_ | ~new_P1_U2382;
  assign new_P1_U5994 = ~new_P1_U2381 | ~new_U320;
  assign new_P1_U5995 = ~new_P1_U5994 | ~new_P1_U5993;
  assign new_P1_U5996 = ~P1_EAX_REG_3_ | ~new_P1_U2382;
  assign new_P1_U5997 = ~new_P1_U2381 | ~new_U321;
  assign new_P1_U5998 = ~new_P1_U5997 | ~new_P1_U5996;
  assign new_P1_U5999 = ~P1_EAX_REG_2_ | ~new_P1_U2382;
  assign new_P1_U6000 = ~new_P1_U2381 | ~new_U324;
  assign new_P1_U6001 = ~new_P1_U6000 | ~new_P1_U5999;
  assign new_P1_U6002 = ~P1_EAX_REG_1_ | ~new_P1_U2382;
  assign new_P1_U6003 = ~new_P1_U2381 | ~new_U335;
  assign new_P1_U6004 = ~new_P1_U6003 | ~new_P1_U6002;
  assign new_P1_U6005 = ~P1_EAX_REG_0_ | ~new_P1_U2382;
  assign new_P1_U6006 = ~new_P1_U2381 | ~new_U346;
  assign new_P1_U6007 = ~new_P1_U6006 | ~new_P1_U6005;
  assign new_P1_U6008 = ~P1_EAX_REG_30_ | ~new_P1_U2382;
  assign new_P1_U6009 = ~new_U341 | ~new_P1_U2381;
  assign new_P1_U6010 = ~new_P1_U6009 | ~new_P1_U6008;
  assign new_P1_U6011 = ~P1_EAX_REG_29_ | ~new_P1_U2382;
  assign new_P1_U6012 = ~new_U342 | ~new_P1_U2381;
  assign new_P1_U6013 = ~new_P1_U6012 | ~new_P1_U6011;
  assign new_P1_U6014 = ~P1_EAX_REG_28_ | ~new_P1_U2382;
  assign new_P1_U6015 = ~new_U343 | ~new_P1_U2381;
  assign new_P1_U6016 = ~new_P1_U6015 | ~new_P1_U6014;
  assign new_P1_U6017 = ~P1_EAX_REG_27_ | ~new_P1_U2382;
  assign new_P1_U6018 = ~new_U344 | ~new_P1_U2381;
  assign new_P1_U6019 = ~new_P1_U6018 | ~new_P1_U6017;
  assign new_P1_U6020 = ~P1_EAX_REG_26_ | ~new_P1_U2382;
  assign new_P1_U6021 = ~new_U345 | ~new_P1_U2381;
  assign new_P1_U6022 = ~new_P1_U6021 | ~new_P1_U6020;
  assign new_P1_U6023 = ~P1_EAX_REG_25_ | ~new_P1_U2382;
  assign new_P1_U6024 = ~new_U315 | ~new_P1_U2381;
  assign new_P1_U6025 = ~new_P1_U6024 | ~new_P1_U6023;
  assign new_P1_U6026 = ~P1_EAX_REG_24_ | ~new_P1_U2382;
  assign new_P1_U6027 = ~new_U316 | ~new_P1_U2381;
  assign new_P1_U6028 = ~new_P1_U6027 | ~new_P1_U6026;
  assign new_P1_U6029 = ~P1_EAX_REG_23_ | ~new_P1_U2382;
  assign new_P1_U6030 = ~new_P1_U2381 | ~new_U317;
  assign new_P1_U6031 = ~new_P1_U6030 | ~new_P1_U6029;
  assign new_P1_U6032 = ~P1_EAX_REG_22_ | ~new_P1_U2382;
  assign new_P1_U6033 = ~new_P1_U2381 | ~new_U318;
  assign new_P1_U6034 = ~new_P1_U6033 | ~new_P1_U6032;
  assign new_P1_U6035 = ~P1_EAX_REG_21_ | ~new_P1_U2382;
  assign new_P1_U6036 = ~new_P1_U2381 | ~new_U319;
  assign new_P1_U6037 = ~new_P1_U6036 | ~new_P1_U6035;
  assign new_P1_U6038 = ~P1_EAX_REG_20_ | ~new_P1_U2382;
  assign new_P1_U6039 = ~new_P1_U2381 | ~new_U320;
  assign new_P1_U6040 = ~new_P1_U6039 | ~new_P1_U6038;
  assign new_P1_U6041 = ~P1_EAX_REG_19_ | ~new_P1_U2382;
  assign new_P1_U6042 = ~new_P1_U2381 | ~new_U321;
  assign new_P1_U6043 = ~new_P1_U6042 | ~new_P1_U6041;
  assign new_P1_U6044 = ~P1_EAX_REG_18_ | ~new_P1_U2382;
  assign new_P1_U6045 = ~new_P1_U2381 | ~new_U324;
  assign new_P1_U6046 = ~new_P1_U6045 | ~new_P1_U6044;
  assign new_P1_U6047 = ~P1_EAX_REG_17_ | ~new_P1_U2382;
  assign new_P1_U6048 = ~new_P1_U2381 | ~new_U335;
  assign new_P1_U6049 = ~new_P1_U6048 | ~new_P1_U6047;
  assign new_P1_U6050 = ~P1_EAX_REG_16_ | ~new_P1_U2382;
  assign new_P1_U6051 = ~new_P1_U2381 | ~new_U346;
  assign new_P1_U6052 = ~new_P1_U6051 | ~new_P1_U6050;
  assign new_P1_U6053 = ~new_P1_U4259 | ~new_P1_U4235 | ~new_P1_U7606;
  assign new_P1_U6054 = ~new_P1_U2428 | ~new_P1_U3294;
  assign new_P1_U6055 = ~new_P1_U3417;
  assign new_P1_U6056 = ~new_P1_U2385 | ~P1_LWORD_REG_0_;
  assign new_P1_U6057 = ~new_P1_U2384 | ~P1_EAX_REG_0_;
  assign new_P1_U6058 = ~P1_DATAO_REG_0_ | ~new_P1_U6055;
  assign new_P1_U6059 = ~new_P1_U2385 | ~P1_LWORD_REG_1_;
  assign new_P1_U6060 = ~new_P1_U2384 | ~P1_EAX_REG_1_;
  assign new_P1_U6061 = ~P1_DATAO_REG_1_ | ~new_P1_U6055;
  assign new_P1_U6062 = ~new_P1_U2385 | ~P1_LWORD_REG_2_;
  assign new_P1_U6063 = ~new_P1_U2384 | ~P1_EAX_REG_2_;
  assign new_P1_U6064 = ~P1_DATAO_REG_2_ | ~new_P1_U6055;
  assign new_P1_U6065 = ~new_P1_U2385 | ~P1_LWORD_REG_3_;
  assign new_P1_U6066 = ~new_P1_U2384 | ~P1_EAX_REG_3_;
  assign new_P1_U6067 = ~P1_DATAO_REG_3_ | ~new_P1_U6055;
  assign new_P1_U6068 = ~new_P1_U2385 | ~P1_LWORD_REG_4_;
  assign new_P1_U6069 = ~new_P1_U2384 | ~P1_EAX_REG_4_;
  assign new_P1_U6070 = ~P1_DATAO_REG_4_ | ~new_P1_U6055;
  assign new_P1_U6071 = ~new_P1_U2385 | ~P1_LWORD_REG_5_;
  assign new_P1_U6072 = ~new_P1_U2384 | ~P1_EAX_REG_5_;
  assign new_P1_U6073 = ~P1_DATAO_REG_5_ | ~new_P1_U6055;
  assign new_P1_U6074 = ~new_P1_U2385 | ~P1_LWORD_REG_6_;
  assign new_P1_U6075 = ~new_P1_U2384 | ~P1_EAX_REG_6_;
  assign new_P1_U6076 = ~P1_DATAO_REG_6_ | ~new_P1_U6055;
  assign new_P1_U6077 = ~new_P1_U2385 | ~P1_LWORD_REG_7_;
  assign new_P1_U6078 = ~new_P1_U2384 | ~P1_EAX_REG_7_;
  assign new_P1_U6079 = ~P1_DATAO_REG_7_ | ~new_P1_U6055;
  assign new_P1_U6080 = ~new_P1_U2385 | ~P1_LWORD_REG_8_;
  assign new_P1_U6081 = ~new_P1_U2384 | ~P1_EAX_REG_8_;
  assign new_P1_U6082 = ~P1_DATAO_REG_8_ | ~new_P1_U6055;
  assign new_P1_U6083 = ~new_P1_U2385 | ~P1_LWORD_REG_9_;
  assign new_P1_U6084 = ~new_P1_U2384 | ~P1_EAX_REG_9_;
  assign new_P1_U6085 = ~P1_DATAO_REG_9_ | ~new_P1_U6055;
  assign new_P1_U6086 = ~new_P1_U2385 | ~P1_LWORD_REG_10_;
  assign new_P1_U6087 = ~new_P1_U2384 | ~P1_EAX_REG_10_;
  assign new_P1_U6088 = ~P1_DATAO_REG_10_ | ~new_P1_U6055;
  assign new_P1_U6089 = ~new_P1_U2385 | ~P1_LWORD_REG_11_;
  assign new_P1_U6090 = ~new_P1_U2384 | ~P1_EAX_REG_11_;
  assign new_P1_U6091 = ~P1_DATAO_REG_11_ | ~new_P1_U6055;
  assign new_P1_U6092 = ~new_P1_U2385 | ~P1_LWORD_REG_12_;
  assign new_P1_U6093 = ~new_P1_U2384 | ~P1_EAX_REG_12_;
  assign new_P1_U6094 = ~P1_DATAO_REG_12_ | ~new_P1_U6055;
  assign new_P1_U6095 = ~new_P1_U2385 | ~P1_LWORD_REG_13_;
  assign new_P1_U6096 = ~new_P1_U2384 | ~P1_EAX_REG_13_;
  assign new_P1_U6097 = ~P1_DATAO_REG_13_ | ~new_P1_U6055;
  assign new_P1_U6098 = ~new_P1_U2385 | ~P1_LWORD_REG_14_;
  assign new_P1_U6099 = ~new_P1_U2384 | ~P1_EAX_REG_14_;
  assign new_P1_U6100 = ~P1_DATAO_REG_14_ | ~new_P1_U6055;
  assign new_P1_U6101 = ~new_P1_U2385 | ~P1_LWORD_REG_15_;
  assign new_P1_U6102 = ~new_P1_U2384 | ~P1_EAX_REG_15_;
  assign new_P1_U6103 = ~P1_DATAO_REG_15_ | ~new_P1_U6055;
  assign new_P1_U6104 = ~new_P1_U2424 | ~P1_EAX_REG_16_;
  assign new_P1_U6105 = ~new_P1_U2385 | ~P1_UWORD_REG_0_;
  assign new_P1_U6106 = ~P1_DATAO_REG_16_ | ~new_P1_U6055;
  assign new_P1_U6107 = ~new_P1_U2424 | ~P1_EAX_REG_17_;
  assign new_P1_U6108 = ~new_P1_U2385 | ~P1_UWORD_REG_1_;
  assign new_P1_U6109 = ~P1_DATAO_REG_17_ | ~new_P1_U6055;
  assign new_P1_U6110 = ~new_P1_U2424 | ~P1_EAX_REG_18_;
  assign new_P1_U6111 = ~new_P1_U2385 | ~P1_UWORD_REG_2_;
  assign new_P1_U6112 = ~P1_DATAO_REG_18_ | ~new_P1_U6055;
  assign new_P1_U6113 = ~new_P1_U2424 | ~P1_EAX_REG_19_;
  assign new_P1_U6114 = ~new_P1_U2385 | ~P1_UWORD_REG_3_;
  assign new_P1_U6115 = ~P1_DATAO_REG_19_ | ~new_P1_U6055;
  assign new_P1_U6116 = ~new_P1_U2424 | ~P1_EAX_REG_20_;
  assign new_P1_U6117 = ~new_P1_U2385 | ~P1_UWORD_REG_4_;
  assign new_P1_U6118 = ~P1_DATAO_REG_20_ | ~new_P1_U6055;
  assign new_P1_U6119 = ~new_P1_U2424 | ~P1_EAX_REG_21_;
  assign new_P1_U6120 = ~new_P1_U2385 | ~P1_UWORD_REG_5_;
  assign new_P1_U6121 = ~P1_DATAO_REG_21_ | ~new_P1_U6055;
  assign new_P1_U6122 = ~new_P1_U2424 | ~P1_EAX_REG_22_;
  assign new_P1_U6123 = ~new_P1_U2385 | ~P1_UWORD_REG_6_;
  assign new_P1_U6124 = ~P1_DATAO_REG_22_ | ~new_P1_U6055;
  assign new_P1_U6125 = ~new_P1_U2424 | ~P1_EAX_REG_23_;
  assign new_P1_U6126 = ~new_P1_U2385 | ~P1_UWORD_REG_7_;
  assign new_P1_U6127 = ~P1_DATAO_REG_23_ | ~new_P1_U6055;
  assign new_P1_U6128 = ~new_P1_U2424 | ~P1_EAX_REG_24_;
  assign new_P1_U6129 = ~new_P1_U2385 | ~P1_UWORD_REG_8_;
  assign new_P1_U6130 = ~P1_DATAO_REG_24_ | ~new_P1_U6055;
  assign new_P1_U6131 = ~new_P1_U2424 | ~P1_EAX_REG_25_;
  assign new_P1_U6132 = ~new_P1_U2385 | ~P1_UWORD_REG_9_;
  assign new_P1_U6133 = ~P1_DATAO_REG_25_ | ~new_P1_U6055;
  assign new_P1_U6134 = ~new_P1_U2424 | ~P1_EAX_REG_26_;
  assign new_P1_U6135 = ~new_P1_U2385 | ~P1_UWORD_REG_10_;
  assign new_P1_U6136 = ~P1_DATAO_REG_26_ | ~new_P1_U6055;
  assign new_P1_U6137 = ~new_P1_U2424 | ~P1_EAX_REG_27_;
  assign new_P1_U6138 = ~new_P1_U2385 | ~P1_UWORD_REG_11_;
  assign new_P1_U6139 = ~P1_DATAO_REG_27_ | ~new_P1_U6055;
  assign new_P1_U6140 = ~new_P1_U2424 | ~P1_EAX_REG_28_;
  assign new_P1_U6141 = ~new_P1_U2385 | ~P1_UWORD_REG_12_;
  assign new_P1_U6142 = ~P1_DATAO_REG_28_ | ~new_P1_U6055;
  assign new_P1_U6143 = ~new_P1_U2424 | ~P1_EAX_REG_29_;
  assign new_P1_U6144 = ~new_P1_U2385 | ~P1_UWORD_REG_13_;
  assign new_P1_U6145 = ~P1_DATAO_REG_29_ | ~new_P1_U6055;
  assign new_P1_U6146 = ~new_P1_U2424 | ~P1_EAX_REG_30_;
  assign new_P1_U6147 = ~new_P1_U2385 | ~P1_UWORD_REG_14_;
  assign new_P1_U6148 = ~P1_DATAO_REG_30_ | ~new_P1_U6055;
  assign new_P1_U6149 = ~new_P1_GTE_485_U6 | ~new_P1_U4194 | ~new_P1_U2447;
  assign new_P1_U6150 = ~new_P1_U4194 | ~new_P1_U4254 | ~new_P1_U4197;
  assign new_P1_U6151 = ~new_P1_R2167_U17 | ~new_P1_U4200 | ~new_P1_U3283;
  assign new_P1_U6152 = ~new_P1_U7503 | ~new_P1_U3257;
  assign new_P1_U6153 = ~new_P1_U3883 | ~new_P1_U6152;
  assign new_P1_U6154 = ~new_P1_U2422 | ~new_U346;
  assign new_P1_U6155 = ~new_P1_U2386 | ~new_P1_R2358_U76;
  assign new_P1_U6156 = ~P1_EAX_REG_0_ | ~new_P1_U3424;
  assign new_P1_U6157 = ~new_P1_U2422 | ~new_U335;
  assign new_P1_U6158 = ~new_P1_U2386 | ~new_P1_R2358_U107;
  assign new_P1_U6159 = ~P1_EAX_REG_1_ | ~new_P1_U3424;
  assign new_P1_U6160 = ~new_P1_U2422 | ~new_U324;
  assign new_P1_U6161 = ~new_P1_U2386 | ~new_P1_R2358_U18;
  assign new_P1_U6162 = ~P1_EAX_REG_2_ | ~new_P1_U3424;
  assign new_P1_U6163 = ~new_P1_U2422 | ~new_U321;
  assign new_P1_U6164 = ~new_P1_U2386 | ~new_P1_R2358_U19;
  assign new_P1_U6165 = ~P1_EAX_REG_3_ | ~new_P1_U3424;
  assign new_P1_U6166 = ~new_P1_U2422 | ~new_U320;
  assign new_P1_U6167 = ~new_P1_U2386 | ~new_P1_R2358_U84;
  assign new_P1_U6168 = ~P1_EAX_REG_4_ | ~new_P1_U3424;
  assign new_P1_U6169 = ~new_P1_U2422 | ~new_U319;
  assign new_P1_U6170 = ~new_P1_U2386 | ~new_P1_R2358_U82;
  assign new_P1_U6171 = ~P1_EAX_REG_5_ | ~new_P1_U3424;
  assign new_P1_U6172 = ~new_P1_U2422 | ~new_U318;
  assign new_P1_U6173 = ~new_P1_U2386 | ~new_P1_R2358_U20;
  assign new_P1_U6174 = ~P1_EAX_REG_6_ | ~new_P1_U3424;
  assign new_P1_U6175 = ~new_P1_U2422 | ~new_U317;
  assign new_P1_U6176 = ~new_P1_U2386 | ~new_P1_R2358_U21;
  assign new_P1_U6177 = ~P1_EAX_REG_7_ | ~new_P1_U3424;
  assign new_P1_U6178 = ~new_P1_U2422 | ~new_U316;
  assign new_P1_U6179 = ~new_P1_U2386 | ~new_P1_R2358_U80;
  assign new_P1_U6180 = ~P1_EAX_REG_8_ | ~new_P1_U3424;
  assign new_P1_U6181 = ~new_P1_U2422 | ~new_U315;
  assign new_P1_U6182 = ~new_P1_U2386 | ~new_P1_R2358_U78;
  assign new_P1_U6183 = ~P1_EAX_REG_9_ | ~new_P1_U3424;
  assign new_P1_U6184 = ~new_P1_U2422 | ~new_U345;
  assign new_P1_U6185 = ~new_P1_U2386 | ~new_P1_R2358_U14;
  assign new_P1_U6186 = ~P1_EAX_REG_10_ | ~new_P1_U3424;
  assign new_P1_U6187 = ~new_P1_U2422 | ~new_U344;
  assign new_P1_U6188 = ~new_P1_U2386 | ~new_P1_R2358_U15;
  assign new_P1_U6189 = ~P1_EAX_REG_11_ | ~new_P1_U3424;
  assign new_P1_U6190 = ~new_P1_U2422 | ~new_U343;
  assign new_P1_U6191 = ~new_P1_U2386 | ~new_P1_R2358_U119;
  assign new_P1_U6192 = ~P1_EAX_REG_12_ | ~new_P1_U3424;
  assign new_P1_U6193 = ~new_P1_U2422 | ~new_U342;
  assign new_P1_U6194 = ~new_P1_U2386 | ~new_P1_R2358_U117;
  assign new_P1_U6195 = ~P1_EAX_REG_13_ | ~new_P1_U3424;
  assign new_P1_U6196 = ~new_P1_U2422 | ~new_U341;
  assign new_P1_U6197 = ~new_P1_U2386 | ~new_P1_R2358_U16;
  assign new_P1_U6198 = ~P1_EAX_REG_14_ | ~new_P1_U3424;
  assign new_P1_U6199 = ~new_P1_U2422 | ~new_U340;
  assign new_P1_U6200 = ~new_P1_U2386 | ~new_P1_R2358_U17;
  assign new_P1_U6201 = ~P1_EAX_REG_15_ | ~new_P1_U3424;
  assign new_P1_U6202 = ~new_P1_U2423 | ~new_U339;
  assign new_P1_U6203 = ~new_P1_U2387 | ~new_U346;
  assign new_P1_U6204 = ~new_P1_U2386 | ~new_P1_R2358_U115;
  assign new_P1_U6205 = ~P1_EAX_REG_16_ | ~new_P1_U3424;
  assign new_P1_U6206 = ~new_P1_U2423 | ~new_U338;
  assign new_P1_U6207 = ~new_P1_U2387 | ~new_U335;
  assign new_P1_U6208 = ~new_P1_U2386 | ~new_P1_R2358_U113;
  assign new_P1_U6209 = ~P1_EAX_REG_17_ | ~new_P1_U3424;
  assign new_P1_U6210 = ~new_P1_U2423 | ~new_U337;
  assign new_P1_U6211 = ~new_P1_U2387 | ~new_U324;
  assign new_P1_U6212 = ~new_P1_U2386 | ~new_P1_R2358_U111;
  assign new_P1_U6213 = ~P1_EAX_REG_18_ | ~new_P1_U3424;
  assign new_P1_U6214 = ~new_P1_U2423 | ~new_U336;
  assign new_P1_U6215 = ~new_P1_U2387 | ~new_U321;
  assign new_P1_U6216 = ~new_P1_U2386 | ~new_P1_R2358_U109;
  assign new_P1_U6217 = ~P1_EAX_REG_19_ | ~new_P1_U3424;
  assign new_P1_U6218 = ~new_P1_U2423 | ~new_U334;
  assign new_P1_U6219 = ~new_P1_U2387 | ~new_U320;
  assign new_P1_U6220 = ~new_P1_U2386 | ~new_P1_R2358_U105;
  assign new_P1_U6221 = ~P1_EAX_REG_20_ | ~new_P1_U3424;
  assign new_P1_U6222 = ~new_P1_U2423 | ~new_U333;
  assign new_P1_U6223 = ~new_P1_U2387 | ~new_U319;
  assign new_P1_U6224 = ~new_P1_U2386 | ~new_P1_R2358_U103;
  assign new_P1_U6225 = ~P1_EAX_REG_21_ | ~new_P1_U3424;
  assign new_P1_U6226 = ~new_P1_U2423 | ~new_U332;
  assign new_P1_U6227 = ~new_P1_U2387 | ~new_U318;
  assign new_P1_U6228 = ~new_P1_U2386 | ~new_P1_R2358_U101;
  assign new_P1_U6229 = ~P1_EAX_REG_22_ | ~new_P1_U3424;
  assign new_P1_U6230 = ~new_P1_U2423 | ~new_U331;
  assign new_P1_U6231 = ~new_P1_U2387 | ~new_U317;
  assign new_P1_U6232 = ~new_P1_U2386 | ~new_P1_R2358_U99;
  assign new_P1_U6233 = ~P1_EAX_REG_23_ | ~new_P1_U3424;
  assign new_P1_U6234 = ~new_P1_U2423 | ~new_U330;
  assign new_P1_U6235 = ~new_P1_U2387 | ~new_U316;
  assign new_P1_U6236 = ~new_P1_U2386 | ~new_P1_R2358_U97;
  assign new_P1_U6237 = ~P1_EAX_REG_24_ | ~new_P1_U3424;
  assign new_P1_U6238 = ~new_P1_U2423 | ~new_U329;
  assign new_P1_U6239 = ~new_P1_U2387 | ~new_U315;
  assign new_P1_U6240 = ~new_P1_U2386 | ~new_P1_R2358_U95;
  assign new_P1_U6241 = ~P1_EAX_REG_25_ | ~new_P1_U3424;
  assign new_P1_U6242 = ~new_P1_U2423 | ~new_U328;
  assign new_P1_U6243 = ~new_P1_U2387 | ~new_U345;
  assign new_P1_U6244 = ~new_P1_U2386 | ~new_P1_R2358_U93;
  assign new_P1_U6245 = ~P1_EAX_REG_26_ | ~new_P1_U3424;
  assign new_P1_U6246 = ~new_P1_U2423 | ~new_U327;
  assign new_P1_U6247 = ~new_P1_U2387 | ~new_U344;
  assign new_P1_U6248 = ~new_P1_U2386 | ~new_P1_R2358_U91;
  assign new_P1_U6249 = ~P1_EAX_REG_27_ | ~new_P1_U3424;
  assign new_P1_U6250 = ~new_P1_U2423 | ~new_U326;
  assign new_P1_U6251 = ~new_P1_U2387 | ~new_U343;
  assign new_P1_U6252 = ~new_P1_U2386 | ~new_P1_R2358_U89;
  assign new_P1_U6253 = ~P1_EAX_REG_28_ | ~new_P1_U3424;
  assign new_P1_U6254 = ~new_P1_U2423 | ~new_U325;
  assign new_P1_U6255 = ~new_P1_U2387 | ~new_U342;
  assign new_P1_U6256 = ~new_P1_U2386 | ~new_P1_R2358_U87;
  assign new_P1_U6257 = ~P1_EAX_REG_29_ | ~new_P1_U3424;
  assign new_P1_U6258 = ~new_P1_U2423 | ~new_U323;
  assign new_P1_U6259 = ~new_P1_U2387 | ~new_U341;
  assign new_P1_U6260 = ~new_P1_U2386 | ~new_P1_R2358_U85;
  assign new_P1_U6261 = ~P1_EAX_REG_30_ | ~new_P1_U3424;
  assign new_P1_U6262 = ~new_P1_U2423 | ~new_U322;
  assign new_P1_U6263 = ~new_P1_U4198 | ~new_P1_U3273;
  assign new_P1_U6264 = ~new_P1_U4205 | ~new_P1_U6263;
  assign new_P1_U6265 = ~new_P1_U2383 | ~new_P1_R2358_U76;
  assign new_P1_U6266 = ~new_P1_U2371 | ~new_P1_R2099_U86;
  assign new_P1_U6267 = ~P1_EBX_REG_0_ | ~new_P1_U3426;
  assign new_P1_U6268 = ~new_P1_U2383 | ~new_P1_R2358_U107;
  assign new_P1_U6269 = ~new_P1_U2371 | ~new_P1_R2099_U87;
  assign new_P1_U6270 = ~P1_EBX_REG_1_ | ~new_P1_U3426;
  assign new_P1_U6271 = ~new_P1_U2383 | ~new_P1_R2358_U18;
  assign new_P1_U6272 = ~new_P1_U2371 | ~new_P1_R2099_U138;
  assign new_P1_U6273 = ~P1_EBX_REG_2_ | ~new_P1_U3426;
  assign new_P1_U6274 = ~new_P1_U2383 | ~new_P1_R2358_U19;
  assign new_P1_U6275 = ~new_P1_U2371 | ~new_P1_R2099_U42;
  assign new_P1_U6276 = ~P1_EBX_REG_3_ | ~new_P1_U3426;
  assign new_P1_U6277 = ~new_P1_U2383 | ~new_P1_R2358_U84;
  assign new_P1_U6278 = ~new_P1_U2371 | ~new_P1_R2099_U41;
  assign new_P1_U6279 = ~P1_EBX_REG_4_ | ~new_P1_U3426;
  assign new_P1_U6280 = ~new_P1_U2383 | ~new_P1_R2358_U82;
  assign new_P1_U6281 = ~new_P1_U2371 | ~new_P1_R2099_U40;
  assign new_P1_U6282 = ~P1_EBX_REG_5_ | ~new_P1_U3426;
  assign new_P1_U6283 = ~new_P1_U2383 | ~new_P1_R2358_U20;
  assign new_P1_U6284 = ~new_P1_U2371 | ~new_P1_R2099_U39;
  assign new_P1_U6285 = ~P1_EBX_REG_6_ | ~new_P1_U3426;
  assign new_P1_U6286 = ~new_P1_U2383 | ~new_P1_R2358_U21;
  assign new_P1_U6287 = ~new_P1_U2371 | ~new_P1_R2099_U38;
  assign new_P1_U6288 = ~P1_EBX_REG_7_ | ~new_P1_U3426;
  assign new_P1_U6289 = ~new_P1_U2383 | ~new_P1_R2358_U80;
  assign new_P1_U6290 = ~new_P1_U2371 | ~new_P1_R2099_U37;
  assign new_P1_U6291 = ~P1_EBX_REG_8_ | ~new_P1_U3426;
  assign new_P1_U6292 = ~new_P1_U2383 | ~new_P1_R2358_U78;
  assign new_P1_U6293 = ~new_P1_U2371 | ~new_P1_R2099_U36;
  assign new_P1_U6294 = ~P1_EBX_REG_9_ | ~new_P1_U3426;
  assign new_P1_U6295 = ~new_P1_U2383 | ~new_P1_R2358_U14;
  assign new_P1_U6296 = ~new_P1_U2371 | ~new_P1_R2099_U85;
  assign new_P1_U6297 = ~P1_EBX_REG_10_ | ~new_P1_U3426;
  assign new_P1_U6298 = ~new_P1_U2383 | ~new_P1_R2358_U15;
  assign new_P1_U6299 = ~new_P1_U2371 | ~new_P1_R2099_U84;
  assign new_P1_U6300 = ~P1_EBX_REG_11_ | ~new_P1_U3426;
  assign new_P1_U6301 = ~new_P1_U2383 | ~new_P1_R2358_U119;
  assign new_P1_U6302 = ~new_P1_U2371 | ~new_P1_R2099_U83;
  assign new_P1_U6303 = ~P1_EBX_REG_12_ | ~new_P1_U3426;
  assign new_P1_U6304 = ~new_P1_U2383 | ~new_P1_R2358_U117;
  assign new_P1_U6305 = ~new_P1_U2371 | ~new_P1_R2099_U82;
  assign new_P1_U6306 = ~P1_EBX_REG_13_ | ~new_P1_U3426;
  assign new_P1_U6307 = ~new_P1_U2383 | ~new_P1_R2358_U16;
  assign new_P1_U6308 = ~new_P1_U2371 | ~new_P1_R2099_U81;
  assign new_P1_U6309 = ~P1_EBX_REG_14_ | ~new_P1_U3426;
  assign new_P1_U6310 = ~new_P1_U2383 | ~new_P1_R2358_U17;
  assign new_P1_U6311 = ~new_P1_U2371 | ~new_P1_R2099_U80;
  assign new_P1_U6312 = ~P1_EBX_REG_15_ | ~new_P1_U3426;
  assign new_P1_U6313 = ~new_P1_U2383 | ~new_P1_R2358_U115;
  assign new_P1_U6314 = ~new_P1_U2371 | ~new_P1_R2099_U79;
  assign new_P1_U6315 = ~P1_EBX_REG_16_ | ~new_P1_U3426;
  assign new_P1_U6316 = ~new_P1_U2383 | ~new_P1_R2358_U113;
  assign new_P1_U6317 = ~new_P1_U2371 | ~new_P1_R2099_U78;
  assign new_P1_U6318 = ~P1_EBX_REG_17_ | ~new_P1_U3426;
  assign new_P1_U6319 = ~new_P1_U2383 | ~new_P1_R2358_U111;
  assign new_P1_U6320 = ~new_P1_U2371 | ~new_P1_R2099_U77;
  assign new_P1_U6321 = ~P1_EBX_REG_18_ | ~new_P1_U3426;
  assign new_P1_U6322 = ~new_P1_U2383 | ~new_P1_R2358_U109;
  assign new_P1_U6323 = ~new_P1_U2371 | ~new_P1_R2099_U76;
  assign new_P1_U6324 = ~P1_EBX_REG_19_ | ~new_P1_U3426;
  assign new_P1_U6325 = ~new_P1_U2383 | ~new_P1_R2358_U105;
  assign new_P1_U6326 = ~new_P1_U2371 | ~new_P1_R2099_U75;
  assign new_P1_U6327 = ~P1_EBX_REG_20_ | ~new_P1_U3426;
  assign new_P1_U6328 = ~new_P1_U2383 | ~new_P1_R2358_U103;
  assign new_P1_U6329 = ~new_P1_U2371 | ~new_P1_R2099_U74;
  assign new_P1_U6330 = ~P1_EBX_REG_21_ | ~new_P1_U3426;
  assign new_P1_U6331 = ~new_P1_U2383 | ~new_P1_R2358_U101;
  assign new_P1_U6332 = ~new_P1_U2371 | ~new_P1_R2099_U73;
  assign new_P1_U6333 = ~P1_EBX_REG_22_ | ~new_P1_U3426;
  assign new_P1_U6334 = ~new_P1_U2383 | ~new_P1_R2358_U99;
  assign new_P1_U6335 = ~new_P1_U2371 | ~new_P1_R2099_U72;
  assign new_P1_U6336 = ~P1_EBX_REG_23_ | ~new_P1_U3426;
  assign new_P1_U6337 = ~new_P1_U2383 | ~new_P1_R2358_U97;
  assign new_P1_U6338 = ~new_P1_U2371 | ~new_P1_R2099_U71;
  assign new_P1_U6339 = ~P1_EBX_REG_24_ | ~new_P1_U3426;
  assign new_P1_U6340 = ~new_P1_U2383 | ~new_P1_R2358_U95;
  assign new_P1_U6341 = ~new_P1_U2371 | ~new_P1_R2099_U70;
  assign new_P1_U6342 = ~P1_EBX_REG_25_ | ~new_P1_U3426;
  assign new_P1_U6343 = ~new_P1_U2383 | ~new_P1_R2358_U93;
  assign new_P1_U6344 = ~new_P1_U2371 | ~new_P1_R2099_U69;
  assign new_P1_U6345 = ~P1_EBX_REG_26_ | ~new_P1_U3426;
  assign new_P1_U6346 = ~new_P1_U2383 | ~new_P1_R2358_U91;
  assign new_P1_U6347 = ~new_P1_U2371 | ~new_P1_R2099_U68;
  assign new_P1_U6348 = ~P1_EBX_REG_27_ | ~new_P1_U3426;
  assign new_P1_U6349 = ~new_P1_U2383 | ~new_P1_R2358_U89;
  assign new_P1_U6350 = ~new_P1_U2371 | ~new_P1_R2099_U67;
  assign new_P1_U6351 = ~P1_EBX_REG_28_ | ~new_P1_U3426;
  assign new_P1_U6352 = ~new_P1_U2383 | ~new_P1_R2358_U87;
  assign new_P1_U6353 = ~new_P1_U2371 | ~new_P1_R2099_U66;
  assign new_P1_U6354 = ~P1_EBX_REG_29_ | ~new_P1_U3426;
  assign new_P1_U6355 = ~new_P1_U2383 | ~new_P1_R2358_U85;
  assign new_P1_U6356 = ~new_P1_U2371 | ~new_P1_R2099_U65;
  assign new_P1_U6357 = ~P1_EBX_REG_30_ | ~new_P1_U3426;
  assign new_P1_U6358 = ~new_P1_U2371 | ~new_P1_R2099_U64;
  assign new_P1_U6359 = ~P1_EBX_REG_31_ | ~new_P1_U3426;
  assign new_P1_U6360 = ~new_P1_U4204 | ~new_P1_GTE_485_U6;
  assign new_P1_U6361 = ~new_P1_U4202 | ~new_P1_R2167_U17;
  assign new_P1_U6362 = ~new_P1_U4203 | ~new_P1_U3263;
  assign new_P1_U6363 = ~new_P1_U3431;
  assign new_P1_U6364 = ~new_P1_U4249 | ~P1_STATE2_REG_2_;
  assign new_P1_U6365 = ~new_P1_R2337_U69 | ~P1_STATE2_REG_1_;
  assign new_P1_U6366 = ~new_P1_U6365 | ~new_P1_U6364;
  assign new_P1_U6367 = P1_STATEBS16_REG | new_U210;
  assign new_P1_U6368 = ~new_P1_U2604 | ~new_P1_R2099_U86;
  assign new_P1_U6369 = ~P1_REIP_REG_0_ | ~new_P1_U7485;
  assign new_P1_U6370 = ~P1_EBX_REG_0_ | ~new_P1_U7484;
  assign new_P1_U6371 = ~new_P1_U2429 | ~new_P1_R2358_U76;
  assign new_P1_U6372 = ~new_P1_U2426 | ~new_P1_R2182_U34;
  assign new_P1_U6373 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_0_;
  assign new_P1_U6374 = ~new_P1_U2366 | ~P1_PHYADDRPOINTER_REG_0_;
  assign new_P1_U6375 = ~new_P1_U6363 | ~P1_REIP_REG_0_;
  assign new_P1_U6376 = ~new_P1_U2604 | ~new_P1_R2099_U87;
  assign new_P1_U6377 = ~new_P1_R2096_U4 | ~new_P1_U7485;
  assign new_P1_U6378 = ~P1_EBX_REG_1_ | ~new_P1_U7484;
  assign new_P1_U6379 = ~new_P1_U2429 | ~new_P1_R2358_U107;
  assign new_P1_U6380 = ~new_P1_U2426 | ~new_P1_R2182_U33;
  assign new_P1_U6381 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_1_;
  assign new_P1_U6382 = ~new_P1_U2366 | ~new_P1_R2337_U4;
  assign new_P1_U6383 = ~new_P1_U6363 | ~P1_REIP_REG_1_;
  assign new_P1_U6384 = ~new_P1_U2604 | ~new_P1_R2099_U138;
  assign new_P1_U6385 = ~new_P1_R2096_U71 | ~new_P1_U7485;
  assign new_P1_U6386 = ~P1_EBX_REG_2_ | ~new_P1_U7484;
  assign new_P1_U6387 = ~new_P1_U2429 | ~new_P1_R2358_U18;
  assign new_P1_U6388 = ~new_P1_U2426 | ~new_P1_R2182_U42;
  assign new_P1_U6389 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_2_;
  assign new_P1_U6390 = ~new_P1_U2366 | ~new_P1_R2337_U71;
  assign new_P1_U6391 = ~new_P1_U6363 | ~P1_REIP_REG_2_;
  assign new_P1_U6392 = ~new_P1_U2604 | ~new_P1_R2099_U42;
  assign new_P1_U6393 = ~new_P1_R2096_U68 | ~new_P1_U7485;
  assign new_P1_U6394 = ~P1_EBX_REG_3_ | ~new_P1_U7484;
  assign new_P1_U6395 = ~new_P1_U2429 | ~new_P1_R2358_U19;
  assign new_P1_U6396 = ~new_P1_U2426 | ~new_P1_R2182_U25;
  assign new_P1_U6397 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_3_;
  assign new_P1_U6398 = ~new_P1_U2366 | ~new_P1_R2337_U68;
  assign new_P1_U6399 = ~new_P1_U6363 | ~P1_REIP_REG_3_;
  assign new_P1_U6400 = ~new_P1_U2604 | ~new_P1_R2099_U41;
  assign new_P1_U6401 = ~new_P1_R2096_U67 | ~new_P1_U7485;
  assign new_P1_U6402 = ~P1_EBX_REG_4_ | ~new_P1_U7484;
  assign new_P1_U6403 = ~new_P1_U2429 | ~new_P1_R2358_U84;
  assign new_P1_U6404 = ~new_P1_U2426 | ~new_P1_R2182_U24;
  assign new_P1_U6405 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_4_;
  assign new_P1_U6406 = ~new_P1_U2366 | ~new_P1_R2337_U67;
  assign new_P1_U6407 = ~new_P1_U6363 | ~P1_REIP_REG_4_;
  assign new_P1_U6408 = ~new_P1_U2604 | ~new_P1_R2099_U40;
  assign new_P1_U6409 = ~new_P1_R2096_U66 | ~new_P1_U7485;
  assign new_P1_U6410 = ~P1_EBX_REG_5_ | ~new_P1_U7484;
  assign new_P1_U6411 = ~new_P1_U2429 | ~new_P1_R2358_U82;
  assign new_P1_U6412 = ~new_P1_R2182_U5 | ~new_P1_U2426;
  assign new_P1_U6413 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_5_;
  assign new_P1_U6414 = ~new_P1_U2366 | ~new_P1_R2337_U66;
  assign new_P1_U6415 = ~new_P1_U6363 | ~P1_REIP_REG_5_;
  assign new_P1_U6416 = ~new_P1_U2604 | ~new_P1_R2099_U39;
  assign new_P1_U6417 = ~new_P1_R2096_U65 | ~new_P1_U7485;
  assign new_P1_U6418 = ~P1_EBX_REG_6_ | ~new_P1_U7484;
  assign new_P1_U6419 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_6_;
  assign new_P1_U6420 = ~new_P1_U2367 | ~new_P1_R2358_U20;
  assign new_P1_U6421 = ~new_P1_U2366 | ~new_P1_R2337_U65;
  assign new_P1_U6422 = ~new_P1_U6363 | ~P1_REIP_REG_6_;
  assign new_P1_U6423 = ~new_P1_U2604 | ~new_P1_R2099_U38;
  assign new_P1_U6424 = ~new_P1_R2096_U64 | ~new_P1_U7485;
  assign new_P1_U6425 = ~P1_EBX_REG_7_ | ~new_P1_U7484;
  assign new_P1_U6426 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_7_;
  assign new_P1_U6427 = ~new_P1_U2367 | ~new_P1_R2358_U21;
  assign new_P1_U6428 = ~new_P1_U2366 | ~new_P1_R2337_U64;
  assign new_P1_U6429 = ~new_P1_U6363 | ~P1_REIP_REG_7_;
  assign new_P1_U6430 = ~new_P1_U2604 | ~new_P1_R2099_U37;
  assign new_P1_U6431 = ~new_P1_R2096_U63 | ~new_P1_U7485;
  assign new_P1_U6432 = ~P1_EBX_REG_8_ | ~new_P1_U7484;
  assign new_P1_U6433 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_8_;
  assign new_P1_U6434 = ~new_P1_U2367 | ~new_P1_R2358_U80;
  assign new_P1_U6435 = ~new_P1_U2366 | ~new_P1_R2337_U63;
  assign new_P1_U6436 = ~new_P1_U6363 | ~P1_REIP_REG_8_;
  assign new_P1_U6437 = ~new_P1_U2604 | ~new_P1_R2099_U36;
  assign new_P1_U6438 = ~new_P1_R2096_U62 | ~new_P1_U7485;
  assign new_P1_U6439 = ~P1_EBX_REG_9_ | ~new_P1_U7484;
  assign new_P1_U6440 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_9_;
  assign new_P1_U6441 = ~new_P1_U2367 | ~new_P1_R2358_U78;
  assign new_P1_U6442 = ~new_P1_U2366 | ~new_P1_R2337_U62;
  assign new_P1_U6443 = ~new_P1_U6363 | ~P1_REIP_REG_9_;
  assign new_P1_U6444 = ~new_P1_U2604 | ~new_P1_R2099_U85;
  assign new_P1_U6445 = ~new_P1_R2096_U91 | ~new_P1_U7485;
  assign new_P1_U6446 = ~P1_EBX_REG_10_ | ~new_P1_U7484;
  assign new_P1_U6447 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_10_;
  assign new_P1_U6448 = ~new_P1_U2367 | ~new_P1_R2358_U14;
  assign new_P1_U6449 = ~new_P1_U2366 | ~new_P1_R2337_U91;
  assign new_P1_U6450 = ~new_P1_U6363 | ~P1_REIP_REG_10_;
  assign new_P1_U6451 = ~new_P1_U2604 | ~new_P1_R2099_U84;
  assign new_P1_U6452 = ~new_P1_R2096_U90 | ~new_P1_U7485;
  assign new_P1_U6453 = ~P1_EBX_REG_11_ | ~new_P1_U7484;
  assign new_P1_U6454 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_11_;
  assign new_P1_U6455 = ~new_P1_U2367 | ~new_P1_R2358_U15;
  assign new_P1_U6456 = ~new_P1_U2366 | ~new_P1_R2337_U90;
  assign new_P1_U6457 = ~new_P1_U6363 | ~P1_REIP_REG_11_;
  assign new_P1_U6458 = ~new_P1_U2604 | ~new_P1_R2099_U83;
  assign new_P1_U6459 = ~new_P1_R2096_U89 | ~new_P1_U7485;
  assign new_P1_U6460 = ~P1_EBX_REG_12_ | ~new_P1_U7484;
  assign new_P1_U6461 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_12_;
  assign new_P1_U6462 = ~new_P1_U2367 | ~new_P1_R2358_U119;
  assign new_P1_U6463 = ~new_P1_U2366 | ~new_P1_R2337_U89;
  assign new_P1_U6464 = ~new_P1_U6363 | ~P1_REIP_REG_12_;
  assign new_P1_U6465 = ~new_P1_U2604 | ~new_P1_R2099_U82;
  assign new_P1_U6466 = ~new_P1_R2096_U88 | ~new_P1_U7485;
  assign new_P1_U6467 = ~P1_EBX_REG_13_ | ~new_P1_U7484;
  assign new_P1_U6468 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_13_;
  assign new_P1_U6469 = ~new_P1_U2367 | ~new_P1_R2358_U117;
  assign new_P1_U6470 = ~new_P1_U2366 | ~new_P1_R2337_U88;
  assign new_P1_U6471 = ~new_P1_U6363 | ~P1_REIP_REG_13_;
  assign new_P1_U6472 = ~new_P1_U2604 | ~new_P1_R2099_U81;
  assign new_P1_U6473 = ~new_P1_R2096_U87 | ~new_P1_U7485;
  assign new_P1_U6474 = ~P1_EBX_REG_14_ | ~new_P1_U7484;
  assign new_P1_U6475 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_14_;
  assign new_P1_U6476 = ~new_P1_U2367 | ~new_P1_R2358_U16;
  assign new_P1_U6477 = ~new_P1_U2366 | ~new_P1_R2337_U87;
  assign new_P1_U6478 = ~new_P1_U6363 | ~P1_REIP_REG_14_;
  assign new_P1_U6479 = ~new_P1_U2604 | ~new_P1_R2099_U80;
  assign new_P1_U6480 = ~new_P1_R2096_U86 | ~new_P1_U7485;
  assign new_P1_U6481 = ~P1_EBX_REG_15_ | ~new_P1_U7484;
  assign new_P1_U6482 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_15_;
  assign new_P1_U6483 = ~new_P1_U2367 | ~new_P1_R2358_U17;
  assign new_P1_U6484 = ~new_P1_U2366 | ~new_P1_R2337_U86;
  assign new_P1_U6485 = ~new_P1_U6363 | ~P1_REIP_REG_15_;
  assign new_P1_U6486 = ~new_P1_U2604 | ~new_P1_R2099_U79;
  assign new_P1_U6487 = ~new_P1_R2096_U85 | ~new_P1_U7485;
  assign new_P1_U6488 = ~P1_EBX_REG_16_ | ~new_P1_U7484;
  assign new_P1_U6489 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_16_;
  assign new_P1_U6490 = ~new_P1_U2367 | ~new_P1_R2358_U115;
  assign new_P1_U6491 = ~new_P1_U2366 | ~new_P1_R2337_U85;
  assign new_P1_U6492 = ~new_P1_U6363 | ~P1_REIP_REG_16_;
  assign new_P1_U6493 = ~new_P1_U2604 | ~new_P1_R2099_U78;
  assign new_P1_U6494 = ~new_P1_R2096_U84 | ~new_P1_U7485;
  assign new_P1_U6495 = ~P1_EBX_REG_17_ | ~new_P1_U7484;
  assign new_P1_U6496 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_17_;
  assign new_P1_U6497 = ~new_P1_U2367 | ~new_P1_R2358_U113;
  assign new_P1_U6498 = ~new_P1_U2366 | ~new_P1_R2337_U84;
  assign new_P1_U6499 = ~new_P1_U6363 | ~P1_REIP_REG_17_;
  assign new_P1_U6500 = ~new_P1_U2604 | ~new_P1_R2099_U77;
  assign new_P1_U6501 = ~new_P1_R2096_U83 | ~new_P1_U7485;
  assign new_P1_U6502 = ~P1_EBX_REG_18_ | ~new_P1_U7484;
  assign new_P1_U6503 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_18_;
  assign new_P1_U6504 = ~new_P1_U2367 | ~new_P1_R2358_U111;
  assign new_P1_U6505 = ~new_P1_U2366 | ~new_P1_R2337_U83;
  assign new_P1_U6506 = ~new_P1_U6363 | ~P1_REIP_REG_18_;
  assign new_P1_U6507 = ~new_P1_U2604 | ~new_P1_R2099_U76;
  assign new_P1_U6508 = ~new_P1_R2096_U82 | ~new_P1_U7485;
  assign new_P1_U6509 = ~P1_EBX_REG_19_ | ~new_P1_U7484;
  assign new_P1_U6510 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_19_;
  assign new_P1_U6511 = ~new_P1_U2367 | ~new_P1_R2358_U109;
  assign new_P1_U6512 = ~new_P1_U2366 | ~new_P1_R2337_U82;
  assign new_P1_U6513 = ~new_P1_U6363 | ~P1_REIP_REG_19_;
  assign new_P1_U6514 = ~new_P1_U2604 | ~new_P1_R2099_U75;
  assign new_P1_U6515 = ~new_P1_R2096_U81 | ~new_P1_U7485;
  assign new_P1_U6516 = ~P1_EBX_REG_20_ | ~new_P1_U7484;
  assign new_P1_U6517 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_20_;
  assign new_P1_U6518 = ~new_P1_U2367 | ~new_P1_R2358_U105;
  assign new_P1_U6519 = ~new_P1_U2366 | ~new_P1_R2337_U81;
  assign new_P1_U6520 = ~new_P1_U6363 | ~P1_REIP_REG_20_;
  assign new_P1_U6521 = ~new_P1_U2604 | ~new_P1_R2099_U74;
  assign new_P1_U6522 = ~new_P1_R2096_U80 | ~new_P1_U7485;
  assign new_P1_U6523 = ~P1_EBX_REG_21_ | ~new_P1_U7484;
  assign new_P1_U6524 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_21_;
  assign new_P1_U6525 = ~new_P1_U2367 | ~new_P1_R2358_U103;
  assign new_P1_U6526 = ~new_P1_U2366 | ~new_P1_R2337_U80;
  assign new_P1_U6527 = ~new_P1_U6363 | ~P1_REIP_REG_21_;
  assign new_P1_U6528 = ~new_P1_U2604 | ~new_P1_R2099_U73;
  assign new_P1_U6529 = ~new_P1_R2096_U79 | ~new_P1_U7485;
  assign new_P1_U6530 = ~P1_EBX_REG_22_ | ~new_P1_U7484;
  assign new_P1_U6531 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_22_;
  assign new_P1_U6532 = ~new_P1_U2367 | ~new_P1_R2358_U101;
  assign new_P1_U6533 = ~new_P1_U2366 | ~new_P1_R2337_U79;
  assign new_P1_U6534 = ~new_P1_U6363 | ~P1_REIP_REG_22_;
  assign new_P1_U6535 = ~new_P1_U2604 | ~new_P1_R2099_U72;
  assign new_P1_U6536 = ~new_P1_R2096_U78 | ~new_P1_U7485;
  assign new_P1_U6537 = ~P1_EBX_REG_23_ | ~new_P1_U7484;
  assign new_P1_U6538 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_23_;
  assign new_P1_U6539 = ~new_P1_U2367 | ~new_P1_R2358_U99;
  assign new_P1_U6540 = ~new_P1_U2366 | ~new_P1_R2337_U78;
  assign new_P1_U6541 = ~new_P1_U6363 | ~P1_REIP_REG_23_;
  assign new_P1_U6542 = ~new_P1_U2604 | ~new_P1_R2099_U71;
  assign new_P1_U6543 = ~new_P1_R2096_U77 | ~new_P1_U7485;
  assign new_P1_U6544 = ~P1_EBX_REG_24_ | ~new_P1_U7484;
  assign new_P1_U6545 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_24_;
  assign new_P1_U6546 = ~new_P1_U2367 | ~new_P1_R2358_U97;
  assign new_P1_U6547 = ~new_P1_U2366 | ~new_P1_R2337_U77;
  assign new_P1_U6548 = ~new_P1_U6363 | ~P1_REIP_REG_24_;
  assign new_P1_U6549 = ~new_P1_U2604 | ~new_P1_R2099_U70;
  assign new_P1_U6550 = ~new_P1_R2096_U76 | ~new_P1_U7485;
  assign new_P1_U6551 = ~P1_EBX_REG_25_ | ~new_P1_U7484;
  assign new_P1_U6552 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_25_;
  assign new_P1_U6553 = ~new_P1_U2367 | ~new_P1_R2358_U95;
  assign new_P1_U6554 = ~new_P1_U2366 | ~new_P1_R2337_U76;
  assign new_P1_U6555 = ~new_P1_U6363 | ~P1_REIP_REG_25_;
  assign new_P1_U6556 = ~new_P1_U2604 | ~new_P1_R2099_U69;
  assign new_P1_U6557 = ~new_P1_R2096_U75 | ~new_P1_U7485;
  assign new_P1_U6558 = ~P1_EBX_REG_26_ | ~new_P1_U7484;
  assign new_P1_U6559 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_26_;
  assign new_P1_U6560 = ~new_P1_U2367 | ~new_P1_R2358_U93;
  assign new_P1_U6561 = ~new_P1_U2366 | ~new_P1_R2337_U75;
  assign new_P1_U6562 = ~new_P1_U6363 | ~P1_REIP_REG_26_;
  assign new_P1_U6563 = ~new_P1_U2604 | ~new_P1_R2099_U68;
  assign new_P1_U6564 = ~new_P1_R2096_U74 | ~new_P1_U7485;
  assign new_P1_U6565 = ~P1_EBX_REG_27_ | ~new_P1_U7484;
  assign new_P1_U6566 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_27_;
  assign new_P1_U6567 = ~new_P1_U2367 | ~new_P1_R2358_U91;
  assign new_P1_U6568 = ~new_P1_U2366 | ~new_P1_R2337_U74;
  assign new_P1_U6569 = ~new_P1_U6363 | ~P1_REIP_REG_27_;
  assign new_P1_U6570 = ~new_P1_U2604 | ~new_P1_R2099_U67;
  assign new_P1_U6571 = ~new_P1_R2096_U73 | ~new_P1_U7485;
  assign new_P1_U6572 = ~P1_EBX_REG_28_ | ~new_P1_U7484;
  assign new_P1_U6573 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_28_;
  assign new_P1_U6574 = ~new_P1_U2367 | ~new_P1_R2358_U89;
  assign new_P1_U6575 = ~new_P1_U2366 | ~new_P1_R2337_U73;
  assign new_P1_U6576 = ~new_P1_U6363 | ~P1_REIP_REG_28_;
  assign new_P1_U6577 = ~new_P1_U2604 | ~new_P1_R2099_U66;
  assign new_P1_U6578 = ~new_P1_R2096_U72 | ~new_P1_U7485;
  assign new_P1_U6579 = ~P1_EBX_REG_29_ | ~new_P1_U7484;
  assign new_P1_U6580 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_29_;
  assign new_P1_U6581 = ~new_P1_U2367 | ~new_P1_R2358_U87;
  assign new_P1_U6582 = ~new_P1_U2366 | ~new_P1_R2337_U72;
  assign new_P1_U6583 = ~new_P1_U6363 | ~P1_REIP_REG_29_;
  assign new_P1_U6584 = ~new_P1_U2604 | ~new_P1_R2099_U65;
  assign new_P1_U6585 = ~new_P1_R2096_U70 | ~new_P1_U7485;
  assign new_P1_U6586 = ~P1_EBX_REG_30_ | ~new_P1_U7484;
  assign new_P1_U6587 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_30_;
  assign new_P1_U6588 = ~new_P1_U2367 | ~new_P1_R2358_U85;
  assign new_P1_U6589 = ~new_P1_U2366 | ~new_P1_R2337_U70;
  assign new_P1_U6590 = ~new_P1_U6363 | ~P1_REIP_REG_30_;
  assign new_P1_U6591 = ~new_P1_U2604 | ~new_P1_R2099_U64;
  assign new_P1_U6592 = ~new_P1_R2096_U69 | ~new_P1_U7485;
  assign new_P1_U6593 = ~P1_EBX_REG_31_ | ~new_P1_U7484;
  assign new_P1_U6594 = ~new_P1_U2373 | ~P1_PHYADDRPOINTER_REG_31_;
  assign new_P1_U6595 = ~new_P1_U2367 | ~new_P1_R2358_U22;
  assign new_P1_U6596 = ~new_P1_U2366 | ~new_P1_R2337_U69;
  assign new_P1_U6597 = ~new_P1_U6363 | ~P1_REIP_REG_31_;
  assign new_P1_U6598 = ~P1_DATAWIDTH_REG_1_ | ~P1_DATAWIDTH_REG_0_;
  assign new_P1_U6599 = P1_REIP_REG_1_ | P1_REIP_REG_0_;
  assign new_P1_U6600 = ~new_P1_U4177;
  assign new_P1_U6601 = ~P1_FLUSH_REG | ~new_P1_U4177;
  assign new_P1_U6602 = ~new_P1_U3966 | ~new_P1_U2428;
  assign new_P1_U6603 = ~new_P1_U4180;
  assign new_P1_U6604 = ~P1_STATEBS16_REG | ~new_P1_U4497;
  assign new_P1_U6605 = ~new_P1_U4208 | ~new_P1_U6604;
  assign new_P1_U6606 = ~new_P1_U3964 | ~new_P1_U6605;
  assign new_P1_U6607 = ~P1_STATE2_REG_0_ | ~new_P1_U6606;
  assign new_P1_U6608 = ~new_P1_U4193 | ~new_P1_U3272;
  assign new_P1_U6609 = ~new_P1_U3965 | ~new_P1_U6607;
  assign new_P1_U6610 = ~new_P1_U2368 | ~new_P1_U2473;
  assign new_P1_U6611 = ~P1_CODEFETCH_REG | ~new_P1_U6610;
  assign new_P1_U6612 = ~new_P1_U4255 | ~P1_STATE2_REG_0_;
  assign new_P1_U6613 = ~P1_ADS_N_REG | ~P1_STATE_REG_0_;
  assign new_P1_U6614 = ~new_P1_U4181;
  assign new_P1_U6615 = ~new_P1_U3968 | ~new_P1_U3291;
  assign new_P1_U6616 = ~new_P1_U3406 | ~new_P1_U4499 | ~new_P1_U3969;
  assign new_P1_U6617 = ~P1_MEMORYFETCH_REG | ~new_P1_U6616;
  assign new_P1_U6618 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__7_;
  assign new_P1_U6619 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__7_;
  assign new_P1_U6620 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__7_;
  assign new_P1_U6621 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__7_;
  assign new_P1_U6622 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__7_;
  assign new_P1_U6623 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__7_;
  assign new_P1_U6624 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__7_;
  assign new_P1_U6625 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__7_;
  assign new_P1_U6626 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__7_;
  assign new_P1_U6627 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__7_;
  assign new_P1_U6628 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__7_;
  assign new_P1_U6629 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__7_;
  assign new_P1_U6630 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__7_;
  assign new_P1_U6631 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__7_;
  assign new_P1_U6632 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__7_;
  assign new_P1_U6633 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__7_;
  assign new_P1_U6634 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__6_;
  assign new_P1_U6635 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__6_;
  assign new_P1_U6636 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__6_;
  assign new_P1_U6637 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__6_;
  assign new_P1_U6638 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__6_;
  assign new_P1_U6639 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__6_;
  assign new_P1_U6640 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__6_;
  assign new_P1_U6641 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__6_;
  assign new_P1_U6642 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__6_;
  assign new_P1_U6643 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__6_;
  assign new_P1_U6644 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__6_;
  assign new_P1_U6645 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__6_;
  assign new_P1_U6646 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__6_;
  assign new_P1_U6647 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__6_;
  assign new_P1_U6648 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__6_;
  assign new_P1_U6649 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__6_;
  assign new_P1_U6650 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__5_;
  assign new_P1_U6651 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__5_;
  assign new_P1_U6652 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__5_;
  assign new_P1_U6653 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__5_;
  assign new_P1_U6654 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__5_;
  assign new_P1_U6655 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__5_;
  assign new_P1_U6656 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__5_;
  assign new_P1_U6657 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__5_;
  assign new_P1_U6658 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__5_;
  assign new_P1_U6659 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__5_;
  assign new_P1_U6660 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__5_;
  assign new_P1_U6661 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__5_;
  assign new_P1_U6662 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__5_;
  assign new_P1_U6663 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__5_;
  assign new_P1_U6664 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__5_;
  assign new_P1_U6665 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__5_;
  assign new_P1_U6666 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__4_;
  assign new_P1_U6667 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__4_;
  assign new_P1_U6668 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__4_;
  assign new_P1_U6669 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__4_;
  assign new_P1_U6670 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__4_;
  assign new_P1_U6671 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__4_;
  assign new_P1_U6672 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__4_;
  assign new_P1_U6673 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__4_;
  assign new_P1_U6674 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__4_;
  assign new_P1_U6675 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__4_;
  assign new_P1_U6676 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__4_;
  assign new_P1_U6677 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__4_;
  assign new_P1_U6678 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__4_;
  assign new_P1_U6679 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__4_;
  assign new_P1_U6680 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__4_;
  assign new_P1_U6681 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__3_;
  assign new_P1_U6682 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__3_;
  assign new_P1_U6683 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__3_;
  assign new_P1_U6684 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__3_;
  assign new_P1_U6685 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__3_;
  assign new_P1_U6686 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__3_;
  assign new_P1_U6687 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__3_;
  assign new_P1_U6688 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__3_;
  assign new_P1_U6689 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__3_;
  assign new_P1_U6690 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__3_;
  assign new_P1_U6691 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__3_;
  assign new_P1_U6692 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__3_;
  assign new_P1_U6693 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__3_;
  assign new_P1_U6694 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__3_;
  assign new_P1_U6695 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__3_;
  assign new_P1_U6696 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__3_;
  assign new_P1_U6697 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__2_;
  assign new_P1_U6698 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__2_;
  assign new_P1_U6699 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__2_;
  assign new_P1_U6700 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__2_;
  assign new_P1_U6701 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__2_;
  assign new_P1_U6702 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__2_;
  assign new_P1_U6703 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__2_;
  assign new_P1_U6704 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__2_;
  assign new_P1_U6705 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__2_;
  assign new_P1_U6706 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__2_;
  assign new_P1_U6707 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__2_;
  assign new_P1_U6708 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__2_;
  assign new_P1_U6709 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__2_;
  assign new_P1_U6710 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__2_;
  assign new_P1_U6711 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__2_;
  assign new_P1_U6712 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__2_;
  assign new_P1_U6713 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__1_;
  assign new_P1_U6714 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__1_;
  assign new_P1_U6715 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__1_;
  assign new_P1_U6716 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__1_;
  assign new_P1_U6717 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__1_;
  assign new_P1_U6718 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__1_;
  assign new_P1_U6719 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__1_;
  assign new_P1_U6720 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__1_;
  assign new_P1_U6721 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__1_;
  assign new_P1_U6722 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__1_;
  assign new_P1_U6723 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__1_;
  assign new_P1_U6724 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__1_;
  assign new_P1_U6725 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__1_;
  assign new_P1_U6726 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__1_;
  assign new_P1_U6727 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__1_;
  assign new_P1_U6728 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__1_;
  assign new_P1_U6729 = ~new_P1_U2544 | ~P1_INSTQUEUE_REG_15__0_;
  assign new_P1_U6730 = ~new_P1_U2543 | ~P1_INSTQUEUE_REG_14__0_;
  assign new_P1_U6731 = ~new_P1_U2542 | ~P1_INSTQUEUE_REG_13__0_;
  assign new_P1_U6732 = ~new_P1_U2541 | ~P1_INSTQUEUE_REG_12__0_;
  assign new_P1_U6733 = ~new_P1_U2539 | ~P1_INSTQUEUE_REG_11__0_;
  assign new_P1_U6734 = ~new_P1_U2538 | ~P1_INSTQUEUE_REG_10__0_;
  assign new_P1_U6735 = ~new_P1_U2537 | ~P1_INSTQUEUE_REG_9__0_;
  assign new_P1_U6736 = ~new_P1_U2536 | ~P1_INSTQUEUE_REG_8__0_;
  assign new_P1_U6737 = ~new_P1_U2534 | ~P1_INSTQUEUE_REG_7__0_;
  assign new_P1_U6738 = ~new_P1_U2533 | ~P1_INSTQUEUE_REG_6__0_;
  assign new_P1_U6739 = ~new_P1_U2532 | ~P1_INSTQUEUE_REG_5__0_;
  assign new_P1_U6740 = ~new_P1_U2531 | ~P1_INSTQUEUE_REG_4__0_;
  assign new_P1_U6741 = ~new_P1_U2529 | ~P1_INSTQUEUE_REG_3__0_;
  assign new_P1_U6742 = ~new_P1_U2527 | ~P1_INSTQUEUE_REG_2__0_;
  assign new_P1_U6743 = ~new_P1_U2525 | ~P1_INSTQUEUE_REG_1__0_;
  assign new_P1_U6744 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__0_;
  assign new_P1_U6745 = ~new_P1_U4460 | ~P1_STATE2_REG_2_;
  assign new_P1_U6746 = ~new_P1_U3412 | ~new_P1_U6745;
  assign new_P1_U6747 = ~new_P1_U4188 | ~P1_EAX_REG_9_;
  assign new_P1_U6748 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_9_;
  assign new_P1_U6749 = ~new_P1_R2337_U62 | ~new_P1_U2352;
  assign new_P1_U6750 = ~new_P1_U4188 | ~P1_EAX_REG_8_;
  assign new_P1_U6751 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_8_;
  assign new_P1_U6752 = ~new_P1_R2337_U63 | ~new_P1_U2352;
  assign new_P1_U6753 = ~new_P1_U4188 | ~P1_EAX_REG_7_;
  assign new_P1_U6754 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_7_;
  assign new_P1_U6755 = ~new_P1_R2337_U64 | ~new_P1_U2352;
  assign new_P1_U6756 = ~new_P1_U4188 | ~P1_EAX_REG_6_;
  assign new_P1_U6757 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_6_;
  assign new_P1_U6758 = ~new_P1_R2337_U65 | ~new_P1_U2352;
  assign new_P1_U6759 = ~new_P1_R2182_U5 | ~new_P1_U6746;
  assign new_P1_U6760 = ~new_P1_U4188 | ~P1_EAX_REG_5_;
  assign new_P1_U6761 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_5_;
  assign new_P1_U6762 = ~new_P1_R2337_U66 | ~new_P1_U2352;
  assign new_P1_U6763 = ~new_P1_R2182_U24 | ~new_P1_U6746;
  assign new_P1_U6764 = ~new_P1_U4188 | ~P1_EAX_REG_4_;
  assign new_P1_U6765 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_4_;
  assign new_P1_U6766 = ~new_P1_R2337_U67 | ~new_P1_U2352;
  assign new_P1_U6767 = ~new_P1_U2353 | ~P1_INSTQUEUERD_ADDR_REG_4_;
  assign new_P1_U6768 = ~new_P1_U4188 | ~P1_EAX_REG_31_;
  assign new_P1_U6769 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_31_;
  assign new_P1_U6770 = ~new_P1_R2337_U69 | ~new_P1_U2352;
  assign new_P1_U6771 = ~new_P1_R2182_U26 | ~new_P1_U6746;
  assign new_P1_U6772 = ~new_P1_U4188 | ~P1_EAX_REG_30_;
  assign new_P1_U6773 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_30_;
  assign new_P1_U6774 = ~new_P1_R2337_U70 | ~new_P1_U2352;
  assign new_P1_U6775 = ~new_P1_R2182_U25 | ~new_P1_U6746;
  assign new_P1_U6776 = ~new_P1_U4188 | ~P1_EAX_REG_3_;
  assign new_P1_U6777 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_3_;
  assign new_P1_U6778 = ~new_P1_R2337_U68 | ~new_P1_U2352;
  assign new_P1_U6779 = ~new_P1_U2353 | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U6780 = ~new_P1_R2182_U27 | ~new_P1_U6746;
  assign new_P1_U6781 = ~new_P1_U4188 | ~P1_EAX_REG_29_;
  assign new_P1_U6782 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_29_;
  assign new_P1_U6783 = ~new_P1_R2337_U72 | ~new_P1_U2352;
  assign new_P1_U6784 = ~new_P1_R2182_U28 | ~new_P1_U6746;
  assign new_P1_U6785 = ~new_P1_U4188 | ~P1_EAX_REG_28_;
  assign new_P1_U6786 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_28_;
  assign new_P1_U6787 = ~new_P1_R2337_U73 | ~new_P1_U2352;
  assign new_P1_U6788 = ~new_P1_R2182_U29 | ~new_P1_U6746;
  assign new_P1_U6789 = ~new_P1_U4188 | ~P1_EAX_REG_27_;
  assign new_P1_U6790 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_27_;
  assign new_P1_U6791 = ~new_P1_R2337_U74 | ~new_P1_U2352;
  assign new_P1_U6792 = ~new_P1_R2182_U30 | ~new_P1_U6746;
  assign new_P1_U6793 = ~new_P1_U4188 | ~P1_EAX_REG_26_;
  assign new_P1_U6794 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_26_;
  assign new_P1_U6795 = ~new_P1_R2337_U75 | ~new_P1_U2352;
  assign new_P1_U6796 = ~new_P1_R2182_U31 | ~new_P1_U6746;
  assign new_P1_U6797 = ~new_P1_U4188 | ~P1_EAX_REG_25_;
  assign new_P1_U6798 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_25_;
  assign new_P1_U6799 = ~new_P1_R2337_U76 | ~new_P1_U2352;
  assign new_P1_U6800 = ~new_P1_R2182_U32 | ~new_P1_U6746;
  assign new_P1_U6801 = ~new_P1_U4188 | ~P1_EAX_REG_24_;
  assign new_P1_U6802 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_24_;
  assign new_P1_U6803 = ~new_P1_R2337_U77 | ~new_P1_U2352;
  assign new_P1_U6804 = ~new_P1_R2182_U6 | ~new_P1_U6746;
  assign new_P1_U6805 = ~new_P1_U4188 | ~P1_EAX_REG_23_;
  assign new_P1_U6806 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_23_;
  assign new_P1_U6807 = ~new_P1_R2337_U78 | ~new_P1_U2352;
  assign new_P1_U6808 = ~new_P1_U2724 | ~new_P1_U6746;
  assign new_P1_U6809 = ~new_P1_U4188 | ~P1_EAX_REG_22_;
  assign new_P1_U6810 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_22_;
  assign new_P1_U6811 = ~new_P1_R2337_U79 | ~new_P1_U2352;
  assign new_P1_U6812 = ~new_P1_U2725 | ~new_P1_U6746;
  assign new_P1_U6813 = ~new_P1_U4188 | ~P1_EAX_REG_21_;
  assign new_P1_U6814 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_21_;
  assign new_P1_U6815 = ~new_P1_R2337_U80 | ~new_P1_U2352;
  assign new_P1_U6816 = ~new_P1_U2726 | ~new_P1_U6746;
  assign new_P1_U6817 = ~new_P1_U4188 | ~P1_EAX_REG_20_;
  assign new_P1_U6818 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_20_;
  assign new_P1_U6819 = ~new_P1_R2337_U81 | ~new_P1_U2352;
  assign new_P1_U6820 = ~new_P1_R2182_U42 | ~new_P1_U6746;
  assign new_P1_U6821 = ~new_P1_U4188 | ~P1_EAX_REG_2_;
  assign new_P1_U6822 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_2_;
  assign new_P1_U6823 = ~new_P1_R2337_U71 | ~new_P1_U2352;
  assign new_P1_U6824 = ~new_P1_U2353 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U6825 = ~new_P1_U2727 | ~new_P1_U6746;
  assign new_P1_U6826 = ~new_P1_U4188 | ~P1_EAX_REG_19_;
  assign new_P1_U6827 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_19_;
  assign new_P1_U6828 = ~new_P1_R2337_U82 | ~new_P1_U2352;
  assign new_P1_U6829 = ~new_P1_U2728 | ~new_P1_U6746;
  assign new_P1_U6830 = ~new_P1_U4188 | ~P1_EAX_REG_18_;
  assign new_P1_U6831 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_18_;
  assign new_P1_U6832 = ~new_P1_R2337_U83 | ~new_P1_U2352;
  assign new_P1_U6833 = ~new_P1_U2729 | ~new_P1_U6746;
  assign new_P1_U6834 = ~new_P1_U4188 | ~P1_EAX_REG_17_;
  assign new_P1_U6835 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_17_;
  assign new_P1_U6836 = ~new_P1_R2337_U84 | ~new_P1_U2352;
  assign new_P1_U6837 = ~new_P1_U2730 | ~new_P1_U6746;
  assign new_P1_U6838 = ~new_P1_U4188 | ~P1_EAX_REG_16_;
  assign new_P1_U6839 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_16_;
  assign new_P1_U6840 = ~new_P1_R2337_U85 | ~new_P1_U2352;
  assign new_P1_U6841 = ~new_P1_U4188 | ~P1_EAX_REG_15_;
  assign new_P1_U6842 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_15_;
  assign new_P1_U6843 = ~new_P1_R2337_U86 | ~new_P1_U2352;
  assign new_P1_U6844 = ~new_P1_U4188 | ~P1_EAX_REG_14_;
  assign new_P1_U6845 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_14_;
  assign new_P1_U6846 = ~new_P1_R2337_U87 | ~new_P1_U2352;
  assign new_P1_U6847 = ~new_P1_U4188 | ~P1_EAX_REG_13_;
  assign new_P1_U6848 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_13_;
  assign new_P1_U6849 = ~new_P1_R2337_U88 | ~new_P1_U2352;
  assign new_P1_U6850 = ~new_P1_U4188 | ~P1_EAX_REG_12_;
  assign new_P1_U6851 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_12_;
  assign new_P1_U6852 = ~new_P1_R2337_U89 | ~new_P1_U2352;
  assign new_P1_U6853 = ~new_P1_U4188 | ~P1_EAX_REG_11_;
  assign new_P1_U6854 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_11_;
  assign new_P1_U6855 = ~new_P1_R2337_U90 | ~new_P1_U2352;
  assign new_P1_U6856 = ~new_P1_U4188 | ~P1_EAX_REG_10_;
  assign new_P1_U6857 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_10_;
  assign new_P1_U6858 = ~new_P1_R2337_U91 | ~new_P1_U2352;
  assign new_P1_U6859 = ~new_P1_R2182_U33 | ~new_P1_U6746;
  assign new_P1_U6860 = ~new_P1_U4188 | ~P1_EAX_REG_1_;
  assign new_P1_U6861 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_1_;
  assign new_P1_U6862 = ~new_P1_R2337_U4 | ~new_P1_U2352;
  assign new_P1_U6863 = ~new_P1_U2353 | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U6864 = ~new_P1_R2182_U34 | ~new_P1_U6746;
  assign new_P1_U6865 = ~new_P1_U4188 | ~P1_EAX_REG_0_;
  assign new_P1_U6866 = ~new_P1_U4187 | ~P1_PHYADDRPOINTER_REG_0_;
  assign new_P1_U6867 = ~P1_PHYADDRPOINTER_REG_0_ | ~new_P1_U2352;
  assign new_P1_U6868 = ~new_P1_U2353 | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U6869 = ~new_P1_R2144_U49 | ~new_P1_U6746;
  assign new_P1_U6870 = ~new_P1_U3309 | ~new_P1_U3439 | ~new_P1_U4460;
  assign new_P1_U6871 = ~new_P1_U4159 | ~new_P1_R2144_U80;
  assign new_P1_U6872 = ~new_P1_ADD_371_U6 | ~new_P1_U4208;
  assign new_P1_U6873 = ~new_P1_U4159 | ~new_P1_R2144_U10;
  assign new_P1_U6874 = ~new_P1_ADD_371_U21 | ~new_P1_U4208;
  assign new_P1_U6875 = ~new_P1_U4159 | ~new_P1_R2144_U9;
  assign new_P1_U6876 = ~new_P1_ADD_371_U17 | ~new_P1_U4208;
  assign new_P1_U6877 = ~new_P1_U4159 | ~new_P1_R2144_U45;
  assign new_P1_U6878 = ~new_P1_ADD_371_U19 | ~new_P1_U4208;
  assign new_P1_U6879 = ~new_P1_U4159 | ~new_P1_R2144_U47;
  assign new_P1_U6880 = ~new_P1_ADD_371_U18 | ~new_P1_U4208;
  assign new_P1_U6881 = ~new_P1_U4159 | ~new_P1_R2144_U8;
  assign new_P1_U6882 = ~new_P1_ADD_371_U24 | ~new_P1_U4208;
  assign new_P1_U6883 = ~new_P1_U4159 | ~new_P1_R2144_U49;
  assign new_P1_U6884 = ~new_P1_ADD_371_U5 | ~new_P1_U4208;
  assign new_P1_U6885 = ~new_P1_U4494 | ~new_P1_U3283;
  assign new_P1_U6886 = ~new_P1_U4159 | ~new_P1_R2144_U50;
  assign new_P1_U6887 = ~new_P1_ADD_371_U20 | ~new_P1_U4208;
  assign new_P1_U6888 = ~new_P1_U2605 | ~new_P1_U3284;
  assign new_P1_U6889 = ~new_P1_U4159 | ~new_P1_R2144_U43;
  assign new_P1_U6890 = ~new_P1_ADD_371_U4 | ~new_P1_U4208;
  assign new_P1_U6891 = ~new_P1_U4494 | ~new_P1_U3283;
  assign new_P1_U6892 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__1_;
  assign new_P1_U6893 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__1_;
  assign new_P1_U6894 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__1_;
  assign new_P1_U6895 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__1_;
  assign new_P1_U6896 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__1_;
  assign new_P1_U6897 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__1_;
  assign new_P1_U6898 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__1_;
  assign new_P1_U6899 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__1_;
  assign new_P1_U6900 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__1_;
  assign new_P1_U6901 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__1_;
  assign new_P1_U6902 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__1_;
  assign new_P1_U6903 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__1_;
  assign new_P1_U6904 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__1_;
  assign new_P1_U6905 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__1_;
  assign new_P1_U6906 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__1_;
  assign new_P1_U6907 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__1_;
  assign new_P1_U6908 = ~new_P1_U4029 | ~new_P1_U4030 | ~new_P1_U4032 | ~new_P1_U4031;
  assign new_P1_U6909 = ~new_P1_U3405 | ~new_P1_U3418;
  assign new_P1_U6910 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__0_;
  assign new_P1_U6911 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__0_;
  assign new_P1_U6912 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__0_;
  assign new_P1_U6913 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__0_;
  assign new_P1_U6914 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__0_;
  assign new_P1_U6915 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__0_;
  assign new_P1_U6916 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__0_;
  assign new_P1_U6917 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__0_;
  assign new_P1_U6918 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__0_;
  assign new_P1_U6919 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__0_;
  assign new_P1_U6920 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__0_;
  assign new_P1_U6921 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__0_;
  assign new_P1_U6922 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__0_;
  assign new_P1_U6923 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__0_;
  assign new_P1_U6924 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__0_;
  assign new_P1_U6925 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__0_;
  assign new_P1_U6926 = ~new_P1_U4033 | ~new_P1_U4034 | ~new_P1_U4036 | ~new_P1_U4035;
  assign new_P1_U6927 = ~new_P1_U4207 | ~new_P1_U3234;
  assign new_P1_U6928 = ~new_P1_U2355 | ~new_P1_SUB_357_U8;
  assign new_P1_U6929 = ~new_P1_U4207 | ~new_P1_U3233;
  assign new_P1_U6930 = ~new_P1_SUB_357_U6 | ~new_P1_U2355;
  assign new_P1_U6931 = ~new_P1_U4207 | ~new_P1_U3232;
  assign new_P1_U6932 = ~new_P1_SUB_357_U9 | ~new_P1_U2355;
  assign new_P1_U6933 = ~new_P1_U4207 | ~new_P1_U3231;
  assign new_P1_U6934 = ~new_P1_SUB_357_U13 | ~new_P1_U2355;
  assign new_P1_U6935 = ~new_P1_U4207 | ~new_P1_U3230;
  assign new_P1_U6936 = ~new_P1_SUB_357_U11 | ~new_P1_U2355;
  assign new_P1_U6937 = ~new_P1_R2182_U25 | ~new_P1_U3294;
  assign new_P1_U6938 = ~new_P1_U4207 | ~new_P1_U3229;
  assign new_P1_U6939 = ~new_P1_SUB_357_U12 | ~new_P1_U2355;
  assign new_P1_U6940 = ~new_P1_R2182_U42 | ~new_P1_U3294;
  assign new_P1_U6941 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__7_;
  assign new_P1_U6942 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__7_;
  assign new_P1_U6943 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__7_;
  assign new_P1_U6944 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__7_;
  assign new_P1_U6945 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__7_;
  assign new_P1_U6946 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__7_;
  assign new_P1_U6947 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__7_;
  assign new_P1_U6948 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__7_;
  assign new_P1_U6949 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__7_;
  assign new_P1_U6950 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__7_;
  assign new_P1_U6951 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__7_;
  assign new_P1_U6952 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__7_;
  assign new_P1_U6953 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__7_;
  assign new_P1_U6954 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__7_;
  assign new_P1_U6955 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__7_;
  assign new_P1_U6956 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__7_;
  assign new_P1_U6957 = ~new_P1_U4037 | ~new_P1_U4038 | ~new_P1_U4040 | ~new_P1_U4039;
  assign new_P1_U6958 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__6_;
  assign new_P1_U6959 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__6_;
  assign new_P1_U6960 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__6_;
  assign new_P1_U6961 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__6_;
  assign new_P1_U6962 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__6_;
  assign new_P1_U6963 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__6_;
  assign new_P1_U6964 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__6_;
  assign new_P1_U6965 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__6_;
  assign new_P1_U6966 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__6_;
  assign new_P1_U6967 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__6_;
  assign new_P1_U6968 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__6_;
  assign new_P1_U6969 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__6_;
  assign new_P1_U6970 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__6_;
  assign new_P1_U6971 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__6_;
  assign new_P1_U6972 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__6_;
  assign new_P1_U6973 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__6_;
  assign new_P1_U6974 = ~new_P1_U4041 | ~new_P1_U4042 | ~new_P1_U4044 | ~new_P1_U4043;
  assign new_P1_U6975 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__5_;
  assign new_P1_U6976 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__5_;
  assign new_P1_U6977 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__5_;
  assign new_P1_U6978 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__5_;
  assign new_P1_U6979 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__5_;
  assign new_P1_U6980 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__5_;
  assign new_P1_U6981 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__5_;
  assign new_P1_U6982 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__5_;
  assign new_P1_U6983 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__5_;
  assign new_P1_U6984 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__5_;
  assign new_P1_U6985 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__5_;
  assign new_P1_U6986 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__5_;
  assign new_P1_U6987 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__5_;
  assign new_P1_U6988 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__5_;
  assign new_P1_U6989 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__5_;
  assign new_P1_U6990 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__5_;
  assign new_P1_U6991 = ~new_P1_U4045 | ~new_P1_U4046 | ~new_P1_U4048 | ~new_P1_U4047;
  assign new_P1_U6992 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__4_;
  assign new_P1_U6993 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__4_;
  assign new_P1_U6994 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__4_;
  assign new_P1_U6995 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__4_;
  assign new_P1_U6996 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__4_;
  assign new_P1_U6997 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__4_;
  assign new_P1_U6998 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__4_;
  assign new_P1_U6999 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__4_;
  assign new_P1_U7000 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__4_;
  assign new_P1_U7001 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__4_;
  assign new_P1_U7002 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__4_;
  assign new_P1_U7003 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__4_;
  assign new_P1_U7004 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__4_;
  assign new_P1_U7005 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__4_;
  assign new_P1_U7006 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__4_;
  assign new_P1_U7007 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__3_;
  assign new_P1_U7008 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__3_;
  assign new_P1_U7009 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__3_;
  assign new_P1_U7010 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__3_;
  assign new_P1_U7011 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__3_;
  assign new_P1_U7012 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__3_;
  assign new_P1_U7013 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__3_;
  assign new_P1_U7014 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__3_;
  assign new_P1_U7015 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__3_;
  assign new_P1_U7016 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__3_;
  assign new_P1_U7017 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__3_;
  assign new_P1_U7018 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__3_;
  assign new_P1_U7019 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__3_;
  assign new_P1_U7020 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__3_;
  assign new_P1_U7021 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__3_;
  assign new_P1_U7022 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__3_;
  assign new_P1_U7023 = ~new_P1_U4053 | ~new_P1_U4054 | ~new_P1_U4056 | ~new_P1_U4055;
  assign new_P1_U7024 = ~new_P1_U2564 | ~P1_INSTQUEUE_REG_15__2_;
  assign new_P1_U7025 = ~new_P1_U2563 | ~P1_INSTQUEUE_REG_14__2_;
  assign new_P1_U7026 = ~new_P1_U2562 | ~P1_INSTQUEUE_REG_13__2_;
  assign new_P1_U7027 = ~new_P1_U2561 | ~P1_INSTQUEUE_REG_12__2_;
  assign new_P1_U7028 = ~new_P1_U2559 | ~P1_INSTQUEUE_REG_11__2_;
  assign new_P1_U7029 = ~new_P1_U2558 | ~P1_INSTQUEUE_REG_10__2_;
  assign new_P1_U7030 = ~new_P1_U2557 | ~P1_INSTQUEUE_REG_9__2_;
  assign new_P1_U7031 = ~new_P1_U2556 | ~P1_INSTQUEUE_REG_8__2_;
  assign new_P1_U7032 = ~new_P1_U2554 | ~P1_INSTQUEUE_REG_7__2_;
  assign new_P1_U7033 = ~new_P1_U2553 | ~P1_INSTQUEUE_REG_6__2_;
  assign new_P1_U7034 = ~new_P1_U2552 | ~P1_INSTQUEUE_REG_5__2_;
  assign new_P1_U7035 = ~new_P1_U2551 | ~P1_INSTQUEUE_REG_4__2_;
  assign new_P1_U7036 = ~new_P1_U2549 | ~P1_INSTQUEUE_REG_3__2_;
  assign new_P1_U7037 = ~new_P1_U2548 | ~P1_INSTQUEUE_REG_2__2_;
  assign new_P1_U7038 = ~new_P1_U2547 | ~P1_INSTQUEUE_REG_1__2_;
  assign new_P1_U7039 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__2_;
  assign new_P1_U7040 = ~new_P1_U4057 | ~new_P1_U4058 | ~new_P1_U4060 | ~new_P1_U4059;
  assign new_P1_U7041 = ~new_P1_U4207 | ~new_P1_U3228;
  assign new_P1_U7042 = ~new_P1_SUB_357_U7 | ~new_P1_U2355;
  assign new_P1_U7043 = ~new_P1_R2182_U33 | ~new_P1_U3294;
  assign new_P1_U7044 = ~new_P1_U4207 | ~new_P1_U3227;
  assign new_P1_U7045 = ~new_P1_SUB_357_U10 | ~new_P1_U2355;
  assign new_P1_U7046 = ~new_P1_R2182_U34 | ~new_P1_U3294;
  assign new_P1_U7047 = ~new_P1_U4206 | ~new_P1_U3234;
  assign new_P1_U7048 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__7_;
  assign new_P1_U7049 = ~new_P1_U4206 | ~new_P1_U3233;
  assign new_P1_U7050 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__6_;
  assign new_P1_U7051 = ~new_P1_U4206 | ~new_P1_U3232;
  assign new_P1_U7052 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__5_;
  assign new_P1_U7053 = ~new_P1_U4206 | ~new_P1_U3231;
  assign new_P1_U7054 = ~new_P1_U4206 | ~new_P1_U3230;
  assign new_P1_U7055 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__3_;
  assign new_P1_U7056 = ~new_P1_U4206 | ~new_P1_U3229;
  assign new_P1_U7057 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__2_;
  assign new_P1_U7058 = ~new_P1_U4206 | ~new_P1_U3228;
  assign new_P1_U7059 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__1_;
  assign new_P1_U7060 = ~new_P1_U4206 | ~new_P1_U3227;
  assign new_P1_U7061 = ~new_P1_U3234 | ~new_P1_U4400;
  assign new_P1_U7062 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__0_;
  assign new_P1_U7063 = ~new_P1_U3428 | ~new_P1_U3427;
  assign new_P1_U7064 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3264;
  assign new_P1_U7065 = ~new_P1_U3445;
  assign new_P1_U7066 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__7_;
  assign new_P1_U7067 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__7_;
  assign new_P1_U7068 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__7_;
  assign new_P1_U7069 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__7_;
  assign new_P1_U7070 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__7_;
  assign new_P1_U7071 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__7_;
  assign new_P1_U7072 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__7_;
  assign new_P1_U7073 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__7_;
  assign new_P1_U7074 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__7_;
  assign new_P1_U7075 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__7_;
  assign new_P1_U7076 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__7_;
  assign new_P1_U7077 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__7_;
  assign new_P1_U7078 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__7_;
  assign new_P1_U7079 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__7_;
  assign new_P1_U7080 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__7_;
  assign new_P1_U7081 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__7_;
  assign new_P1_U7082 = ~new_P1_U4063 | ~new_P1_U4064 | ~new_P1_U4066 | ~new_P1_U4065;
  assign new_P1_U7083 = ~new_P1_U3425 | ~new_P1_U3421;
  assign new_P1_U7084 = ~new_P1_U4073 | ~new_P1_U4191;
  assign new_P1_U7085 = ~new_P1_U7084 | ~new_P1_U3422;
  assign new_P1_U7086 = ~new_P1_U4503 | ~new_P1_U3278;
  assign new_P1_U7087 = ~new_P1_U3245;
  assign new_P1_U7088 = ~new_P1_U3394 | ~new_P1_U4154 | ~new_P1_U4400 | ~new_P1_U4503;
  assign new_P1_U7089 = ~new_P1_U4189 | ~P1_STATE2_REG_0_;
  assign new_P1_U7090 = ~new_P1_U4067 | ~new_P1_U3245;
  assign new_P1_U7091 = ~new_P1_U3451;
  assign new_P1_U7092 = ~new_P1_U7629 | ~new_P1_U3451 | ~new_P1_U5492;
  assign new_P1_U7093 = ~new_P1_U4194 | ~new_P1_U7092;
  assign new_P1_U7094 = ~new_P1_U3450;
  assign new_P1_U7095 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_U3297;
  assign new_P1_U7096 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3450;
  assign new_P1_U7097 = ~new_P1_U4203 | ~new_P1_U3360;
  assign new_P1_U7098 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__6_;
  assign new_P1_U7099 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__6_;
  assign new_P1_U7100 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__6_;
  assign new_P1_U7101 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__6_;
  assign new_P1_U7102 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__6_;
  assign new_P1_U7103 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__6_;
  assign new_P1_U7104 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__6_;
  assign new_P1_U7105 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__6_;
  assign new_P1_U7106 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__6_;
  assign new_P1_U7107 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__6_;
  assign new_P1_U7108 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__6_;
  assign new_P1_U7109 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__6_;
  assign new_P1_U7110 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__6_;
  assign new_P1_U7111 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__6_;
  assign new_P1_U7112 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__6_;
  assign new_P1_U7113 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__6_;
  assign new_P1_U7114 = ~new_P1_U4079 | ~new_P1_U4080 | ~new_P1_U4082 | ~new_P1_U4081;
  assign new_P1_U7115 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__5_;
  assign new_P1_U7116 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__5_;
  assign new_P1_U7117 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__5_;
  assign new_P1_U7118 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__5_;
  assign new_P1_U7119 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__5_;
  assign new_P1_U7120 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__5_;
  assign new_P1_U7121 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__5_;
  assign new_P1_U7122 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__5_;
  assign new_P1_U7123 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__5_;
  assign new_P1_U7124 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__5_;
  assign new_P1_U7125 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__5_;
  assign new_P1_U7126 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__5_;
  assign new_P1_U7127 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__5_;
  assign new_P1_U7128 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__5_;
  assign new_P1_U7129 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__5_;
  assign new_P1_U7130 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__5_;
  assign new_P1_U7131 = ~new_P1_U4083 | ~new_P1_U4084 | ~new_P1_U4086 | ~new_P1_U4085;
  assign new_P1_U7132 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__4_;
  assign new_P1_U7133 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__4_;
  assign new_P1_U7134 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__4_;
  assign new_P1_U7135 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__4_;
  assign new_P1_U7136 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__4_;
  assign new_P1_U7137 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__4_;
  assign new_P1_U7138 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__4_;
  assign new_P1_U7139 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__4_;
  assign new_P1_U7140 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__4_;
  assign new_P1_U7141 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__4_;
  assign new_P1_U7142 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__4_;
  assign new_P1_U7143 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__4_;
  assign new_P1_U7144 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__4_;
  assign new_P1_U7145 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__4_;
  assign new_P1_U7146 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__4_;
  assign new_P1_U7147 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__3_;
  assign new_P1_U7148 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__3_;
  assign new_P1_U7149 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__3_;
  assign new_P1_U7150 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__3_;
  assign new_P1_U7151 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__3_;
  assign new_P1_U7152 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__3_;
  assign new_P1_U7153 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__3_;
  assign new_P1_U7154 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__3_;
  assign new_P1_U7155 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__3_;
  assign new_P1_U7156 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__3_;
  assign new_P1_U7157 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__3_;
  assign new_P1_U7158 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__3_;
  assign new_P1_U7159 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__3_;
  assign new_P1_U7160 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__3_;
  assign new_P1_U7161 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__3_;
  assign new_P1_U7162 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__3_;
  assign new_P1_U7163 = ~new_P1_U4092 | ~new_P1_U4093 | ~new_P1_U4095 | ~new_P1_U4094;
  assign new_P1_U7164 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__2_;
  assign new_P1_U7165 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__2_;
  assign new_P1_U7166 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__2_;
  assign new_P1_U7167 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__2_;
  assign new_P1_U7168 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__2_;
  assign new_P1_U7169 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__2_;
  assign new_P1_U7170 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__2_;
  assign new_P1_U7171 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__2_;
  assign new_P1_U7172 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__2_;
  assign new_P1_U7173 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__2_;
  assign new_P1_U7174 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__2_;
  assign new_P1_U7175 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__2_;
  assign new_P1_U7176 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__2_;
  assign new_P1_U7177 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__2_;
  assign new_P1_U7178 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__2_;
  assign new_P1_U7179 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__2_;
  assign new_P1_U7180 = ~new_P1_U4096 | ~new_P1_U4097 | ~new_P1_U4099 | ~new_P1_U4098;
  assign new_P1_U7181 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__1_;
  assign new_P1_U7182 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__1_;
  assign new_P1_U7183 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__1_;
  assign new_P1_U7184 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__1_;
  assign new_P1_U7185 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__1_;
  assign new_P1_U7186 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__1_;
  assign new_P1_U7187 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__1_;
  assign new_P1_U7188 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__1_;
  assign new_P1_U7189 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__1_;
  assign new_P1_U7190 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__1_;
  assign new_P1_U7191 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__1_;
  assign new_P1_U7192 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__1_;
  assign new_P1_U7193 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__1_;
  assign new_P1_U7194 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__1_;
  assign new_P1_U7195 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__1_;
  assign new_P1_U7196 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__1_;
  assign new_P1_U7197 = ~new_P1_U4100 | ~new_P1_U4101 | ~new_P1_U4103 | ~new_P1_U4102;
  assign new_P1_U7198 = ~new_P1_U2582 | ~P1_INSTQUEUE_REG_8__0_;
  assign new_P1_U7199 = ~new_P1_U2581 | ~P1_INSTQUEUE_REG_9__0_;
  assign new_P1_U7200 = ~new_P1_U2580 | ~P1_INSTQUEUE_REG_10__0_;
  assign new_P1_U7201 = ~new_P1_U2579 | ~P1_INSTQUEUE_REG_11__0_;
  assign new_P1_U7202 = ~new_P1_U2577 | ~P1_INSTQUEUE_REG_12__0_;
  assign new_P1_U7203 = ~new_P1_U2576 | ~P1_INSTQUEUE_REG_13__0_;
  assign new_P1_U7204 = ~new_P1_U2575 | ~P1_INSTQUEUE_REG_14__0_;
  assign new_P1_U7205 = ~new_P1_U2574 | ~P1_INSTQUEUE_REG_15__0_;
  assign new_P1_U7206 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__0_;
  assign new_P1_U7207 = ~new_P1_U2572 | ~P1_INSTQUEUE_REG_1__0_;
  assign new_P1_U7208 = ~new_P1_U2571 | ~P1_INSTQUEUE_REG_2__0_;
  assign new_P1_U7209 = ~new_P1_U2570 | ~P1_INSTQUEUE_REG_3__0_;
  assign new_P1_U7210 = ~new_P1_U2568 | ~P1_INSTQUEUE_REG_4__0_;
  assign new_P1_U7211 = ~new_P1_U2567 | ~P1_INSTQUEUE_REG_5__0_;
  assign new_P1_U7212 = ~new_P1_U2566 | ~P1_INSTQUEUE_REG_6__0_;
  assign new_P1_U7213 = ~new_P1_U2565 | ~P1_INSTQUEUE_REG_7__0_;
  assign new_P1_U7214 = ~new_P1_U4104 | ~new_P1_U4105 | ~new_P1_U4107 | ~new_P1_U4106;
  assign new_P1_U7215 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_U3297;
  assign new_P1_U7216 = ~new_P1_U4203 | ~new_P1_U3455;
  assign new_P1_U7217 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_U3297;
  assign new_P1_U7218 = ~new_P1_U4203 | ~new_P1_U3235;
  assign new_P1_U7219 = ~new_P1_U4183;
  assign new_P1_U7220 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__7_;
  assign new_P1_U7221 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__7_;
  assign new_P1_U7222 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__7_;
  assign new_P1_U7223 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__7_;
  assign new_P1_U7224 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__7_;
  assign new_P1_U7225 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__7_;
  assign new_P1_U7226 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__7_;
  assign new_P1_U7227 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__7_;
  assign new_P1_U7228 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__7_;
  assign new_P1_U7229 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__7_;
  assign new_P1_U7230 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__7_;
  assign new_P1_U7231 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__7_;
  assign new_P1_U7232 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__7_;
  assign new_P1_U7233 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__7_;
  assign new_P1_U7234 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__7_;
  assign new_P1_U7235 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__7_;
  assign new_P1_U7236 = ~new_P1_U4121 | ~new_P1_U4122 | ~new_P1_U4124 | ~new_P1_U4123;
  assign new_P1_U7237 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__6_;
  assign new_P1_U7238 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__6_;
  assign new_P1_U7239 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__6_;
  assign new_P1_U7240 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__6_;
  assign new_P1_U7241 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__6_;
  assign new_P1_U7242 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__6_;
  assign new_P1_U7243 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__6_;
  assign new_P1_U7244 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__6_;
  assign new_P1_U7245 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__6_;
  assign new_P1_U7246 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__6_;
  assign new_P1_U7247 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__6_;
  assign new_P1_U7248 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__6_;
  assign new_P1_U7249 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__6_;
  assign new_P1_U7250 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__6_;
  assign new_P1_U7251 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__6_;
  assign new_P1_U7252 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__6_;
  assign new_P1_U7253 = ~new_P1_U4125 | ~new_P1_U4126 | ~new_P1_U4128 | ~new_P1_U4127;
  assign new_P1_U7254 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__5_;
  assign new_P1_U7255 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__5_;
  assign new_P1_U7256 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__5_;
  assign new_P1_U7257 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__5_;
  assign new_P1_U7258 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__5_;
  assign new_P1_U7259 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__5_;
  assign new_P1_U7260 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__5_;
  assign new_P1_U7261 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__5_;
  assign new_P1_U7262 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__5_;
  assign new_P1_U7263 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__5_;
  assign new_P1_U7264 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__5_;
  assign new_P1_U7265 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__5_;
  assign new_P1_U7266 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__5_;
  assign new_P1_U7267 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__5_;
  assign new_P1_U7268 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__5_;
  assign new_P1_U7269 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__5_;
  assign new_P1_U7270 = ~new_P1_U4129 | ~new_P1_U4130 | ~new_P1_U4132 | ~new_P1_U4131;
  assign new_P1_U7271 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__4_;
  assign new_P1_U7272 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__4_;
  assign new_P1_U7273 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__4_;
  assign new_P1_U7274 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__4_;
  assign new_P1_U7275 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__4_;
  assign new_P1_U7276 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__4_;
  assign new_P1_U7277 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__4_;
  assign new_P1_U7278 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__4_;
  assign new_P1_U7279 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__4_;
  assign new_P1_U7280 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__4_;
  assign new_P1_U7281 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__4_;
  assign new_P1_U7282 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__4_;
  assign new_P1_U7283 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__4_;
  assign new_P1_U7284 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__4_;
  assign new_P1_U7285 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__4_;
  assign new_P1_U7286 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__3_;
  assign new_P1_U7287 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__3_;
  assign new_P1_U7288 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__3_;
  assign new_P1_U7289 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__3_;
  assign new_P1_U7290 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__3_;
  assign new_P1_U7291 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__3_;
  assign new_P1_U7292 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__3_;
  assign new_P1_U7293 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__3_;
  assign new_P1_U7294 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__3_;
  assign new_P1_U7295 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__3_;
  assign new_P1_U7296 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__3_;
  assign new_P1_U7297 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__3_;
  assign new_P1_U7298 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__3_;
  assign new_P1_U7299 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__3_;
  assign new_P1_U7300 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__3_;
  assign new_P1_U7301 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__3_;
  assign new_P1_U7302 = ~new_P1_U4137 | ~new_P1_U4138 | ~new_P1_U4140 | ~new_P1_U4139;
  assign new_P1_U7303 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__2_;
  assign new_P1_U7304 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__2_;
  assign new_P1_U7305 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__2_;
  assign new_P1_U7306 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__2_;
  assign new_P1_U7307 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__2_;
  assign new_P1_U7308 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__2_;
  assign new_P1_U7309 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__2_;
  assign new_P1_U7310 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__2_;
  assign new_P1_U7311 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__2_;
  assign new_P1_U7312 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__2_;
  assign new_P1_U7313 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__2_;
  assign new_P1_U7314 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__2_;
  assign new_P1_U7315 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__2_;
  assign new_P1_U7316 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__2_;
  assign new_P1_U7317 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__2_;
  assign new_P1_U7318 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__2_;
  assign new_P1_U7319 = ~new_P1_U4141 | ~new_P1_U4142 | ~new_P1_U4144 | ~new_P1_U4143;
  assign new_P1_U7320 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__1_;
  assign new_P1_U7321 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__1_;
  assign new_P1_U7322 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__1_;
  assign new_P1_U7323 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__1_;
  assign new_P1_U7324 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__1_;
  assign new_P1_U7325 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__1_;
  assign new_P1_U7326 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__1_;
  assign new_P1_U7327 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__1_;
  assign new_P1_U7328 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__1_;
  assign new_P1_U7329 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__1_;
  assign new_P1_U7330 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__1_;
  assign new_P1_U7331 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__1_;
  assign new_P1_U7332 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__1_;
  assign new_P1_U7333 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__1_;
  assign new_P1_U7334 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__1_;
  assign new_P1_U7335 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__1_;
  assign new_P1_U7336 = ~new_P1_U4145 | ~new_P1_U4146 | ~new_P1_U4148 | ~new_P1_U4147;
  assign new_P1_U7337 = ~new_P1_U2602 | ~P1_INSTQUEUE_REG_8__0_;
  assign new_P1_U7338 = ~new_P1_U2601 | ~P1_INSTQUEUE_REG_9__0_;
  assign new_P1_U7339 = ~new_P1_U2600 | ~P1_INSTQUEUE_REG_10__0_;
  assign new_P1_U7340 = ~new_P1_U2599 | ~P1_INSTQUEUE_REG_11__0_;
  assign new_P1_U7341 = ~new_P1_U2597 | ~P1_INSTQUEUE_REG_12__0_;
  assign new_P1_U7342 = ~new_P1_U2596 | ~P1_INSTQUEUE_REG_13__0_;
  assign new_P1_U7343 = ~new_P1_U2595 | ~P1_INSTQUEUE_REG_14__0_;
  assign new_P1_U7344 = ~new_P1_U2594 | ~P1_INSTQUEUE_REG_15__0_;
  assign new_P1_U7345 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__0_;
  assign new_P1_U7346 = ~new_P1_U2591 | ~P1_INSTQUEUE_REG_1__0_;
  assign new_P1_U7347 = ~new_P1_U2590 | ~P1_INSTQUEUE_REG_2__0_;
  assign new_P1_U7348 = ~new_P1_U2589 | ~P1_INSTQUEUE_REG_3__0_;
  assign new_P1_U7349 = ~new_P1_U2587 | ~P1_INSTQUEUE_REG_4__0_;
  assign new_P1_U7350 = ~new_P1_U2586 | ~P1_INSTQUEUE_REG_5__0_;
  assign new_P1_U7351 = ~new_P1_U2585 | ~P1_INSTQUEUE_REG_6__0_;
  assign new_P1_U7352 = ~new_P1_U2584 | ~P1_INSTQUEUE_REG_7__0_;
  assign new_P1_U7353 = ~new_P1_U4149 | ~new_P1_U4150 | ~new_P1_U4152 | ~new_P1_U4151;
  assign new_P1_U7354 = ~new_P1_U4234 | ~new_P1_U4231 | ~new_P1_U2354;
  assign new_P1_U7355 = ~new_P1_U4153 | ~new_P1_U7087;
  assign new_P1_U7356 = ~new_P1_U3396 | ~new_P1_U3410;
  assign new_P1_U7357 = ~new_P1_U4234 | ~new_P1_U7356;
  assign new_P1_U7358 = ~new_P1_U4190 | ~new_P1_U2452;
  assign new_P1_U7359 = ~new_P1_U7355 | ~new_P1_U3271;
  assign new_P1_U7360 = ~new_P1_U4208 | ~new_P1_U7088;
  assign new_P1_U7361 = ~new_P1_U4160 | ~new_P1_U4208;
  assign new_P1_U7362 = ~new_P1_U2451 | ~new_P1_U4210;
  assign new_P1_U7363 = ~new_P1_U7361 | ~new_P1_U7362 | ~new_P1_U4195 | ~new_P1_U3420 | ~new_P1_U3434;
  assign new_P1_U7364 = ~new_P1_R2238_U6 | ~new_P1_U7363;
  assign new_P1_U7365 = ~new_P1_SUB_450_U6 | ~new_P1_U2354;
  assign new_P1_U7366 = ~new_P1_R2238_U19 | ~new_P1_U7363;
  assign new_P1_U7367 = ~new_P1_SUB_450_U19 | ~new_P1_U2354;
  assign new_P1_U7368 = ~new_P1_R2238_U20 | ~new_P1_U7363;
  assign new_P1_U7369 = ~new_P1_SUB_450_U20 | ~new_P1_U2354;
  assign new_P1_U7370 = ~new_P1_R2238_U21 | ~new_P1_U7363;
  assign new_P1_U7371 = ~new_P1_SUB_450_U21 | ~new_P1_U2354;
  assign new_P1_U7372 = ~new_P1_R2238_U22 | ~new_P1_U7363;
  assign new_P1_U7373 = ~new_P1_SUB_450_U22 | ~new_P1_U2354;
  assign new_P1_U7374 = ~new_P1_R2238_U7 | ~new_P1_U7363;
  assign new_P1_U7375 = ~new_P1_SUB_450_U7 | ~new_P1_U2354;
  assign new_P1_U7376 = ~new_P1_R2238_U19 | ~new_P1_U4192;
  assign new_P1_U7377 = ~P1_INSTQUEUERD_ADDR_REG_4_ | ~new_P1_U3294;
  assign new_P1_U7378 = ~new_P1_R2238_U20 | ~new_P1_U4192;
  assign new_P1_U7379 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3294;
  assign new_P1_U7380 = ~P1_STATE2_REG_0_ | ~new_P1_U4173;
  assign new_P1_U7381 = ~new_P1_U3420 | ~new_P1_U7380;
  assign new_P1_U7382 = ~new_P1_R2238_U21 | ~new_P1_U4192;
  assign new_P1_U7383 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3294;
  assign new_P1_U7384 = ~new_P1_U2450 | ~new_P1_U3271;
  assign new_P1_U7385 = ~new_P1_R2238_U22 | ~new_P1_U4192;
  assign new_P1_U7386 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3294;
  assign new_P1_U7387 = ~new_P1_U2451 | ~new_P1_U3284;
  assign new_P1_U7388 = ~new_P1_R2238_U7 | ~new_P1_U4192;
  assign new_P1_U7389 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~new_P1_U3294;
  assign new_P1_U7390 = ~new_P1_U3393 | ~new_P1_U3290;
  assign new_P1_U7391 = ~new_P1_U3284 | ~new_P1_U3449;
  assign new_P1_U7392 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_U7391;
  assign new_P1_U7393 = ~P1_EBX_REG_9_ | ~new_P1_U7390;
  assign new_P1_U7394 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_U7391;
  assign new_P1_U7395 = ~P1_EBX_REG_8_ | ~new_P1_U7390;
  assign new_P1_U7396 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_U7391;
  assign new_P1_U7397 = ~P1_EBX_REG_7_ | ~new_P1_U7390;
  assign new_P1_U7398 = ~P1_INSTADDRPOINTER_REG_6_ | ~new_P1_U7391;
  assign new_P1_U7399 = ~P1_EBX_REG_6_ | ~new_P1_U7390;
  assign new_P1_U7400 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_U7391;
  assign new_P1_U7401 = ~P1_EBX_REG_5_ | ~new_P1_U7390;
  assign new_P1_U7402 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_U7391;
  assign new_P1_U7403 = ~P1_EBX_REG_4_ | ~new_P1_U7390;
  assign new_P1_U7404 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_U7391;
  assign new_P1_U7405 = ~P1_EBX_REG_31_ | ~new_P1_U7390;
  assign new_P1_U7406 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_U7391;
  assign new_P1_U7407 = ~P1_EBX_REG_30_ | ~new_P1_U7390;
  assign new_P1_U7408 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_U7391;
  assign new_P1_U7409 = ~P1_EBX_REG_3_ | ~new_P1_U7390;
  assign new_P1_U7410 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_U7391;
  assign new_P1_U7411 = ~P1_EBX_REG_29_ | ~new_P1_U7390;
  assign new_P1_U7412 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_U7391;
  assign new_P1_U7413 = ~P1_EBX_REG_28_ | ~new_P1_U7390;
  assign new_P1_U7414 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_U7391;
  assign new_P1_U7415 = ~P1_EBX_REG_27_ | ~new_P1_U7390;
  assign new_P1_U7416 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_U7391;
  assign new_P1_U7417 = ~P1_EBX_REG_26_ | ~new_P1_U7390;
  assign new_P1_U7418 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_U7391;
  assign new_P1_U7419 = ~P1_EBX_REG_25_ | ~new_P1_U7390;
  assign new_P1_U7420 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_U7391;
  assign new_P1_U7421 = ~P1_EBX_REG_24_ | ~new_P1_U7390;
  assign new_P1_U7422 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_U7391;
  assign new_P1_U7423 = ~P1_EBX_REG_23_ | ~new_P1_U7390;
  assign new_P1_U7424 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_U7391;
  assign new_P1_U7425 = ~P1_EBX_REG_22_ | ~new_P1_U7390;
  assign new_P1_U7426 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_U7391;
  assign new_P1_U7427 = ~P1_EBX_REG_21_ | ~new_P1_U7390;
  assign new_P1_U7428 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_U7391;
  assign new_P1_U7429 = ~P1_EBX_REG_20_ | ~new_P1_U7390;
  assign new_P1_U7430 = ~P1_INSTADDRPOINTER_REG_2_ | ~new_P1_U7391;
  assign new_P1_U7431 = ~P1_EBX_REG_2_ | ~new_P1_U7390;
  assign new_P1_U7432 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_U7391;
  assign new_P1_U7433 = ~P1_EBX_REG_19_ | ~new_P1_U7390;
  assign new_P1_U7434 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_U7391;
  assign new_P1_U7435 = ~P1_EBX_REG_18_ | ~new_P1_U7390;
  assign new_P1_U7436 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_U7391;
  assign new_P1_U7437 = ~P1_EBX_REG_17_ | ~new_P1_U7390;
  assign new_P1_U7438 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_U7391;
  assign new_P1_U7439 = ~P1_EBX_REG_16_ | ~new_P1_U7390;
  assign new_P1_U7440 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_U7391;
  assign new_P1_U7441 = ~P1_EBX_REG_15_ | ~new_P1_U7390;
  assign new_P1_U7442 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_U7391;
  assign new_P1_U7443 = ~P1_EBX_REG_14_ | ~new_P1_U7390;
  assign new_P1_U7444 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_U7391;
  assign new_P1_U7445 = ~P1_EBX_REG_13_ | ~new_P1_U7390;
  assign new_P1_U7446 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_U7391;
  assign new_P1_U7447 = ~P1_EBX_REG_12_ | ~new_P1_U7390;
  assign new_P1_U7448 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_U7391;
  assign new_P1_U7449 = ~P1_EBX_REG_11_ | ~new_P1_U7390;
  assign new_P1_U7450 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_U7391;
  assign new_P1_U7451 = ~P1_EBX_REG_10_ | ~new_P1_U7390;
  assign new_P1_U7452 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_U7391;
  assign new_P1_U7453 = ~P1_EBX_REG_1_ | ~new_P1_U7390;
  assign new_P1_U7454 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_U7391;
  assign new_P1_U7455 = ~P1_EBX_REG_0_ | ~new_P1_U7390;
  assign new_P1_U7456 = ~new_P1_U4477 | ~new_P1_U4496;
  assign new_P1_U7457 = ~new_P1_U2430 | ~P1_INSTQUEUERD_ADDR_REG_4_;
  assign new_P1_U7458 = ~new_P1_U3489 | ~new_P1_U3262;
  assign new_P1_U7459 = ~new_P1_U2430 | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7460 = ~new_P1_U3490 | ~new_P1_U3262;
  assign new_P1_U7461 = ~new_P1_U3470 | ~P1_FLUSH_REG | ~new_P1_U2446;
  assign new_P1_U7462 = ~new_P1_U2430 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U7463 = ~new_P1_U3491 | ~new_P1_U3262;
  assign new_P1_U7464 = ~new_P1_U7712 | ~new_P1_U2446 | ~P1_FLUSH_REG;
  assign new_P1_U7465 = ~new_P1_U2430 | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U7466 = ~new_P1_U3492 | ~new_P1_U3262;
  assign new_P1_U7467 = ~new_P1_U2430 | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7468 = ~P1_STATE_REG_0_ | ~new_P1_U4185;
  assign new_P1_U7469 = new_U210 | P1_STATE2_REG_2_;
  assign new_P1_U7470 = ~new_P1_U4110 | ~new_P1_U7218;
  assign new_P1_U7471 = ~new_P1_U7084 | ~new_P1_U3422;
  assign new_P1_U7472 = ~new_P1_U4211 | ~P1_STATE2_REG_0_;
  assign new_P1_U7473 = ~new_P1_U4212 | ~P1_STATE2_REG_0_;
  assign new_P1_U7474 = ~new_P1_U4213 | ~P1_STATE2_REG_0_;
  assign new_P1_U7475 = ~new_P1_U4236 | ~P1_STATE2_REG_0_;
  assign new_P1_U7476 = ~new_P1_U4264 | ~P1_STATE2_REG_0_;
  assign new_P1_U7477 = ~P1_STATE2_REG_0_ | ~new_P1_U7632;
  assign new_P1_U7478 = ~new_P1_U2608 | ~new_P1_U3266;
  assign new_P1_U7479 = ~new_P1_U4120 | ~new_P1_U4118 | ~new_P1_U4117 | ~new_P1_U7093;
  assign new_P1_U7480 = ~P1_STATE2_REG_0_ | ~new_P1_U7632;
  assign new_P1_U7481 = ~new_P1_U2379 | ~new_P1_U3429;
  assign new_P1_U7482 = ~new_P1_U2369 | ~new_P1_U6367;
  assign new_P1_U7483 = ~new_P1_U3888 | ~new_P1_U2369;
  assign new_P1_U7484 = ~new_P1_U7482 | ~new_P1_U7481 | ~new_P1_U4229;
  assign new_P1_U7485 = ~new_P1_U7483 | ~new_P1_U4230;
  assign new_P1_U7486 = ~new_P1_U4194 | ~new_P1_U5491 | ~new_P1_U4171;
  assign new_P1_U7487 = ~new_P1_U7091 | ~new_P1_U4194;
  assign new_P1_U7488 = ~new_P1_U4194 | ~new_P1_U3392;
  assign new_P1_U7489 = ~new_P1_U4236 | ~P1_STATE2_REG_0_;
  assign new_P1_U7490 = ~new_P1_U4072 | ~new_P1_U7785 | ~new_P1_U7784;
  assign new_P1_U7491 = ~new_P1_U4108 | ~new_P1_U7216;
  assign new_P1_U7492 = ~new_P1_U4109 | ~new_P1_U7094;
  assign new_P1_U7493 = ~new_P1_U3279;
  assign new_P1_U7494 = ~new_P1_U3276;
  assign new_P1_U7495 = ~new_P1_U4068 | ~new_P1_U4069 | ~new_P1_U4070 | ~new_P1_U4071 | ~new_P1_U2607;
  assign new_P1_U7496 = ~new_P1_U3734 | ~new_P1_U7493;
  assign new_P1_U7497 = ~new_P1_U3735 | ~new_P1_U5469;
  assign new_P1_U7498 = ~new_P1_U2425 | ~new_P1_U7493;
  assign new_P1_U7499 = ~new_P1_U2425 | ~new_P1_U7493;
  assign new_P1_U7500 = ~new_P1_U7499 | ~new_P1_U6361 | ~new_P1_U6360;
  assign new_P1_U7501 = ~new_P1_U7493 | ~new_P1_R2167_U17;
  assign new_P1_U7502 = ~new_P1_R2167_U17 | ~new_P1_U7493 | ~new_P1_U4201;
  assign new_P1_U7503 = ~new_P1_U7502 | ~new_P1_U6149;
  assign new_P1_U7504 = ~new_P1_U7493 | ~new_P1_U7085;
  assign new_P1_U7505 = ~new_P1_U7493 | ~new_P1_U7471;
  assign new_P1_U7506 = ~new_P1_U4114 | ~new_P1_U4116 | ~new_P1_U4115;
  assign new_P1_U7507 = ~new_P1_U3759 | ~new_P1_U7493;
  assign new_P1_U7508 = ~new_P1_U3760 | ~new_P1_U3761 | ~new_P1_U5565;
  assign new_P1_U7509 = ~new_P1_U3746 | ~new_P1_U2519;
  assign new_P1_U7510 = ~new_P1_U7493 | ~new_P1_U5962;
  assign new_P1_U7511 = ~new_P1_U7493 | ~new_P1_U5965;
  assign new_P1_U7512 = ~new_P1_U7493 | ~new_P1_U5968;
  assign new_P1_U7513 = ~new_P1_U7493 | ~new_P1_U5971;
  assign new_P1_U7514 = ~new_P1_U7493 | ~new_P1_U5974;
  assign new_P1_U7515 = ~new_P1_U7493 | ~new_P1_U5977;
  assign new_P1_U7516 = ~new_P1_U7493 | ~new_P1_U5980;
  assign new_P1_U7517 = ~new_P1_U7493 | ~new_P1_U5983;
  assign new_P1_U7518 = ~new_P1_U7493 | ~new_P1_U5986;
  assign new_P1_U7519 = ~new_P1_U7493 | ~new_P1_U5989;
  assign new_P1_U7520 = ~new_P1_U7493 | ~new_P1_U5992;
  assign new_P1_U7521 = ~new_P1_U7493 | ~new_P1_U5995;
  assign new_P1_U7522 = ~new_P1_U7493 | ~new_P1_U5998;
  assign new_P1_U7523 = ~new_P1_U7493 | ~new_P1_U6001;
  assign new_P1_U7524 = ~new_P1_U7493 | ~new_P1_U6004;
  assign new_P1_U7525 = ~new_P1_U7493 | ~new_P1_U6007;
  assign new_P1_U7526 = ~new_P1_U7493 | ~new_P1_U6010;
  assign new_P1_U7527 = ~new_P1_U7493 | ~new_P1_U6013;
  assign new_P1_U7528 = ~new_P1_U7493 | ~new_P1_U6016;
  assign new_P1_U7529 = ~new_P1_U7493 | ~new_P1_U6019;
  assign new_P1_U7530 = ~new_P1_U7493 | ~new_P1_U6022;
  assign new_P1_U7531 = ~new_P1_U7493 | ~new_P1_U6025;
  assign new_P1_U7532 = ~new_P1_U7493 | ~new_P1_U6028;
  assign new_P1_U7533 = ~new_P1_U7493 | ~new_P1_U6031;
  assign new_P1_U7534 = ~new_P1_U7493 | ~new_P1_U6034;
  assign new_P1_U7535 = ~new_P1_U7493 | ~new_P1_U6037;
  assign new_P1_U7536 = ~new_P1_U7493 | ~new_P1_U6040;
  assign new_P1_U7537 = ~new_P1_U7493 | ~new_P1_U6043;
  assign new_P1_U7538 = ~new_P1_U7493 | ~new_P1_U6046;
  assign new_P1_U7539 = ~new_P1_U7493 | ~new_P1_U6049;
  assign new_P1_U7540 = ~new_P1_U7493 | ~new_P1_U6052;
  assign new_P1_U7541 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7542 = ~P1_UWORD_REG_0_ | ~new_P1_U7541;
  assign new_P1_U7543 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7544 = ~P1_UWORD_REG_1_ | ~new_P1_U7543;
  assign new_P1_U7545 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7546 = ~P1_UWORD_REG_2_ | ~new_P1_U7545;
  assign new_P1_U7547 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7548 = ~P1_UWORD_REG_3_ | ~new_P1_U7547;
  assign new_P1_U7549 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7550 = ~P1_UWORD_REG_4_ | ~new_P1_U7549;
  assign new_P1_U7551 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7552 = ~P1_UWORD_REG_5_ | ~new_P1_U7551;
  assign new_P1_U7553 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7554 = ~P1_UWORD_REG_6_ | ~new_P1_U7553;
  assign new_P1_U7555 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7556 = ~P1_UWORD_REG_7_ | ~new_P1_U7555;
  assign new_P1_U7557 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7558 = ~P1_UWORD_REG_8_ | ~new_P1_U7557;
  assign new_P1_U7559 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7560 = ~P1_UWORD_REG_9_ | ~new_P1_U7559;
  assign new_P1_U7561 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7562 = ~P1_UWORD_REG_10_ | ~new_P1_U7561;
  assign new_P1_U7563 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7564 = ~P1_UWORD_REG_11_ | ~new_P1_U7563;
  assign new_P1_U7565 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7566 = ~P1_UWORD_REG_12_ | ~new_P1_U7565;
  assign new_P1_U7567 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7568 = ~P1_UWORD_REG_13_ | ~new_P1_U7567;
  assign new_P1_U7569 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7570 = ~P1_UWORD_REG_14_ | ~new_P1_U7569;
  assign new_P1_U7571 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7572 = ~P1_LWORD_REG_0_ | ~new_P1_U7571;
  assign new_P1_U7573 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7574 = ~P1_LWORD_REG_1_ | ~new_P1_U7573;
  assign new_P1_U7575 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7576 = ~P1_LWORD_REG_2_ | ~new_P1_U7575;
  assign new_P1_U7577 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7578 = ~P1_LWORD_REG_3_ | ~new_P1_U7577;
  assign new_P1_U7579 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7580 = ~P1_LWORD_REG_4_ | ~new_P1_U7579;
  assign new_P1_U7581 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7582 = ~P1_LWORD_REG_5_ | ~new_P1_U7581;
  assign new_P1_U7583 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7584 = ~P1_LWORD_REG_6_ | ~new_P1_U7583;
  assign new_P1_U7585 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7586 = ~P1_LWORD_REG_7_ | ~new_P1_U7585;
  assign new_P1_U7587 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7588 = ~P1_LWORD_REG_8_ | ~new_P1_U7587;
  assign new_P1_U7589 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7590 = ~P1_LWORD_REG_9_ | ~new_P1_U7589;
  assign new_P1_U7591 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7592 = ~P1_LWORD_REG_10_ | ~new_P1_U7591;
  assign new_P1_U7593 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7594 = ~P1_LWORD_REG_11_ | ~new_P1_U7593;
  assign new_P1_U7595 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7596 = ~P1_LWORD_REG_12_ | ~new_P1_U7595;
  assign new_P1_U7597 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7598 = ~P1_LWORD_REG_13_ | ~new_P1_U7597;
  assign new_P1_U7599 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7600 = ~P1_LWORD_REG_14_ | ~new_P1_U7599;
  assign new_P1_U7601 = ~new_P1_U2357 | ~new_P1_U7493;
  assign new_P1_U7602 = ~P1_LWORD_REG_15_ | ~new_P1_U7601;
  assign new_P1_U7603 = ~new_P1_U4259 | ~new_P1_U7493 | ~new_P1_U3568;
  assign new_P1_U7604 = ~new_P1_U3581 | ~new_P1_U7684 | ~new_P1_U7683;
  assign new_P1_U7605 = ~new_P1_U3867 | ~new_P1_U7493;
  assign new_P1_U7606 = ~new_P1_U7605 | ~new_P1_U3428;
  assign new_P1_U7607 = ~new_P1_U4208 | ~new_P1_U7493;
  assign new_P1_U7608 = ~new_P1_U7607 | ~new_P1_U3447;
  assign new_P1_U7609 = ~new_P1_U3279 | ~new_P1_U3400;
  assign new_P1_U7610 = ~new_P1_U3754 | ~new_P1_U7493;
  assign new_P1_U7611 = ~new_P1_U3755 | ~new_P1_U7610;
  assign new_P1_U7612 = ~P1_INSTQUEUE_REG_0__4_ | ~new_P1_U5416;
  assign new_P1_U7613 = ~new_P1_U2523 | ~P1_INSTQUEUE_REG_0__4_;
  assign new_P1_U7614 = ~new_P1_U2546 | ~P1_INSTQUEUE_REG_0__4_;
  assign new_P1_U7615 = ~new_P1_U4049 | ~new_P1_U4050 | ~new_P1_U4052 | ~new_P1_U4051;
  assign new_P1_U7616 = ~new_P1_U4192 | ~P1_INSTQUEUE_REG_0__4_;
  assign new_P1_U7617 = ~new_P1_U2573 | ~P1_INSTQUEUE_REG_0__4_;
  assign new_P1_U7618 = ~new_P1_U4087 | ~new_P1_U4088 | ~new_P1_U4091 | ~new_P1_U4089;
  assign new_P1_U7619 = ~new_P1_U2592 | ~P1_INSTQUEUE_REG_0__4_;
  assign new_P1_U7620 = ~new_P1_U4133 | ~new_P1_U4134 | ~new_P1_U4136 | ~new_P1_U4135;
  assign new_P1_U7621 = ~new_P1_U3259;
  assign new_P1_U7622 = ~new_P1_U7621 | ~new_P1_U3261;
  assign new_P1_U7623 = ~new_P1_U4358 | ~new_P1_U4361 | ~P1_STATE_REG_1_;
  assign new_P1_U7624 = ~P1_STATE_REG_2_ | ~new_P1_U7468;
  assign new_P1_U7625 = ~P1_STATE_REG_1_ | ~new_P1_U4358;
  assign new_P1_U7626 = ~new_P1_U4502 | ~new_P1_U4510;
  assign new_P1_U7627 = ~new_P1_U5487 | ~new_P1_U4171;
  assign new_P1_U7628 = ~new_P1_U3283 | ~new_P1_U3289;
  assign new_P1_U7629 = ~new_P1_U3392;
  assign new_P1_U7630 = ~new_P1_U4208 | ~new_P1_U7490;
  assign new_P1_U7631 = ~new_P1_U5487 | ~new_P1_U4171;
  assign new_P1_U7632 = ~new_P1_U7631 | ~new_P1_U7630;
  assign new_P1_U7633 = ~P1_BE_N_REG_3_ | ~new_P1_U3249;
  assign new_P1_U7634 = ~P1_BYTEENABLE_REG_3_ | ~new_P1_U4221;
  assign new_P1_U7635 = ~P1_BE_N_REG_2_ | ~new_P1_U3249;
  assign new_P1_U7636 = ~P1_BYTEENABLE_REG_2_ | ~new_P1_U4221;
  assign new_P1_U7637 = ~P1_BE_N_REG_1_ | ~new_P1_U3249;
  assign new_P1_U7638 = ~P1_BYTEENABLE_REG_1_ | ~new_P1_U4221;
  assign new_P1_U7639 = ~P1_BE_N_REG_0_ | ~new_P1_U3249;
  assign new_P1_U7640 = ~P1_BYTEENABLE_REG_0_ | ~new_P1_U4221;
  assign new_P1_U7641 = ~new_P1_U3251 | ~P1_STATE_REG_0_ | ~P1_REQUESTPENDING_REG;
  assign new_P1_U7642 = ~P1_STATE_REG_2_ | ~new_P1_U3259;
  assign new_P1_U7643 = ~new_P1_U7642 | ~new_P1_U7641;
  assign new_P1_U7644 = ~P1_STATE_REG_1_ | ~new_P1_U7624 | ~new_P1_U4361;
  assign new_P1_U7645 = ~new_P1_U7643 | ~new_P1_U3248;
  assign new_P1_U7646 = ~P1_STATE_REG_2_ | ~P1_STATE_REG_0_ | ~new_P1_U3260;
  assign new_P1_U7647 = ~new_P1_U4371 | ~new_P1_U3251;
  assign new_P1_U7648 = P1_STATE_REG_0_ | P1_STATE_REG_1_;
  assign new_P1_U7649 = ~P1_STATE_REG_0_ | ~new_P1_U4258;
  assign new_P1_U7650 = ~new_P1_U3462;
  assign new_P1_U7651 = ~new_P1_U7650 | ~P1_DATAWIDTH_REG_0_;
  assign new_P1_U7652 = ~new_P1_U3463 | ~new_P1_U3462;
  assign new_P1_U7653 = ~new_P1_U3462 | ~new_P1_U4376;
  assign new_P1_U7654 = ~new_P1_U7650 | ~P1_DATAWIDTH_REG_1_;
  assign new_P1_U7655 = ~new_P1_U3265 | ~new_P1_U3541 | ~new_P1_U3540;
  assign new_P1_U7656 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3270 | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~P1_INSTQUEUE_REG_7__4_ | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7657 = ~new_P1_U3265 | ~new_P1_U3270 | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~P1_INSTQUEUE_REG_5__4_ | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7658 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3266 | ~new_P1_U3264 | ~P1_INSTQUEUE_REG_2__4_ | ~new_P1_U3270;
  assign new_P1_U7659 = ~new_P1_U3270 | ~new_P1_U3543 | ~new_P1_U3542;
  assign new_P1_U7660 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3545 | ~new_P1_U3544;
  assign new_P1_U7661 = ~new_P1_U3265 | ~new_P1_U3547 | ~new_P1_U3546;
  assign new_P1_U7662 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3549 | ~new_P1_U3548;
  assign new_P1_U7663 = ~new_P1_U3266 | ~new_P1_U3551 | ~new_P1_U3550;
  assign new_P1_U7664 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUERD_ADDR_REG_2_ | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_15__4_ | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7665 = ~new_P1_U3270 | ~new_P1_U3266 | ~new_P1_U3265 | ~P1_INSTQUEUE_REG_0__4_ | ~new_P1_U3264;
  assign new_P1_U7666 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3266 | ~new_P1_U3265 | ~P1_INSTQUEUE_REG_8__4_ | ~new_P1_U3264;
  assign new_P1_U7667 = ~new_P1_U3266 | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_10__4_ | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7668 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~new_P1_U3553 | ~new_P1_U3552;
  assign new_P1_U7669 = ~new_P1_U3270 | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_3__4_ | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7670 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_11__4_ | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7671 = ~new_P1_U3270 | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_3__5_ | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7672 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3529 | ~new_P1_U3528;
  assign new_P1_U7673 = ~new_P1_U3265 | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_0_ | ~P1_INSTQUEUE_REG_9__6_ | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7674 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3535 | ~new_P1_U3534;
  assign new_P1_U7675 = ~new_P1_U3266 | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_10__6_ | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7676 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~new_P1_U3264 | ~P1_INSTQUEUERD_ADDR_REG_1_ | ~P1_INSTQUEUE_REG_11__6_ | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7677 = ~new_P1_U3270 | ~new_P1_U3266 | ~new_P1_U3265 | ~P1_INSTQUEUE_REG_0__6_ | ~new_P1_U3264;
  assign new_P1_U7678 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U3266 | ~new_P1_U3265 | ~P1_INSTQUEUE_REG_8__6_ | ~new_P1_U3264;
  assign new_P1_U7679 = ~new_P1_U4494 | ~new_P1_U3437;
  assign new_P1_U7680 = ~new_P1_U7501 | ~new_P1_U3284;
  assign new_P1_U7681 = ~new_P1_U4216 | ~new_P1_R2167_U17;
  assign new_P1_U7682 = ~new_P1_U4506 | ~new_P1_U3273;
  assign new_P1_U7683 = ~P1_STATE2_REG_0_ | ~new_P1_U4512;
  assign new_P1_U7684 = ~new_P1_U4513 | ~new_P1_U3294;
  assign new_P1_U7685 = ~P1_STATE2_REG_3_ | ~new_P1_U3295;
  assign new_P1_U7686 = ~new_P1_U2428 | ~new_P1_U4514;
  assign new_P1_U7687 = P1_STATEBS16_REG | P1_STATE2_REG_0_;
  assign new_P1_U7688 = ~P1_STATE2_REG_0_ | ~new_P1_U7469;
  assign new_P1_U7689 = ~P1_STATE2_REG_0_ | ~new_P1_U4522;
  assign new_P1_U7690 = ~new_P1_U3294 | ~new_P1_U7604 | ~new_P1_U4521;
  assign new_P1_U7691 = ~new_P1_R2144_U49 | ~new_P1_U3313;
  assign new_P1_U7692 = ~new_P1_U4528 | ~new_P1_U3311;
  assign new_P1_U7693 = ~new_P1_U3454;
  assign new_P1_U7694 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_U3305;
  assign new_P1_U7695 = ~new_P1_U4533 | ~new_P1_U3304;
  assign new_P1_U7696 = ~new_P1_U3455;
  assign new_P1_U7697 = ~new_P1_U4216 | ~new_P1_U3273;
  assign new_P1_U7698 = ~new_P1_R2167_U17 | ~new_P1_U7497;
  assign new_P1_U7699 = ~new_P1_U4432 | ~new_P1_U5466;
  assign new_P1_U7700 = ~new_P1_U5467 | ~new_P1_U4171;
  assign new_P1_U7701 = ~new_P1_U3467 | ~new_P1_U4172;
  assign new_P1_U7702 = ~new_P1_U5476 | ~P1_INSTQUEUERD_ADDR_REG_4_;
  assign new_P1_U7703 = ~new_P1_U4460 | ~new_P1_U3278;
  assign new_P1_U7704 = ~new_P1_U4415 | ~new_P1_U3277;
  assign new_P1_U7705 = ~new_P1_U3271 | ~new_P1_U3415;
  assign new_P1_U7706 = ~new_P1_U4477 | ~new_P1_U5493;
  assign new_P1_U7707 = ~new_P1_U7706 | ~new_P1_U7705;
  assign new_P1_U7708 = ~new_P1_U5476 | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7709 = ~new_P1_U5509 | ~new_P1_U4172;
  assign new_P1_U7710 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_U4174;
  assign new_P1_U7711 = ~new_P1_SUB_580_U6 | ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_U7712 = ~new_P1_U3470;
  assign new_P1_U7713 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_U4174;
  assign new_P1_U7714 = ~P1_INSTADDRPOINTER_REG_0_ | ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_U7715 = ~new_P1_U3471;
  assign new_P1_U7716 = ~new_P1_U5511 | ~new_P1_U5501;
  assign new_P1_U7717 = ~new_P1_U4218 | ~new_P1_U3401;
  assign new_P1_U7718 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_U3264;
  assign new_P1_U7719 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_U3265;
  assign new_P1_U7720 = ~new_P1_U3456;
  assign new_P1_U7721 = ~new_P1_U5476 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U7722 = ~new_P1_U5518 | ~new_P1_U4172;
  assign new_P1_U7723 = ~new_P1_U5476 | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U7724 = ~new_P1_U5529 | ~new_P1_U4172;
  assign new_P1_U7725 = ~new_P1_U4214 | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7726 = ~new_P1_U5521 | ~new_P1_U3266;
  assign new_P1_U7727 = ~new_P1_U5476 | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7728 = ~new_P1_U5535 | ~new_P1_U4172;
  assign new_P1_U7729 = ~new_P1_U5537 | ~P1_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P1_U7730 = ~new_P1_U5545 | ~new_P1_U3404;
  assign new_P1_U7731 = ~new_P1_U7693 | ~new_P1_U4527;
  assign new_P1_U7732 = ~new_P1_U3454 | ~new_P1_U3314;
  assign new_P1_U7733 = ~new_P1_U7732 | ~new_P1_U7731;
  assign new_P1_U7734 = ~new_P1_U5537 | ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P1_U7735 = ~new_P1_U5549 | ~new_P1_U3404;
  assign new_P1_U7736 = ~new_P1_U5537 | ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P1_U7737 = ~new_P1_U5554 | ~new_P1_U3404;
  assign new_P1_U7738 = ~new_P1_U5537 | ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P1_U7739 = ~new_P1_U5557 | ~new_P1_U3404;
  assign new_P1_U7740 = ~new_P1_U4477 | ~new_P1_U3388;
  assign new_P1_U7741 = ~new_P1_U3271 | ~new_P1_U3281;
  assign new_P1_U7742 = ~new_P1_U4171 | ~new_P1_U3257 | ~new_P1_U7741 | ~new_P1_U7740;
  assign new_P1_U7743 = ~new_P1_U4432 | ~new_P1_R2167_U17 | ~new_P1_U7611;
  assign new_P1_U7744 = ~P1_EAX_REG_31_ | ~new_P1_U3424;
  assign new_P1_U7745 = ~new_P1_U3479 | ~new_P1_U4223;
  assign new_P1_U7746 = ~P1_BYTEENABLE_REG_3_ | ~new_P1_U3433;
  assign new_P1_U7747 = ~new_P1_U3480 | ~new_P1_U4220;
  assign new_P1_U7748 = P1_DATAWIDTH_REG_0_ | P1_DATAWIDTH_REG_1_;
  assign new_P1_U7749 = ~P1_DATAWIDTH_REG_0_ | ~new_P1_U3413;
  assign new_P1_U7750 = ~new_P1_U7749 | ~new_P1_U7748;
  assign new_P1_U7751 = ~new_P1_U7750 | ~new_P1_U3253;
  assign new_P1_U7752 = ~P1_REIP_REG_0_ | ~P1_REIP_REG_1_;
  assign new_P1_U7753 = ~new_P1_U7752 | ~new_P1_U7751;
  assign new_P1_U7754 = ~P1_BYTEENABLE_REG_2_ | ~new_P1_U3433;
  assign new_P1_U7755 = ~new_P1_U7753 | ~new_P1_U4220;
  assign new_P1_U7756 = ~P1_BYTEENABLE_REG_1_ | ~new_P1_U3433;
  assign new_P1_U7757 = ~new_P1_U4220 | ~P1_REIP_REG_1_;
  assign new_P1_U7758 = ~P1_BYTEENABLE_REG_0_ | ~new_P1_U3433;
  assign new_P1_U7759 = ~new_P1_U4220 | ~new_P1_U6599;
  assign new_P1_U7760 = ~new_P1_U4221 | ~new_P1_U3436;
  assign new_P1_U7761 = ~P1_W_R_N_REG | ~new_P1_U3249;
  assign new_P1_U7762 = ~P1_MORE_REG | ~new_P1_U4177;
  assign new_P1_U7763 = ~new_P1_U4237 | ~new_P1_U6600;
  assign new_P1_U7764 = ~new_P1_U7650 | ~P1_STATEBS16_REG;
  assign new_P1_U7765 = ~BS16 | ~new_P1_U3462;
  assign new_P1_U7766 = ~new_P1_U6603 | ~P1_REQUESTPENDING_REG;
  assign new_P1_U7767 = ~new_P1_U6609 | ~new_P1_U4180;
  assign new_P1_U7768 = ~new_P1_U4221 | ~new_P1_U3435;
  assign new_P1_U7769 = ~P1_D_C_N_REG | ~new_P1_U3249;
  assign new_P1_U7770 = ~P1_M_IO_N_REG | ~new_P1_U3249;
  assign new_P1_U7771 = ~P1_MEMORYFETCH_REG | ~new_P1_U4221;
  assign new_P1_U7772 = ~new_P1_U6614 | ~P1_READREQUEST_REG;
  assign new_P1_U7773 = ~new_P1_U6615 | ~new_P1_U4181;
  assign new_P1_U7774 = ~new_P1_U3488 | ~new_P1_U4182;
  assign new_P1_U7775 = ~new_P1_U5473 | ~P1_INSTQUEUERD_ADDR_REG_4_;
  assign new_P1_U7776 = ~new_P1_U5473 | ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_U7777 = ~new_P1_U5506 | ~new_P1_U4182;
  assign new_P1_U7778 = ~new_P1_U5473 | ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_U7779 = ~new_P1_U5514 | ~new_P1_U4182;
  assign new_P1_U7780 = ~new_P1_U5473 | ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_U7781 = ~new_P1_U5525 | ~new_P1_U4182;
  assign new_P1_U7782 = ~new_P1_U5473 | ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_U7783 = ~new_P1_U5531 | ~new_P1_U4182;
  assign new_P1_U7784 = ~new_P1_U2605 | ~new_P1_U3277;
  assign new_P1_U7785 = ~new_P1_U4460 | ~new_P1_U7495;
  assign new_P1_U7786 = ~new_P1_U4203 | ~new_P1_U3301;
  assign new_P1_U7787 = ~P1_INSTQUEUEWR_ADDR_REG_0_ | ~new_P1_U3297;
  assign new_P1_U7788 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_U4183;
  assign new_P1_U7789 = ~new_P1_U7219 | ~new_P1_U3270;
  assign new_P1_U7790 = ~new_P1_U3457;
  assign new_P1_U7791 = ~new_P1_U3276 | ~new_P1_U3284;
  assign new_P1_U7792 = ~new_P1_U7707 | ~new_P1_U4494;
  assign new_P1_U7793 = ~new_P1_U3493 | ~new_P1_U3262;
  assign new_P1_U7794 = ~P1_STATE2_REG_1_ | ~P1_FLUSH_REG | ~new_P1_U7715;
  assign new_P1_ADD_405_U113 = ~new_P1_ADD_405_U38;
  assign new_P1_ADD_405_U112 = ~new_P1_ADD_405_U36;
  assign new_P1_ADD_405_U111 = ~new_P1_ADD_405_U34;
  assign new_P1_ADD_405_U110 = ~new_P1_ADD_405_U32;
  assign new_P1_ADD_405_U109 = ~new_P1_ADD_405_U30;
  assign new_P1_ADD_405_U108 = ~new_P1_ADD_405_U28;
  assign new_P1_ADD_405_U107 = ~new_P1_ADD_405_U26;
  assign new_P1_ADD_405_U106 = ~new_P1_ADD_405_U24;
  assign new_P1_ADD_405_U105 = ~new_P1_ADD_405_U22;
  assign new_P1_ADD_405_U104 = ~new_P1_ADD_405_U20;
  assign new_P1_ADD_405_U103 = ~new_P1_ADD_405_U18;
  assign new_P1_ADD_405_U102 = ~new_P1_ADD_405_U16;
  assign new_P1_ADD_405_U101 = ~new_P1_ADD_405_U14;
  assign new_P1_ADD_405_U100 = ~new_P1_ADD_405_U13;
  assign new_P1_ADD_405_U99 = ~new_P1_ADD_405_U10;
  assign new_P1_ADD_405_U98 = ~new_P1_ADD_405_U8;
  assign new_P1_ADD_405_U97 = ~new_P1_ADD_405_U94;
  assign new_P1_ADD_405_U96 = ~P1_INSTADDRPOINTER_REG_1_ | ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_ADD_405_U95 = new_P1_ADD_405_U172 & new_P1_ADD_405_U171;
  assign new_P1_ADD_405_U94 = ~new_P1_ADD_405_U62 | ~new_P1_ADD_405_U96;
  assign new_P1_ADD_405_U93 = ~new_P1_ADD_405_U124 | ~P1_INSTADDRPOINTER_REG_30_;
  assign new_P1_ADD_405_U92 = ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_ADD_405_U91 = ~new_P1_ADD_405_U186 | ~new_P1_ADD_405_U185;
  assign new_P1_ADD_405_U90 = ~new_P1_ADD_405_U184 | ~new_P1_ADD_405_U183;
  assign new_P1_ADD_405_U89 = ~new_P1_ADD_405_U182 | ~new_P1_ADD_405_U181;
  assign new_P1_ADD_405_U88 = ~new_P1_ADD_405_U180 | ~new_P1_ADD_405_U179;
  assign new_P1_ADD_405_U87 = ~new_P1_ADD_405_U178 | ~new_P1_ADD_405_U177;
  assign new_LT_782_120_U6 = ~P3_DATAO_REG_30_ | ~new_LT_782_120_U7;
  assign new_LT_782_120_U7 = ~P3_DATAO_REG_31_;
  assign new_LT_782_U6 = ~P1_DATAO_REG_30_ | ~new_LT_782_U7;
  assign new_LT_782_U7 = ~P1_DATAO_REG_31_;
  assign new_LT_748_U6 = ~P2_ADDRESS_REG_29_;
  assign new_R170_U6 = P2_ADDRESS_REG_29_ & new_R170_U15;
  assign new_R170_U7 = P2_ADDRESS_REG_22_ | P2_ADDRESS_REG_7_ | P2_ADDRESS_REG_17_ | P2_ADDRESS_REG_9_;
  assign new_R170_U8 = ~P2_ADDRESS_REG_24_ & ~P2_ADDRESS_REG_25_ & ~P2_ADDRESS_REG_19_ & ~new_R170_U7 & ~P2_ADDRESS_REG_10_;
  assign new_R170_U9 = P2_ADDRESS_REG_8_ | P2_ADDRESS_REG_18_ | P2_ADDRESS_REG_16_ | P2_ADDRESS_REG_0_;
  assign new_R170_U10 = ~P2_ADDRESS_REG_11_ & ~P2_ADDRESS_REG_1_ & ~new_R170_U9 & ~P2_ADDRESS_REG_23_;
  assign new_R170_U11 = P2_ADDRESS_REG_6_ | P2_ADDRESS_REG_28_ | P2_ADDRESS_REG_26_ | P2_ADDRESS_REG_21_;
  assign new_R170_U12 = ~P2_ADDRESS_REG_4_ & ~P2_ADDRESS_REG_14_ & ~new_R170_U11 & ~P2_ADDRESS_REG_12_;
  assign new_R170_U13 = P2_ADDRESS_REG_27_ | P2_ADDRESS_REG_3_ | P2_ADDRESS_REG_13_ | P2_ADDRESS_REG_20_;
  assign new_R170_U14 = ~P2_ADDRESS_REG_15_ & ~P2_ADDRESS_REG_5_ & ~new_R170_U13 & ~P2_ADDRESS_REG_2_;
  assign new_R170_U15 = ~new_R170_U8 | ~new_R170_U10 | ~new_R170_U14 | ~new_R170_U12;
  assign new_R165_U6 = P1_ADDRESS_REG_29_ & new_R165_U15;
  assign new_R165_U7 = P1_ADDRESS_REG_22_ | P1_ADDRESS_REG_7_ | P1_ADDRESS_REG_17_ | P1_ADDRESS_REG_9_;
  assign new_R165_U8 = ~P1_ADDRESS_REG_24_ & ~P1_ADDRESS_REG_25_ & ~P1_ADDRESS_REG_19_ & ~new_R165_U7 & ~P1_ADDRESS_REG_10_;
  assign new_R165_U9 = P1_ADDRESS_REG_8_ | P1_ADDRESS_REG_18_ | P1_ADDRESS_REG_16_ | P1_ADDRESS_REG_0_;
  assign new_R165_U10 = ~P1_ADDRESS_REG_11_ & ~P1_ADDRESS_REG_1_ & ~new_R165_U9 & ~P1_ADDRESS_REG_23_;
  assign new_R165_U11 = P1_ADDRESS_REG_6_ | P1_ADDRESS_REG_28_ | P1_ADDRESS_REG_26_ | P1_ADDRESS_REG_21_;
  assign new_R165_U12 = ~P1_ADDRESS_REG_4_ & ~P1_ADDRESS_REG_14_ & ~new_R165_U11 & ~P1_ADDRESS_REG_12_;
  assign new_R165_U13 = P1_ADDRESS_REG_27_ | P1_ADDRESS_REG_3_ | P1_ADDRESS_REG_13_ | P1_ADDRESS_REG_20_;
  assign new_R165_U14 = ~P1_ADDRESS_REG_15_ & ~P1_ADDRESS_REG_5_ & ~new_R165_U13 & ~P1_ADDRESS_REG_2_;
  assign new_R165_U15 = ~new_R165_U8 | ~new_R165_U10 | ~new_R165_U14 | ~new_R165_U12;
  assign new_LT_782_119_U6 = ~P2_DATAO_REG_30_ | ~new_LT_782_119_U7;
  assign new_LT_782_119_U7 = ~P2_DATAO_REG_31_;
  assign new_P3_ADD_526_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_526_U6 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_526_U7 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_526_U8 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_526_U9 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_526_U10 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_526_U11 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_526_U12 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_526_U13 = ~new_P3_ADD_526_U82 | ~new_P3_ADD_526_U111;
  assign new_P3_ADD_526_U14 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_526_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_526_U16 = ~new_P3_ADD_526_U83 | ~new_P3_ADD_526_U112;
  assign new_P3_ADD_526_U17 = ~new_P3_ADD_526_U84 | ~new_P3_ADD_526_U118;
  assign new_P3_ADD_526_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_526_U19 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_526_U20 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_526_U21 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_526_U22 = ~new_P3_ADD_526_U85 | ~new_P3_ADD_526_U120;
  assign new_P3_ADD_526_U23 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_526_U24 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_526_U25 = ~new_P3_ADD_526_U86 | ~new_P3_ADD_526_U113;
  assign new_P3_ADD_526_U26 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_526_U27 = ~new_P3_ADD_526_U87 | ~new_P3_ADD_526_U119;
  assign new_P3_ADD_526_U28 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_526_U29 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_526_U30 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_526_U31 = ~new_P3_ADD_526_U88 | ~new_P3_ADD_526_U124;
  assign new_P3_ADD_526_U32 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_526_U33 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_526_U34 = ~new_P3_ADD_526_U89 | ~new_P3_ADD_526_U117;
  assign new_P3_ADD_526_U35 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_526_U36 = ~new_P3_ADD_526_U90 | ~new_P3_ADD_526_U114;
  assign new_P3_ADD_526_U37 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_526_U38 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_526_U39 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_526_U40 = ~new_P3_ADD_526_U91 | ~new_P3_ADD_526_U121;
  assign new_P3_ADD_526_U41 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_526_U42 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_526_U43 = ~new_P3_ADD_526_U92 | ~new_P3_ADD_526_U115;
  assign new_P3_ADD_526_U44 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_526_U45 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_526_U46 = ~new_P3_ADD_526_U93 | ~new_P3_ADD_526_U116;
  assign new_P3_ADD_526_U47 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_526_U48 = ~new_P3_ADD_526_U94 | ~new_P3_ADD_526_U122;
  assign new_P3_ADD_526_U49 = ~new_P3_ADD_526_U123 | ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_526_U50 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_526_U51 = ~new_P3_ADD_526_U142 | ~new_P3_ADD_526_U141;
  assign new_P3_ADD_526_U52 = ~new_P3_ADD_526_U144 | ~new_P3_ADD_526_U143;
  assign new_P3_ADD_526_U53 = ~new_P3_ADD_526_U146 | ~new_P3_ADD_526_U145;
  assign new_P3_ADD_526_U54 = ~new_P3_ADD_526_U148 | ~new_P3_ADD_526_U147;
  assign new_P3_ADD_526_U55 = ~new_P3_ADD_526_U150 | ~new_P3_ADD_526_U149;
  assign new_P3_ADD_526_U56 = ~new_P3_ADD_526_U152 | ~new_P3_ADD_526_U151;
  assign new_P3_ADD_526_U57 = ~new_P3_ADD_526_U154 | ~new_P3_ADD_526_U153;
  assign new_P3_ADD_526_U58 = ~new_P3_ADD_526_U156 | ~new_P3_ADD_526_U155;
  assign new_P3_ADD_526_U59 = ~new_P3_ADD_526_U158 | ~new_P3_ADD_526_U157;
  assign new_P3_ADD_526_U60 = ~new_P3_ADD_526_U160 | ~new_P3_ADD_526_U159;
  assign new_P3_ADD_526_U61 = ~new_P3_ADD_526_U162 | ~new_P3_ADD_526_U161;
  assign new_P3_ADD_526_U62 = ~new_P3_ADD_526_U164 | ~new_P3_ADD_526_U163;
  assign new_P3_ADD_526_U63 = ~new_P3_ADD_526_U166 | ~new_P3_ADD_526_U165;
  assign new_P3_ADD_526_U64 = ~new_P3_ADD_526_U168 | ~new_P3_ADD_526_U167;
  assign new_P3_ADD_526_U65 = ~new_P3_ADD_526_U170 | ~new_P3_ADD_526_U169;
  assign new_P3_ADD_526_U66 = ~new_P3_ADD_526_U172 | ~new_P3_ADD_526_U171;
  assign new_P3_ADD_526_U67 = ~new_P3_ADD_526_U174 | ~new_P3_ADD_526_U173;
  assign new_P3_ADD_526_U68 = ~new_P3_ADD_526_U176 | ~new_P3_ADD_526_U175;
  assign new_P3_ADD_526_U69 = ~new_P3_ADD_526_U178 | ~new_P3_ADD_526_U177;
  assign new_P3_ADD_526_U70 = ~new_P3_ADD_526_U180 | ~new_P3_ADD_526_U179;
  assign new_P3_ADD_526_U71 = ~new_P3_ADD_526_U182 | ~new_P3_ADD_526_U181;
  assign new_P3_ADD_526_U72 = ~new_P3_ADD_526_U184 | ~new_P3_ADD_526_U183;
  assign new_P3_ADD_526_U73 = ~new_P3_ADD_526_U186 | ~new_P3_ADD_526_U185;
  assign new_P3_ADD_526_U74 = ~new_P3_ADD_526_U188 | ~new_P3_ADD_526_U187;
  assign new_P3_ADD_526_U75 = ~new_P3_ADD_526_U190 | ~new_P3_ADD_526_U189;
  assign new_P3_ADD_526_U76 = ~new_P3_ADD_526_U192 | ~new_P3_ADD_526_U191;
  assign new_P3_ADD_526_U77 = ~new_P3_ADD_526_U194 | ~new_P3_ADD_526_U193;
  assign new_P3_ADD_526_U78 = ~new_P3_ADD_526_U196 | ~new_P3_ADD_526_U195;
  assign new_P3_ADD_526_U79 = ~new_P3_ADD_526_U198 | ~new_P3_ADD_526_U197;
  assign new_P3_ADD_526_U80 = ~new_P3_ADD_526_U200 | ~new_P3_ADD_526_U199;
  assign new_P3_ADD_526_U81 = ~new_P3_ADD_526_U202 | ~new_P3_ADD_526_U201;
  assign new_P3_ADD_526_U82 = P3_INSTADDRPOINTER_REG_3_ & P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_526_U83 = P3_INSTADDRPOINTER_REG_5_ & P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_526_U84 = P3_INSTADDRPOINTER_REG_7_ & P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_526_U85 = P3_INSTADDRPOINTER_REG_9_ & P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_526_U86 = P3_INSTADDRPOINTER_REG_11_ & P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_526_U87 = P3_INSTADDRPOINTER_REG_13_ & P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_526_U88 = P3_INSTADDRPOINTER_REG_16_ & P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_526_U89 = P3_INSTADDRPOINTER_REG_17_ & P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_526_U90 = P3_INSTADDRPOINTER_REG_19_ & P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_526_U91 = P3_INSTADDRPOINTER_REG_22_ & P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_526_U92 = P3_INSTADDRPOINTER_REG_23_ & P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_526_U93 = P3_INSTADDRPOINTER_REG_25_ & P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_526_U94 = P3_INSTADDRPOINTER_REG_28_ & P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_526_U95 = ~new_P3_ADD_526_U118 | ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_526_U96 = ~new_P3_ADD_526_U112 | ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_526_U97 = ~new_P3_ADD_526_U111 | ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_526_U98 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_526_U99 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_526_U128;
  assign new_P3_ADD_526_U100 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_526_U101 = ~new_P3_ADD_526_U122 | ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_526_U102 = ~new_P3_ADD_526_U116 | ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_526_U103 = ~new_P3_ADD_526_U115 | ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_526_U104 = ~new_P3_ADD_526_U121 | ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_526_U105 = ~new_P3_ADD_526_U114 | ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_526_U106 = ~new_P3_ADD_526_U117 | ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_526_U107 = ~new_P3_ADD_526_U124 | ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_526_U108 = ~new_P3_ADD_526_U119 | ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_526_U109 = ~new_P3_ADD_526_U113 | ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_526_U110 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_526_U120;
  assign new_P3_ADD_526_U111 = ~new_P3_ADD_526_U10;
  assign new_P3_ADD_526_U112 = ~new_P3_ADD_526_U13;
  assign new_P3_ADD_526_U113 = ~new_P3_ADD_526_U22;
  assign new_P3_ADD_526_U114 = ~new_P3_ADD_526_U34;
  assign new_P3_ADD_526_U115 = ~new_P3_ADD_526_U40;
  assign new_P3_ADD_526_U116 = ~new_P3_ADD_526_U43;
  assign new_P3_ADD_526_U117 = ~new_P3_ADD_526_U31;
  assign new_P3_ADD_526_U118 = ~new_P3_ADD_526_U16;
  assign new_P3_ADD_526_U119 = ~new_P3_ADD_526_U25;
  assign new_P3_ADD_526_U120 = ~new_P3_ADD_526_U17;
  assign new_P3_ADD_526_U121 = ~new_P3_ADD_526_U36;
  assign new_P3_ADD_526_U122 = ~new_P3_ADD_526_U46;
  assign new_P3_ADD_526_U123 = ~new_P3_ADD_526_U48;
  assign new_P3_ADD_526_U124 = ~new_P3_ADD_526_U27;
  assign new_P3_ADD_526_U125 = ~new_P3_ADD_526_U95;
  assign new_P3_ADD_526_U126 = ~new_P3_ADD_526_U96;
  assign new_P3_ADD_526_U127 = ~new_P3_ADD_526_U97;
  assign new_P3_ADD_526_U128 = ~new_P3_ADD_526_U49;
  assign new_P3_ADD_526_U129 = ~new_P3_ADD_526_U99;
  assign new_P3_ADD_526_U130 = ~new_P3_ADD_526_U100;
  assign new_P3_ADD_526_U131 = ~new_P3_ADD_526_U101;
  assign new_P3_ADD_526_U132 = ~new_P3_ADD_526_U102;
  assign new_P3_ADD_526_U133 = ~new_P3_ADD_526_U103;
  assign new_P3_ADD_526_U134 = ~new_P3_ADD_526_U104;
  assign new_P3_ADD_526_U135 = ~new_P3_ADD_526_U105;
  assign new_P3_ADD_526_U136 = ~new_P3_ADD_526_U106;
  assign new_P3_ADD_526_U137 = ~new_P3_ADD_526_U107;
  assign new_P3_ADD_526_U138 = ~new_P3_ADD_526_U108;
  assign new_P3_ADD_526_U139 = ~new_P3_ADD_526_U109;
  assign new_P3_ADD_526_U140 = ~new_P3_ADD_526_U110;
  assign new_P3_ADD_526_U141 = ~new_P3_ADD_526_U120 | ~new_P3_ADD_526_U18;
  assign new_P3_ADD_526_U142 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_526_U17;
  assign new_P3_ADD_526_U143 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_526_U95;
  assign new_P3_ADD_526_U144 = ~new_P3_ADD_526_U125 | ~new_P3_ADD_526_U14;
  assign new_P3_ADD_526_U145 = ~new_P3_ADD_526_U118 | ~new_P3_ADD_526_U15;
  assign new_P3_ADD_526_U146 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_526_U16;
  assign new_P3_ADD_526_U147 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_526_U96;
  assign new_P3_ADD_526_U148 = ~new_P3_ADD_526_U126 | ~new_P3_ADD_526_U11;
  assign new_P3_ADD_526_U149 = ~new_P3_ADD_526_U112 | ~new_P3_ADD_526_U12;
  assign new_P3_ADD_526_U150 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_526_U13;
  assign new_P3_ADD_526_U151 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_526_U97;
  assign new_P3_ADD_526_U152 = ~new_P3_ADD_526_U127 | ~new_P3_ADD_526_U8;
  assign new_P3_ADD_526_U153 = ~new_P3_ADD_526_U111 | ~new_P3_ADD_526_U9;
  assign new_P3_ADD_526_U154 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_526_U10;
  assign new_P3_ADD_526_U155 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_526_U99;
  assign new_P3_ADD_526_U156 = ~new_P3_ADD_526_U129 | ~new_P3_ADD_526_U98;
  assign new_P3_ADD_526_U157 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_526_U49;
  assign new_P3_ADD_526_U158 = ~new_P3_ADD_526_U128 | ~new_P3_ADD_526_U50;
  assign new_P3_ADD_526_U159 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_526_U100;
  assign new_P3_ADD_526_U160 = ~new_P3_ADD_526_U130 | ~new_P3_ADD_526_U6;
  assign new_P3_ADD_526_U161 = ~new_P3_ADD_526_U123 | ~new_P3_ADD_526_U47;
  assign new_P3_ADD_526_U162 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_526_U48;
  assign new_P3_ADD_526_U163 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_526_U101;
  assign new_P3_ADD_526_U164 = ~new_P3_ADD_526_U131 | ~new_P3_ADD_526_U45;
  assign new_P3_ADD_526_U165 = ~new_P3_ADD_526_U122 | ~new_P3_ADD_526_U44;
  assign new_P3_ADD_526_U166 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_526_U46;
  assign new_P3_ADD_526_U167 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_526_U102;
  assign new_P3_ADD_526_U168 = ~new_P3_ADD_526_U132 | ~new_P3_ADD_526_U41;
  assign new_P3_ADD_526_U169 = ~new_P3_ADD_526_U116 | ~new_P3_ADD_526_U42;
  assign new_P3_ADD_526_U170 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_526_U43;
  assign new_P3_ADD_526_U171 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_526_U103;
  assign new_P3_ADD_526_U172 = ~new_P3_ADD_526_U133 | ~new_P3_ADD_526_U38;
  assign new_P3_ADD_526_U173 = ~new_P3_ADD_526_U115 | ~new_P3_ADD_526_U39;
  assign new_P3_ADD_526_U174 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_526_U40;
  assign new_P3_ADD_526_U175 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_526_U104;
  assign new_P3_ADD_526_U176 = ~new_P3_ADD_526_U134 | ~new_P3_ADD_526_U37;
  assign new_P3_ADD_526_U177 = ~new_P3_ADD_526_U121 | ~new_P3_ADD_526_U35;
  assign new_P3_ADD_526_U178 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_526_U36;
  assign new_P3_ADD_526_U179 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_526_U105;
  assign new_P3_ADD_526_U180 = ~new_P3_ADD_526_U135 | ~new_P3_ADD_526_U32;
  assign new_P3_ADD_526_U181 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_526_U7;
  assign new_P3_ADD_526_U182 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_526_U5;
  assign new_P3_ADD_526_U183 = ~new_P3_ADD_526_U114 | ~new_P3_ADD_526_U33;
  assign new_P3_ADD_526_U184 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_526_U34;
  assign new_P3_ADD_526_U185 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_526_U106;
  assign new_P3_ADD_526_U186 = ~new_P3_ADD_526_U136 | ~new_P3_ADD_526_U29;
  assign new_P3_ADD_526_U187 = ~new_P3_ADD_526_U117 | ~new_P3_ADD_526_U30;
  assign new_P3_ADD_526_U188 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_526_U31;
  assign new_P3_ADD_526_U189 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_526_U107;
  assign new_P3_ADD_526_U190 = ~new_P3_ADD_526_U137 | ~new_P3_ADD_526_U28;
  assign new_P3_ADD_526_U191 = ~new_P3_ADD_526_U124 | ~new_P3_ADD_526_U26;
  assign new_P3_ADD_526_U192 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_526_U27;
  assign new_P3_ADD_526_U193 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_526_U108;
  assign new_P3_ADD_526_U194 = ~new_P3_ADD_526_U138 | ~new_P3_ADD_526_U23;
  assign new_P3_ADD_526_U195 = ~new_P3_ADD_526_U119 | ~new_P3_ADD_526_U24;
  assign new_P3_ADD_526_U196 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_526_U25;
  assign new_P3_ADD_526_U197 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_526_U109;
  assign new_P3_ADD_526_U198 = ~new_P3_ADD_526_U139 | ~new_P3_ADD_526_U20;
  assign new_P3_ADD_526_U199 = ~new_P3_ADD_526_U113 | ~new_P3_ADD_526_U21;
  assign new_P3_ADD_526_U200 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_526_U22;
  assign new_P3_ADD_526_U201 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_526_U110;
  assign new_P3_ADD_526_U202 = ~new_P3_ADD_526_U140 | ~new_P3_ADD_526_U19;
  assign new_P3_ADD_552_U5 = ~P3_EBX_REG_0_;
  assign new_P3_ADD_552_U6 = ~P3_EBX_REG_2_;
  assign new_P3_ADD_552_U7 = ~P3_EBX_REG_1_;
  assign new_P3_ADD_552_U8 = ~P3_EBX_REG_4_;
  assign new_P3_ADD_552_U9 = ~P3_EBX_REG_3_;
  assign new_P3_ADD_552_U10 = ~P3_EBX_REG_1_ | ~P3_EBX_REG_2_ | ~P3_EBX_REG_0_;
  assign new_P3_ADD_552_U11 = ~P3_EBX_REG_6_;
  assign new_P3_ADD_552_U12 = ~P3_EBX_REG_5_;
  assign new_P3_ADD_552_U13 = ~new_P3_ADD_552_U82 | ~new_P3_ADD_552_U111;
  assign new_P3_ADD_552_U14 = ~P3_EBX_REG_8_;
  assign new_P3_ADD_552_U15 = ~P3_EBX_REG_7_;
  assign new_P3_ADD_552_U16 = ~new_P3_ADD_552_U83 | ~new_P3_ADD_552_U112;
  assign new_P3_ADD_552_U17 = ~new_P3_ADD_552_U84 | ~new_P3_ADD_552_U118;
  assign new_P3_ADD_552_U18 = ~P3_EBX_REG_9_;
  assign new_P3_ADD_552_U19 = ~P3_EBX_REG_10_;
  assign new_P3_ADD_552_U20 = ~P3_EBX_REG_12_;
  assign new_P3_ADD_552_U21 = ~P3_EBX_REG_11_;
  assign new_P3_ADD_552_U22 = ~new_P3_ADD_552_U85 | ~new_P3_ADD_552_U120;
  assign new_P3_ADD_552_U23 = ~P3_EBX_REG_14_;
  assign new_P3_ADD_552_U24 = ~P3_EBX_REG_13_;
  assign new_P3_ADD_552_U25 = ~new_P3_ADD_552_U86 | ~new_P3_ADD_552_U113;
  assign new_P3_ADD_552_U26 = ~P3_EBX_REG_15_;
  assign new_P3_ADD_552_U27 = ~new_P3_ADD_552_U87 | ~new_P3_ADD_552_U119;
  assign new_P3_ADD_552_U28 = ~P3_EBX_REG_16_;
  assign new_P3_ADD_552_U29 = ~P3_EBX_REG_18_;
  assign new_P3_ADD_552_U30 = ~P3_EBX_REG_17_;
  assign new_P3_ADD_552_U31 = ~new_P3_ADD_552_U88 | ~new_P3_ADD_552_U124;
  assign new_P3_ADD_552_U32 = ~P3_EBX_REG_20_;
  assign new_P3_ADD_552_U33 = ~P3_EBX_REG_19_;
  assign new_P3_ADD_552_U34 = ~new_P3_ADD_552_U89 | ~new_P3_ADD_552_U117;
  assign new_P3_ADD_552_U35 = ~P3_EBX_REG_21_;
  assign new_P3_ADD_552_U36 = ~new_P3_ADD_552_U90 | ~new_P3_ADD_552_U114;
  assign new_P3_ADD_552_U37 = ~P3_EBX_REG_22_;
  assign new_P3_ADD_552_U38 = ~P3_EBX_REG_24_;
  assign new_P3_ADD_552_U39 = ~P3_EBX_REG_23_;
  assign new_P3_ADD_552_U40 = ~new_P3_ADD_552_U91 | ~new_P3_ADD_552_U121;
  assign new_P3_ADD_552_U41 = ~P3_EBX_REG_26_;
  assign new_P3_ADD_552_U42 = ~P3_EBX_REG_25_;
  assign new_P3_ADD_552_U43 = ~new_P3_ADD_552_U92 | ~new_P3_ADD_552_U115;
  assign new_P3_ADD_552_U44 = ~P3_EBX_REG_27_;
  assign new_P3_ADD_552_U45 = ~P3_EBX_REG_28_;
  assign new_P3_ADD_552_U46 = ~new_P3_ADD_552_U93 | ~new_P3_ADD_552_U116;
  assign new_P3_ADD_552_U47 = ~P3_EBX_REG_29_;
  assign new_P3_ADD_552_U48 = ~new_P3_ADD_552_U94 | ~new_P3_ADD_552_U122;
  assign new_P3_ADD_552_U49 = ~new_P3_ADD_552_U123 | ~P3_EBX_REG_29_;
  assign new_P3_ADD_552_U50 = ~P3_EBX_REG_30_;
  assign new_P3_ADD_552_U51 = ~new_P3_ADD_552_U142 | ~new_P3_ADD_552_U141;
  assign new_P3_ADD_552_U52 = ~new_P3_ADD_552_U144 | ~new_P3_ADD_552_U143;
  assign new_P3_ADD_552_U53 = ~new_P3_ADD_552_U146 | ~new_P3_ADD_552_U145;
  assign new_P3_ADD_552_U54 = ~new_P3_ADD_552_U148 | ~new_P3_ADD_552_U147;
  assign new_P3_ADD_552_U55 = ~new_P3_ADD_552_U150 | ~new_P3_ADD_552_U149;
  assign new_P3_ADD_552_U56 = ~new_P3_ADD_552_U152 | ~new_P3_ADD_552_U151;
  assign new_P3_ADD_552_U57 = ~new_P3_ADD_552_U154 | ~new_P3_ADD_552_U153;
  assign new_P3_ADD_552_U58 = ~new_P3_ADD_552_U156 | ~new_P3_ADD_552_U155;
  assign new_P3_ADD_552_U59 = ~new_P3_ADD_552_U158 | ~new_P3_ADD_552_U157;
  assign new_P3_ADD_552_U60 = ~new_P3_ADD_552_U160 | ~new_P3_ADD_552_U159;
  assign new_P3_ADD_552_U61 = ~new_P3_ADD_552_U162 | ~new_P3_ADD_552_U161;
  assign new_P3_ADD_552_U62 = ~new_P3_ADD_552_U164 | ~new_P3_ADD_552_U163;
  assign new_P3_ADD_552_U63 = ~new_P3_ADD_552_U166 | ~new_P3_ADD_552_U165;
  assign new_P3_ADD_552_U64 = ~new_P3_ADD_552_U168 | ~new_P3_ADD_552_U167;
  assign new_P3_ADD_552_U65 = ~new_P3_ADD_552_U170 | ~new_P3_ADD_552_U169;
  assign new_P3_ADD_552_U66 = ~new_P3_ADD_552_U172 | ~new_P3_ADD_552_U171;
  assign new_P3_ADD_552_U67 = ~new_P3_ADD_552_U174 | ~new_P3_ADD_552_U173;
  assign new_P3_ADD_552_U68 = ~new_P3_ADD_552_U176 | ~new_P3_ADD_552_U175;
  assign new_P3_ADD_552_U69 = ~new_P3_ADD_552_U178 | ~new_P3_ADD_552_U177;
  assign new_P3_ADD_552_U70 = ~new_P3_ADD_552_U180 | ~new_P3_ADD_552_U179;
  assign new_P3_ADD_552_U71 = ~new_P3_ADD_552_U182 | ~new_P3_ADD_552_U181;
  assign new_P3_ADD_552_U72 = ~new_P3_ADD_552_U184 | ~new_P3_ADD_552_U183;
  assign new_P3_ADD_552_U73 = ~new_P3_ADD_552_U186 | ~new_P3_ADD_552_U185;
  assign new_P3_ADD_552_U74 = ~new_P3_ADD_552_U188 | ~new_P3_ADD_552_U187;
  assign new_P3_ADD_552_U75 = ~new_P3_ADD_552_U190 | ~new_P3_ADD_552_U189;
  assign new_P3_ADD_552_U76 = ~new_P3_ADD_552_U192 | ~new_P3_ADD_552_U191;
  assign new_P3_ADD_552_U77 = ~new_P3_ADD_552_U194 | ~new_P3_ADD_552_U193;
  assign new_P3_ADD_552_U78 = ~new_P3_ADD_552_U196 | ~new_P3_ADD_552_U195;
  assign new_P3_ADD_552_U79 = ~new_P3_ADD_552_U198 | ~new_P3_ADD_552_U197;
  assign new_P3_ADD_552_U80 = ~new_P3_ADD_552_U200 | ~new_P3_ADD_552_U199;
  assign new_P3_ADD_552_U81 = ~new_P3_ADD_552_U202 | ~new_P3_ADD_552_U201;
  assign new_P3_ADD_552_U82 = P3_EBX_REG_3_ & P3_EBX_REG_4_;
  assign new_P3_ADD_552_U83 = P3_EBX_REG_5_ & P3_EBX_REG_6_;
  assign new_P3_ADD_552_U84 = P3_EBX_REG_7_ & P3_EBX_REG_8_;
  assign new_P3_ADD_552_U85 = P3_EBX_REG_9_ & P3_EBX_REG_10_;
  assign new_P3_ADD_552_U86 = P3_EBX_REG_11_ & P3_EBX_REG_12_;
  assign new_P3_ADD_552_U87 = P3_EBX_REG_13_ & P3_EBX_REG_14_;
  assign new_P3_ADD_552_U88 = P3_EBX_REG_16_ & P3_EBX_REG_15_;
  assign new_P3_ADD_552_U89 = P3_EBX_REG_17_ & P3_EBX_REG_18_;
  assign new_P3_ADD_552_U90 = P3_EBX_REG_19_ & P3_EBX_REG_20_;
  assign new_P3_ADD_552_U91 = P3_EBX_REG_22_ & P3_EBX_REG_21_;
  assign new_P3_ADD_552_U92 = P3_EBX_REG_23_ & P3_EBX_REG_24_;
  assign new_P3_ADD_552_U93 = P3_EBX_REG_25_ & P3_EBX_REG_26_;
  assign new_P3_ADD_552_U94 = P3_EBX_REG_28_ & P3_EBX_REG_27_;
  assign new_P3_ADD_552_U95 = ~new_P3_ADD_552_U118 | ~P3_EBX_REG_7_;
  assign new_P3_ADD_552_U96 = ~new_P3_ADD_552_U112 | ~P3_EBX_REG_5_;
  assign new_P3_ADD_552_U97 = ~new_P3_ADD_552_U111 | ~P3_EBX_REG_3_;
  assign new_P3_ADD_552_U98 = ~P3_EBX_REG_31_;
  assign new_P3_ADD_552_U99 = ~P3_EBX_REG_30_ | ~new_P3_ADD_552_U128;
  assign new_P3_ADD_552_U100 = ~P3_EBX_REG_1_ | ~P3_EBX_REG_0_;
  assign new_P3_ADD_552_U101 = ~new_P3_ADD_552_U122 | ~P3_EBX_REG_27_;
  assign new_P3_ADD_552_U102 = ~new_P3_ADD_552_U116 | ~P3_EBX_REG_25_;
  assign new_P3_ADD_552_U103 = ~new_P3_ADD_552_U115 | ~P3_EBX_REG_23_;
  assign new_P3_ADD_552_U104 = ~new_P3_ADD_552_U121 | ~P3_EBX_REG_21_;
  assign new_P3_ADD_552_U105 = ~new_P3_ADD_552_U114 | ~P3_EBX_REG_19_;
  assign new_P3_ADD_552_U106 = ~new_P3_ADD_552_U117 | ~P3_EBX_REG_17_;
  assign new_P3_ADD_552_U107 = ~new_P3_ADD_552_U124 | ~P3_EBX_REG_15_;
  assign new_P3_ADD_552_U108 = ~new_P3_ADD_552_U119 | ~P3_EBX_REG_13_;
  assign new_P3_ADD_552_U109 = ~new_P3_ADD_552_U113 | ~P3_EBX_REG_11_;
  assign new_P3_ADD_552_U110 = ~P3_EBX_REG_9_ | ~new_P3_ADD_552_U120;
  assign new_P3_ADD_552_U111 = ~new_P3_ADD_552_U10;
  assign new_P3_ADD_552_U112 = ~new_P3_ADD_552_U13;
  assign new_P3_ADD_552_U113 = ~new_P3_ADD_552_U22;
  assign new_P3_ADD_552_U114 = ~new_P3_ADD_552_U34;
  assign new_P3_ADD_552_U115 = ~new_P3_ADD_552_U40;
  assign new_P3_ADD_552_U116 = ~new_P3_ADD_552_U43;
  assign new_P3_ADD_552_U117 = ~new_P3_ADD_552_U31;
  assign new_P3_ADD_552_U118 = ~new_P3_ADD_552_U16;
  assign new_P3_ADD_552_U119 = ~new_P3_ADD_552_U25;
  assign new_P3_ADD_552_U120 = ~new_P3_ADD_552_U17;
  assign new_P3_ADD_552_U121 = ~new_P3_ADD_552_U36;
  assign new_P3_ADD_552_U122 = ~new_P3_ADD_552_U46;
  assign new_P3_ADD_552_U123 = ~new_P3_ADD_552_U48;
  assign new_P3_ADD_552_U124 = ~new_P3_ADD_552_U27;
  assign new_P3_ADD_552_U125 = ~new_P3_ADD_552_U95;
  assign new_P3_ADD_552_U126 = ~new_P3_ADD_552_U96;
  assign new_P3_ADD_552_U127 = ~new_P3_ADD_552_U97;
  assign new_P3_ADD_552_U128 = ~new_P3_ADD_552_U49;
  assign new_P3_ADD_552_U129 = ~new_P3_ADD_552_U99;
  assign new_P3_ADD_552_U130 = ~new_P3_ADD_552_U100;
  assign new_P3_ADD_552_U131 = ~new_P3_ADD_552_U101;
  assign new_P3_ADD_552_U132 = ~new_P3_ADD_552_U102;
  assign new_P3_ADD_552_U133 = ~new_P3_ADD_552_U103;
  assign new_P3_ADD_552_U134 = ~new_P3_ADD_552_U104;
  assign new_P3_ADD_552_U135 = ~new_P3_ADD_552_U105;
  assign new_P3_ADD_552_U136 = ~new_P3_ADD_552_U106;
  assign new_P3_ADD_552_U137 = ~new_P3_ADD_552_U107;
  assign new_P3_ADD_552_U138 = ~new_P3_ADD_552_U108;
  assign new_P3_ADD_552_U139 = ~new_P3_ADD_552_U109;
  assign new_P3_ADD_552_U140 = ~new_P3_ADD_552_U110;
  assign new_P3_ADD_552_U141 = ~new_P3_ADD_552_U120 | ~new_P3_ADD_552_U18;
  assign new_P3_ADD_552_U142 = ~P3_EBX_REG_9_ | ~new_P3_ADD_552_U17;
  assign new_P3_ADD_552_U143 = ~P3_EBX_REG_8_ | ~new_P3_ADD_552_U95;
  assign new_P3_ADD_552_U144 = ~new_P3_ADD_552_U125 | ~new_P3_ADD_552_U14;
  assign new_P3_ADD_552_U145 = ~new_P3_ADD_552_U118 | ~new_P3_ADD_552_U15;
  assign new_P3_ADD_552_U146 = ~P3_EBX_REG_7_ | ~new_P3_ADD_552_U16;
  assign new_P3_ADD_552_U147 = ~P3_EBX_REG_6_ | ~new_P3_ADD_552_U96;
  assign new_P3_ADD_552_U148 = ~new_P3_ADD_552_U126 | ~new_P3_ADD_552_U11;
  assign new_P3_ADD_552_U149 = ~new_P3_ADD_552_U112 | ~new_P3_ADD_552_U12;
  assign new_P3_ADD_552_U150 = ~P3_EBX_REG_5_ | ~new_P3_ADD_552_U13;
  assign new_P3_ADD_552_U151 = ~P3_EBX_REG_4_ | ~new_P3_ADD_552_U97;
  assign new_P3_ADD_552_U152 = ~new_P3_ADD_552_U127 | ~new_P3_ADD_552_U8;
  assign new_P3_ADD_552_U153 = ~new_P3_ADD_552_U111 | ~new_P3_ADD_552_U9;
  assign new_P3_ADD_552_U154 = ~P3_EBX_REG_3_ | ~new_P3_ADD_552_U10;
  assign new_P3_ADD_552_U155 = ~P3_EBX_REG_31_ | ~new_P3_ADD_552_U99;
  assign new_P3_ADD_552_U156 = ~new_P3_ADD_552_U129 | ~new_P3_ADD_552_U98;
  assign new_P3_ADD_552_U157 = ~P3_EBX_REG_30_ | ~new_P3_ADD_552_U49;
  assign new_P3_ADD_552_U158 = ~new_P3_ADD_552_U128 | ~new_P3_ADD_552_U50;
  assign new_P3_ADD_552_U159 = ~P3_EBX_REG_2_ | ~new_P3_ADD_552_U100;
  assign new_P3_ADD_552_U160 = ~new_P3_ADD_552_U130 | ~new_P3_ADD_552_U6;
  assign new_P3_ADD_552_U161 = ~new_P3_ADD_552_U123 | ~new_P3_ADD_552_U47;
  assign new_P3_ADD_552_U162 = ~P3_EBX_REG_29_ | ~new_P3_ADD_552_U48;
  assign new_P3_ADD_552_U163 = ~P3_EBX_REG_28_ | ~new_P3_ADD_552_U101;
  assign new_P3_ADD_552_U164 = ~new_P3_ADD_552_U131 | ~new_P3_ADD_552_U45;
  assign new_P3_ADD_552_U165 = ~new_P3_ADD_552_U122 | ~new_P3_ADD_552_U44;
  assign new_P3_ADD_552_U166 = ~P3_EBX_REG_27_ | ~new_P3_ADD_552_U46;
  assign new_P3_ADD_552_U167 = ~P3_EBX_REG_26_ | ~new_P3_ADD_552_U102;
  assign new_P3_ADD_552_U168 = ~new_P3_ADD_552_U132 | ~new_P3_ADD_552_U41;
  assign new_P3_ADD_552_U169 = ~new_P3_ADD_552_U116 | ~new_P3_ADD_552_U42;
  assign new_P3_ADD_552_U170 = ~P3_EBX_REG_25_ | ~new_P3_ADD_552_U43;
  assign new_P3_ADD_552_U171 = ~P3_EBX_REG_24_ | ~new_P3_ADD_552_U103;
  assign new_P3_ADD_552_U172 = ~new_P3_ADD_552_U133 | ~new_P3_ADD_552_U38;
  assign new_P3_ADD_552_U173 = ~new_P3_ADD_552_U115 | ~new_P3_ADD_552_U39;
  assign new_P3_ADD_552_U174 = ~P3_EBX_REG_23_ | ~new_P3_ADD_552_U40;
  assign new_P3_ADD_552_U175 = ~P3_EBX_REG_22_ | ~new_P3_ADD_552_U104;
  assign new_P3_ADD_552_U176 = ~new_P3_ADD_552_U134 | ~new_P3_ADD_552_U37;
  assign new_P3_ADD_552_U177 = ~new_P3_ADD_552_U121 | ~new_P3_ADD_552_U35;
  assign new_P3_ADD_552_U178 = ~P3_EBX_REG_21_ | ~new_P3_ADD_552_U36;
  assign new_P3_ADD_552_U179 = ~P3_EBX_REG_20_ | ~new_P3_ADD_552_U105;
  assign new_P3_ADD_552_U180 = ~new_P3_ADD_552_U135 | ~new_P3_ADD_552_U32;
  assign new_P3_ADD_552_U181 = ~P3_EBX_REG_0_ | ~new_P3_ADD_552_U7;
  assign new_P3_ADD_552_U182 = ~P3_EBX_REG_1_ | ~new_P3_ADD_552_U5;
  assign new_P3_ADD_552_U183 = ~new_P3_ADD_552_U114 | ~new_P3_ADD_552_U33;
  assign new_P3_ADD_552_U184 = ~P3_EBX_REG_19_ | ~new_P3_ADD_552_U34;
  assign new_P3_ADD_552_U185 = ~P3_EBX_REG_18_ | ~new_P3_ADD_552_U106;
  assign new_P3_ADD_552_U186 = ~new_P3_ADD_552_U136 | ~new_P3_ADD_552_U29;
  assign new_P3_ADD_552_U187 = ~new_P3_ADD_552_U117 | ~new_P3_ADD_552_U30;
  assign new_P3_ADD_552_U188 = ~P3_EBX_REG_17_ | ~new_P3_ADD_552_U31;
  assign new_P3_ADD_552_U189 = ~P3_EBX_REG_16_ | ~new_P3_ADD_552_U107;
  assign new_P3_ADD_552_U190 = ~new_P3_ADD_552_U137 | ~new_P3_ADD_552_U28;
  assign new_P3_ADD_552_U191 = ~new_P3_ADD_552_U124 | ~new_P3_ADD_552_U26;
  assign new_P3_ADD_552_U192 = ~P3_EBX_REG_15_ | ~new_P3_ADD_552_U27;
  assign new_P3_ADD_552_U193 = ~P3_EBX_REG_14_ | ~new_P3_ADD_552_U108;
  assign new_P3_ADD_552_U194 = ~new_P3_ADD_552_U138 | ~new_P3_ADD_552_U23;
  assign new_P3_ADD_552_U195 = ~new_P3_ADD_552_U119 | ~new_P3_ADD_552_U24;
  assign new_P3_ADD_552_U196 = ~P3_EBX_REG_13_ | ~new_P3_ADD_552_U25;
  assign new_P3_ADD_552_U197 = ~P3_EBX_REG_12_ | ~new_P3_ADD_552_U109;
  assign new_P3_ADD_552_U198 = ~new_P3_ADD_552_U139 | ~new_P3_ADD_552_U20;
  assign new_P3_ADD_552_U199 = ~new_P3_ADD_552_U113 | ~new_P3_ADD_552_U21;
  assign new_P3_ADD_552_U200 = ~P3_EBX_REG_11_ | ~new_P3_ADD_552_U22;
  assign new_P3_ADD_552_U201 = ~P3_EBX_REG_10_ | ~new_P3_ADD_552_U110;
  assign new_P3_ADD_552_U202 = ~new_P3_ADD_552_U140 | ~new_P3_ADD_552_U19;
  assign new_P3_ADD_546_U5 = ~P3_EAX_REG_0_;
  assign new_P3_ADD_546_U6 = ~P3_EAX_REG_2_;
  assign new_P3_ADD_546_U7 = ~P3_EAX_REG_1_;
  assign new_P3_ADD_546_U8 = ~P3_EAX_REG_4_;
  assign new_P3_ADD_546_U9 = ~P3_EAX_REG_3_;
  assign new_P3_ADD_546_U10 = ~P3_EAX_REG_1_ | ~P3_EAX_REG_2_ | ~P3_EAX_REG_0_;
  assign new_P3_ADD_546_U11 = ~P3_EAX_REG_6_;
  assign new_P3_ADD_546_U12 = ~P3_EAX_REG_5_;
  assign new_P3_ADD_546_U13 = ~new_P3_ADD_546_U82 | ~new_P3_ADD_546_U111;
  assign new_P3_ADD_546_U14 = ~P3_EAX_REG_8_;
  assign new_P3_ADD_546_U15 = ~P3_EAX_REG_7_;
  assign new_P3_ADD_546_U16 = ~new_P3_ADD_546_U83 | ~new_P3_ADD_546_U112;
  assign new_P3_ADD_546_U17 = ~new_P3_ADD_546_U84 | ~new_P3_ADD_546_U118;
  assign new_P3_ADD_546_U18 = ~P3_EAX_REG_9_;
  assign new_P3_ADD_546_U19 = ~P3_EAX_REG_10_;
  assign new_P3_ADD_546_U20 = ~P3_EAX_REG_12_;
  assign new_P3_ADD_546_U21 = ~P3_EAX_REG_11_;
  assign new_P3_ADD_546_U22 = ~new_P3_ADD_546_U85 | ~new_P3_ADD_546_U120;
  assign new_P3_ADD_546_U23 = ~P3_EAX_REG_14_;
  assign new_P3_ADD_546_U24 = ~P3_EAX_REG_13_;
  assign new_P3_ADD_546_U25 = ~new_P3_ADD_546_U86 | ~new_P3_ADD_546_U113;
  assign new_P3_ADD_546_U26 = ~P3_EAX_REG_15_;
  assign new_P3_ADD_546_U27 = ~new_P3_ADD_546_U87 | ~new_P3_ADD_546_U119;
  assign new_P3_ADD_546_U28 = ~P3_EAX_REG_16_;
  assign new_P3_ADD_546_U29 = ~P3_EAX_REG_18_;
  assign new_P3_ADD_546_U30 = ~P3_EAX_REG_17_;
  assign new_P3_ADD_546_U31 = ~new_P3_ADD_546_U88 | ~new_P3_ADD_546_U124;
  assign new_P3_ADD_546_U32 = ~P3_EAX_REG_20_;
  assign new_P3_ADD_546_U33 = ~P3_EAX_REG_19_;
  assign new_P3_ADD_546_U34 = ~new_P3_ADD_546_U89 | ~new_P3_ADD_546_U117;
  assign new_P3_ADD_546_U35 = ~P3_EAX_REG_21_;
  assign new_P3_ADD_546_U36 = ~new_P3_ADD_546_U90 | ~new_P3_ADD_546_U114;
  assign new_P3_ADD_546_U37 = ~P3_EAX_REG_22_;
  assign new_P3_ADD_546_U38 = ~P3_EAX_REG_24_;
  assign new_P3_ADD_546_U39 = ~P3_EAX_REG_23_;
  assign new_P3_ADD_546_U40 = ~new_P3_ADD_546_U91 | ~new_P3_ADD_546_U121;
  assign new_P3_ADD_546_U41 = ~P3_EAX_REG_26_;
  assign new_P3_ADD_546_U42 = ~P3_EAX_REG_25_;
  assign new_P3_ADD_546_U43 = ~new_P3_ADD_546_U92 | ~new_P3_ADD_546_U115;
  assign new_P3_ADD_546_U44 = ~P3_EAX_REG_27_;
  assign new_P3_ADD_546_U45 = ~P3_EAX_REG_28_;
  assign new_P3_ADD_546_U46 = ~new_P3_ADD_546_U93 | ~new_P3_ADD_546_U116;
  assign new_P3_ADD_546_U47 = ~P3_EAX_REG_29_;
  assign new_P3_ADD_546_U48 = ~new_P3_ADD_546_U94 | ~new_P3_ADD_546_U122;
  assign new_P3_ADD_546_U49 = ~new_P3_ADD_546_U123 | ~P3_EAX_REG_29_;
  assign new_P3_ADD_546_U50 = ~P3_EAX_REG_30_;
  assign new_P3_ADD_546_U51 = ~new_P3_ADD_546_U142 | ~new_P3_ADD_546_U141;
  assign new_P3_ADD_546_U52 = ~new_P3_ADD_546_U144 | ~new_P3_ADD_546_U143;
  assign new_P3_ADD_546_U53 = ~new_P3_ADD_546_U146 | ~new_P3_ADD_546_U145;
  assign new_P3_ADD_546_U54 = ~new_P3_ADD_546_U148 | ~new_P3_ADD_546_U147;
  assign new_P3_ADD_546_U55 = ~new_P3_ADD_546_U150 | ~new_P3_ADD_546_U149;
  assign new_P3_ADD_546_U56 = ~new_P3_ADD_546_U152 | ~new_P3_ADD_546_U151;
  assign new_P3_ADD_546_U57 = ~new_P3_ADD_546_U154 | ~new_P3_ADD_546_U153;
  assign new_P3_ADD_546_U58 = ~new_P3_ADD_546_U156 | ~new_P3_ADD_546_U155;
  assign new_P3_ADD_546_U59 = ~new_P3_ADD_546_U158 | ~new_P3_ADD_546_U157;
  assign new_P3_ADD_546_U60 = ~new_P3_ADD_546_U160 | ~new_P3_ADD_546_U159;
  assign new_P3_ADD_546_U61 = ~new_P3_ADD_546_U162 | ~new_P3_ADD_546_U161;
  assign new_P3_ADD_546_U62 = ~new_P3_ADD_546_U164 | ~new_P3_ADD_546_U163;
  assign new_P3_ADD_546_U63 = ~new_P3_ADD_546_U166 | ~new_P3_ADD_546_U165;
  assign new_P3_ADD_546_U64 = ~new_P3_ADD_546_U168 | ~new_P3_ADD_546_U167;
  assign new_P3_ADD_546_U65 = ~new_P3_ADD_546_U170 | ~new_P3_ADD_546_U169;
  assign new_P3_ADD_546_U66 = ~new_P3_ADD_546_U172 | ~new_P3_ADD_546_U171;
  assign new_P3_ADD_546_U67 = ~new_P3_ADD_546_U174 | ~new_P3_ADD_546_U173;
  assign new_P3_ADD_546_U68 = ~new_P3_ADD_546_U176 | ~new_P3_ADD_546_U175;
  assign new_P3_ADD_546_U69 = ~new_P3_ADD_546_U178 | ~new_P3_ADD_546_U177;
  assign new_P3_ADD_546_U70 = ~new_P3_ADD_546_U180 | ~new_P3_ADD_546_U179;
  assign new_P3_ADD_546_U71 = ~new_P3_ADD_546_U182 | ~new_P3_ADD_546_U181;
  assign new_P3_ADD_546_U72 = ~new_P3_ADD_546_U184 | ~new_P3_ADD_546_U183;
  assign new_P3_ADD_546_U73 = ~new_P3_ADD_546_U186 | ~new_P3_ADD_546_U185;
  assign new_P3_ADD_546_U74 = ~new_P3_ADD_546_U188 | ~new_P3_ADD_546_U187;
  assign new_P3_ADD_546_U75 = ~new_P3_ADD_546_U190 | ~new_P3_ADD_546_U189;
  assign new_P3_ADD_546_U76 = ~new_P3_ADD_546_U192 | ~new_P3_ADD_546_U191;
  assign new_P3_ADD_546_U77 = ~new_P3_ADD_546_U194 | ~new_P3_ADD_546_U193;
  assign new_P3_ADD_546_U78 = ~new_P3_ADD_546_U196 | ~new_P3_ADD_546_U195;
  assign new_P3_ADD_546_U79 = ~new_P3_ADD_546_U198 | ~new_P3_ADD_546_U197;
  assign new_P3_ADD_546_U80 = ~new_P3_ADD_546_U200 | ~new_P3_ADD_546_U199;
  assign new_P3_ADD_546_U81 = ~new_P3_ADD_546_U202 | ~new_P3_ADD_546_U201;
  assign new_P3_ADD_546_U82 = P3_EAX_REG_3_ & P3_EAX_REG_4_;
  assign new_P3_ADD_546_U83 = P3_EAX_REG_5_ & P3_EAX_REG_6_;
  assign new_P3_ADD_546_U84 = P3_EAX_REG_7_ & P3_EAX_REG_8_;
  assign new_P3_ADD_546_U85 = P3_EAX_REG_9_ & P3_EAX_REG_10_;
  assign new_P3_ADD_546_U86 = P3_EAX_REG_11_ & P3_EAX_REG_12_;
  assign new_P3_ADD_546_U87 = P3_EAX_REG_13_ & P3_EAX_REG_14_;
  assign new_P3_ADD_546_U88 = P3_EAX_REG_16_ & P3_EAX_REG_15_;
  assign new_P3_ADD_546_U89 = P3_EAX_REG_17_ & P3_EAX_REG_18_;
  assign new_P3_ADD_546_U90 = P3_EAX_REG_19_ & P3_EAX_REG_20_;
  assign new_P3_ADD_546_U91 = P3_EAX_REG_22_ & P3_EAX_REG_21_;
  assign new_P3_ADD_546_U92 = P3_EAX_REG_23_ & P3_EAX_REG_24_;
  assign new_P3_ADD_546_U93 = P3_EAX_REG_25_ & P3_EAX_REG_26_;
  assign new_P3_ADD_546_U94 = P3_EAX_REG_28_ & P3_EAX_REG_27_;
  assign new_P3_ADD_546_U95 = ~new_P3_ADD_546_U118 | ~P3_EAX_REG_7_;
  assign new_P3_ADD_546_U96 = ~new_P3_ADD_546_U112 | ~P3_EAX_REG_5_;
  assign new_P3_ADD_546_U97 = ~new_P3_ADD_546_U111 | ~P3_EAX_REG_3_;
  assign new_P3_ADD_546_U98 = ~P3_EAX_REG_31_;
  assign new_P3_ADD_546_U99 = ~P3_EAX_REG_30_ | ~new_P3_ADD_546_U128;
  assign new_P3_ADD_546_U100 = ~P3_EAX_REG_1_ | ~P3_EAX_REG_0_;
  assign new_P3_ADD_546_U101 = ~new_P3_ADD_546_U122 | ~P3_EAX_REG_27_;
  assign new_P3_ADD_546_U102 = ~new_P3_ADD_546_U116 | ~P3_EAX_REG_25_;
  assign new_P3_ADD_546_U103 = ~new_P3_ADD_546_U115 | ~P3_EAX_REG_23_;
  assign new_P3_ADD_546_U104 = ~new_P3_ADD_546_U121 | ~P3_EAX_REG_21_;
  assign new_P3_ADD_546_U105 = ~new_P3_ADD_546_U114 | ~P3_EAX_REG_19_;
  assign new_P3_ADD_546_U106 = ~new_P3_ADD_546_U117 | ~P3_EAX_REG_17_;
  assign new_P3_ADD_546_U107 = ~new_P3_ADD_546_U124 | ~P3_EAX_REG_15_;
  assign new_P3_ADD_546_U108 = ~new_P3_ADD_546_U119 | ~P3_EAX_REG_13_;
  assign new_P3_ADD_546_U109 = ~new_P3_ADD_546_U113 | ~P3_EAX_REG_11_;
  assign new_P3_ADD_546_U110 = ~P3_EAX_REG_9_ | ~new_P3_ADD_546_U120;
  assign new_P3_ADD_546_U111 = ~new_P3_ADD_546_U10;
  assign new_P3_ADD_546_U112 = ~new_P3_ADD_546_U13;
  assign new_P3_ADD_546_U113 = ~new_P3_ADD_546_U22;
  assign new_P3_ADD_546_U114 = ~new_P3_ADD_546_U34;
  assign new_P3_ADD_546_U115 = ~new_P3_ADD_546_U40;
  assign new_P3_ADD_546_U116 = ~new_P3_ADD_546_U43;
  assign new_P3_ADD_546_U117 = ~new_P3_ADD_546_U31;
  assign new_P3_ADD_546_U118 = ~new_P3_ADD_546_U16;
  assign new_P3_ADD_546_U119 = ~new_P3_ADD_546_U25;
  assign new_P3_ADD_546_U120 = ~new_P3_ADD_546_U17;
  assign new_P3_ADD_546_U121 = ~new_P3_ADD_546_U36;
  assign new_P3_ADD_546_U122 = ~new_P3_ADD_546_U46;
  assign new_P3_ADD_546_U123 = ~new_P3_ADD_546_U48;
  assign new_P3_ADD_546_U124 = ~new_P3_ADD_546_U27;
  assign new_P3_ADD_546_U125 = ~new_P3_ADD_546_U95;
  assign new_P3_ADD_546_U126 = ~new_P3_ADD_546_U96;
  assign new_P3_ADD_546_U127 = ~new_P3_ADD_546_U97;
  assign new_P3_ADD_546_U128 = ~new_P3_ADD_546_U49;
  assign new_P3_ADD_546_U129 = ~new_P3_ADD_546_U99;
  assign new_P3_ADD_546_U130 = ~new_P3_ADD_546_U100;
  assign new_P3_ADD_546_U131 = ~new_P3_ADD_546_U101;
  assign new_P3_ADD_546_U132 = ~new_P3_ADD_546_U102;
  assign new_P3_ADD_546_U133 = ~new_P3_ADD_546_U103;
  assign new_P3_ADD_546_U134 = ~new_P3_ADD_546_U104;
  assign new_P3_ADD_546_U135 = ~new_P3_ADD_546_U105;
  assign new_P3_ADD_546_U136 = ~new_P3_ADD_546_U106;
  assign new_P3_ADD_546_U137 = ~new_P3_ADD_546_U107;
  assign new_P3_ADD_546_U138 = ~new_P3_ADD_546_U108;
  assign new_P3_ADD_546_U139 = ~new_P3_ADD_546_U109;
  assign new_P3_ADD_546_U140 = ~new_P3_ADD_546_U110;
  assign new_P3_ADD_546_U141 = ~new_P3_ADD_546_U120 | ~new_P3_ADD_546_U18;
  assign new_P3_ADD_546_U142 = ~P3_EAX_REG_9_ | ~new_P3_ADD_546_U17;
  assign new_P3_ADD_546_U143 = ~P3_EAX_REG_8_ | ~new_P3_ADD_546_U95;
  assign new_P3_ADD_546_U144 = ~new_P3_ADD_546_U125 | ~new_P3_ADD_546_U14;
  assign new_P3_ADD_546_U145 = ~new_P3_ADD_546_U118 | ~new_P3_ADD_546_U15;
  assign new_P3_ADD_546_U146 = ~P3_EAX_REG_7_ | ~new_P3_ADD_546_U16;
  assign new_P3_ADD_546_U147 = ~P3_EAX_REG_6_ | ~new_P3_ADD_546_U96;
  assign new_P3_ADD_546_U148 = ~new_P3_ADD_546_U126 | ~new_P3_ADD_546_U11;
  assign new_P3_ADD_546_U149 = ~new_P3_ADD_546_U112 | ~new_P3_ADD_546_U12;
  assign new_P3_ADD_546_U150 = ~P3_EAX_REG_5_ | ~new_P3_ADD_546_U13;
  assign new_P3_ADD_546_U151 = ~P3_EAX_REG_4_ | ~new_P3_ADD_546_U97;
  assign new_P3_ADD_546_U152 = ~new_P3_ADD_546_U127 | ~new_P3_ADD_546_U8;
  assign new_P3_ADD_546_U153 = ~new_P3_ADD_546_U111 | ~new_P3_ADD_546_U9;
  assign new_P3_ADD_546_U154 = ~P3_EAX_REG_3_ | ~new_P3_ADD_546_U10;
  assign new_P3_ADD_546_U155 = ~P3_EAX_REG_31_ | ~new_P3_ADD_546_U99;
  assign new_P3_ADD_546_U156 = ~new_P3_ADD_546_U129 | ~new_P3_ADD_546_U98;
  assign new_P3_ADD_546_U157 = ~P3_EAX_REG_30_ | ~new_P3_ADD_546_U49;
  assign new_P3_ADD_546_U158 = ~new_P3_ADD_546_U128 | ~new_P3_ADD_546_U50;
  assign new_P3_ADD_546_U159 = ~P3_EAX_REG_2_ | ~new_P3_ADD_546_U100;
  assign new_P3_ADD_546_U160 = ~new_P3_ADD_546_U130 | ~new_P3_ADD_546_U6;
  assign new_P3_ADD_546_U161 = ~new_P3_ADD_546_U123 | ~new_P3_ADD_546_U47;
  assign new_P3_ADD_546_U162 = ~P3_EAX_REG_29_ | ~new_P3_ADD_546_U48;
  assign new_P3_ADD_546_U163 = ~P3_EAX_REG_28_ | ~new_P3_ADD_546_U101;
  assign new_P3_ADD_546_U164 = ~new_P3_ADD_546_U131 | ~new_P3_ADD_546_U45;
  assign new_P3_ADD_546_U165 = ~new_P3_ADD_546_U122 | ~new_P3_ADD_546_U44;
  assign new_P3_ADD_546_U166 = ~P3_EAX_REG_27_ | ~new_P3_ADD_546_U46;
  assign new_P3_ADD_546_U167 = ~P3_EAX_REG_26_ | ~new_P3_ADD_546_U102;
  assign new_P3_ADD_546_U168 = ~new_P3_ADD_546_U132 | ~new_P3_ADD_546_U41;
  assign new_P3_ADD_546_U169 = ~new_P3_ADD_546_U116 | ~new_P3_ADD_546_U42;
  assign new_P3_ADD_546_U170 = ~P3_EAX_REG_25_ | ~new_P3_ADD_546_U43;
  assign new_P3_ADD_546_U171 = ~P3_EAX_REG_24_ | ~new_P3_ADD_546_U103;
  assign new_P3_ADD_546_U172 = ~new_P3_ADD_546_U133 | ~new_P3_ADD_546_U38;
  assign new_P3_ADD_546_U173 = ~new_P3_ADD_546_U115 | ~new_P3_ADD_546_U39;
  assign new_P3_ADD_546_U174 = ~P3_EAX_REG_23_ | ~new_P3_ADD_546_U40;
  assign new_P3_ADD_546_U175 = ~P3_EAX_REG_22_ | ~new_P3_ADD_546_U104;
  assign new_P3_ADD_546_U176 = ~new_P3_ADD_546_U134 | ~new_P3_ADD_546_U37;
  assign new_P3_ADD_546_U177 = ~new_P3_ADD_546_U121 | ~new_P3_ADD_546_U35;
  assign new_P3_ADD_546_U178 = ~P3_EAX_REG_21_ | ~new_P3_ADD_546_U36;
  assign new_P3_ADD_546_U179 = ~P3_EAX_REG_20_ | ~new_P3_ADD_546_U105;
  assign new_P3_ADD_546_U180 = ~new_P3_ADD_546_U135 | ~new_P3_ADD_546_U32;
  assign new_P3_ADD_546_U181 = ~P3_EAX_REG_0_ | ~new_P3_ADD_546_U7;
  assign new_P3_ADD_546_U182 = ~P3_EAX_REG_1_ | ~new_P3_ADD_546_U5;
  assign new_P3_ADD_546_U183 = ~new_P3_ADD_546_U114 | ~new_P3_ADD_546_U33;
  assign new_P3_ADD_546_U184 = ~P3_EAX_REG_19_ | ~new_P3_ADD_546_U34;
  assign new_P3_ADD_546_U185 = ~P3_EAX_REG_18_ | ~new_P3_ADD_546_U106;
  assign new_P3_ADD_546_U186 = ~new_P3_ADD_546_U136 | ~new_P3_ADD_546_U29;
  assign new_P3_ADD_546_U187 = ~new_P3_ADD_546_U117 | ~new_P3_ADD_546_U30;
  assign new_P3_ADD_546_U188 = ~P3_EAX_REG_17_ | ~new_P3_ADD_546_U31;
  assign new_P3_ADD_546_U189 = ~P3_EAX_REG_16_ | ~new_P3_ADD_546_U107;
  assign new_P3_ADD_546_U190 = ~new_P3_ADD_546_U137 | ~new_P3_ADD_546_U28;
  assign new_P3_ADD_546_U191 = ~new_P3_ADD_546_U124 | ~new_P3_ADD_546_U26;
  assign new_P3_ADD_546_U192 = ~P3_EAX_REG_15_ | ~new_P3_ADD_546_U27;
  assign new_P3_ADD_546_U193 = ~P3_EAX_REG_14_ | ~new_P3_ADD_546_U108;
  assign new_P3_ADD_546_U194 = ~new_P3_ADD_546_U138 | ~new_P3_ADD_546_U23;
  assign new_P3_ADD_546_U195 = ~new_P3_ADD_546_U119 | ~new_P3_ADD_546_U24;
  assign new_P3_ADD_546_U196 = ~P3_EAX_REG_13_ | ~new_P3_ADD_546_U25;
  assign new_P3_ADD_546_U197 = ~P3_EAX_REG_12_ | ~new_P3_ADD_546_U109;
  assign new_P3_ADD_546_U198 = ~new_P3_ADD_546_U139 | ~new_P3_ADD_546_U20;
  assign new_P3_ADD_546_U199 = ~new_P3_ADD_546_U113 | ~new_P3_ADD_546_U21;
  assign new_P3_ADD_546_U200 = ~P3_EAX_REG_11_ | ~new_P3_ADD_546_U22;
  assign new_P3_ADD_546_U201 = ~P3_EAX_REG_10_ | ~new_P3_ADD_546_U110;
  assign new_P3_ADD_546_U202 = ~new_P3_ADD_546_U140 | ~new_P3_ADD_546_U19;
  assign new_P3_GTE_401_U6 = ~new_P3_SUB_401_U6 & ~new_P3_GTE_401_U8;
  assign new_P3_GTE_401_U7 = new_P3_SUB_401_U21 & new_P3_GTE_401_U9;
  assign new_P3_GTE_401_U8 = ~new_P3_GTE_401_U7 & ~new_P3_SUB_401_U19 & ~new_P3_SUB_401_U20;
  assign new_P3_GTE_401_U9 = new_P3_SUB_401_U7 | new_P3_SUB_401_U22;
  assign new_P3_ADD_391_1180_U4 = ~new_P3_U2613;
  assign new_P3_ADD_391_1180_U5 = ~new_P3_U3069;
  assign new_P3_ADD_391_1180_U6 = ~new_P3_U3069 | ~new_P3_U2613;
  assign new_P3_ADD_391_1180_U7 = ~new_P3_U2614;
  assign new_P3_ADD_391_1180_U8 = ~new_P3_U2614 | ~new_P3_ADD_391_1180_U28;
  assign new_P3_ADD_391_1180_U9 = ~new_P3_U2615;
  assign new_P3_ADD_391_1180_U10 = ~new_P3_U2615 | ~new_P3_ADD_391_1180_U29;
  assign new_P3_ADD_391_1180_U11 = ~new_P3_U2616;
  assign new_P3_ADD_391_1180_U12 = ~new_P3_U2616 | ~new_P3_ADD_391_1180_U30;
  assign new_P3_ADD_391_1180_U13 = ~new_P3_U2617;
  assign new_P3_ADD_391_1180_U14 = ~new_P3_U2617 | ~new_P3_ADD_391_1180_U31;
  assign new_P3_ADD_391_1180_U15 = ~new_P3_U2618;
  assign new_P3_ADD_391_1180_U16 = ~new_P3_U2618 | ~new_P3_ADD_391_1180_U32;
  assign new_P3_ADD_391_1180_U17 = ~new_P3_U2619;
  assign new_P3_ADD_391_1180_U18 = ~new_P3_ADD_391_1180_U36 | ~new_P3_ADD_391_1180_U35;
  assign new_P3_ADD_391_1180_U19 = ~new_P3_ADD_391_1180_U38 | ~new_P3_ADD_391_1180_U37;
  assign new_P3_ADD_391_1180_U20 = ~new_P3_ADD_391_1180_U40 | ~new_P3_ADD_391_1180_U39;
  assign new_P3_ADD_391_1180_U21 = ~new_P3_ADD_391_1180_U42 | ~new_P3_ADD_391_1180_U41;
  assign new_P3_ADD_391_1180_U22 = ~new_P3_ADD_391_1180_U44 | ~new_P3_ADD_391_1180_U43;
  assign new_P3_ADD_391_1180_U23 = ~new_P3_ADD_391_1180_U46 | ~new_P3_ADD_391_1180_U45;
  assign new_P3_ADD_391_1180_U24 = ~new_P3_ADD_391_1180_U48 | ~new_P3_ADD_391_1180_U47;
  assign new_P3_ADD_391_1180_U25 = ~new_P3_ADD_391_1180_U50 | ~new_P3_ADD_391_1180_U49;
  assign new_P3_ADD_391_1180_U26 = ~new_P3_U2620;
  assign new_P3_ADD_391_1180_U27 = ~new_P3_U2619 | ~new_P3_ADD_391_1180_U33;
  assign new_P3_ADD_391_1180_U28 = ~new_P3_ADD_391_1180_U6;
  assign new_P3_ADD_391_1180_U29 = ~new_P3_ADD_391_1180_U8;
  assign new_P3_ADD_391_1180_U30 = ~new_P3_ADD_391_1180_U10;
  assign new_P3_ADD_391_1180_U31 = ~new_P3_ADD_391_1180_U12;
  assign new_P3_ADD_391_1180_U32 = ~new_P3_ADD_391_1180_U14;
  assign new_P3_ADD_391_1180_U33 = ~new_P3_ADD_391_1180_U16;
  assign new_P3_ADD_391_1180_U34 = ~new_P3_ADD_391_1180_U27;
  assign new_P3_ADD_391_1180_U35 = ~new_P3_U2620 | ~new_P3_ADD_391_1180_U27;
  assign new_P3_ADD_391_1180_U36 = ~new_P3_ADD_391_1180_U34 | ~new_P3_ADD_391_1180_U26;
  assign new_P3_ADD_391_1180_U37 = ~new_P3_U2619 | ~new_P3_ADD_391_1180_U16;
  assign new_P3_ADD_391_1180_U38 = ~new_P3_ADD_391_1180_U33 | ~new_P3_ADD_391_1180_U17;
  assign new_P3_ADD_391_1180_U39 = ~new_P3_U2618 | ~new_P3_ADD_391_1180_U14;
  assign new_P3_ADD_391_1180_U40 = ~new_P3_ADD_391_1180_U32 | ~new_P3_ADD_391_1180_U15;
  assign new_P3_ADD_391_1180_U41 = ~new_P3_U2617 | ~new_P3_ADD_391_1180_U12;
  assign new_P3_ADD_391_1180_U42 = ~new_P3_ADD_391_1180_U31 | ~new_P3_ADD_391_1180_U13;
  assign new_P3_ADD_391_1180_U43 = ~new_P3_U2616 | ~new_P3_ADD_391_1180_U10;
  assign new_P3_ADD_391_1180_U44 = ~new_P3_ADD_391_1180_U30 | ~new_P3_ADD_391_1180_U11;
  assign new_P3_ADD_391_1180_U45 = ~new_P3_U2615 | ~new_P3_ADD_391_1180_U8;
  assign new_P3_ADD_391_1180_U46 = ~new_P3_ADD_391_1180_U29 | ~new_P3_ADD_391_1180_U9;
  assign new_P3_ADD_391_1180_U47 = ~new_P3_U2614 | ~new_P3_ADD_391_1180_U6;
  assign new_P3_ADD_391_1180_U48 = ~new_P3_ADD_391_1180_U28 | ~new_P3_ADD_391_1180_U7;
  assign new_P3_ADD_391_1180_U49 = ~new_P3_U3069 | ~new_P3_ADD_391_1180_U4;
  assign new_P3_ADD_391_1180_U50 = ~new_P3_U2613 | ~new_P3_ADD_391_1180_U5;
  assign new_P3_ADD_476_U4 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_476_U5 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_476_U6 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_476_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_476_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_476_U94;
  assign new_P3_ADD_476_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_476_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_476_U95;
  assign new_P3_ADD_476_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_476_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_476_U96;
  assign new_P3_ADD_476_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_476_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_476_U97;
  assign new_P3_ADD_476_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_476_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_476_U98;
  assign new_P3_ADD_476_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_476_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_476_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_476_U99;
  assign new_P3_ADD_476_U20 = ~new_P3_ADD_476_U100 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_476_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_476_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_476_U101;
  assign new_P3_ADD_476_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_476_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_476_U102;
  assign new_P3_ADD_476_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_476_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_476_U103;
  assign new_P3_ADD_476_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_476_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_476_U104;
  assign new_P3_ADD_476_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_476_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_476_U105;
  assign new_P3_ADD_476_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_476_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_476_U106;
  assign new_P3_ADD_476_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_476_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_476_U107;
  assign new_P3_ADD_476_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_476_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_476_U108;
  assign new_P3_ADD_476_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_476_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_476_U109;
  assign new_P3_ADD_476_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_476_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_476_U110;
  assign new_P3_ADD_476_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_476_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_476_U111;
  assign new_P3_ADD_476_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_476_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_476_U112;
  assign new_P3_ADD_476_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_476_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_476_U113;
  assign new_P3_ADD_476_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_476_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_476_U114;
  assign new_P3_ADD_476_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_476_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_476_U115;
  assign new_P3_ADD_476_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_476_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_476_U116;
  assign new_P3_ADD_476_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_476_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_476_U117;
  assign new_P3_ADD_476_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_476_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_476_U118;
  assign new_P3_ADD_476_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_476_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_476_U119;
  assign new_P3_ADD_476_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_476_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_476_U120;
  assign new_P3_ADD_476_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_476_U62 = ~new_P3_ADD_476_U124 | ~new_P3_ADD_476_U123;
  assign new_P3_ADD_476_U63 = ~new_P3_ADD_476_U126 | ~new_P3_ADD_476_U125;
  assign new_P3_ADD_476_U64 = ~new_P3_ADD_476_U128 | ~new_P3_ADD_476_U127;
  assign new_P3_ADD_476_U65 = ~new_P3_ADD_476_U130 | ~new_P3_ADD_476_U129;
  assign new_P3_ADD_476_U66 = ~new_P3_ADD_476_U132 | ~new_P3_ADD_476_U131;
  assign new_P3_ADD_476_U67 = ~new_P3_ADD_476_U134 | ~new_P3_ADD_476_U133;
  assign new_P3_ADD_476_U68 = ~new_P3_ADD_476_U136 | ~new_P3_ADD_476_U135;
  assign new_P3_ADD_476_U69 = ~new_P3_ADD_476_U138 | ~new_P3_ADD_476_U137;
  assign new_P3_ADD_476_U70 = ~new_P3_ADD_476_U140 | ~new_P3_ADD_476_U139;
  assign new_P3_ADD_476_U71 = ~new_P3_ADD_476_U142 | ~new_P3_ADD_476_U141;
  assign new_P3_ADD_476_U72 = ~new_P3_ADD_476_U144 | ~new_P3_ADD_476_U143;
  assign new_P3_ADD_476_U73 = ~new_P3_ADD_476_U146 | ~new_P3_ADD_476_U145;
  assign new_P3_ADD_476_U74 = ~new_P3_ADD_476_U148 | ~new_P3_ADD_476_U147;
  assign new_P3_ADD_476_U75 = ~new_P3_ADD_476_U150 | ~new_P3_ADD_476_U149;
  assign new_P3_ADD_476_U76 = ~new_P3_ADD_476_U152 | ~new_P3_ADD_476_U151;
  assign new_P3_ADD_476_U77 = ~new_P3_ADD_476_U154 | ~new_P3_ADD_476_U153;
  assign new_P3_ADD_476_U78 = ~new_P3_ADD_476_U156 | ~new_P3_ADD_476_U155;
  assign new_P3_ADD_476_U79 = ~new_P3_ADD_476_U158 | ~new_P3_ADD_476_U157;
  assign new_P3_ADD_476_U80 = ~new_P3_ADD_476_U160 | ~new_P3_ADD_476_U159;
  assign new_P3_ADD_476_U81 = ~new_P3_ADD_476_U162 | ~new_P3_ADD_476_U161;
  assign new_P3_ADD_476_U82 = ~new_P3_ADD_476_U164 | ~new_P3_ADD_476_U163;
  assign new_P3_ADD_476_U83 = ~new_P3_ADD_476_U166 | ~new_P3_ADD_476_U165;
  assign new_P3_ADD_476_U84 = ~new_P3_ADD_476_U168 | ~new_P3_ADD_476_U167;
  assign new_P3_ADD_476_U85 = ~new_P3_ADD_476_U170 | ~new_P3_ADD_476_U169;
  assign new_P3_ADD_476_U86 = ~new_P3_ADD_476_U172 | ~new_P3_ADD_476_U171;
  assign new_P3_ADD_476_U87 = ~new_P3_ADD_476_U174 | ~new_P3_ADD_476_U173;
  assign new_P3_ADD_476_U88 = ~new_P3_ADD_476_U176 | ~new_P3_ADD_476_U175;
  assign new_P3_ADD_476_U89 = ~new_P3_ADD_476_U178 | ~new_P3_ADD_476_U177;
  assign new_P3_ADD_476_U90 = ~new_P3_ADD_476_U180 | ~new_P3_ADD_476_U179;
  assign new_P3_ADD_476_U91 = ~new_P3_ADD_476_U182 | ~new_P3_ADD_476_U181;
  assign new_P3_ADD_476_U92 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_476_U93 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_476_U121;
  assign new_P3_ADD_476_U94 = ~new_P3_ADD_476_U6;
  assign new_P3_ADD_476_U95 = ~new_P3_ADD_476_U8;
  assign new_P3_ADD_476_U96 = ~new_P3_ADD_476_U10;
  assign new_P3_ADD_476_U97 = ~new_P3_ADD_476_U12;
  assign new_P3_ADD_476_U98 = ~new_P3_ADD_476_U14;
  assign new_P3_ADD_476_U99 = ~new_P3_ADD_476_U16;
  assign new_P3_ADD_476_U100 = ~new_P3_ADD_476_U19;
  assign new_P3_ADD_476_U101 = ~new_P3_ADD_476_U20;
  assign new_P3_ADD_476_U102 = ~new_P3_ADD_476_U22;
  assign new_P3_ADD_476_U103 = ~new_P3_ADD_476_U24;
  assign new_P3_ADD_476_U104 = ~new_P3_ADD_476_U26;
  assign new_P3_ADD_476_U105 = ~new_P3_ADD_476_U28;
  assign new_P3_ADD_476_U106 = ~new_P3_ADD_476_U30;
  assign new_P3_ADD_476_U107 = ~new_P3_ADD_476_U32;
  assign new_P3_ADD_476_U108 = ~new_P3_ADD_476_U34;
  assign new_P3_ADD_476_U109 = ~new_P3_ADD_476_U36;
  assign new_P3_ADD_476_U110 = ~new_P3_ADD_476_U38;
  assign new_P3_ADD_476_U111 = ~new_P3_ADD_476_U40;
  assign new_P3_ADD_476_U112 = ~new_P3_ADD_476_U42;
  assign new_P3_ADD_476_U113 = ~new_P3_ADD_476_U44;
  assign new_P3_ADD_476_U114 = ~new_P3_ADD_476_U46;
  assign new_P3_ADD_476_U115 = ~new_P3_ADD_476_U48;
  assign new_P3_ADD_476_U116 = ~new_P3_ADD_476_U50;
  assign new_P3_ADD_476_U117 = ~new_P3_ADD_476_U52;
  assign new_P3_ADD_476_U118 = ~new_P3_ADD_476_U54;
  assign new_P3_ADD_476_U119 = ~new_P3_ADD_476_U56;
  assign new_P3_ADD_476_U120 = ~new_P3_ADD_476_U58;
  assign new_P3_ADD_476_U121 = ~new_P3_ADD_476_U60;
  assign new_P3_ADD_476_U122 = ~new_P3_ADD_476_U93;
  assign new_P3_ADD_476_U123 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_476_U19;
  assign new_P3_ADD_476_U124 = ~new_P3_ADD_476_U100 | ~new_P3_ADD_476_U18;
  assign new_P3_ADD_476_U125 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_476_U16;
  assign new_P3_ADD_476_U126 = ~new_P3_ADD_476_U99 | ~new_P3_ADD_476_U17;
  assign new_P3_ADD_476_U127 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_476_U14;
  assign new_P3_ADD_476_U128 = ~new_P3_ADD_476_U98 | ~new_P3_ADD_476_U15;
  assign new_P3_ADD_476_U129 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_476_U12;
  assign new_P3_ADD_476_U130 = ~new_P3_ADD_476_U97 | ~new_P3_ADD_476_U13;
  assign new_P3_ADD_476_U131 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_476_U10;
  assign new_P3_ADD_476_U132 = ~new_P3_ADD_476_U96 | ~new_P3_ADD_476_U11;
  assign new_P3_ADD_476_U133 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_476_U8;
  assign new_P3_ADD_476_U134 = ~new_P3_ADD_476_U95 | ~new_P3_ADD_476_U9;
  assign new_P3_ADD_476_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_476_U6;
  assign new_P3_ADD_476_U136 = ~new_P3_ADD_476_U94 | ~new_P3_ADD_476_U7;
  assign new_P3_ADD_476_U137 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_476_U93;
  assign new_P3_ADD_476_U138 = ~new_P3_ADD_476_U122 | ~new_P3_ADD_476_U92;
  assign new_P3_ADD_476_U139 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_476_U60;
  assign new_P3_ADD_476_U140 = ~new_P3_ADD_476_U121 | ~new_P3_ADD_476_U61;
  assign new_P3_ADD_476_U141 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_476_U4;
  assign new_P3_ADD_476_U142 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_476_U5;
  assign new_P3_ADD_476_U143 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_476_U58;
  assign new_P3_ADD_476_U144 = ~new_P3_ADD_476_U120 | ~new_P3_ADD_476_U59;
  assign new_P3_ADD_476_U145 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_476_U56;
  assign new_P3_ADD_476_U146 = ~new_P3_ADD_476_U119 | ~new_P3_ADD_476_U57;
  assign new_P3_ADD_476_U147 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_476_U54;
  assign new_P3_ADD_476_U148 = ~new_P3_ADD_476_U118 | ~new_P3_ADD_476_U55;
  assign new_P3_ADD_476_U149 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_476_U52;
  assign new_P3_ADD_476_U150 = ~new_P3_ADD_476_U117 | ~new_P3_ADD_476_U53;
  assign new_P3_ADD_476_U151 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_476_U50;
  assign new_P3_ADD_476_U152 = ~new_P3_ADD_476_U116 | ~new_P3_ADD_476_U51;
  assign new_P3_ADD_476_U153 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_476_U48;
  assign new_P3_ADD_476_U154 = ~new_P3_ADD_476_U115 | ~new_P3_ADD_476_U49;
  assign new_P3_ADD_476_U155 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_476_U46;
  assign new_P3_ADD_476_U156 = ~new_P3_ADD_476_U114 | ~new_P3_ADD_476_U47;
  assign new_P3_ADD_476_U157 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_476_U44;
  assign new_P3_ADD_476_U158 = ~new_P3_ADD_476_U113 | ~new_P3_ADD_476_U45;
  assign new_P3_ADD_476_U159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_476_U42;
  assign new_P3_ADD_476_U160 = ~new_P3_ADD_476_U112 | ~new_P3_ADD_476_U43;
  assign new_P3_ADD_476_U161 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_476_U40;
  assign new_P3_ADD_476_U162 = ~new_P3_ADD_476_U111 | ~new_P3_ADD_476_U41;
  assign new_P3_ADD_476_U163 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_476_U38;
  assign new_P3_ADD_476_U164 = ~new_P3_ADD_476_U110 | ~new_P3_ADD_476_U39;
  assign new_P3_ADD_476_U165 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_476_U36;
  assign new_P3_ADD_476_U166 = ~new_P3_ADD_476_U109 | ~new_P3_ADD_476_U37;
  assign new_P3_ADD_476_U167 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_476_U34;
  assign new_P3_ADD_476_U168 = ~new_P3_ADD_476_U108 | ~new_P3_ADD_476_U35;
  assign new_P3_ADD_476_U169 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_476_U32;
  assign new_P3_ADD_476_U170 = ~new_P3_ADD_476_U107 | ~new_P3_ADD_476_U33;
  assign new_P3_ADD_476_U171 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_476_U30;
  assign new_P3_ADD_476_U172 = ~new_P3_ADD_476_U106 | ~new_P3_ADD_476_U31;
  assign new_P3_ADD_476_U173 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_476_U28;
  assign new_P3_ADD_476_U174 = ~new_P3_ADD_476_U105 | ~new_P3_ADD_476_U29;
  assign new_P3_ADD_476_U175 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_476_U26;
  assign new_P3_ADD_476_U176 = ~new_P3_ADD_476_U104 | ~new_P3_ADD_476_U27;
  assign new_P3_ADD_476_U177 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_476_U24;
  assign new_P3_ADD_476_U178 = ~new_P3_ADD_476_U103 | ~new_P3_ADD_476_U25;
  assign new_P3_ADD_476_U179 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_476_U22;
  assign new_P3_ADD_476_U180 = ~new_P3_ADD_476_U102 | ~new_P3_ADD_476_U23;
  assign new_P3_ADD_476_U181 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_476_U20;
  assign new_P3_ADD_476_U182 = ~new_P3_ADD_476_U101 | ~new_P3_ADD_476_U21;
  assign new_P3_GTE_390_U6 = ~new_P3_SUB_390_U6 & ~new_P3_GTE_390_U8;
  assign new_P3_GTE_390_U7 = new_P3_SUB_390_U21 & new_P3_GTE_390_U9;
  assign new_P3_GTE_390_U8 = ~new_P3_GTE_390_U7 & ~new_P3_SUB_390_U19 & ~new_P3_SUB_390_U20;
  assign new_P3_GTE_390_U9 = new_P3_SUB_390_U7 | new_P3_SUB_390_U22;
  assign new_P3_ADD_531_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_531_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_531_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_531_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_531_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_531_U98;
  assign new_P3_ADD_531_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_531_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_531_U99;
  assign new_P3_ADD_531_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_531_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_531_U100;
  assign new_P3_ADD_531_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_531_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_531_U101;
  assign new_P3_ADD_531_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_531_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_531_U102;
  assign new_P3_ADD_531_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_531_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_531_U103;
  assign new_P3_ADD_531_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_531_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_531_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_531_U104;
  assign new_P3_ADD_531_U23 = ~new_P3_ADD_531_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_531_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_531_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_531_U106;
  assign new_P3_ADD_531_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_531_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_531_U107;
  assign new_P3_ADD_531_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_531_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_531_U108;
  assign new_P3_ADD_531_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_531_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_531_U109;
  assign new_P3_ADD_531_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_531_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_531_U110;
  assign new_P3_ADD_531_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_531_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_531_U111;
  assign new_P3_ADD_531_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_531_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_531_U112;
  assign new_P3_ADD_531_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_531_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_531_U113;
  assign new_P3_ADD_531_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_531_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_531_U114;
  assign new_P3_ADD_531_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_531_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_531_U115;
  assign new_P3_ADD_531_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_531_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_531_U116;
  assign new_P3_ADD_531_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_531_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_531_U117;
  assign new_P3_ADD_531_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_531_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_531_U118;
  assign new_P3_ADD_531_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_531_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_531_U119;
  assign new_P3_ADD_531_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_531_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_531_U120;
  assign new_P3_ADD_531_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_531_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_531_U121;
  assign new_P3_ADD_531_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_531_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_531_U122;
  assign new_P3_ADD_531_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_531_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_531_U123;
  assign new_P3_ADD_531_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_531_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_531_U124;
  assign new_P3_ADD_531_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_531_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_531_U125;
  assign new_P3_ADD_531_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_531_U65 = ~new_P3_ADD_531_U129 | ~new_P3_ADD_531_U128;
  assign new_P3_ADD_531_U66 = ~new_P3_ADD_531_U131 | ~new_P3_ADD_531_U130;
  assign new_P3_ADD_531_U67 = ~new_P3_ADD_531_U133 | ~new_P3_ADD_531_U132;
  assign new_P3_ADD_531_U68 = ~new_P3_ADD_531_U135 | ~new_P3_ADD_531_U134;
  assign new_P3_ADD_531_U69 = ~new_P3_ADD_531_U137 | ~new_P3_ADD_531_U136;
  assign new_P3_ADD_531_U70 = ~new_P3_ADD_531_U139 | ~new_P3_ADD_531_U138;
  assign new_P3_ADD_531_U71 = ~new_P3_ADD_531_U141 | ~new_P3_ADD_531_U140;
  assign new_P3_ADD_531_U72 = ~new_P3_ADD_531_U143 | ~new_P3_ADD_531_U142;
  assign new_P3_ADD_531_U73 = ~new_P3_ADD_531_U145 | ~new_P3_ADD_531_U144;
  assign new_P3_ADD_531_U74 = ~new_P3_ADD_531_U147 | ~new_P3_ADD_531_U146;
  assign new_P3_ADD_531_U75 = ~new_P3_ADD_531_U149 | ~new_P3_ADD_531_U148;
  assign new_P3_ADD_531_U76 = ~new_P3_ADD_531_U151 | ~new_P3_ADD_531_U150;
  assign new_P3_ADD_531_U77 = ~new_P3_ADD_531_U153 | ~new_P3_ADD_531_U152;
  assign new_P3_ADD_531_U78 = ~new_P3_ADD_531_U155 | ~new_P3_ADD_531_U154;
  assign new_P3_ADD_531_U79 = ~new_P3_ADD_531_U157 | ~new_P3_ADD_531_U156;
  assign new_P3_ADD_531_U80 = ~new_P3_ADD_531_U159 | ~new_P3_ADD_531_U158;
  assign new_P3_ADD_531_U81 = ~new_P3_ADD_531_U161 | ~new_P3_ADD_531_U160;
  assign new_P3_ADD_531_U82 = ~new_P3_ADD_531_U163 | ~new_P3_ADD_531_U162;
  assign new_P3_ADD_531_U83 = ~new_P3_ADD_531_U165 | ~new_P3_ADD_531_U164;
  assign new_P3_ADD_531_U84 = ~new_P3_ADD_531_U167 | ~new_P3_ADD_531_U166;
  assign new_P3_ADD_531_U85 = ~new_P3_ADD_531_U169 | ~new_P3_ADD_531_U168;
  assign new_P3_ADD_531_U86 = ~new_P3_ADD_531_U171 | ~new_P3_ADD_531_U170;
  assign new_P3_ADD_531_U87 = ~new_P3_ADD_531_U173 | ~new_P3_ADD_531_U172;
  assign new_P3_ADD_531_U88 = ~new_P3_ADD_531_U175 | ~new_P3_ADD_531_U174;
  assign new_P3_ADD_531_U89 = ~new_P3_ADD_531_U177 | ~new_P3_ADD_531_U176;
  assign new_P3_ADD_531_U90 = ~new_P3_ADD_531_U179 | ~new_P3_ADD_531_U178;
  assign new_P3_ADD_531_U91 = ~new_P3_ADD_531_U181 | ~new_P3_ADD_531_U180;
  assign new_P3_ADD_531_U92 = ~new_P3_ADD_531_U183 | ~new_P3_ADD_531_U182;
  assign new_P3_ADD_531_U93 = ~new_P3_ADD_531_U185 | ~new_P3_ADD_531_U184;
  assign new_P3_ADD_531_U94 = ~new_P3_ADD_531_U187 | ~new_P3_ADD_531_U186;
  assign new_P3_ADD_531_U95 = ~new_P3_ADD_531_U189 | ~new_P3_ADD_531_U188;
  assign new_P3_ADD_531_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_531_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_531_U126;
  assign new_P3_ADD_531_U98 = ~new_P3_ADD_531_U7;
  assign new_P3_ADD_531_U99 = ~new_P3_ADD_531_U9;
  assign new_P3_ADD_531_U100 = ~new_P3_ADD_531_U11;
  assign new_P3_ADD_531_U101 = ~new_P3_ADD_531_U13;
  assign new_P3_ADD_531_U102 = ~new_P3_ADD_531_U15;
  assign new_P3_ADD_531_U103 = ~new_P3_ADD_531_U17;
  assign new_P3_ADD_531_U104 = ~new_P3_ADD_531_U19;
  assign new_P3_ADD_531_U105 = ~new_P3_ADD_531_U22;
  assign new_P3_ADD_531_U106 = ~new_P3_ADD_531_U23;
  assign new_P3_ADD_531_U107 = ~new_P3_ADD_531_U25;
  assign new_P3_ADD_531_U108 = ~new_P3_ADD_531_U27;
  assign new_P3_ADD_531_U109 = ~new_P3_ADD_531_U29;
  assign new_P3_ADD_531_U110 = ~new_P3_ADD_531_U31;
  assign new_P3_ADD_531_U111 = ~new_P3_ADD_531_U33;
  assign new_P3_ADD_531_U112 = ~new_P3_ADD_531_U35;
  assign new_P3_ADD_531_U113 = ~new_P3_ADD_531_U37;
  assign new_P3_ADD_531_U114 = ~new_P3_ADD_531_U39;
  assign new_P3_ADD_531_U115 = ~new_P3_ADD_531_U41;
  assign new_P3_ADD_531_U116 = ~new_P3_ADD_531_U43;
  assign new_P3_ADD_531_U117 = ~new_P3_ADD_531_U45;
  assign new_P3_ADD_531_U118 = ~new_P3_ADD_531_U47;
  assign new_P3_ADD_531_U119 = ~new_P3_ADD_531_U49;
  assign new_P3_ADD_531_U120 = ~new_P3_ADD_531_U51;
  assign new_P3_ADD_531_U121 = ~new_P3_ADD_531_U53;
  assign new_P3_ADD_531_U122 = ~new_P3_ADD_531_U55;
  assign new_P3_ADD_531_U123 = ~new_P3_ADD_531_U57;
  assign new_P3_ADD_531_U124 = ~new_P3_ADD_531_U59;
  assign new_P3_ADD_531_U125 = ~new_P3_ADD_531_U61;
  assign new_P3_ADD_531_U126 = ~new_P3_ADD_531_U63;
  assign new_P3_ADD_531_U127 = ~new_P3_ADD_531_U97;
  assign new_P3_ADD_531_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_531_U22;
  assign new_P3_ADD_531_U129 = ~new_P3_ADD_531_U105 | ~new_P3_ADD_531_U21;
  assign new_P3_ADD_531_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_531_U19;
  assign new_P3_ADD_531_U131 = ~new_P3_ADD_531_U104 | ~new_P3_ADD_531_U20;
  assign new_P3_ADD_531_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_531_U17;
  assign new_P3_ADD_531_U133 = ~new_P3_ADD_531_U103 | ~new_P3_ADD_531_U18;
  assign new_P3_ADD_531_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_531_U15;
  assign new_P3_ADD_531_U135 = ~new_P3_ADD_531_U102 | ~new_P3_ADD_531_U16;
  assign new_P3_ADD_531_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_531_U13;
  assign new_P3_ADD_531_U137 = ~new_P3_ADD_531_U101 | ~new_P3_ADD_531_U14;
  assign new_P3_ADD_531_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_531_U11;
  assign new_P3_ADD_531_U139 = ~new_P3_ADD_531_U100 | ~new_P3_ADD_531_U12;
  assign new_P3_ADD_531_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_531_U9;
  assign new_P3_ADD_531_U141 = ~new_P3_ADD_531_U99 | ~new_P3_ADD_531_U10;
  assign new_P3_ADD_531_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_531_U97;
  assign new_P3_ADD_531_U143 = ~new_P3_ADD_531_U127 | ~new_P3_ADD_531_U96;
  assign new_P3_ADD_531_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_531_U63;
  assign new_P3_ADD_531_U145 = ~new_P3_ADD_531_U126 | ~new_P3_ADD_531_U64;
  assign new_P3_ADD_531_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_531_U7;
  assign new_P3_ADD_531_U147 = ~new_P3_ADD_531_U98 | ~new_P3_ADD_531_U8;
  assign new_P3_ADD_531_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_531_U61;
  assign new_P3_ADD_531_U149 = ~new_P3_ADD_531_U125 | ~new_P3_ADD_531_U62;
  assign new_P3_ADD_531_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_531_U59;
  assign new_P3_ADD_531_U151 = ~new_P3_ADD_531_U124 | ~new_P3_ADD_531_U60;
  assign new_P3_ADD_531_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_531_U57;
  assign new_P3_ADD_531_U153 = ~new_P3_ADD_531_U123 | ~new_P3_ADD_531_U58;
  assign new_P3_ADD_531_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_531_U55;
  assign new_P3_ADD_531_U155 = ~new_P3_ADD_531_U122 | ~new_P3_ADD_531_U56;
  assign new_P3_ADD_531_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_531_U53;
  assign new_P3_ADD_531_U157 = ~new_P3_ADD_531_U121 | ~new_P3_ADD_531_U54;
  assign new_P3_ADD_531_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_531_U51;
  assign new_P3_ADD_531_U159 = ~new_P3_ADD_531_U120 | ~new_P3_ADD_531_U52;
  assign new_P3_ADD_531_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_531_U49;
  assign new_P3_ADD_531_U161 = ~new_P3_ADD_531_U119 | ~new_P3_ADD_531_U50;
  assign new_P3_ADD_531_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_531_U47;
  assign new_P3_ADD_531_U163 = ~new_P3_ADD_531_U118 | ~new_P3_ADD_531_U48;
  assign new_P3_ADD_531_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_531_U45;
  assign new_P3_ADD_531_U165 = ~new_P3_ADD_531_U117 | ~new_P3_ADD_531_U46;
  assign new_P3_ADD_531_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_531_U43;
  assign new_P3_ADD_531_U167 = ~new_P3_ADD_531_U116 | ~new_P3_ADD_531_U44;
  assign new_P3_ADD_531_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_531_U5;
  assign new_P3_ADD_531_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_531_U6;
  assign new_P3_ADD_531_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_531_U41;
  assign new_P3_ADD_531_U171 = ~new_P3_ADD_531_U115 | ~new_P3_ADD_531_U42;
  assign new_P3_ADD_531_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_531_U39;
  assign new_P3_ADD_531_U173 = ~new_P3_ADD_531_U114 | ~new_P3_ADD_531_U40;
  assign new_P3_ADD_531_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_531_U37;
  assign new_P3_ADD_531_U175 = ~new_P3_ADD_531_U113 | ~new_P3_ADD_531_U38;
  assign new_P3_ADD_531_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_531_U35;
  assign new_P3_ADD_531_U177 = ~new_P3_ADD_531_U112 | ~new_P3_ADD_531_U36;
  assign new_P3_ADD_531_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_531_U33;
  assign new_P3_ADD_531_U179 = ~new_P3_ADD_531_U111 | ~new_P3_ADD_531_U34;
  assign new_P3_ADD_531_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_531_U31;
  assign new_P3_ADD_531_U181 = ~new_P3_ADD_531_U110 | ~new_P3_ADD_531_U32;
  assign new_P3_ADD_531_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_531_U29;
  assign new_P3_ADD_531_U183 = ~new_P3_ADD_531_U109 | ~new_P3_ADD_531_U30;
  assign new_P3_ADD_531_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_531_U27;
  assign new_P3_ADD_531_U185 = ~new_P3_ADD_531_U108 | ~new_P3_ADD_531_U28;
  assign new_P3_ADD_531_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_531_U25;
  assign new_P3_ADD_531_U187 = ~new_P3_ADD_531_U107 | ~new_P3_ADD_531_U26;
  assign new_P3_ADD_531_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_531_U23;
  assign new_P3_ADD_531_U189 = ~new_P3_ADD_531_U106 | ~new_P3_ADD_531_U24;
  assign new_P3_SUB_320_U6 = new_P3_SUB_320_U126 & new_P3_SUB_320_U28;
  assign new_P3_SUB_320_U7 = new_P3_SUB_320_U124 & new_P3_SUB_320_U29;
  assign new_P3_SUB_320_U8 = new_P3_SUB_320_U122 & new_P3_SUB_320_U30;
  assign new_P3_SUB_320_U9 = new_P3_SUB_320_U120 & new_P3_SUB_320_U31;
  assign new_P3_SUB_320_U10 = new_P3_SUB_320_U118 & new_P3_SUB_320_U32;
  assign new_P3_SUB_320_U11 = new_P3_SUB_320_U116 & new_P3_SUB_320_U33;
  assign new_P3_SUB_320_U12 = new_P3_SUB_320_U114 & new_P3_SUB_320_U34;
  assign new_P3_SUB_320_U13 = new_P3_SUB_320_U112 & new_P3_SUB_320_U35;
  assign new_P3_SUB_320_U14 = new_P3_SUB_320_U110 & new_P3_SUB_320_U36;
  assign new_P3_SUB_320_U15 = new_P3_SUB_320_U108 & new_P3_SUB_320_U37;
  assign new_P3_SUB_320_U16 = new_P3_SUB_320_U106 & new_P3_SUB_320_U38;
  assign new_P3_SUB_320_U17 = new_P3_SUB_320_U105 & new_P3_SUB_320_U21;
  assign new_P3_SUB_320_U18 = new_P3_SUB_320_U92 & new_P3_SUB_320_U22;
  assign new_P3_SUB_320_U19 = new_P3_SUB_320_U90 & new_P3_SUB_320_U23;
  assign new_P3_SUB_320_U20 = new_P3_SUB_320_U88 & new_P3_SUB_320_U24;
  assign new_P3_SUB_320_U21 = new_P3_ADD_318_U71 | new_P3_ADD_318_U4 | P3_PHYADDRPOINTER_REG_0_;
  assign new_P3_SUB_320_U22 = ~new_P3_SUB_320_U83 | ~new_P3_SUB_320_U27 | ~new_P3_SUB_320_U58;
  assign new_P3_SUB_320_U23 = ~new_P3_SUB_320_U84 | ~new_P3_SUB_320_U26 | ~new_P3_SUB_320_U56;
  assign new_P3_SUB_320_U24 = ~new_P3_SUB_320_U85 | ~new_P3_SUB_320_U25 | ~new_P3_SUB_320_U54;
  assign new_P3_SUB_320_U25 = ~new_P3_ADD_318_U63;
  assign new_P3_SUB_320_U26 = ~new_P3_ADD_318_U65;
  assign new_P3_SUB_320_U27 = ~new_P3_ADD_318_U67;
  assign new_P3_SUB_320_U28 = ~new_P3_SUB_320_U86 | ~new_P3_SUB_320_U52 | ~new_P3_SUB_320_U49;
  assign new_P3_SUB_320_U29 = ~new_P3_SUB_320_U93 | ~new_P3_SUB_320_U48 | ~new_P3_SUB_320_U81;
  assign new_P3_SUB_320_U30 = ~new_P3_SUB_320_U94 | ~new_P3_SUB_320_U47 | ~new_P3_SUB_320_U79;
  assign new_P3_SUB_320_U31 = ~new_P3_SUB_320_U95 | ~new_P3_SUB_320_U46 | ~new_P3_SUB_320_U77;
  assign new_P3_SUB_320_U32 = ~new_P3_SUB_320_U96 | ~new_P3_SUB_320_U45 | ~new_P3_SUB_320_U75;
  assign new_P3_SUB_320_U33 = ~new_P3_SUB_320_U97 | ~new_P3_SUB_320_U44 | ~new_P3_SUB_320_U73;
  assign new_P3_SUB_320_U34 = ~new_P3_SUB_320_U98 | ~new_P3_SUB_320_U43 | ~new_P3_SUB_320_U69;
  assign new_P3_SUB_320_U35 = ~new_P3_SUB_320_U99 | ~new_P3_SUB_320_U42 | ~new_P3_SUB_320_U67;
  assign new_P3_SUB_320_U36 = ~new_P3_SUB_320_U100 | ~new_P3_SUB_320_U41 | ~new_P3_SUB_320_U65;
  assign new_P3_SUB_320_U37 = ~new_P3_SUB_320_U101 | ~new_P3_SUB_320_U40 | ~new_P3_SUB_320_U63;
  assign new_P3_SUB_320_U38 = ~new_P3_SUB_320_U102 | ~new_P3_SUB_320_U39;
  assign new_P3_SUB_320_U39 = ~new_P3_ADD_318_U72;
  assign new_P3_SUB_320_U40 = ~new_P3_ADD_318_U73;
  assign new_P3_SUB_320_U41 = ~new_P3_ADD_318_U75;
  assign new_P3_SUB_320_U42 = ~new_P3_ADD_318_U77;
  assign new_P3_SUB_320_U43 = ~new_P3_ADD_318_U79;
  assign new_P3_SUB_320_U44 = ~new_P3_ADD_318_U81;
  assign new_P3_SUB_320_U45 = ~new_P3_ADD_318_U83;
  assign new_P3_SUB_320_U46 = ~new_P3_ADD_318_U85;
  assign new_P3_SUB_320_U47 = ~new_P3_ADD_318_U87;
  assign new_P3_SUB_320_U48 = ~new_P3_ADD_318_U89;
  assign new_P3_SUB_320_U49 = ~new_P3_ADD_318_U91;
  assign new_P3_SUB_320_U50 = ~new_P3_SUB_320_U149 | ~new_P3_SUB_320_U148;
  assign new_P3_SUB_320_U51 = ~new_P3_SUB_320_U137 | ~new_P3_SUB_320_U136;
  assign new_P3_SUB_320_U52 = ~new_P3_ADD_318_U62;
  assign new_P3_SUB_320_U53 = new_P3_SUB_320_U129 & new_P3_SUB_320_U128;
  assign new_P3_SUB_320_U54 = ~new_P3_ADD_318_U64;
  assign new_P3_SUB_320_U55 = new_P3_SUB_320_U131 & new_P3_SUB_320_U130;
  assign new_P3_SUB_320_U56 = ~new_P3_ADD_318_U66;
  assign new_P3_SUB_320_U57 = new_P3_SUB_320_U133 & new_P3_SUB_320_U132;
  assign new_P3_SUB_320_U58 = ~new_P3_ADD_318_U68;
  assign new_P3_SUB_320_U59 = new_P3_SUB_320_U135 & new_P3_SUB_320_U134;
  assign new_P3_SUB_320_U60 = ~new_P3_ADD_318_U69;
  assign new_P3_SUB_320_U61 = ~new_P3_ADD_318_U70;
  assign new_P3_SUB_320_U62 = new_P3_SUB_320_U139 & new_P3_SUB_320_U138;
  assign new_P3_SUB_320_U63 = ~new_P3_ADD_318_U74;
  assign new_P3_SUB_320_U64 = new_P3_SUB_320_U141 & new_P3_SUB_320_U140;
  assign new_P3_SUB_320_U65 = ~new_P3_ADD_318_U76;
  assign new_P3_SUB_320_U66 = new_P3_SUB_320_U143 & new_P3_SUB_320_U142;
  assign new_P3_SUB_320_U67 = ~new_P3_ADD_318_U78;
  assign new_P3_SUB_320_U68 = new_P3_SUB_320_U145 & new_P3_SUB_320_U144;
  assign new_P3_SUB_320_U69 = ~new_P3_ADD_318_U80;
  assign new_P3_SUB_320_U70 = new_P3_SUB_320_U147 & new_P3_SUB_320_U146;
  assign new_P3_SUB_320_U71 = ~new_P3_ADD_318_U4;
  assign new_P3_SUB_320_U72 = ~P3_PHYADDRPOINTER_REG_0_;
  assign new_P3_SUB_320_U73 = ~new_P3_ADD_318_U82;
  assign new_P3_SUB_320_U74 = new_P3_SUB_320_U151 & new_P3_SUB_320_U150;
  assign new_P3_SUB_320_U75 = ~new_P3_ADD_318_U84;
  assign new_P3_SUB_320_U76 = new_P3_SUB_320_U153 & new_P3_SUB_320_U152;
  assign new_P3_SUB_320_U77 = ~new_P3_ADD_318_U86;
  assign new_P3_SUB_320_U78 = new_P3_SUB_320_U155 & new_P3_SUB_320_U154;
  assign new_P3_SUB_320_U79 = ~new_P3_ADD_318_U88;
  assign new_P3_SUB_320_U80 = new_P3_SUB_320_U157 & new_P3_SUB_320_U156;
  assign new_P3_SUB_320_U81 = ~new_P3_ADD_318_U90;
  assign new_P3_SUB_320_U82 = new_P3_SUB_320_U159 & new_P3_SUB_320_U158;
  assign new_P3_SUB_320_U83 = ~new_P3_SUB_320_U21;
  assign new_P3_SUB_320_U84 = ~new_P3_SUB_320_U22;
  assign new_P3_SUB_320_U85 = ~new_P3_SUB_320_U23;
  assign new_P3_SUB_320_U86 = ~new_P3_SUB_320_U24;
  assign new_P3_SUB_320_U87 = ~new_P3_SUB_320_U85 | ~new_P3_SUB_320_U54;
  assign new_P3_SUB_320_U88 = ~new_P3_ADD_318_U63 | ~new_P3_SUB_320_U87;
  assign new_P3_SUB_320_U89 = ~new_P3_SUB_320_U84 | ~new_P3_SUB_320_U56;
  assign new_P3_SUB_320_U90 = ~new_P3_ADD_318_U65 | ~new_P3_SUB_320_U89;
  assign new_P3_SUB_320_U91 = ~new_P3_SUB_320_U83 | ~new_P3_SUB_320_U58;
  assign new_P3_SUB_320_U92 = ~new_P3_ADD_318_U67 | ~new_P3_SUB_320_U91;
  assign new_P3_SUB_320_U93 = ~new_P3_SUB_320_U28;
  assign new_P3_SUB_320_U94 = ~new_P3_SUB_320_U29;
  assign new_P3_SUB_320_U95 = ~new_P3_SUB_320_U30;
  assign new_P3_SUB_320_U96 = ~new_P3_SUB_320_U31;
  assign new_P3_SUB_320_U97 = ~new_P3_SUB_320_U32;
  assign new_P3_SUB_320_U98 = ~new_P3_SUB_320_U33;
  assign new_P3_SUB_320_U99 = ~new_P3_SUB_320_U34;
  assign new_P3_SUB_320_U100 = ~new_P3_SUB_320_U35;
  assign new_P3_SUB_320_U101 = ~new_P3_SUB_320_U36;
  assign new_P3_SUB_320_U102 = ~new_P3_SUB_320_U37;
  assign new_P3_SUB_320_U103 = ~new_P3_SUB_320_U38;
  assign new_P3_SUB_320_U104 = new_P3_ADD_318_U4 | P3_PHYADDRPOINTER_REG_0_;
  assign new_P3_SUB_320_U105 = ~new_P3_ADD_318_U71 | ~new_P3_SUB_320_U104;
  assign new_P3_SUB_320_U106 = ~new_P3_ADD_318_U72 | ~new_P3_SUB_320_U37;
  assign new_P3_SUB_320_U107 = ~new_P3_SUB_320_U101 | ~new_P3_SUB_320_U63;
  assign new_P3_SUB_320_U108 = ~new_P3_ADD_318_U73 | ~new_P3_SUB_320_U107;
  assign new_P3_SUB_320_U109 = ~new_P3_SUB_320_U100 | ~new_P3_SUB_320_U65;
  assign new_P3_SUB_320_U110 = ~new_P3_ADD_318_U75 | ~new_P3_SUB_320_U109;
  assign new_P3_SUB_320_U111 = ~new_P3_SUB_320_U99 | ~new_P3_SUB_320_U67;
  assign new_P3_SUB_320_U112 = ~new_P3_ADD_318_U77 | ~new_P3_SUB_320_U111;
  assign new_P3_SUB_320_U113 = ~new_P3_SUB_320_U98 | ~new_P3_SUB_320_U69;
  assign new_P3_SUB_320_U114 = ~new_P3_ADD_318_U79 | ~new_P3_SUB_320_U113;
  assign new_P3_SUB_320_U115 = ~new_P3_SUB_320_U97 | ~new_P3_SUB_320_U73;
  assign new_P3_SUB_320_U116 = ~new_P3_ADD_318_U81 | ~new_P3_SUB_320_U115;
  assign new_P3_SUB_320_U117 = ~new_P3_SUB_320_U96 | ~new_P3_SUB_320_U75;
  assign new_P3_SUB_320_U118 = ~new_P3_ADD_318_U83 | ~new_P3_SUB_320_U117;
  assign new_P3_SUB_320_U119 = ~new_P3_SUB_320_U95 | ~new_P3_SUB_320_U77;
  assign new_P3_SUB_320_U120 = ~new_P3_ADD_318_U85 | ~new_P3_SUB_320_U119;
  assign new_P3_SUB_320_U121 = ~new_P3_SUB_320_U94 | ~new_P3_SUB_320_U79;
  assign new_P3_SUB_320_U122 = ~new_P3_ADD_318_U87 | ~new_P3_SUB_320_U121;
  assign new_P3_SUB_320_U123 = ~new_P3_SUB_320_U93 | ~new_P3_SUB_320_U81;
  assign new_P3_SUB_320_U124 = ~new_P3_ADD_318_U89 | ~new_P3_SUB_320_U123;
  assign new_P3_SUB_320_U125 = ~new_P3_SUB_320_U86 | ~new_P3_SUB_320_U52;
  assign new_P3_SUB_320_U126 = ~new_P3_ADD_318_U91 | ~new_P3_SUB_320_U125;
  assign new_P3_SUB_320_U127 = ~new_P3_SUB_320_U103 | ~new_P3_SUB_320_U61;
  assign new_P3_SUB_320_U128 = ~new_P3_ADD_318_U62 | ~new_P3_SUB_320_U24;
  assign new_P3_SUB_320_U129 = ~new_P3_SUB_320_U86 | ~new_P3_SUB_320_U52;
  assign new_P3_SUB_320_U130 = ~new_P3_ADD_318_U64 | ~new_P3_SUB_320_U23;
  assign new_P3_SUB_320_U131 = ~new_P3_SUB_320_U85 | ~new_P3_SUB_320_U54;
  assign new_P3_SUB_320_U132 = ~new_P3_ADD_318_U66 | ~new_P3_SUB_320_U22;
  assign new_P3_SUB_320_U133 = ~new_P3_SUB_320_U84 | ~new_P3_SUB_320_U56;
  assign new_P3_SUB_320_U134 = ~new_P3_ADD_318_U68 | ~new_P3_SUB_320_U21;
  assign new_P3_SUB_320_U135 = ~new_P3_SUB_320_U83 | ~new_P3_SUB_320_U58;
  assign new_P3_SUB_320_U136 = ~new_P3_SUB_320_U127 | ~new_P3_SUB_320_U60;
  assign new_P3_SUB_320_U137 = ~new_P3_ADD_318_U69 | ~new_P3_SUB_320_U103 | ~new_P3_SUB_320_U61;
  assign new_P3_SUB_320_U138 = ~new_P3_ADD_318_U70 | ~new_P3_SUB_320_U38;
  assign new_P3_SUB_320_U139 = ~new_P3_SUB_320_U103 | ~new_P3_SUB_320_U61;
  assign new_P3_SUB_320_U140 = ~new_P3_ADD_318_U74 | ~new_P3_SUB_320_U36;
  assign new_P3_SUB_320_U141 = ~new_P3_SUB_320_U101 | ~new_P3_SUB_320_U63;
  assign new_P3_SUB_320_U142 = ~new_P3_ADD_318_U76 | ~new_P3_SUB_320_U35;
  assign new_P3_SUB_320_U143 = ~new_P3_SUB_320_U100 | ~new_P3_SUB_320_U65;
  assign new_P3_SUB_320_U144 = ~new_P3_ADD_318_U78 | ~new_P3_SUB_320_U34;
  assign new_P3_SUB_320_U145 = ~new_P3_SUB_320_U99 | ~new_P3_SUB_320_U67;
  assign new_P3_SUB_320_U146 = ~new_P3_ADD_318_U80 | ~new_P3_SUB_320_U33;
  assign new_P3_SUB_320_U147 = ~new_P3_SUB_320_U98 | ~new_P3_SUB_320_U69;
  assign new_P3_SUB_320_U148 = ~new_P3_ADD_318_U4 | ~new_P3_SUB_320_U72;
  assign new_P3_SUB_320_U149 = ~P3_PHYADDRPOINTER_REG_0_ | ~new_P3_SUB_320_U71;
  assign new_P3_SUB_320_U150 = ~new_P3_ADD_318_U82 | ~new_P3_SUB_320_U32;
  assign new_P3_SUB_320_U151 = ~new_P3_SUB_320_U97 | ~new_P3_SUB_320_U73;
  assign new_P3_SUB_320_U152 = ~new_P3_ADD_318_U84 | ~new_P3_SUB_320_U31;
  assign new_P3_SUB_320_U153 = ~new_P3_SUB_320_U96 | ~new_P3_SUB_320_U75;
  assign new_P3_SUB_320_U154 = ~new_P3_ADD_318_U86 | ~new_P3_SUB_320_U30;
  assign new_P3_SUB_320_U155 = ~new_P3_SUB_320_U95 | ~new_P3_SUB_320_U77;
  assign new_P3_SUB_320_U156 = ~new_P3_ADD_318_U88 | ~new_P3_SUB_320_U29;
  assign new_P3_SUB_320_U157 = ~new_P3_SUB_320_U94 | ~new_P3_SUB_320_U79;
  assign new_P3_SUB_320_U158 = ~new_P3_ADD_318_U90 | ~new_P3_SUB_320_U28;
  assign new_P3_SUB_320_U159 = ~new_P3_SUB_320_U93 | ~new_P3_SUB_320_U81;
  assign new_P3_ADD_505_U5 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_ADD_505_U6 = P3_INSTQUEUERD_ADDR_REG_4_ & new_P3_ADD_505_U20;
  assign new_P3_ADD_505_U7 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_ADD_505_U8 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_ADD_505_U9 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_ADD_505_U10 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_ADD_505_U18;
  assign new_P3_ADD_505_U11 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_ADD_505_U12 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_ADD_505_U19;
  assign new_P3_ADD_505_U13 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_ADD_505_U14 = ~new_P3_ADD_505_U22 | ~new_P3_ADD_505_U21;
  assign new_P3_ADD_505_U15 = ~new_P3_ADD_505_U24 | ~new_P3_ADD_505_U23;
  assign new_P3_ADD_505_U16 = ~new_P3_ADD_505_U26 | ~new_P3_ADD_505_U25;
  assign new_P3_ADD_505_U17 = ~new_P3_ADD_505_U28 | ~new_P3_ADD_505_U27;
  assign new_P3_ADD_505_U18 = ~new_P3_ADD_505_U8;
  assign new_P3_ADD_505_U19 = ~new_P3_ADD_505_U10;
  assign new_P3_ADD_505_U20 = ~new_P3_ADD_505_U12;
  assign new_P3_ADD_505_U21 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_ADD_505_U12;
  assign new_P3_ADD_505_U22 = ~new_P3_ADD_505_U20 | ~new_P3_ADD_505_U13;
  assign new_P3_ADD_505_U23 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_ADD_505_U10;
  assign new_P3_ADD_505_U24 = ~new_P3_ADD_505_U19 | ~new_P3_ADD_505_U11;
  assign new_P3_ADD_505_U25 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_ADD_505_U8;
  assign new_P3_ADD_505_U26 = ~new_P3_ADD_505_U18 | ~new_P3_ADD_505_U9;
  assign new_P3_ADD_505_U27 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_ADD_505_U5;
  assign new_P3_ADD_505_U28 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_ADD_505_U7;
  assign new_P3_GTE_485_U6 = ~new_P3_SUB_485_U6 & ~new_P3_GTE_485_U7;
  assign new_P3_GTE_485_U7 = ~new_P3_SUB_485_U18 & ~new_P3_SUB_485_U19 & ~new_P3_SUB_485_U16 & ~new_P3_SUB_485_U17;
  assign new_P3_ADD_318_U4 = ~P3_PHYADDRPOINTER_REG_1_;
  assign new_P3_ADD_318_U5 = ~P3_PHYADDRPOINTER_REG_2_;
  assign new_P3_ADD_318_U6 = ~P3_PHYADDRPOINTER_REG_2_ | ~P3_PHYADDRPOINTER_REG_1_;
  assign new_P3_ADD_318_U7 = ~P3_PHYADDRPOINTER_REG_3_;
  assign new_P3_ADD_318_U8 = ~P3_PHYADDRPOINTER_REG_3_ | ~new_P3_ADD_318_U94;
  assign new_P3_ADD_318_U9 = ~P3_PHYADDRPOINTER_REG_4_;
  assign new_P3_ADD_318_U10 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_ADD_318_U95;
  assign new_P3_ADD_318_U11 = ~P3_PHYADDRPOINTER_REG_5_;
  assign new_P3_ADD_318_U12 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_ADD_318_U96;
  assign new_P3_ADD_318_U13 = ~P3_PHYADDRPOINTER_REG_6_;
  assign new_P3_ADD_318_U14 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_ADD_318_U97;
  assign new_P3_ADD_318_U15 = ~P3_PHYADDRPOINTER_REG_7_;
  assign new_P3_ADD_318_U16 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_ADD_318_U98;
  assign new_P3_ADD_318_U17 = ~P3_PHYADDRPOINTER_REG_8_;
  assign new_P3_ADD_318_U18 = ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_ADD_318_U19 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_ADD_318_U99;
  assign new_P3_ADD_318_U20 = ~new_P3_ADD_318_U100 | ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_ADD_318_U21 = ~P3_PHYADDRPOINTER_REG_10_;
  assign new_P3_ADD_318_U22 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_ADD_318_U101;
  assign new_P3_ADD_318_U23 = ~P3_PHYADDRPOINTER_REG_11_;
  assign new_P3_ADD_318_U24 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_ADD_318_U102;
  assign new_P3_ADD_318_U25 = ~P3_PHYADDRPOINTER_REG_12_;
  assign new_P3_ADD_318_U26 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_ADD_318_U103;
  assign new_P3_ADD_318_U27 = ~P3_PHYADDRPOINTER_REG_13_;
  assign new_P3_ADD_318_U28 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_ADD_318_U104;
  assign new_P3_ADD_318_U29 = ~P3_PHYADDRPOINTER_REG_14_;
  assign new_P3_ADD_318_U30 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_ADD_318_U105;
  assign new_P3_ADD_318_U31 = ~P3_PHYADDRPOINTER_REG_15_;
  assign new_P3_ADD_318_U32 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_ADD_318_U106;
  assign new_P3_ADD_318_U33 = ~P3_PHYADDRPOINTER_REG_16_;
  assign new_P3_ADD_318_U34 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_ADD_318_U107;
  assign new_P3_ADD_318_U35 = ~P3_PHYADDRPOINTER_REG_17_;
  assign new_P3_ADD_318_U36 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_ADD_318_U108;
  assign new_P3_ADD_318_U37 = ~P3_PHYADDRPOINTER_REG_18_;
  assign new_P3_ADD_318_U38 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_ADD_318_U109;
  assign new_P3_ADD_318_U39 = ~P3_PHYADDRPOINTER_REG_19_;
  assign new_P3_ADD_318_U40 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_ADD_318_U110;
  assign new_P3_ADD_318_U41 = ~P3_PHYADDRPOINTER_REG_20_;
  assign new_P3_ADD_318_U42 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_ADD_318_U111;
  assign new_P3_ADD_318_U43 = ~P3_PHYADDRPOINTER_REG_21_;
  assign new_P3_ADD_318_U44 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_ADD_318_U112;
  assign new_P3_ADD_318_U45 = ~P3_PHYADDRPOINTER_REG_22_;
  assign new_P3_ADD_318_U46 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_ADD_318_U113;
  assign new_P3_ADD_318_U47 = ~P3_PHYADDRPOINTER_REG_23_;
  assign new_P3_ADD_318_U48 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_ADD_318_U114;
  assign new_P3_ADD_318_U49 = ~P3_PHYADDRPOINTER_REG_24_;
  assign new_P3_ADD_318_U50 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_ADD_318_U115;
  assign new_P3_ADD_318_U51 = ~P3_PHYADDRPOINTER_REG_25_;
  assign new_P3_ADD_318_U52 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_ADD_318_U116;
  assign new_P3_ADD_318_U53 = ~P3_PHYADDRPOINTER_REG_26_;
  assign new_P3_ADD_318_U54 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_ADD_318_U117;
  assign new_P3_ADD_318_U55 = ~P3_PHYADDRPOINTER_REG_27_;
  assign new_P3_ADD_318_U56 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_ADD_318_U118;
  assign new_P3_ADD_318_U57 = ~P3_PHYADDRPOINTER_REG_28_;
  assign new_P3_ADD_318_U58 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_ADD_318_U119;
  assign new_P3_ADD_318_U59 = ~P3_PHYADDRPOINTER_REG_29_;
  assign new_P3_ADD_318_U60 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_ADD_318_U120;
  assign new_P3_ADD_318_U61 = ~P3_PHYADDRPOINTER_REG_30_;
  assign new_P3_ADD_318_U62 = ~new_P3_ADD_318_U124 | ~new_P3_ADD_318_U123;
  assign new_P3_ADD_318_U63 = ~new_P3_ADD_318_U126 | ~new_P3_ADD_318_U125;
  assign new_P3_ADD_318_U64 = ~new_P3_ADD_318_U128 | ~new_P3_ADD_318_U127;
  assign new_P3_ADD_318_U65 = ~new_P3_ADD_318_U130 | ~new_P3_ADD_318_U129;
  assign new_P3_ADD_318_U66 = ~new_P3_ADD_318_U132 | ~new_P3_ADD_318_U131;
  assign new_P3_ADD_318_U67 = ~new_P3_ADD_318_U134 | ~new_P3_ADD_318_U133;
  assign new_P3_ADD_318_U68 = ~new_P3_ADD_318_U136 | ~new_P3_ADD_318_U135;
  assign new_P3_ADD_318_U69 = ~new_P3_ADD_318_U138 | ~new_P3_ADD_318_U137;
  assign new_P3_ADD_318_U70 = ~new_P3_ADD_318_U140 | ~new_P3_ADD_318_U139;
  assign new_P3_ADD_318_U71 = ~new_P3_ADD_318_U142 | ~new_P3_ADD_318_U141;
  assign new_P3_ADD_318_U72 = ~new_P3_ADD_318_U144 | ~new_P3_ADD_318_U143;
  assign new_P3_ADD_318_U73 = ~new_P3_ADD_318_U146 | ~new_P3_ADD_318_U145;
  assign new_P3_ADD_318_U74 = ~new_P3_ADD_318_U148 | ~new_P3_ADD_318_U147;
  assign new_P3_ADD_318_U75 = ~new_P3_ADD_318_U150 | ~new_P3_ADD_318_U149;
  assign new_P3_ADD_318_U76 = ~new_P3_ADD_318_U152 | ~new_P3_ADD_318_U151;
  assign new_P3_ADD_318_U77 = ~new_P3_ADD_318_U154 | ~new_P3_ADD_318_U153;
  assign new_P3_ADD_318_U78 = ~new_P3_ADD_318_U156 | ~new_P3_ADD_318_U155;
  assign new_P3_ADD_318_U79 = ~new_P3_ADD_318_U158 | ~new_P3_ADD_318_U157;
  assign new_P3_ADD_318_U80 = ~new_P3_ADD_318_U160 | ~new_P3_ADD_318_U159;
  assign new_P3_ADD_318_U81 = ~new_P3_ADD_318_U162 | ~new_P3_ADD_318_U161;
  assign new_P3_ADD_318_U82 = ~new_P3_ADD_318_U164 | ~new_P3_ADD_318_U163;
  assign new_P3_ADD_318_U83 = ~new_P3_ADD_318_U166 | ~new_P3_ADD_318_U165;
  assign new_P3_ADD_318_U84 = ~new_P3_ADD_318_U168 | ~new_P3_ADD_318_U167;
  assign new_P3_ADD_318_U85 = ~new_P3_ADD_318_U170 | ~new_P3_ADD_318_U169;
  assign new_P3_ADD_318_U86 = ~new_P3_ADD_318_U172 | ~new_P3_ADD_318_U171;
  assign new_P3_ADD_318_U87 = ~new_P3_ADD_318_U174 | ~new_P3_ADD_318_U173;
  assign new_P3_ADD_318_U88 = ~new_P3_ADD_318_U176 | ~new_P3_ADD_318_U175;
  assign new_P3_ADD_318_U89 = ~new_P3_ADD_318_U178 | ~new_P3_ADD_318_U177;
  assign new_P3_ADD_318_U90 = ~new_P3_ADD_318_U180 | ~new_P3_ADD_318_U179;
  assign new_P3_ADD_318_U91 = ~new_P3_ADD_318_U182 | ~new_P3_ADD_318_U181;
  assign new_P3_ADD_318_U92 = ~P3_PHYADDRPOINTER_REG_31_;
  assign new_P3_ADD_318_U93 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_ADD_318_U121;
  assign new_P3_ADD_318_U94 = ~new_P3_ADD_318_U6;
  assign new_P3_ADD_318_U95 = ~new_P3_ADD_318_U8;
  assign new_P3_ADD_318_U96 = ~new_P3_ADD_318_U10;
  assign new_P3_ADD_318_U97 = ~new_P3_ADD_318_U12;
  assign new_P3_ADD_318_U98 = ~new_P3_ADD_318_U14;
  assign new_P3_ADD_318_U99 = ~new_P3_ADD_318_U16;
  assign new_P3_ADD_318_U100 = ~new_P3_ADD_318_U19;
  assign new_P3_ADD_318_U101 = ~new_P3_ADD_318_U20;
  assign new_P3_ADD_318_U102 = ~new_P3_ADD_318_U22;
  assign new_P3_ADD_318_U103 = ~new_P3_ADD_318_U24;
  assign new_P3_ADD_318_U104 = ~new_P3_ADD_318_U26;
  assign new_P3_ADD_318_U105 = ~new_P3_ADD_318_U28;
  assign new_P3_ADD_318_U106 = ~new_P3_ADD_318_U30;
  assign new_P3_ADD_318_U107 = ~new_P3_ADD_318_U32;
  assign new_P3_ADD_318_U108 = ~new_P3_ADD_318_U34;
  assign new_P3_ADD_318_U109 = ~new_P3_ADD_318_U36;
  assign new_P3_ADD_318_U110 = ~new_P3_ADD_318_U38;
  assign new_P3_ADD_318_U111 = ~new_P3_ADD_318_U40;
  assign new_P3_ADD_318_U112 = ~new_P3_ADD_318_U42;
  assign new_P3_ADD_318_U113 = ~new_P3_ADD_318_U44;
  assign new_P3_ADD_318_U114 = ~new_P3_ADD_318_U46;
  assign new_P3_ADD_318_U115 = ~new_P3_ADD_318_U48;
  assign new_P3_ADD_318_U116 = ~new_P3_ADD_318_U50;
  assign new_P3_ADD_318_U117 = ~new_P3_ADD_318_U52;
  assign new_P3_ADD_318_U118 = ~new_P3_ADD_318_U54;
  assign new_P3_ADD_318_U119 = ~new_P3_ADD_318_U56;
  assign new_P3_ADD_318_U120 = ~new_P3_ADD_318_U58;
  assign new_P3_ADD_318_U121 = ~new_P3_ADD_318_U60;
  assign new_P3_ADD_318_U122 = ~new_P3_ADD_318_U93;
  assign new_P3_ADD_318_U123 = ~P3_PHYADDRPOINTER_REG_9_ | ~new_P3_ADD_318_U19;
  assign new_P3_ADD_318_U124 = ~new_P3_ADD_318_U100 | ~new_P3_ADD_318_U18;
  assign new_P3_ADD_318_U125 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_ADD_318_U16;
  assign new_P3_ADD_318_U126 = ~new_P3_ADD_318_U99 | ~new_P3_ADD_318_U17;
  assign new_P3_ADD_318_U127 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_ADD_318_U14;
  assign new_P3_ADD_318_U128 = ~new_P3_ADD_318_U98 | ~new_P3_ADD_318_U15;
  assign new_P3_ADD_318_U129 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_ADD_318_U12;
  assign new_P3_ADD_318_U130 = ~new_P3_ADD_318_U97 | ~new_P3_ADD_318_U13;
  assign new_P3_ADD_318_U131 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_ADD_318_U10;
  assign new_P3_ADD_318_U132 = ~new_P3_ADD_318_U96 | ~new_P3_ADD_318_U11;
  assign new_P3_ADD_318_U133 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_ADD_318_U8;
  assign new_P3_ADD_318_U134 = ~new_P3_ADD_318_U95 | ~new_P3_ADD_318_U9;
  assign new_P3_ADD_318_U135 = ~P3_PHYADDRPOINTER_REG_3_ | ~new_P3_ADD_318_U6;
  assign new_P3_ADD_318_U136 = ~new_P3_ADD_318_U94 | ~new_P3_ADD_318_U7;
  assign new_P3_ADD_318_U137 = ~P3_PHYADDRPOINTER_REG_31_ | ~new_P3_ADD_318_U93;
  assign new_P3_ADD_318_U138 = ~new_P3_ADD_318_U122 | ~new_P3_ADD_318_U92;
  assign new_P3_ADD_318_U139 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_ADD_318_U60;
  assign new_P3_ADD_318_U140 = ~new_P3_ADD_318_U121 | ~new_P3_ADD_318_U61;
  assign new_P3_ADD_318_U141 = ~P3_PHYADDRPOINTER_REG_2_ | ~new_P3_ADD_318_U4;
  assign new_P3_ADD_318_U142 = ~P3_PHYADDRPOINTER_REG_1_ | ~new_P3_ADD_318_U5;
  assign new_P3_ADD_318_U143 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_ADD_318_U58;
  assign new_P3_ADD_318_U144 = ~new_P3_ADD_318_U120 | ~new_P3_ADD_318_U59;
  assign new_P3_ADD_318_U145 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_ADD_318_U56;
  assign new_P3_ADD_318_U146 = ~new_P3_ADD_318_U119 | ~new_P3_ADD_318_U57;
  assign new_P3_ADD_318_U147 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_ADD_318_U54;
  assign new_P3_ADD_318_U148 = ~new_P3_ADD_318_U118 | ~new_P3_ADD_318_U55;
  assign new_P3_ADD_318_U149 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_ADD_318_U52;
  assign new_P3_ADD_318_U150 = ~new_P3_ADD_318_U117 | ~new_P3_ADD_318_U53;
  assign new_P3_ADD_318_U151 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_ADD_318_U50;
  assign new_P3_ADD_318_U152 = ~new_P3_ADD_318_U116 | ~new_P3_ADD_318_U51;
  assign new_P3_ADD_318_U153 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_ADD_318_U48;
  assign new_P3_ADD_318_U154 = ~new_P3_ADD_318_U115 | ~new_P3_ADD_318_U49;
  assign new_P3_ADD_318_U155 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_ADD_318_U46;
  assign new_P3_ADD_318_U156 = ~new_P3_ADD_318_U114 | ~new_P3_ADD_318_U47;
  assign new_P3_ADD_318_U157 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_ADD_318_U44;
  assign new_P3_ADD_318_U158 = ~new_P3_ADD_318_U113 | ~new_P3_ADD_318_U45;
  assign new_P3_ADD_318_U159 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_ADD_318_U42;
  assign new_P3_ADD_318_U160 = ~new_P3_ADD_318_U112 | ~new_P3_ADD_318_U43;
  assign new_P3_ADD_318_U161 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_ADD_318_U40;
  assign new_P3_ADD_318_U162 = ~new_P3_ADD_318_U111 | ~new_P3_ADD_318_U41;
  assign new_P3_ADD_318_U163 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_ADD_318_U38;
  assign new_P3_ADD_318_U164 = ~new_P3_ADD_318_U110 | ~new_P3_ADD_318_U39;
  assign new_P3_ADD_318_U165 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_ADD_318_U36;
  assign new_P3_ADD_318_U166 = ~new_P3_ADD_318_U109 | ~new_P3_ADD_318_U37;
  assign new_P3_ADD_318_U167 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_ADD_318_U34;
  assign new_P3_ADD_318_U168 = ~new_P3_ADD_318_U108 | ~new_P3_ADD_318_U35;
  assign new_P3_ADD_318_U169 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_ADD_318_U32;
  assign new_P3_ADD_318_U170 = ~new_P3_ADD_318_U107 | ~new_P3_ADD_318_U33;
  assign new_P3_ADD_318_U171 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_ADD_318_U30;
  assign new_P3_ADD_318_U172 = ~new_P3_ADD_318_U106 | ~new_P3_ADD_318_U31;
  assign new_P3_ADD_318_U173 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_ADD_318_U28;
  assign new_P3_ADD_318_U174 = ~new_P3_ADD_318_U105 | ~new_P3_ADD_318_U29;
  assign new_P3_ADD_318_U175 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_ADD_318_U26;
  assign new_P3_ADD_318_U176 = ~new_P3_ADD_318_U104 | ~new_P3_ADD_318_U27;
  assign new_P3_ADD_318_U177 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_ADD_318_U24;
  assign new_P3_ADD_318_U178 = ~new_P3_ADD_318_U103 | ~new_P3_ADD_318_U25;
  assign new_P3_ADD_318_U179 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_ADD_318_U22;
  assign new_P3_ADD_318_U180 = ~new_P3_ADD_318_U102 | ~new_P3_ADD_318_U23;
  assign new_P3_ADD_318_U181 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_ADD_318_U20;
  assign new_P3_ADD_318_U182 = ~new_P3_ADD_318_U101 | ~new_P3_ADD_318_U21;
  assign new_P3_SUB_370_U6 = ~new_P3_SUB_370_U45 | ~new_P3_SUB_370_U44;
  assign new_P3_SUB_370_U7 = ~new_P3_SUB_370_U9 | ~new_P3_SUB_370_U46;
  assign new_P3_SUB_370_U8 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_SUB_370_U9 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_370_U18;
  assign new_P3_SUB_370_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_370_U11 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_370_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_370_U13 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_370_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_370_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_370_U16 = ~new_P3_SUB_370_U41 | ~new_P3_SUB_370_U40;
  assign new_P3_SUB_370_U17 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_370_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_370_U19 = ~new_P3_SUB_370_U51 | ~new_P3_SUB_370_U50;
  assign new_P3_SUB_370_U20 = ~new_P3_SUB_370_U56 | ~new_P3_SUB_370_U55;
  assign new_P3_SUB_370_U21 = ~new_P3_SUB_370_U61 | ~new_P3_SUB_370_U60;
  assign new_P3_SUB_370_U22 = ~new_P3_SUB_370_U66 | ~new_P3_SUB_370_U65;
  assign new_P3_SUB_370_U23 = ~new_P3_SUB_370_U48 | ~new_P3_SUB_370_U47;
  assign new_P3_SUB_370_U24 = ~new_P3_SUB_370_U53 | ~new_P3_SUB_370_U52;
  assign new_P3_SUB_370_U25 = ~new_P3_SUB_370_U58 | ~new_P3_SUB_370_U57;
  assign new_P3_SUB_370_U26 = ~new_P3_SUB_370_U63 | ~new_P3_SUB_370_U62;
  assign new_P3_SUB_370_U27 = ~new_P3_SUB_370_U37 | ~new_P3_SUB_370_U36;
  assign new_P3_SUB_370_U28 = ~new_P3_SUB_370_U33 | ~new_P3_SUB_370_U32;
  assign new_P3_SUB_370_U29 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_370_U30 = ~new_P3_SUB_370_U9;
  assign new_P3_SUB_370_U31 = ~new_P3_SUB_370_U30 | ~new_P3_SUB_370_U10;
  assign new_P3_SUB_370_U32 = ~new_P3_SUB_370_U31 | ~new_P3_SUB_370_U29;
  assign new_P3_SUB_370_U33 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_370_U9;
  assign new_P3_SUB_370_U34 = ~new_P3_SUB_370_U28;
  assign new_P3_SUB_370_U35 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_370_U12;
  assign new_P3_SUB_370_U36 = ~new_P3_SUB_370_U35 | ~new_P3_SUB_370_U28;
  assign new_P3_SUB_370_U37 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_370_U11;
  assign new_P3_SUB_370_U38 = ~new_P3_SUB_370_U27;
  assign new_P3_SUB_370_U39 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_370_U14;
  assign new_P3_SUB_370_U40 = ~new_P3_SUB_370_U39 | ~new_P3_SUB_370_U27;
  assign new_P3_SUB_370_U41 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_370_U13;
  assign new_P3_SUB_370_U42 = ~new_P3_SUB_370_U16;
  assign new_P3_SUB_370_U43 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_370_U17;
  assign new_P3_SUB_370_U44 = ~new_P3_SUB_370_U42 | ~new_P3_SUB_370_U43;
  assign new_P3_SUB_370_U45 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_370_U15;
  assign new_P3_SUB_370_U46 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_SUB_370_U8;
  assign new_P3_SUB_370_U47 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_370_U15;
  assign new_P3_SUB_370_U48 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_370_U17;
  assign new_P3_SUB_370_U49 = ~new_P3_SUB_370_U23;
  assign new_P3_SUB_370_U50 = ~new_P3_SUB_370_U49 | ~new_P3_SUB_370_U42;
  assign new_P3_SUB_370_U51 = ~new_P3_SUB_370_U23 | ~new_P3_SUB_370_U16;
  assign new_P3_SUB_370_U52 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_370_U14;
  assign new_P3_SUB_370_U53 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_370_U13;
  assign new_P3_SUB_370_U54 = ~new_P3_SUB_370_U24;
  assign new_P3_SUB_370_U55 = ~new_P3_SUB_370_U38 | ~new_P3_SUB_370_U54;
  assign new_P3_SUB_370_U56 = ~new_P3_SUB_370_U24 | ~new_P3_SUB_370_U27;
  assign new_P3_SUB_370_U57 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_370_U12;
  assign new_P3_SUB_370_U58 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_370_U11;
  assign new_P3_SUB_370_U59 = ~new_P3_SUB_370_U25;
  assign new_P3_SUB_370_U60 = ~new_P3_SUB_370_U34 | ~new_P3_SUB_370_U59;
  assign new_P3_SUB_370_U61 = ~new_P3_SUB_370_U25 | ~new_P3_SUB_370_U28;
  assign new_P3_SUB_370_U62 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_370_U10;
  assign new_P3_SUB_370_U63 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_370_U29;
  assign new_P3_SUB_370_U64 = ~new_P3_SUB_370_U26;
  assign new_P3_SUB_370_U65 = ~new_P3_SUB_370_U64 | ~new_P3_SUB_370_U30;
  assign new_P3_SUB_370_U66 = ~new_P3_SUB_370_U26 | ~new_P3_SUB_370_U9;
  assign new_P3_ADD_315_U4 = ~P3_PHYADDRPOINTER_REG_2_;
  assign new_P3_ADD_315_U5 = ~P3_PHYADDRPOINTER_REG_3_;
  assign new_P3_ADD_315_U6 = ~P3_PHYADDRPOINTER_REG_3_ | ~P3_PHYADDRPOINTER_REG_2_;
  assign new_P3_ADD_315_U7 = ~P3_PHYADDRPOINTER_REG_4_;
  assign new_P3_ADD_315_U8 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_ADD_315_U91;
  assign new_P3_ADD_315_U9 = ~P3_PHYADDRPOINTER_REG_5_;
  assign new_P3_ADD_315_U10 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_ADD_315_U92;
  assign new_P3_ADD_315_U11 = ~P3_PHYADDRPOINTER_REG_6_;
  assign new_P3_ADD_315_U12 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_ADD_315_U93;
  assign new_P3_ADD_315_U13 = ~P3_PHYADDRPOINTER_REG_7_;
  assign new_P3_ADD_315_U14 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_ADD_315_U94;
  assign new_P3_ADD_315_U15 = ~P3_PHYADDRPOINTER_REG_8_;
  assign new_P3_ADD_315_U16 = ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_ADD_315_U17 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_ADD_315_U95;
  assign new_P3_ADD_315_U18 = ~new_P3_ADD_315_U96 | ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_ADD_315_U19 = ~P3_PHYADDRPOINTER_REG_10_;
  assign new_P3_ADD_315_U20 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_ADD_315_U97;
  assign new_P3_ADD_315_U21 = ~P3_PHYADDRPOINTER_REG_11_;
  assign new_P3_ADD_315_U22 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_ADD_315_U98;
  assign new_P3_ADD_315_U23 = ~P3_PHYADDRPOINTER_REG_12_;
  assign new_P3_ADD_315_U24 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_ADD_315_U99;
  assign new_P3_ADD_315_U25 = ~P3_PHYADDRPOINTER_REG_13_;
  assign new_P3_ADD_315_U26 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_ADD_315_U100;
  assign new_P3_ADD_315_U27 = ~P3_PHYADDRPOINTER_REG_14_;
  assign new_P3_ADD_315_U28 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_ADD_315_U101;
  assign new_P3_ADD_315_U29 = ~P3_PHYADDRPOINTER_REG_15_;
  assign new_P3_ADD_315_U30 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_ADD_315_U102;
  assign new_P3_ADD_315_U31 = ~P3_PHYADDRPOINTER_REG_16_;
  assign new_P3_ADD_315_U32 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_ADD_315_U103;
  assign new_P3_ADD_315_U33 = ~P3_PHYADDRPOINTER_REG_17_;
  assign new_P3_ADD_315_U34 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_ADD_315_U104;
  assign new_P3_ADD_315_U35 = ~P3_PHYADDRPOINTER_REG_18_;
  assign new_P3_ADD_315_U36 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_ADD_315_U105;
  assign new_P3_ADD_315_U37 = ~P3_PHYADDRPOINTER_REG_19_;
  assign new_P3_ADD_315_U38 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_ADD_315_U106;
  assign new_P3_ADD_315_U39 = ~P3_PHYADDRPOINTER_REG_20_;
  assign new_P3_ADD_315_U40 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_ADD_315_U107;
  assign new_P3_ADD_315_U41 = ~P3_PHYADDRPOINTER_REG_21_;
  assign new_P3_ADD_315_U42 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_ADD_315_U108;
  assign new_P3_ADD_315_U43 = ~P3_PHYADDRPOINTER_REG_22_;
  assign new_P3_ADD_315_U44 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_ADD_315_U109;
  assign new_P3_ADD_315_U45 = ~P3_PHYADDRPOINTER_REG_23_;
  assign new_P3_ADD_315_U46 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_ADD_315_U110;
  assign new_P3_ADD_315_U47 = ~P3_PHYADDRPOINTER_REG_24_;
  assign new_P3_ADD_315_U48 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_ADD_315_U111;
  assign new_P3_ADD_315_U49 = ~P3_PHYADDRPOINTER_REG_25_;
  assign new_P3_ADD_315_U50 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_ADD_315_U112;
  assign new_P3_ADD_315_U51 = ~P3_PHYADDRPOINTER_REG_26_;
  assign new_P3_ADD_315_U52 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_ADD_315_U113;
  assign new_P3_ADD_315_U53 = ~P3_PHYADDRPOINTER_REG_27_;
  assign new_P3_ADD_315_U54 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_ADD_315_U114;
  assign new_P3_ADD_315_U55 = ~P3_PHYADDRPOINTER_REG_28_;
  assign new_P3_ADD_315_U56 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_ADD_315_U115;
  assign new_P3_ADD_315_U57 = ~P3_PHYADDRPOINTER_REG_29_;
  assign new_P3_ADD_315_U58 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_ADD_315_U116;
  assign new_P3_ADD_315_U59 = ~P3_PHYADDRPOINTER_REG_30_;
  assign new_P3_ADD_315_U60 = ~new_P3_ADD_315_U120 | ~new_P3_ADD_315_U119;
  assign new_P3_ADD_315_U61 = ~new_P3_ADD_315_U122 | ~new_P3_ADD_315_U121;
  assign new_P3_ADD_315_U62 = ~new_P3_ADD_315_U124 | ~new_P3_ADD_315_U123;
  assign new_P3_ADD_315_U63 = ~new_P3_ADD_315_U126 | ~new_P3_ADD_315_U125;
  assign new_P3_ADD_315_U64 = ~new_P3_ADD_315_U128 | ~new_P3_ADD_315_U127;
  assign new_P3_ADD_315_U65 = ~new_P3_ADD_315_U130 | ~new_P3_ADD_315_U129;
  assign new_P3_ADD_315_U66 = ~new_P3_ADD_315_U132 | ~new_P3_ADD_315_U131;
  assign new_P3_ADD_315_U67 = ~new_P3_ADD_315_U134 | ~new_P3_ADD_315_U133;
  assign new_P3_ADD_315_U68 = ~new_P3_ADD_315_U136 | ~new_P3_ADD_315_U135;
  assign new_P3_ADD_315_U69 = ~new_P3_ADD_315_U138 | ~new_P3_ADD_315_U137;
  assign new_P3_ADD_315_U70 = ~new_P3_ADD_315_U140 | ~new_P3_ADD_315_U139;
  assign new_P3_ADD_315_U71 = ~new_P3_ADD_315_U142 | ~new_P3_ADD_315_U141;
  assign new_P3_ADD_315_U72 = ~new_P3_ADD_315_U144 | ~new_P3_ADD_315_U143;
  assign new_P3_ADD_315_U73 = ~new_P3_ADD_315_U146 | ~new_P3_ADD_315_U145;
  assign new_P3_ADD_315_U74 = ~new_P3_ADD_315_U148 | ~new_P3_ADD_315_U147;
  assign new_P3_ADD_315_U75 = ~new_P3_ADD_315_U150 | ~new_P3_ADD_315_U149;
  assign new_P3_ADD_315_U76 = ~new_P3_ADD_315_U152 | ~new_P3_ADD_315_U151;
  assign new_P3_ADD_315_U77 = ~new_P3_ADD_315_U154 | ~new_P3_ADD_315_U153;
  assign new_P3_ADD_315_U78 = ~new_P3_ADD_315_U156 | ~new_P3_ADD_315_U155;
  assign new_P3_ADD_315_U79 = ~new_P3_ADD_315_U158 | ~new_P3_ADD_315_U157;
  assign new_P3_ADD_315_U80 = ~new_P3_ADD_315_U160 | ~new_P3_ADD_315_U159;
  assign new_P3_ADD_315_U81 = ~new_P3_ADD_315_U162 | ~new_P3_ADD_315_U161;
  assign new_P3_ADD_315_U82 = ~new_P3_ADD_315_U164 | ~new_P3_ADD_315_U163;
  assign new_P3_ADD_315_U83 = ~new_P3_ADD_315_U166 | ~new_P3_ADD_315_U165;
  assign new_P3_ADD_315_U84 = ~new_P3_ADD_315_U168 | ~new_P3_ADD_315_U167;
  assign new_P3_ADD_315_U85 = ~new_P3_ADD_315_U170 | ~new_P3_ADD_315_U169;
  assign new_P3_ADD_315_U86 = ~new_P3_ADD_315_U172 | ~new_P3_ADD_315_U171;
  assign new_P3_ADD_315_U87 = ~new_P3_ADD_315_U174 | ~new_P3_ADD_315_U173;
  assign new_P3_ADD_315_U88 = ~new_P3_ADD_315_U176 | ~new_P3_ADD_315_U175;
  assign new_P3_ADD_315_U89 = ~P3_PHYADDRPOINTER_REG_31_;
  assign new_P3_ADD_315_U90 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_ADD_315_U117;
  assign new_P3_ADD_315_U91 = ~new_P3_ADD_315_U6;
  assign new_P3_ADD_315_U92 = ~new_P3_ADD_315_U8;
  assign new_P3_ADD_315_U93 = ~new_P3_ADD_315_U10;
  assign new_P3_ADD_315_U94 = ~new_P3_ADD_315_U12;
  assign new_P3_ADD_315_U95 = ~new_P3_ADD_315_U14;
  assign new_P3_ADD_315_U96 = ~new_P3_ADD_315_U17;
  assign new_P3_ADD_315_U97 = ~new_P3_ADD_315_U18;
  assign new_P3_ADD_315_U98 = ~new_P3_ADD_315_U20;
  assign new_P3_ADD_315_U99 = ~new_P3_ADD_315_U22;
  assign new_P3_ADD_315_U100 = ~new_P3_ADD_315_U24;
  assign new_P3_ADD_315_U101 = ~new_P3_ADD_315_U26;
  assign new_P3_ADD_315_U102 = ~new_P3_ADD_315_U28;
  assign new_P3_ADD_315_U103 = ~new_P3_ADD_315_U30;
  assign new_P3_ADD_315_U104 = ~new_P3_ADD_315_U32;
  assign new_P3_ADD_315_U105 = ~new_P3_ADD_315_U34;
  assign new_P3_ADD_315_U106 = ~new_P3_ADD_315_U36;
  assign new_P3_ADD_315_U107 = ~new_P3_ADD_315_U38;
  assign new_P3_ADD_315_U108 = ~new_P3_ADD_315_U40;
  assign new_P3_ADD_315_U109 = ~new_P3_ADD_315_U42;
  assign new_P3_ADD_315_U110 = ~new_P3_ADD_315_U44;
  assign new_P3_ADD_315_U111 = ~new_P3_ADD_315_U46;
  assign new_P3_ADD_315_U112 = ~new_P3_ADD_315_U48;
  assign new_P3_ADD_315_U113 = ~new_P3_ADD_315_U50;
  assign new_P3_ADD_315_U114 = ~new_P3_ADD_315_U52;
  assign new_P3_ADD_315_U115 = ~new_P3_ADD_315_U54;
  assign new_P3_ADD_315_U116 = ~new_P3_ADD_315_U56;
  assign new_P3_ADD_315_U117 = ~new_P3_ADD_315_U58;
  assign new_P3_ADD_315_U118 = ~new_P3_ADD_315_U90;
  assign new_P3_ADD_315_U119 = ~P3_PHYADDRPOINTER_REG_9_ | ~new_P3_ADD_315_U17;
  assign new_P3_ADD_315_U120 = ~new_P3_ADD_315_U96 | ~new_P3_ADD_315_U16;
  assign new_P3_ADD_315_U121 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_ADD_315_U14;
  assign new_P3_ADD_315_U122 = ~new_P3_ADD_315_U95 | ~new_P3_ADD_315_U15;
  assign new_P3_ADD_315_U123 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_ADD_315_U12;
  assign new_P3_ADD_315_U124 = ~new_P3_ADD_315_U94 | ~new_P3_ADD_315_U13;
  assign new_P3_ADD_315_U125 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_ADD_315_U10;
  assign new_P3_ADD_315_U126 = ~new_P3_ADD_315_U93 | ~new_P3_ADD_315_U11;
  assign new_P3_ADD_315_U127 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_ADD_315_U8;
  assign new_P3_ADD_315_U128 = ~new_P3_ADD_315_U92 | ~new_P3_ADD_315_U9;
  assign new_P3_ADD_315_U129 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_ADD_315_U6;
  assign new_P3_ADD_315_U130 = ~new_P3_ADD_315_U91 | ~new_P3_ADD_315_U7;
  assign new_P3_ADD_315_U131 = ~P3_PHYADDRPOINTER_REG_3_ | ~new_P3_ADD_315_U4;
  assign new_P3_ADD_315_U132 = ~P3_PHYADDRPOINTER_REG_2_ | ~new_P3_ADD_315_U5;
  assign new_P3_ADD_315_U133 = ~P3_PHYADDRPOINTER_REG_31_ | ~new_P3_ADD_315_U90;
  assign new_P3_ADD_315_U134 = ~new_P3_ADD_315_U118 | ~new_P3_ADD_315_U89;
  assign new_P3_ADD_315_U135 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_ADD_315_U58;
  assign new_P3_ADD_315_U136 = ~new_P3_ADD_315_U117 | ~new_P3_ADD_315_U59;
  assign new_P3_ADD_315_U137 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_ADD_315_U56;
  assign new_P3_ADD_315_U138 = ~new_P3_ADD_315_U116 | ~new_P3_ADD_315_U57;
  assign new_P3_ADD_315_U139 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_ADD_315_U54;
  assign new_P3_ADD_315_U140 = ~new_P3_ADD_315_U115 | ~new_P3_ADD_315_U55;
  assign new_P3_ADD_315_U141 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_ADD_315_U52;
  assign new_P3_ADD_315_U142 = ~new_P3_ADD_315_U114 | ~new_P3_ADD_315_U53;
  assign new_P3_ADD_315_U143 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_ADD_315_U50;
  assign new_P3_ADD_315_U144 = ~new_P3_ADD_315_U113 | ~new_P3_ADD_315_U51;
  assign new_P3_ADD_315_U145 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_ADD_315_U48;
  assign new_P3_ADD_315_U146 = ~new_P3_ADD_315_U112 | ~new_P3_ADD_315_U49;
  assign new_P3_ADD_315_U147 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_ADD_315_U46;
  assign new_P3_ADD_315_U148 = ~new_P3_ADD_315_U111 | ~new_P3_ADD_315_U47;
  assign new_P3_ADD_315_U149 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_ADD_315_U44;
  assign new_P3_ADD_315_U150 = ~new_P3_ADD_315_U110 | ~new_P3_ADD_315_U45;
  assign new_P3_ADD_315_U151 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_ADD_315_U42;
  assign new_P3_ADD_315_U152 = ~new_P3_ADD_315_U109 | ~new_P3_ADD_315_U43;
  assign new_P3_ADD_315_U153 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_ADD_315_U40;
  assign new_P3_ADD_315_U154 = ~new_P3_ADD_315_U108 | ~new_P3_ADD_315_U41;
  assign new_P3_ADD_315_U155 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_ADD_315_U38;
  assign new_P3_ADD_315_U156 = ~new_P3_ADD_315_U107 | ~new_P3_ADD_315_U39;
  assign new_P3_ADD_315_U157 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_ADD_315_U36;
  assign new_P3_ADD_315_U158 = ~new_P3_ADD_315_U106 | ~new_P3_ADD_315_U37;
  assign new_P3_ADD_315_U159 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_ADD_315_U34;
  assign new_P3_ADD_315_U160 = ~new_P3_ADD_315_U105 | ~new_P3_ADD_315_U35;
  assign new_P3_ADD_315_U161 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_ADD_315_U32;
  assign new_P3_ADD_315_U162 = ~new_P3_ADD_315_U104 | ~new_P3_ADD_315_U33;
  assign new_P3_ADD_315_U163 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_ADD_315_U30;
  assign new_P3_ADD_315_U164 = ~new_P3_ADD_315_U103 | ~new_P3_ADD_315_U31;
  assign new_P3_ADD_315_U165 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_ADD_315_U28;
  assign new_P3_ADD_315_U166 = ~new_P3_ADD_315_U102 | ~new_P3_ADD_315_U29;
  assign new_P3_ADD_315_U167 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_ADD_315_U26;
  assign new_P3_ADD_315_U168 = ~new_P3_ADD_315_U101 | ~new_P3_ADD_315_U27;
  assign new_P3_ADD_315_U169 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_ADD_315_U24;
  assign new_P3_ADD_315_U170 = ~new_P3_ADD_315_U100 | ~new_P3_ADD_315_U25;
  assign new_P3_ADD_315_U171 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_ADD_315_U22;
  assign new_P3_ADD_315_U172 = ~new_P3_ADD_315_U99 | ~new_P3_ADD_315_U23;
  assign new_P3_ADD_315_U173 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_ADD_315_U20;
  assign new_P3_ADD_315_U174 = ~new_P3_ADD_315_U98 | ~new_P3_ADD_315_U21;
  assign new_P3_ADD_315_U175 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_ADD_315_U18;
  assign new_P3_ADD_315_U176 = ~new_P3_ADD_315_U97 | ~new_P3_ADD_315_U19;
  assign new_P3_GTE_355_U6 = ~new_P3_SUB_355_U6 & ~new_P3_GTE_355_U8;
  assign new_P3_GTE_355_U7 = new_P3_SUB_355_U7 & new_P3_SUB_355_U22;
  assign new_P3_GTE_355_U8 = ~new_P3_SUB_355_U21 & ~new_P3_GTE_355_U7 & ~new_P3_SUB_355_U19 & ~new_P3_SUB_355_U20;
  assign new_P3_ADD_360_1242_U4 = new_P3_ADD_360_1242_U186 & new_P3_ADD_360_1242_U45;
  assign new_P3_ADD_360_1242_U5 = new_P3_ADD_360_1242_U184 & new_P3_ADD_360_1242_U46;
  assign new_P3_ADD_360_1242_U6 = new_P3_ADD_360_1242_U182 & new_P3_ADD_360_1242_U76;
  assign new_P3_ADD_360_1242_U7 = new_P3_ADD_360_1242_U181 & new_P3_ADD_360_1242_U50;
  assign new_P3_ADD_360_1242_U8 = new_P3_ADD_360_1242_U179 & new_P3_ADD_360_1242_U53;
  assign new_P3_ADD_360_1242_U9 = new_P3_ADD_360_1242_U177 & new_P3_ADD_360_1242_U56;
  assign new_P3_ADD_360_1242_U10 = new_P3_ADD_360_1242_U175 & new_P3_ADD_360_1242_U58;
  assign new_P3_ADD_360_1242_U11 = new_P3_ADD_360_1242_U174 & new_P3_ADD_360_1242_U60;
  assign new_P3_ADD_360_1242_U12 = new_P3_ADD_360_1242_U173 & new_P3_ADD_360_1242_U63;
  assign new_P3_ADD_360_1242_U13 = new_P3_ADD_360_1242_U171 & new_P3_ADD_360_1242_U66;
  assign new_P3_ADD_360_1242_U14 = new_P3_ADD_360_1242_U169 & new_P3_ADD_360_1242_U68;
  assign new_P3_ADD_360_1242_U15 = new_P3_ADD_360_1242_U168 & new_P3_ADD_360_1242_U71;
  assign new_P3_ADD_360_1242_U16 = new_P3_ADD_360_1242_U166 & new_P3_ADD_360_1242_U73;
  assign new_P3_ADD_360_1242_U17 = new_P3_ADD_360_1242_U153 & new_P3_ADD_360_1242_U152;
  assign new_P3_ADD_360_1242_U18 = new_P3_ADD_360_1242_U151 & new_P3_ADD_360_1242_U149;
  assign new_P3_ADD_360_1242_U19 = ~new_P3_ADD_360_1242_U192 | ~new_P3_ADD_360_1242_U248 | ~new_P3_ADD_360_1242_U247;
  assign new_P3_ADD_360_1242_U20 = ~new_P3_ADD_360_U19;
  assign new_P3_ADD_360_1242_U21 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_360_1242_U22 = ~new_P3_ADD_360_U20;
  assign new_P3_ADD_360_1242_U23 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_360_1242_U24 = ~new_P3_U2621;
  assign new_P3_ADD_360_1242_U25 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_360_1242_U26 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_360_1242_U27 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_U2621;
  assign new_P3_ADD_360_1242_U28 = ~new_P3_ADD_360_U4;
  assign new_P3_ADD_360_1242_U29 = ~new_P3_ADD_360_U21;
  assign new_P3_ADD_360_1242_U30 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_360_1242_U31 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_360_1242_U32 = ~new_P3_ADD_360_U18;
  assign new_P3_ADD_360_1242_U33 = ~new_P3_ADD_360_U17;
  assign new_P3_ADD_360_1242_U34 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_360_1242_U35 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_360_1242_U36 = ~new_P3_ADD_360_U16;
  assign new_P3_ADD_360_1242_U37 = ~new_P3_ADD_360_U5;
  assign new_P3_ADD_360_1242_U38 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_360_1242_U39 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_360_1242_U40 = ~new_P3_ADD_360_1242_U131 | ~new_P3_ADD_360_1242_U130;
  assign new_P3_ADD_360_1242_U41 = ~new_P3_ADD_360_1242_U40 | ~new_P3_ADD_360_1242_U133;
  assign new_P3_ADD_360_1242_U42 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_360_1242_U43 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_360_1242_U44 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_360_1242_U45 = ~new_P3_ADD_360_1242_U97 | ~new_P3_ADD_360_1242_U105;
  assign new_P3_ADD_360_1242_U46 = ~new_P3_ADD_360_1242_U98 | ~new_P3_ADD_360_1242_U119;
  assign new_P3_ADD_360_1242_U47 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_360_1242_U48 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_360_1242_U49 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_360_1242_U50 = ~new_P3_ADD_360_1242_U154 | ~new_P3_ADD_360_1242_U99;
  assign new_P3_ADD_360_1242_U51 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_360_1242_U52 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_360_1242_U53 = ~new_P3_ADD_360_1242_U100 | ~new_P3_ADD_360_1242_U156;
  assign new_P3_ADD_360_1242_U54 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_360_1242_U55 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_360_1242_U56 = ~new_P3_ADD_360_1242_U101 | ~new_P3_ADD_360_1242_U157;
  assign new_P3_ADD_360_1242_U57 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_360_1242_U58 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_360_1242_U158;
  assign new_P3_ADD_360_1242_U59 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_360_1242_U60 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_360_1242_U159;
  assign new_P3_ADD_360_1242_U61 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_360_1242_U62 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_360_1242_U63 = ~new_P3_ADD_360_1242_U102 | ~new_P3_ADD_360_1242_U160;
  assign new_P3_ADD_360_1242_U64 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_360_1242_U65 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_360_1242_U66 = ~new_P3_ADD_360_1242_U103 | ~new_P3_ADD_360_1242_U161;
  assign new_P3_ADD_360_1242_U67 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_360_1242_U68 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_360_1242_U162;
  assign new_P3_ADD_360_1242_U69 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_360_1242_U70 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_360_1242_U71 = ~new_P3_ADD_360_1242_U104 | ~new_P3_ADD_360_1242_U163;
  assign new_P3_ADD_360_1242_U72 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_360_1242_U73 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_360_1242_U164;
  assign new_P3_ADD_360_1242_U74 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_360_1242_U75 = ~new_P3_ADD_360_U4 | ~new_P3_ADD_360_1242_U124;
  assign new_P3_ADD_360_1242_U76 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_360_1242_U154;
  assign new_P3_ADD_360_1242_U77 = ~new_P3_ADD_360_1242_U230 | ~new_P3_ADD_360_1242_U229;
  assign new_P3_ADD_360_1242_U78 = ~new_P3_ADD_360_1242_U239 | ~new_P3_ADD_360_1242_U238;
  assign new_P3_ADD_360_1242_U79 = ~new_P3_ADD_360_1242_U241 | ~new_P3_ADD_360_1242_U240;
  assign new_P3_ADD_360_1242_U80 = ~new_P3_ADD_360_1242_U243 | ~new_P3_ADD_360_1242_U242;
  assign new_P3_ADD_360_1242_U81 = ~new_P3_ADD_360_1242_U250 | ~new_P3_ADD_360_1242_U249;
  assign new_P3_ADD_360_1242_U82 = ~new_P3_ADD_360_1242_U252 | ~new_P3_ADD_360_1242_U251;
  assign new_P3_ADD_360_1242_U83 = ~new_P3_ADD_360_1242_U254 | ~new_P3_ADD_360_1242_U253;
  assign new_P3_ADD_360_1242_U84 = ~new_P3_ADD_360_1242_U256 | ~new_P3_ADD_360_1242_U255;
  assign new_P3_ADD_360_1242_U85 = ~new_P3_ADD_360_1242_U258 | ~new_P3_ADD_360_1242_U257;
  assign new_P3_ADD_360_1242_U86 = ~new_P3_ADD_360_1242_U201 | ~new_P3_ADD_360_1242_U200;
  assign new_P3_ADD_360_1242_U87 = ~new_P3_ADD_360_1242_U208 | ~new_P3_ADD_360_1242_U207;
  assign new_P3_ADD_360_1242_U88 = ~new_P3_ADD_360_1242_U215 | ~new_P3_ADD_360_1242_U214;
  assign new_P3_ADD_360_1242_U89 = ~new_P3_ADD_360_1242_U222 | ~new_P3_ADD_360_1242_U221;
  assign new_P3_ADD_360_1242_U90 = ~new_P3_ADD_360_1242_U228 | ~new_P3_ADD_360_1242_U227;
  assign new_P3_ADD_360_1242_U91 = ~new_P3_ADD_360_1242_U237 | ~new_P3_ADD_360_1242_U236;
  assign new_P3_ADD_360_1242_U92 = new_P3_ADD_360_U20 & P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_360_1242_U93 = new_P3_ADD_360_1242_U133 & new_P3_ADD_360_1242_U123;
  assign new_P3_ADD_360_1242_U94 = new_P3_ADD_360_1242_U190 & new_P3_ADD_360_1242_U125;
  assign new_P3_ADD_360_1242_U95 = new_P3_ADD_360_1242_U135 & new_P3_ADD_360_1242_U224 & new_P3_ADD_360_1242_U223;
  assign new_P3_ADD_360_1242_U96 = new_P3_ADD_360_1242_U125 & new_P3_ADD_360_1242_U123;
  assign new_P3_ADD_360_1242_U97 = P3_INSTADDRPOINTER_REG_9_ & P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_360_1242_U98 = P3_INSTADDRPOINTER_REG_12_ & P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_360_1242_U99 = P3_INSTADDRPOINTER_REG_13_ & P3_INSTADDRPOINTER_REG_14_ & P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_360_1242_U100 = P3_INSTADDRPOINTER_REG_17_ & P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_360_1242_U101 = P3_INSTADDRPOINTER_REG_18_ & P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_360_1242_U102 = P3_INSTADDRPOINTER_REG_23_ & P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_360_1242_U103 = P3_INSTADDRPOINTER_REG_25_ & P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_360_1242_U104 = P3_INSTADDRPOINTER_REG_28_ & P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_360_1242_U105 = ~new_P3_ADD_360_1242_U147 | ~new_P3_ADD_360_1242_U146;
  assign new_P3_ADD_360_1242_U106 = new_P3_ADD_360_1242_U194 & new_P3_ADD_360_1242_U193;
  assign new_P3_ADD_360_1242_U107 = new_P3_ADD_360_1242_U196 & new_P3_ADD_360_1242_U195;
  assign new_P3_ADD_360_1242_U108 = ~new_P3_ADD_360_1242_U189 | ~new_P3_ADD_360_1242_U143 | ~new_P3_ADD_360_1242_U120;
  assign new_P3_ADD_360_1242_U109 = new_P3_ADD_360_1242_U203 & new_P3_ADD_360_1242_U202;
  assign new_P3_ADD_360_1242_U110 = ~new_P3_ADD_360_1242_U141 | ~new_P3_ADD_360_1242_U140;
  assign new_P3_ADD_360_1242_U111 = new_P3_ADD_360_1242_U210 & new_P3_ADD_360_1242_U209;
  assign new_P3_ADD_360_1242_U112 = ~new_P3_ADD_360_1242_U188 | ~new_P3_ADD_360_1242_U137 | ~new_P3_ADD_360_1242_U121;
  assign new_P3_ADD_360_1242_U113 = new_P3_ADD_360_1242_U217 & new_P3_ADD_360_1242_U216;
  assign new_P3_ADD_360_1242_U114 = ~new_P3_ADD_360_1242_U94 | ~new_P3_ADD_360_1242_U191;
  assign new_P3_ADD_360_1242_U115 = new_P3_ADD_360_1242_U226 & new_P3_ADD_360_1242_U225;
  assign new_P3_ADD_360_1242_U116 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_360_1242_U117 = new_P3_ADD_360_1242_U232 & new_P3_ADD_360_1242_U231;
  assign new_P3_ADD_360_1242_U118 = ~new_P3_ADD_360_1242_U75 | ~new_P3_ADD_360_1242_U127;
  assign new_P3_ADD_360_1242_U119 = ~new_P3_ADD_360_1242_U45;
  assign new_P3_ADD_360_1242_U120 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_360_1242_U110;
  assign new_P3_ADD_360_1242_U121 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_360_1242_U114;
  assign new_P3_ADD_360_1242_U122 = ~new_P3_ADD_360_1242_U75;
  assign new_P3_ADD_360_1242_U123 = P3_INSTADDRPOINTER_REG_4_ | new_P3_ADD_360_U19;
  assign new_P3_ADD_360_1242_U124 = ~new_P3_ADD_360_1242_U27;
  assign new_P3_ADD_360_1242_U125 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_360_U19;
  assign new_P3_ADD_360_1242_U126 = ~new_P3_ADD_360_1242_U28 | ~new_P3_ADD_360_1242_U27;
  assign new_P3_ADD_360_1242_U127 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_360_1242_U126;
  assign new_P3_ADD_360_1242_U128 = ~new_P3_ADD_360_1242_U118;
  assign new_P3_ADD_360_1242_U129 = new_P3_ADD_360_U21 | P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_360_1242_U130 = ~new_P3_ADD_360_1242_U129 | ~new_P3_ADD_360_1242_U118;
  assign new_P3_ADD_360_1242_U131 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_360_U21;
  assign new_P3_ADD_360_1242_U132 = ~new_P3_ADD_360_1242_U40;
  assign new_P3_ADD_360_1242_U133 = P3_INSTADDRPOINTER_REG_3_ | new_P3_ADD_360_U20;
  assign new_P3_ADD_360_1242_U134 = ~new_P3_ADD_360_1242_U41;
  assign new_P3_ADD_360_1242_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_360_U20;
  assign new_P3_ADD_360_1242_U136 = ~new_P3_ADD_360_1242_U114;
  assign new_P3_ADD_360_1242_U137 = ~new_P3_ADD_360_U18 | ~new_P3_ADD_360_1242_U114;
  assign new_P3_ADD_360_1242_U138 = ~new_P3_ADD_360_1242_U112;
  assign new_P3_ADD_360_1242_U139 = new_P3_ADD_360_U17 | P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_360_1242_U140 = ~new_P3_ADD_360_1242_U139 | ~new_P3_ADD_360_1242_U112;
  assign new_P3_ADD_360_1242_U141 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_360_U17;
  assign new_P3_ADD_360_1242_U142 = ~new_P3_ADD_360_1242_U110;
  assign new_P3_ADD_360_1242_U143 = ~new_P3_ADD_360_U16 | ~new_P3_ADD_360_1242_U110;
  assign new_P3_ADD_360_1242_U144 = ~new_P3_ADD_360_1242_U108;
  assign new_P3_ADD_360_1242_U145 = new_P3_ADD_360_U5 | P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_360_1242_U146 = ~new_P3_ADD_360_1242_U145 | ~new_P3_ADD_360_1242_U108;
  assign new_P3_ADD_360_1242_U147 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_360_U5;
  assign new_P3_ADD_360_1242_U148 = ~new_P3_ADD_360_1242_U105;
  assign new_P3_ADD_360_1242_U149 = ~new_P3_ADD_360_1242_U95 | ~new_P3_ADD_360_1242_U41;
  assign new_P3_ADD_360_1242_U150 = ~new_P3_ADD_360_1242_U135 | ~new_P3_ADD_360_1242_U41;
  assign new_P3_ADD_360_1242_U151 = ~new_P3_ADD_360_1242_U96 | ~new_P3_ADD_360_1242_U150;
  assign new_P3_ADD_360_1242_U152 = ~new_P3_ADD_360_1242_U115 | ~new_P3_ADD_360_1242_U132;
  assign new_P3_ADD_360_1242_U153 = ~new_P3_ADD_360_1242_U134 | ~new_P3_ADD_360_1242_U135;
  assign new_P3_ADD_360_1242_U154 = ~new_P3_ADD_360_1242_U46;
  assign new_P3_ADD_360_1242_U155 = ~new_P3_ADD_360_1242_U76;
  assign new_P3_ADD_360_1242_U156 = ~new_P3_ADD_360_1242_U50;
  assign new_P3_ADD_360_1242_U157 = ~new_P3_ADD_360_1242_U53;
  assign new_P3_ADD_360_1242_U158 = ~new_P3_ADD_360_1242_U56;
  assign new_P3_ADD_360_1242_U159 = ~new_P3_ADD_360_1242_U58;
  assign new_P3_ADD_360_1242_U160 = ~new_P3_ADD_360_1242_U60;
  assign new_P3_ADD_360_1242_U161 = ~new_P3_ADD_360_1242_U63;
  assign new_P3_ADD_360_1242_U162 = ~new_P3_ADD_360_1242_U66;
  assign new_P3_ADD_360_1242_U163 = ~new_P3_ADD_360_1242_U68;
  assign new_P3_ADD_360_1242_U164 = ~new_P3_ADD_360_1242_U71;
  assign new_P3_ADD_360_1242_U165 = ~new_P3_ADD_360_1242_U73;
  assign new_P3_ADD_360_1242_U166 = ~new_P3_ADD_360_1242_U72 | ~new_P3_ADD_360_1242_U71;
  assign new_P3_ADD_360_1242_U167 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_360_1242_U163;
  assign new_P3_ADD_360_1242_U168 = ~new_P3_ADD_360_1242_U69 | ~new_P3_ADD_360_1242_U167;
  assign new_P3_ADD_360_1242_U169 = ~new_P3_ADD_360_1242_U67 | ~new_P3_ADD_360_1242_U66;
  assign new_P3_ADD_360_1242_U170 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_360_1242_U161;
  assign new_P3_ADD_360_1242_U171 = ~new_P3_ADD_360_1242_U64 | ~new_P3_ADD_360_1242_U170;
  assign new_P3_ADD_360_1242_U172 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_360_1242_U160;
  assign new_P3_ADD_360_1242_U173 = ~new_P3_ADD_360_1242_U61 | ~new_P3_ADD_360_1242_U172;
  assign new_P3_ADD_360_1242_U174 = ~new_P3_ADD_360_1242_U59 | ~new_P3_ADD_360_1242_U58;
  assign new_P3_ADD_360_1242_U175 = ~new_P3_ADD_360_1242_U57 | ~new_P3_ADD_360_1242_U56;
  assign new_P3_ADD_360_1242_U176 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_360_1242_U157;
  assign new_P3_ADD_360_1242_U177 = ~new_P3_ADD_360_1242_U55 | ~new_P3_ADD_360_1242_U176;
  assign new_P3_ADD_360_1242_U178 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_360_1242_U156;
  assign new_P3_ADD_360_1242_U179 = ~new_P3_ADD_360_1242_U51 | ~new_P3_ADD_360_1242_U178;
  assign new_P3_ADD_360_1242_U180 = ~new_P3_ADD_360_1242_U155 | ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_360_1242_U181 = ~new_P3_ADD_360_1242_U48 | ~new_P3_ADD_360_1242_U180;
  assign new_P3_ADD_360_1242_U182 = ~new_P3_ADD_360_1242_U47 | ~new_P3_ADD_360_1242_U46;
  assign new_P3_ADD_360_1242_U183 = ~new_P3_ADD_360_1242_U119 | ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_360_1242_U184 = ~new_P3_ADD_360_1242_U44 | ~new_P3_ADD_360_1242_U183;
  assign new_P3_ADD_360_1242_U185 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_360_1242_U105;
  assign new_P3_ADD_360_1242_U186 = ~new_P3_ADD_360_1242_U42 | ~new_P3_ADD_360_1242_U185;
  assign new_P3_ADD_360_1242_U187 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_360_1242_U165;
  assign new_P3_ADD_360_1242_U188 = ~new_P3_ADD_360_U18 | ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_360_1242_U189 = ~new_P3_ADD_360_U16 | ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_360_1242_U190 = ~new_P3_ADD_360_1242_U92 | ~new_P3_ADD_360_1242_U123;
  assign new_P3_ADD_360_1242_U191 = ~new_P3_ADD_360_1242_U93 | ~new_P3_ADD_360_1242_U40;
  assign new_P3_ADD_360_1242_U192 = ~new_P3_ADD_360_1242_U122 | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_360_1242_U193 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_360_1242_U105;
  assign new_P3_ADD_360_1242_U194 = ~new_P3_ADD_360_1242_U148 | ~new_P3_ADD_360_1242_U39;
  assign new_P3_ADD_360_1242_U195 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_360_1242_U37;
  assign new_P3_ADD_360_1242_U196 = ~new_P3_ADD_360_U5 | ~new_P3_ADD_360_1242_U38;
  assign new_P3_ADD_360_1242_U197 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_360_1242_U37;
  assign new_P3_ADD_360_1242_U198 = ~new_P3_ADD_360_U5 | ~new_P3_ADD_360_1242_U38;
  assign new_P3_ADD_360_1242_U199 = ~new_P3_ADD_360_1242_U198 | ~new_P3_ADD_360_1242_U197;
  assign new_P3_ADD_360_1242_U200 = ~new_P3_ADD_360_1242_U107 | ~new_P3_ADD_360_1242_U108;
  assign new_P3_ADD_360_1242_U201 = ~new_P3_ADD_360_1242_U144 | ~new_P3_ADD_360_1242_U199;
  assign new_P3_ADD_360_1242_U202 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_360_1242_U36;
  assign new_P3_ADD_360_1242_U203 = ~new_P3_ADD_360_U16 | ~new_P3_ADD_360_1242_U35;
  assign new_P3_ADD_360_1242_U204 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_360_1242_U36;
  assign new_P3_ADD_360_1242_U205 = ~new_P3_ADD_360_U16 | ~new_P3_ADD_360_1242_U35;
  assign new_P3_ADD_360_1242_U206 = ~new_P3_ADD_360_1242_U205 | ~new_P3_ADD_360_1242_U204;
  assign new_P3_ADD_360_1242_U207 = ~new_P3_ADD_360_1242_U109 | ~new_P3_ADD_360_1242_U110;
  assign new_P3_ADD_360_1242_U208 = ~new_P3_ADD_360_1242_U142 | ~new_P3_ADD_360_1242_U206;
  assign new_P3_ADD_360_1242_U209 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_360_1242_U33;
  assign new_P3_ADD_360_1242_U210 = ~new_P3_ADD_360_U17 | ~new_P3_ADD_360_1242_U34;
  assign new_P3_ADD_360_1242_U211 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_360_1242_U33;
  assign new_P3_ADD_360_1242_U212 = ~new_P3_ADD_360_U17 | ~new_P3_ADD_360_1242_U34;
  assign new_P3_ADD_360_1242_U213 = ~new_P3_ADD_360_1242_U212 | ~new_P3_ADD_360_1242_U211;
  assign new_P3_ADD_360_1242_U214 = ~new_P3_ADD_360_1242_U111 | ~new_P3_ADD_360_1242_U112;
  assign new_P3_ADD_360_1242_U215 = ~new_P3_ADD_360_1242_U138 | ~new_P3_ADD_360_1242_U213;
  assign new_P3_ADD_360_1242_U216 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_360_1242_U32;
  assign new_P3_ADD_360_1242_U217 = ~new_P3_ADD_360_U18 | ~new_P3_ADD_360_1242_U31;
  assign new_P3_ADD_360_1242_U218 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_360_1242_U32;
  assign new_P3_ADD_360_1242_U219 = ~new_P3_ADD_360_U18 | ~new_P3_ADD_360_1242_U31;
  assign new_P3_ADD_360_1242_U220 = ~new_P3_ADD_360_1242_U219 | ~new_P3_ADD_360_1242_U218;
  assign new_P3_ADD_360_1242_U221 = ~new_P3_ADD_360_1242_U113 | ~new_P3_ADD_360_1242_U114;
  assign new_P3_ADD_360_1242_U222 = ~new_P3_ADD_360_1242_U136 | ~new_P3_ADD_360_1242_U220;
  assign new_P3_ADD_360_1242_U223 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_360_1242_U20;
  assign new_P3_ADD_360_1242_U224 = ~new_P3_ADD_360_U19 | ~new_P3_ADD_360_1242_U21;
  assign new_P3_ADD_360_1242_U225 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_360_1242_U22;
  assign new_P3_ADD_360_1242_U226 = ~new_P3_ADD_360_U20 | ~new_P3_ADD_360_1242_U23;
  assign new_P3_ADD_360_1242_U227 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_360_1242_U187;
  assign new_P3_ADD_360_1242_U228 = ~new_P3_ADD_360_1242_U116 | ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_360_1242_U165;
  assign new_P3_ADD_360_1242_U229 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_360_1242_U73;
  assign new_P3_ADD_360_1242_U230 = ~new_P3_ADD_360_1242_U165 | ~new_P3_ADD_360_1242_U74;
  assign new_P3_ADD_360_1242_U231 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_360_1242_U29;
  assign new_P3_ADD_360_1242_U232 = ~new_P3_ADD_360_U21 | ~new_P3_ADD_360_1242_U30;
  assign new_P3_ADD_360_1242_U233 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_360_1242_U29;
  assign new_P3_ADD_360_1242_U234 = ~new_P3_ADD_360_U21 | ~new_P3_ADD_360_1242_U30;
  assign new_P3_ADD_360_1242_U235 = ~new_P3_ADD_360_1242_U234 | ~new_P3_ADD_360_1242_U233;
  assign new_P3_ADD_360_1242_U236 = ~new_P3_ADD_360_1242_U117 | ~new_P3_ADD_360_1242_U118;
  assign new_P3_ADD_360_1242_U237 = ~new_P3_ADD_360_1242_U128 | ~new_P3_ADD_360_1242_U235;
  assign new_P3_ADD_360_1242_U238 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_360_1242_U68;
  assign new_P3_ADD_360_1242_U239 = ~new_P3_ADD_360_1242_U163 | ~new_P3_ADD_360_1242_U70;
  assign new_P3_ADD_360_1242_U240 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_360_1242_U63;
  assign new_P3_ADD_360_1242_U241 = ~new_P3_ADD_360_1242_U161 | ~new_P3_ADD_360_1242_U65;
  assign new_P3_ADD_360_1242_U242 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_360_1242_U60;
  assign new_P3_ADD_360_1242_U243 = ~new_P3_ADD_360_1242_U160 | ~new_P3_ADD_360_1242_U62;
  assign new_P3_ADD_360_1242_U244 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_360_1242_U27;
  assign new_P3_ADD_360_1242_U245 = ~new_P3_ADD_360_1242_U124 | ~new_P3_ADD_360_1242_U26;
  assign new_P3_ADD_360_1242_U246 = ~new_P3_ADD_360_1242_U245 | ~new_P3_ADD_360_1242_U244;
  assign new_P3_ADD_360_1242_U247 = ~new_P3_ADD_360_U4 | ~new_P3_ADD_360_1242_U27 | ~new_P3_ADD_360_1242_U26;
  assign new_P3_ADD_360_1242_U248 = ~new_P3_ADD_360_1242_U246 | ~new_P3_ADD_360_1242_U28;
  assign new_P3_ADD_360_1242_U249 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_360_1242_U53;
  assign new_P3_ADD_360_1242_U250 = ~new_P3_ADD_360_1242_U157 | ~new_P3_ADD_360_1242_U54;
  assign new_P3_ADD_360_1242_U251 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_360_1242_U50;
  assign new_P3_ADD_360_1242_U252 = ~new_P3_ADD_360_1242_U156 | ~new_P3_ADD_360_1242_U52;
  assign new_P3_ADD_360_1242_U253 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_360_1242_U76;
  assign new_P3_ADD_360_1242_U254 = ~new_P3_ADD_360_1242_U155 | ~new_P3_ADD_360_1242_U49;
  assign new_P3_ADD_360_1242_U255 = ~new_P3_ADD_360_1242_U119 | ~new_P3_ADD_360_1242_U43;
  assign new_P3_ADD_360_1242_U256 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_360_1242_U45;
  assign new_P3_ADD_360_1242_U257 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_360_1242_U24;
  assign new_P3_ADD_360_1242_U258 = ~new_P3_U2621 | ~new_P3_ADD_360_1242_U25;
  assign new_P3_LT_563_1260_U6 = new_P3_LT_563_1260_U7 | new_P3_U3304;
  assign new_P3_LT_563_1260_U7 = ~new_P3_SUB_563_U7 & ~new_P3_SUB_563_U6;
  assign new_P3_SUB_589_U6 = ~new_P3_U3301;
  assign new_P3_SUB_589_U7 = ~new_P3_U3302;
  assign new_P3_SUB_589_U8 = ~new_P3_U2632;
  assign new_P3_SUB_589_U9 = ~new_P3_U3300;
  assign new_P3_ADD_467_U4 = ~P3_REIP_REG_1_;
  assign new_P3_ADD_467_U5 = ~P3_REIP_REG_2_;
  assign new_P3_ADD_467_U6 = ~P3_REIP_REG_2_ | ~P3_REIP_REG_1_;
  assign new_P3_ADD_467_U7 = ~P3_REIP_REG_3_;
  assign new_P3_ADD_467_U8 = ~P3_REIP_REG_3_ | ~new_P3_ADD_467_U94;
  assign new_P3_ADD_467_U9 = ~P3_REIP_REG_4_;
  assign new_P3_ADD_467_U10 = ~P3_REIP_REG_4_ | ~new_P3_ADD_467_U95;
  assign new_P3_ADD_467_U11 = ~P3_REIP_REG_5_;
  assign new_P3_ADD_467_U12 = ~P3_REIP_REG_5_ | ~new_P3_ADD_467_U96;
  assign new_P3_ADD_467_U13 = ~P3_REIP_REG_6_;
  assign new_P3_ADD_467_U14 = ~P3_REIP_REG_6_ | ~new_P3_ADD_467_U97;
  assign new_P3_ADD_467_U15 = ~P3_REIP_REG_7_;
  assign new_P3_ADD_467_U16 = ~P3_REIP_REG_7_ | ~new_P3_ADD_467_U98;
  assign new_P3_ADD_467_U17 = ~P3_REIP_REG_8_;
  assign new_P3_ADD_467_U18 = ~P3_REIP_REG_9_;
  assign new_P3_ADD_467_U19 = ~P3_REIP_REG_8_ | ~new_P3_ADD_467_U99;
  assign new_P3_ADD_467_U20 = ~new_P3_ADD_467_U100 | ~P3_REIP_REG_9_;
  assign new_P3_ADD_467_U21 = ~P3_REIP_REG_10_;
  assign new_P3_ADD_467_U22 = ~P3_REIP_REG_10_ | ~new_P3_ADD_467_U101;
  assign new_P3_ADD_467_U23 = ~P3_REIP_REG_11_;
  assign new_P3_ADD_467_U24 = ~P3_REIP_REG_11_ | ~new_P3_ADD_467_U102;
  assign new_P3_ADD_467_U25 = ~P3_REIP_REG_12_;
  assign new_P3_ADD_467_U26 = ~P3_REIP_REG_12_ | ~new_P3_ADD_467_U103;
  assign new_P3_ADD_467_U27 = ~P3_REIP_REG_13_;
  assign new_P3_ADD_467_U28 = ~P3_REIP_REG_13_ | ~new_P3_ADD_467_U104;
  assign new_P3_ADD_467_U29 = ~P3_REIP_REG_14_;
  assign new_P3_ADD_467_U30 = ~P3_REIP_REG_14_ | ~new_P3_ADD_467_U105;
  assign new_P3_ADD_467_U31 = ~P3_REIP_REG_15_;
  assign new_P3_ADD_467_U32 = ~P3_REIP_REG_15_ | ~new_P3_ADD_467_U106;
  assign new_P3_ADD_467_U33 = ~P3_REIP_REG_16_;
  assign new_P3_ADD_467_U34 = ~P3_REIP_REG_16_ | ~new_P3_ADD_467_U107;
  assign new_P3_ADD_467_U35 = ~P3_REIP_REG_17_;
  assign new_P3_ADD_467_U36 = ~P3_REIP_REG_17_ | ~new_P3_ADD_467_U108;
  assign new_P3_ADD_467_U37 = ~P3_REIP_REG_18_;
  assign new_P3_ADD_467_U38 = ~P3_REIP_REG_18_ | ~new_P3_ADD_467_U109;
  assign new_P3_ADD_467_U39 = ~P3_REIP_REG_19_;
  assign new_P3_ADD_467_U40 = ~P3_REIP_REG_19_ | ~new_P3_ADD_467_U110;
  assign new_P3_ADD_467_U41 = ~P3_REIP_REG_20_;
  assign new_P3_ADD_467_U42 = ~P3_REIP_REG_20_ | ~new_P3_ADD_467_U111;
  assign new_P3_ADD_467_U43 = ~P3_REIP_REG_21_;
  assign new_P3_ADD_467_U44 = ~P3_REIP_REG_21_ | ~new_P3_ADD_467_U112;
  assign new_P3_ADD_467_U45 = ~P3_REIP_REG_22_;
  assign new_P3_ADD_467_U46 = ~P3_REIP_REG_22_ | ~new_P3_ADD_467_U113;
  assign new_P3_ADD_467_U47 = ~P3_REIP_REG_23_;
  assign new_P3_ADD_467_U48 = ~P3_REIP_REG_23_ | ~new_P3_ADD_467_U114;
  assign new_P3_ADD_467_U49 = ~P3_REIP_REG_24_;
  assign new_P3_ADD_467_U50 = ~P3_REIP_REG_24_ | ~new_P3_ADD_467_U115;
  assign new_P3_ADD_467_U51 = ~P3_REIP_REG_25_;
  assign new_P3_ADD_467_U52 = ~P3_REIP_REG_25_ | ~new_P3_ADD_467_U116;
  assign new_P3_ADD_467_U53 = ~P3_REIP_REG_26_;
  assign new_P3_ADD_467_U54 = ~P3_REIP_REG_26_ | ~new_P3_ADD_467_U117;
  assign new_P3_ADD_467_U55 = ~P3_REIP_REG_27_;
  assign new_P3_ADD_467_U56 = ~P3_REIP_REG_27_ | ~new_P3_ADD_467_U118;
  assign new_P3_ADD_467_U57 = ~P3_REIP_REG_28_;
  assign new_P3_ADD_467_U58 = ~P3_REIP_REG_28_ | ~new_P3_ADD_467_U119;
  assign new_P3_ADD_467_U59 = ~P3_REIP_REG_29_;
  assign new_P3_ADD_467_U60 = ~P3_REIP_REG_29_ | ~new_P3_ADD_467_U120;
  assign new_P3_ADD_467_U61 = ~P3_REIP_REG_30_;
  assign new_P3_ADD_467_U62 = ~new_P3_ADD_467_U124 | ~new_P3_ADD_467_U123;
  assign new_P3_ADD_467_U63 = ~new_P3_ADD_467_U126 | ~new_P3_ADD_467_U125;
  assign new_P3_ADD_467_U64 = ~new_P3_ADD_467_U128 | ~new_P3_ADD_467_U127;
  assign new_P3_ADD_467_U65 = ~new_P3_ADD_467_U130 | ~new_P3_ADD_467_U129;
  assign new_P3_ADD_467_U66 = ~new_P3_ADD_467_U132 | ~new_P3_ADD_467_U131;
  assign new_P3_ADD_467_U67 = ~new_P3_ADD_467_U134 | ~new_P3_ADD_467_U133;
  assign new_P3_ADD_467_U68 = ~new_P3_ADD_467_U136 | ~new_P3_ADD_467_U135;
  assign new_P3_ADD_467_U69 = ~new_P3_ADD_467_U138 | ~new_P3_ADD_467_U137;
  assign new_P3_ADD_467_U70 = ~new_P3_ADD_467_U140 | ~new_P3_ADD_467_U139;
  assign new_P3_ADD_467_U71 = ~new_P3_ADD_467_U142 | ~new_P3_ADD_467_U141;
  assign new_P3_ADD_467_U72 = ~new_P3_ADD_467_U144 | ~new_P3_ADD_467_U143;
  assign new_P3_ADD_467_U73 = ~new_P3_ADD_467_U146 | ~new_P3_ADD_467_U145;
  assign new_P3_ADD_467_U74 = ~new_P3_ADD_467_U148 | ~new_P3_ADD_467_U147;
  assign new_P3_ADD_467_U75 = ~new_P3_ADD_467_U150 | ~new_P3_ADD_467_U149;
  assign new_P3_ADD_467_U76 = ~new_P3_ADD_467_U152 | ~new_P3_ADD_467_U151;
  assign new_P3_ADD_467_U77 = ~new_P3_ADD_467_U154 | ~new_P3_ADD_467_U153;
  assign new_P3_ADD_467_U78 = ~new_P3_ADD_467_U156 | ~new_P3_ADD_467_U155;
  assign new_P3_ADD_467_U79 = ~new_P3_ADD_467_U158 | ~new_P3_ADD_467_U157;
  assign new_P3_ADD_467_U80 = ~new_P3_ADD_467_U160 | ~new_P3_ADD_467_U159;
  assign new_P3_ADD_467_U81 = ~new_P3_ADD_467_U162 | ~new_P3_ADD_467_U161;
  assign new_P3_ADD_467_U82 = ~new_P3_ADD_467_U164 | ~new_P3_ADD_467_U163;
  assign new_P3_ADD_467_U83 = ~new_P3_ADD_467_U166 | ~new_P3_ADD_467_U165;
  assign new_P3_ADD_467_U84 = ~new_P3_ADD_467_U168 | ~new_P3_ADD_467_U167;
  assign new_P3_ADD_467_U85 = ~new_P3_ADD_467_U170 | ~new_P3_ADD_467_U169;
  assign new_P3_ADD_467_U86 = ~new_P3_ADD_467_U172 | ~new_P3_ADD_467_U171;
  assign new_P3_ADD_467_U87 = ~new_P3_ADD_467_U174 | ~new_P3_ADD_467_U173;
  assign new_P3_ADD_467_U88 = ~new_P3_ADD_467_U176 | ~new_P3_ADD_467_U175;
  assign new_P3_ADD_467_U89 = ~new_P3_ADD_467_U178 | ~new_P3_ADD_467_U177;
  assign new_P3_ADD_467_U90 = ~new_P3_ADD_467_U180 | ~new_P3_ADD_467_U179;
  assign new_P3_ADD_467_U91 = ~new_P3_ADD_467_U182 | ~new_P3_ADD_467_U181;
  assign new_P3_ADD_467_U92 = ~P3_REIP_REG_31_;
  assign new_P3_ADD_467_U93 = ~P3_REIP_REG_30_ | ~new_P3_ADD_467_U121;
  assign new_P3_ADD_467_U94 = ~new_P3_ADD_467_U6;
  assign new_P3_ADD_467_U95 = ~new_P3_ADD_467_U8;
  assign new_P3_ADD_467_U96 = ~new_P3_ADD_467_U10;
  assign new_P3_ADD_467_U97 = ~new_P3_ADD_467_U12;
  assign new_P3_ADD_467_U98 = ~new_P3_ADD_467_U14;
  assign new_P3_ADD_467_U99 = ~new_P3_ADD_467_U16;
  assign new_P3_ADD_467_U100 = ~new_P3_ADD_467_U19;
  assign new_P3_ADD_467_U101 = ~new_P3_ADD_467_U20;
  assign new_P3_ADD_467_U102 = ~new_P3_ADD_467_U22;
  assign new_P3_ADD_467_U103 = ~new_P3_ADD_467_U24;
  assign new_P3_ADD_467_U104 = ~new_P3_ADD_467_U26;
  assign new_P3_ADD_467_U105 = ~new_P3_ADD_467_U28;
  assign new_P3_ADD_467_U106 = ~new_P3_ADD_467_U30;
  assign new_P3_ADD_467_U107 = ~new_P3_ADD_467_U32;
  assign new_P3_ADD_467_U108 = ~new_P3_ADD_467_U34;
  assign new_P3_ADD_467_U109 = ~new_P3_ADD_467_U36;
  assign new_P3_ADD_467_U110 = ~new_P3_ADD_467_U38;
  assign new_P3_ADD_467_U111 = ~new_P3_ADD_467_U40;
  assign new_P3_ADD_467_U112 = ~new_P3_ADD_467_U42;
  assign new_P3_ADD_467_U113 = ~new_P3_ADD_467_U44;
  assign new_P3_ADD_467_U114 = ~new_P3_ADD_467_U46;
  assign new_P3_ADD_467_U115 = ~new_P3_ADD_467_U48;
  assign new_P3_ADD_467_U116 = ~new_P3_ADD_467_U50;
  assign new_P3_ADD_467_U117 = ~new_P3_ADD_467_U52;
  assign new_P3_ADD_467_U118 = ~new_P3_ADD_467_U54;
  assign new_P3_ADD_467_U119 = ~new_P3_ADD_467_U56;
  assign new_P3_ADD_467_U120 = ~new_P3_ADD_467_U58;
  assign new_P3_ADD_467_U121 = ~new_P3_ADD_467_U60;
  assign new_P3_ADD_467_U122 = ~new_P3_ADD_467_U93;
  assign new_P3_ADD_467_U123 = ~P3_REIP_REG_9_ | ~new_P3_ADD_467_U19;
  assign new_P3_ADD_467_U124 = ~new_P3_ADD_467_U100 | ~new_P3_ADD_467_U18;
  assign new_P3_ADD_467_U125 = ~P3_REIP_REG_8_ | ~new_P3_ADD_467_U16;
  assign new_P3_ADD_467_U126 = ~new_P3_ADD_467_U99 | ~new_P3_ADD_467_U17;
  assign new_P3_ADD_467_U127 = ~P3_REIP_REG_7_ | ~new_P3_ADD_467_U14;
  assign new_P3_ADD_467_U128 = ~new_P3_ADD_467_U98 | ~new_P3_ADD_467_U15;
  assign new_P3_ADD_467_U129 = ~P3_REIP_REG_6_ | ~new_P3_ADD_467_U12;
  assign new_P3_ADD_467_U130 = ~new_P3_ADD_467_U97 | ~new_P3_ADD_467_U13;
  assign new_P3_ADD_467_U131 = ~P3_REIP_REG_5_ | ~new_P3_ADD_467_U10;
  assign new_P3_ADD_467_U132 = ~new_P3_ADD_467_U96 | ~new_P3_ADD_467_U11;
  assign new_P3_ADD_467_U133 = ~P3_REIP_REG_4_ | ~new_P3_ADD_467_U8;
  assign new_P3_ADD_467_U134 = ~new_P3_ADD_467_U95 | ~new_P3_ADD_467_U9;
  assign new_P3_ADD_467_U135 = ~P3_REIP_REG_3_ | ~new_P3_ADD_467_U6;
  assign new_P3_ADD_467_U136 = ~new_P3_ADD_467_U94 | ~new_P3_ADD_467_U7;
  assign new_P3_ADD_467_U137 = ~P3_REIP_REG_31_ | ~new_P3_ADD_467_U93;
  assign new_P3_ADD_467_U138 = ~new_P3_ADD_467_U122 | ~new_P3_ADD_467_U92;
  assign new_P3_ADD_467_U139 = ~P3_REIP_REG_30_ | ~new_P3_ADD_467_U60;
  assign new_P3_ADD_467_U140 = ~new_P3_ADD_467_U121 | ~new_P3_ADD_467_U61;
  assign new_P3_ADD_467_U141 = ~P3_REIP_REG_2_ | ~new_P3_ADD_467_U4;
  assign new_P3_ADD_467_U142 = ~P3_REIP_REG_1_ | ~new_P3_ADD_467_U5;
  assign new_P3_ADD_467_U143 = ~P3_REIP_REG_29_ | ~new_P3_ADD_467_U58;
  assign new_P3_ADD_467_U144 = ~new_P3_ADD_467_U120 | ~new_P3_ADD_467_U59;
  assign new_P3_ADD_467_U145 = ~P3_REIP_REG_28_ | ~new_P3_ADD_467_U56;
  assign new_P3_ADD_467_U146 = ~new_P3_ADD_467_U119 | ~new_P3_ADD_467_U57;
  assign new_P3_ADD_467_U147 = ~P3_REIP_REG_27_ | ~new_P3_ADD_467_U54;
  assign new_P3_ADD_467_U148 = ~new_P3_ADD_467_U118 | ~new_P3_ADD_467_U55;
  assign new_P3_ADD_467_U149 = ~P3_REIP_REG_26_ | ~new_P3_ADD_467_U52;
  assign new_P3_ADD_467_U150 = ~new_P3_ADD_467_U117 | ~new_P3_ADD_467_U53;
  assign new_P3_ADD_467_U151 = ~P3_REIP_REG_25_ | ~new_P3_ADD_467_U50;
  assign new_P3_ADD_467_U152 = ~new_P3_ADD_467_U116 | ~new_P3_ADD_467_U51;
  assign new_P3_ADD_467_U153 = ~P3_REIP_REG_24_ | ~new_P3_ADD_467_U48;
  assign new_P3_ADD_467_U154 = ~new_P3_ADD_467_U115 | ~new_P3_ADD_467_U49;
  assign new_P3_ADD_467_U155 = ~P3_REIP_REG_23_ | ~new_P3_ADD_467_U46;
  assign new_P3_ADD_467_U156 = ~new_P3_ADD_467_U114 | ~new_P3_ADD_467_U47;
  assign new_P3_ADD_467_U157 = ~P3_REIP_REG_22_ | ~new_P3_ADD_467_U44;
  assign new_P3_ADD_467_U158 = ~new_P3_ADD_467_U113 | ~new_P3_ADD_467_U45;
  assign new_P3_ADD_467_U159 = ~P3_REIP_REG_21_ | ~new_P3_ADD_467_U42;
  assign new_P3_ADD_467_U160 = ~new_P3_ADD_467_U112 | ~new_P3_ADD_467_U43;
  assign new_P3_ADD_467_U161 = ~P3_REIP_REG_20_ | ~new_P3_ADD_467_U40;
  assign new_P3_ADD_467_U162 = ~new_P3_ADD_467_U111 | ~new_P3_ADD_467_U41;
  assign new_P3_ADD_467_U163 = ~P3_REIP_REG_19_ | ~new_P3_ADD_467_U38;
  assign new_P3_ADD_467_U164 = ~new_P3_ADD_467_U110 | ~new_P3_ADD_467_U39;
  assign new_P3_ADD_467_U165 = ~P3_REIP_REG_18_ | ~new_P3_ADD_467_U36;
  assign new_P3_ADD_467_U166 = ~new_P3_ADD_467_U109 | ~new_P3_ADD_467_U37;
  assign new_P3_ADD_467_U167 = ~P3_REIP_REG_17_ | ~new_P3_ADD_467_U34;
  assign new_P3_ADD_467_U168 = ~new_P3_ADD_467_U108 | ~new_P3_ADD_467_U35;
  assign new_P3_ADD_467_U169 = ~P3_REIP_REG_16_ | ~new_P3_ADD_467_U32;
  assign new_P3_ADD_467_U170 = ~new_P3_ADD_467_U107 | ~new_P3_ADD_467_U33;
  assign new_P3_ADD_467_U171 = ~P3_REIP_REG_15_ | ~new_P3_ADD_467_U30;
  assign new_P3_ADD_467_U172 = ~new_P3_ADD_467_U106 | ~new_P3_ADD_467_U31;
  assign new_P3_ADD_467_U173 = ~P3_REIP_REG_14_ | ~new_P3_ADD_467_U28;
  assign new_P3_ADD_467_U174 = ~new_P3_ADD_467_U105 | ~new_P3_ADD_467_U29;
  assign new_P3_ADD_467_U175 = ~P3_REIP_REG_13_ | ~new_P3_ADD_467_U26;
  assign new_P3_ADD_467_U176 = ~new_P3_ADD_467_U104 | ~new_P3_ADD_467_U27;
  assign new_P3_ADD_467_U177 = ~P3_REIP_REG_12_ | ~new_P3_ADD_467_U24;
  assign new_P3_ADD_467_U178 = ~new_P3_ADD_467_U103 | ~new_P3_ADD_467_U25;
  assign new_P3_ADD_467_U179 = ~P3_REIP_REG_11_ | ~new_P3_ADD_467_U22;
  assign new_P3_ADD_467_U180 = ~new_P3_ADD_467_U102 | ~new_P3_ADD_467_U23;
  assign new_P3_ADD_467_U181 = ~P3_REIP_REG_10_ | ~new_P3_ADD_467_U20;
  assign new_P3_ADD_467_U182 = ~new_P3_ADD_467_U101 | ~new_P3_ADD_467_U21;
  assign new_P3_ADD_430_U4 = ~P3_REIP_REG_1_;
  assign new_P3_ADD_430_U5 = ~P3_REIP_REG_2_;
  assign new_P3_ADD_430_U6 = ~P3_REIP_REG_2_ | ~P3_REIP_REG_1_;
  assign new_P3_ADD_430_U7 = ~P3_REIP_REG_3_;
  assign new_P3_ADD_430_U8 = ~P3_REIP_REG_3_ | ~new_P3_ADD_430_U94;
  assign new_P3_ADD_430_U9 = ~P3_REIP_REG_4_;
  assign new_P3_ADD_430_U10 = ~P3_REIP_REG_4_ | ~new_P3_ADD_430_U95;
  assign new_P3_ADD_430_U11 = ~P3_REIP_REG_5_;
  assign new_P3_ADD_430_U12 = ~P3_REIP_REG_5_ | ~new_P3_ADD_430_U96;
  assign new_P3_ADD_430_U13 = ~P3_REIP_REG_6_;
  assign new_P3_ADD_430_U14 = ~P3_REIP_REG_6_ | ~new_P3_ADD_430_U97;
  assign new_P3_ADD_430_U15 = ~P3_REIP_REG_7_;
  assign new_P3_ADD_430_U16 = ~P3_REIP_REG_7_ | ~new_P3_ADD_430_U98;
  assign new_P3_ADD_430_U17 = ~P3_REIP_REG_8_;
  assign new_P3_ADD_430_U18 = ~P3_REIP_REG_9_;
  assign new_P3_ADD_430_U19 = ~P3_REIP_REG_8_ | ~new_P3_ADD_430_U99;
  assign new_P3_ADD_430_U20 = ~new_P3_ADD_430_U100 | ~P3_REIP_REG_9_;
  assign new_P3_ADD_430_U21 = ~P3_REIP_REG_10_;
  assign new_P3_ADD_430_U22 = ~P3_REIP_REG_10_ | ~new_P3_ADD_430_U101;
  assign new_P3_ADD_430_U23 = ~P3_REIP_REG_11_;
  assign new_P3_ADD_430_U24 = ~P3_REIP_REG_11_ | ~new_P3_ADD_430_U102;
  assign new_P3_ADD_430_U25 = ~P3_REIP_REG_12_;
  assign new_P3_ADD_430_U26 = ~P3_REIP_REG_12_ | ~new_P3_ADD_430_U103;
  assign new_P3_ADD_430_U27 = ~P3_REIP_REG_13_;
  assign new_P3_ADD_430_U28 = ~P3_REIP_REG_13_ | ~new_P3_ADD_430_U104;
  assign new_P3_ADD_430_U29 = ~P3_REIP_REG_14_;
  assign new_P3_ADD_430_U30 = ~P3_REIP_REG_14_ | ~new_P3_ADD_430_U105;
  assign new_P3_ADD_430_U31 = ~P3_REIP_REG_15_;
  assign new_P3_ADD_430_U32 = ~P3_REIP_REG_15_ | ~new_P3_ADD_430_U106;
  assign new_P3_ADD_430_U33 = ~P3_REIP_REG_16_;
  assign new_P3_ADD_430_U34 = ~P3_REIP_REG_16_ | ~new_P3_ADD_430_U107;
  assign new_P3_ADD_430_U35 = ~P3_REIP_REG_17_;
  assign new_P3_ADD_430_U36 = ~P3_REIP_REG_17_ | ~new_P3_ADD_430_U108;
  assign new_P3_ADD_430_U37 = ~P3_REIP_REG_18_;
  assign new_P3_ADD_430_U38 = ~P3_REIP_REG_18_ | ~new_P3_ADD_430_U109;
  assign new_P3_ADD_430_U39 = ~P3_REIP_REG_19_;
  assign new_P3_ADD_430_U40 = ~P3_REIP_REG_19_ | ~new_P3_ADD_430_U110;
  assign new_P3_ADD_430_U41 = ~P3_REIP_REG_20_;
  assign new_P3_ADD_430_U42 = ~P3_REIP_REG_20_ | ~new_P3_ADD_430_U111;
  assign new_P3_ADD_430_U43 = ~P3_REIP_REG_21_;
  assign new_P3_ADD_430_U44 = ~P3_REIP_REG_21_ | ~new_P3_ADD_430_U112;
  assign new_P3_ADD_430_U45 = ~P3_REIP_REG_22_;
  assign new_P3_ADD_430_U46 = ~P3_REIP_REG_22_ | ~new_P3_ADD_430_U113;
  assign new_P3_ADD_430_U47 = ~P3_REIP_REG_23_;
  assign new_P3_ADD_430_U48 = ~P3_REIP_REG_23_ | ~new_P3_ADD_430_U114;
  assign new_P3_ADD_430_U49 = ~P3_REIP_REG_24_;
  assign new_P3_ADD_430_U50 = ~P3_REIP_REG_24_ | ~new_P3_ADD_430_U115;
  assign new_P3_ADD_430_U51 = ~P3_REIP_REG_25_;
  assign new_P3_ADD_430_U52 = ~P3_REIP_REG_25_ | ~new_P3_ADD_430_U116;
  assign new_P3_ADD_430_U53 = ~P3_REIP_REG_26_;
  assign new_P3_ADD_430_U54 = ~P3_REIP_REG_26_ | ~new_P3_ADD_430_U117;
  assign new_P3_ADD_430_U55 = ~P3_REIP_REG_27_;
  assign new_P3_ADD_430_U56 = ~P3_REIP_REG_27_ | ~new_P3_ADD_430_U118;
  assign new_P3_ADD_430_U57 = ~P3_REIP_REG_28_;
  assign new_P3_ADD_430_U58 = ~P3_REIP_REG_28_ | ~new_P3_ADD_430_U119;
  assign new_P3_ADD_430_U59 = ~P3_REIP_REG_29_;
  assign new_P3_ADD_430_U60 = ~P3_REIP_REG_29_ | ~new_P3_ADD_430_U120;
  assign new_P3_ADD_430_U61 = ~P3_REIP_REG_30_;
  assign new_P3_ADD_430_U62 = ~new_P3_ADD_430_U124 | ~new_P3_ADD_430_U123;
  assign new_P3_ADD_430_U63 = ~new_P3_ADD_430_U126 | ~new_P3_ADD_430_U125;
  assign new_P3_ADD_430_U64 = ~new_P3_ADD_430_U128 | ~new_P3_ADD_430_U127;
  assign new_P3_ADD_430_U65 = ~new_P3_ADD_430_U130 | ~new_P3_ADD_430_U129;
  assign new_P3_ADD_430_U66 = ~new_P3_ADD_430_U132 | ~new_P3_ADD_430_U131;
  assign new_P3_ADD_430_U67 = ~new_P3_ADD_430_U134 | ~new_P3_ADD_430_U133;
  assign new_P3_ADD_430_U68 = ~new_P3_ADD_430_U136 | ~new_P3_ADD_430_U135;
  assign new_P3_ADD_430_U69 = ~new_P3_ADD_430_U138 | ~new_P3_ADD_430_U137;
  assign new_P3_ADD_430_U70 = ~new_P3_ADD_430_U140 | ~new_P3_ADD_430_U139;
  assign new_P3_ADD_430_U71 = ~new_P3_ADD_430_U142 | ~new_P3_ADD_430_U141;
  assign new_P3_ADD_430_U72 = ~new_P3_ADD_430_U144 | ~new_P3_ADD_430_U143;
  assign new_P3_ADD_430_U73 = ~new_P3_ADD_430_U146 | ~new_P3_ADD_430_U145;
  assign new_P3_ADD_430_U74 = ~new_P3_ADD_430_U148 | ~new_P3_ADD_430_U147;
  assign new_P3_ADD_430_U75 = ~new_P3_ADD_430_U150 | ~new_P3_ADD_430_U149;
  assign new_P3_ADD_430_U76 = ~new_P3_ADD_430_U152 | ~new_P3_ADD_430_U151;
  assign new_P3_ADD_430_U77 = ~new_P3_ADD_430_U154 | ~new_P3_ADD_430_U153;
  assign new_P3_ADD_430_U78 = ~new_P3_ADD_430_U156 | ~new_P3_ADD_430_U155;
  assign new_P3_ADD_430_U79 = ~new_P3_ADD_430_U158 | ~new_P3_ADD_430_U157;
  assign new_P3_ADD_430_U80 = ~new_P3_ADD_430_U160 | ~new_P3_ADD_430_U159;
  assign new_P3_ADD_430_U81 = ~new_P3_ADD_430_U162 | ~new_P3_ADD_430_U161;
  assign new_P3_ADD_430_U82 = ~new_P3_ADD_430_U164 | ~new_P3_ADD_430_U163;
  assign new_P3_ADD_430_U83 = ~new_P3_ADD_430_U166 | ~new_P3_ADD_430_U165;
  assign new_P3_ADD_430_U84 = ~new_P3_ADD_430_U168 | ~new_P3_ADD_430_U167;
  assign new_P3_ADD_430_U85 = ~new_P3_ADD_430_U170 | ~new_P3_ADD_430_U169;
  assign new_P3_ADD_430_U86 = ~new_P3_ADD_430_U172 | ~new_P3_ADD_430_U171;
  assign new_P3_ADD_430_U87 = ~new_P3_ADD_430_U174 | ~new_P3_ADD_430_U173;
  assign new_P3_ADD_430_U88 = ~new_P3_ADD_430_U176 | ~new_P3_ADD_430_U175;
  assign new_P3_ADD_430_U89 = ~new_P3_ADD_430_U178 | ~new_P3_ADD_430_U177;
  assign new_P3_ADD_430_U90 = ~new_P3_ADD_430_U180 | ~new_P3_ADD_430_U179;
  assign new_P3_ADD_430_U91 = ~new_P3_ADD_430_U182 | ~new_P3_ADD_430_U181;
  assign new_P3_ADD_430_U92 = ~P3_REIP_REG_31_;
  assign new_P3_ADD_430_U93 = ~P3_REIP_REG_30_ | ~new_P3_ADD_430_U121;
  assign new_P3_ADD_430_U94 = ~new_P3_ADD_430_U6;
  assign new_P3_ADD_430_U95 = ~new_P3_ADD_430_U8;
  assign new_P3_ADD_430_U96 = ~new_P3_ADD_430_U10;
  assign new_P3_ADD_430_U97 = ~new_P3_ADD_430_U12;
  assign new_P3_ADD_430_U98 = ~new_P3_ADD_430_U14;
  assign new_P3_ADD_430_U99 = ~new_P3_ADD_430_U16;
  assign new_P3_ADD_430_U100 = ~new_P3_ADD_430_U19;
  assign new_P3_ADD_430_U101 = ~new_P3_ADD_430_U20;
  assign new_P3_ADD_430_U102 = ~new_P3_ADD_430_U22;
  assign new_P3_ADD_430_U103 = ~new_P3_ADD_430_U24;
  assign new_P3_ADD_430_U104 = ~new_P3_ADD_430_U26;
  assign new_P3_ADD_430_U105 = ~new_P3_ADD_430_U28;
  assign new_P3_ADD_430_U106 = ~new_P3_ADD_430_U30;
  assign new_P3_ADD_430_U107 = ~new_P3_ADD_430_U32;
  assign new_P3_ADD_430_U108 = ~new_P3_ADD_430_U34;
  assign new_P3_ADD_430_U109 = ~new_P3_ADD_430_U36;
  assign new_P3_ADD_430_U110 = ~new_P3_ADD_430_U38;
  assign new_P3_ADD_430_U111 = ~new_P3_ADD_430_U40;
  assign new_P3_ADD_430_U112 = ~new_P3_ADD_430_U42;
  assign new_P3_ADD_430_U113 = ~new_P3_ADD_430_U44;
  assign new_P3_ADD_430_U114 = ~new_P3_ADD_430_U46;
  assign new_P3_ADD_430_U115 = ~new_P3_ADD_430_U48;
  assign new_P3_ADD_430_U116 = ~new_P3_ADD_430_U50;
  assign new_P3_ADD_430_U117 = ~new_P3_ADD_430_U52;
  assign new_P3_ADD_430_U118 = ~new_P3_ADD_430_U54;
  assign new_P3_ADD_430_U119 = ~new_P3_ADD_430_U56;
  assign new_P3_ADD_430_U120 = ~new_P3_ADD_430_U58;
  assign new_P3_ADD_430_U121 = ~new_P3_ADD_430_U60;
  assign new_P3_ADD_430_U122 = ~new_P3_ADD_430_U93;
  assign new_P3_ADD_430_U123 = ~P3_REIP_REG_9_ | ~new_P3_ADD_430_U19;
  assign new_P3_ADD_430_U124 = ~new_P3_ADD_430_U100 | ~new_P3_ADD_430_U18;
  assign new_P3_ADD_430_U125 = ~P3_REIP_REG_8_ | ~new_P3_ADD_430_U16;
  assign new_P3_ADD_430_U126 = ~new_P3_ADD_430_U99 | ~new_P3_ADD_430_U17;
  assign new_P3_ADD_430_U127 = ~P3_REIP_REG_7_ | ~new_P3_ADD_430_U14;
  assign new_P3_ADD_430_U128 = ~new_P3_ADD_430_U98 | ~new_P3_ADD_430_U15;
  assign new_P3_ADD_430_U129 = ~P3_REIP_REG_6_ | ~new_P3_ADD_430_U12;
  assign new_P3_ADD_430_U130 = ~new_P3_ADD_430_U97 | ~new_P3_ADD_430_U13;
  assign new_P3_ADD_430_U131 = ~P3_REIP_REG_5_ | ~new_P3_ADD_430_U10;
  assign new_P3_ADD_430_U132 = ~new_P3_ADD_430_U96 | ~new_P3_ADD_430_U11;
  assign new_P3_ADD_430_U133 = ~P3_REIP_REG_4_ | ~new_P3_ADD_430_U8;
  assign new_P3_ADD_430_U134 = ~new_P3_ADD_430_U95 | ~new_P3_ADD_430_U9;
  assign new_P3_ADD_430_U135 = ~P3_REIP_REG_3_ | ~new_P3_ADD_430_U6;
  assign new_P3_ADD_430_U136 = ~new_P3_ADD_430_U94 | ~new_P3_ADD_430_U7;
  assign new_P3_ADD_430_U137 = ~P3_REIP_REG_31_ | ~new_P3_ADD_430_U93;
  assign new_P3_ADD_430_U138 = ~new_P3_ADD_430_U122 | ~new_P3_ADD_430_U92;
  assign new_P3_ADD_430_U139 = ~P3_REIP_REG_30_ | ~new_P3_ADD_430_U60;
  assign new_P3_ADD_430_U140 = ~new_P3_ADD_430_U121 | ~new_P3_ADD_430_U61;
  assign new_P3_ADD_430_U141 = ~P3_REIP_REG_2_ | ~new_P3_ADD_430_U4;
  assign new_P3_ADD_430_U142 = ~P3_REIP_REG_1_ | ~new_P3_ADD_430_U5;
  assign new_P3_ADD_430_U143 = ~P3_REIP_REG_29_ | ~new_P3_ADD_430_U58;
  assign new_P3_ADD_430_U144 = ~new_P3_ADD_430_U120 | ~new_P3_ADD_430_U59;
  assign new_P3_ADD_430_U145 = ~P3_REIP_REG_28_ | ~new_P3_ADD_430_U56;
  assign new_P3_ADD_430_U146 = ~new_P3_ADD_430_U119 | ~new_P3_ADD_430_U57;
  assign new_P3_ADD_430_U147 = ~P3_REIP_REG_27_ | ~new_P3_ADD_430_U54;
  assign new_P3_ADD_430_U148 = ~new_P3_ADD_430_U118 | ~new_P3_ADD_430_U55;
  assign new_P3_ADD_430_U149 = ~P3_REIP_REG_26_ | ~new_P3_ADD_430_U52;
  assign new_P3_ADD_430_U150 = ~new_P3_ADD_430_U117 | ~new_P3_ADD_430_U53;
  assign new_P3_ADD_430_U151 = ~P3_REIP_REG_25_ | ~new_P3_ADD_430_U50;
  assign new_P3_ADD_430_U152 = ~new_P3_ADD_430_U116 | ~new_P3_ADD_430_U51;
  assign new_P3_ADD_430_U153 = ~P3_REIP_REG_24_ | ~new_P3_ADD_430_U48;
  assign new_P3_ADD_430_U154 = ~new_P3_ADD_430_U115 | ~new_P3_ADD_430_U49;
  assign new_P3_ADD_430_U155 = ~P3_REIP_REG_23_ | ~new_P3_ADD_430_U46;
  assign new_P3_ADD_430_U156 = ~new_P3_ADD_430_U114 | ~new_P3_ADD_430_U47;
  assign new_P3_ADD_430_U157 = ~P3_REIP_REG_22_ | ~new_P3_ADD_430_U44;
  assign new_P3_ADD_430_U158 = ~new_P3_ADD_430_U113 | ~new_P3_ADD_430_U45;
  assign new_P3_ADD_430_U159 = ~P3_REIP_REG_21_ | ~new_P3_ADD_430_U42;
  assign new_P3_ADD_430_U160 = ~new_P3_ADD_430_U112 | ~new_P3_ADD_430_U43;
  assign new_P3_ADD_430_U161 = ~P3_REIP_REG_20_ | ~new_P3_ADD_430_U40;
  assign new_P3_ADD_430_U162 = ~new_P3_ADD_430_U111 | ~new_P3_ADD_430_U41;
  assign new_P3_ADD_430_U163 = ~P3_REIP_REG_19_ | ~new_P3_ADD_430_U38;
  assign new_P3_ADD_430_U164 = ~new_P3_ADD_430_U110 | ~new_P3_ADD_430_U39;
  assign new_P3_ADD_430_U165 = ~P3_REIP_REG_18_ | ~new_P3_ADD_430_U36;
  assign new_P3_ADD_430_U166 = ~new_P3_ADD_430_U109 | ~new_P3_ADD_430_U37;
  assign new_P3_ADD_430_U167 = ~P3_REIP_REG_17_ | ~new_P3_ADD_430_U34;
  assign new_P3_ADD_430_U168 = ~new_P3_ADD_430_U108 | ~new_P3_ADD_430_U35;
  assign new_P3_ADD_430_U169 = ~P3_REIP_REG_16_ | ~new_P3_ADD_430_U32;
  assign new_P3_ADD_430_U170 = ~new_P3_ADD_430_U107 | ~new_P3_ADD_430_U33;
  assign new_P3_ADD_430_U171 = ~P3_REIP_REG_15_ | ~new_P3_ADD_430_U30;
  assign new_P3_ADD_430_U172 = ~new_P3_ADD_430_U106 | ~new_P3_ADD_430_U31;
  assign new_P3_ADD_430_U173 = ~P3_REIP_REG_14_ | ~new_P3_ADD_430_U28;
  assign new_P3_ADD_430_U174 = ~new_P3_ADD_430_U105 | ~new_P3_ADD_430_U29;
  assign new_P3_ADD_430_U175 = ~P3_REIP_REG_13_ | ~new_P3_ADD_430_U26;
  assign new_P3_ADD_430_U176 = ~new_P3_ADD_430_U104 | ~new_P3_ADD_430_U27;
  assign new_P3_ADD_430_U177 = ~P3_REIP_REG_12_ | ~new_P3_ADD_430_U24;
  assign new_P3_ADD_430_U178 = ~new_P3_ADD_430_U103 | ~new_P3_ADD_430_U25;
  assign new_P3_ADD_430_U179 = ~P3_REIP_REG_11_ | ~new_P3_ADD_430_U22;
  assign new_P3_ADD_430_U180 = ~new_P3_ADD_430_U102 | ~new_P3_ADD_430_U23;
  assign new_P3_ADD_430_U181 = ~P3_REIP_REG_10_ | ~new_P3_ADD_430_U20;
  assign new_P3_ADD_430_U182 = ~new_P3_ADD_430_U101 | ~new_P3_ADD_430_U21;
  assign new_P3_ADD_380_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_380_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_380_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_380_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_380_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_380_U98;
  assign new_P3_ADD_380_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_380_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_380_U99;
  assign new_P3_ADD_380_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_380_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_380_U100;
  assign new_P3_ADD_380_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_380_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_380_U101;
  assign new_P3_ADD_380_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_380_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_380_U102;
  assign new_P3_ADD_380_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_380_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_380_U103;
  assign new_P3_ADD_380_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_380_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_380_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_380_U104;
  assign new_P3_ADD_380_U23 = ~new_P3_ADD_380_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_380_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_380_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_380_U106;
  assign new_P3_ADD_380_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_380_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_380_U107;
  assign new_P3_ADD_380_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_380_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_380_U108;
  assign new_P3_ADD_380_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_380_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_380_U109;
  assign new_P3_ADD_380_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_380_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_380_U110;
  assign new_P3_ADD_380_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_380_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_380_U111;
  assign new_P3_ADD_380_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_380_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_380_U112;
  assign new_P3_ADD_380_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_380_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_380_U113;
  assign new_P3_ADD_380_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_380_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_380_U114;
  assign new_P3_ADD_380_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_380_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_380_U115;
  assign new_P3_ADD_380_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_380_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_380_U116;
  assign new_P3_ADD_380_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_380_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_380_U117;
  assign new_P3_ADD_380_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_380_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_380_U118;
  assign new_P3_ADD_380_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_380_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_380_U119;
  assign new_P3_ADD_380_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_380_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_380_U120;
  assign new_P3_ADD_380_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_380_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_380_U121;
  assign new_P3_ADD_380_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_380_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_380_U122;
  assign new_P3_ADD_380_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_380_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_380_U123;
  assign new_P3_ADD_380_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_380_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_380_U124;
  assign new_P3_ADD_380_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_380_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_380_U125;
  assign new_P3_ADD_380_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_380_U65 = ~new_P3_ADD_380_U129 | ~new_P3_ADD_380_U128;
  assign new_P3_ADD_380_U66 = ~new_P3_ADD_380_U131 | ~new_P3_ADD_380_U130;
  assign new_P3_ADD_380_U67 = ~new_P3_ADD_380_U133 | ~new_P3_ADD_380_U132;
  assign new_P3_ADD_380_U68 = ~new_P3_ADD_380_U135 | ~new_P3_ADD_380_U134;
  assign new_P3_ADD_380_U69 = ~new_P3_ADD_380_U137 | ~new_P3_ADD_380_U136;
  assign new_P3_ADD_380_U70 = ~new_P3_ADD_380_U139 | ~new_P3_ADD_380_U138;
  assign new_P3_ADD_380_U71 = ~new_P3_ADD_380_U141 | ~new_P3_ADD_380_U140;
  assign new_P3_ADD_380_U72 = ~new_P3_ADD_380_U143 | ~new_P3_ADD_380_U142;
  assign new_P3_ADD_380_U73 = ~new_P3_ADD_380_U145 | ~new_P3_ADD_380_U144;
  assign new_P3_ADD_380_U74 = ~new_P3_ADD_380_U147 | ~new_P3_ADD_380_U146;
  assign new_P3_ADD_380_U75 = ~new_P3_ADD_380_U149 | ~new_P3_ADD_380_U148;
  assign new_P3_ADD_380_U76 = ~new_P3_ADD_380_U151 | ~new_P3_ADD_380_U150;
  assign new_P3_ADD_380_U77 = ~new_P3_ADD_380_U153 | ~new_P3_ADD_380_U152;
  assign new_P3_ADD_380_U78 = ~new_P3_ADD_380_U155 | ~new_P3_ADD_380_U154;
  assign new_P3_ADD_380_U79 = ~new_P3_ADD_380_U157 | ~new_P3_ADD_380_U156;
  assign new_P3_ADD_380_U80 = ~new_P3_ADD_380_U159 | ~new_P3_ADD_380_U158;
  assign new_P3_ADD_380_U81 = ~new_P3_ADD_380_U161 | ~new_P3_ADD_380_U160;
  assign new_P3_ADD_380_U82 = ~new_P3_ADD_380_U163 | ~new_P3_ADD_380_U162;
  assign new_P3_ADD_380_U83 = ~new_P3_ADD_380_U165 | ~new_P3_ADD_380_U164;
  assign new_P3_ADD_380_U84 = ~new_P3_ADD_380_U167 | ~new_P3_ADD_380_U166;
  assign new_P3_ADD_380_U85 = ~new_P3_ADD_380_U169 | ~new_P3_ADD_380_U168;
  assign new_P3_ADD_380_U86 = ~new_P3_ADD_380_U171 | ~new_P3_ADD_380_U170;
  assign new_P3_ADD_380_U87 = ~new_P3_ADD_380_U173 | ~new_P3_ADD_380_U172;
  assign new_P3_ADD_380_U88 = ~new_P3_ADD_380_U175 | ~new_P3_ADD_380_U174;
  assign new_P3_ADD_380_U89 = ~new_P3_ADD_380_U177 | ~new_P3_ADD_380_U176;
  assign new_P3_ADD_380_U90 = ~new_P3_ADD_380_U179 | ~new_P3_ADD_380_U178;
  assign new_P3_ADD_380_U91 = ~new_P3_ADD_380_U181 | ~new_P3_ADD_380_U180;
  assign new_P3_ADD_380_U92 = ~new_P3_ADD_380_U183 | ~new_P3_ADD_380_U182;
  assign new_P3_ADD_380_U93 = ~new_P3_ADD_380_U185 | ~new_P3_ADD_380_U184;
  assign new_P3_ADD_380_U94 = ~new_P3_ADD_380_U187 | ~new_P3_ADD_380_U186;
  assign new_P3_ADD_380_U95 = ~new_P3_ADD_380_U189 | ~new_P3_ADD_380_U188;
  assign new_P3_ADD_380_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_380_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_380_U126;
  assign new_P3_ADD_380_U98 = ~new_P3_ADD_380_U7;
  assign new_P3_ADD_380_U99 = ~new_P3_ADD_380_U9;
  assign new_P3_ADD_380_U100 = ~new_P3_ADD_380_U11;
  assign new_P3_ADD_380_U101 = ~new_P3_ADD_380_U13;
  assign new_P3_ADD_380_U102 = ~new_P3_ADD_380_U15;
  assign new_P3_ADD_380_U103 = ~new_P3_ADD_380_U17;
  assign new_P3_ADD_380_U104 = ~new_P3_ADD_380_U19;
  assign new_P3_ADD_380_U105 = ~new_P3_ADD_380_U22;
  assign new_P3_ADD_380_U106 = ~new_P3_ADD_380_U23;
  assign new_P3_ADD_380_U107 = ~new_P3_ADD_380_U25;
  assign new_P3_ADD_380_U108 = ~new_P3_ADD_380_U27;
  assign new_P3_ADD_380_U109 = ~new_P3_ADD_380_U29;
  assign new_P3_ADD_380_U110 = ~new_P3_ADD_380_U31;
  assign new_P3_ADD_380_U111 = ~new_P3_ADD_380_U33;
  assign new_P3_ADD_380_U112 = ~new_P3_ADD_380_U35;
  assign new_P3_ADD_380_U113 = ~new_P3_ADD_380_U37;
  assign new_P3_ADD_380_U114 = ~new_P3_ADD_380_U39;
  assign new_P3_ADD_380_U115 = ~new_P3_ADD_380_U41;
  assign new_P3_ADD_380_U116 = ~new_P3_ADD_380_U43;
  assign new_P3_ADD_380_U117 = ~new_P3_ADD_380_U45;
  assign new_P3_ADD_380_U118 = ~new_P3_ADD_380_U47;
  assign new_P3_ADD_380_U119 = ~new_P3_ADD_380_U49;
  assign new_P3_ADD_380_U120 = ~new_P3_ADD_380_U51;
  assign new_P3_ADD_380_U121 = ~new_P3_ADD_380_U53;
  assign new_P3_ADD_380_U122 = ~new_P3_ADD_380_U55;
  assign new_P3_ADD_380_U123 = ~new_P3_ADD_380_U57;
  assign new_P3_ADD_380_U124 = ~new_P3_ADD_380_U59;
  assign new_P3_ADD_380_U125 = ~new_P3_ADD_380_U61;
  assign new_P3_ADD_380_U126 = ~new_P3_ADD_380_U63;
  assign new_P3_ADD_380_U127 = ~new_P3_ADD_380_U97;
  assign new_P3_ADD_380_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_380_U22;
  assign new_P3_ADD_380_U129 = ~new_P3_ADD_380_U105 | ~new_P3_ADD_380_U21;
  assign new_P3_ADD_380_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_380_U19;
  assign new_P3_ADD_380_U131 = ~new_P3_ADD_380_U104 | ~new_P3_ADD_380_U20;
  assign new_P3_ADD_380_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_380_U17;
  assign new_P3_ADD_380_U133 = ~new_P3_ADD_380_U103 | ~new_P3_ADD_380_U18;
  assign new_P3_ADD_380_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_380_U15;
  assign new_P3_ADD_380_U135 = ~new_P3_ADD_380_U102 | ~new_P3_ADD_380_U16;
  assign new_P3_ADD_380_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_380_U13;
  assign new_P3_ADD_380_U137 = ~new_P3_ADD_380_U101 | ~new_P3_ADD_380_U14;
  assign new_P3_ADD_380_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_380_U11;
  assign new_P3_ADD_380_U139 = ~new_P3_ADD_380_U100 | ~new_P3_ADD_380_U12;
  assign new_P3_ADD_380_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_380_U9;
  assign new_P3_ADD_380_U141 = ~new_P3_ADD_380_U99 | ~new_P3_ADD_380_U10;
  assign new_P3_ADD_380_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_380_U97;
  assign new_P3_ADD_380_U143 = ~new_P3_ADD_380_U127 | ~new_P3_ADD_380_U96;
  assign new_P3_ADD_380_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_380_U63;
  assign new_P3_ADD_380_U145 = ~new_P3_ADD_380_U126 | ~new_P3_ADD_380_U64;
  assign new_P3_ADD_380_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_380_U7;
  assign new_P3_ADD_380_U147 = ~new_P3_ADD_380_U98 | ~new_P3_ADD_380_U8;
  assign new_P3_ADD_380_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_380_U61;
  assign new_P3_ADD_380_U149 = ~new_P3_ADD_380_U125 | ~new_P3_ADD_380_U62;
  assign new_P3_ADD_380_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_380_U59;
  assign new_P3_ADD_380_U151 = ~new_P3_ADD_380_U124 | ~new_P3_ADD_380_U60;
  assign new_P3_ADD_380_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_380_U57;
  assign new_P3_ADD_380_U153 = ~new_P3_ADD_380_U123 | ~new_P3_ADD_380_U58;
  assign new_P3_ADD_380_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_380_U55;
  assign new_P3_ADD_380_U155 = ~new_P3_ADD_380_U122 | ~new_P3_ADD_380_U56;
  assign new_P3_ADD_380_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_380_U53;
  assign new_P3_ADD_380_U157 = ~new_P3_ADD_380_U121 | ~new_P3_ADD_380_U54;
  assign new_P3_ADD_380_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_380_U51;
  assign new_P3_ADD_380_U159 = ~new_P3_ADD_380_U120 | ~new_P3_ADD_380_U52;
  assign new_P3_ADD_380_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_380_U49;
  assign new_P3_ADD_380_U161 = ~new_P3_ADD_380_U119 | ~new_P3_ADD_380_U50;
  assign new_P3_ADD_380_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_380_U47;
  assign new_P3_ADD_380_U163 = ~new_P3_ADD_380_U118 | ~new_P3_ADD_380_U48;
  assign new_P3_ADD_380_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_380_U45;
  assign new_P3_ADD_380_U165 = ~new_P3_ADD_380_U117 | ~new_P3_ADD_380_U46;
  assign new_P3_ADD_380_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_380_U43;
  assign new_P3_ADD_380_U167 = ~new_P3_ADD_380_U116 | ~new_P3_ADD_380_U44;
  assign new_P3_ADD_380_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_380_U5;
  assign new_P3_ADD_380_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_380_U6;
  assign new_P3_ADD_380_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_380_U41;
  assign new_P3_ADD_380_U171 = ~new_P3_ADD_380_U115 | ~new_P3_ADD_380_U42;
  assign new_P3_ADD_380_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_380_U39;
  assign new_P3_ADD_380_U173 = ~new_P3_ADD_380_U114 | ~new_P3_ADD_380_U40;
  assign new_P3_ADD_380_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_380_U37;
  assign new_P3_ADD_380_U175 = ~new_P3_ADD_380_U113 | ~new_P3_ADD_380_U38;
  assign new_P3_ADD_380_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_380_U35;
  assign new_P3_ADD_380_U177 = ~new_P3_ADD_380_U112 | ~new_P3_ADD_380_U36;
  assign new_P3_ADD_380_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_380_U33;
  assign new_P3_ADD_380_U179 = ~new_P3_ADD_380_U111 | ~new_P3_ADD_380_U34;
  assign new_P3_ADD_380_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_380_U31;
  assign new_P3_ADD_380_U181 = ~new_P3_ADD_380_U110 | ~new_P3_ADD_380_U32;
  assign new_P3_ADD_380_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_380_U29;
  assign new_P3_ADD_380_U183 = ~new_P3_ADD_380_U109 | ~new_P3_ADD_380_U30;
  assign new_P3_ADD_380_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_380_U27;
  assign new_P3_ADD_380_U185 = ~new_P3_ADD_380_U108 | ~new_P3_ADD_380_U28;
  assign new_P3_ADD_380_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_380_U25;
  assign new_P3_ADD_380_U187 = ~new_P3_ADD_380_U107 | ~new_P3_ADD_380_U26;
  assign new_P3_ADD_380_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_380_U23;
  assign new_P3_ADD_380_U189 = ~new_P3_ADD_380_U106 | ~new_P3_ADD_380_U24;
  assign new_P3_GTE_370_U6 = ~new_P3_SUB_370_U6 & ~new_P3_GTE_370_U8;
  assign new_P3_GTE_370_U7 = new_P3_SUB_370_U21 & new_P3_GTE_370_U9;
  assign new_P3_GTE_370_U8 = ~new_P3_SUB_370_U20 & ~new_P3_SUB_370_U19 & ~new_P3_GTE_370_U7;
  assign new_P3_GTE_370_U9 = new_P3_SUB_370_U7 | new_P3_SUB_370_U22;
  assign new_P3_ADD_344_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_344_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_344_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_344_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_344_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_344_U98;
  assign new_P3_ADD_344_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_344_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_344_U99;
  assign new_P3_ADD_344_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_344_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_344_U100;
  assign new_P3_ADD_344_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_344_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_344_U101;
  assign new_P3_ADD_344_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_344_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_344_U102;
  assign new_P3_ADD_344_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_344_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_344_U103;
  assign new_P3_ADD_344_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_344_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_344_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_344_U104;
  assign new_P3_ADD_344_U23 = ~new_P3_ADD_344_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_344_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_344_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_344_U106;
  assign new_P3_ADD_344_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_344_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_344_U107;
  assign new_P3_ADD_344_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_344_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_344_U108;
  assign new_P3_ADD_344_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_344_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_344_U109;
  assign new_P3_ADD_344_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_344_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_344_U110;
  assign new_P3_ADD_344_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_344_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_344_U111;
  assign new_P3_ADD_344_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_344_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_344_U112;
  assign new_P3_ADD_344_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_344_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_344_U113;
  assign new_P3_ADD_344_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_344_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_344_U114;
  assign new_P3_ADD_344_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_344_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_344_U115;
  assign new_P3_ADD_344_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_344_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_344_U116;
  assign new_P3_ADD_344_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_344_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_344_U117;
  assign new_P3_ADD_344_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_344_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_344_U118;
  assign new_P3_ADD_344_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_344_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_344_U119;
  assign new_P3_ADD_344_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_344_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_344_U120;
  assign new_P3_ADD_344_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_344_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_344_U121;
  assign new_P3_ADD_344_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_344_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_344_U122;
  assign new_P3_ADD_344_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_344_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_344_U123;
  assign new_P3_ADD_344_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_344_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_344_U124;
  assign new_P3_ADD_344_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_344_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_344_U125;
  assign new_P3_ADD_344_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_344_U65 = ~new_P3_ADD_344_U129 | ~new_P3_ADD_344_U128;
  assign new_P3_ADD_344_U66 = ~new_P3_ADD_344_U131 | ~new_P3_ADD_344_U130;
  assign new_P3_ADD_344_U67 = ~new_P3_ADD_344_U133 | ~new_P3_ADD_344_U132;
  assign new_P3_ADD_344_U68 = ~new_P3_ADD_344_U135 | ~new_P3_ADD_344_U134;
  assign new_P3_ADD_344_U69 = ~new_P3_ADD_344_U137 | ~new_P3_ADD_344_U136;
  assign new_P3_ADD_344_U70 = ~new_P3_ADD_344_U139 | ~new_P3_ADD_344_U138;
  assign new_P3_ADD_344_U71 = ~new_P3_ADD_344_U141 | ~new_P3_ADD_344_U140;
  assign new_P3_ADD_344_U72 = ~new_P3_ADD_344_U143 | ~new_P3_ADD_344_U142;
  assign new_P3_ADD_344_U73 = ~new_P3_ADD_344_U145 | ~new_P3_ADD_344_U144;
  assign new_P3_ADD_344_U74 = ~new_P3_ADD_344_U147 | ~new_P3_ADD_344_U146;
  assign new_P3_ADD_344_U75 = ~new_P3_ADD_344_U149 | ~new_P3_ADD_344_U148;
  assign new_P3_ADD_344_U76 = ~new_P3_ADD_344_U151 | ~new_P3_ADD_344_U150;
  assign new_P3_ADD_344_U77 = ~new_P3_ADD_344_U153 | ~new_P3_ADD_344_U152;
  assign new_P3_ADD_344_U78 = ~new_P3_ADD_344_U155 | ~new_P3_ADD_344_U154;
  assign new_P3_ADD_344_U79 = ~new_P3_ADD_344_U157 | ~new_P3_ADD_344_U156;
  assign new_P3_ADD_344_U80 = ~new_P3_ADD_344_U159 | ~new_P3_ADD_344_U158;
  assign new_P3_ADD_344_U81 = ~new_P3_ADD_344_U161 | ~new_P3_ADD_344_U160;
  assign new_P3_ADD_344_U82 = ~new_P3_ADD_344_U163 | ~new_P3_ADD_344_U162;
  assign new_P3_ADD_344_U83 = ~new_P3_ADD_344_U165 | ~new_P3_ADD_344_U164;
  assign new_P3_ADD_344_U84 = ~new_P3_ADD_344_U167 | ~new_P3_ADD_344_U166;
  assign new_P3_ADD_344_U85 = ~new_P3_ADD_344_U169 | ~new_P3_ADD_344_U168;
  assign new_P3_ADD_344_U86 = ~new_P3_ADD_344_U171 | ~new_P3_ADD_344_U170;
  assign new_P3_ADD_344_U87 = ~new_P3_ADD_344_U173 | ~new_P3_ADD_344_U172;
  assign new_P3_ADD_344_U88 = ~new_P3_ADD_344_U175 | ~new_P3_ADD_344_U174;
  assign new_P3_ADD_344_U89 = ~new_P3_ADD_344_U177 | ~new_P3_ADD_344_U176;
  assign new_P3_ADD_344_U90 = ~new_P3_ADD_344_U179 | ~new_P3_ADD_344_U178;
  assign new_P3_ADD_344_U91 = ~new_P3_ADD_344_U181 | ~new_P3_ADD_344_U180;
  assign new_P3_ADD_344_U92 = ~new_P3_ADD_344_U183 | ~new_P3_ADD_344_U182;
  assign new_P3_ADD_344_U93 = ~new_P3_ADD_344_U185 | ~new_P3_ADD_344_U184;
  assign new_P3_ADD_344_U94 = ~new_P3_ADD_344_U187 | ~new_P3_ADD_344_U186;
  assign new_P3_ADD_344_U95 = ~new_P3_ADD_344_U189 | ~new_P3_ADD_344_U188;
  assign new_P3_ADD_344_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_344_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_344_U126;
  assign new_P3_ADD_344_U98 = ~new_P3_ADD_344_U7;
  assign new_P3_ADD_344_U99 = ~new_P3_ADD_344_U9;
  assign new_P3_ADD_344_U100 = ~new_P3_ADD_344_U11;
  assign new_P3_ADD_344_U101 = ~new_P3_ADD_344_U13;
  assign new_P3_ADD_344_U102 = ~new_P3_ADD_344_U15;
  assign new_P3_ADD_344_U103 = ~new_P3_ADD_344_U17;
  assign new_P3_ADD_344_U104 = ~new_P3_ADD_344_U19;
  assign new_P3_ADD_344_U105 = ~new_P3_ADD_344_U22;
  assign new_P3_ADD_344_U106 = ~new_P3_ADD_344_U23;
  assign new_P3_ADD_344_U107 = ~new_P3_ADD_344_U25;
  assign new_P3_ADD_344_U108 = ~new_P3_ADD_344_U27;
  assign new_P3_ADD_344_U109 = ~new_P3_ADD_344_U29;
  assign new_P3_ADD_344_U110 = ~new_P3_ADD_344_U31;
  assign new_P3_ADD_344_U111 = ~new_P3_ADD_344_U33;
  assign new_P3_ADD_344_U112 = ~new_P3_ADD_344_U35;
  assign new_P3_ADD_344_U113 = ~new_P3_ADD_344_U37;
  assign new_P3_ADD_344_U114 = ~new_P3_ADD_344_U39;
  assign new_P3_ADD_344_U115 = ~new_P3_ADD_344_U41;
  assign new_P3_ADD_344_U116 = ~new_P3_ADD_344_U43;
  assign new_P3_ADD_344_U117 = ~new_P3_ADD_344_U45;
  assign new_P3_ADD_344_U118 = ~new_P3_ADD_344_U47;
  assign new_P3_ADD_344_U119 = ~new_P3_ADD_344_U49;
  assign new_P3_ADD_344_U120 = ~new_P3_ADD_344_U51;
  assign new_P3_ADD_344_U121 = ~new_P3_ADD_344_U53;
  assign new_P3_ADD_344_U122 = ~new_P3_ADD_344_U55;
  assign new_P3_ADD_344_U123 = ~new_P3_ADD_344_U57;
  assign new_P3_ADD_344_U124 = ~new_P3_ADD_344_U59;
  assign new_P3_ADD_344_U125 = ~new_P3_ADD_344_U61;
  assign new_P3_ADD_344_U126 = ~new_P3_ADD_344_U63;
  assign new_P3_ADD_344_U127 = ~new_P3_ADD_344_U97;
  assign new_P3_ADD_344_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_344_U22;
  assign new_P3_ADD_344_U129 = ~new_P3_ADD_344_U105 | ~new_P3_ADD_344_U21;
  assign new_P3_ADD_344_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_344_U19;
  assign new_P3_ADD_344_U131 = ~new_P3_ADD_344_U104 | ~new_P3_ADD_344_U20;
  assign new_P3_ADD_344_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_344_U17;
  assign new_P3_ADD_344_U133 = ~new_P3_ADD_344_U103 | ~new_P3_ADD_344_U18;
  assign new_P3_ADD_344_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_344_U15;
  assign new_P3_ADD_344_U135 = ~new_P3_ADD_344_U102 | ~new_P3_ADD_344_U16;
  assign new_P3_ADD_344_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_344_U13;
  assign new_P3_ADD_344_U137 = ~new_P3_ADD_344_U101 | ~new_P3_ADD_344_U14;
  assign new_P3_ADD_344_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_344_U11;
  assign new_P3_ADD_344_U139 = ~new_P3_ADD_344_U100 | ~new_P3_ADD_344_U12;
  assign new_P3_ADD_344_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_344_U9;
  assign new_P3_ADD_344_U141 = ~new_P3_ADD_344_U99 | ~new_P3_ADD_344_U10;
  assign new_P3_ADD_344_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_344_U97;
  assign new_P3_ADD_344_U143 = ~new_P3_ADD_344_U127 | ~new_P3_ADD_344_U96;
  assign new_P3_ADD_344_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_344_U63;
  assign new_P3_ADD_344_U145 = ~new_P3_ADD_344_U126 | ~new_P3_ADD_344_U64;
  assign new_P3_ADD_344_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_344_U7;
  assign new_P3_ADD_344_U147 = ~new_P3_ADD_344_U98 | ~new_P3_ADD_344_U8;
  assign new_P3_ADD_344_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_344_U61;
  assign new_P3_ADD_344_U149 = ~new_P3_ADD_344_U125 | ~new_P3_ADD_344_U62;
  assign new_P3_ADD_344_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_344_U59;
  assign new_P3_ADD_344_U151 = ~new_P3_ADD_344_U124 | ~new_P3_ADD_344_U60;
  assign new_P3_ADD_344_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_344_U57;
  assign new_P3_ADD_344_U153 = ~new_P3_ADD_344_U123 | ~new_P3_ADD_344_U58;
  assign new_P3_ADD_344_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_344_U55;
  assign new_P3_ADD_344_U155 = ~new_P3_ADD_344_U122 | ~new_P3_ADD_344_U56;
  assign new_P3_ADD_344_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_344_U53;
  assign new_P3_ADD_344_U157 = ~new_P3_ADD_344_U121 | ~new_P3_ADD_344_U54;
  assign new_P3_ADD_344_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_344_U51;
  assign new_P3_ADD_344_U159 = ~new_P3_ADD_344_U120 | ~new_P3_ADD_344_U52;
  assign new_P3_ADD_344_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_344_U49;
  assign new_P3_ADD_344_U161 = ~new_P3_ADD_344_U119 | ~new_P3_ADD_344_U50;
  assign new_P3_ADD_344_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_344_U47;
  assign new_P3_ADD_344_U163 = ~new_P3_ADD_344_U118 | ~new_P3_ADD_344_U48;
  assign new_P3_ADD_344_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_344_U45;
  assign new_P3_ADD_344_U165 = ~new_P3_ADD_344_U117 | ~new_P3_ADD_344_U46;
  assign new_P3_ADD_344_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_344_U43;
  assign new_P3_ADD_344_U167 = ~new_P3_ADD_344_U116 | ~new_P3_ADD_344_U44;
  assign new_P3_ADD_344_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_344_U5;
  assign new_P3_ADD_344_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_344_U6;
  assign new_P3_ADD_344_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_344_U41;
  assign new_P3_ADD_344_U171 = ~new_P3_ADD_344_U115 | ~new_P3_ADD_344_U42;
  assign new_P3_ADD_344_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_344_U39;
  assign new_P3_ADD_344_U173 = ~new_P3_ADD_344_U114 | ~new_P3_ADD_344_U40;
  assign new_P3_ADD_344_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_344_U37;
  assign new_P3_ADD_344_U175 = ~new_P3_ADD_344_U113 | ~new_P3_ADD_344_U38;
  assign new_P3_ADD_344_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_344_U35;
  assign new_P3_ADD_344_U177 = ~new_P3_ADD_344_U112 | ~new_P3_ADD_344_U36;
  assign new_P3_ADD_344_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_344_U33;
  assign new_P3_ADD_344_U179 = ~new_P3_ADD_344_U111 | ~new_P3_ADD_344_U34;
  assign new_P3_ADD_344_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_344_U31;
  assign new_P3_ADD_344_U181 = ~new_P3_ADD_344_U110 | ~new_P3_ADD_344_U32;
  assign new_P3_ADD_344_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_344_U29;
  assign new_P3_ADD_344_U183 = ~new_P3_ADD_344_U109 | ~new_P3_ADD_344_U30;
  assign new_P3_ADD_344_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_344_U27;
  assign new_P3_ADD_344_U185 = ~new_P3_ADD_344_U108 | ~new_P3_ADD_344_U28;
  assign new_P3_ADD_344_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_344_U25;
  assign new_P3_ADD_344_U187 = ~new_P3_ADD_344_U107 | ~new_P3_ADD_344_U26;
  assign new_P3_ADD_344_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_344_U23;
  assign new_P3_ADD_344_U189 = ~new_P3_ADD_344_U106 | ~new_P3_ADD_344_U24;
  assign new_P3_LT_563_U6 = ~new_P3_LT_563_U27 | ~new_P3_LT_563_U28;
  assign new_P3_LT_563_U7 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_LT_563_U8 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_LT_563_U15;
  assign new_P3_LT_563_U9 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_LT_563_U10 = ~new_P3_U3306;
  assign new_P3_LT_563_U11 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_LT_563_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_LT_563_U13 = ~new_P3_U3305;
  assign new_P3_LT_563_U14 = ~new_P3_U3304;
  assign new_P3_LT_563_U15 = ~new_P3_U3308;
  assign new_P3_LT_563_U16 = ~new_P3_LT_563_U8;
  assign new_P3_LT_563_U17 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_LT_563_U16;
  assign new_P3_LT_563_U18 = ~new_P3_U3307 | ~new_P3_LT_563_U17;
  assign new_P3_LT_563_U19 = ~new_P3_LT_563_U8 | ~new_P3_LT_563_U9;
  assign new_P3_LT_563_U20 = ~new_P3_U3306 | ~new_P3_LT_563_U11;
  assign new_P3_LT_563_U21 = ~new_P3_LT_563_U18 | ~new_P3_LT_563_U19 | ~new_P3_LT_563_U20;
  assign new_P3_LT_563_U22 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_LT_563_U10;
  assign new_P3_LT_563_U23 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_LT_563_U13;
  assign new_P3_LT_563_U24 = ~new_P3_LT_563_U21 | ~new_P3_LT_563_U22 | ~new_P3_LT_563_U23;
  assign new_P3_LT_563_U25 = ~new_P3_U3305 | ~new_P3_LT_563_U12;
  assign new_P3_LT_563_U26 = ~new_P3_U3304 | ~new_P3_LT_563_U7;
  assign new_P3_LT_563_U27 = ~new_P3_LT_563_U24 | ~new_P3_LT_563_U25 | ~new_P3_LT_563_U26;
  assign new_P3_LT_563_U28 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_LT_563_U14;
  assign new_P3_ADD_339_U4 = ~P3_PHYADDRPOINTER_REG_1_;
  assign new_P3_ADD_339_U5 = ~P3_PHYADDRPOINTER_REG_2_;
  assign new_P3_ADD_339_U6 = ~P3_PHYADDRPOINTER_REG_2_ | ~P3_PHYADDRPOINTER_REG_1_;
  assign new_P3_ADD_339_U7 = ~P3_PHYADDRPOINTER_REG_3_;
  assign new_P3_ADD_339_U8 = ~P3_PHYADDRPOINTER_REG_3_ | ~new_P3_ADD_339_U94;
  assign new_P3_ADD_339_U9 = ~P3_PHYADDRPOINTER_REG_4_;
  assign new_P3_ADD_339_U10 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_ADD_339_U95;
  assign new_P3_ADD_339_U11 = ~P3_PHYADDRPOINTER_REG_5_;
  assign new_P3_ADD_339_U12 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_ADD_339_U96;
  assign new_P3_ADD_339_U13 = ~P3_PHYADDRPOINTER_REG_6_;
  assign new_P3_ADD_339_U14 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_ADD_339_U97;
  assign new_P3_ADD_339_U15 = ~P3_PHYADDRPOINTER_REG_7_;
  assign new_P3_ADD_339_U16 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_ADD_339_U98;
  assign new_P3_ADD_339_U17 = ~P3_PHYADDRPOINTER_REG_8_;
  assign new_P3_ADD_339_U18 = ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_ADD_339_U19 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_ADD_339_U99;
  assign new_P3_ADD_339_U20 = ~new_P3_ADD_339_U100 | ~P3_PHYADDRPOINTER_REG_9_;
  assign new_P3_ADD_339_U21 = ~P3_PHYADDRPOINTER_REG_10_;
  assign new_P3_ADD_339_U22 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_ADD_339_U101;
  assign new_P3_ADD_339_U23 = ~P3_PHYADDRPOINTER_REG_11_;
  assign new_P3_ADD_339_U24 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_ADD_339_U102;
  assign new_P3_ADD_339_U25 = ~P3_PHYADDRPOINTER_REG_12_;
  assign new_P3_ADD_339_U26 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_ADD_339_U103;
  assign new_P3_ADD_339_U27 = ~P3_PHYADDRPOINTER_REG_13_;
  assign new_P3_ADD_339_U28 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_ADD_339_U104;
  assign new_P3_ADD_339_U29 = ~P3_PHYADDRPOINTER_REG_14_;
  assign new_P3_ADD_339_U30 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_ADD_339_U105;
  assign new_P3_ADD_339_U31 = ~P3_PHYADDRPOINTER_REG_15_;
  assign new_P3_ADD_339_U32 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_ADD_339_U106;
  assign new_P3_ADD_339_U33 = ~P3_PHYADDRPOINTER_REG_16_;
  assign new_P3_ADD_339_U34 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_ADD_339_U107;
  assign new_P3_ADD_339_U35 = ~P3_PHYADDRPOINTER_REG_17_;
  assign new_P3_ADD_339_U36 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_ADD_339_U108;
  assign new_P3_ADD_339_U37 = ~P3_PHYADDRPOINTER_REG_18_;
  assign new_P3_ADD_339_U38 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_ADD_339_U109;
  assign new_P3_ADD_339_U39 = ~P3_PHYADDRPOINTER_REG_19_;
  assign new_P3_ADD_339_U40 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_ADD_339_U110;
  assign new_P3_ADD_339_U41 = ~P3_PHYADDRPOINTER_REG_20_;
  assign new_P3_ADD_339_U42 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_ADD_339_U111;
  assign new_P3_ADD_339_U43 = ~P3_PHYADDRPOINTER_REG_21_;
  assign new_P3_ADD_339_U44 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_ADD_339_U112;
  assign new_P3_ADD_339_U45 = ~P3_PHYADDRPOINTER_REG_22_;
  assign new_P3_ADD_339_U46 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_ADD_339_U113;
  assign new_P3_ADD_339_U47 = ~P3_PHYADDRPOINTER_REG_23_;
  assign new_P3_ADD_339_U48 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_ADD_339_U114;
  assign new_P3_ADD_339_U49 = ~P3_PHYADDRPOINTER_REG_24_;
  assign new_P3_ADD_339_U50 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_ADD_339_U115;
  assign new_P3_ADD_339_U51 = ~P3_PHYADDRPOINTER_REG_25_;
  assign new_P3_ADD_339_U52 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_ADD_339_U116;
  assign new_P3_ADD_339_U53 = ~P3_PHYADDRPOINTER_REG_26_;
  assign new_P3_ADD_339_U54 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_ADD_339_U117;
  assign new_P3_ADD_339_U55 = ~P3_PHYADDRPOINTER_REG_27_;
  assign new_P3_ADD_339_U56 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_ADD_339_U118;
  assign new_P3_ADD_339_U57 = ~P3_PHYADDRPOINTER_REG_28_;
  assign new_P3_ADD_339_U58 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_ADD_339_U119;
  assign new_P3_ADD_339_U59 = ~P3_PHYADDRPOINTER_REG_29_;
  assign new_P3_ADD_339_U60 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_ADD_339_U120;
  assign new_P3_ADD_339_U61 = ~P3_PHYADDRPOINTER_REG_30_;
  assign new_P3_ADD_339_U62 = ~new_P3_ADD_339_U124 | ~new_P3_ADD_339_U123;
  assign new_P3_ADD_339_U63 = ~new_P3_ADD_339_U126 | ~new_P3_ADD_339_U125;
  assign new_P3_ADD_339_U64 = ~new_P3_ADD_339_U128 | ~new_P3_ADD_339_U127;
  assign new_P3_ADD_339_U65 = ~new_P3_ADD_339_U130 | ~new_P3_ADD_339_U129;
  assign new_P3_ADD_339_U66 = ~new_P3_ADD_339_U132 | ~new_P3_ADD_339_U131;
  assign new_P3_ADD_339_U67 = ~new_P3_ADD_339_U134 | ~new_P3_ADD_339_U133;
  assign new_P3_ADD_339_U68 = ~new_P3_ADD_339_U136 | ~new_P3_ADD_339_U135;
  assign new_P3_ADD_339_U69 = ~new_P3_ADD_339_U138 | ~new_P3_ADD_339_U137;
  assign new_P3_ADD_339_U70 = ~new_P3_ADD_339_U140 | ~new_P3_ADD_339_U139;
  assign new_P3_ADD_339_U71 = ~new_P3_ADD_339_U142 | ~new_P3_ADD_339_U141;
  assign new_P3_ADD_339_U72 = ~new_P3_ADD_339_U144 | ~new_P3_ADD_339_U143;
  assign new_P3_ADD_339_U73 = ~new_P3_ADD_339_U146 | ~new_P3_ADD_339_U145;
  assign new_P3_ADD_339_U74 = ~new_P3_ADD_339_U148 | ~new_P3_ADD_339_U147;
  assign new_P3_ADD_339_U75 = ~new_P3_ADD_339_U150 | ~new_P3_ADD_339_U149;
  assign new_P3_ADD_339_U76 = ~new_P3_ADD_339_U152 | ~new_P3_ADD_339_U151;
  assign new_P3_ADD_339_U77 = ~new_P3_ADD_339_U154 | ~new_P3_ADD_339_U153;
  assign new_P3_ADD_339_U78 = ~new_P3_ADD_339_U156 | ~new_P3_ADD_339_U155;
  assign new_P3_ADD_339_U79 = ~new_P3_ADD_339_U158 | ~new_P3_ADD_339_U157;
  assign new_P3_ADD_339_U80 = ~new_P3_ADD_339_U160 | ~new_P3_ADD_339_U159;
  assign new_P3_ADD_339_U81 = ~new_P3_ADD_339_U162 | ~new_P3_ADD_339_U161;
  assign new_P3_ADD_339_U82 = ~new_P3_ADD_339_U164 | ~new_P3_ADD_339_U163;
  assign new_P3_ADD_339_U83 = ~new_P3_ADD_339_U166 | ~new_P3_ADD_339_U165;
  assign new_P3_ADD_339_U84 = ~new_P3_ADD_339_U168 | ~new_P3_ADD_339_U167;
  assign new_P3_ADD_339_U85 = ~new_P3_ADD_339_U170 | ~new_P3_ADD_339_U169;
  assign new_P3_ADD_339_U86 = ~new_P3_ADD_339_U172 | ~new_P3_ADD_339_U171;
  assign new_P3_ADD_339_U87 = ~new_P3_ADD_339_U174 | ~new_P3_ADD_339_U173;
  assign new_P3_ADD_339_U88 = ~new_P3_ADD_339_U176 | ~new_P3_ADD_339_U175;
  assign new_P3_ADD_339_U89 = ~new_P3_ADD_339_U178 | ~new_P3_ADD_339_U177;
  assign new_P3_ADD_339_U90 = ~new_P3_ADD_339_U180 | ~new_P3_ADD_339_U179;
  assign new_P3_ADD_339_U91 = ~new_P3_ADD_339_U182 | ~new_P3_ADD_339_U181;
  assign new_P3_ADD_339_U92 = ~P3_PHYADDRPOINTER_REG_31_;
  assign new_P3_ADD_339_U93 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_ADD_339_U121;
  assign new_P3_ADD_339_U94 = ~new_P3_ADD_339_U6;
  assign new_P3_ADD_339_U95 = ~new_P3_ADD_339_U8;
  assign new_P3_ADD_339_U96 = ~new_P3_ADD_339_U10;
  assign new_P3_ADD_339_U97 = ~new_P3_ADD_339_U12;
  assign new_P3_ADD_339_U98 = ~new_P3_ADD_339_U14;
  assign new_P3_ADD_339_U99 = ~new_P3_ADD_339_U16;
  assign new_P3_ADD_339_U100 = ~new_P3_ADD_339_U19;
  assign new_P3_ADD_339_U101 = ~new_P3_ADD_339_U20;
  assign new_P3_ADD_339_U102 = ~new_P3_ADD_339_U22;
  assign new_P3_ADD_339_U103 = ~new_P3_ADD_339_U24;
  assign new_P3_ADD_339_U104 = ~new_P3_ADD_339_U26;
  assign new_P3_ADD_339_U105 = ~new_P3_ADD_339_U28;
  assign new_P3_ADD_339_U106 = ~new_P3_ADD_339_U30;
  assign new_P3_ADD_339_U107 = ~new_P3_ADD_339_U32;
  assign new_P3_ADD_339_U108 = ~new_P3_ADD_339_U34;
  assign new_P3_ADD_339_U109 = ~new_P3_ADD_339_U36;
  assign new_P3_ADD_339_U110 = ~new_P3_ADD_339_U38;
  assign new_P3_ADD_339_U111 = ~new_P3_ADD_339_U40;
  assign new_P3_ADD_339_U112 = ~new_P3_ADD_339_U42;
  assign new_P3_ADD_339_U113 = ~new_P3_ADD_339_U44;
  assign new_P3_ADD_339_U114 = ~new_P3_ADD_339_U46;
  assign new_P3_ADD_339_U115 = ~new_P3_ADD_339_U48;
  assign new_P3_ADD_339_U116 = ~new_P3_ADD_339_U50;
  assign new_P3_ADD_339_U117 = ~new_P3_ADD_339_U52;
  assign new_P3_ADD_339_U118 = ~new_P3_ADD_339_U54;
  assign new_P3_ADD_339_U119 = ~new_P3_ADD_339_U56;
  assign new_P3_ADD_339_U120 = ~new_P3_ADD_339_U58;
  assign new_P3_ADD_339_U121 = ~new_P3_ADD_339_U60;
  assign new_P3_ADD_339_U122 = ~new_P3_ADD_339_U93;
  assign new_P3_ADD_339_U123 = ~P3_PHYADDRPOINTER_REG_9_ | ~new_P3_ADD_339_U19;
  assign new_P3_ADD_339_U124 = ~new_P3_ADD_339_U100 | ~new_P3_ADD_339_U18;
  assign new_P3_ADD_339_U125 = ~P3_PHYADDRPOINTER_REG_8_ | ~new_P3_ADD_339_U16;
  assign new_P3_ADD_339_U126 = ~new_P3_ADD_339_U99 | ~new_P3_ADD_339_U17;
  assign new_P3_ADD_339_U127 = ~P3_PHYADDRPOINTER_REG_7_ | ~new_P3_ADD_339_U14;
  assign new_P3_ADD_339_U128 = ~new_P3_ADD_339_U98 | ~new_P3_ADD_339_U15;
  assign new_P3_ADD_339_U129 = ~P3_PHYADDRPOINTER_REG_6_ | ~new_P3_ADD_339_U12;
  assign new_P3_ADD_339_U130 = ~new_P3_ADD_339_U97 | ~new_P3_ADD_339_U13;
  assign new_P3_ADD_339_U131 = ~P3_PHYADDRPOINTER_REG_5_ | ~new_P3_ADD_339_U10;
  assign new_P3_ADD_339_U132 = ~new_P3_ADD_339_U96 | ~new_P3_ADD_339_U11;
  assign new_P3_ADD_339_U133 = ~P3_PHYADDRPOINTER_REG_4_ | ~new_P3_ADD_339_U8;
  assign new_P3_ADD_339_U134 = ~new_P3_ADD_339_U95 | ~new_P3_ADD_339_U9;
  assign new_P3_ADD_339_U135 = ~P3_PHYADDRPOINTER_REG_3_ | ~new_P3_ADD_339_U6;
  assign new_P3_ADD_339_U136 = ~new_P3_ADD_339_U94 | ~new_P3_ADD_339_U7;
  assign new_P3_ADD_339_U137 = ~P3_PHYADDRPOINTER_REG_31_ | ~new_P3_ADD_339_U93;
  assign new_P3_ADD_339_U138 = ~new_P3_ADD_339_U122 | ~new_P3_ADD_339_U92;
  assign new_P3_ADD_339_U139 = ~P3_PHYADDRPOINTER_REG_30_ | ~new_P3_ADD_339_U60;
  assign new_P3_ADD_339_U140 = ~new_P3_ADD_339_U121 | ~new_P3_ADD_339_U61;
  assign new_P3_ADD_339_U141 = ~P3_PHYADDRPOINTER_REG_2_ | ~new_P3_ADD_339_U4;
  assign new_P3_ADD_339_U142 = ~P3_PHYADDRPOINTER_REG_1_ | ~new_P3_ADD_339_U5;
  assign new_P3_ADD_339_U143 = ~P3_PHYADDRPOINTER_REG_29_ | ~new_P3_ADD_339_U58;
  assign new_P3_ADD_339_U144 = ~new_P3_ADD_339_U120 | ~new_P3_ADD_339_U59;
  assign new_P3_ADD_339_U145 = ~P3_PHYADDRPOINTER_REG_28_ | ~new_P3_ADD_339_U56;
  assign new_P3_ADD_339_U146 = ~new_P3_ADD_339_U119 | ~new_P3_ADD_339_U57;
  assign new_P3_ADD_339_U147 = ~P3_PHYADDRPOINTER_REG_27_ | ~new_P3_ADD_339_U54;
  assign new_P3_ADD_339_U148 = ~new_P3_ADD_339_U118 | ~new_P3_ADD_339_U55;
  assign new_P3_ADD_339_U149 = ~P3_PHYADDRPOINTER_REG_26_ | ~new_P3_ADD_339_U52;
  assign new_P3_ADD_339_U150 = ~new_P3_ADD_339_U117 | ~new_P3_ADD_339_U53;
  assign new_P3_ADD_339_U151 = ~P3_PHYADDRPOINTER_REG_25_ | ~new_P3_ADD_339_U50;
  assign new_P3_ADD_339_U152 = ~new_P3_ADD_339_U116 | ~new_P3_ADD_339_U51;
  assign new_P3_ADD_339_U153 = ~P3_PHYADDRPOINTER_REG_24_ | ~new_P3_ADD_339_U48;
  assign new_P3_ADD_339_U154 = ~new_P3_ADD_339_U115 | ~new_P3_ADD_339_U49;
  assign new_P3_ADD_339_U155 = ~P3_PHYADDRPOINTER_REG_23_ | ~new_P3_ADD_339_U46;
  assign new_P3_ADD_339_U156 = ~new_P3_ADD_339_U114 | ~new_P3_ADD_339_U47;
  assign new_P3_ADD_339_U157 = ~P3_PHYADDRPOINTER_REG_22_ | ~new_P3_ADD_339_U44;
  assign new_P3_ADD_339_U158 = ~new_P3_ADD_339_U113 | ~new_P3_ADD_339_U45;
  assign new_P3_ADD_339_U159 = ~P3_PHYADDRPOINTER_REG_21_ | ~new_P3_ADD_339_U42;
  assign new_P3_ADD_339_U160 = ~new_P3_ADD_339_U112 | ~new_P3_ADD_339_U43;
  assign new_P3_ADD_339_U161 = ~P3_PHYADDRPOINTER_REG_20_ | ~new_P3_ADD_339_U40;
  assign new_P3_ADD_339_U162 = ~new_P3_ADD_339_U111 | ~new_P3_ADD_339_U41;
  assign new_P3_ADD_339_U163 = ~P3_PHYADDRPOINTER_REG_19_ | ~new_P3_ADD_339_U38;
  assign new_P3_ADD_339_U164 = ~new_P3_ADD_339_U110 | ~new_P3_ADD_339_U39;
  assign new_P3_ADD_339_U165 = ~P3_PHYADDRPOINTER_REG_18_ | ~new_P3_ADD_339_U36;
  assign new_P3_ADD_339_U166 = ~new_P3_ADD_339_U109 | ~new_P3_ADD_339_U37;
  assign new_P3_ADD_339_U167 = ~P3_PHYADDRPOINTER_REG_17_ | ~new_P3_ADD_339_U34;
  assign new_P3_ADD_339_U168 = ~new_P3_ADD_339_U108 | ~new_P3_ADD_339_U35;
  assign new_P3_ADD_339_U169 = ~P3_PHYADDRPOINTER_REG_16_ | ~new_P3_ADD_339_U32;
  assign new_P3_ADD_339_U170 = ~new_P3_ADD_339_U107 | ~new_P3_ADD_339_U33;
  assign new_P3_ADD_339_U171 = ~P3_PHYADDRPOINTER_REG_15_ | ~new_P3_ADD_339_U30;
  assign new_P3_ADD_339_U172 = ~new_P3_ADD_339_U106 | ~new_P3_ADD_339_U31;
  assign new_P3_ADD_339_U173 = ~P3_PHYADDRPOINTER_REG_14_ | ~new_P3_ADD_339_U28;
  assign new_P3_ADD_339_U174 = ~new_P3_ADD_339_U105 | ~new_P3_ADD_339_U29;
  assign new_P3_ADD_339_U175 = ~P3_PHYADDRPOINTER_REG_13_ | ~new_P3_ADD_339_U26;
  assign new_P3_ADD_339_U176 = ~new_P3_ADD_339_U104 | ~new_P3_ADD_339_U27;
  assign new_P3_ADD_339_U177 = ~P3_PHYADDRPOINTER_REG_12_ | ~new_P3_ADD_339_U24;
  assign new_P3_ADD_339_U178 = ~new_P3_ADD_339_U103 | ~new_P3_ADD_339_U25;
  assign new_P3_ADD_339_U179 = ~P3_PHYADDRPOINTER_REG_11_ | ~new_P3_ADD_339_U22;
  assign new_P3_ADD_339_U180 = ~new_P3_ADD_339_U102 | ~new_P3_ADD_339_U23;
  assign new_P3_ADD_339_U181 = ~P3_PHYADDRPOINTER_REG_10_ | ~new_P3_ADD_339_U20;
  assign new_P3_ADD_339_U182 = ~new_P3_ADD_339_U101 | ~new_P3_ADD_339_U21;
  assign new_P3_ADD_360_U4 = ~new_P3_U2622;
  assign new_P3_ADD_360_U5 = new_P3_ADD_360_U22 & new_P3_ADD_360_U27;
  assign new_P3_ADD_360_U6 = ~new_P3_U2623;
  assign new_P3_ADD_360_U7 = ~new_P3_U2623 | ~new_P3_U2622;
  assign new_P3_ADD_360_U8 = ~new_P3_U2624;
  assign new_P3_ADD_360_U9 = ~new_P3_U2624 | ~new_P3_ADD_360_U24;
  assign new_P3_ADD_360_U10 = ~new_P3_U2625;
  assign new_P3_ADD_360_U11 = ~new_P3_U2625 | ~new_P3_ADD_360_U25;
  assign new_P3_ADD_360_U12 = ~new_P3_U2626;
  assign new_P3_ADD_360_U13 = ~new_P3_U2626 | ~new_P3_ADD_360_U26;
  assign new_P3_ADD_360_U14 = ~new_P3_U2628;
  assign new_P3_ADD_360_U15 = ~new_P3_U2627;
  assign new_P3_ADD_360_U16 = ~new_P3_ADD_360_U30 | ~new_P3_ADD_360_U29;
  assign new_P3_ADD_360_U17 = ~new_P3_ADD_360_U32 | ~new_P3_ADD_360_U31;
  assign new_P3_ADD_360_U18 = ~new_P3_ADD_360_U34 | ~new_P3_ADD_360_U33;
  assign new_P3_ADD_360_U19 = ~new_P3_ADD_360_U36 | ~new_P3_ADD_360_U35;
  assign new_P3_ADD_360_U20 = ~new_P3_ADD_360_U38 | ~new_P3_ADD_360_U37;
  assign new_P3_ADD_360_U21 = ~new_P3_ADD_360_U40 | ~new_P3_ADD_360_U39;
  assign new_P3_ADD_360_U22 = new_P3_U2628 & new_P3_U2627;
  assign new_P3_ADD_360_U23 = ~new_P3_U2627 | ~new_P3_ADD_360_U27;
  assign new_P3_ADD_360_U24 = ~new_P3_ADD_360_U7;
  assign new_P3_ADD_360_U25 = ~new_P3_ADD_360_U9;
  assign new_P3_ADD_360_U26 = ~new_P3_ADD_360_U11;
  assign new_P3_ADD_360_U27 = ~new_P3_ADD_360_U13;
  assign new_P3_ADD_360_U28 = ~new_P3_ADD_360_U23;
  assign new_P3_ADD_360_U29 = ~new_P3_U2628 | ~new_P3_ADD_360_U23;
  assign new_P3_ADD_360_U30 = ~new_P3_ADD_360_U28 | ~new_P3_ADD_360_U14;
  assign new_P3_ADD_360_U31 = ~new_P3_U2627 | ~new_P3_ADD_360_U13;
  assign new_P3_ADD_360_U32 = ~new_P3_ADD_360_U27 | ~new_P3_ADD_360_U15;
  assign new_P3_ADD_360_U33 = ~new_P3_U2626 | ~new_P3_ADD_360_U11;
  assign new_P3_ADD_360_U34 = ~new_P3_ADD_360_U26 | ~new_P3_ADD_360_U12;
  assign new_P3_ADD_360_U35 = ~new_P3_U2625 | ~new_P3_ADD_360_U9;
  assign new_P3_ADD_360_U36 = ~new_P3_ADD_360_U25 | ~new_P3_ADD_360_U10;
  assign new_P3_ADD_360_U37 = ~new_P3_U2624 | ~new_P3_ADD_360_U7;
  assign new_P3_ADD_360_U38 = ~new_P3_ADD_360_U24 | ~new_P3_ADD_360_U8;
  assign new_P3_ADD_360_U39 = ~new_P3_U2623 | ~new_P3_ADD_360_U4;
  assign new_P3_ADD_360_U40 = ~new_P3_U2622 | ~new_P3_ADD_360_U6;
  assign new_P3_LTE_597_U6 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_580_U6 = ~new_P3_SUB_580_U10 | ~new_P3_SUB_580_U9;
  assign new_P3_SUB_580_U7 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_SUB_580_U8 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_SUB_580_U9 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_SUB_580_U8;
  assign new_P3_SUB_580_U10 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_SUB_580_U7;
  assign new_P3_LT_589_U6 = new_P3_LT_589_U8 | new_P3_U2629;
  assign new_P3_LT_589_U7 = new_P3_SUB_589_U7 & new_P3_SUB_589_U6;
  assign new_P3_LT_589_U8 = ~new_P3_SUB_589_U9 & ~new_P3_LT_589_U7 & ~new_P3_SUB_589_U8;
  assign new_P3_ADD_541_U4 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_541_U5 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_541_U6 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_541_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_541_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_541_U94;
  assign new_P3_ADD_541_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_541_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_541_U95;
  assign new_P3_ADD_541_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_541_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_541_U96;
  assign new_P3_ADD_541_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_541_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_541_U97;
  assign new_P3_ADD_541_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_541_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_541_U98;
  assign new_P3_ADD_541_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_541_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_541_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_541_U99;
  assign new_P3_ADD_541_U20 = ~new_P3_ADD_541_U100 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_541_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_541_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_541_U101;
  assign new_P3_ADD_541_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_541_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_541_U102;
  assign new_P3_ADD_541_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_541_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_541_U103;
  assign new_P3_ADD_541_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_541_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_541_U104;
  assign new_P3_ADD_541_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_541_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_541_U105;
  assign new_P3_ADD_541_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_541_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_541_U106;
  assign new_P3_ADD_541_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_541_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_541_U107;
  assign new_P3_ADD_541_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_541_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_541_U108;
  assign new_P3_ADD_541_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_541_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_541_U109;
  assign new_P3_ADD_541_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_541_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_541_U110;
  assign new_P3_ADD_541_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_541_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_541_U111;
  assign new_P3_ADD_541_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_541_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_541_U112;
  assign new_P3_ADD_541_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_541_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_541_U113;
  assign new_P3_ADD_541_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_541_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_541_U114;
  assign new_P3_ADD_541_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_541_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_541_U115;
  assign new_P3_ADD_541_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_541_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_541_U116;
  assign new_P3_ADD_541_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_541_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_541_U117;
  assign new_P3_ADD_541_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_541_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_541_U118;
  assign new_P3_ADD_541_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_541_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_541_U119;
  assign new_P3_ADD_541_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_541_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_541_U120;
  assign new_P3_ADD_541_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_541_U62 = ~new_P3_ADD_541_U124 | ~new_P3_ADD_541_U123;
  assign new_P3_ADD_541_U63 = ~new_P3_ADD_541_U126 | ~new_P3_ADD_541_U125;
  assign new_P3_ADD_541_U64 = ~new_P3_ADD_541_U128 | ~new_P3_ADD_541_U127;
  assign new_P3_ADD_541_U65 = ~new_P3_ADD_541_U130 | ~new_P3_ADD_541_U129;
  assign new_P3_ADD_541_U66 = ~new_P3_ADD_541_U132 | ~new_P3_ADD_541_U131;
  assign new_P3_ADD_541_U67 = ~new_P3_ADD_541_U134 | ~new_P3_ADD_541_U133;
  assign new_P3_ADD_541_U68 = ~new_P3_ADD_541_U136 | ~new_P3_ADD_541_U135;
  assign new_P3_ADD_541_U69 = ~new_P3_ADD_541_U138 | ~new_P3_ADD_541_U137;
  assign new_P3_ADD_541_U70 = ~new_P3_ADD_541_U140 | ~new_P3_ADD_541_U139;
  assign new_P3_ADD_541_U71 = ~new_P3_ADD_541_U142 | ~new_P3_ADD_541_U141;
  assign new_P3_ADD_541_U72 = ~new_P3_ADD_541_U144 | ~new_P3_ADD_541_U143;
  assign new_P3_ADD_541_U73 = ~new_P3_ADD_541_U146 | ~new_P3_ADD_541_U145;
  assign new_P3_ADD_541_U74 = ~new_P3_ADD_541_U148 | ~new_P3_ADD_541_U147;
  assign new_P3_ADD_541_U75 = ~new_P3_ADD_541_U150 | ~new_P3_ADD_541_U149;
  assign new_P3_ADD_541_U76 = ~new_P3_ADD_541_U152 | ~new_P3_ADD_541_U151;
  assign new_P3_ADD_541_U77 = ~new_P3_ADD_541_U154 | ~new_P3_ADD_541_U153;
  assign new_P3_ADD_541_U78 = ~new_P3_ADD_541_U156 | ~new_P3_ADD_541_U155;
  assign new_P3_ADD_541_U79 = ~new_P3_ADD_541_U158 | ~new_P3_ADD_541_U157;
  assign new_P3_ADD_541_U80 = ~new_P3_ADD_541_U160 | ~new_P3_ADD_541_U159;
  assign new_P3_ADD_541_U81 = ~new_P3_ADD_541_U162 | ~new_P3_ADD_541_U161;
  assign new_P3_ADD_541_U82 = ~new_P3_ADD_541_U164 | ~new_P3_ADD_541_U163;
  assign new_P3_ADD_541_U83 = ~new_P3_ADD_541_U166 | ~new_P3_ADD_541_U165;
  assign new_P3_ADD_541_U84 = ~new_P3_ADD_541_U168 | ~new_P3_ADD_541_U167;
  assign new_P3_ADD_541_U85 = ~new_P3_ADD_541_U170 | ~new_P3_ADD_541_U169;
  assign new_P3_ADD_541_U86 = ~new_P3_ADD_541_U172 | ~new_P3_ADD_541_U171;
  assign new_P3_ADD_541_U87 = ~new_P3_ADD_541_U174 | ~new_P3_ADD_541_U173;
  assign new_P3_ADD_541_U88 = ~new_P3_ADD_541_U176 | ~new_P3_ADD_541_U175;
  assign new_P3_ADD_541_U89 = ~new_P3_ADD_541_U178 | ~new_P3_ADD_541_U177;
  assign new_P3_ADD_541_U90 = ~new_P3_ADD_541_U180 | ~new_P3_ADD_541_U179;
  assign new_P3_ADD_541_U91 = ~new_P3_ADD_541_U182 | ~new_P3_ADD_541_U181;
  assign new_P3_ADD_541_U92 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_541_U93 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_541_U121;
  assign new_P3_ADD_541_U94 = ~new_P3_ADD_541_U6;
  assign new_P3_ADD_541_U95 = ~new_P3_ADD_541_U8;
  assign new_P3_ADD_541_U96 = ~new_P3_ADD_541_U10;
  assign new_P3_ADD_541_U97 = ~new_P3_ADD_541_U12;
  assign new_P3_ADD_541_U98 = ~new_P3_ADD_541_U14;
  assign new_P3_ADD_541_U99 = ~new_P3_ADD_541_U16;
  assign new_P3_ADD_541_U100 = ~new_P3_ADD_541_U19;
  assign new_P3_ADD_541_U101 = ~new_P3_ADD_541_U20;
  assign new_P3_ADD_541_U102 = ~new_P3_ADD_541_U22;
  assign new_P3_ADD_541_U103 = ~new_P3_ADD_541_U24;
  assign new_P3_ADD_541_U104 = ~new_P3_ADD_541_U26;
  assign new_P3_ADD_541_U105 = ~new_P3_ADD_541_U28;
  assign new_P3_ADD_541_U106 = ~new_P3_ADD_541_U30;
  assign new_P3_ADD_541_U107 = ~new_P3_ADD_541_U32;
  assign new_P3_ADD_541_U108 = ~new_P3_ADD_541_U34;
  assign new_P3_ADD_541_U109 = ~new_P3_ADD_541_U36;
  assign new_P3_ADD_541_U110 = ~new_P3_ADD_541_U38;
  assign new_P3_ADD_541_U111 = ~new_P3_ADD_541_U40;
  assign new_P3_ADD_541_U112 = ~new_P3_ADD_541_U42;
  assign new_P3_ADD_541_U113 = ~new_P3_ADD_541_U44;
  assign new_P3_ADD_541_U114 = ~new_P3_ADD_541_U46;
  assign new_P3_ADD_541_U115 = ~new_P3_ADD_541_U48;
  assign new_P3_ADD_541_U116 = ~new_P3_ADD_541_U50;
  assign new_P3_ADD_541_U117 = ~new_P3_ADD_541_U52;
  assign new_P3_ADD_541_U118 = ~new_P3_ADD_541_U54;
  assign new_P3_ADD_541_U119 = ~new_P3_ADD_541_U56;
  assign new_P3_ADD_541_U120 = ~new_P3_ADD_541_U58;
  assign new_P3_ADD_541_U121 = ~new_P3_ADD_541_U60;
  assign new_P3_ADD_541_U122 = ~new_P3_ADD_541_U93;
  assign new_P3_ADD_541_U123 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_541_U19;
  assign new_P3_ADD_541_U124 = ~new_P3_ADD_541_U100 | ~new_P3_ADD_541_U18;
  assign new_P3_ADD_541_U125 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_541_U16;
  assign new_P3_ADD_541_U126 = ~new_P3_ADD_541_U99 | ~new_P3_ADD_541_U17;
  assign new_P3_ADD_541_U127 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_541_U14;
  assign new_P3_ADD_541_U128 = ~new_P3_ADD_541_U98 | ~new_P3_ADD_541_U15;
  assign new_P3_ADD_541_U129 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_541_U12;
  assign new_P3_ADD_541_U130 = ~new_P3_ADD_541_U97 | ~new_P3_ADD_541_U13;
  assign new_P3_ADD_541_U131 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_541_U10;
  assign new_P3_ADD_541_U132 = ~new_P3_ADD_541_U96 | ~new_P3_ADD_541_U11;
  assign new_P3_ADD_541_U133 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_541_U8;
  assign new_P3_ADD_541_U134 = ~new_P3_ADD_541_U95 | ~new_P3_ADD_541_U9;
  assign new_P3_ADD_541_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_541_U6;
  assign new_P3_ADD_541_U136 = ~new_P3_ADD_541_U94 | ~new_P3_ADD_541_U7;
  assign new_P3_ADD_541_U137 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_541_U93;
  assign new_P3_ADD_541_U138 = ~new_P3_ADD_541_U122 | ~new_P3_ADD_541_U92;
  assign new_P3_ADD_541_U139 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_541_U60;
  assign new_P3_ADD_541_U140 = ~new_P3_ADD_541_U121 | ~new_P3_ADD_541_U61;
  assign new_P3_ADD_541_U141 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_541_U4;
  assign new_P3_ADD_541_U142 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_541_U5;
  assign new_P3_ADD_541_U143 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_541_U58;
  assign new_P3_ADD_541_U144 = ~new_P3_ADD_541_U120 | ~new_P3_ADD_541_U59;
  assign new_P3_ADD_541_U145 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_541_U56;
  assign new_P3_ADD_541_U146 = ~new_P3_ADD_541_U119 | ~new_P3_ADD_541_U57;
  assign new_P3_ADD_541_U147 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_541_U54;
  assign new_P3_ADD_541_U148 = ~new_P3_ADD_541_U118 | ~new_P3_ADD_541_U55;
  assign new_P3_ADD_541_U149 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_541_U52;
  assign new_P3_ADD_541_U150 = ~new_P3_ADD_541_U117 | ~new_P3_ADD_541_U53;
  assign new_P3_ADD_541_U151 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_541_U50;
  assign new_P3_ADD_541_U152 = ~new_P3_ADD_541_U116 | ~new_P3_ADD_541_U51;
  assign new_P3_ADD_541_U153 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_541_U48;
  assign new_P3_ADD_541_U154 = ~new_P3_ADD_541_U115 | ~new_P3_ADD_541_U49;
  assign new_P3_ADD_541_U155 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_541_U46;
  assign new_P3_ADD_541_U156 = ~new_P3_ADD_541_U114 | ~new_P3_ADD_541_U47;
  assign new_P3_ADD_541_U157 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_541_U44;
  assign new_P3_ADD_541_U158 = ~new_P3_ADD_541_U113 | ~new_P3_ADD_541_U45;
  assign new_P3_ADD_541_U159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_541_U42;
  assign new_P3_ADD_541_U160 = ~new_P3_ADD_541_U112 | ~new_P3_ADD_541_U43;
  assign new_P3_ADD_541_U161 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_541_U40;
  assign new_P3_ADD_541_U162 = ~new_P3_ADD_541_U111 | ~new_P3_ADD_541_U41;
  assign new_P3_ADD_541_U163 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_541_U38;
  assign new_P3_ADD_541_U164 = ~new_P3_ADD_541_U110 | ~new_P3_ADD_541_U39;
  assign new_P3_ADD_541_U165 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_541_U36;
  assign new_P3_ADD_541_U166 = ~new_P3_ADD_541_U109 | ~new_P3_ADD_541_U37;
  assign new_P3_ADD_541_U167 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_541_U34;
  assign new_P3_ADD_541_U168 = ~new_P3_ADD_541_U108 | ~new_P3_ADD_541_U35;
  assign new_P3_ADD_541_U169 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_541_U32;
  assign new_P3_ADD_541_U170 = ~new_P3_ADD_541_U107 | ~new_P3_ADD_541_U33;
  assign new_P3_ADD_541_U171 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_541_U30;
  assign new_P3_ADD_541_U172 = ~new_P3_ADD_541_U106 | ~new_P3_ADD_541_U31;
  assign new_P3_ADD_541_U173 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_541_U28;
  assign new_P3_ADD_541_U174 = ~new_P3_ADD_541_U105 | ~new_P3_ADD_541_U29;
  assign new_P3_ADD_541_U175 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_541_U26;
  assign new_P3_ADD_541_U176 = ~new_P3_ADD_541_U104 | ~new_P3_ADD_541_U27;
  assign new_P3_ADD_541_U177 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_541_U24;
  assign new_P3_ADD_541_U178 = ~new_P3_ADD_541_U103 | ~new_P3_ADD_541_U25;
  assign new_P3_ADD_541_U179 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_541_U22;
  assign new_P3_ADD_541_U180 = ~new_P3_ADD_541_U102 | ~new_P3_ADD_541_U23;
  assign new_P3_ADD_541_U181 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_541_U20;
  assign new_P3_ADD_541_U182 = ~new_P3_ADD_541_U101 | ~new_P3_ADD_541_U21;
  assign new_P3_SUB_355_U6 = ~new_P3_SUB_355_U45 | ~new_P3_SUB_355_U44;
  assign new_P3_SUB_355_U7 = ~new_P3_SUB_355_U9 | ~new_P3_SUB_355_U46;
  assign new_P3_SUB_355_U8 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_SUB_355_U9 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_355_U18;
  assign new_P3_SUB_355_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_355_U11 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_355_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_355_U13 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_355_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_355_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_355_U16 = ~new_P3_SUB_355_U41 | ~new_P3_SUB_355_U40;
  assign new_P3_SUB_355_U17 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_355_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_355_U19 = ~new_P3_SUB_355_U51 | ~new_P3_SUB_355_U50;
  assign new_P3_SUB_355_U20 = ~new_P3_SUB_355_U56 | ~new_P3_SUB_355_U55;
  assign new_P3_SUB_355_U21 = ~new_P3_SUB_355_U61 | ~new_P3_SUB_355_U60;
  assign new_P3_SUB_355_U22 = ~new_P3_SUB_355_U66 | ~new_P3_SUB_355_U65;
  assign new_P3_SUB_355_U23 = ~new_P3_SUB_355_U48 | ~new_P3_SUB_355_U47;
  assign new_P3_SUB_355_U24 = ~new_P3_SUB_355_U53 | ~new_P3_SUB_355_U52;
  assign new_P3_SUB_355_U25 = ~new_P3_SUB_355_U58 | ~new_P3_SUB_355_U57;
  assign new_P3_SUB_355_U26 = ~new_P3_SUB_355_U63 | ~new_P3_SUB_355_U62;
  assign new_P3_SUB_355_U27 = ~new_P3_SUB_355_U37 | ~new_P3_SUB_355_U36;
  assign new_P3_SUB_355_U28 = ~new_P3_SUB_355_U33 | ~new_P3_SUB_355_U32;
  assign new_P3_SUB_355_U29 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_355_U30 = ~new_P3_SUB_355_U9;
  assign new_P3_SUB_355_U31 = ~new_P3_SUB_355_U30 | ~new_P3_SUB_355_U10;
  assign new_P3_SUB_355_U32 = ~new_P3_SUB_355_U31 | ~new_P3_SUB_355_U29;
  assign new_P3_SUB_355_U33 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_355_U9;
  assign new_P3_SUB_355_U34 = ~new_P3_SUB_355_U28;
  assign new_P3_SUB_355_U35 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_355_U12;
  assign new_P3_SUB_355_U36 = ~new_P3_SUB_355_U35 | ~new_P3_SUB_355_U28;
  assign new_P3_SUB_355_U37 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_355_U11;
  assign new_P3_SUB_355_U38 = ~new_P3_SUB_355_U27;
  assign new_P3_SUB_355_U39 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_355_U14;
  assign new_P3_SUB_355_U40 = ~new_P3_SUB_355_U39 | ~new_P3_SUB_355_U27;
  assign new_P3_SUB_355_U41 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_355_U13;
  assign new_P3_SUB_355_U42 = ~new_P3_SUB_355_U16;
  assign new_P3_SUB_355_U43 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_355_U17;
  assign new_P3_SUB_355_U44 = ~new_P3_SUB_355_U42 | ~new_P3_SUB_355_U43;
  assign new_P3_SUB_355_U45 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_355_U15;
  assign new_P3_SUB_355_U46 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_SUB_355_U8;
  assign new_P3_SUB_355_U47 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_355_U15;
  assign new_P3_SUB_355_U48 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_355_U17;
  assign new_P3_SUB_355_U49 = ~new_P3_SUB_355_U23;
  assign new_P3_SUB_355_U50 = ~new_P3_SUB_355_U49 | ~new_P3_SUB_355_U42;
  assign new_P3_SUB_355_U51 = ~new_P3_SUB_355_U23 | ~new_P3_SUB_355_U16;
  assign new_P3_SUB_355_U52 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_355_U14;
  assign new_P3_SUB_355_U53 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_355_U13;
  assign new_P3_SUB_355_U54 = ~new_P3_SUB_355_U24;
  assign new_P3_SUB_355_U55 = ~new_P3_SUB_355_U38 | ~new_P3_SUB_355_U54;
  assign new_P3_SUB_355_U56 = ~new_P3_SUB_355_U24 | ~new_P3_SUB_355_U27;
  assign new_P3_SUB_355_U57 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_355_U12;
  assign new_P3_SUB_355_U58 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_355_U11;
  assign new_P3_SUB_355_U59 = ~new_P3_SUB_355_U25;
  assign new_P3_SUB_355_U60 = ~new_P3_SUB_355_U34 | ~new_P3_SUB_355_U59;
  assign new_P3_SUB_355_U61 = ~new_P3_SUB_355_U25 | ~new_P3_SUB_355_U28;
  assign new_P3_SUB_355_U62 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_355_U10;
  assign new_P3_SUB_355_U63 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_355_U29;
  assign new_P3_SUB_355_U64 = ~new_P3_SUB_355_U26;
  assign new_P3_SUB_355_U65 = ~new_P3_SUB_355_U64 | ~new_P3_SUB_355_U30;
  assign new_P3_SUB_355_U66 = ~new_P3_SUB_355_U26 | ~new_P3_SUB_355_U9;
  assign new_P3_SUB_450_U6 = ~new_P3_SUB_450_U43 | ~new_P3_SUB_450_U42;
  assign new_P3_SUB_450_U7 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_450_U27;
  assign new_P3_SUB_450_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_450_U9 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_450_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_450_U11 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_450_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_450_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_450_U14 = ~new_P3_SUB_450_U39 | ~new_P3_SUB_450_U38;
  assign new_P3_SUB_450_U15 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_450_U16 = ~new_P3_SUB_450_U48 | ~new_P3_SUB_450_U47;
  assign new_P3_SUB_450_U17 = ~new_P3_SUB_450_U53 | ~new_P3_SUB_450_U52;
  assign new_P3_SUB_450_U18 = ~new_P3_SUB_450_U58 | ~new_P3_SUB_450_U57;
  assign new_P3_SUB_450_U19 = ~new_P3_SUB_450_U63 | ~new_P3_SUB_450_U62;
  assign new_P3_SUB_450_U20 = ~new_P3_SUB_450_U45 | ~new_P3_SUB_450_U44;
  assign new_P3_SUB_450_U21 = ~new_P3_SUB_450_U50 | ~new_P3_SUB_450_U49;
  assign new_P3_SUB_450_U22 = ~new_P3_SUB_450_U55 | ~new_P3_SUB_450_U54;
  assign new_P3_SUB_450_U23 = ~new_P3_SUB_450_U60 | ~new_P3_SUB_450_U59;
  assign new_P3_SUB_450_U24 = ~new_P3_SUB_450_U35 | ~new_P3_SUB_450_U34;
  assign new_P3_SUB_450_U25 = ~new_P3_SUB_450_U31 | ~new_P3_SUB_450_U30;
  assign new_P3_SUB_450_U26 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_450_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_450_U28 = ~new_P3_SUB_450_U7;
  assign new_P3_SUB_450_U29 = ~new_P3_SUB_450_U28 | ~new_P3_SUB_450_U8;
  assign new_P3_SUB_450_U30 = ~new_P3_SUB_450_U29 | ~new_P3_SUB_450_U26;
  assign new_P3_SUB_450_U31 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_450_U7;
  assign new_P3_SUB_450_U32 = ~new_P3_SUB_450_U25;
  assign new_P3_SUB_450_U33 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_450_U10;
  assign new_P3_SUB_450_U34 = ~new_P3_SUB_450_U33 | ~new_P3_SUB_450_U25;
  assign new_P3_SUB_450_U35 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_450_U9;
  assign new_P3_SUB_450_U36 = ~new_P3_SUB_450_U24;
  assign new_P3_SUB_450_U37 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_450_U12;
  assign new_P3_SUB_450_U38 = ~new_P3_SUB_450_U37 | ~new_P3_SUB_450_U24;
  assign new_P3_SUB_450_U39 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_450_U11;
  assign new_P3_SUB_450_U40 = ~new_P3_SUB_450_U14;
  assign new_P3_SUB_450_U41 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_450_U15;
  assign new_P3_SUB_450_U42 = ~new_P3_SUB_450_U40 | ~new_P3_SUB_450_U41;
  assign new_P3_SUB_450_U43 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_450_U13;
  assign new_P3_SUB_450_U44 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_450_U13;
  assign new_P3_SUB_450_U45 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_450_U15;
  assign new_P3_SUB_450_U46 = ~new_P3_SUB_450_U20;
  assign new_P3_SUB_450_U47 = ~new_P3_SUB_450_U46 | ~new_P3_SUB_450_U40;
  assign new_P3_SUB_450_U48 = ~new_P3_SUB_450_U20 | ~new_P3_SUB_450_U14;
  assign new_P3_SUB_450_U49 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_450_U12;
  assign new_P3_SUB_450_U50 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_450_U11;
  assign new_P3_SUB_450_U51 = ~new_P3_SUB_450_U21;
  assign new_P3_SUB_450_U52 = ~new_P3_SUB_450_U36 | ~new_P3_SUB_450_U51;
  assign new_P3_SUB_450_U53 = ~new_P3_SUB_450_U21 | ~new_P3_SUB_450_U24;
  assign new_P3_SUB_450_U54 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_450_U10;
  assign new_P3_SUB_450_U55 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_450_U9;
  assign new_P3_SUB_450_U56 = ~new_P3_SUB_450_U22;
  assign new_P3_SUB_450_U57 = ~new_P3_SUB_450_U32 | ~new_P3_SUB_450_U56;
  assign new_P3_SUB_450_U58 = ~new_P3_SUB_450_U22 | ~new_P3_SUB_450_U25;
  assign new_P3_SUB_450_U59 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_450_U8;
  assign new_P3_SUB_450_U60 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_450_U26;
  assign new_P3_SUB_450_U61 = ~new_P3_SUB_450_U23;
  assign new_P3_SUB_450_U62 = ~new_P3_SUB_450_U61 | ~new_P3_SUB_450_U28;
  assign new_P3_SUB_450_U63 = ~new_P3_SUB_450_U23 | ~new_P3_SUB_450_U7;
  assign new_P3_SUB_357_1258_U4 = P3_INSTADDRPOINTER_REG_27_ & P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_SUB_357_1258_U5 = new_P3_SUB_357_1258_U188 & new_P3_SUB_357_1258_U186;
  assign new_P3_SUB_357_1258_U6 = new_P3_SUB_357_1258_U187 & new_P3_SUB_357_1258_U178;
  assign new_P3_SUB_357_1258_U7 = new_P3_SUB_357_1258_U6 & new_P3_SUB_357_1258_U189;
  assign new_P3_SUB_357_1258_U8 = new_P3_SUB_357_1258_U5 & new_P3_SUB_357_1258_U190;
  assign new_P3_SUB_357_1258_U9 = new_P3_SUB_357_1258_U209 & new_P3_SUB_357_1258_U204;
  assign new_P3_SUB_357_1258_U10 = new_P3_SUB_357_1258_U156 & new_P3_SUB_357_1258_U206 & new_P3_SUB_357_1258_U210 & new_P3_SUB_357_1258_U205;
  assign new_P3_SUB_357_1258_U11 = new_P3_SUB_357_1258_U9 & new_P3_SUB_357_1258_U211;
  assign new_P3_SUB_357_1258_U12 = new_P3_SUB_357_1258_U10 & new_P3_SUB_357_1258_U212;
  assign new_P3_SUB_357_1258_U13 = new_P3_SUB_357_1258_U11 & new_P3_SUB_357_1258_U213;
  assign new_P3_SUB_357_1258_U14 = new_P3_SUB_357_1258_U12 & new_P3_SUB_357_1258_U214;
  assign new_P3_SUB_357_1258_U15 = new_P3_SUB_357_1258_U255 & new_P3_SUB_357_1258_U252;
  assign new_P3_SUB_357_1258_U16 = new_P3_SUB_357_1258_U249 & new_P3_SUB_357_1258_U248;
  assign new_P3_SUB_357_1258_U17 = new_P3_SUB_357_1258_U244 & new_P3_SUB_357_1258_U241;
  assign new_P3_SUB_357_1258_U18 = new_P3_SUB_357_1258_U233 & new_P3_SUB_357_1258_U230;
  assign new_P3_SUB_357_1258_U19 = new_P3_SUB_357_1258_U227 & new_P3_SUB_357_1258_U303;
  assign new_P3_SUB_357_1258_U20 = new_P3_SUB_357_1258_U225 & new_P3_SUB_357_1258_U296;
  assign new_P3_SUB_357_1258_U21 = ~new_P3_SUB_357_1258_U307 | ~new_P3_SUB_357_1258_U426 | ~new_P3_SUB_357_1258_U425;
  assign new_P3_SUB_357_1258_U22 = ~new_P3_ADD_357_U9;
  assign new_P3_SUB_357_1258_U23 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_SUB_357_1258_U24 = ~new_P3_ADD_357_U8;
  assign new_P3_SUB_357_1258_U25 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_SUB_357_1258_U26 = ~new_P3_ADD_357_U19;
  assign new_P3_SUB_357_1258_U27 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_SUB_357_1258_U28 = ~new_P3_ADD_357_U10;
  assign new_P3_SUB_357_1258_U29 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_SUB_357_1258_U30 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_357_U10;
  assign new_P3_SUB_357_1258_U31 = ~new_P3_SUB_357_U7;
  assign new_P3_SUB_357_1258_U32 = ~new_P3_ADD_357_U13;
  assign new_P3_SUB_357_1258_U33 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_SUB_357_1258_U34 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_SUB_357_1258_U35 = ~new_P3_ADD_357_U7;
  assign new_P3_SUB_357_1258_U36 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_SUB_357_1258_U37 = ~new_P3_ADD_357_U17;
  assign new_P3_SUB_357_1258_U38 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_SUB_357_1258_U39 = ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U40 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_SUB_357_1258_U41 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_SUB_357_1258_U42 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_SUB_357_1258_U43 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_SUB_357_1258_U44 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_SUB_357_1258_U45 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_SUB_357_1258_U46 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_SUB_357_1258_U47 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_SUB_357_1258_U48 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_SUB_357_1258_U49 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_SUB_357_1258_U50 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_SUB_357_1258_U51 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_SUB_357_1258_U52 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_SUB_357_1258_U53 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_SUB_357_1258_U54 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_SUB_357_1258_U55 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_SUB_357_1258_U56 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_SUB_357_1258_U57 = ~P3_INSTADDRPOINTER_REG_19_ | ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_SUB_357_1258_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_SUB_357_1258_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_SUB_357_1258_U60 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_SUB_357_1258_U61 = ~new_P3_SUB_357_1258_U269 | ~new_P3_SUB_357_1258_U222 | ~new_P3_SUB_357_1258_U151;
  assign new_P3_SUB_357_1258_U62 = ~new_P3_SUB_357_1258_U105 | ~new_P3_SUB_357_1258_U218;
  assign new_P3_SUB_357_1258_U63 = ~new_P3_SUB_357_1258_U104 | ~new_P3_SUB_357_1258_U284;
  assign new_P3_SUB_357_1258_U64 = ~new_P3_SUB_357_1258_U276 | ~new_P3_SUB_357_1258_U205;
  assign new_P3_SUB_357_1258_U65 = ~new_P3_SUB_357_1258_U277 | ~new_P3_SUB_357_1258_U47;
  assign new_P3_SUB_357_1258_U66 = ~new_P3_SUB_357_U7 | ~new_P3_SUB_357_1258_U161;
  assign new_P3_SUB_357_1258_U67 = ~new_P3_SUB_357_1258_U102 | ~new_P3_SUB_357_1258_U198;
  assign new_P3_SUB_357_1258_U68 = ~new_P3_SUB_357_1258_U290 | ~new_P3_SUB_357_1258_U8;
  assign new_P3_SUB_357_1258_U69 = ~new_P3_SUB_357_1258_U484 | ~new_P3_SUB_357_1258_U483;
  assign new_P3_SUB_357_1258_U70 = ~new_P3_SUB_357_1258_U312 | ~new_P3_SUB_357_1258_U311;
  assign new_P3_SUB_357_1258_U71 = ~new_P3_SUB_357_1258_U319 | ~new_P3_SUB_357_1258_U318;
  assign new_P3_SUB_357_1258_U72 = ~new_P3_SUB_357_1258_U326 | ~new_P3_SUB_357_1258_U325;
  assign new_P3_SUB_357_1258_U73 = ~new_P3_SUB_357_1258_U333 | ~new_P3_SUB_357_1258_U332;
  assign new_P3_SUB_357_1258_U74 = ~new_P3_SUB_357_1258_U340 | ~new_P3_SUB_357_1258_U339;
  assign new_P3_SUB_357_1258_U75 = ~new_P3_SUB_357_1258_U345 | ~new_P3_SUB_357_1258_U344;
  assign new_P3_SUB_357_1258_U76 = ~new_P3_SUB_357_1258_U350 | ~new_P3_SUB_357_1258_U349;
  assign new_P3_SUB_357_1258_U77 = ~new_P3_SUB_357_1258_U361 | ~new_P3_SUB_357_1258_U360;
  assign new_P3_SUB_357_1258_U78 = ~new_P3_SUB_357_1258_U366 | ~new_P3_SUB_357_1258_U365;
  assign new_P3_SUB_357_1258_U79 = ~new_P3_SUB_357_1258_U373 | ~new_P3_SUB_357_1258_U372;
  assign new_P3_SUB_357_1258_U80 = ~new_P3_SUB_357_1258_U384 | ~new_P3_SUB_357_1258_U383;
  assign new_P3_SUB_357_1258_U81 = ~new_P3_SUB_357_1258_U391 | ~new_P3_SUB_357_1258_U390;
  assign new_P3_SUB_357_1258_U82 = ~new_P3_SUB_357_1258_U398 | ~new_P3_SUB_357_1258_U397;
  assign new_P3_SUB_357_1258_U83 = ~new_P3_SUB_357_1258_U405 | ~new_P3_SUB_357_1258_U404;
  assign new_P3_SUB_357_1258_U84 = ~new_P3_SUB_357_1258_U412 | ~new_P3_SUB_357_1258_U411;
  assign new_P3_SUB_357_1258_U85 = ~new_P3_SUB_357_1258_U419 | ~new_P3_SUB_357_1258_U418;
  assign new_P3_SUB_357_1258_U86 = ~new_P3_SUB_357_1258_U431 | ~new_P3_SUB_357_1258_U430;
  assign new_P3_SUB_357_1258_U87 = ~new_P3_SUB_357_1258_U438 | ~new_P3_SUB_357_1258_U437;
  assign new_P3_SUB_357_1258_U88 = ~new_P3_SUB_357_1258_U449 | ~new_P3_SUB_357_1258_U448;
  assign new_P3_SUB_357_1258_U89 = ~new_P3_SUB_357_1258_U456 | ~new_P3_SUB_357_1258_U455;
  assign new_P3_SUB_357_1258_U90 = ~new_P3_SUB_357_1258_U463 | ~new_P3_SUB_357_1258_U462;
  assign new_P3_SUB_357_1258_U91 = ~new_P3_SUB_357_1258_U470 | ~new_P3_SUB_357_1258_U469;
  assign new_P3_SUB_357_1258_U92 = ~new_P3_SUB_357_1258_U477 | ~new_P3_SUB_357_1258_U476;
  assign new_P3_SUB_357_1258_U93 = ~new_P3_SUB_357_1258_U482 | ~new_P3_SUB_357_1258_U481;
  assign new_P3_SUB_357_1258_U94 = new_P3_SUB_357_1258_U160 & new_P3_SUB_357_1258_U163 & new_P3_SUB_357_1258_U164;
  assign new_P3_SUB_357_1258_U95 = new_P3_ADD_357_U7 & P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_SUB_357_1258_U96 = new_P3_SUB_357_1258_U168 & new_P3_SUB_357_1258_U162;
  assign new_P3_SUB_357_1258_U97 = new_P3_SUB_357_1258_U164 & new_P3_SUB_357_1258_U163;
  assign new_P3_SUB_357_1258_U98 = new_P3_SUB_357_1258_U7 & new_P3_SUB_357_1258_U154;
  assign new_P3_SUB_357_1258_U99 = new_P3_SUB_357_1258_U192 & new_P3_SUB_357_1258_U155;
  assign new_P3_SUB_357_1258_U100 = new_P3_SUB_357_1258_U99 & new_P3_SUB_357_1258_U8;
  assign new_P3_SUB_357_1258_U101 = P3_INSTADDRPOINTER_REG_17_ & P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_SUB_357_1258_U102 = new_P3_SUB_357_1258_U199 & new_P3_SUB_357_1258_U56;
  assign new_P3_SUB_357_1258_U103 = new_P3_SUB_357_1258_U215 & new_P3_SUB_357_1258_U13;
  assign new_P3_SUB_357_1258_U104 = new_P3_SUB_357_1258_U14 & new_P3_SUB_357_1258_U216;
  assign new_P3_SUB_357_1258_U105 = new_P3_SUB_357_1258_U219 & new_P3_SUB_357_1258_U157 & new_P3_SUB_357_1258_U58;
  assign new_P3_SUB_357_1258_U106 = new_P3_SUB_357_1258_U219 & new_P3_SUB_357_1258_U157;
  assign new_P3_SUB_357_1258_U107 = new_P3_SUB_357_1258_U269 & P3_INSTADDRPOINTER_REG_31_ & new_P3_SUB_357_1258_U60;
  assign new_P3_SUB_357_1258_U108 = P3_INSTADDRPOINTER_REG_30_ & P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_SUB_357_1258_U109 = new_P3_SUB_357_1258_U157 & new_P3_SUB_357_1258_U386 & new_P3_SUB_357_1258_U385;
  assign new_P3_SUB_357_1258_U110 = new_P3_SUB_357_1258_U232 & new_P3_SUB_357_1258_U153;
  assign new_P3_SUB_357_1258_U111 = new_P3_SUB_357_1258_U237 & new_P3_SUB_357_1258_U156;
  assign new_P3_SUB_357_1258_U112 = new_P3_SUB_357_1258_U243 & new_P3_SUB_357_1258_U156;
  assign new_P3_SUB_357_1258_U113 = new_P3_SUB_357_1258_U155 & new_P3_SUB_357_1258_U465 & new_P3_SUB_357_1258_U464;
  assign new_P3_SUB_357_1258_U114 = new_P3_SUB_357_1258_U254 & new_P3_SUB_357_1258_U154;
  assign new_P3_SUB_357_1258_U115 = ~new_P3_SUB_357_1258_U268 | ~new_P3_SUB_357_1258_U176 | ~new_P3_SUB_357_1258_U152;
  assign new_P3_SUB_357_1258_U116 = new_P3_SUB_357_1258_U314 & new_P3_SUB_357_1258_U313;
  assign new_P3_SUB_357_1258_U117 = ~new_P3_SUB_357_1258_U300 | ~new_P3_SUB_357_1258_U267;
  assign new_P3_SUB_357_1258_U118 = new_P3_SUB_357_1258_U321 & new_P3_SUB_357_1258_U320;
  assign new_P3_SUB_357_1258_U119 = ~new_P3_SUB_357_1258_U173 | ~new_P3_SUB_357_1258_U172;
  assign new_P3_SUB_357_1258_U120 = new_P3_SUB_357_1258_U328 & new_P3_SUB_357_1258_U327;
  assign new_P3_SUB_357_1258_U121 = ~new_P3_SUB_357_1258_U298 | ~new_P3_SUB_357_1258_U266;
  assign new_P3_SUB_357_1258_U122 = new_P3_SUB_357_1258_U335 & new_P3_SUB_357_1258_U334;
  assign new_P3_SUB_357_1258_U123 = ~new_P3_SUB_357_1258_U96 | ~new_P3_SUB_357_1258_U167;
  assign new_P3_SUB_357_1258_U124 = ~new_P3_SUB_357_1258_U181 | ~new_P3_SUB_357_1258_U180;
  assign new_P3_SUB_357_1258_U125 = ~new_P3_SUB_357_1258_U159 | ~new_P3_SUB_357_1258_U183;
  assign new_P3_SUB_357_1258_U126 = new_P3_SUB_357_1258_U356 & new_P3_SUB_357_1258_U355;
  assign new_P3_SUB_357_1258_U127 = ~new_P3_SUB_357_1258_U271 | ~new_P3_SUB_357_1258_U270 | ~new_P3_SUB_357_1258_U66;
  assign new_P3_SUB_357_1258_U128 = new_P3_SUB_357_1258_U368 & new_P3_SUB_357_1258_U367;
  assign new_P3_SUB_357_1258_U129 = ~new_P3_SUB_357_1258_U304 | ~new_P3_SUB_357_1258_U275 | ~new_P3_SUB_357_1258_U274;
  assign new_P3_SUB_357_1258_U130 = new_P3_SUB_357_1258_U379 & new_P3_SUB_357_1258_U378;
  assign new_P3_SUB_357_1258_U131 = ~new_P3_SUB_357_1258_U106 | ~new_P3_SUB_357_1258_U218;
  assign new_P3_SUB_357_1258_U132 = new_P3_SUB_357_1258_U393 & new_P3_SUB_357_1258_U392;
  assign new_P3_SUB_357_1258_U133 = ~new_P3_SUB_357_1258_U282 | ~new_P3_SUB_357_1258_U14;
  assign new_P3_SUB_357_1258_U134 = new_P3_SUB_357_1258_U400 & new_P3_SUB_357_1258_U399;
  assign new_P3_SUB_357_1258_U135 = ~new_P3_SUB_357_1258_U280 | ~new_P3_SUB_357_1258_U12;
  assign new_P3_SUB_357_1258_U136 = new_P3_SUB_357_1258_U407 & new_P3_SUB_357_1258_U406;
  assign new_P3_SUB_357_1258_U137 = ~new_P3_SUB_357_1258_U278 | ~new_P3_SUB_357_1258_U10;
  assign new_P3_SUB_357_1258_U138 = new_P3_SUB_357_1258_U414 & new_P3_SUB_357_1258_U413;
  assign new_P3_SUB_357_1258_U139 = ~new_P3_SUB_357_1258_U111 | ~new_P3_SUB_357_1258_U236;
  assign new_P3_SUB_357_1258_U140 = new_P3_SUB_357_1258_U433 & new_P3_SUB_357_1258_U432;
  assign new_P3_SUB_357_1258_U141 = ~new_P3_SUB_357_1258_U273 | ~new_P3_SUB_357_1258_U272 | ~new_P3_SUB_357_1258_U201;
  assign new_P3_SUB_357_1258_U142 = new_P3_SUB_357_1258_U444 & new_P3_SUB_357_1258_U443;
  assign new_P3_SUB_357_1258_U143 = ~new_P3_SUB_357_1258_U199 | ~new_P3_SUB_357_1258_U198;
  assign new_P3_SUB_357_1258_U144 = new_P3_SUB_357_1258_U451 & new_P3_SUB_357_1258_U450;
  assign new_P3_SUB_357_1258_U145 = ~new_P3_SUB_357_1258_U195 | ~new_P3_SUB_357_1258_U194;
  assign new_P3_SUB_357_1258_U146 = new_P3_SUB_357_1258_U458 & new_P3_SUB_357_1258_U457;
  assign new_P3_SUB_357_1258_U147 = ~new_P3_SUB_357_1258_U100 | ~new_P3_SUB_357_1258_U292;
  assign new_P3_SUB_357_1258_U148 = new_P3_SUB_357_1258_U472 & new_P3_SUB_357_1258_U471;
  assign new_P3_SUB_357_1258_U149 = ~new_P3_SUB_357_1258_U288 | ~new_P3_SUB_357_1258_U5;
  assign new_P3_SUB_357_1258_U150 = ~new_P3_SUB_357_1258_U286 | ~new_P3_SUB_357_1258_U186;
  assign new_P3_SUB_357_1258_U151 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U129;
  assign new_P3_SUB_357_1258_U152 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U117;
  assign new_P3_SUB_357_1258_U153 = ~new_P3_SUB_357_1258_U217 | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U154 = ~new_P3_SUB_357_1258_U191 | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U155 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U156 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U157 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U158 = ~new_P3_SUB_357_1258_U66;
  assign new_P3_SUB_357_1258_U159 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_357_U13;
  assign new_P3_SUB_357_1258_U160 = P3_INSTADDRPOINTER_REG_4_ | new_P3_ADD_357_U19;
  assign new_P3_SUB_357_1258_U161 = ~new_P3_SUB_357_1258_U30;
  assign new_P3_SUB_357_1258_U162 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_357_U19;
  assign new_P3_SUB_357_1258_U163 = new_P3_ADD_357_U7 | P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_SUB_357_1258_U164 = new_P3_ADD_357_U13 | P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_SUB_357_1258_U165 = ~new_P3_SUB_357_1258_U127;
  assign new_P3_SUB_357_1258_U166 = ~new_P3_SUB_357_1258_U66 | ~new_P3_SUB_357_1258_U159 | ~new_P3_SUB_357_1258_U271 | ~new_P3_SUB_357_1258_U270;
  assign new_P3_SUB_357_1258_U167 = ~new_P3_SUB_357_1258_U94 | ~new_P3_SUB_357_1258_U166;
  assign new_P3_SUB_357_1258_U168 = ~new_P3_SUB_357_1258_U95 | ~new_P3_SUB_357_1258_U160;
  assign new_P3_SUB_357_1258_U169 = ~new_P3_SUB_357_1258_U123;
  assign new_P3_SUB_357_1258_U170 = P3_INSTADDRPOINTER_REG_5_ | new_P3_ADD_357_U8;
  assign new_P3_SUB_357_1258_U171 = new_P3_ADD_357_U17 | P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_SUB_357_1258_U172 = ~new_P3_SUB_357_1258_U171 | ~new_P3_SUB_357_1258_U121;
  assign new_P3_SUB_357_1258_U173 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_357_U17;
  assign new_P3_SUB_357_1258_U174 = ~new_P3_SUB_357_1258_U119;
  assign new_P3_SUB_357_1258_U175 = P3_INSTADDRPOINTER_REG_7_ | new_P3_ADD_357_U9;
  assign new_P3_SUB_357_1258_U176 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_SUB_357_1258_U117;
  assign new_P3_SUB_357_1258_U177 = ~new_P3_SUB_357_1258_U115;
  assign new_P3_SUB_357_1258_U178 = P3_INSTADDRPOINTER_REG_9_ | new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U179 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U180 = ~new_P3_SUB_357_1258_U97 | ~new_P3_SUB_357_1258_U166;
  assign new_P3_SUB_357_1258_U181 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_357_U7;
  assign new_P3_SUB_357_1258_U182 = ~new_P3_SUB_357_1258_U124;
  assign new_P3_SUB_357_1258_U183 = ~new_P3_SUB_357_1258_U127 | ~new_P3_SUB_357_1258_U164;
  assign new_P3_SUB_357_1258_U184 = ~new_P3_SUB_357_1258_U125;
  assign new_P3_SUB_357_1258_U185 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_357_U7;
  assign new_P3_SUB_357_1258_U186 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U187 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_SUB_357_1258_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U189 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_SUB_357_1258_U190 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U191 = ~P3_INSTADDRPOINTER_REG_13_ | ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_SUB_357_1258_U192 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U193 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_SUB_357_1258_U194 = ~new_P3_SUB_357_1258_U193 | ~new_P3_SUB_357_1258_U147;
  assign new_P3_SUB_357_1258_U195 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U196 = ~new_P3_SUB_357_1258_U145;
  assign new_P3_SUB_357_1258_U197 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_SUB_357_1258_U198 = ~new_P3_SUB_357_1258_U197 | ~new_P3_SUB_357_1258_U145;
  assign new_P3_SUB_357_1258_U199 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U200 = ~new_P3_SUB_357_1258_U143;
  assign new_P3_SUB_357_1258_U201 = ~new_P3_SUB_357_1258_U101 | ~new_P3_SUB_357_1258_U143;
  assign new_P3_SUB_357_1258_U202 = ~new_P3_SUB_357_1258_U67;
  assign new_P3_SUB_357_1258_U203 = ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U204 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_SUB_357_1258_U205 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U206 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U207 = ~new_P3_SUB_357_1258_U57;
  assign new_P3_SUB_357_1258_U208 = ~new_P3_SUB_357_1258_U207 | ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_SUB_357_1258_U209 = ~new_P3_SUB_357_1258_U39 | ~new_P3_SUB_357_1258_U208;
  assign new_P3_SUB_357_1258_U210 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U211 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_SUB_357_1258_U212 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U213 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_SUB_357_1258_U214 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U215 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_SUB_357_1258_U216 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U217 = ~P3_INSTADDRPOINTER_REG_26_ | ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_SUB_357_1258_U218 = ~new_P3_SUB_357_1258_U63 | ~new_P3_SUB_357_1258_U153;
  assign new_P3_SUB_357_1258_U219 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U220 = ~new_P3_SUB_357_1258_U131;
  assign new_P3_SUB_357_1258_U221 = ~new_P3_SUB_357_1258_U62;
  assign new_P3_SUB_357_1258_U222 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_SUB_357_1258_U129;
  assign new_P3_SUB_357_1258_U223 = ~new_P3_SUB_357_1258_U61;
  assign new_P3_SUB_357_1258_U224 = ~new_P3_SUB_357_1258_U151 | ~new_P3_SUB_357_1258_U107;
  assign new_P3_SUB_357_1258_U225 = ~new_P3_SUB_357_1258_U294 | ~new_P3_SUB_357_1258_U354 | ~new_P3_SUB_357_1258_U353;
  assign new_P3_SUB_357_1258_U226 = ~new_P3_SUB_357_1258_U221 | ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_SUB_357_1258_U227 = ~new_P3_SUB_357_1258_U62 | ~new_P3_SUB_357_1258_U377 | ~new_P3_SUB_357_1258_U376;
  assign new_P3_SUB_357_1258_U228 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_SUB_357_1258_U229 = ~new_P3_SUB_357_1258_U228 | ~new_P3_SUB_357_1258_U63;
  assign new_P3_SUB_357_1258_U230 = ~new_P3_SUB_357_1258_U109 | ~new_P3_SUB_357_1258_U229;
  assign new_P3_SUB_357_1258_U231 = ~new_P3_SUB_357_1258_U285 | ~new_P3_SUB_357_1258_U157;
  assign new_P3_SUB_357_1258_U232 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U233 = ~new_P3_SUB_357_1258_U110 | ~new_P3_SUB_357_1258_U231;
  assign new_P3_SUB_357_1258_U234 = P3_INSTADDRPOINTER_REG_25_ | new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U235 = ~new_P3_SUB_357_1258_U65;
  assign new_P3_SUB_357_1258_U236 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U65;
  assign new_P3_SUB_357_1258_U237 = ~new_P3_SUB_357_1258_U207 | ~new_P3_SUB_357_1258_U64;
  assign new_P3_SUB_357_1258_U238 = ~new_P3_SUB_357_1258_U139;
  assign new_P3_SUB_357_1258_U239 = ~new_P3_SUB_357_1258_U235 | ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_SUB_357_1258_U240 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_SUB_357_1258_U64;
  assign new_P3_SUB_357_1258_U241 = ~new_P3_SUB_357_1258_U240 | ~new_P3_SUB_357_1258_U421 | ~new_P3_SUB_357_1258_U420;
  assign new_P3_SUB_357_1258_U242 = ~new_P3_SUB_357_1258_U277 | ~new_P3_SUB_357_1258_U206;
  assign new_P3_SUB_357_1258_U243 = ~new_P3_SUB_357_1258_U57 | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U244 = ~new_P3_SUB_357_1258_U112 | ~new_P3_SUB_357_1258_U242;
  assign new_P3_SUB_357_1258_U245 = P3_INSTADDRPOINTER_REG_19_ | new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U246 = ~new_P3_SUB_357_1258_U202 | ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_SUB_357_1258_U247 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_SUB_357_1258_U143;
  assign new_P3_SUB_357_1258_U248 = ~new_P3_SUB_357_1258_U247 | ~new_P3_SUB_357_1258_U440 | ~new_P3_SUB_357_1258_U439;
  assign new_P3_SUB_357_1258_U249 = ~new_P3_SUB_357_1258_U67 | ~new_P3_SUB_357_1258_U442 | ~new_P3_SUB_357_1258_U441;
  assign new_P3_SUB_357_1258_U250 = new_P3_ADD_357_U6 | P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_SUB_357_1258_U251 = ~new_P3_SUB_357_1258_U250 | ~new_P3_SUB_357_1258_U68;
  assign new_P3_SUB_357_1258_U252 = ~new_P3_SUB_357_1258_U113 | ~new_P3_SUB_357_1258_U251;
  assign new_P3_SUB_357_1258_U253 = ~new_P3_SUB_357_1258_U291 | ~new_P3_SUB_357_1258_U155;
  assign new_P3_SUB_357_1258_U254 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U255 = ~new_P3_SUB_357_1258_U114 | ~new_P3_SUB_357_1258_U253;
  assign new_P3_SUB_357_1258_U256 = P3_INSTADDRPOINTER_REG_12_ | new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U257 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U258 = ~new_P3_SUB_357_1258_U179 | ~new_P3_SUB_357_1258_U178;
  assign new_P3_SUB_357_1258_U259 = ~new_P3_SUB_357_1258_U162 | ~new_P3_SUB_357_1258_U160;
  assign new_P3_SUB_357_1258_U260 = ~new_P3_SUB_357_1258_U185 | ~new_P3_SUB_357_1258_U163;
  assign new_P3_SUB_357_1258_U261 = ~new_P3_SUB_357_1258_U164 | ~new_P3_SUB_357_1258_U159;
  assign new_P3_SUB_357_1258_U262 = ~new_P3_SUB_357_1258_U234 | ~new_P3_SUB_357_1258_U157;
  assign new_P3_SUB_357_1258_U263 = ~new_P3_SUB_357_1258_U245 | ~new_P3_SUB_357_1258_U206;
  assign new_P3_SUB_357_1258_U264 = ~new_P3_SUB_357_1258_U256 | ~new_P3_SUB_357_1258_U155;
  assign new_P3_SUB_357_1258_U265 = ~new_P3_SUB_357_1258_U257 | ~new_P3_SUB_357_1258_U187;
  assign new_P3_SUB_357_1258_U266 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_357_U8;
  assign new_P3_SUB_357_1258_U267 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_357_U9;
  assign new_P3_SUB_357_1258_U268 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U269 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U270 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_SUB_357_1258_U161;
  assign new_P3_SUB_357_1258_U271 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_SUB_357_U7;
  assign new_P3_SUB_357_1258_U272 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U67;
  assign new_P3_SUB_357_1258_U273 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U274 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U62;
  assign new_P3_SUB_357_1258_U275 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U276 = ~new_P3_SUB_357_1258_U204 | ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U277 = ~new_P3_SUB_357_1258_U64;
  assign new_P3_SUB_357_1258_U278 = ~new_P3_SUB_357_1258_U9 | ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U279 = ~new_P3_SUB_357_1258_U137;
  assign new_P3_SUB_357_1258_U280 = ~new_P3_SUB_357_1258_U11 | ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U281 = ~new_P3_SUB_357_1258_U135;
  assign new_P3_SUB_357_1258_U282 = ~new_P3_SUB_357_1258_U13 | ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U283 = ~new_P3_SUB_357_1258_U133;
  assign new_P3_SUB_357_1258_U284 = ~new_P3_SUB_357_1258_U103 | ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U285 = ~new_P3_SUB_357_1258_U63;
  assign new_P3_SUB_357_1258_U286 = ~new_P3_SUB_357_1258_U178 | ~new_P3_SUB_357_1258_U115;
  assign new_P3_SUB_357_1258_U287 = ~new_P3_SUB_357_1258_U150;
  assign new_P3_SUB_357_1258_U288 = ~new_P3_SUB_357_1258_U6 | ~new_P3_SUB_357_1258_U115;
  assign new_P3_SUB_357_1258_U289 = ~new_P3_SUB_357_1258_U149;
  assign new_P3_SUB_357_1258_U290 = ~new_P3_SUB_357_1258_U7 | ~new_P3_SUB_357_1258_U115;
  assign new_P3_SUB_357_1258_U291 = ~new_P3_SUB_357_1258_U68;
  assign new_P3_SUB_357_1258_U292 = ~new_P3_SUB_357_1258_U98 | ~new_P3_SUB_357_1258_U115;
  assign new_P3_SUB_357_1258_U293 = ~new_P3_SUB_357_1258_U147;
  assign new_P3_SUB_357_1258_U294 = ~new_P3_SUB_357_1258_U223 | ~new_P3_SUB_357_1258_U60;
  assign new_P3_SUB_357_1258_U295 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_SUB_357_1258_U61;
  assign new_P3_SUB_357_1258_U296 = ~new_P3_SUB_357_1258_U295 | ~new_P3_SUB_357_1258_U352 | ~new_P3_SUB_357_1258_U351;
  assign new_P3_SUB_357_1258_U297 = ~new_P3_SUB_357_1258_U108 | ~new_P3_SUB_357_1258_U61;
  assign new_P3_SUB_357_1258_U298 = ~new_P3_SUB_357_1258_U170 | ~new_P3_SUB_357_1258_U123;
  assign new_P3_SUB_357_1258_U299 = ~new_P3_SUB_357_1258_U121;
  assign new_P3_SUB_357_1258_U300 = ~new_P3_SUB_357_1258_U175 | ~new_P3_SUB_357_1258_U119;
  assign new_P3_SUB_357_1258_U301 = ~new_P3_SUB_357_1258_U117;
  assign new_P3_SUB_357_1258_U302 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_SUB_357_1258_U131;
  assign new_P3_SUB_357_1258_U303 = ~new_P3_SUB_357_1258_U302 | ~new_P3_SUB_357_1258_U375 | ~new_P3_SUB_357_1258_U374;
  assign new_P3_SUB_357_1258_U304 = ~new_P3_SUB_357_1258_U4 | ~new_P3_SUB_357_1258_U131;
  assign new_P3_SUB_357_1258_U305 = ~new_P3_SUB_357_1258_U129;
  assign new_P3_SUB_357_1258_U306 = ~new_P3_SUB_357_1258_U4 | ~new_P3_SUB_357_1258_U131;
  assign new_P3_SUB_357_1258_U307 = ~new_P3_SUB_357_1258_U158 | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_SUB_357_1258_U308 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U41;
  assign new_P3_SUB_357_1258_U309 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U310 = ~new_P3_SUB_357_1258_U309 | ~new_P3_SUB_357_1258_U308;
  assign new_P3_SUB_357_1258_U311 = ~new_P3_SUB_357_1258_U258 | ~new_P3_SUB_357_1258_U115;
  assign new_P3_SUB_357_1258_U312 = ~new_P3_SUB_357_1258_U177 | ~new_P3_SUB_357_1258_U310;
  assign new_P3_SUB_357_1258_U313 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U40;
  assign new_P3_SUB_357_1258_U314 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U315 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U40;
  assign new_P3_SUB_357_1258_U316 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U317 = ~new_P3_SUB_357_1258_U316 | ~new_P3_SUB_357_1258_U315;
  assign new_P3_SUB_357_1258_U318 = ~new_P3_SUB_357_1258_U116 | ~new_P3_SUB_357_1258_U117;
  assign new_P3_SUB_357_1258_U319 = ~new_P3_SUB_357_1258_U301 | ~new_P3_SUB_357_1258_U317;
  assign new_P3_SUB_357_1258_U320 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_SUB_357_1258_U22;
  assign new_P3_SUB_357_1258_U321 = ~new_P3_ADD_357_U9 | ~new_P3_SUB_357_1258_U23;
  assign new_P3_SUB_357_1258_U322 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_SUB_357_1258_U22;
  assign new_P3_SUB_357_1258_U323 = ~new_P3_ADD_357_U9 | ~new_P3_SUB_357_1258_U23;
  assign new_P3_SUB_357_1258_U324 = ~new_P3_SUB_357_1258_U323 | ~new_P3_SUB_357_1258_U322;
  assign new_P3_SUB_357_1258_U325 = ~new_P3_SUB_357_1258_U118 | ~new_P3_SUB_357_1258_U119;
  assign new_P3_SUB_357_1258_U326 = ~new_P3_SUB_357_1258_U174 | ~new_P3_SUB_357_1258_U324;
  assign new_P3_SUB_357_1258_U327 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_SUB_357_1258_U37;
  assign new_P3_SUB_357_1258_U328 = ~new_P3_ADD_357_U17 | ~new_P3_SUB_357_1258_U38;
  assign new_P3_SUB_357_1258_U329 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_SUB_357_1258_U37;
  assign new_P3_SUB_357_1258_U330 = ~new_P3_ADD_357_U17 | ~new_P3_SUB_357_1258_U38;
  assign new_P3_SUB_357_1258_U331 = ~new_P3_SUB_357_1258_U330 | ~new_P3_SUB_357_1258_U329;
  assign new_P3_SUB_357_1258_U332 = ~new_P3_SUB_357_1258_U120 | ~new_P3_SUB_357_1258_U121;
  assign new_P3_SUB_357_1258_U333 = ~new_P3_SUB_357_1258_U299 | ~new_P3_SUB_357_1258_U331;
  assign new_P3_SUB_357_1258_U334 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_SUB_357_1258_U24;
  assign new_P3_SUB_357_1258_U335 = ~new_P3_ADD_357_U8 | ~new_P3_SUB_357_1258_U25;
  assign new_P3_SUB_357_1258_U336 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_SUB_357_1258_U24;
  assign new_P3_SUB_357_1258_U337 = ~new_P3_ADD_357_U8 | ~new_P3_SUB_357_1258_U25;
  assign new_P3_SUB_357_1258_U338 = ~new_P3_SUB_357_1258_U337 | ~new_P3_SUB_357_1258_U336;
  assign new_P3_SUB_357_1258_U339 = ~new_P3_SUB_357_1258_U122 | ~new_P3_SUB_357_1258_U123;
  assign new_P3_SUB_357_1258_U340 = ~new_P3_SUB_357_1258_U169 | ~new_P3_SUB_357_1258_U338;
  assign new_P3_SUB_357_1258_U341 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_SUB_357_1258_U26;
  assign new_P3_SUB_357_1258_U342 = ~new_P3_ADD_357_U19 | ~new_P3_SUB_357_1258_U27;
  assign new_P3_SUB_357_1258_U343 = ~new_P3_SUB_357_1258_U342 | ~new_P3_SUB_357_1258_U341;
  assign new_P3_SUB_357_1258_U344 = ~new_P3_SUB_357_1258_U259 | ~new_P3_SUB_357_1258_U124;
  assign new_P3_SUB_357_1258_U345 = ~new_P3_SUB_357_1258_U182 | ~new_P3_SUB_357_1258_U343;
  assign new_P3_SUB_357_1258_U346 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_SUB_357_1258_U35;
  assign new_P3_SUB_357_1258_U347 = ~new_P3_ADD_357_U7 | ~new_P3_SUB_357_1258_U36;
  assign new_P3_SUB_357_1258_U348 = ~new_P3_SUB_357_1258_U347 | ~new_P3_SUB_357_1258_U346;
  assign new_P3_SUB_357_1258_U349 = ~new_P3_SUB_357_1258_U260 | ~new_P3_SUB_357_1258_U125;
  assign new_P3_SUB_357_1258_U350 = ~new_P3_SUB_357_1258_U184 | ~new_P3_SUB_357_1258_U348;
  assign new_P3_SUB_357_1258_U351 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U352 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U224;
  assign new_P3_SUB_357_1258_U353 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U354 = ~new_P3_SUB_357_1258_U297 | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U355 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U60;
  assign new_P3_SUB_357_1258_U356 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U357 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U60;
  assign new_P3_SUB_357_1258_U358 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U359 = ~new_P3_SUB_357_1258_U358 | ~new_P3_SUB_357_1258_U357;
  assign new_P3_SUB_357_1258_U360 = ~new_P3_SUB_357_1258_U126 | ~new_P3_SUB_357_1258_U61;
  assign new_P3_SUB_357_1258_U361 = ~new_P3_SUB_357_1258_U359 | ~new_P3_SUB_357_1258_U223;
  assign new_P3_SUB_357_1258_U362 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_SUB_357_1258_U32;
  assign new_P3_SUB_357_1258_U363 = ~new_P3_ADD_357_U13 | ~new_P3_SUB_357_1258_U33;
  assign new_P3_SUB_357_1258_U364 = ~new_P3_SUB_357_1258_U363 | ~new_P3_SUB_357_1258_U362;
  assign new_P3_SUB_357_1258_U365 = ~new_P3_SUB_357_1258_U261 | ~new_P3_SUB_357_1258_U127;
  assign new_P3_SUB_357_1258_U366 = ~new_P3_SUB_357_1258_U165 | ~new_P3_SUB_357_1258_U364;
  assign new_P3_SUB_357_1258_U367 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U59;
  assign new_P3_SUB_357_1258_U368 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U369 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U59;
  assign new_P3_SUB_357_1258_U370 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U371 = ~new_P3_SUB_357_1258_U370 | ~new_P3_SUB_357_1258_U369;
  assign new_P3_SUB_357_1258_U372 = ~new_P3_SUB_357_1258_U128 | ~new_P3_SUB_357_1258_U129;
  assign new_P3_SUB_357_1258_U373 = ~new_P3_SUB_357_1258_U305 | ~new_P3_SUB_357_1258_U371;
  assign new_P3_SUB_357_1258_U374 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U375 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U226;
  assign new_P3_SUB_357_1258_U376 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U377 = ~new_P3_SUB_357_1258_U306 | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U378 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U379 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U58;
  assign new_P3_SUB_357_1258_U380 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U381 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U58;
  assign new_P3_SUB_357_1258_U382 = ~new_P3_SUB_357_1258_U381 | ~new_P3_SUB_357_1258_U380;
  assign new_P3_SUB_357_1258_U383 = ~new_P3_SUB_357_1258_U130 | ~new_P3_SUB_357_1258_U131;
  assign new_P3_SUB_357_1258_U384 = ~new_P3_SUB_357_1258_U220 | ~new_P3_SUB_357_1258_U382;
  assign new_P3_SUB_357_1258_U385 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U386 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U43;
  assign new_P3_SUB_357_1258_U387 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U388 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U42;
  assign new_P3_SUB_357_1258_U389 = ~new_P3_SUB_357_1258_U388 | ~new_P3_SUB_357_1258_U387;
  assign new_P3_SUB_357_1258_U390 = ~new_P3_SUB_357_1258_U63 | ~new_P3_SUB_357_1258_U262;
  assign new_P3_SUB_357_1258_U391 = ~new_P3_SUB_357_1258_U389 | ~new_P3_SUB_357_1258_U285;
  assign new_P3_SUB_357_1258_U392 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U393 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U44;
  assign new_P3_SUB_357_1258_U394 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U395 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U44;
  assign new_P3_SUB_357_1258_U396 = ~new_P3_SUB_357_1258_U395 | ~new_P3_SUB_357_1258_U394;
  assign new_P3_SUB_357_1258_U397 = ~new_P3_SUB_357_1258_U132 | ~new_P3_SUB_357_1258_U133;
  assign new_P3_SUB_357_1258_U398 = ~new_P3_SUB_357_1258_U283 | ~new_P3_SUB_357_1258_U396;
  assign new_P3_SUB_357_1258_U399 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U400 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U45;
  assign new_P3_SUB_357_1258_U401 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U402 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U45;
  assign new_P3_SUB_357_1258_U403 = ~new_P3_SUB_357_1258_U402 | ~new_P3_SUB_357_1258_U401;
  assign new_P3_SUB_357_1258_U404 = ~new_P3_SUB_357_1258_U134 | ~new_P3_SUB_357_1258_U135;
  assign new_P3_SUB_357_1258_U405 = ~new_P3_SUB_357_1258_U281 | ~new_P3_SUB_357_1258_U403;
  assign new_P3_SUB_357_1258_U406 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U407 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U46;
  assign new_P3_SUB_357_1258_U408 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U409 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U46;
  assign new_P3_SUB_357_1258_U410 = ~new_P3_SUB_357_1258_U409 | ~new_P3_SUB_357_1258_U408;
  assign new_P3_SUB_357_1258_U411 = ~new_P3_SUB_357_1258_U136 | ~new_P3_SUB_357_1258_U137;
  assign new_P3_SUB_357_1258_U412 = ~new_P3_SUB_357_1258_U279 | ~new_P3_SUB_357_1258_U410;
  assign new_P3_SUB_357_1258_U413 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U414 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U48;
  assign new_P3_SUB_357_1258_U415 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U416 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U48;
  assign new_P3_SUB_357_1258_U417 = ~new_P3_SUB_357_1258_U416 | ~new_P3_SUB_357_1258_U415;
  assign new_P3_SUB_357_1258_U418 = ~new_P3_SUB_357_1258_U138 | ~new_P3_SUB_357_1258_U139;
  assign new_P3_SUB_357_1258_U419 = ~new_P3_SUB_357_1258_U238 | ~new_P3_SUB_357_1258_U417;
  assign new_P3_SUB_357_1258_U420 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U421 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U239;
  assign new_P3_SUB_357_1258_U422 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_SUB_357_1258_U30;
  assign new_P3_SUB_357_1258_U423 = ~new_P3_SUB_357_1258_U161 | ~new_P3_SUB_357_1258_U34;
  assign new_P3_SUB_357_1258_U424 = ~new_P3_SUB_357_1258_U423 | ~new_P3_SUB_357_1258_U422;
  assign new_P3_SUB_357_1258_U425 = ~new_P3_SUB_357_U7 | ~new_P3_SUB_357_1258_U30 | ~new_P3_SUB_357_1258_U34;
  assign new_P3_SUB_357_1258_U426 = ~new_P3_SUB_357_1258_U424 | ~new_P3_SUB_357_1258_U31;
  assign new_P3_SUB_357_1258_U427 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U428 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U47;
  assign new_P3_SUB_357_1258_U429 = ~new_P3_SUB_357_1258_U428 | ~new_P3_SUB_357_1258_U427;
  assign new_P3_SUB_357_1258_U430 = ~new_P3_SUB_357_1258_U64 | ~new_P3_SUB_357_1258_U263;
  assign new_P3_SUB_357_1258_U431 = ~new_P3_SUB_357_1258_U429 | ~new_P3_SUB_357_1258_U277;
  assign new_P3_SUB_357_1258_U432 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U433 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U49;
  assign new_P3_SUB_357_1258_U434 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U435 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U49;
  assign new_P3_SUB_357_1258_U436 = ~new_P3_SUB_357_1258_U435 | ~new_P3_SUB_357_1258_U434;
  assign new_P3_SUB_357_1258_U437 = ~new_P3_SUB_357_1258_U140 | ~new_P3_SUB_357_1258_U141;
  assign new_P3_SUB_357_1258_U438 = ~new_P3_SUB_357_1258_U203 | ~new_P3_SUB_357_1258_U436;
  assign new_P3_SUB_357_1258_U439 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U440 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U246;
  assign new_P3_SUB_357_1258_U441 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_357_U6;
  assign new_P3_SUB_357_1258_U442 = ~new_P3_SUB_357_1258_U201 | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U443 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U444 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U56;
  assign new_P3_SUB_357_1258_U445 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U446 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U56;
  assign new_P3_SUB_357_1258_U447 = ~new_P3_SUB_357_1258_U446 | ~new_P3_SUB_357_1258_U445;
  assign new_P3_SUB_357_1258_U448 = ~new_P3_SUB_357_1258_U142 | ~new_P3_SUB_357_1258_U143;
  assign new_P3_SUB_357_1258_U449 = ~new_P3_SUB_357_1258_U200 | ~new_P3_SUB_357_1258_U447;
  assign new_P3_SUB_357_1258_U450 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U451 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U55;
  assign new_P3_SUB_357_1258_U452 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U453 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U55;
  assign new_P3_SUB_357_1258_U454 = ~new_P3_SUB_357_1258_U453 | ~new_P3_SUB_357_1258_U452;
  assign new_P3_SUB_357_1258_U455 = ~new_P3_SUB_357_1258_U144 | ~new_P3_SUB_357_1258_U145;
  assign new_P3_SUB_357_1258_U456 = ~new_P3_SUB_357_1258_U196 | ~new_P3_SUB_357_1258_U454;
  assign new_P3_SUB_357_1258_U457 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U458 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U54;
  assign new_P3_SUB_357_1258_U459 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U460 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U54;
  assign new_P3_SUB_357_1258_U461 = ~new_P3_SUB_357_1258_U460 | ~new_P3_SUB_357_1258_U459;
  assign new_P3_SUB_357_1258_U462 = ~new_P3_SUB_357_1258_U146 | ~new_P3_SUB_357_1258_U147;
  assign new_P3_SUB_357_1258_U463 = ~new_P3_SUB_357_1258_U293 | ~new_P3_SUB_357_1258_U461;
  assign new_P3_SUB_357_1258_U464 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U465 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U51;
  assign new_P3_SUB_357_1258_U466 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U467 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U50;
  assign new_P3_SUB_357_1258_U468 = ~new_P3_SUB_357_1258_U467 | ~new_P3_SUB_357_1258_U466;
  assign new_P3_SUB_357_1258_U469 = ~new_P3_SUB_357_1258_U68 | ~new_P3_SUB_357_1258_U264;
  assign new_P3_SUB_357_1258_U470 = ~new_P3_SUB_357_1258_U468 | ~new_P3_SUB_357_1258_U291;
  assign new_P3_SUB_357_1258_U471 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U472 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U52;
  assign new_P3_SUB_357_1258_U473 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U474 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U52;
  assign new_P3_SUB_357_1258_U475 = ~new_P3_SUB_357_1258_U474 | ~new_P3_SUB_357_1258_U473;
  assign new_P3_SUB_357_1258_U476 = ~new_P3_SUB_357_1258_U148 | ~new_P3_SUB_357_1258_U149;
  assign new_P3_SUB_357_1258_U477 = ~new_P3_SUB_357_1258_U289 | ~new_P3_SUB_357_1258_U475;
  assign new_P3_SUB_357_1258_U478 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_SUB_357_1258_U39;
  assign new_P3_SUB_357_1258_U479 = ~new_P3_ADD_357_U6 | ~new_P3_SUB_357_1258_U53;
  assign new_P3_SUB_357_1258_U480 = ~new_P3_SUB_357_1258_U479 | ~new_P3_SUB_357_1258_U478;
  assign new_P3_SUB_357_1258_U481 = ~new_P3_SUB_357_1258_U150 | ~new_P3_SUB_357_1258_U265;
  assign new_P3_SUB_357_1258_U482 = ~new_P3_SUB_357_1258_U287 | ~new_P3_SUB_357_1258_U480;
  assign new_P3_SUB_357_1258_U483 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_SUB_357_1258_U28;
  assign new_P3_SUB_357_1258_U484 = ~new_P3_ADD_357_U10 | ~new_P3_SUB_357_1258_U29;
  assign new_P3_ADD_486_U5 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_ADD_486_U6 = P3_INSTQUEUERD_ADDR_REG_4_ & new_P3_ADD_486_U20;
  assign new_P3_ADD_486_U7 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_ADD_486_U8 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_ADD_486_U9 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_ADD_486_U10 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_ADD_486_U18;
  assign new_P3_ADD_486_U11 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_ADD_486_U12 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_ADD_486_U19;
  assign new_P3_ADD_486_U13 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_ADD_486_U14 = ~new_P3_ADD_486_U22 | ~new_P3_ADD_486_U21;
  assign new_P3_ADD_486_U15 = ~new_P3_ADD_486_U24 | ~new_P3_ADD_486_U23;
  assign new_P3_ADD_486_U16 = ~new_P3_ADD_486_U26 | ~new_P3_ADD_486_U25;
  assign new_P3_ADD_486_U17 = ~new_P3_ADD_486_U28 | ~new_P3_ADD_486_U27;
  assign new_P3_ADD_486_U18 = ~new_P3_ADD_486_U8;
  assign new_P3_ADD_486_U19 = ~new_P3_ADD_486_U10;
  assign new_P3_ADD_486_U20 = ~new_P3_ADD_486_U12;
  assign new_P3_ADD_486_U21 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_ADD_486_U12;
  assign new_P3_ADD_486_U22 = ~new_P3_ADD_486_U20 | ~new_P3_ADD_486_U13;
  assign new_P3_ADD_486_U23 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_ADD_486_U10;
  assign new_P3_ADD_486_U24 = ~new_P3_ADD_486_U19 | ~new_P3_ADD_486_U11;
  assign new_P3_ADD_486_U25 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_ADD_486_U8;
  assign new_P3_ADD_486_U26 = ~new_P3_ADD_486_U18 | ~new_P3_ADD_486_U9;
  assign new_P3_ADD_486_U27 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_ADD_486_U5;
  assign new_P3_ADD_486_U28 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_ADD_486_U7;
  assign new_P3_SUB_485_U6 = ~new_P3_SUB_485_U43 | ~new_P3_SUB_485_U42;
  assign new_P3_SUB_485_U7 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_485_U27;
  assign new_P3_SUB_485_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_485_U9 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_485_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_485_U11 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_485_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_485_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_485_U14 = ~new_P3_SUB_485_U39 | ~new_P3_SUB_485_U38;
  assign new_P3_SUB_485_U15 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_485_U16 = ~new_P3_SUB_485_U48 | ~new_P3_SUB_485_U47;
  assign new_P3_SUB_485_U17 = ~new_P3_SUB_485_U53 | ~new_P3_SUB_485_U52;
  assign new_P3_SUB_485_U18 = ~new_P3_SUB_485_U58 | ~new_P3_SUB_485_U57;
  assign new_P3_SUB_485_U19 = ~new_P3_SUB_485_U63 | ~new_P3_SUB_485_U62;
  assign new_P3_SUB_485_U20 = ~new_P3_SUB_485_U45 | ~new_P3_SUB_485_U44;
  assign new_P3_SUB_485_U21 = ~new_P3_SUB_485_U50 | ~new_P3_SUB_485_U49;
  assign new_P3_SUB_485_U22 = ~new_P3_SUB_485_U55 | ~new_P3_SUB_485_U54;
  assign new_P3_SUB_485_U23 = ~new_P3_SUB_485_U60 | ~new_P3_SUB_485_U59;
  assign new_P3_SUB_485_U24 = ~new_P3_SUB_485_U35 | ~new_P3_SUB_485_U34;
  assign new_P3_SUB_485_U25 = ~new_P3_SUB_485_U31 | ~new_P3_SUB_485_U30;
  assign new_P3_SUB_485_U26 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_485_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_485_U28 = ~new_P3_SUB_485_U7;
  assign new_P3_SUB_485_U29 = ~new_P3_SUB_485_U28 | ~new_P3_SUB_485_U8;
  assign new_P3_SUB_485_U30 = ~new_P3_SUB_485_U29 | ~new_P3_SUB_485_U26;
  assign new_P3_SUB_485_U31 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_485_U7;
  assign new_P3_SUB_485_U32 = ~new_P3_SUB_485_U25;
  assign new_P3_SUB_485_U33 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_485_U10;
  assign new_P3_SUB_485_U34 = ~new_P3_SUB_485_U33 | ~new_P3_SUB_485_U25;
  assign new_P3_SUB_485_U35 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_485_U9;
  assign new_P3_SUB_485_U36 = ~new_P3_SUB_485_U24;
  assign new_P3_SUB_485_U37 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_485_U12;
  assign new_P3_SUB_485_U38 = ~new_P3_SUB_485_U37 | ~new_P3_SUB_485_U24;
  assign new_P3_SUB_485_U39 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_485_U11;
  assign new_P3_SUB_485_U40 = ~new_P3_SUB_485_U14;
  assign new_P3_SUB_485_U41 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_485_U15;
  assign new_P3_SUB_485_U42 = ~new_P3_SUB_485_U40 | ~new_P3_SUB_485_U41;
  assign new_P3_SUB_485_U43 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_485_U13;
  assign new_P3_SUB_485_U44 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_485_U13;
  assign new_P3_SUB_485_U45 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_485_U15;
  assign new_P3_SUB_485_U46 = ~new_P3_SUB_485_U20;
  assign new_P3_SUB_485_U47 = ~new_P3_SUB_485_U46 | ~new_P3_SUB_485_U40;
  assign new_P3_SUB_485_U48 = ~new_P3_SUB_485_U20 | ~new_P3_SUB_485_U14;
  assign new_P3_SUB_485_U49 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_485_U12;
  assign new_P3_SUB_485_U50 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_485_U11;
  assign new_P3_SUB_485_U51 = ~new_P3_SUB_485_U21;
  assign new_P3_SUB_485_U52 = ~new_P3_SUB_485_U36 | ~new_P3_SUB_485_U51;
  assign new_P3_SUB_485_U53 = ~new_P3_SUB_485_U21 | ~new_P3_SUB_485_U24;
  assign new_P3_SUB_485_U54 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_485_U10;
  assign new_P3_SUB_485_U55 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_485_U9;
  assign new_P3_SUB_485_U56 = ~new_P3_SUB_485_U22;
  assign new_P3_SUB_485_U57 = ~new_P3_SUB_485_U32 | ~new_P3_SUB_485_U56;
  assign new_P3_SUB_485_U58 = ~new_P3_SUB_485_U22 | ~new_P3_SUB_485_U25;
  assign new_P3_SUB_485_U59 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_485_U8;
  assign new_P3_SUB_485_U60 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_485_U26;
  assign new_P3_SUB_485_U61 = ~new_P3_SUB_485_U23;
  assign new_P3_SUB_485_U62 = ~new_P3_SUB_485_U61 | ~new_P3_SUB_485_U28;
  assign new_P3_SUB_485_U63 = ~new_P3_SUB_485_U23 | ~new_P3_SUB_485_U7;
  assign new_P3_SUB_563_U6 = ~new_P3_U3305;
  assign new_P3_SUB_563_U7 = ~new_P3_U3306;
  assign new_P3_ADD_515_U4 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_515_U5 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_515_U6 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_515_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_515_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_515_U94;
  assign new_P3_ADD_515_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_515_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_515_U95;
  assign new_P3_ADD_515_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_515_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_515_U96;
  assign new_P3_ADD_515_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_515_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_515_U97;
  assign new_P3_ADD_515_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_515_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_515_U98;
  assign new_P3_ADD_515_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_515_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_515_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_515_U99;
  assign new_P3_ADD_515_U20 = ~new_P3_ADD_515_U100 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_515_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_515_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_515_U101;
  assign new_P3_ADD_515_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_515_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_515_U102;
  assign new_P3_ADD_515_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_515_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_515_U103;
  assign new_P3_ADD_515_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_515_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_515_U104;
  assign new_P3_ADD_515_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_515_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_515_U105;
  assign new_P3_ADD_515_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_515_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_515_U106;
  assign new_P3_ADD_515_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_515_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_515_U107;
  assign new_P3_ADD_515_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_515_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_515_U108;
  assign new_P3_ADD_515_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_515_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_515_U109;
  assign new_P3_ADD_515_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_515_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_515_U110;
  assign new_P3_ADD_515_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_515_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_515_U111;
  assign new_P3_ADD_515_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_515_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_515_U112;
  assign new_P3_ADD_515_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_515_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_515_U113;
  assign new_P3_ADD_515_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_515_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_515_U114;
  assign new_P3_ADD_515_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_515_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_515_U115;
  assign new_P3_ADD_515_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_515_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_515_U116;
  assign new_P3_ADD_515_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_515_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_515_U117;
  assign new_P3_ADD_515_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_515_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_515_U118;
  assign new_P3_ADD_515_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_515_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_515_U119;
  assign new_P3_ADD_515_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_515_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_515_U120;
  assign new_P3_ADD_515_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_515_U62 = ~new_P3_ADD_515_U124 | ~new_P3_ADD_515_U123;
  assign new_P3_ADD_515_U63 = ~new_P3_ADD_515_U126 | ~new_P3_ADD_515_U125;
  assign new_P3_ADD_515_U64 = ~new_P3_ADD_515_U128 | ~new_P3_ADD_515_U127;
  assign new_P3_ADD_515_U65 = ~new_P3_ADD_515_U130 | ~new_P3_ADD_515_U129;
  assign new_P3_ADD_515_U66 = ~new_P3_ADD_515_U132 | ~new_P3_ADD_515_U131;
  assign new_P3_ADD_515_U67 = ~new_P3_ADD_515_U134 | ~new_P3_ADD_515_U133;
  assign new_P3_ADD_515_U68 = ~new_P3_ADD_515_U136 | ~new_P3_ADD_515_U135;
  assign new_P3_ADD_515_U69 = ~new_P3_ADD_515_U138 | ~new_P3_ADD_515_U137;
  assign new_P3_ADD_515_U70 = ~new_P3_ADD_515_U140 | ~new_P3_ADD_515_U139;
  assign new_P3_ADD_515_U71 = ~new_P3_ADD_515_U142 | ~new_P3_ADD_515_U141;
  assign new_P3_ADD_515_U72 = ~new_P3_ADD_515_U144 | ~new_P3_ADD_515_U143;
  assign new_P3_ADD_515_U73 = ~new_P3_ADD_515_U146 | ~new_P3_ADD_515_U145;
  assign new_P3_ADD_515_U74 = ~new_P3_ADD_515_U148 | ~new_P3_ADD_515_U147;
  assign new_P3_ADD_515_U75 = ~new_P3_ADD_515_U150 | ~new_P3_ADD_515_U149;
  assign new_P3_ADD_515_U76 = ~new_P3_ADD_515_U152 | ~new_P3_ADD_515_U151;
  assign new_P3_ADD_515_U77 = ~new_P3_ADD_515_U154 | ~new_P3_ADD_515_U153;
  assign new_P3_ADD_515_U78 = ~new_P3_ADD_515_U156 | ~new_P3_ADD_515_U155;
  assign new_P3_ADD_515_U79 = ~new_P3_ADD_515_U158 | ~new_P3_ADD_515_U157;
  assign new_P3_ADD_515_U80 = ~new_P3_ADD_515_U160 | ~new_P3_ADD_515_U159;
  assign new_P3_ADD_515_U81 = ~new_P3_ADD_515_U162 | ~new_P3_ADD_515_U161;
  assign new_P3_ADD_515_U82 = ~new_P3_ADD_515_U164 | ~new_P3_ADD_515_U163;
  assign new_P3_ADD_515_U83 = ~new_P3_ADD_515_U166 | ~new_P3_ADD_515_U165;
  assign new_P3_ADD_515_U84 = ~new_P3_ADD_515_U168 | ~new_P3_ADD_515_U167;
  assign new_P3_ADD_515_U85 = ~new_P3_ADD_515_U170 | ~new_P3_ADD_515_U169;
  assign new_P3_ADD_515_U86 = ~new_P3_ADD_515_U172 | ~new_P3_ADD_515_U171;
  assign new_P3_ADD_515_U87 = ~new_P3_ADD_515_U174 | ~new_P3_ADD_515_U173;
  assign new_P3_ADD_515_U88 = ~new_P3_ADD_515_U176 | ~new_P3_ADD_515_U175;
  assign new_P3_ADD_515_U89 = ~new_P3_ADD_515_U178 | ~new_P3_ADD_515_U177;
  assign new_P3_ADD_515_U90 = ~new_P3_ADD_515_U180 | ~new_P3_ADD_515_U179;
  assign new_P3_ADD_515_U91 = ~new_P3_ADD_515_U182 | ~new_P3_ADD_515_U181;
  assign new_P3_ADD_515_U92 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_515_U93 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_515_U121;
  assign new_P3_ADD_515_U94 = ~new_P3_ADD_515_U6;
  assign new_P3_ADD_515_U95 = ~new_P3_ADD_515_U8;
  assign new_P3_ADD_515_U96 = ~new_P3_ADD_515_U10;
  assign new_P3_ADD_515_U97 = ~new_P3_ADD_515_U12;
  assign new_P3_ADD_515_U98 = ~new_P3_ADD_515_U14;
  assign new_P3_ADD_515_U99 = ~new_P3_ADD_515_U16;
  assign new_P3_ADD_515_U100 = ~new_P3_ADD_515_U19;
  assign new_P3_ADD_515_U101 = ~new_P3_ADD_515_U20;
  assign new_P3_ADD_515_U102 = ~new_P3_ADD_515_U22;
  assign new_P3_ADD_515_U103 = ~new_P3_ADD_515_U24;
  assign new_P3_ADD_515_U104 = ~new_P3_ADD_515_U26;
  assign new_P3_ADD_515_U105 = ~new_P3_ADD_515_U28;
  assign new_P3_ADD_515_U106 = ~new_P3_ADD_515_U30;
  assign new_P3_ADD_515_U107 = ~new_P3_ADD_515_U32;
  assign new_P3_ADD_515_U108 = ~new_P3_ADD_515_U34;
  assign new_P3_ADD_515_U109 = ~new_P3_ADD_515_U36;
  assign new_P3_ADD_515_U110 = ~new_P3_ADD_515_U38;
  assign new_P3_ADD_515_U111 = ~new_P3_ADD_515_U40;
  assign new_P3_ADD_515_U112 = ~new_P3_ADD_515_U42;
  assign new_P3_ADD_515_U113 = ~new_P3_ADD_515_U44;
  assign new_P3_ADD_515_U114 = ~new_P3_ADD_515_U46;
  assign new_P3_ADD_515_U115 = ~new_P3_ADD_515_U48;
  assign new_P3_ADD_515_U116 = ~new_P3_ADD_515_U50;
  assign new_P3_ADD_515_U117 = ~new_P3_ADD_515_U52;
  assign new_P3_ADD_515_U118 = ~new_P3_ADD_515_U54;
  assign new_P3_ADD_515_U119 = ~new_P3_ADD_515_U56;
  assign new_P3_ADD_515_U120 = ~new_P3_ADD_515_U58;
  assign new_P3_ADD_515_U121 = ~new_P3_ADD_515_U60;
  assign new_P3_ADD_515_U122 = ~new_P3_ADD_515_U93;
  assign new_P3_ADD_515_U123 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_515_U19;
  assign new_P3_ADD_515_U124 = ~new_P3_ADD_515_U100 | ~new_P3_ADD_515_U18;
  assign new_P3_ADD_515_U125 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_515_U16;
  assign new_P3_ADD_515_U126 = ~new_P3_ADD_515_U99 | ~new_P3_ADD_515_U17;
  assign new_P3_ADD_515_U127 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_515_U14;
  assign new_P3_ADD_515_U128 = ~new_P3_ADD_515_U98 | ~new_P3_ADD_515_U15;
  assign new_P3_ADD_515_U129 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_515_U12;
  assign new_P3_ADD_515_U130 = ~new_P3_ADD_515_U97 | ~new_P3_ADD_515_U13;
  assign new_P3_ADD_515_U131 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_515_U10;
  assign new_P3_ADD_515_U132 = ~new_P3_ADD_515_U96 | ~new_P3_ADD_515_U11;
  assign new_P3_ADD_515_U133 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_515_U8;
  assign new_P3_ADD_515_U134 = ~new_P3_ADD_515_U95 | ~new_P3_ADD_515_U9;
  assign new_P3_ADD_515_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_515_U6;
  assign new_P3_ADD_515_U136 = ~new_P3_ADD_515_U94 | ~new_P3_ADD_515_U7;
  assign new_P3_ADD_515_U137 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_515_U93;
  assign new_P3_ADD_515_U138 = ~new_P3_ADD_515_U122 | ~new_P3_ADD_515_U92;
  assign new_P3_ADD_515_U139 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_515_U60;
  assign new_P3_ADD_515_U140 = ~new_P3_ADD_515_U121 | ~new_P3_ADD_515_U61;
  assign new_P3_ADD_515_U141 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_515_U4;
  assign new_P3_ADD_515_U142 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_515_U5;
  assign new_P3_ADD_515_U143 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_515_U58;
  assign new_P3_ADD_515_U144 = ~new_P3_ADD_515_U120 | ~new_P3_ADD_515_U59;
  assign new_P3_ADD_515_U145 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_515_U56;
  assign new_P3_ADD_515_U146 = ~new_P3_ADD_515_U119 | ~new_P3_ADD_515_U57;
  assign new_P3_ADD_515_U147 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_515_U54;
  assign new_P3_ADD_515_U148 = ~new_P3_ADD_515_U118 | ~new_P3_ADD_515_U55;
  assign new_P3_ADD_515_U149 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_515_U52;
  assign new_P3_ADD_515_U150 = ~new_P3_ADD_515_U117 | ~new_P3_ADD_515_U53;
  assign new_P3_ADD_515_U151 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_515_U50;
  assign new_P3_ADD_515_U152 = ~new_P3_ADD_515_U116 | ~new_P3_ADD_515_U51;
  assign new_P3_ADD_515_U153 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_515_U48;
  assign new_P3_ADD_515_U154 = ~new_P3_ADD_515_U115 | ~new_P3_ADD_515_U49;
  assign new_P3_ADD_515_U155 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_515_U46;
  assign new_P3_ADD_515_U156 = ~new_P3_ADD_515_U114 | ~new_P3_ADD_515_U47;
  assign new_P3_ADD_515_U157 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_515_U44;
  assign new_P3_ADD_515_U158 = ~new_P3_ADD_515_U113 | ~new_P3_ADD_515_U45;
  assign new_P3_ADD_515_U159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_515_U42;
  assign new_P3_ADD_515_U160 = ~new_P3_ADD_515_U112 | ~new_P3_ADD_515_U43;
  assign new_P3_ADD_515_U161 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_515_U40;
  assign new_P3_ADD_515_U162 = ~new_P3_ADD_515_U111 | ~new_P3_ADD_515_U41;
  assign new_P3_ADD_515_U163 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_515_U38;
  assign new_P3_ADD_515_U164 = ~new_P3_ADD_515_U110 | ~new_P3_ADD_515_U39;
  assign new_P3_ADD_515_U165 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_515_U36;
  assign new_P3_ADD_515_U166 = ~new_P3_ADD_515_U109 | ~new_P3_ADD_515_U37;
  assign new_P3_ADD_515_U167 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_515_U34;
  assign new_P3_ADD_515_U168 = ~new_P3_ADD_515_U108 | ~new_P3_ADD_515_U35;
  assign new_P3_ADD_515_U169 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_515_U32;
  assign new_P3_ADD_515_U170 = ~new_P3_ADD_515_U107 | ~new_P3_ADD_515_U33;
  assign new_P3_ADD_515_U171 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_515_U30;
  assign new_P3_ADD_515_U172 = ~new_P3_ADD_515_U106 | ~new_P3_ADD_515_U31;
  assign new_P3_ADD_515_U173 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_515_U28;
  assign new_P3_ADD_515_U174 = ~new_P3_ADD_515_U105 | ~new_P3_ADD_515_U29;
  assign new_P3_ADD_515_U175 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_515_U26;
  assign new_P3_ADD_515_U176 = ~new_P3_ADD_515_U104 | ~new_P3_ADD_515_U27;
  assign new_P3_ADD_515_U177 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_515_U24;
  assign new_P3_ADD_515_U178 = ~new_P3_ADD_515_U103 | ~new_P3_ADD_515_U25;
  assign new_P3_ADD_515_U179 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_515_U22;
  assign new_P3_ADD_515_U180 = ~new_P3_ADD_515_U102 | ~new_P3_ADD_515_U23;
  assign new_P3_ADD_515_U181 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_515_U20;
  assign new_P3_ADD_515_U182 = ~new_P3_ADD_515_U101 | ~new_P3_ADD_515_U21;
  assign new_P3_ADD_394_U4 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_394_U5 = ~new_P3_ADD_394_U92 | ~new_P3_ADD_394_U126;
  assign new_P3_ADD_394_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_394_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_394_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_394_U92;
  assign new_P3_ADD_394_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_394_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_394_U98;
  assign new_P3_ADD_394_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_394_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_394_U99;
  assign new_P3_ADD_394_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_394_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_394_U100;
  assign new_P3_ADD_394_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_394_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_394_U101;
  assign new_P3_ADD_394_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_394_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_394_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_394_U102;
  assign new_P3_ADD_394_U20 = ~new_P3_ADD_394_U103 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_394_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_394_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_394_U104;
  assign new_P3_ADD_394_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_394_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_394_U105;
  assign new_P3_ADD_394_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_394_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_394_U106;
  assign new_P3_ADD_394_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_394_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_394_U107;
  assign new_P3_ADD_394_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_394_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_394_U108;
  assign new_P3_ADD_394_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_394_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_394_U109;
  assign new_P3_ADD_394_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_394_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_394_U110;
  assign new_P3_ADD_394_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_394_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_394_U111;
  assign new_P3_ADD_394_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_394_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_394_U112;
  assign new_P3_ADD_394_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_394_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_394_U113;
  assign new_P3_ADD_394_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_394_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_394_U114;
  assign new_P3_ADD_394_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_394_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_394_U115;
  assign new_P3_ADD_394_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_394_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_394_U116;
  assign new_P3_ADD_394_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_394_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_394_U117;
  assign new_P3_ADD_394_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_394_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_394_U118;
  assign new_P3_ADD_394_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_394_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_394_U119;
  assign new_P3_ADD_394_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_394_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_394_U120;
  assign new_P3_ADD_394_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_394_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_394_U121;
  assign new_P3_ADD_394_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_394_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_394_U122;
  assign new_P3_ADD_394_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_394_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_394_U123;
  assign new_P3_ADD_394_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_394_U62 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_394_U63 = ~new_P3_ADD_394_U128 | ~new_P3_ADD_394_U127;
  assign new_P3_ADD_394_U64 = ~new_P3_ADD_394_U130 | ~new_P3_ADD_394_U129;
  assign new_P3_ADD_394_U65 = ~new_P3_ADD_394_U132 | ~new_P3_ADD_394_U131;
  assign new_P3_ADD_394_U66 = ~new_P3_ADD_394_U134 | ~new_P3_ADD_394_U133;
  assign new_P3_ADD_394_U67 = ~new_P3_ADD_394_U136 | ~new_P3_ADD_394_U135;
  assign new_P3_ADD_394_U68 = ~new_P3_ADD_394_U138 | ~new_P3_ADD_394_U137;
  assign new_P3_ADD_394_U69 = ~new_P3_ADD_394_U142 | ~new_P3_ADD_394_U141;
  assign new_P3_ADD_394_U70 = ~new_P3_ADD_394_U144 | ~new_P3_ADD_394_U143;
  assign new_P3_ADD_394_U71 = ~new_P3_ADD_394_U146 | ~new_P3_ADD_394_U145;
  assign new_P3_ADD_394_U72 = ~new_P3_ADD_394_U148 | ~new_P3_ADD_394_U147;
  assign new_P3_ADD_394_U73 = ~new_P3_ADD_394_U150 | ~new_P3_ADD_394_U149;
  assign new_P3_ADD_394_U74 = ~new_P3_ADD_394_U152 | ~new_P3_ADD_394_U151;
  assign new_P3_ADD_394_U75 = ~new_P3_ADD_394_U154 | ~new_P3_ADD_394_U153;
  assign new_P3_ADD_394_U76 = ~new_P3_ADD_394_U156 | ~new_P3_ADD_394_U155;
  assign new_P3_ADD_394_U77 = ~new_P3_ADD_394_U158 | ~new_P3_ADD_394_U157;
  assign new_P3_ADD_394_U78 = ~new_P3_ADD_394_U160 | ~new_P3_ADD_394_U159;
  assign new_P3_ADD_394_U79 = ~new_P3_ADD_394_U162 | ~new_P3_ADD_394_U161;
  assign new_P3_ADD_394_U80 = ~new_P3_ADD_394_U164 | ~new_P3_ADD_394_U163;
  assign new_P3_ADD_394_U81 = ~new_P3_ADD_394_U166 | ~new_P3_ADD_394_U165;
  assign new_P3_ADD_394_U82 = ~new_P3_ADD_394_U168 | ~new_P3_ADD_394_U167;
  assign new_P3_ADD_394_U83 = ~new_P3_ADD_394_U170 | ~new_P3_ADD_394_U169;
  assign new_P3_ADD_394_U84 = ~new_P3_ADD_394_U172 | ~new_P3_ADD_394_U171;
  assign new_P3_ADD_394_U85 = ~new_P3_ADD_394_U174 | ~new_P3_ADD_394_U173;
  assign new_P3_ADD_394_U86 = ~new_P3_ADD_394_U176 | ~new_P3_ADD_394_U175;
  assign new_P3_ADD_394_U87 = ~new_P3_ADD_394_U178 | ~new_P3_ADD_394_U177;
  assign new_P3_ADD_394_U88 = ~new_P3_ADD_394_U180 | ~new_P3_ADD_394_U179;
  assign new_P3_ADD_394_U89 = ~new_P3_ADD_394_U182 | ~new_P3_ADD_394_U181;
  assign new_P3_ADD_394_U90 = ~new_P3_ADD_394_U184 | ~new_P3_ADD_394_U183;
  assign new_P3_ADD_394_U91 = ~new_P3_ADD_394_U186 | ~new_P3_ADD_394_U185;
  assign new_P3_ADD_394_U92 = ~new_P3_ADD_394_U62 | ~new_P3_ADD_394_U96;
  assign new_P3_ADD_394_U93 = new_P3_ADD_394_U140 & new_P3_ADD_394_U139;
  assign new_P3_ADD_394_U94 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_394_U95 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_394_U124;
  assign new_P3_ADD_394_U96 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_394_U97 = ~new_P3_ADD_394_U92;
  assign new_P3_ADD_394_U98 = ~new_P3_ADD_394_U8;
  assign new_P3_ADD_394_U99 = ~new_P3_ADD_394_U10;
  assign new_P3_ADD_394_U100 = ~new_P3_ADD_394_U12;
  assign new_P3_ADD_394_U101 = ~new_P3_ADD_394_U14;
  assign new_P3_ADD_394_U102 = ~new_P3_ADD_394_U16;
  assign new_P3_ADD_394_U103 = ~new_P3_ADD_394_U19;
  assign new_P3_ADD_394_U104 = ~new_P3_ADD_394_U20;
  assign new_P3_ADD_394_U105 = ~new_P3_ADD_394_U22;
  assign new_P3_ADD_394_U106 = ~new_P3_ADD_394_U24;
  assign new_P3_ADD_394_U107 = ~new_P3_ADD_394_U26;
  assign new_P3_ADD_394_U108 = ~new_P3_ADD_394_U28;
  assign new_P3_ADD_394_U109 = ~new_P3_ADD_394_U30;
  assign new_P3_ADD_394_U110 = ~new_P3_ADD_394_U32;
  assign new_P3_ADD_394_U111 = ~new_P3_ADD_394_U34;
  assign new_P3_ADD_394_U112 = ~new_P3_ADD_394_U36;
  assign new_P3_ADD_394_U113 = ~new_P3_ADD_394_U38;
  assign new_P3_ADD_394_U114 = ~new_P3_ADD_394_U40;
  assign new_P3_ADD_394_U115 = ~new_P3_ADD_394_U42;
  assign new_P3_ADD_394_U116 = ~new_P3_ADD_394_U44;
  assign new_P3_ADD_394_U117 = ~new_P3_ADD_394_U46;
  assign new_P3_ADD_394_U118 = ~new_P3_ADD_394_U48;
  assign new_P3_ADD_394_U119 = ~new_P3_ADD_394_U50;
  assign new_P3_ADD_394_U120 = ~new_P3_ADD_394_U52;
  assign new_P3_ADD_394_U121 = ~new_P3_ADD_394_U54;
  assign new_P3_ADD_394_U122 = ~new_P3_ADD_394_U56;
  assign new_P3_ADD_394_U123 = ~new_P3_ADD_394_U58;
  assign new_P3_ADD_394_U124 = ~new_P3_ADD_394_U60;
  assign new_P3_ADD_394_U125 = ~new_P3_ADD_394_U95;
  assign new_P3_ADD_394_U126 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_394_U127 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_394_U19;
  assign new_P3_ADD_394_U128 = ~new_P3_ADD_394_U103 | ~new_P3_ADD_394_U18;
  assign new_P3_ADD_394_U129 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_394_U16;
  assign new_P3_ADD_394_U130 = ~new_P3_ADD_394_U102 | ~new_P3_ADD_394_U17;
  assign new_P3_ADD_394_U131 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_394_U14;
  assign new_P3_ADD_394_U132 = ~new_P3_ADD_394_U101 | ~new_P3_ADD_394_U15;
  assign new_P3_ADD_394_U133 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_394_U12;
  assign new_P3_ADD_394_U134 = ~new_P3_ADD_394_U100 | ~new_P3_ADD_394_U13;
  assign new_P3_ADD_394_U135 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_394_U10;
  assign new_P3_ADD_394_U136 = ~new_P3_ADD_394_U99 | ~new_P3_ADD_394_U11;
  assign new_P3_ADD_394_U137 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_394_U8;
  assign new_P3_ADD_394_U138 = ~new_P3_ADD_394_U98 | ~new_P3_ADD_394_U9;
  assign new_P3_ADD_394_U139 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_394_U92;
  assign new_P3_ADD_394_U140 = ~new_P3_ADD_394_U97 | ~new_P3_ADD_394_U7;
  assign new_P3_ADD_394_U141 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_394_U95;
  assign new_P3_ADD_394_U142 = ~new_P3_ADD_394_U125 | ~new_P3_ADD_394_U94;
  assign new_P3_ADD_394_U143 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_394_U60;
  assign new_P3_ADD_394_U144 = ~new_P3_ADD_394_U124 | ~new_P3_ADD_394_U61;
  assign new_P3_ADD_394_U145 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_394_U58;
  assign new_P3_ADD_394_U146 = ~new_P3_ADD_394_U123 | ~new_P3_ADD_394_U59;
  assign new_P3_ADD_394_U147 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_394_U56;
  assign new_P3_ADD_394_U148 = ~new_P3_ADD_394_U122 | ~new_P3_ADD_394_U57;
  assign new_P3_ADD_394_U149 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_394_U54;
  assign new_P3_ADD_394_U150 = ~new_P3_ADD_394_U121 | ~new_P3_ADD_394_U55;
  assign new_P3_ADD_394_U151 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_394_U52;
  assign new_P3_ADD_394_U152 = ~new_P3_ADD_394_U120 | ~new_P3_ADD_394_U53;
  assign new_P3_ADD_394_U153 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_394_U50;
  assign new_P3_ADD_394_U154 = ~new_P3_ADD_394_U119 | ~new_P3_ADD_394_U51;
  assign new_P3_ADD_394_U155 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_394_U48;
  assign new_P3_ADD_394_U156 = ~new_P3_ADD_394_U118 | ~new_P3_ADD_394_U49;
  assign new_P3_ADD_394_U157 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_394_U46;
  assign new_P3_ADD_394_U158 = ~new_P3_ADD_394_U117 | ~new_P3_ADD_394_U47;
  assign new_P3_ADD_394_U159 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_394_U44;
  assign new_P3_ADD_394_U160 = ~new_P3_ADD_394_U116 | ~new_P3_ADD_394_U45;
  assign new_P3_ADD_394_U161 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_394_U42;
  assign new_P3_ADD_394_U162 = ~new_P3_ADD_394_U115 | ~new_P3_ADD_394_U43;
  assign new_P3_ADD_394_U163 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_394_U40;
  assign new_P3_ADD_394_U164 = ~new_P3_ADD_394_U114 | ~new_P3_ADD_394_U41;
  assign new_P3_ADD_394_U165 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_394_U4;
  assign new_P3_ADD_394_U166 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_394_U6;
  assign new_P3_ADD_394_U167 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_394_U38;
  assign new_P3_ADD_394_U168 = ~new_P3_ADD_394_U113 | ~new_P3_ADD_394_U39;
  assign new_P3_ADD_394_U169 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_394_U36;
  assign new_P3_ADD_394_U170 = ~new_P3_ADD_394_U112 | ~new_P3_ADD_394_U37;
  assign new_P3_ADD_394_U171 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_394_U34;
  assign new_P3_ADD_394_U172 = ~new_P3_ADD_394_U111 | ~new_P3_ADD_394_U35;
  assign new_P3_ADD_394_U173 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_394_U32;
  assign new_P3_ADD_394_U174 = ~new_P3_ADD_394_U110 | ~new_P3_ADD_394_U33;
  assign new_P3_ADD_394_U175 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_394_U30;
  assign new_P3_ADD_394_U176 = ~new_P3_ADD_394_U109 | ~new_P3_ADD_394_U31;
  assign new_P3_ADD_394_U177 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_394_U28;
  assign new_P3_ADD_394_U178 = ~new_P3_ADD_394_U108 | ~new_P3_ADD_394_U29;
  assign new_P3_ADD_394_U179 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_394_U26;
  assign new_P3_ADD_394_U180 = ~new_P3_ADD_394_U107 | ~new_P3_ADD_394_U27;
  assign new_P3_ADD_394_U181 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_394_U24;
  assign new_P3_ADD_394_U182 = ~new_P3_ADD_394_U106 | ~new_P3_ADD_394_U25;
  assign new_P3_ADD_394_U183 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_394_U22;
  assign new_P3_ADD_394_U184 = ~new_P3_ADD_394_U105 | ~new_P3_ADD_394_U23;
  assign new_P3_ADD_394_U185 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_394_U20;
  assign new_P3_ADD_394_U186 = ~new_P3_ADD_394_U104 | ~new_P3_ADD_394_U21;
  assign new_P3_GTE_450_U6 = ~new_P3_SUB_450_U6 & ~new_P3_GTE_450_U7;
  assign new_P3_GTE_450_U7 = ~new_P3_SUB_450_U18 & ~new_P3_SUB_450_U19 & ~new_P3_SUB_450_U16 & ~new_P3_SUB_450_U17;
  assign new_P3_SUB_414_U6 = new_P3_SUB_414_U126 & new_P3_SUB_414_U28;
  assign new_P3_SUB_414_U7 = new_P3_SUB_414_U124 & new_P3_SUB_414_U29;
  assign new_P3_SUB_414_U8 = new_P3_SUB_414_U122 & new_P3_SUB_414_U30;
  assign new_P3_SUB_414_U9 = new_P3_SUB_414_U120 & new_P3_SUB_414_U31;
  assign new_P3_SUB_414_U10 = new_P3_SUB_414_U118 & new_P3_SUB_414_U32;
  assign new_P3_SUB_414_U11 = new_P3_SUB_414_U116 & new_P3_SUB_414_U33;
  assign new_P3_SUB_414_U12 = new_P3_SUB_414_U114 & new_P3_SUB_414_U34;
  assign new_P3_SUB_414_U13 = new_P3_SUB_414_U112 & new_P3_SUB_414_U35;
  assign new_P3_SUB_414_U14 = new_P3_SUB_414_U110 & new_P3_SUB_414_U36;
  assign new_P3_SUB_414_U15 = new_P3_SUB_414_U108 & new_P3_SUB_414_U37;
  assign new_P3_SUB_414_U16 = new_P3_SUB_414_U106 & new_P3_SUB_414_U38;
  assign new_P3_SUB_414_U17 = new_P3_SUB_414_U105 & new_P3_SUB_414_U21;
  assign new_P3_SUB_414_U18 = new_P3_SUB_414_U92 & new_P3_SUB_414_U22;
  assign new_P3_SUB_414_U19 = new_P3_SUB_414_U90 & new_P3_SUB_414_U23;
  assign new_P3_SUB_414_U20 = new_P3_SUB_414_U88 & new_P3_SUB_414_U24;
  assign new_P3_SUB_414_U21 = P3_EBX_REG_2_ | P3_EBX_REG_1_ | P3_EBX_REG_0_;
  assign new_P3_SUB_414_U22 = ~new_P3_SUB_414_U83 | ~new_P3_SUB_414_U27 | ~new_P3_SUB_414_U58;
  assign new_P3_SUB_414_U23 = ~new_P3_SUB_414_U84 | ~new_P3_SUB_414_U26 | ~new_P3_SUB_414_U56;
  assign new_P3_SUB_414_U24 = ~new_P3_SUB_414_U85 | ~new_P3_SUB_414_U25 | ~new_P3_SUB_414_U54;
  assign new_P3_SUB_414_U25 = ~P3_EBX_REG_8_;
  assign new_P3_SUB_414_U26 = ~P3_EBX_REG_6_;
  assign new_P3_SUB_414_U27 = ~P3_EBX_REG_4_;
  assign new_P3_SUB_414_U28 = ~new_P3_SUB_414_U86 | ~new_P3_SUB_414_U52 | ~new_P3_SUB_414_U49;
  assign new_P3_SUB_414_U29 = ~new_P3_SUB_414_U93 | ~new_P3_SUB_414_U48 | ~new_P3_SUB_414_U81;
  assign new_P3_SUB_414_U30 = ~new_P3_SUB_414_U94 | ~new_P3_SUB_414_U47 | ~new_P3_SUB_414_U79;
  assign new_P3_SUB_414_U31 = ~new_P3_SUB_414_U95 | ~new_P3_SUB_414_U46 | ~new_P3_SUB_414_U77;
  assign new_P3_SUB_414_U32 = ~new_P3_SUB_414_U96 | ~new_P3_SUB_414_U45 | ~new_P3_SUB_414_U75;
  assign new_P3_SUB_414_U33 = ~new_P3_SUB_414_U97 | ~new_P3_SUB_414_U44 | ~new_P3_SUB_414_U73;
  assign new_P3_SUB_414_U34 = ~new_P3_SUB_414_U98 | ~new_P3_SUB_414_U43 | ~new_P3_SUB_414_U69;
  assign new_P3_SUB_414_U35 = ~new_P3_SUB_414_U99 | ~new_P3_SUB_414_U42 | ~new_P3_SUB_414_U67;
  assign new_P3_SUB_414_U36 = ~new_P3_SUB_414_U100 | ~new_P3_SUB_414_U41 | ~new_P3_SUB_414_U65;
  assign new_P3_SUB_414_U37 = ~new_P3_SUB_414_U101 | ~new_P3_SUB_414_U40 | ~new_P3_SUB_414_U63;
  assign new_P3_SUB_414_U38 = ~new_P3_SUB_414_U102 | ~new_P3_SUB_414_U39;
  assign new_P3_SUB_414_U39 = ~P3_EBX_REG_29_;
  assign new_P3_SUB_414_U40 = ~P3_EBX_REG_28_;
  assign new_P3_SUB_414_U41 = ~P3_EBX_REG_26_;
  assign new_P3_SUB_414_U42 = ~P3_EBX_REG_24_;
  assign new_P3_SUB_414_U43 = ~P3_EBX_REG_22_;
  assign new_P3_SUB_414_U44 = ~P3_EBX_REG_20_;
  assign new_P3_SUB_414_U45 = ~P3_EBX_REG_18_;
  assign new_P3_SUB_414_U46 = ~P3_EBX_REG_16_;
  assign new_P3_SUB_414_U47 = ~P3_EBX_REG_14_;
  assign new_P3_SUB_414_U48 = ~P3_EBX_REG_12_;
  assign new_P3_SUB_414_U49 = ~P3_EBX_REG_10_;
  assign new_P3_SUB_414_U50 = ~new_P3_SUB_414_U149 | ~new_P3_SUB_414_U148;
  assign new_P3_SUB_414_U51 = ~new_P3_SUB_414_U137 | ~new_P3_SUB_414_U136;
  assign new_P3_SUB_414_U52 = ~P3_EBX_REG_9_;
  assign new_P3_SUB_414_U53 = new_P3_SUB_414_U129 & new_P3_SUB_414_U128;
  assign new_P3_SUB_414_U54 = ~P3_EBX_REG_7_;
  assign new_P3_SUB_414_U55 = new_P3_SUB_414_U131 & new_P3_SUB_414_U130;
  assign new_P3_SUB_414_U56 = ~P3_EBX_REG_5_;
  assign new_P3_SUB_414_U57 = new_P3_SUB_414_U133 & new_P3_SUB_414_U132;
  assign new_P3_SUB_414_U58 = ~P3_EBX_REG_3_;
  assign new_P3_SUB_414_U59 = new_P3_SUB_414_U135 & new_P3_SUB_414_U134;
  assign new_P3_SUB_414_U60 = ~P3_EBX_REG_31_;
  assign new_P3_SUB_414_U61 = ~P3_EBX_REG_30_;
  assign new_P3_SUB_414_U62 = new_P3_SUB_414_U139 & new_P3_SUB_414_U138;
  assign new_P3_SUB_414_U63 = ~P3_EBX_REG_27_;
  assign new_P3_SUB_414_U64 = new_P3_SUB_414_U141 & new_P3_SUB_414_U140;
  assign new_P3_SUB_414_U65 = ~P3_EBX_REG_25_;
  assign new_P3_SUB_414_U66 = new_P3_SUB_414_U143 & new_P3_SUB_414_U142;
  assign new_P3_SUB_414_U67 = ~P3_EBX_REG_23_;
  assign new_P3_SUB_414_U68 = new_P3_SUB_414_U145 & new_P3_SUB_414_U144;
  assign new_P3_SUB_414_U69 = ~P3_EBX_REG_21_;
  assign new_P3_SUB_414_U70 = new_P3_SUB_414_U147 & new_P3_SUB_414_U146;
  assign new_P3_SUB_414_U71 = ~P3_EBX_REG_1_;
  assign new_P3_SUB_414_U72 = ~P3_EBX_REG_0_;
  assign new_P3_SUB_414_U73 = ~P3_EBX_REG_19_;
  assign new_P3_SUB_414_U74 = new_P3_SUB_414_U151 & new_P3_SUB_414_U150;
  assign new_P3_SUB_414_U75 = ~P3_EBX_REG_17_;
  assign new_P3_SUB_414_U76 = new_P3_SUB_414_U153 & new_P3_SUB_414_U152;
  assign new_P3_SUB_414_U77 = ~P3_EBX_REG_15_;
  assign new_P3_SUB_414_U78 = new_P3_SUB_414_U155 & new_P3_SUB_414_U154;
  assign new_P3_SUB_414_U79 = ~P3_EBX_REG_13_;
  assign new_P3_SUB_414_U80 = new_P3_SUB_414_U157 & new_P3_SUB_414_U156;
  assign new_P3_SUB_414_U81 = ~P3_EBX_REG_11_;
  assign new_P3_SUB_414_U82 = new_P3_SUB_414_U159 & new_P3_SUB_414_U158;
  assign new_P3_SUB_414_U83 = ~new_P3_SUB_414_U21;
  assign new_P3_SUB_414_U84 = ~new_P3_SUB_414_U22;
  assign new_P3_SUB_414_U85 = ~new_P3_SUB_414_U23;
  assign new_P3_SUB_414_U86 = ~new_P3_SUB_414_U24;
  assign new_P3_SUB_414_U87 = ~new_P3_SUB_414_U85 | ~new_P3_SUB_414_U54;
  assign new_P3_SUB_414_U88 = ~P3_EBX_REG_8_ | ~new_P3_SUB_414_U87;
  assign new_P3_SUB_414_U89 = ~new_P3_SUB_414_U84 | ~new_P3_SUB_414_U56;
  assign new_P3_SUB_414_U90 = ~P3_EBX_REG_6_ | ~new_P3_SUB_414_U89;
  assign new_P3_SUB_414_U91 = ~new_P3_SUB_414_U83 | ~new_P3_SUB_414_U58;
  assign new_P3_SUB_414_U92 = ~P3_EBX_REG_4_ | ~new_P3_SUB_414_U91;
  assign new_P3_SUB_414_U93 = ~new_P3_SUB_414_U28;
  assign new_P3_SUB_414_U94 = ~new_P3_SUB_414_U29;
  assign new_P3_SUB_414_U95 = ~new_P3_SUB_414_U30;
  assign new_P3_SUB_414_U96 = ~new_P3_SUB_414_U31;
  assign new_P3_SUB_414_U97 = ~new_P3_SUB_414_U32;
  assign new_P3_SUB_414_U98 = ~new_P3_SUB_414_U33;
  assign new_P3_SUB_414_U99 = ~new_P3_SUB_414_U34;
  assign new_P3_SUB_414_U100 = ~new_P3_SUB_414_U35;
  assign new_P3_SUB_414_U101 = ~new_P3_SUB_414_U36;
  assign new_P3_SUB_414_U102 = ~new_P3_SUB_414_U37;
  assign new_P3_SUB_414_U103 = ~new_P3_SUB_414_U38;
  assign new_P3_SUB_414_U104 = P3_EBX_REG_1_ | P3_EBX_REG_0_;
  assign new_P3_SUB_414_U105 = ~P3_EBX_REG_2_ | ~new_P3_SUB_414_U104;
  assign new_P3_SUB_414_U106 = ~P3_EBX_REG_29_ | ~new_P3_SUB_414_U37;
  assign new_P3_SUB_414_U107 = ~new_P3_SUB_414_U101 | ~new_P3_SUB_414_U63;
  assign new_P3_SUB_414_U108 = ~P3_EBX_REG_28_ | ~new_P3_SUB_414_U107;
  assign new_P3_SUB_414_U109 = ~new_P3_SUB_414_U100 | ~new_P3_SUB_414_U65;
  assign new_P3_SUB_414_U110 = ~P3_EBX_REG_26_ | ~new_P3_SUB_414_U109;
  assign new_P3_SUB_414_U111 = ~new_P3_SUB_414_U99 | ~new_P3_SUB_414_U67;
  assign new_P3_SUB_414_U112 = ~P3_EBX_REG_24_ | ~new_P3_SUB_414_U111;
  assign new_P3_SUB_414_U113 = ~new_P3_SUB_414_U98 | ~new_P3_SUB_414_U69;
  assign new_P3_SUB_414_U114 = ~P3_EBX_REG_22_ | ~new_P3_SUB_414_U113;
  assign new_P3_SUB_414_U115 = ~new_P3_SUB_414_U97 | ~new_P3_SUB_414_U73;
  assign new_P3_SUB_414_U116 = ~P3_EBX_REG_20_ | ~new_P3_SUB_414_U115;
  assign new_P3_SUB_414_U117 = ~new_P3_SUB_414_U96 | ~new_P3_SUB_414_U75;
  assign new_P3_SUB_414_U118 = ~P3_EBX_REG_18_ | ~new_P3_SUB_414_U117;
  assign new_P3_SUB_414_U119 = ~new_P3_SUB_414_U95 | ~new_P3_SUB_414_U77;
  assign new_P3_SUB_414_U120 = ~P3_EBX_REG_16_ | ~new_P3_SUB_414_U119;
  assign new_P3_SUB_414_U121 = ~new_P3_SUB_414_U94 | ~new_P3_SUB_414_U79;
  assign new_P3_SUB_414_U122 = ~P3_EBX_REG_14_ | ~new_P3_SUB_414_U121;
  assign new_P3_SUB_414_U123 = ~new_P3_SUB_414_U93 | ~new_P3_SUB_414_U81;
  assign new_P3_SUB_414_U124 = ~P3_EBX_REG_12_ | ~new_P3_SUB_414_U123;
  assign new_P3_SUB_414_U125 = ~new_P3_SUB_414_U86 | ~new_P3_SUB_414_U52;
  assign new_P3_SUB_414_U126 = ~P3_EBX_REG_10_ | ~new_P3_SUB_414_U125;
  assign new_P3_SUB_414_U127 = ~new_P3_SUB_414_U103 | ~new_P3_SUB_414_U61;
  assign new_P3_SUB_414_U128 = ~P3_EBX_REG_9_ | ~new_P3_SUB_414_U24;
  assign new_P3_SUB_414_U129 = ~new_P3_SUB_414_U86 | ~new_P3_SUB_414_U52;
  assign new_P3_SUB_414_U130 = ~P3_EBX_REG_7_ | ~new_P3_SUB_414_U23;
  assign new_P3_SUB_414_U131 = ~new_P3_SUB_414_U85 | ~new_P3_SUB_414_U54;
  assign new_P3_SUB_414_U132 = ~P3_EBX_REG_5_ | ~new_P3_SUB_414_U22;
  assign new_P3_SUB_414_U133 = ~new_P3_SUB_414_U84 | ~new_P3_SUB_414_U56;
  assign new_P3_SUB_414_U134 = ~P3_EBX_REG_3_ | ~new_P3_SUB_414_U21;
  assign new_P3_SUB_414_U135 = ~new_P3_SUB_414_U83 | ~new_P3_SUB_414_U58;
  assign new_P3_SUB_414_U136 = ~new_P3_SUB_414_U127 | ~new_P3_SUB_414_U60;
  assign new_P3_SUB_414_U137 = ~P3_EBX_REG_31_ | ~new_P3_SUB_414_U103 | ~new_P3_SUB_414_U61;
  assign new_P3_SUB_414_U138 = ~P3_EBX_REG_30_ | ~new_P3_SUB_414_U38;
  assign new_P3_SUB_414_U139 = ~new_P3_SUB_414_U103 | ~new_P3_SUB_414_U61;
  assign new_P3_SUB_414_U140 = ~P3_EBX_REG_27_ | ~new_P3_SUB_414_U36;
  assign new_P3_SUB_414_U141 = ~new_P3_SUB_414_U101 | ~new_P3_SUB_414_U63;
  assign new_P3_SUB_414_U142 = ~P3_EBX_REG_25_ | ~new_P3_SUB_414_U35;
  assign new_P3_SUB_414_U143 = ~new_P3_SUB_414_U100 | ~new_P3_SUB_414_U65;
  assign new_P3_SUB_414_U144 = ~P3_EBX_REG_23_ | ~new_P3_SUB_414_U34;
  assign new_P3_SUB_414_U145 = ~new_P3_SUB_414_U99 | ~new_P3_SUB_414_U67;
  assign new_P3_SUB_414_U146 = ~P3_EBX_REG_21_ | ~new_P3_SUB_414_U33;
  assign new_P3_SUB_414_U147 = ~new_P3_SUB_414_U98 | ~new_P3_SUB_414_U69;
  assign new_P3_SUB_414_U148 = ~P3_EBX_REG_1_ | ~new_P3_SUB_414_U72;
  assign new_P3_SUB_414_U149 = ~P3_EBX_REG_0_ | ~new_P3_SUB_414_U71;
  assign new_P3_SUB_414_U150 = ~P3_EBX_REG_19_ | ~new_P3_SUB_414_U32;
  assign new_P3_SUB_414_U151 = ~new_P3_SUB_414_U97 | ~new_P3_SUB_414_U73;
  assign new_P3_SUB_414_U152 = ~P3_EBX_REG_17_ | ~new_P3_SUB_414_U31;
  assign new_P3_SUB_414_U153 = ~new_P3_SUB_414_U96 | ~new_P3_SUB_414_U75;
  assign new_P3_SUB_414_U154 = ~P3_EBX_REG_15_ | ~new_P3_SUB_414_U30;
  assign new_P3_SUB_414_U155 = ~new_P3_SUB_414_U95 | ~new_P3_SUB_414_U77;
  assign new_P3_SUB_414_U156 = ~P3_EBX_REG_13_ | ~new_P3_SUB_414_U29;
  assign new_P3_SUB_414_U157 = ~new_P3_SUB_414_U94 | ~new_P3_SUB_414_U79;
  assign new_P3_SUB_414_U158 = ~P3_EBX_REG_11_ | ~new_P3_SUB_414_U28;
  assign new_P3_SUB_414_U159 = ~new_P3_SUB_414_U93 | ~new_P3_SUB_414_U81;
  assign new_P3_ADD_441_U4 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_441_U5 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_441_U6 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_441_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_441_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_441_U94;
  assign new_P3_ADD_441_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_441_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_441_U95;
  assign new_P3_ADD_441_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_441_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_441_U96;
  assign new_P3_ADD_441_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_441_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_441_U97;
  assign new_P3_ADD_441_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_441_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_441_U98;
  assign new_P3_ADD_441_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_441_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_441_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_441_U99;
  assign new_P3_ADD_441_U20 = ~new_P3_ADD_441_U100 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_441_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_441_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_441_U101;
  assign new_P3_ADD_441_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_441_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_441_U102;
  assign new_P3_ADD_441_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_441_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_441_U103;
  assign new_P3_ADD_441_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_441_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_441_U104;
  assign new_P3_ADD_441_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_441_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_441_U105;
  assign new_P3_ADD_441_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_441_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_441_U106;
  assign new_P3_ADD_441_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_441_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_441_U107;
  assign new_P3_ADD_441_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_441_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_441_U108;
  assign new_P3_ADD_441_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_441_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_441_U109;
  assign new_P3_ADD_441_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_441_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_441_U110;
  assign new_P3_ADD_441_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_441_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_441_U111;
  assign new_P3_ADD_441_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_441_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_441_U112;
  assign new_P3_ADD_441_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_441_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_441_U113;
  assign new_P3_ADD_441_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_441_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_441_U114;
  assign new_P3_ADD_441_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_441_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_441_U115;
  assign new_P3_ADD_441_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_441_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_441_U116;
  assign new_P3_ADD_441_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_441_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_441_U117;
  assign new_P3_ADD_441_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_441_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_441_U118;
  assign new_P3_ADD_441_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_441_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_441_U119;
  assign new_P3_ADD_441_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_441_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_441_U120;
  assign new_P3_ADD_441_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_441_U62 = ~new_P3_ADD_441_U124 | ~new_P3_ADD_441_U123;
  assign new_P3_ADD_441_U63 = ~new_P3_ADD_441_U126 | ~new_P3_ADD_441_U125;
  assign new_P3_ADD_441_U64 = ~new_P3_ADD_441_U128 | ~new_P3_ADD_441_U127;
  assign new_P3_ADD_441_U65 = ~new_P3_ADD_441_U130 | ~new_P3_ADD_441_U129;
  assign new_P3_ADD_441_U66 = ~new_P3_ADD_441_U132 | ~new_P3_ADD_441_U131;
  assign new_P3_ADD_441_U67 = ~new_P3_ADD_441_U134 | ~new_P3_ADD_441_U133;
  assign new_P3_ADD_441_U68 = ~new_P3_ADD_441_U136 | ~new_P3_ADD_441_U135;
  assign new_P3_ADD_441_U69 = ~new_P3_ADD_441_U138 | ~new_P3_ADD_441_U137;
  assign new_P3_ADD_441_U70 = ~new_P3_ADD_441_U140 | ~new_P3_ADD_441_U139;
  assign new_P3_ADD_441_U71 = ~new_P3_ADD_441_U142 | ~new_P3_ADD_441_U141;
  assign new_P3_ADD_441_U72 = ~new_P3_ADD_441_U144 | ~new_P3_ADD_441_U143;
  assign new_P3_ADD_441_U73 = ~new_P3_ADD_441_U146 | ~new_P3_ADD_441_U145;
  assign new_P3_ADD_441_U74 = ~new_P3_ADD_441_U148 | ~new_P3_ADD_441_U147;
  assign new_P3_ADD_441_U75 = ~new_P3_ADD_441_U150 | ~new_P3_ADD_441_U149;
  assign new_P3_ADD_441_U76 = ~new_P3_ADD_441_U152 | ~new_P3_ADD_441_U151;
  assign new_P3_ADD_441_U77 = ~new_P3_ADD_441_U154 | ~new_P3_ADD_441_U153;
  assign new_P3_ADD_441_U78 = ~new_P3_ADD_441_U156 | ~new_P3_ADD_441_U155;
  assign new_P3_ADD_441_U79 = ~new_P3_ADD_441_U158 | ~new_P3_ADD_441_U157;
  assign new_P3_ADD_441_U80 = ~new_P3_ADD_441_U160 | ~new_P3_ADD_441_U159;
  assign new_P3_ADD_441_U81 = ~new_P3_ADD_441_U162 | ~new_P3_ADD_441_U161;
  assign new_P3_ADD_441_U82 = ~new_P3_ADD_441_U164 | ~new_P3_ADD_441_U163;
  assign new_P3_ADD_441_U83 = ~new_P3_ADD_441_U166 | ~new_P3_ADD_441_U165;
  assign new_P3_ADD_441_U84 = ~new_P3_ADD_441_U168 | ~new_P3_ADD_441_U167;
  assign new_P3_ADD_441_U85 = ~new_P3_ADD_441_U170 | ~new_P3_ADD_441_U169;
  assign new_P3_ADD_441_U86 = ~new_P3_ADD_441_U172 | ~new_P3_ADD_441_U171;
  assign new_P3_ADD_441_U87 = ~new_P3_ADD_441_U174 | ~new_P3_ADD_441_U173;
  assign new_P3_ADD_441_U88 = ~new_P3_ADD_441_U176 | ~new_P3_ADD_441_U175;
  assign new_P3_ADD_441_U89 = ~new_P3_ADD_441_U178 | ~new_P3_ADD_441_U177;
  assign new_P3_ADD_441_U90 = ~new_P3_ADD_441_U180 | ~new_P3_ADD_441_U179;
  assign new_P3_ADD_441_U91 = ~new_P3_ADD_441_U182 | ~new_P3_ADD_441_U181;
  assign new_P3_ADD_441_U92 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_441_U93 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_441_U121;
  assign new_P3_ADD_441_U94 = ~new_P3_ADD_441_U6;
  assign new_P3_ADD_441_U95 = ~new_P3_ADD_441_U8;
  assign new_P3_ADD_441_U96 = ~new_P3_ADD_441_U10;
  assign new_P3_ADD_441_U97 = ~new_P3_ADD_441_U12;
  assign new_P3_ADD_441_U98 = ~new_P3_ADD_441_U14;
  assign new_P3_ADD_441_U99 = ~new_P3_ADD_441_U16;
  assign new_P3_ADD_441_U100 = ~new_P3_ADD_441_U19;
  assign new_P3_ADD_441_U101 = ~new_P3_ADD_441_U20;
  assign new_P3_ADD_441_U102 = ~new_P3_ADD_441_U22;
  assign new_P3_ADD_441_U103 = ~new_P3_ADD_441_U24;
  assign new_P3_ADD_441_U104 = ~new_P3_ADD_441_U26;
  assign new_P3_ADD_441_U105 = ~new_P3_ADD_441_U28;
  assign new_P3_ADD_441_U106 = ~new_P3_ADD_441_U30;
  assign new_P3_ADD_441_U107 = ~new_P3_ADD_441_U32;
  assign new_P3_ADD_441_U108 = ~new_P3_ADD_441_U34;
  assign new_P3_ADD_441_U109 = ~new_P3_ADD_441_U36;
  assign new_P3_ADD_441_U110 = ~new_P3_ADD_441_U38;
  assign new_P3_ADD_441_U111 = ~new_P3_ADD_441_U40;
  assign new_P3_ADD_441_U112 = ~new_P3_ADD_441_U42;
  assign new_P3_ADD_441_U113 = ~new_P3_ADD_441_U44;
  assign new_P3_ADD_441_U114 = ~new_P3_ADD_441_U46;
  assign new_P3_ADD_441_U115 = ~new_P3_ADD_441_U48;
  assign new_P3_ADD_441_U116 = ~new_P3_ADD_441_U50;
  assign new_P3_ADD_441_U117 = ~new_P3_ADD_441_U52;
  assign new_P3_ADD_441_U118 = ~new_P3_ADD_441_U54;
  assign new_P3_ADD_441_U119 = ~new_P3_ADD_441_U56;
  assign new_P3_ADD_441_U120 = ~new_P3_ADD_441_U58;
  assign new_P3_ADD_441_U121 = ~new_P3_ADD_441_U60;
  assign new_P3_ADD_441_U122 = ~new_P3_ADD_441_U93;
  assign new_P3_ADD_441_U123 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_441_U19;
  assign new_P3_ADD_441_U124 = ~new_P3_ADD_441_U100 | ~new_P3_ADD_441_U18;
  assign new_P3_ADD_441_U125 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_441_U16;
  assign new_P3_ADD_441_U126 = ~new_P3_ADD_441_U99 | ~new_P3_ADD_441_U17;
  assign new_P3_ADD_441_U127 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_441_U14;
  assign new_P3_ADD_441_U128 = ~new_P3_ADD_441_U98 | ~new_P3_ADD_441_U15;
  assign new_P3_ADD_441_U129 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_441_U12;
  assign new_P3_ADD_441_U130 = ~new_P3_ADD_441_U97 | ~new_P3_ADD_441_U13;
  assign new_P3_ADD_441_U131 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_441_U10;
  assign new_P3_ADD_441_U132 = ~new_P3_ADD_441_U96 | ~new_P3_ADD_441_U11;
  assign new_P3_ADD_441_U133 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_441_U8;
  assign new_P3_ADD_441_U134 = ~new_P3_ADD_441_U95 | ~new_P3_ADD_441_U9;
  assign new_P3_ADD_441_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_441_U6;
  assign new_P3_ADD_441_U136 = ~new_P3_ADD_441_U94 | ~new_P3_ADD_441_U7;
  assign new_P3_ADD_441_U137 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_441_U93;
  assign new_P3_ADD_441_U138 = ~new_P3_ADD_441_U122 | ~new_P3_ADD_441_U92;
  assign new_P3_ADD_441_U139 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_441_U60;
  assign new_P3_ADD_441_U140 = ~new_P3_ADD_441_U121 | ~new_P3_ADD_441_U61;
  assign new_P3_ADD_441_U141 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_441_U4;
  assign new_P3_ADD_441_U142 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_441_U5;
  assign new_P3_ADD_441_U143 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_441_U58;
  assign new_P3_ADD_441_U144 = ~new_P3_ADD_441_U120 | ~new_P3_ADD_441_U59;
  assign new_P3_ADD_441_U145 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_441_U56;
  assign new_P3_ADD_441_U146 = ~new_P3_ADD_441_U119 | ~new_P3_ADD_441_U57;
  assign new_P3_ADD_441_U147 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_441_U54;
  assign new_P3_ADD_441_U148 = ~new_P3_ADD_441_U118 | ~new_P3_ADD_441_U55;
  assign new_P3_ADD_441_U149 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_441_U52;
  assign new_P3_ADD_441_U150 = ~new_P3_ADD_441_U117 | ~new_P3_ADD_441_U53;
  assign new_P3_ADD_441_U151 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_441_U50;
  assign new_P3_ADD_441_U152 = ~new_P3_ADD_441_U116 | ~new_P3_ADD_441_U51;
  assign new_P3_ADD_441_U153 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_441_U48;
  assign new_P3_ADD_441_U154 = ~new_P3_ADD_441_U115 | ~new_P3_ADD_441_U49;
  assign new_P3_ADD_441_U155 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_441_U46;
  assign new_P3_ADD_441_U156 = ~new_P3_ADD_441_U114 | ~new_P3_ADD_441_U47;
  assign new_P3_ADD_441_U157 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_441_U44;
  assign new_P3_ADD_441_U158 = ~new_P3_ADD_441_U113 | ~new_P3_ADD_441_U45;
  assign new_P3_ADD_441_U159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_441_U42;
  assign new_P3_ADD_441_U160 = ~new_P3_ADD_441_U112 | ~new_P3_ADD_441_U43;
  assign new_P3_ADD_441_U161 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_441_U40;
  assign new_P3_ADD_441_U162 = ~new_P3_ADD_441_U111 | ~new_P3_ADD_441_U41;
  assign new_P3_ADD_441_U163 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_441_U38;
  assign new_P3_ADD_441_U164 = ~new_P3_ADD_441_U110 | ~new_P3_ADD_441_U39;
  assign new_P3_ADD_441_U165 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_441_U36;
  assign new_P3_ADD_441_U166 = ~new_P3_ADD_441_U109 | ~new_P3_ADD_441_U37;
  assign new_P3_ADD_441_U167 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_441_U34;
  assign new_P3_ADD_441_U168 = ~new_P3_ADD_441_U108 | ~new_P3_ADD_441_U35;
  assign new_P3_ADD_441_U169 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_441_U32;
  assign new_P3_ADD_441_U170 = ~new_P3_ADD_441_U107 | ~new_P3_ADD_441_U33;
  assign new_P3_ADD_441_U171 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_441_U30;
  assign new_P3_ADD_441_U172 = ~new_P3_ADD_441_U106 | ~new_P3_ADD_441_U31;
  assign new_P3_ADD_441_U173 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_441_U28;
  assign new_P3_ADD_441_U174 = ~new_P3_ADD_441_U105 | ~new_P3_ADD_441_U29;
  assign new_P3_ADD_441_U175 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_441_U26;
  assign new_P3_ADD_441_U176 = ~new_P3_ADD_441_U104 | ~new_P3_ADD_441_U27;
  assign new_P3_ADD_441_U177 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_441_U24;
  assign new_P3_ADD_441_U178 = ~new_P3_ADD_441_U103 | ~new_P3_ADD_441_U25;
  assign new_P3_ADD_441_U179 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_441_U22;
  assign new_P3_ADD_441_U180 = ~new_P3_ADD_441_U102 | ~new_P3_ADD_441_U23;
  assign new_P3_ADD_441_U181 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_441_U20;
  assign new_P3_ADD_441_U182 = ~new_P3_ADD_441_U101 | ~new_P3_ADD_441_U21;
  assign new_P3_ADD_349_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_349_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_349_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_349_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_349_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_349_U98;
  assign new_P3_ADD_349_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_349_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_349_U99;
  assign new_P3_ADD_349_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_349_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_349_U100;
  assign new_P3_ADD_349_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_349_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_349_U101;
  assign new_P3_ADD_349_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_349_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_349_U102;
  assign new_P3_ADD_349_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_349_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_349_U103;
  assign new_P3_ADD_349_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_349_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_349_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_349_U104;
  assign new_P3_ADD_349_U23 = ~new_P3_ADD_349_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_349_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_349_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_349_U106;
  assign new_P3_ADD_349_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_349_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_349_U107;
  assign new_P3_ADD_349_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_349_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_349_U108;
  assign new_P3_ADD_349_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_349_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_349_U109;
  assign new_P3_ADD_349_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_349_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_349_U110;
  assign new_P3_ADD_349_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_349_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_349_U111;
  assign new_P3_ADD_349_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_349_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_349_U112;
  assign new_P3_ADD_349_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_349_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_349_U113;
  assign new_P3_ADD_349_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_349_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_349_U114;
  assign new_P3_ADD_349_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_349_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_349_U115;
  assign new_P3_ADD_349_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_349_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_349_U116;
  assign new_P3_ADD_349_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_349_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_349_U117;
  assign new_P3_ADD_349_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_349_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_349_U118;
  assign new_P3_ADD_349_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_349_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_349_U119;
  assign new_P3_ADD_349_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_349_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_349_U120;
  assign new_P3_ADD_349_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_349_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_349_U121;
  assign new_P3_ADD_349_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_349_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_349_U122;
  assign new_P3_ADD_349_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_349_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_349_U123;
  assign new_P3_ADD_349_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_349_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_349_U124;
  assign new_P3_ADD_349_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_349_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_349_U125;
  assign new_P3_ADD_349_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_349_U65 = ~new_P3_ADD_349_U129 | ~new_P3_ADD_349_U128;
  assign new_P3_ADD_349_U66 = ~new_P3_ADD_349_U131 | ~new_P3_ADD_349_U130;
  assign new_P3_ADD_349_U67 = ~new_P3_ADD_349_U133 | ~new_P3_ADD_349_U132;
  assign new_P3_ADD_349_U68 = ~new_P3_ADD_349_U135 | ~new_P3_ADD_349_U134;
  assign new_P3_ADD_349_U69 = ~new_P3_ADD_349_U137 | ~new_P3_ADD_349_U136;
  assign new_P3_ADD_349_U70 = ~new_P3_ADD_349_U139 | ~new_P3_ADD_349_U138;
  assign new_P3_ADD_349_U71 = ~new_P3_ADD_349_U141 | ~new_P3_ADD_349_U140;
  assign new_P3_ADD_349_U72 = ~new_P3_ADD_349_U143 | ~new_P3_ADD_349_U142;
  assign new_P3_ADD_349_U73 = ~new_P3_ADD_349_U145 | ~new_P3_ADD_349_U144;
  assign new_P3_ADD_349_U74 = ~new_P3_ADD_349_U147 | ~new_P3_ADD_349_U146;
  assign new_P3_ADD_349_U75 = ~new_P3_ADD_349_U149 | ~new_P3_ADD_349_U148;
  assign new_P3_ADD_349_U76 = ~new_P3_ADD_349_U151 | ~new_P3_ADD_349_U150;
  assign new_P3_ADD_349_U77 = ~new_P3_ADD_349_U153 | ~new_P3_ADD_349_U152;
  assign new_P3_ADD_349_U78 = ~new_P3_ADD_349_U155 | ~new_P3_ADD_349_U154;
  assign new_P3_ADD_349_U79 = ~new_P3_ADD_349_U157 | ~new_P3_ADD_349_U156;
  assign new_P3_ADD_349_U80 = ~new_P3_ADD_349_U159 | ~new_P3_ADD_349_U158;
  assign new_P3_ADD_349_U81 = ~new_P3_ADD_349_U161 | ~new_P3_ADD_349_U160;
  assign new_P3_ADD_349_U82 = ~new_P3_ADD_349_U163 | ~new_P3_ADD_349_U162;
  assign new_P3_ADD_349_U83 = ~new_P3_ADD_349_U165 | ~new_P3_ADD_349_U164;
  assign new_P3_ADD_349_U84 = ~new_P3_ADD_349_U167 | ~new_P3_ADD_349_U166;
  assign new_P3_ADD_349_U85 = ~new_P3_ADD_349_U169 | ~new_P3_ADD_349_U168;
  assign new_P3_ADD_349_U86 = ~new_P3_ADD_349_U171 | ~new_P3_ADD_349_U170;
  assign new_P3_ADD_349_U87 = ~new_P3_ADD_349_U173 | ~new_P3_ADD_349_U172;
  assign new_P3_ADD_349_U88 = ~new_P3_ADD_349_U175 | ~new_P3_ADD_349_U174;
  assign new_P3_ADD_349_U89 = ~new_P3_ADD_349_U177 | ~new_P3_ADD_349_U176;
  assign new_P3_ADD_349_U90 = ~new_P3_ADD_349_U179 | ~new_P3_ADD_349_U178;
  assign new_P3_ADD_349_U91 = ~new_P3_ADD_349_U181 | ~new_P3_ADD_349_U180;
  assign new_P3_ADD_349_U92 = ~new_P3_ADD_349_U183 | ~new_P3_ADD_349_U182;
  assign new_P3_ADD_349_U93 = ~new_P3_ADD_349_U185 | ~new_P3_ADD_349_U184;
  assign new_P3_ADD_349_U94 = ~new_P3_ADD_349_U187 | ~new_P3_ADD_349_U186;
  assign new_P3_ADD_349_U95 = ~new_P3_ADD_349_U189 | ~new_P3_ADD_349_U188;
  assign new_P3_ADD_349_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_349_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_349_U126;
  assign new_P3_ADD_349_U98 = ~new_P3_ADD_349_U7;
  assign new_P3_ADD_349_U99 = ~new_P3_ADD_349_U9;
  assign new_P3_ADD_349_U100 = ~new_P3_ADD_349_U11;
  assign new_P3_ADD_349_U101 = ~new_P3_ADD_349_U13;
  assign new_P3_ADD_349_U102 = ~new_P3_ADD_349_U15;
  assign new_P3_ADD_349_U103 = ~new_P3_ADD_349_U17;
  assign new_P3_ADD_349_U104 = ~new_P3_ADD_349_U19;
  assign new_P3_ADD_349_U105 = ~new_P3_ADD_349_U22;
  assign new_P3_ADD_349_U106 = ~new_P3_ADD_349_U23;
  assign new_P3_ADD_349_U107 = ~new_P3_ADD_349_U25;
  assign new_P3_ADD_349_U108 = ~new_P3_ADD_349_U27;
  assign new_P3_ADD_349_U109 = ~new_P3_ADD_349_U29;
  assign new_P3_ADD_349_U110 = ~new_P3_ADD_349_U31;
  assign new_P3_ADD_349_U111 = ~new_P3_ADD_349_U33;
  assign new_P3_ADD_349_U112 = ~new_P3_ADD_349_U35;
  assign new_P3_ADD_349_U113 = ~new_P3_ADD_349_U37;
  assign new_P3_ADD_349_U114 = ~new_P3_ADD_349_U39;
  assign new_P3_ADD_349_U115 = ~new_P3_ADD_349_U41;
  assign new_P3_ADD_349_U116 = ~new_P3_ADD_349_U43;
  assign new_P3_ADD_349_U117 = ~new_P3_ADD_349_U45;
  assign new_P3_ADD_349_U118 = ~new_P3_ADD_349_U47;
  assign new_P3_ADD_349_U119 = ~new_P3_ADD_349_U49;
  assign new_P3_ADD_349_U120 = ~new_P3_ADD_349_U51;
  assign new_P3_ADD_349_U121 = ~new_P3_ADD_349_U53;
  assign new_P3_ADD_349_U122 = ~new_P3_ADD_349_U55;
  assign new_P3_ADD_349_U123 = ~new_P3_ADD_349_U57;
  assign new_P3_ADD_349_U124 = ~new_P3_ADD_349_U59;
  assign new_P3_ADD_349_U125 = ~new_P3_ADD_349_U61;
  assign new_P3_ADD_349_U126 = ~new_P3_ADD_349_U63;
  assign new_P3_ADD_349_U127 = ~new_P3_ADD_349_U97;
  assign new_P3_ADD_349_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_349_U22;
  assign new_P3_ADD_349_U129 = ~new_P3_ADD_349_U105 | ~new_P3_ADD_349_U21;
  assign new_P3_ADD_349_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_349_U19;
  assign new_P3_ADD_349_U131 = ~new_P3_ADD_349_U104 | ~new_P3_ADD_349_U20;
  assign new_P3_ADD_349_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_349_U17;
  assign new_P3_ADD_349_U133 = ~new_P3_ADD_349_U103 | ~new_P3_ADD_349_U18;
  assign new_P3_ADD_349_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_349_U15;
  assign new_P3_ADD_349_U135 = ~new_P3_ADD_349_U102 | ~new_P3_ADD_349_U16;
  assign new_P3_ADD_349_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_349_U13;
  assign new_P3_ADD_349_U137 = ~new_P3_ADD_349_U101 | ~new_P3_ADD_349_U14;
  assign new_P3_ADD_349_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_349_U11;
  assign new_P3_ADD_349_U139 = ~new_P3_ADD_349_U100 | ~new_P3_ADD_349_U12;
  assign new_P3_ADD_349_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_349_U9;
  assign new_P3_ADD_349_U141 = ~new_P3_ADD_349_U99 | ~new_P3_ADD_349_U10;
  assign new_P3_ADD_349_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_349_U97;
  assign new_P3_ADD_349_U143 = ~new_P3_ADD_349_U127 | ~new_P3_ADD_349_U96;
  assign new_P3_ADD_349_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_349_U63;
  assign new_P3_ADD_349_U145 = ~new_P3_ADD_349_U126 | ~new_P3_ADD_349_U64;
  assign new_P3_ADD_349_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_349_U7;
  assign new_P3_ADD_349_U147 = ~new_P3_ADD_349_U98 | ~new_P3_ADD_349_U8;
  assign new_P3_ADD_349_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_349_U61;
  assign new_P3_ADD_349_U149 = ~new_P3_ADD_349_U125 | ~new_P3_ADD_349_U62;
  assign new_P3_ADD_349_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_349_U59;
  assign new_P3_ADD_349_U151 = ~new_P3_ADD_349_U124 | ~new_P3_ADD_349_U60;
  assign new_P3_ADD_349_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_349_U57;
  assign new_P3_ADD_349_U153 = ~new_P3_ADD_349_U123 | ~new_P3_ADD_349_U58;
  assign new_P3_ADD_349_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_349_U55;
  assign new_P3_ADD_349_U155 = ~new_P3_ADD_349_U122 | ~new_P3_ADD_349_U56;
  assign new_P3_ADD_349_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_349_U53;
  assign new_P3_ADD_349_U157 = ~new_P3_ADD_349_U121 | ~new_P3_ADD_349_U54;
  assign new_P3_ADD_349_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_349_U51;
  assign new_P3_ADD_349_U159 = ~new_P3_ADD_349_U120 | ~new_P3_ADD_349_U52;
  assign new_P3_ADD_349_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_349_U49;
  assign new_P3_ADD_349_U161 = ~new_P3_ADD_349_U119 | ~new_P3_ADD_349_U50;
  assign new_P3_ADD_349_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_349_U47;
  assign new_P3_ADD_349_U163 = ~new_P3_ADD_349_U118 | ~new_P3_ADD_349_U48;
  assign new_P3_ADD_349_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_349_U45;
  assign new_P3_ADD_349_U165 = ~new_P3_ADD_349_U117 | ~new_P3_ADD_349_U46;
  assign new_P3_ADD_349_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_349_U43;
  assign new_P3_ADD_349_U167 = ~new_P3_ADD_349_U116 | ~new_P3_ADD_349_U44;
  assign new_P3_ADD_349_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_349_U5;
  assign new_P3_ADD_349_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_349_U6;
  assign new_P3_ADD_349_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_349_U41;
  assign new_P3_ADD_349_U171 = ~new_P3_ADD_349_U115 | ~new_P3_ADD_349_U42;
  assign new_P3_ADD_349_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_349_U39;
  assign new_P3_ADD_349_U173 = ~new_P3_ADD_349_U114 | ~new_P3_ADD_349_U40;
  assign new_P3_ADD_349_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_349_U37;
  assign new_P3_ADD_349_U175 = ~new_P3_ADD_349_U113 | ~new_P3_ADD_349_U38;
  assign new_P3_ADD_349_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_349_U35;
  assign new_P3_ADD_349_U177 = ~new_P3_ADD_349_U112 | ~new_P3_ADD_349_U36;
  assign new_P3_ADD_349_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_349_U33;
  assign new_P3_ADD_349_U179 = ~new_P3_ADD_349_U111 | ~new_P3_ADD_349_U34;
  assign new_P3_ADD_349_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_349_U31;
  assign new_P3_ADD_349_U181 = ~new_P3_ADD_349_U110 | ~new_P3_ADD_349_U32;
  assign new_P3_ADD_349_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_349_U29;
  assign new_P3_ADD_349_U183 = ~new_P3_ADD_349_U109 | ~new_P3_ADD_349_U30;
  assign new_P3_ADD_349_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_349_U27;
  assign new_P3_ADD_349_U185 = ~new_P3_ADD_349_U108 | ~new_P3_ADD_349_U28;
  assign new_P3_ADD_349_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_349_U25;
  assign new_P3_ADD_349_U187 = ~new_P3_ADD_349_U107 | ~new_P3_ADD_349_U26;
  assign new_P3_ADD_349_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_349_U23;
  assign new_P3_ADD_349_U189 = ~new_P3_ADD_349_U106 | ~new_P3_ADD_349_U24;
  assign new_P3_ADD_405_U4 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_405_U5 = ~new_P3_ADD_405_U92 | ~new_P3_ADD_405_U126;
  assign new_P3_ADD_405_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_405_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_405_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_405_U92;
  assign new_P3_ADD_405_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_405_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_405_U98;
  assign new_P3_ADD_405_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_405_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_405_U99;
  assign new_P3_ADD_405_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_405_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_405_U100;
  assign new_P3_ADD_405_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_405_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_405_U101;
  assign new_P3_ADD_405_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_405_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_405_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_405_U102;
  assign new_P3_ADD_405_U20 = ~new_P3_ADD_405_U103 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_405_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_405_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_405_U104;
  assign new_P3_ADD_405_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_405_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_405_U105;
  assign new_P3_ADD_405_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_405_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_405_U106;
  assign new_P3_ADD_405_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_405_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_405_U107;
  assign new_P3_ADD_405_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_405_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_405_U108;
  assign new_P3_ADD_405_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_405_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_405_U109;
  assign new_P3_ADD_405_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_405_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_405_U110;
  assign new_P3_ADD_405_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_405_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_405_U111;
  assign new_P3_ADD_405_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_405_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_405_U112;
  assign new_P3_ADD_405_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_405_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_405_U113;
  assign new_P3_ADD_405_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_405_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_405_U114;
  assign new_P3_ADD_405_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_405_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_405_U115;
  assign new_P3_ADD_405_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_405_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_405_U116;
  assign new_P3_ADD_405_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_405_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_405_U117;
  assign new_P3_ADD_405_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_405_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_405_U118;
  assign new_P3_ADD_405_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_405_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_405_U119;
  assign new_P3_ADD_405_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_405_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_405_U120;
  assign new_P3_ADD_405_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_405_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_405_U121;
  assign new_P3_ADD_405_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_405_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_405_U122;
  assign new_P3_ADD_405_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_405_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_405_U123;
  assign new_P3_ADD_405_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_405_U62 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_405_U63 = ~new_P3_ADD_405_U128 | ~new_P3_ADD_405_U127;
  assign new_P3_ADD_405_U64 = ~new_P3_ADD_405_U130 | ~new_P3_ADD_405_U129;
  assign new_P3_ADD_405_U65 = ~new_P3_ADD_405_U132 | ~new_P3_ADD_405_U131;
  assign new_P3_ADD_405_U66 = ~new_P3_ADD_405_U134 | ~new_P3_ADD_405_U133;
  assign new_P3_ADD_405_U67 = ~new_P3_ADD_405_U136 | ~new_P3_ADD_405_U135;
  assign new_P3_ADD_405_U68 = ~new_P3_ADD_405_U138 | ~new_P3_ADD_405_U137;
  assign new_P3_ADD_405_U69 = ~new_P3_ADD_405_U142 | ~new_P3_ADD_405_U141;
  assign new_P3_ADD_405_U70 = ~new_P3_ADD_405_U144 | ~new_P3_ADD_405_U143;
  assign new_P3_ADD_405_U71 = ~new_P3_ADD_405_U146 | ~new_P3_ADD_405_U145;
  assign new_P3_ADD_405_U72 = ~new_P3_ADD_405_U148 | ~new_P3_ADD_405_U147;
  assign new_P3_ADD_405_U73 = ~new_P3_ADD_405_U150 | ~new_P3_ADD_405_U149;
  assign new_P3_ADD_405_U74 = ~new_P3_ADD_405_U152 | ~new_P3_ADD_405_U151;
  assign new_P3_ADD_405_U75 = ~new_P3_ADD_405_U154 | ~new_P3_ADD_405_U153;
  assign new_P3_ADD_405_U76 = ~new_P3_ADD_405_U156 | ~new_P3_ADD_405_U155;
  assign new_P3_ADD_405_U77 = ~new_P3_ADD_405_U158 | ~new_P3_ADD_405_U157;
  assign new_P3_ADD_405_U78 = ~new_P3_ADD_405_U160 | ~new_P3_ADD_405_U159;
  assign new_P3_ADD_405_U79 = ~new_P3_ADD_405_U162 | ~new_P3_ADD_405_U161;
  assign new_P3_ADD_405_U80 = ~new_P3_ADD_405_U164 | ~new_P3_ADD_405_U163;
  assign new_P3_ADD_405_U81 = ~new_P3_ADD_405_U166 | ~new_P3_ADD_405_U165;
  assign new_P3_ADD_405_U82 = ~new_P3_ADD_405_U168 | ~new_P3_ADD_405_U167;
  assign new_P3_ADD_405_U83 = ~new_P3_ADD_405_U170 | ~new_P3_ADD_405_U169;
  assign new_P3_ADD_405_U84 = ~new_P3_ADD_405_U172 | ~new_P3_ADD_405_U171;
  assign new_P3_ADD_405_U85 = ~new_P3_ADD_405_U174 | ~new_P3_ADD_405_U173;
  assign new_P3_ADD_405_U86 = ~new_P3_ADD_405_U176 | ~new_P3_ADD_405_U175;
  assign new_P3_ADD_405_U87 = ~new_P3_ADD_405_U178 | ~new_P3_ADD_405_U177;
  assign new_P3_ADD_405_U88 = ~new_P3_ADD_405_U180 | ~new_P3_ADD_405_U179;
  assign new_P3_ADD_405_U89 = ~new_P3_ADD_405_U182 | ~new_P3_ADD_405_U181;
  assign new_P3_ADD_405_U90 = ~new_P3_ADD_405_U184 | ~new_P3_ADD_405_U183;
  assign new_P3_ADD_405_U91 = ~new_P3_ADD_405_U186 | ~new_P3_ADD_405_U185;
  assign new_P3_ADD_405_U92 = ~new_P3_ADD_405_U62 | ~new_P3_ADD_405_U96;
  assign new_P3_ADD_405_U93 = new_P3_ADD_405_U140 & new_P3_ADD_405_U139;
  assign new_P3_ADD_405_U94 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_405_U95 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_405_U124;
  assign new_P3_ADD_405_U96 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_405_U97 = ~new_P3_ADD_405_U92;
  assign new_P3_ADD_405_U98 = ~new_P3_ADD_405_U8;
  assign new_P3_ADD_405_U99 = ~new_P3_ADD_405_U10;
  assign new_P3_ADD_405_U100 = ~new_P3_ADD_405_U12;
  assign new_P3_ADD_405_U101 = ~new_P3_ADD_405_U14;
  assign new_P3_ADD_405_U102 = ~new_P3_ADD_405_U16;
  assign new_P3_ADD_405_U103 = ~new_P3_ADD_405_U19;
  assign new_P3_ADD_405_U104 = ~new_P3_ADD_405_U20;
  assign new_P3_ADD_405_U105 = ~new_P3_ADD_405_U22;
  assign new_P3_ADD_405_U106 = ~new_P3_ADD_405_U24;
  assign new_P3_ADD_405_U107 = ~new_P3_ADD_405_U26;
  assign new_P3_ADD_405_U108 = ~new_P3_ADD_405_U28;
  assign new_P3_ADD_405_U109 = ~new_P3_ADD_405_U30;
  assign new_P3_ADD_405_U110 = ~new_P3_ADD_405_U32;
  assign new_P3_ADD_405_U111 = ~new_P3_ADD_405_U34;
  assign new_P3_ADD_405_U112 = ~new_P3_ADD_405_U36;
  assign new_P3_ADD_405_U113 = ~new_P3_ADD_405_U38;
  assign new_P3_ADD_405_U114 = ~new_P3_ADD_405_U40;
  assign new_P3_ADD_405_U115 = ~new_P3_ADD_405_U42;
  assign new_P3_ADD_405_U116 = ~new_P3_ADD_405_U44;
  assign new_P3_ADD_405_U117 = ~new_P3_ADD_405_U46;
  assign new_P3_ADD_405_U118 = ~new_P3_ADD_405_U48;
  assign new_P3_ADD_405_U119 = ~new_P3_ADD_405_U50;
  assign new_P3_ADD_405_U120 = ~new_P3_ADD_405_U52;
  assign new_P3_ADD_405_U121 = ~new_P3_ADD_405_U54;
  assign new_P3_ADD_405_U122 = ~new_P3_ADD_405_U56;
  assign new_P3_ADD_405_U123 = ~new_P3_ADD_405_U58;
  assign new_P3_ADD_405_U124 = ~new_P3_ADD_405_U60;
  assign new_P3_ADD_405_U125 = ~new_P3_ADD_405_U95;
  assign new_P3_ADD_405_U126 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_405_U127 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_405_U19;
  assign new_P3_ADD_405_U128 = ~new_P3_ADD_405_U103 | ~new_P3_ADD_405_U18;
  assign new_P3_ADD_405_U129 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_405_U16;
  assign new_P3_ADD_405_U130 = ~new_P3_ADD_405_U102 | ~new_P3_ADD_405_U17;
  assign new_P3_ADD_405_U131 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_405_U14;
  assign new_P3_ADD_405_U132 = ~new_P3_ADD_405_U101 | ~new_P3_ADD_405_U15;
  assign new_P3_ADD_405_U133 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_405_U12;
  assign new_P3_ADD_405_U134 = ~new_P3_ADD_405_U100 | ~new_P3_ADD_405_U13;
  assign new_P3_ADD_405_U135 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_405_U10;
  assign new_P3_ADD_405_U136 = ~new_P3_ADD_405_U99 | ~new_P3_ADD_405_U11;
  assign new_P3_ADD_405_U137 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_405_U8;
  assign new_P3_ADD_405_U138 = ~new_P3_ADD_405_U98 | ~new_P3_ADD_405_U9;
  assign new_P3_ADD_405_U139 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_405_U92;
  assign new_P3_ADD_405_U140 = ~new_P3_ADD_405_U97 | ~new_P3_ADD_405_U7;
  assign new_P3_ADD_405_U141 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_405_U95;
  assign new_P3_ADD_405_U142 = ~new_P3_ADD_405_U125 | ~new_P3_ADD_405_U94;
  assign new_P3_ADD_405_U143 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_405_U60;
  assign new_P3_ADD_405_U144 = ~new_P3_ADD_405_U124 | ~new_P3_ADD_405_U61;
  assign new_P3_ADD_405_U145 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_405_U58;
  assign new_P3_ADD_405_U146 = ~new_P3_ADD_405_U123 | ~new_P3_ADD_405_U59;
  assign new_P3_ADD_405_U147 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_405_U56;
  assign new_P3_ADD_405_U148 = ~new_P3_ADD_405_U122 | ~new_P3_ADD_405_U57;
  assign new_P3_ADD_405_U149 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_405_U54;
  assign new_P3_ADD_405_U150 = ~new_P3_ADD_405_U121 | ~new_P3_ADD_405_U55;
  assign new_P3_ADD_405_U151 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_405_U52;
  assign new_P3_ADD_405_U152 = ~new_P3_ADD_405_U120 | ~new_P3_ADD_405_U53;
  assign new_P3_ADD_405_U153 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_405_U50;
  assign new_P3_ADD_405_U154 = ~new_P3_ADD_405_U119 | ~new_P3_ADD_405_U51;
  assign new_P3_ADD_405_U155 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_405_U48;
  assign new_P3_ADD_405_U156 = ~new_P3_ADD_405_U118 | ~new_P3_ADD_405_U49;
  assign new_P3_ADD_405_U157 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_405_U46;
  assign new_P3_ADD_405_U158 = ~new_P3_ADD_405_U117 | ~new_P3_ADD_405_U47;
  assign new_P3_ADD_405_U159 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_405_U44;
  assign new_P3_ADD_405_U160 = ~new_P3_ADD_405_U116 | ~new_P3_ADD_405_U45;
  assign new_P3_ADD_405_U161 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_405_U42;
  assign new_P3_ADD_405_U162 = ~new_P3_ADD_405_U115 | ~new_P3_ADD_405_U43;
  assign new_P3_ADD_405_U163 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_405_U40;
  assign new_P3_ADD_405_U164 = ~new_P3_ADD_405_U114 | ~new_P3_ADD_405_U41;
  assign new_P3_ADD_405_U165 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_405_U4;
  assign new_P3_ADD_405_U166 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_405_U6;
  assign new_P3_ADD_405_U167 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_405_U38;
  assign new_P3_ADD_405_U168 = ~new_P3_ADD_405_U113 | ~new_P3_ADD_405_U39;
  assign new_P3_ADD_405_U169 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_405_U36;
  assign new_P3_ADD_405_U170 = ~new_P3_ADD_405_U112 | ~new_P3_ADD_405_U37;
  assign new_P3_ADD_405_U171 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_405_U34;
  assign new_P3_ADD_405_U172 = ~new_P3_ADD_405_U111 | ~new_P3_ADD_405_U35;
  assign new_P3_ADD_405_U173 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_405_U32;
  assign new_P3_ADD_405_U174 = ~new_P3_ADD_405_U110 | ~new_P3_ADD_405_U33;
  assign new_P3_ADD_405_U175 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_405_U30;
  assign new_P3_ADD_405_U176 = ~new_P3_ADD_405_U109 | ~new_P3_ADD_405_U31;
  assign new_P3_ADD_405_U177 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_405_U28;
  assign new_P3_ADD_405_U178 = ~new_P3_ADD_405_U108 | ~new_P3_ADD_405_U29;
  assign new_P3_ADD_405_U179 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_405_U26;
  assign new_P3_ADD_405_U180 = ~new_P3_ADD_405_U107 | ~new_P3_ADD_405_U27;
  assign new_P3_ADD_405_U181 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_405_U24;
  assign new_P3_ADD_405_U182 = ~new_P3_ADD_405_U106 | ~new_P3_ADD_405_U25;
  assign new_P3_ADD_405_U183 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_405_U22;
  assign new_P3_ADD_405_U184 = ~new_P3_ADD_405_U105 | ~new_P3_ADD_405_U23;
  assign new_P3_ADD_405_U185 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_405_U20;
  assign new_P3_ADD_405_U186 = ~new_P3_ADD_405_U104 | ~new_P3_ADD_405_U21;
  assign new_P3_ADD_553_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_553_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_553_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_553_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_553_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_553_U98;
  assign new_P3_ADD_553_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_553_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_553_U99;
  assign new_P3_ADD_553_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_553_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_553_U100;
  assign new_P3_ADD_553_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_553_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_553_U101;
  assign new_P3_ADD_553_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_553_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_553_U102;
  assign new_P3_ADD_553_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_553_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_553_U103;
  assign new_P3_ADD_553_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_553_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_553_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_553_U104;
  assign new_P3_ADD_553_U23 = ~new_P3_ADD_553_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_553_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_553_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_553_U106;
  assign new_P3_ADD_553_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_553_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_553_U107;
  assign new_P3_ADD_553_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_553_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_553_U108;
  assign new_P3_ADD_553_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_553_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_553_U109;
  assign new_P3_ADD_553_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_553_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_553_U110;
  assign new_P3_ADD_553_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_553_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_553_U111;
  assign new_P3_ADD_553_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_553_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_553_U112;
  assign new_P3_ADD_553_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_553_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_553_U113;
  assign new_P3_ADD_553_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_553_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_553_U114;
  assign new_P3_ADD_553_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_553_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_553_U115;
  assign new_P3_ADD_553_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_553_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_553_U116;
  assign new_P3_ADD_553_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_553_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_553_U117;
  assign new_P3_ADD_553_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_553_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_553_U118;
  assign new_P3_ADD_553_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_553_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_553_U119;
  assign new_P3_ADD_553_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_553_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_553_U120;
  assign new_P3_ADD_553_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_553_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_553_U121;
  assign new_P3_ADD_553_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_553_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_553_U122;
  assign new_P3_ADD_553_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_553_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_553_U123;
  assign new_P3_ADD_553_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_553_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_553_U124;
  assign new_P3_ADD_553_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_553_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_553_U125;
  assign new_P3_ADD_553_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_553_U65 = ~new_P3_ADD_553_U129 | ~new_P3_ADD_553_U128;
  assign new_P3_ADD_553_U66 = ~new_P3_ADD_553_U131 | ~new_P3_ADD_553_U130;
  assign new_P3_ADD_553_U67 = ~new_P3_ADD_553_U133 | ~new_P3_ADD_553_U132;
  assign new_P3_ADD_553_U68 = ~new_P3_ADD_553_U135 | ~new_P3_ADD_553_U134;
  assign new_P3_ADD_553_U69 = ~new_P3_ADD_553_U137 | ~new_P3_ADD_553_U136;
  assign new_P3_ADD_553_U70 = ~new_P3_ADD_553_U139 | ~new_P3_ADD_553_U138;
  assign new_P3_ADD_553_U71 = ~new_P3_ADD_553_U141 | ~new_P3_ADD_553_U140;
  assign new_P3_ADD_553_U72 = ~new_P3_ADD_553_U143 | ~new_P3_ADD_553_U142;
  assign new_P3_ADD_553_U73 = ~new_P3_ADD_553_U145 | ~new_P3_ADD_553_U144;
  assign new_P3_ADD_553_U74 = ~new_P3_ADD_553_U147 | ~new_P3_ADD_553_U146;
  assign new_P3_ADD_553_U75 = ~new_P3_ADD_553_U149 | ~new_P3_ADD_553_U148;
  assign new_P3_ADD_553_U76 = ~new_P3_ADD_553_U151 | ~new_P3_ADD_553_U150;
  assign new_P3_ADD_553_U77 = ~new_P3_ADD_553_U153 | ~new_P3_ADD_553_U152;
  assign new_P3_ADD_553_U78 = ~new_P3_ADD_553_U155 | ~new_P3_ADD_553_U154;
  assign new_P3_ADD_553_U79 = ~new_P3_ADD_553_U157 | ~new_P3_ADD_553_U156;
  assign new_P3_ADD_553_U80 = ~new_P3_ADD_553_U159 | ~new_P3_ADD_553_U158;
  assign new_P3_ADD_553_U81 = ~new_P3_ADD_553_U161 | ~new_P3_ADD_553_U160;
  assign new_P3_ADD_553_U82 = ~new_P3_ADD_553_U163 | ~new_P3_ADD_553_U162;
  assign new_P3_ADD_553_U83 = ~new_P3_ADD_553_U165 | ~new_P3_ADD_553_U164;
  assign new_P3_ADD_553_U84 = ~new_P3_ADD_553_U167 | ~new_P3_ADD_553_U166;
  assign new_P3_ADD_553_U85 = ~new_P3_ADD_553_U169 | ~new_P3_ADD_553_U168;
  assign new_P3_ADD_553_U86 = ~new_P3_ADD_553_U171 | ~new_P3_ADD_553_U170;
  assign new_P3_ADD_553_U87 = ~new_P3_ADD_553_U173 | ~new_P3_ADD_553_U172;
  assign new_P3_ADD_553_U88 = ~new_P3_ADD_553_U175 | ~new_P3_ADD_553_U174;
  assign new_P3_ADD_553_U89 = ~new_P3_ADD_553_U177 | ~new_P3_ADD_553_U176;
  assign new_P3_ADD_553_U90 = ~new_P3_ADD_553_U179 | ~new_P3_ADD_553_U178;
  assign new_P3_ADD_553_U91 = ~new_P3_ADD_553_U181 | ~new_P3_ADD_553_U180;
  assign new_P3_ADD_553_U92 = ~new_P3_ADD_553_U183 | ~new_P3_ADD_553_U182;
  assign new_P3_ADD_553_U93 = ~new_P3_ADD_553_U185 | ~new_P3_ADD_553_U184;
  assign new_P3_ADD_553_U94 = ~new_P3_ADD_553_U187 | ~new_P3_ADD_553_U186;
  assign new_P3_ADD_553_U95 = ~new_P3_ADD_553_U189 | ~new_P3_ADD_553_U188;
  assign new_P3_ADD_553_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_553_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_553_U126;
  assign new_P3_ADD_553_U98 = ~new_P3_ADD_553_U7;
  assign new_P3_ADD_553_U99 = ~new_P3_ADD_553_U9;
  assign new_P3_ADD_553_U100 = ~new_P3_ADD_553_U11;
  assign new_P3_ADD_553_U101 = ~new_P3_ADD_553_U13;
  assign new_P3_ADD_553_U102 = ~new_P3_ADD_553_U15;
  assign new_P3_ADD_553_U103 = ~new_P3_ADD_553_U17;
  assign new_P3_ADD_553_U104 = ~new_P3_ADD_553_U19;
  assign new_P3_ADD_553_U105 = ~new_P3_ADD_553_U22;
  assign new_P3_ADD_553_U106 = ~new_P3_ADD_553_U23;
  assign new_P3_ADD_553_U107 = ~new_P3_ADD_553_U25;
  assign new_P3_ADD_553_U108 = ~new_P3_ADD_553_U27;
  assign new_P3_ADD_553_U109 = ~new_P3_ADD_553_U29;
  assign new_P3_ADD_553_U110 = ~new_P3_ADD_553_U31;
  assign new_P3_ADD_553_U111 = ~new_P3_ADD_553_U33;
  assign new_P3_ADD_553_U112 = ~new_P3_ADD_553_U35;
  assign new_P3_ADD_553_U113 = ~new_P3_ADD_553_U37;
  assign new_P3_ADD_553_U114 = ~new_P3_ADD_553_U39;
  assign new_P3_ADD_553_U115 = ~new_P3_ADD_553_U41;
  assign new_P3_ADD_553_U116 = ~new_P3_ADD_553_U43;
  assign new_P3_ADD_553_U117 = ~new_P3_ADD_553_U45;
  assign new_P3_ADD_553_U118 = ~new_P3_ADD_553_U47;
  assign new_P3_ADD_553_U119 = ~new_P3_ADD_553_U49;
  assign new_P3_ADD_553_U120 = ~new_P3_ADD_553_U51;
  assign new_P3_ADD_553_U121 = ~new_P3_ADD_553_U53;
  assign new_P3_ADD_553_U122 = ~new_P3_ADD_553_U55;
  assign new_P3_ADD_553_U123 = ~new_P3_ADD_553_U57;
  assign new_P3_ADD_553_U124 = ~new_P3_ADD_553_U59;
  assign new_P3_ADD_553_U125 = ~new_P3_ADD_553_U61;
  assign new_P3_ADD_553_U126 = ~new_P3_ADD_553_U63;
  assign new_P3_ADD_553_U127 = ~new_P3_ADD_553_U97;
  assign new_P3_ADD_553_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_553_U22;
  assign new_P3_ADD_553_U129 = ~new_P3_ADD_553_U105 | ~new_P3_ADD_553_U21;
  assign new_P3_ADD_553_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_553_U19;
  assign new_P3_ADD_553_U131 = ~new_P3_ADD_553_U104 | ~new_P3_ADD_553_U20;
  assign new_P3_ADD_553_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_553_U17;
  assign new_P3_ADD_553_U133 = ~new_P3_ADD_553_U103 | ~new_P3_ADD_553_U18;
  assign new_P3_ADD_553_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_553_U15;
  assign new_P3_ADD_553_U135 = ~new_P3_ADD_553_U102 | ~new_P3_ADD_553_U16;
  assign new_P3_ADD_553_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_553_U13;
  assign new_P3_ADD_553_U137 = ~new_P3_ADD_553_U101 | ~new_P3_ADD_553_U14;
  assign new_P3_ADD_553_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_553_U11;
  assign new_P3_ADD_553_U139 = ~new_P3_ADD_553_U100 | ~new_P3_ADD_553_U12;
  assign new_P3_ADD_553_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_553_U9;
  assign new_P3_ADD_553_U141 = ~new_P3_ADD_553_U99 | ~new_P3_ADD_553_U10;
  assign new_P3_ADD_553_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_553_U97;
  assign new_P3_ADD_553_U143 = ~new_P3_ADD_553_U127 | ~new_P3_ADD_553_U96;
  assign new_P3_ADD_553_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_553_U63;
  assign new_P3_ADD_553_U145 = ~new_P3_ADD_553_U126 | ~new_P3_ADD_553_U64;
  assign new_P3_ADD_553_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_553_U7;
  assign new_P3_ADD_553_U147 = ~new_P3_ADD_553_U98 | ~new_P3_ADD_553_U8;
  assign new_P3_ADD_553_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_553_U61;
  assign new_P3_ADD_553_U149 = ~new_P3_ADD_553_U125 | ~new_P3_ADD_553_U62;
  assign new_P3_ADD_553_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_553_U59;
  assign new_P3_ADD_553_U151 = ~new_P3_ADD_553_U124 | ~new_P3_ADD_553_U60;
  assign new_P3_ADD_553_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_553_U57;
  assign new_P3_ADD_553_U153 = ~new_P3_ADD_553_U123 | ~new_P3_ADD_553_U58;
  assign new_P3_ADD_553_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_553_U55;
  assign new_P3_ADD_553_U155 = ~new_P3_ADD_553_U122 | ~new_P3_ADD_553_U56;
  assign new_P3_ADD_553_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_553_U53;
  assign new_P3_ADD_553_U157 = ~new_P3_ADD_553_U121 | ~new_P3_ADD_553_U54;
  assign new_P3_ADD_553_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_553_U51;
  assign new_P3_ADD_553_U159 = ~new_P3_ADD_553_U120 | ~new_P3_ADD_553_U52;
  assign new_P3_ADD_553_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_553_U49;
  assign new_P3_ADD_553_U161 = ~new_P3_ADD_553_U119 | ~new_P3_ADD_553_U50;
  assign new_P3_ADD_553_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_553_U47;
  assign new_P3_ADD_553_U163 = ~new_P3_ADD_553_U118 | ~new_P3_ADD_553_U48;
  assign new_P3_ADD_553_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_553_U45;
  assign new_P3_ADD_553_U165 = ~new_P3_ADD_553_U117 | ~new_P3_ADD_553_U46;
  assign new_P3_ADD_553_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_553_U43;
  assign new_P3_ADD_553_U167 = ~new_P3_ADD_553_U116 | ~new_P3_ADD_553_U44;
  assign new_P3_ADD_553_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_553_U5;
  assign new_P3_ADD_553_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_553_U6;
  assign new_P3_ADD_553_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_553_U41;
  assign new_P3_ADD_553_U171 = ~new_P3_ADD_553_U115 | ~new_P3_ADD_553_U42;
  assign new_P3_ADD_553_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_553_U39;
  assign new_P3_ADD_553_U173 = ~new_P3_ADD_553_U114 | ~new_P3_ADD_553_U40;
  assign new_P3_ADD_553_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_553_U37;
  assign new_P3_ADD_553_U175 = ~new_P3_ADD_553_U113 | ~new_P3_ADD_553_U38;
  assign new_P3_ADD_553_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_553_U35;
  assign new_P3_ADD_553_U177 = ~new_P3_ADD_553_U112 | ~new_P3_ADD_553_U36;
  assign new_P3_ADD_553_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_553_U33;
  assign new_P3_ADD_553_U179 = ~new_P3_ADD_553_U111 | ~new_P3_ADD_553_U34;
  assign new_P3_ADD_553_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_553_U31;
  assign new_P3_ADD_553_U181 = ~new_P3_ADD_553_U110 | ~new_P3_ADD_553_U32;
  assign new_P3_ADD_553_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_553_U29;
  assign new_P3_ADD_553_U183 = ~new_P3_ADD_553_U109 | ~new_P3_ADD_553_U30;
  assign new_P3_ADD_553_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_553_U27;
  assign new_P3_ADD_553_U185 = ~new_P3_ADD_553_U108 | ~new_P3_ADD_553_U28;
  assign new_P3_ADD_553_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_553_U25;
  assign new_P3_ADD_553_U187 = ~new_P3_ADD_553_U107 | ~new_P3_ADD_553_U26;
  assign new_P3_ADD_553_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_553_U23;
  assign new_P3_ADD_553_U189 = ~new_P3_ADD_553_U106 | ~new_P3_ADD_553_U24;
  assign new_P3_ADD_558_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_558_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_558_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_558_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_558_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_558_U98;
  assign new_P3_ADD_558_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_558_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_558_U99;
  assign new_P3_ADD_558_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_558_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_558_U100;
  assign new_P3_ADD_558_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_558_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_558_U101;
  assign new_P3_ADD_558_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_558_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_558_U102;
  assign new_P3_ADD_558_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_558_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_558_U103;
  assign new_P3_ADD_558_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_558_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_558_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_558_U104;
  assign new_P3_ADD_558_U23 = ~new_P3_ADD_558_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_558_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_558_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_558_U106;
  assign new_P3_ADD_558_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_558_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_558_U107;
  assign new_P3_ADD_558_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_558_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_558_U108;
  assign new_P3_ADD_558_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_558_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_558_U109;
  assign new_P3_ADD_558_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_558_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_558_U110;
  assign new_P3_ADD_558_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_558_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_558_U111;
  assign new_P3_ADD_558_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_558_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_558_U112;
  assign new_P3_ADD_558_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_558_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_558_U113;
  assign new_P3_ADD_558_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_558_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_558_U114;
  assign new_P3_ADD_558_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_558_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_558_U115;
  assign new_P3_ADD_558_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_558_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_558_U116;
  assign new_P3_ADD_558_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_558_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_558_U117;
  assign new_P3_ADD_558_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_558_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_558_U118;
  assign new_P3_ADD_558_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_558_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_558_U119;
  assign new_P3_ADD_558_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_558_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_558_U120;
  assign new_P3_ADD_558_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_558_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_558_U121;
  assign new_P3_ADD_558_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_558_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_558_U122;
  assign new_P3_ADD_558_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_558_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_558_U123;
  assign new_P3_ADD_558_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_558_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_558_U124;
  assign new_P3_ADD_558_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_558_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_558_U125;
  assign new_P3_ADD_558_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_558_U65 = ~new_P3_ADD_558_U129 | ~new_P3_ADD_558_U128;
  assign new_P3_ADD_558_U66 = ~new_P3_ADD_558_U131 | ~new_P3_ADD_558_U130;
  assign new_P3_ADD_558_U67 = ~new_P3_ADD_558_U133 | ~new_P3_ADD_558_U132;
  assign new_P3_ADD_558_U68 = ~new_P3_ADD_558_U135 | ~new_P3_ADD_558_U134;
  assign new_P3_ADD_558_U69 = ~new_P3_ADD_558_U137 | ~new_P3_ADD_558_U136;
  assign new_P3_ADD_558_U70 = ~new_P3_ADD_558_U139 | ~new_P3_ADD_558_U138;
  assign new_P3_ADD_558_U71 = ~new_P3_ADD_558_U141 | ~new_P3_ADD_558_U140;
  assign new_P3_ADD_558_U72 = ~new_P3_ADD_558_U143 | ~new_P3_ADD_558_U142;
  assign new_P3_ADD_558_U73 = ~new_P3_ADD_558_U145 | ~new_P3_ADD_558_U144;
  assign new_P3_ADD_558_U74 = ~new_P3_ADD_558_U147 | ~new_P3_ADD_558_U146;
  assign new_P3_ADD_558_U75 = ~new_P3_ADD_558_U149 | ~new_P3_ADD_558_U148;
  assign new_P3_ADD_558_U76 = ~new_P3_ADD_558_U151 | ~new_P3_ADD_558_U150;
  assign new_P3_ADD_558_U77 = ~new_P3_ADD_558_U153 | ~new_P3_ADD_558_U152;
  assign new_P3_ADD_558_U78 = ~new_P3_ADD_558_U155 | ~new_P3_ADD_558_U154;
  assign new_P3_ADD_558_U79 = ~new_P3_ADD_558_U157 | ~new_P3_ADD_558_U156;
  assign new_P3_ADD_558_U80 = ~new_P3_ADD_558_U159 | ~new_P3_ADD_558_U158;
  assign new_P3_ADD_558_U81 = ~new_P3_ADD_558_U161 | ~new_P3_ADD_558_U160;
  assign new_P3_ADD_558_U82 = ~new_P3_ADD_558_U163 | ~new_P3_ADD_558_U162;
  assign new_P3_ADD_558_U83 = ~new_P3_ADD_558_U165 | ~new_P3_ADD_558_U164;
  assign new_P3_ADD_558_U84 = ~new_P3_ADD_558_U167 | ~new_P3_ADD_558_U166;
  assign new_P3_ADD_558_U85 = ~new_P3_ADD_558_U169 | ~new_P3_ADD_558_U168;
  assign new_P3_ADD_558_U86 = ~new_P3_ADD_558_U171 | ~new_P3_ADD_558_U170;
  assign new_P3_ADD_558_U87 = ~new_P3_ADD_558_U173 | ~new_P3_ADD_558_U172;
  assign new_P3_ADD_558_U88 = ~new_P3_ADD_558_U175 | ~new_P3_ADD_558_U174;
  assign new_P3_ADD_558_U89 = ~new_P3_ADD_558_U177 | ~new_P3_ADD_558_U176;
  assign new_P3_ADD_558_U90 = ~new_P3_ADD_558_U179 | ~new_P3_ADD_558_U178;
  assign new_P3_ADD_558_U91 = ~new_P3_ADD_558_U181 | ~new_P3_ADD_558_U180;
  assign new_P3_ADD_558_U92 = ~new_P3_ADD_558_U183 | ~new_P3_ADD_558_U182;
  assign new_P3_ADD_558_U93 = ~new_P3_ADD_558_U185 | ~new_P3_ADD_558_U184;
  assign new_P3_ADD_558_U94 = ~new_P3_ADD_558_U187 | ~new_P3_ADD_558_U186;
  assign new_P3_ADD_558_U95 = ~new_P3_ADD_558_U189 | ~new_P3_ADD_558_U188;
  assign new_P3_ADD_558_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_558_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_558_U126;
  assign new_P3_ADD_558_U98 = ~new_P3_ADD_558_U7;
  assign new_P3_ADD_558_U99 = ~new_P3_ADD_558_U9;
  assign new_P3_ADD_558_U100 = ~new_P3_ADD_558_U11;
  assign new_P3_ADD_558_U101 = ~new_P3_ADD_558_U13;
  assign new_P3_ADD_558_U102 = ~new_P3_ADD_558_U15;
  assign new_P3_ADD_558_U103 = ~new_P3_ADD_558_U17;
  assign new_P3_ADD_558_U104 = ~new_P3_ADD_558_U19;
  assign new_P3_ADD_558_U105 = ~new_P3_ADD_558_U22;
  assign new_P3_ADD_558_U106 = ~new_P3_ADD_558_U23;
  assign new_P3_ADD_558_U107 = ~new_P3_ADD_558_U25;
  assign new_P3_ADD_558_U108 = ~new_P3_ADD_558_U27;
  assign new_P3_ADD_558_U109 = ~new_P3_ADD_558_U29;
  assign new_P3_ADD_558_U110 = ~new_P3_ADD_558_U31;
  assign new_P3_ADD_558_U111 = ~new_P3_ADD_558_U33;
  assign new_P3_ADD_558_U112 = ~new_P3_ADD_558_U35;
  assign new_P3_ADD_558_U113 = ~new_P3_ADD_558_U37;
  assign new_P3_ADD_558_U114 = ~new_P3_ADD_558_U39;
  assign new_P3_ADD_558_U115 = ~new_P3_ADD_558_U41;
  assign new_P3_ADD_558_U116 = ~new_P3_ADD_558_U43;
  assign new_P3_ADD_558_U117 = ~new_P3_ADD_558_U45;
  assign new_P3_ADD_558_U118 = ~new_P3_ADD_558_U47;
  assign new_P3_ADD_558_U119 = ~new_P3_ADD_558_U49;
  assign new_P3_ADD_558_U120 = ~new_P3_ADD_558_U51;
  assign new_P3_ADD_558_U121 = ~new_P3_ADD_558_U53;
  assign new_P3_ADD_558_U122 = ~new_P3_ADD_558_U55;
  assign new_P3_ADD_558_U123 = ~new_P3_ADD_558_U57;
  assign new_P3_ADD_558_U124 = ~new_P3_ADD_558_U59;
  assign new_P3_ADD_558_U125 = ~new_P3_ADD_558_U61;
  assign new_P3_ADD_558_U126 = ~new_P3_ADD_558_U63;
  assign new_P3_ADD_558_U127 = ~new_P3_ADD_558_U97;
  assign new_P3_ADD_558_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_558_U22;
  assign new_P3_ADD_558_U129 = ~new_P3_ADD_558_U105 | ~new_P3_ADD_558_U21;
  assign new_P3_ADD_558_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_558_U19;
  assign new_P3_ADD_558_U131 = ~new_P3_ADD_558_U104 | ~new_P3_ADD_558_U20;
  assign new_P3_ADD_558_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_558_U17;
  assign new_P3_ADD_558_U133 = ~new_P3_ADD_558_U103 | ~new_P3_ADD_558_U18;
  assign new_P3_ADD_558_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_558_U15;
  assign new_P3_ADD_558_U135 = ~new_P3_ADD_558_U102 | ~new_P3_ADD_558_U16;
  assign new_P3_ADD_558_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_558_U13;
  assign new_P3_ADD_558_U137 = ~new_P3_ADD_558_U101 | ~new_P3_ADD_558_U14;
  assign new_P3_ADD_558_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_558_U11;
  assign new_P3_ADD_558_U139 = ~new_P3_ADD_558_U100 | ~new_P3_ADD_558_U12;
  assign new_P3_ADD_558_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_558_U9;
  assign new_P3_ADD_558_U141 = ~new_P3_ADD_558_U99 | ~new_P3_ADD_558_U10;
  assign new_P3_ADD_558_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_558_U97;
  assign new_P3_ADD_558_U143 = ~new_P3_ADD_558_U127 | ~new_P3_ADD_558_U96;
  assign new_P3_ADD_558_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_558_U63;
  assign new_P3_ADD_558_U145 = ~new_P3_ADD_558_U126 | ~new_P3_ADD_558_U64;
  assign new_P3_ADD_558_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_558_U7;
  assign new_P3_ADD_558_U147 = ~new_P3_ADD_558_U98 | ~new_P3_ADD_558_U8;
  assign new_P3_ADD_558_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_558_U61;
  assign new_P3_ADD_558_U149 = ~new_P3_ADD_558_U125 | ~new_P3_ADD_558_U62;
  assign new_P3_ADD_558_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_558_U59;
  assign new_P3_ADD_558_U151 = ~new_P3_ADD_558_U124 | ~new_P3_ADD_558_U60;
  assign new_P3_ADD_558_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_558_U57;
  assign new_P3_ADD_558_U153 = ~new_P3_ADD_558_U123 | ~new_P3_ADD_558_U58;
  assign new_P3_ADD_558_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_558_U55;
  assign new_P3_ADD_558_U155 = ~new_P3_ADD_558_U122 | ~new_P3_ADD_558_U56;
  assign new_P3_ADD_558_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_558_U53;
  assign new_P3_ADD_558_U157 = ~new_P3_ADD_558_U121 | ~new_P3_ADD_558_U54;
  assign new_P3_ADD_558_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_558_U51;
  assign new_P3_ADD_558_U159 = ~new_P3_ADD_558_U120 | ~new_P3_ADD_558_U52;
  assign new_P3_ADD_558_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_558_U49;
  assign new_P3_ADD_558_U161 = ~new_P3_ADD_558_U119 | ~new_P3_ADD_558_U50;
  assign new_P3_ADD_558_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_558_U47;
  assign new_P3_ADD_558_U163 = ~new_P3_ADD_558_U118 | ~new_P3_ADD_558_U48;
  assign new_P3_ADD_558_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_558_U45;
  assign new_P3_ADD_558_U165 = ~new_P3_ADD_558_U117 | ~new_P3_ADD_558_U46;
  assign new_P3_ADD_558_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_558_U43;
  assign new_P3_ADD_558_U167 = ~new_P3_ADD_558_U116 | ~new_P3_ADD_558_U44;
  assign new_P3_ADD_558_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_558_U5;
  assign new_P3_ADD_558_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_558_U6;
  assign new_P3_ADD_558_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_558_U41;
  assign new_P3_ADD_558_U171 = ~new_P3_ADD_558_U115 | ~new_P3_ADD_558_U42;
  assign new_P3_ADD_558_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_558_U39;
  assign new_P3_ADD_558_U173 = ~new_P3_ADD_558_U114 | ~new_P3_ADD_558_U40;
  assign new_P3_ADD_558_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_558_U37;
  assign new_P3_ADD_558_U175 = ~new_P3_ADD_558_U113 | ~new_P3_ADD_558_U38;
  assign new_P3_ADD_558_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_558_U35;
  assign new_P3_ADD_558_U177 = ~new_P3_ADD_558_U112 | ~new_P3_ADD_558_U36;
  assign new_P3_ADD_558_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_558_U33;
  assign new_P3_ADD_558_U179 = ~new_P3_ADD_558_U111 | ~new_P3_ADD_558_U34;
  assign new_P3_ADD_558_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_558_U31;
  assign new_P3_ADD_558_U181 = ~new_P3_ADD_558_U110 | ~new_P3_ADD_558_U32;
  assign new_P3_ADD_558_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_558_U29;
  assign new_P3_ADD_558_U183 = ~new_P3_ADD_558_U109 | ~new_P3_ADD_558_U30;
  assign new_P3_ADD_558_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_558_U27;
  assign new_P3_ADD_558_U185 = ~new_P3_ADD_558_U108 | ~new_P3_ADD_558_U28;
  assign new_P3_ADD_558_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_558_U25;
  assign new_P3_ADD_558_U187 = ~new_P3_ADD_558_U107 | ~new_P3_ADD_558_U26;
  assign new_P3_ADD_558_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_558_U23;
  assign new_P3_ADD_558_U189 = ~new_P3_ADD_558_U106 | ~new_P3_ADD_558_U24;
  assign new_P3_ADD_385_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_385_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_385_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_385_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_385_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_385_U98;
  assign new_P3_ADD_385_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_385_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_385_U99;
  assign new_P3_ADD_385_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_385_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_385_U100;
  assign new_P3_ADD_385_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_385_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_385_U101;
  assign new_P3_ADD_385_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_385_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_385_U102;
  assign new_P3_ADD_385_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_385_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_385_U103;
  assign new_P3_ADD_385_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_385_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_385_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_385_U104;
  assign new_P3_ADD_385_U23 = ~new_P3_ADD_385_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_385_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_385_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_385_U106;
  assign new_P3_ADD_385_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_385_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_385_U107;
  assign new_P3_ADD_385_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_385_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_385_U108;
  assign new_P3_ADD_385_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_385_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_385_U109;
  assign new_P3_ADD_385_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_385_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_385_U110;
  assign new_P3_ADD_385_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_385_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_385_U111;
  assign new_P3_ADD_385_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_385_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_385_U112;
  assign new_P3_ADD_385_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_385_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_385_U113;
  assign new_P3_ADD_385_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_385_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_385_U114;
  assign new_P3_ADD_385_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_385_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_385_U115;
  assign new_P3_ADD_385_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_385_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_385_U116;
  assign new_P3_ADD_385_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_385_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_385_U117;
  assign new_P3_ADD_385_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_385_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_385_U118;
  assign new_P3_ADD_385_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_385_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_385_U119;
  assign new_P3_ADD_385_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_385_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_385_U120;
  assign new_P3_ADD_385_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_385_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_385_U121;
  assign new_P3_ADD_385_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_385_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_385_U122;
  assign new_P3_ADD_385_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_385_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_385_U123;
  assign new_P3_ADD_385_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_385_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_385_U124;
  assign new_P3_ADD_385_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_385_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_385_U125;
  assign new_P3_ADD_385_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_385_U65 = ~new_P3_ADD_385_U129 | ~new_P3_ADD_385_U128;
  assign new_P3_ADD_385_U66 = ~new_P3_ADD_385_U131 | ~new_P3_ADD_385_U130;
  assign new_P3_ADD_385_U67 = ~new_P3_ADD_385_U133 | ~new_P3_ADD_385_U132;
  assign new_P3_ADD_385_U68 = ~new_P3_ADD_385_U135 | ~new_P3_ADD_385_U134;
  assign new_P3_ADD_385_U69 = ~new_P3_ADD_385_U137 | ~new_P3_ADD_385_U136;
  assign new_P3_ADD_385_U70 = ~new_P3_ADD_385_U139 | ~new_P3_ADD_385_U138;
  assign new_P3_ADD_385_U71 = ~new_P3_ADD_385_U141 | ~new_P3_ADD_385_U140;
  assign new_P3_ADD_385_U72 = ~new_P3_ADD_385_U143 | ~new_P3_ADD_385_U142;
  assign new_P3_ADD_385_U73 = ~new_P3_ADD_385_U145 | ~new_P3_ADD_385_U144;
  assign new_P3_ADD_385_U74 = ~new_P3_ADD_385_U147 | ~new_P3_ADD_385_U146;
  assign new_P3_ADD_385_U75 = ~new_P3_ADD_385_U149 | ~new_P3_ADD_385_U148;
  assign new_P3_ADD_385_U76 = ~new_P3_ADD_385_U151 | ~new_P3_ADD_385_U150;
  assign new_P3_ADD_385_U77 = ~new_P3_ADD_385_U153 | ~new_P3_ADD_385_U152;
  assign new_P3_ADD_385_U78 = ~new_P3_ADD_385_U155 | ~new_P3_ADD_385_U154;
  assign new_P3_ADD_385_U79 = ~new_P3_ADD_385_U157 | ~new_P3_ADD_385_U156;
  assign new_P3_ADD_385_U80 = ~new_P3_ADD_385_U159 | ~new_P3_ADD_385_U158;
  assign new_P3_ADD_385_U81 = ~new_P3_ADD_385_U161 | ~new_P3_ADD_385_U160;
  assign new_P3_ADD_385_U82 = ~new_P3_ADD_385_U163 | ~new_P3_ADD_385_U162;
  assign new_P3_ADD_385_U83 = ~new_P3_ADD_385_U165 | ~new_P3_ADD_385_U164;
  assign new_P3_ADD_385_U84 = ~new_P3_ADD_385_U167 | ~new_P3_ADD_385_U166;
  assign new_P3_ADD_385_U85 = ~new_P3_ADD_385_U169 | ~new_P3_ADD_385_U168;
  assign new_P3_ADD_385_U86 = ~new_P3_ADD_385_U171 | ~new_P3_ADD_385_U170;
  assign new_P3_ADD_385_U87 = ~new_P3_ADD_385_U173 | ~new_P3_ADD_385_U172;
  assign new_P3_ADD_385_U88 = ~new_P3_ADD_385_U175 | ~new_P3_ADD_385_U174;
  assign new_P3_ADD_385_U89 = ~new_P3_ADD_385_U177 | ~new_P3_ADD_385_U176;
  assign new_P3_ADD_385_U90 = ~new_P3_ADD_385_U179 | ~new_P3_ADD_385_U178;
  assign new_P3_ADD_385_U91 = ~new_P3_ADD_385_U181 | ~new_P3_ADD_385_U180;
  assign new_P3_ADD_385_U92 = ~new_P3_ADD_385_U183 | ~new_P3_ADD_385_U182;
  assign new_P3_ADD_385_U93 = ~new_P3_ADD_385_U185 | ~new_P3_ADD_385_U184;
  assign new_P3_ADD_385_U94 = ~new_P3_ADD_385_U187 | ~new_P3_ADD_385_U186;
  assign new_P3_ADD_385_U95 = ~new_P3_ADD_385_U189 | ~new_P3_ADD_385_U188;
  assign new_P3_ADD_385_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_385_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_385_U126;
  assign new_P3_ADD_385_U98 = ~new_P3_ADD_385_U7;
  assign new_P3_ADD_385_U99 = ~new_P3_ADD_385_U9;
  assign new_P3_ADD_385_U100 = ~new_P3_ADD_385_U11;
  assign new_P3_ADD_385_U101 = ~new_P3_ADD_385_U13;
  assign new_P3_ADD_385_U102 = ~new_P3_ADD_385_U15;
  assign new_P3_ADD_385_U103 = ~new_P3_ADD_385_U17;
  assign new_P3_ADD_385_U104 = ~new_P3_ADD_385_U19;
  assign new_P3_ADD_385_U105 = ~new_P3_ADD_385_U22;
  assign new_P3_ADD_385_U106 = ~new_P3_ADD_385_U23;
  assign new_P3_ADD_385_U107 = ~new_P3_ADD_385_U25;
  assign new_P3_ADD_385_U108 = ~new_P3_ADD_385_U27;
  assign new_P3_ADD_385_U109 = ~new_P3_ADD_385_U29;
  assign new_P3_ADD_385_U110 = ~new_P3_ADD_385_U31;
  assign new_P3_ADD_385_U111 = ~new_P3_ADD_385_U33;
  assign new_P3_ADD_385_U112 = ~new_P3_ADD_385_U35;
  assign new_P3_ADD_385_U113 = ~new_P3_ADD_385_U37;
  assign new_P3_ADD_385_U114 = ~new_P3_ADD_385_U39;
  assign new_P3_ADD_385_U115 = ~new_P3_ADD_385_U41;
  assign new_P3_ADD_385_U116 = ~new_P3_ADD_385_U43;
  assign new_P3_ADD_385_U117 = ~new_P3_ADD_385_U45;
  assign new_P3_ADD_385_U118 = ~new_P3_ADD_385_U47;
  assign new_P3_ADD_385_U119 = ~new_P3_ADD_385_U49;
  assign new_P3_ADD_385_U120 = ~new_P3_ADD_385_U51;
  assign new_P3_ADD_385_U121 = ~new_P3_ADD_385_U53;
  assign new_P3_ADD_385_U122 = ~new_P3_ADD_385_U55;
  assign new_P3_ADD_385_U123 = ~new_P3_ADD_385_U57;
  assign new_P3_ADD_385_U124 = ~new_P3_ADD_385_U59;
  assign new_P3_ADD_385_U125 = ~new_P3_ADD_385_U61;
  assign new_P3_ADD_385_U126 = ~new_P3_ADD_385_U63;
  assign new_P3_ADD_385_U127 = ~new_P3_ADD_385_U97;
  assign new_P3_ADD_385_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_385_U22;
  assign new_P3_ADD_385_U129 = ~new_P3_ADD_385_U105 | ~new_P3_ADD_385_U21;
  assign new_P3_ADD_385_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_385_U19;
  assign new_P3_ADD_385_U131 = ~new_P3_ADD_385_U104 | ~new_P3_ADD_385_U20;
  assign new_P3_ADD_385_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_385_U17;
  assign new_P3_ADD_385_U133 = ~new_P3_ADD_385_U103 | ~new_P3_ADD_385_U18;
  assign new_P3_ADD_385_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_385_U15;
  assign new_P3_ADD_385_U135 = ~new_P3_ADD_385_U102 | ~new_P3_ADD_385_U16;
  assign new_P3_ADD_385_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_385_U13;
  assign new_P3_ADD_385_U137 = ~new_P3_ADD_385_U101 | ~new_P3_ADD_385_U14;
  assign new_P3_ADD_385_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_385_U11;
  assign new_P3_ADD_385_U139 = ~new_P3_ADD_385_U100 | ~new_P3_ADD_385_U12;
  assign new_P3_ADD_385_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_385_U9;
  assign new_P3_ADD_385_U141 = ~new_P3_ADD_385_U99 | ~new_P3_ADD_385_U10;
  assign new_P3_ADD_385_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_385_U97;
  assign new_P3_ADD_385_U143 = ~new_P3_ADD_385_U127 | ~new_P3_ADD_385_U96;
  assign new_P3_ADD_385_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_385_U63;
  assign new_P3_ADD_385_U145 = ~new_P3_ADD_385_U126 | ~new_P3_ADD_385_U64;
  assign new_P3_ADD_385_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_385_U7;
  assign new_P3_ADD_385_U147 = ~new_P3_ADD_385_U98 | ~new_P3_ADD_385_U8;
  assign new_P3_ADD_385_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_385_U61;
  assign new_P3_ADD_385_U149 = ~new_P3_ADD_385_U125 | ~new_P3_ADD_385_U62;
  assign new_P3_ADD_385_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_385_U59;
  assign new_P3_ADD_385_U151 = ~new_P3_ADD_385_U124 | ~new_P3_ADD_385_U60;
  assign new_P3_ADD_385_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_385_U57;
  assign new_P3_ADD_385_U153 = ~new_P3_ADD_385_U123 | ~new_P3_ADD_385_U58;
  assign new_P3_ADD_385_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_385_U55;
  assign new_P3_ADD_385_U155 = ~new_P3_ADD_385_U122 | ~new_P3_ADD_385_U56;
  assign new_P3_ADD_385_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_385_U53;
  assign new_P3_ADD_385_U157 = ~new_P3_ADD_385_U121 | ~new_P3_ADD_385_U54;
  assign new_P3_ADD_385_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_385_U51;
  assign new_P3_ADD_385_U159 = ~new_P3_ADD_385_U120 | ~new_P3_ADD_385_U52;
  assign new_P3_ADD_385_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_385_U49;
  assign new_P3_ADD_385_U161 = ~new_P3_ADD_385_U119 | ~new_P3_ADD_385_U50;
  assign new_P3_ADD_385_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_385_U47;
  assign new_P3_ADD_385_U163 = ~new_P3_ADD_385_U118 | ~new_P3_ADD_385_U48;
  assign new_P3_ADD_385_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_385_U45;
  assign new_P3_ADD_385_U165 = ~new_P3_ADD_385_U117 | ~new_P3_ADD_385_U46;
  assign new_P3_ADD_385_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_385_U43;
  assign new_P3_ADD_385_U167 = ~new_P3_ADD_385_U116 | ~new_P3_ADD_385_U44;
  assign new_P3_ADD_385_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_385_U5;
  assign new_P3_ADD_385_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_385_U6;
  assign new_P3_ADD_385_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_385_U41;
  assign new_P3_ADD_385_U171 = ~new_P3_ADD_385_U115 | ~new_P3_ADD_385_U42;
  assign new_P3_ADD_385_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_385_U39;
  assign new_P3_ADD_385_U173 = ~new_P3_ADD_385_U114 | ~new_P3_ADD_385_U40;
  assign new_P3_ADD_385_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_385_U37;
  assign new_P3_ADD_385_U175 = ~new_P3_ADD_385_U113 | ~new_P3_ADD_385_U38;
  assign new_P3_ADD_385_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_385_U35;
  assign new_P3_ADD_385_U177 = ~new_P3_ADD_385_U112 | ~new_P3_ADD_385_U36;
  assign new_P3_ADD_385_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_385_U33;
  assign new_P3_ADD_385_U179 = ~new_P3_ADD_385_U111 | ~new_P3_ADD_385_U34;
  assign new_P3_ADD_385_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_385_U31;
  assign new_P3_ADD_385_U181 = ~new_P3_ADD_385_U110 | ~new_P3_ADD_385_U32;
  assign new_P3_ADD_385_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_385_U29;
  assign new_P3_ADD_385_U183 = ~new_P3_ADD_385_U109 | ~new_P3_ADD_385_U30;
  assign new_P3_ADD_385_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_385_U27;
  assign new_P3_ADD_385_U185 = ~new_P3_ADD_385_U108 | ~new_P3_ADD_385_U28;
  assign new_P3_ADD_385_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_385_U25;
  assign new_P3_ADD_385_U187 = ~new_P3_ADD_385_U107 | ~new_P3_ADD_385_U26;
  assign new_P3_ADD_385_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_385_U23;
  assign new_P3_ADD_385_U189 = ~new_P3_ADD_385_U106 | ~new_P3_ADD_385_U24;
  assign new_P3_ADD_357_U6 = ~new_P3_ADD_357_U15 | ~new_P3_ADD_357_U23;
  assign new_P3_ADD_357_U7 = new_P3_ADD_357_U29 & new_P3_ADD_357_U11;
  assign new_P3_ADD_357_U8 = new_P3_ADD_357_U27 & new_P3_ADD_357_U12;
  assign new_P3_ADD_357_U9 = new_P3_ADD_357_U25 & new_P3_ADD_357_U6;
  assign new_P3_ADD_357_U10 = ~new_P3_SUB_357_U10;
  assign new_P3_ADD_357_U11 = new_P3_SUB_357_U11 | new_P3_SUB_357_U7 | new_P3_SUB_357_U12;
  assign new_P3_ADD_357_U12 = ~new_P3_ADD_357_U14 | ~new_P3_ADD_357_U22;
  assign new_P3_ADD_357_U13 = ~new_P3_ADD_357_U35 | ~new_P3_ADD_357_U34;
  assign new_P3_ADD_357_U14 = ~new_P3_SUB_357_U13 & ~new_P3_SUB_357_U9;
  assign new_P3_ADD_357_U15 = ~new_P3_SUB_357_U6 & ~new_P3_SUB_357_U8;
  assign new_P3_ADD_357_U16 = ~new_P3_SUB_357_U6;
  assign new_P3_ADD_357_U17 = new_P3_ADD_357_U31 & new_P3_ADD_357_U30;
  assign new_P3_ADD_357_U18 = ~new_P3_SUB_357_U13;
  assign new_P3_ADD_357_U19 = new_P3_ADD_357_U33 & new_P3_ADD_357_U32;
  assign new_P3_ADD_357_U20 = ~new_P3_SUB_357_U7;
  assign new_P3_ADD_357_U21 = ~new_P3_SUB_357_U12;
  assign new_P3_ADD_357_U22 = ~new_P3_ADD_357_U11;
  assign new_P3_ADD_357_U23 = ~new_P3_ADD_357_U12;
  assign new_P3_ADD_357_U24 = ~new_P3_ADD_357_U23 | ~new_P3_ADD_357_U16;
  assign new_P3_ADD_357_U25 = ~new_P3_SUB_357_U8 | ~new_P3_ADD_357_U24;
  assign new_P3_ADD_357_U26 = ~new_P3_ADD_357_U22 | ~new_P3_ADD_357_U18;
  assign new_P3_ADD_357_U27 = ~new_P3_SUB_357_U9 | ~new_P3_ADD_357_U26;
  assign new_P3_ADD_357_U28 = new_P3_SUB_357_U7 | new_P3_SUB_357_U12;
  assign new_P3_ADD_357_U29 = ~new_P3_SUB_357_U11 | ~new_P3_ADD_357_U28;
  assign new_P3_ADD_357_U30 = ~new_P3_SUB_357_U6 | ~new_P3_ADD_357_U12;
  assign new_P3_ADD_357_U31 = ~new_P3_ADD_357_U23 | ~new_P3_ADD_357_U16;
  assign new_P3_ADD_357_U32 = ~new_P3_SUB_357_U13 | ~new_P3_ADD_357_U11;
  assign new_P3_ADD_357_U33 = ~new_P3_ADD_357_U22 | ~new_P3_ADD_357_U18;
  assign new_P3_ADD_357_U34 = ~new_P3_SUB_357_U7 | ~new_P3_ADD_357_U21;
  assign new_P3_ADD_357_U35 = ~new_P3_SUB_357_U12 | ~new_P3_ADD_357_U20;
  assign new_P3_ADD_547_U5 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_547_U6 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_547_U7 = ~P3_INSTADDRPOINTER_REG_1_ | ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_547_U8 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_547_U9 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_547_U98;
  assign new_P3_ADD_547_U10 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_547_U11 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_547_U99;
  assign new_P3_ADD_547_U12 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_547_U13 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_547_U100;
  assign new_P3_ADD_547_U14 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_547_U15 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_547_U101;
  assign new_P3_ADD_547_U16 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_547_U17 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_547_U102;
  assign new_P3_ADD_547_U18 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_547_U19 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_547_U103;
  assign new_P3_ADD_547_U20 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_547_U21 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_547_U22 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_547_U104;
  assign new_P3_ADD_547_U23 = ~new_P3_ADD_547_U105 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_547_U24 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_547_U25 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_547_U106;
  assign new_P3_ADD_547_U26 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_547_U27 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_547_U107;
  assign new_P3_ADD_547_U28 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_547_U29 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_547_U108;
  assign new_P3_ADD_547_U30 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_547_U31 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_547_U109;
  assign new_P3_ADD_547_U32 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_547_U33 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_547_U110;
  assign new_P3_ADD_547_U34 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_547_U35 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_547_U111;
  assign new_P3_ADD_547_U36 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_547_U37 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_547_U112;
  assign new_P3_ADD_547_U38 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_547_U39 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_547_U113;
  assign new_P3_ADD_547_U40 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_547_U41 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_547_U114;
  assign new_P3_ADD_547_U42 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_547_U43 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_547_U115;
  assign new_P3_ADD_547_U44 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_547_U45 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_547_U116;
  assign new_P3_ADD_547_U46 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_547_U47 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_547_U117;
  assign new_P3_ADD_547_U48 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_547_U49 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_547_U118;
  assign new_P3_ADD_547_U50 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_547_U51 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_547_U119;
  assign new_P3_ADD_547_U52 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_547_U53 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_547_U120;
  assign new_P3_ADD_547_U54 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_547_U55 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_547_U121;
  assign new_P3_ADD_547_U56 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_547_U57 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_547_U122;
  assign new_P3_ADD_547_U58 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_547_U59 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_547_U123;
  assign new_P3_ADD_547_U60 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_547_U61 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_547_U124;
  assign new_P3_ADD_547_U62 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_547_U63 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_547_U125;
  assign new_P3_ADD_547_U64 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_547_U65 = ~new_P3_ADD_547_U129 | ~new_P3_ADD_547_U128;
  assign new_P3_ADD_547_U66 = ~new_P3_ADD_547_U131 | ~new_P3_ADD_547_U130;
  assign new_P3_ADD_547_U67 = ~new_P3_ADD_547_U133 | ~new_P3_ADD_547_U132;
  assign new_P3_ADD_547_U68 = ~new_P3_ADD_547_U135 | ~new_P3_ADD_547_U134;
  assign new_P3_ADD_547_U69 = ~new_P3_ADD_547_U137 | ~new_P3_ADD_547_U136;
  assign new_P3_ADD_547_U70 = ~new_P3_ADD_547_U139 | ~new_P3_ADD_547_U138;
  assign new_P3_ADD_547_U71 = ~new_P3_ADD_547_U141 | ~new_P3_ADD_547_U140;
  assign new_P3_ADD_547_U72 = ~new_P3_ADD_547_U143 | ~new_P3_ADD_547_U142;
  assign new_P3_ADD_547_U73 = ~new_P3_ADD_547_U145 | ~new_P3_ADD_547_U144;
  assign new_P3_ADD_547_U74 = ~new_P3_ADD_547_U147 | ~new_P3_ADD_547_U146;
  assign new_P3_ADD_547_U75 = ~new_P3_ADD_547_U149 | ~new_P3_ADD_547_U148;
  assign new_P3_ADD_547_U76 = ~new_P3_ADD_547_U151 | ~new_P3_ADD_547_U150;
  assign new_P3_ADD_547_U77 = ~new_P3_ADD_547_U153 | ~new_P3_ADD_547_U152;
  assign new_P3_ADD_547_U78 = ~new_P3_ADD_547_U155 | ~new_P3_ADD_547_U154;
  assign new_P3_ADD_547_U79 = ~new_P3_ADD_547_U157 | ~new_P3_ADD_547_U156;
  assign new_P3_ADD_547_U80 = ~new_P3_ADD_547_U159 | ~new_P3_ADD_547_U158;
  assign new_P3_ADD_547_U81 = ~new_P3_ADD_547_U161 | ~new_P3_ADD_547_U160;
  assign new_P3_ADD_547_U82 = ~new_P3_ADD_547_U163 | ~new_P3_ADD_547_U162;
  assign new_P3_ADD_547_U83 = ~new_P3_ADD_547_U165 | ~new_P3_ADD_547_U164;
  assign new_P3_ADD_547_U84 = ~new_P3_ADD_547_U167 | ~new_P3_ADD_547_U166;
  assign new_P3_ADD_547_U85 = ~new_P3_ADD_547_U169 | ~new_P3_ADD_547_U168;
  assign new_P3_ADD_547_U86 = ~new_P3_ADD_547_U171 | ~new_P3_ADD_547_U170;
  assign new_P3_ADD_547_U87 = ~new_P3_ADD_547_U173 | ~new_P3_ADD_547_U172;
  assign new_P3_ADD_547_U88 = ~new_P3_ADD_547_U175 | ~new_P3_ADD_547_U174;
  assign new_P3_ADD_547_U89 = ~new_P3_ADD_547_U177 | ~new_P3_ADD_547_U176;
  assign new_P3_ADD_547_U90 = ~new_P3_ADD_547_U179 | ~new_P3_ADD_547_U178;
  assign new_P3_ADD_547_U91 = ~new_P3_ADD_547_U181 | ~new_P3_ADD_547_U180;
  assign new_P3_ADD_547_U92 = ~new_P3_ADD_547_U183 | ~new_P3_ADD_547_U182;
  assign new_P3_ADD_547_U93 = ~new_P3_ADD_547_U185 | ~new_P3_ADD_547_U184;
  assign new_P3_ADD_547_U94 = ~new_P3_ADD_547_U187 | ~new_P3_ADD_547_U186;
  assign new_P3_ADD_547_U95 = ~new_P3_ADD_547_U189 | ~new_P3_ADD_547_U188;
  assign new_P3_ADD_547_U96 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_547_U97 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_547_U126;
  assign new_P3_ADD_547_U98 = ~new_P3_ADD_547_U7;
  assign new_P3_ADD_547_U99 = ~new_P3_ADD_547_U9;
  assign new_P3_ADD_547_U100 = ~new_P3_ADD_547_U11;
  assign new_P3_ADD_547_U101 = ~new_P3_ADD_547_U13;
  assign new_P3_ADD_547_U102 = ~new_P3_ADD_547_U15;
  assign new_P3_ADD_547_U103 = ~new_P3_ADD_547_U17;
  assign new_P3_ADD_547_U104 = ~new_P3_ADD_547_U19;
  assign new_P3_ADD_547_U105 = ~new_P3_ADD_547_U22;
  assign new_P3_ADD_547_U106 = ~new_P3_ADD_547_U23;
  assign new_P3_ADD_547_U107 = ~new_P3_ADD_547_U25;
  assign new_P3_ADD_547_U108 = ~new_P3_ADD_547_U27;
  assign new_P3_ADD_547_U109 = ~new_P3_ADD_547_U29;
  assign new_P3_ADD_547_U110 = ~new_P3_ADD_547_U31;
  assign new_P3_ADD_547_U111 = ~new_P3_ADD_547_U33;
  assign new_P3_ADD_547_U112 = ~new_P3_ADD_547_U35;
  assign new_P3_ADD_547_U113 = ~new_P3_ADD_547_U37;
  assign new_P3_ADD_547_U114 = ~new_P3_ADD_547_U39;
  assign new_P3_ADD_547_U115 = ~new_P3_ADD_547_U41;
  assign new_P3_ADD_547_U116 = ~new_P3_ADD_547_U43;
  assign new_P3_ADD_547_U117 = ~new_P3_ADD_547_U45;
  assign new_P3_ADD_547_U118 = ~new_P3_ADD_547_U47;
  assign new_P3_ADD_547_U119 = ~new_P3_ADD_547_U49;
  assign new_P3_ADD_547_U120 = ~new_P3_ADD_547_U51;
  assign new_P3_ADD_547_U121 = ~new_P3_ADD_547_U53;
  assign new_P3_ADD_547_U122 = ~new_P3_ADD_547_U55;
  assign new_P3_ADD_547_U123 = ~new_P3_ADD_547_U57;
  assign new_P3_ADD_547_U124 = ~new_P3_ADD_547_U59;
  assign new_P3_ADD_547_U125 = ~new_P3_ADD_547_U61;
  assign new_P3_ADD_547_U126 = ~new_P3_ADD_547_U63;
  assign new_P3_ADD_547_U127 = ~new_P3_ADD_547_U97;
  assign new_P3_ADD_547_U128 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_547_U22;
  assign new_P3_ADD_547_U129 = ~new_P3_ADD_547_U105 | ~new_P3_ADD_547_U21;
  assign new_P3_ADD_547_U130 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_547_U19;
  assign new_P3_ADD_547_U131 = ~new_P3_ADD_547_U104 | ~new_P3_ADD_547_U20;
  assign new_P3_ADD_547_U132 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_547_U17;
  assign new_P3_ADD_547_U133 = ~new_P3_ADD_547_U103 | ~new_P3_ADD_547_U18;
  assign new_P3_ADD_547_U134 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_547_U15;
  assign new_P3_ADD_547_U135 = ~new_P3_ADD_547_U102 | ~new_P3_ADD_547_U16;
  assign new_P3_ADD_547_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_547_U13;
  assign new_P3_ADD_547_U137 = ~new_P3_ADD_547_U101 | ~new_P3_ADD_547_U14;
  assign new_P3_ADD_547_U138 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_547_U11;
  assign new_P3_ADD_547_U139 = ~new_P3_ADD_547_U100 | ~new_P3_ADD_547_U12;
  assign new_P3_ADD_547_U140 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_547_U9;
  assign new_P3_ADD_547_U141 = ~new_P3_ADD_547_U99 | ~new_P3_ADD_547_U10;
  assign new_P3_ADD_547_U142 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_547_U97;
  assign new_P3_ADD_547_U143 = ~new_P3_ADD_547_U127 | ~new_P3_ADD_547_U96;
  assign new_P3_ADD_547_U144 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_547_U63;
  assign new_P3_ADD_547_U145 = ~new_P3_ADD_547_U126 | ~new_P3_ADD_547_U64;
  assign new_P3_ADD_547_U146 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_547_U7;
  assign new_P3_ADD_547_U147 = ~new_P3_ADD_547_U98 | ~new_P3_ADD_547_U8;
  assign new_P3_ADD_547_U148 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_547_U61;
  assign new_P3_ADD_547_U149 = ~new_P3_ADD_547_U125 | ~new_P3_ADD_547_U62;
  assign new_P3_ADD_547_U150 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_547_U59;
  assign new_P3_ADD_547_U151 = ~new_P3_ADD_547_U124 | ~new_P3_ADD_547_U60;
  assign new_P3_ADD_547_U152 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_547_U57;
  assign new_P3_ADD_547_U153 = ~new_P3_ADD_547_U123 | ~new_P3_ADD_547_U58;
  assign new_P3_ADD_547_U154 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_547_U55;
  assign new_P3_ADD_547_U155 = ~new_P3_ADD_547_U122 | ~new_P3_ADD_547_U56;
  assign new_P3_ADD_547_U156 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_547_U53;
  assign new_P3_ADD_547_U157 = ~new_P3_ADD_547_U121 | ~new_P3_ADD_547_U54;
  assign new_P3_ADD_547_U158 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_547_U51;
  assign new_P3_ADD_547_U159 = ~new_P3_ADD_547_U120 | ~new_P3_ADD_547_U52;
  assign new_P3_ADD_547_U160 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_547_U49;
  assign new_P3_ADD_547_U161 = ~new_P3_ADD_547_U119 | ~new_P3_ADD_547_U50;
  assign new_P3_ADD_547_U162 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_547_U47;
  assign new_P3_ADD_547_U163 = ~new_P3_ADD_547_U118 | ~new_P3_ADD_547_U48;
  assign new_P3_ADD_547_U164 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_547_U45;
  assign new_P3_ADD_547_U165 = ~new_P3_ADD_547_U117 | ~new_P3_ADD_547_U46;
  assign new_P3_ADD_547_U166 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_547_U43;
  assign new_P3_ADD_547_U167 = ~new_P3_ADD_547_U116 | ~new_P3_ADD_547_U44;
  assign new_P3_ADD_547_U168 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_547_U5;
  assign new_P3_ADD_547_U169 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_547_U6;
  assign new_P3_ADD_547_U170 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_547_U41;
  assign new_P3_ADD_547_U171 = ~new_P3_ADD_547_U115 | ~new_P3_ADD_547_U42;
  assign new_P3_ADD_547_U172 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_547_U39;
  assign new_P3_ADD_547_U173 = ~new_P3_ADD_547_U114 | ~new_P3_ADD_547_U40;
  assign new_P3_ADD_547_U174 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_547_U37;
  assign new_P3_ADD_547_U175 = ~new_P3_ADD_547_U113 | ~new_P3_ADD_547_U38;
  assign new_P3_ADD_547_U176 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_547_U35;
  assign new_P3_ADD_547_U177 = ~new_P3_ADD_547_U112 | ~new_P3_ADD_547_U36;
  assign new_P3_ADD_547_U178 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_547_U33;
  assign new_P3_ADD_547_U179 = ~new_P3_ADD_547_U111 | ~new_P3_ADD_547_U34;
  assign new_P3_ADD_547_U180 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_547_U31;
  assign new_P3_ADD_547_U181 = ~new_P3_ADD_547_U110 | ~new_P3_ADD_547_U32;
  assign new_P3_ADD_547_U182 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_547_U29;
  assign new_P3_ADD_547_U183 = ~new_P3_ADD_547_U109 | ~new_P3_ADD_547_U30;
  assign new_P3_ADD_547_U184 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_547_U27;
  assign new_P3_ADD_547_U185 = ~new_P3_ADD_547_U108 | ~new_P3_ADD_547_U28;
  assign new_P3_ADD_547_U186 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_547_U25;
  assign new_P3_ADD_547_U187 = ~new_P3_ADD_547_U107 | ~new_P3_ADD_547_U26;
  assign new_P3_ADD_547_U188 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_547_U23;
  assign new_P3_ADD_547_U189 = ~new_P3_ADD_547_U106 | ~new_P3_ADD_547_U24;
  assign new_P3_SUB_412_U6 = ~new_P3_SUB_412_U43 | ~new_P3_SUB_412_U42;
  assign new_P3_SUB_412_U7 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_412_U27;
  assign new_P3_SUB_412_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_412_U9 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_412_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_412_U11 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_412_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_412_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_412_U14 = ~new_P3_SUB_412_U39 | ~new_P3_SUB_412_U38;
  assign new_P3_SUB_412_U15 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_412_U16 = ~new_P3_SUB_412_U48 | ~new_P3_SUB_412_U47;
  assign new_P3_SUB_412_U17 = ~new_P3_SUB_412_U53 | ~new_P3_SUB_412_U52;
  assign new_P3_SUB_412_U18 = ~new_P3_SUB_412_U58 | ~new_P3_SUB_412_U57;
  assign new_P3_SUB_412_U19 = ~new_P3_SUB_412_U63 | ~new_P3_SUB_412_U62;
  assign new_P3_SUB_412_U20 = ~new_P3_SUB_412_U45 | ~new_P3_SUB_412_U44;
  assign new_P3_SUB_412_U21 = ~new_P3_SUB_412_U50 | ~new_P3_SUB_412_U49;
  assign new_P3_SUB_412_U22 = ~new_P3_SUB_412_U55 | ~new_P3_SUB_412_U54;
  assign new_P3_SUB_412_U23 = ~new_P3_SUB_412_U60 | ~new_P3_SUB_412_U59;
  assign new_P3_SUB_412_U24 = ~new_P3_SUB_412_U35 | ~new_P3_SUB_412_U34;
  assign new_P3_SUB_412_U25 = ~new_P3_SUB_412_U31 | ~new_P3_SUB_412_U30;
  assign new_P3_SUB_412_U26 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_412_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_412_U28 = ~new_P3_SUB_412_U7;
  assign new_P3_SUB_412_U29 = ~new_P3_SUB_412_U28 | ~new_P3_SUB_412_U8;
  assign new_P3_SUB_412_U30 = ~new_P3_SUB_412_U29 | ~new_P3_SUB_412_U26;
  assign new_P3_SUB_412_U31 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_412_U7;
  assign new_P3_SUB_412_U32 = ~new_P3_SUB_412_U25;
  assign new_P3_SUB_412_U33 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_412_U10;
  assign new_P3_SUB_412_U34 = ~new_P3_SUB_412_U33 | ~new_P3_SUB_412_U25;
  assign new_P3_SUB_412_U35 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_412_U9;
  assign new_P3_SUB_412_U36 = ~new_P3_SUB_412_U24;
  assign new_P3_SUB_412_U37 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_412_U12;
  assign new_P3_SUB_412_U38 = ~new_P3_SUB_412_U37 | ~new_P3_SUB_412_U24;
  assign new_P3_SUB_412_U39 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_412_U11;
  assign new_P3_SUB_412_U40 = ~new_P3_SUB_412_U14;
  assign new_P3_SUB_412_U41 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_412_U15;
  assign new_P3_SUB_412_U42 = ~new_P3_SUB_412_U40 | ~new_P3_SUB_412_U41;
  assign new_P3_SUB_412_U43 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_412_U13;
  assign new_P3_SUB_412_U44 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_412_U13;
  assign new_P3_SUB_412_U45 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_412_U15;
  assign new_P3_SUB_412_U46 = ~new_P3_SUB_412_U20;
  assign new_P3_SUB_412_U47 = ~new_P3_SUB_412_U46 | ~new_P3_SUB_412_U40;
  assign new_P3_SUB_412_U48 = ~new_P3_SUB_412_U20 | ~new_P3_SUB_412_U14;
  assign new_P3_SUB_412_U49 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_412_U12;
  assign new_P3_SUB_412_U50 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_412_U11;
  assign new_P3_SUB_412_U51 = ~new_P3_SUB_412_U21;
  assign new_P3_SUB_412_U52 = ~new_P3_SUB_412_U36 | ~new_P3_SUB_412_U51;
  assign new_P3_SUB_412_U53 = ~new_P3_SUB_412_U21 | ~new_P3_SUB_412_U24;
  assign new_P3_SUB_412_U54 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_412_U10;
  assign new_P3_SUB_412_U55 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_412_U9;
  assign new_P3_SUB_412_U56 = ~new_P3_SUB_412_U22;
  assign new_P3_SUB_412_U57 = ~new_P3_SUB_412_U32 | ~new_P3_SUB_412_U56;
  assign new_P3_SUB_412_U58 = ~new_P3_SUB_412_U22 | ~new_P3_SUB_412_U25;
  assign new_P3_SUB_412_U59 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_412_U8;
  assign new_P3_SUB_412_U60 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_412_U26;
  assign new_P3_SUB_412_U61 = ~new_P3_SUB_412_U23;
  assign new_P3_SUB_412_U62 = ~new_P3_SUB_412_U61 | ~new_P3_SUB_412_U28;
  assign new_P3_SUB_412_U63 = ~new_P3_SUB_412_U23 | ~new_P3_SUB_412_U7;
  assign new_P3_ADD_371_1212_U4 = new_P3_ADD_371_1212_U133 & new_P3_ADD_371_1212_U132;
  assign new_P3_ADD_371_1212_U5 = new_P3_ADD_371_1212_U196 & new_P3_ADD_371_1212_U48;
  assign new_P3_ADD_371_1212_U6 = new_P3_ADD_371_1212_U194 & new_P3_ADD_371_1212_U49;
  assign new_P3_ADD_371_1212_U7 = new_P3_ADD_371_1212_U192 & new_P3_ADD_371_1212_U78;
  assign new_P3_ADD_371_1212_U8 = new_P3_ADD_371_1212_U191 & new_P3_ADD_371_1212_U53;
  assign new_P3_ADD_371_1212_U9 = new_P3_ADD_371_1212_U189 & new_P3_ADD_371_1212_U56;
  assign new_P3_ADD_371_1212_U10 = new_P3_ADD_371_1212_U187 & new_P3_ADD_371_1212_U59;
  assign new_P3_ADD_371_1212_U11 = new_P3_ADD_371_1212_U185 & new_P3_ADD_371_1212_U168;
  assign new_P3_ADD_371_1212_U12 = new_P3_ADD_371_1212_U184 & new_P3_ADD_371_1212_U62;
  assign new_P3_ADD_371_1212_U13 = new_P3_ADD_371_1212_U183 & new_P3_ADD_371_1212_U65;
  assign new_P3_ADD_371_1212_U14 = new_P3_ADD_371_1212_U181 & new_P3_ADD_371_1212_U68;
  assign new_P3_ADD_371_1212_U15 = new_P3_ADD_371_1212_U179 & new_P3_ADD_371_1212_U70;
  assign new_P3_ADD_371_1212_U16 = new_P3_ADD_371_1212_U178 & new_P3_ADD_371_1212_U73;
  assign new_P3_ADD_371_1212_U17 = new_P3_ADD_371_1212_U176 & new_P3_ADD_371_1212_U75;
  assign new_P3_ADD_371_1212_U18 = new_P3_ADD_371_1212_U162 & new_P3_ADD_371_1212_U159;
  assign new_P3_ADD_371_1212_U19 = new_P3_ADD_371_1212_U155 & new_P3_ADD_371_1212_U152;
  assign new_P3_ADD_371_1212_U20 = ~new_P3_ADD_371_1212_U203 | ~new_P3_ADD_371_1212_U255 | ~new_P3_ADD_371_1212_U254;
  assign new_P3_ADD_371_1212_U21 = ~new_P3_ADD_371_U20;
  assign new_P3_ADD_371_1212_U22 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_371_1212_U23 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_371_1212_U24 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_371_U20;
  assign new_P3_ADD_371_1212_U25 = ~new_P3_ADD_371_U19;
  assign new_P3_ADD_371_1212_U26 = ~new_P3_ADD_371_U5;
  assign new_P3_ADD_371_1212_U27 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_371_1212_U28 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_371_1212_U29 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_371_U5;
  assign new_P3_ADD_371_1212_U30 = ~new_P3_ADD_371_U25;
  assign new_P3_ADD_371_1212_U31 = ~new_P3_ADD_371_U4;
  assign new_P3_ADD_371_1212_U32 = ~P3_INSTADDRPOINTER_REG_0_;
  assign new_P3_ADD_371_1212_U33 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_371_1212_U34 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_371_U4;
  assign new_P3_ADD_371_1212_U35 = ~new_P3_ADD_371_U21;
  assign new_P3_ADD_371_1212_U36 = ~new_P3_ADD_371_U18;
  assign new_P3_ADD_371_1212_U37 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_371_1212_U38 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_371_1212_U39 = ~new_P3_ADD_371_U17;
  assign new_P3_ADD_371_1212_U40 = ~new_P3_ADD_371_U6;
  assign new_P3_ADD_371_1212_U41 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_371_1212_U42 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_371_1212_U43 = ~new_P3_ADD_371_1212_U94 | ~new_P3_ADD_371_1212_U130;
  assign new_P3_ADD_371_1212_U44 = ~new_P3_ADD_371_1212_U77 | ~new_P3_ADD_371_1212_U123;
  assign new_P3_ADD_371_1212_U45 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_371_1212_U46 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_371_1212_U47 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_371_1212_U48 = ~new_P3_ADD_371_1212_U99 | ~new_P3_ADD_371_1212_U108;
  assign new_P3_ADD_371_1212_U49 = ~new_P3_ADD_371_1212_U100 | ~new_P3_ADD_371_1212_U117;
  assign new_P3_ADD_371_1212_U50 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_371_1212_U51 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_371_1212_U52 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_371_1212_U53 = ~new_P3_ADD_371_1212_U163 | ~new_P3_ADD_371_1212_U101;
  assign new_P3_ADD_371_1212_U54 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_371_1212_U55 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_371_1212_U56 = ~new_P3_ADD_371_1212_U102 | ~new_P3_ADD_371_1212_U165;
  assign new_P3_ADD_371_1212_U57 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_371_1212_U58 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_371_1212_U59 = ~new_P3_ADD_371_1212_U103 | ~new_P3_ADD_371_1212_U166;
  assign new_P3_ADD_371_1212_U60 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_371_1212_U61 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_371_1212_U62 = ~new_P3_ADD_371_1212_U104 | ~new_P3_ADD_371_1212_U167;
  assign new_P3_ADD_371_1212_U63 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_371_1212_U64 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_371_1212_U65 = ~new_P3_ADD_371_1212_U105 | ~new_P3_ADD_371_1212_U169;
  assign new_P3_ADD_371_1212_U66 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_371_1212_U67 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_371_1212_U68 = ~new_P3_ADD_371_1212_U106 | ~new_P3_ADD_371_1212_U170;
  assign new_P3_ADD_371_1212_U69 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_371_1212_U70 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_371_1212_U171;
  assign new_P3_ADD_371_1212_U71 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_371_1212_U72 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_371_1212_U73 = ~new_P3_ADD_371_1212_U107 | ~new_P3_ADD_371_1212_U172;
  assign new_P3_ADD_371_1212_U74 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_371_1212_U75 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_371_1212_U173;
  assign new_P3_ADD_371_1212_U76 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_371_1212_U77 = ~new_P3_ADD_371_U21 | ~new_P3_ADD_371_1212_U121;
  assign new_P3_ADD_371_1212_U78 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_371_1212_U163;
  assign new_P3_ADD_371_1212_U79 = ~new_P3_ADD_371_1212_U239 | ~new_P3_ADD_371_1212_U238;
  assign new_P3_ADD_371_1212_U80 = ~new_P3_ADD_371_1212_U246 | ~new_P3_ADD_371_1212_U245;
  assign new_P3_ADD_371_1212_U81 = ~new_P3_ADD_371_1212_U248 | ~new_P3_ADD_371_1212_U247;
  assign new_P3_ADD_371_1212_U82 = ~new_P3_ADD_371_1212_U250 | ~new_P3_ADD_371_1212_U249;
  assign new_P3_ADD_371_1212_U83 = ~new_P3_ADD_371_1212_U257 | ~new_P3_ADD_371_1212_U256;
  assign new_P3_ADD_371_1212_U84 = ~new_P3_ADD_371_1212_U259 | ~new_P3_ADD_371_1212_U258;
  assign new_P3_ADD_371_1212_U85 = ~new_P3_ADD_371_1212_U261 | ~new_P3_ADD_371_1212_U260;
  assign new_P3_ADD_371_1212_U86 = ~new_P3_ADD_371_1212_U263 | ~new_P3_ADD_371_1212_U262;
  assign new_P3_ADD_371_1212_U87 = ~new_P3_ADD_371_1212_U265 | ~new_P3_ADD_371_1212_U264;
  assign new_P3_ADD_371_1212_U88 = ~new_P3_ADD_371_1212_U212 | ~new_P3_ADD_371_1212_U211;
  assign new_P3_ADD_371_1212_U89 = ~new_P3_ADD_371_1212_U219 | ~new_P3_ADD_371_1212_U218;
  assign new_P3_ADD_371_1212_U90 = ~new_P3_ADD_371_1212_U226 | ~new_P3_ADD_371_1212_U225;
  assign new_P3_ADD_371_1212_U91 = ~new_P3_ADD_371_1212_U233 | ~new_P3_ADD_371_1212_U232;
  assign new_P3_ADD_371_1212_U92 = ~new_P3_ADD_371_1212_U237 | ~new_P3_ADD_371_1212_U236;
  assign new_P3_ADD_371_1212_U93 = ~new_P3_ADD_371_1212_U244 | ~new_P3_ADD_371_1212_U243;
  assign new_P3_ADD_371_1212_U94 = new_P3_ADD_371_1212_U129 & new_P3_ADD_371_1212_U128;
  assign new_P3_ADD_371_1212_U95 = new_P3_ADD_371_1212_U137 & new_P3_ADD_371_1212_U136;
  assign new_P3_ADD_371_1212_U96 = new_P3_ADD_371_1212_U24 & new_P3_ADD_371_1212_U228 & new_P3_ADD_371_1212_U227;
  assign new_P3_ADD_371_1212_U97 = new_P3_ADD_371_1212_U154 & new_P3_ADD_371_1212_U4;
  assign new_P3_ADD_371_1212_U98 = new_P3_ADD_371_1212_U29 & new_P3_ADD_371_1212_U235 & new_P3_ADD_371_1212_U234;
  assign new_P3_ADD_371_1212_U99 = P3_INSTADDRPOINTER_REG_9_ & P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_371_1212_U100 = P3_INSTADDRPOINTER_REG_12_ & P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_371_1212_U101 = P3_INSTADDRPOINTER_REG_13_ & P3_INSTADDRPOINTER_REG_14_ & P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_371_1212_U102 = P3_INSTADDRPOINTER_REG_17_ & P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_371_1212_U103 = P3_INSTADDRPOINTER_REG_18_ & P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_371_1212_U104 = P3_INSTADDRPOINTER_REG_20_ & P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_371_1212_U105 = P3_INSTADDRPOINTER_REG_23_ & P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_371_1212_U106 = P3_INSTADDRPOINTER_REG_25_ & P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_371_1212_U107 = P3_INSTADDRPOINTER_REG_28_ & P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_371_1212_U108 = ~new_P3_ADD_371_1212_U148 | ~new_P3_ADD_371_1212_U147;
  assign new_P3_ADD_371_1212_U109 = new_P3_ADD_371_1212_U205 & new_P3_ADD_371_1212_U204;
  assign new_P3_ADD_371_1212_U110 = new_P3_ADD_371_1212_U207 & new_P3_ADD_371_1212_U206;
  assign new_P3_ADD_371_1212_U111 = ~new_P3_ADD_371_1212_U200 | ~new_P3_ADD_371_1212_U144 | ~new_P3_ADD_371_1212_U118;
  assign new_P3_ADD_371_1212_U112 = new_P3_ADD_371_1212_U214 & new_P3_ADD_371_1212_U213;
  assign new_P3_ADD_371_1212_U113 = ~new_P3_ADD_371_1212_U142 | ~new_P3_ADD_371_1212_U141;
  assign new_P3_ADD_371_1212_U114 = new_P3_ADD_371_1212_U221 & new_P3_ADD_371_1212_U220;
  assign new_P3_ADD_371_1212_U115 = ~new_P3_ADD_371_1212_U95 | ~new_P3_ADD_371_1212_U138;
  assign new_P3_ADD_371_1212_U116 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_371_1212_U117 = ~new_P3_ADD_371_1212_U48;
  assign new_P3_ADD_371_1212_U118 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_371_1212_U113;
  assign new_P3_ADD_371_1212_U119 = ~new_P3_ADD_371_1212_U202 | ~new_P3_ADD_371_1212_U201;
  assign new_P3_ADD_371_1212_U120 = ~new_P3_ADD_371_1212_U77;
  assign new_P3_ADD_371_1212_U121 = ~new_P3_ADD_371_1212_U34;
  assign new_P3_ADD_371_1212_U122 = ~new_P3_ADD_371_1212_U35 | ~new_P3_ADD_371_1212_U34;
  assign new_P3_ADD_371_1212_U123 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_371_1212_U122;
  assign new_P3_ADD_371_1212_U124 = ~new_P3_ADD_371_1212_U44;
  assign new_P3_ADD_371_1212_U125 = P3_INSTADDRPOINTER_REG_2_ | new_P3_ADD_371_U5;
  assign new_P3_ADD_371_1212_U126 = ~new_P3_ADD_371_1212_U29;
  assign new_P3_ADD_371_1212_U127 = ~new_P3_ADD_371_1212_U30 | ~new_P3_ADD_371_1212_U29;
  assign new_P3_ADD_371_1212_U128 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_371_1212_U127;
  assign new_P3_ADD_371_1212_U129 = ~new_P3_ADD_371_U25 | ~new_P3_ADD_371_1212_U126;
  assign new_P3_ADD_371_1212_U130 = ~new_P3_ADD_371_1212_U44 | ~new_P3_ADD_371_1212_U119;
  assign new_P3_ADD_371_1212_U131 = ~new_P3_ADD_371_1212_U43;
  assign new_P3_ADD_371_1212_U132 = P3_INSTADDRPOINTER_REG_5_ | new_P3_ADD_371_U19;
  assign new_P3_ADD_371_1212_U133 = P3_INSTADDRPOINTER_REG_4_ | new_P3_ADD_371_U20;
  assign new_P3_ADD_371_1212_U134 = ~new_P3_ADD_371_1212_U24;
  assign new_P3_ADD_371_1212_U135 = ~new_P3_ADD_371_1212_U25 | ~new_P3_ADD_371_1212_U24;
  assign new_P3_ADD_371_1212_U136 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_371_1212_U135;
  assign new_P3_ADD_371_1212_U137 = ~new_P3_ADD_371_U19 | ~new_P3_ADD_371_1212_U134;
  assign new_P3_ADD_371_1212_U138 = ~new_P3_ADD_371_1212_U4 | ~new_P3_ADD_371_1212_U43;
  assign new_P3_ADD_371_1212_U139 = ~new_P3_ADD_371_1212_U115;
  assign new_P3_ADD_371_1212_U140 = new_P3_ADD_371_U18 | P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_371_1212_U141 = ~new_P3_ADD_371_1212_U140 | ~new_P3_ADD_371_1212_U115;
  assign new_P3_ADD_371_1212_U142 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_371_U18;
  assign new_P3_ADD_371_1212_U143 = ~new_P3_ADD_371_1212_U113;
  assign new_P3_ADD_371_1212_U144 = ~new_P3_ADD_371_U17 | ~new_P3_ADD_371_1212_U113;
  assign new_P3_ADD_371_1212_U145 = ~new_P3_ADD_371_1212_U111;
  assign new_P3_ADD_371_1212_U146 = new_P3_ADD_371_U6 | P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_371_1212_U147 = ~new_P3_ADD_371_1212_U146 | ~new_P3_ADD_371_1212_U111;
  assign new_P3_ADD_371_1212_U148 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_371_U6;
  assign new_P3_ADD_371_1212_U149 = ~new_P3_ADD_371_1212_U108;
  assign new_P3_ADD_371_1212_U150 = new_P3_ADD_371_U20 | P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_371_1212_U151 = ~new_P3_ADD_371_1212_U150 | ~new_P3_ADD_371_1212_U43;
  assign new_P3_ADD_371_1212_U152 = ~new_P3_ADD_371_1212_U96 | ~new_P3_ADD_371_1212_U151;
  assign new_P3_ADD_371_1212_U153 = ~new_P3_ADD_371_1212_U131 | ~new_P3_ADD_371_1212_U24;
  assign new_P3_ADD_371_1212_U154 = ~new_P3_ADD_371_U19 | ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_371_1212_U155 = ~new_P3_ADD_371_1212_U97 | ~new_P3_ADD_371_1212_U153;
  assign new_P3_ADD_371_1212_U156 = P3_INSTADDRPOINTER_REG_4_ | new_P3_ADD_371_U20;
  assign new_P3_ADD_371_1212_U157 = new_P3_ADD_371_U5 | P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_371_1212_U158 = ~new_P3_ADD_371_1212_U157 | ~new_P3_ADD_371_1212_U44;
  assign new_P3_ADD_371_1212_U159 = ~new_P3_ADD_371_1212_U98 | ~new_P3_ADD_371_1212_U158;
  assign new_P3_ADD_371_1212_U160 = ~new_P3_ADD_371_1212_U124 | ~new_P3_ADD_371_1212_U29;
  assign new_P3_ADD_371_1212_U161 = ~new_P3_ADD_371_U25 | ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_371_1212_U162 = ~new_P3_ADD_371_1212_U119 | ~new_P3_ADD_371_1212_U160 | ~new_P3_ADD_371_1212_U161;
  assign new_P3_ADD_371_1212_U163 = ~new_P3_ADD_371_1212_U49;
  assign new_P3_ADD_371_1212_U164 = ~new_P3_ADD_371_1212_U78;
  assign new_P3_ADD_371_1212_U165 = ~new_P3_ADD_371_1212_U53;
  assign new_P3_ADD_371_1212_U166 = ~new_P3_ADD_371_1212_U56;
  assign new_P3_ADD_371_1212_U167 = ~new_P3_ADD_371_1212_U59;
  assign new_P3_ADD_371_1212_U168 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_371_1212_U167;
  assign new_P3_ADD_371_1212_U169 = ~new_P3_ADD_371_1212_U62;
  assign new_P3_ADD_371_1212_U170 = ~new_P3_ADD_371_1212_U65;
  assign new_P3_ADD_371_1212_U171 = ~new_P3_ADD_371_1212_U68;
  assign new_P3_ADD_371_1212_U172 = ~new_P3_ADD_371_1212_U70;
  assign new_P3_ADD_371_1212_U173 = ~new_P3_ADD_371_1212_U73;
  assign new_P3_ADD_371_1212_U174 = ~new_P3_ADD_371_1212_U75;
  assign new_P3_ADD_371_1212_U175 = P3_INSTADDRPOINTER_REG_2_ | new_P3_ADD_371_U5;
  assign new_P3_ADD_371_1212_U176 = ~new_P3_ADD_371_1212_U74 | ~new_P3_ADD_371_1212_U73;
  assign new_P3_ADD_371_1212_U177 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_371_1212_U172;
  assign new_P3_ADD_371_1212_U178 = ~new_P3_ADD_371_1212_U71 | ~new_P3_ADD_371_1212_U177;
  assign new_P3_ADD_371_1212_U179 = ~new_P3_ADD_371_1212_U69 | ~new_P3_ADD_371_1212_U68;
  assign new_P3_ADD_371_1212_U180 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_371_1212_U170;
  assign new_P3_ADD_371_1212_U181 = ~new_P3_ADD_371_1212_U66 | ~new_P3_ADD_371_1212_U180;
  assign new_P3_ADD_371_1212_U182 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_371_1212_U169;
  assign new_P3_ADD_371_1212_U183 = ~new_P3_ADD_371_1212_U63 | ~new_P3_ADD_371_1212_U182;
  assign new_P3_ADD_371_1212_U184 = ~new_P3_ADD_371_1212_U61 | ~new_P3_ADD_371_1212_U168;
  assign new_P3_ADD_371_1212_U185 = ~new_P3_ADD_371_1212_U60 | ~new_P3_ADD_371_1212_U59;
  assign new_P3_ADD_371_1212_U186 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_371_1212_U166;
  assign new_P3_ADD_371_1212_U187 = ~new_P3_ADD_371_1212_U58 | ~new_P3_ADD_371_1212_U186;
  assign new_P3_ADD_371_1212_U188 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_371_1212_U165;
  assign new_P3_ADD_371_1212_U189 = ~new_P3_ADD_371_1212_U54 | ~new_P3_ADD_371_1212_U188;
  assign new_P3_ADD_371_1212_U190 = ~new_P3_ADD_371_1212_U164 | ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_371_1212_U191 = ~new_P3_ADD_371_1212_U51 | ~new_P3_ADD_371_1212_U190;
  assign new_P3_ADD_371_1212_U192 = ~new_P3_ADD_371_1212_U50 | ~new_P3_ADD_371_1212_U49;
  assign new_P3_ADD_371_1212_U193 = ~new_P3_ADD_371_1212_U117 | ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_371_1212_U194 = ~new_P3_ADD_371_1212_U47 | ~new_P3_ADD_371_1212_U193;
  assign new_P3_ADD_371_1212_U195 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_371_1212_U108;
  assign new_P3_ADD_371_1212_U196 = ~new_P3_ADD_371_1212_U45 | ~new_P3_ADD_371_1212_U195;
  assign new_P3_ADD_371_1212_U197 = ~new_P3_ADD_371_1212_U156 | ~new_P3_ADD_371_1212_U24;
  assign new_P3_ADD_371_1212_U198 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_371_1212_U174;
  assign new_P3_ADD_371_1212_U199 = ~new_P3_ADD_371_1212_U175 | ~new_P3_ADD_371_1212_U29;
  assign new_P3_ADD_371_1212_U200 = ~new_P3_ADD_371_U17 | ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_371_1212_U201 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_371_1212_U125;
  assign new_P3_ADD_371_1212_U202 = ~new_P3_ADD_371_U25 | ~new_P3_ADD_371_1212_U125;
  assign new_P3_ADD_371_1212_U203 = ~new_P3_ADD_371_1212_U120 | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_371_1212_U204 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_371_1212_U108;
  assign new_P3_ADD_371_1212_U205 = ~new_P3_ADD_371_1212_U149 | ~new_P3_ADD_371_1212_U42;
  assign new_P3_ADD_371_1212_U206 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_371_1212_U40;
  assign new_P3_ADD_371_1212_U207 = ~new_P3_ADD_371_U6 | ~new_P3_ADD_371_1212_U41;
  assign new_P3_ADD_371_1212_U208 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_371_1212_U40;
  assign new_P3_ADD_371_1212_U209 = ~new_P3_ADD_371_U6 | ~new_P3_ADD_371_1212_U41;
  assign new_P3_ADD_371_1212_U210 = ~new_P3_ADD_371_1212_U209 | ~new_P3_ADD_371_1212_U208;
  assign new_P3_ADD_371_1212_U211 = ~new_P3_ADD_371_1212_U110 | ~new_P3_ADD_371_1212_U111;
  assign new_P3_ADD_371_1212_U212 = ~new_P3_ADD_371_1212_U145 | ~new_P3_ADD_371_1212_U210;
  assign new_P3_ADD_371_1212_U213 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_371_1212_U39;
  assign new_P3_ADD_371_1212_U214 = ~new_P3_ADD_371_U17 | ~new_P3_ADD_371_1212_U38;
  assign new_P3_ADD_371_1212_U215 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_371_1212_U39;
  assign new_P3_ADD_371_1212_U216 = ~new_P3_ADD_371_U17 | ~new_P3_ADD_371_1212_U38;
  assign new_P3_ADD_371_1212_U217 = ~new_P3_ADD_371_1212_U216 | ~new_P3_ADD_371_1212_U215;
  assign new_P3_ADD_371_1212_U218 = ~new_P3_ADD_371_1212_U112 | ~new_P3_ADD_371_1212_U113;
  assign new_P3_ADD_371_1212_U219 = ~new_P3_ADD_371_1212_U143 | ~new_P3_ADD_371_1212_U217;
  assign new_P3_ADD_371_1212_U220 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_371_1212_U36;
  assign new_P3_ADD_371_1212_U221 = ~new_P3_ADD_371_U18 | ~new_P3_ADD_371_1212_U37;
  assign new_P3_ADD_371_1212_U222 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_371_1212_U36;
  assign new_P3_ADD_371_1212_U223 = ~new_P3_ADD_371_U18 | ~new_P3_ADD_371_1212_U37;
  assign new_P3_ADD_371_1212_U224 = ~new_P3_ADD_371_1212_U223 | ~new_P3_ADD_371_1212_U222;
  assign new_P3_ADD_371_1212_U225 = ~new_P3_ADD_371_1212_U114 | ~new_P3_ADD_371_1212_U115;
  assign new_P3_ADD_371_1212_U226 = ~new_P3_ADD_371_1212_U139 | ~new_P3_ADD_371_1212_U224;
  assign new_P3_ADD_371_1212_U227 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_371_1212_U25;
  assign new_P3_ADD_371_1212_U228 = ~new_P3_ADD_371_U19 | ~new_P3_ADD_371_1212_U23;
  assign new_P3_ADD_371_1212_U229 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_371_1212_U21;
  assign new_P3_ADD_371_1212_U230 = ~new_P3_ADD_371_U20 | ~new_P3_ADD_371_1212_U22;
  assign new_P3_ADD_371_1212_U231 = ~new_P3_ADD_371_1212_U230 | ~new_P3_ADD_371_1212_U229;
  assign new_P3_ADD_371_1212_U232 = ~new_P3_ADD_371_1212_U197 | ~new_P3_ADD_371_1212_U43;
  assign new_P3_ADD_371_1212_U233 = ~new_P3_ADD_371_1212_U231 | ~new_P3_ADD_371_1212_U131;
  assign new_P3_ADD_371_1212_U234 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_371_1212_U30;
  assign new_P3_ADD_371_1212_U235 = ~new_P3_ADD_371_U25 | ~new_P3_ADD_371_1212_U28;
  assign new_P3_ADD_371_1212_U236 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_371_1212_U198;
  assign new_P3_ADD_371_1212_U237 = ~new_P3_ADD_371_1212_U116 | ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_371_1212_U174;
  assign new_P3_ADD_371_1212_U238 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_371_1212_U75;
  assign new_P3_ADD_371_1212_U239 = ~new_P3_ADD_371_1212_U174 | ~new_P3_ADD_371_1212_U76;
  assign new_P3_ADD_371_1212_U240 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_371_1212_U26;
  assign new_P3_ADD_371_1212_U241 = ~new_P3_ADD_371_U5 | ~new_P3_ADD_371_1212_U27;
  assign new_P3_ADD_371_1212_U242 = ~new_P3_ADD_371_1212_U241 | ~new_P3_ADD_371_1212_U240;
  assign new_P3_ADD_371_1212_U243 = ~new_P3_ADD_371_1212_U199 | ~new_P3_ADD_371_1212_U44;
  assign new_P3_ADD_371_1212_U244 = ~new_P3_ADD_371_1212_U242 | ~new_P3_ADD_371_1212_U124;
  assign new_P3_ADD_371_1212_U245 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_371_1212_U70;
  assign new_P3_ADD_371_1212_U246 = ~new_P3_ADD_371_1212_U172 | ~new_P3_ADD_371_1212_U72;
  assign new_P3_ADD_371_1212_U247 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_371_1212_U65;
  assign new_P3_ADD_371_1212_U248 = ~new_P3_ADD_371_1212_U170 | ~new_P3_ADD_371_1212_U67;
  assign new_P3_ADD_371_1212_U249 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_371_1212_U62;
  assign new_P3_ADD_371_1212_U250 = ~new_P3_ADD_371_1212_U169 | ~new_P3_ADD_371_1212_U64;
  assign new_P3_ADD_371_1212_U251 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_371_1212_U34;
  assign new_P3_ADD_371_1212_U252 = ~new_P3_ADD_371_1212_U121 | ~new_P3_ADD_371_1212_U33;
  assign new_P3_ADD_371_1212_U253 = ~new_P3_ADD_371_1212_U252 | ~new_P3_ADD_371_1212_U251;
  assign new_P3_ADD_371_1212_U254 = ~new_P3_ADD_371_U21 | ~new_P3_ADD_371_1212_U34 | ~new_P3_ADD_371_1212_U33;
  assign new_P3_ADD_371_1212_U255 = ~new_P3_ADD_371_1212_U253 | ~new_P3_ADD_371_1212_U35;
  assign new_P3_ADD_371_1212_U256 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_371_1212_U56;
  assign new_P3_ADD_371_1212_U257 = ~new_P3_ADD_371_1212_U166 | ~new_P3_ADD_371_1212_U57;
  assign new_P3_ADD_371_1212_U258 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_371_1212_U53;
  assign new_P3_ADD_371_1212_U259 = ~new_P3_ADD_371_1212_U165 | ~new_P3_ADD_371_1212_U55;
  assign new_P3_ADD_371_1212_U260 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_371_1212_U78;
  assign new_P3_ADD_371_1212_U261 = ~new_P3_ADD_371_1212_U164 | ~new_P3_ADD_371_1212_U52;
  assign new_P3_ADD_371_1212_U262 = ~new_P3_ADD_371_1212_U117 | ~new_P3_ADD_371_1212_U46;
  assign new_P3_ADD_371_1212_U263 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_371_1212_U48;
  assign new_P3_ADD_371_1212_U264 = ~P3_INSTADDRPOINTER_REG_0_ | ~new_P3_ADD_371_1212_U31;
  assign new_P3_ADD_371_1212_U265 = ~new_P3_ADD_371_U4 | ~new_P3_ADD_371_1212_U32;
  assign new_P3_SUB_504_U6 = ~new_P3_SUB_504_U43 | ~new_P3_SUB_504_U42;
  assign new_P3_SUB_504_U7 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_504_U27;
  assign new_P3_SUB_504_U8 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_504_U9 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_504_U10 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_504_U11 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_504_U12 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_504_U13 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_504_U14 = ~new_P3_SUB_504_U39 | ~new_P3_SUB_504_U38;
  assign new_P3_SUB_504_U15 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_504_U16 = ~new_P3_SUB_504_U48 | ~new_P3_SUB_504_U47;
  assign new_P3_SUB_504_U17 = ~new_P3_SUB_504_U53 | ~new_P3_SUB_504_U52;
  assign new_P3_SUB_504_U18 = ~new_P3_SUB_504_U58 | ~new_P3_SUB_504_U57;
  assign new_P3_SUB_504_U19 = ~new_P3_SUB_504_U63 | ~new_P3_SUB_504_U62;
  assign new_P3_SUB_504_U20 = ~new_P3_SUB_504_U45 | ~new_P3_SUB_504_U44;
  assign new_P3_SUB_504_U21 = ~new_P3_SUB_504_U50 | ~new_P3_SUB_504_U49;
  assign new_P3_SUB_504_U22 = ~new_P3_SUB_504_U55 | ~new_P3_SUB_504_U54;
  assign new_P3_SUB_504_U23 = ~new_P3_SUB_504_U60 | ~new_P3_SUB_504_U59;
  assign new_P3_SUB_504_U24 = ~new_P3_SUB_504_U35 | ~new_P3_SUB_504_U34;
  assign new_P3_SUB_504_U25 = ~new_P3_SUB_504_U31 | ~new_P3_SUB_504_U30;
  assign new_P3_SUB_504_U26 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_504_U27 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_504_U28 = ~new_P3_SUB_504_U7;
  assign new_P3_SUB_504_U29 = ~new_P3_SUB_504_U28 | ~new_P3_SUB_504_U8;
  assign new_P3_SUB_504_U30 = ~new_P3_SUB_504_U29 | ~new_P3_SUB_504_U26;
  assign new_P3_SUB_504_U31 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_504_U7;
  assign new_P3_SUB_504_U32 = ~new_P3_SUB_504_U25;
  assign new_P3_SUB_504_U33 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_504_U10;
  assign new_P3_SUB_504_U34 = ~new_P3_SUB_504_U33 | ~new_P3_SUB_504_U25;
  assign new_P3_SUB_504_U35 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_504_U9;
  assign new_P3_SUB_504_U36 = ~new_P3_SUB_504_U24;
  assign new_P3_SUB_504_U37 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_504_U12;
  assign new_P3_SUB_504_U38 = ~new_P3_SUB_504_U37 | ~new_P3_SUB_504_U24;
  assign new_P3_SUB_504_U39 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_504_U11;
  assign new_P3_SUB_504_U40 = ~new_P3_SUB_504_U14;
  assign new_P3_SUB_504_U41 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_504_U15;
  assign new_P3_SUB_504_U42 = ~new_P3_SUB_504_U40 | ~new_P3_SUB_504_U41;
  assign new_P3_SUB_504_U43 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_504_U13;
  assign new_P3_SUB_504_U44 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_504_U13;
  assign new_P3_SUB_504_U45 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_504_U15;
  assign new_P3_SUB_504_U46 = ~new_P3_SUB_504_U20;
  assign new_P3_SUB_504_U47 = ~new_P3_SUB_504_U46 | ~new_P3_SUB_504_U40;
  assign new_P3_SUB_504_U48 = ~new_P3_SUB_504_U20 | ~new_P3_SUB_504_U14;
  assign new_P3_SUB_504_U49 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_504_U12;
  assign new_P3_SUB_504_U50 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_504_U11;
  assign new_P3_SUB_504_U51 = ~new_P3_SUB_504_U21;
  assign new_P3_SUB_504_U52 = ~new_P3_SUB_504_U36 | ~new_P3_SUB_504_U51;
  assign new_P3_SUB_504_U53 = ~new_P3_SUB_504_U21 | ~new_P3_SUB_504_U24;
  assign new_P3_SUB_504_U54 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_504_U10;
  assign new_P3_SUB_504_U55 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_504_U9;
  assign new_P3_SUB_504_U56 = ~new_P3_SUB_504_U22;
  assign new_P3_SUB_504_U57 = ~new_P3_SUB_504_U32 | ~new_P3_SUB_504_U56;
  assign new_P3_SUB_504_U58 = ~new_P3_SUB_504_U22 | ~new_P3_SUB_504_U25;
  assign new_P3_SUB_504_U59 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_504_U8;
  assign new_P3_SUB_504_U60 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_504_U26;
  assign new_P3_SUB_504_U61 = ~new_P3_SUB_504_U23;
  assign new_P3_SUB_504_U62 = ~new_P3_SUB_504_U61 | ~new_P3_SUB_504_U28;
  assign new_P3_SUB_504_U63 = ~new_P3_SUB_504_U23 | ~new_P3_SUB_504_U7;
  assign new_P3_SUB_401_U6 = ~new_P3_SUB_401_U45 | ~new_P3_SUB_401_U44;
  assign new_P3_SUB_401_U7 = ~new_P3_SUB_401_U9 | ~new_P3_SUB_401_U46;
  assign new_P3_SUB_401_U8 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_SUB_401_U9 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_401_U18;
  assign new_P3_SUB_401_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_401_U11 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_401_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_401_U13 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_401_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_401_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_401_U16 = ~new_P3_SUB_401_U41 | ~new_P3_SUB_401_U40;
  assign new_P3_SUB_401_U17 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_401_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_401_U19 = ~new_P3_SUB_401_U51 | ~new_P3_SUB_401_U50;
  assign new_P3_SUB_401_U20 = ~new_P3_SUB_401_U56 | ~new_P3_SUB_401_U55;
  assign new_P3_SUB_401_U21 = ~new_P3_SUB_401_U61 | ~new_P3_SUB_401_U60;
  assign new_P3_SUB_401_U22 = ~new_P3_SUB_401_U66 | ~new_P3_SUB_401_U65;
  assign new_P3_SUB_401_U23 = ~new_P3_SUB_401_U48 | ~new_P3_SUB_401_U47;
  assign new_P3_SUB_401_U24 = ~new_P3_SUB_401_U53 | ~new_P3_SUB_401_U52;
  assign new_P3_SUB_401_U25 = ~new_P3_SUB_401_U58 | ~new_P3_SUB_401_U57;
  assign new_P3_SUB_401_U26 = ~new_P3_SUB_401_U63 | ~new_P3_SUB_401_U62;
  assign new_P3_SUB_401_U27 = ~new_P3_SUB_401_U37 | ~new_P3_SUB_401_U36;
  assign new_P3_SUB_401_U28 = ~new_P3_SUB_401_U33 | ~new_P3_SUB_401_U32;
  assign new_P3_SUB_401_U29 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_401_U30 = ~new_P3_SUB_401_U9;
  assign new_P3_SUB_401_U31 = ~new_P3_SUB_401_U30 | ~new_P3_SUB_401_U10;
  assign new_P3_SUB_401_U32 = ~new_P3_SUB_401_U31 | ~new_P3_SUB_401_U29;
  assign new_P3_SUB_401_U33 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_401_U9;
  assign new_P3_SUB_401_U34 = ~new_P3_SUB_401_U28;
  assign new_P3_SUB_401_U35 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_401_U12;
  assign new_P3_SUB_401_U36 = ~new_P3_SUB_401_U35 | ~new_P3_SUB_401_U28;
  assign new_P3_SUB_401_U37 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_401_U11;
  assign new_P3_SUB_401_U38 = ~new_P3_SUB_401_U27;
  assign new_P3_SUB_401_U39 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_401_U14;
  assign new_P3_SUB_401_U40 = ~new_P3_SUB_401_U39 | ~new_P3_SUB_401_U27;
  assign new_P3_SUB_401_U41 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_401_U13;
  assign new_P3_SUB_401_U42 = ~new_P3_SUB_401_U16;
  assign new_P3_SUB_401_U43 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_401_U17;
  assign new_P3_SUB_401_U44 = ~new_P3_SUB_401_U42 | ~new_P3_SUB_401_U43;
  assign new_P3_SUB_401_U45 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_401_U15;
  assign new_P3_SUB_401_U46 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_SUB_401_U8;
  assign new_P3_SUB_401_U47 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_401_U15;
  assign new_P3_SUB_401_U48 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_401_U17;
  assign new_P3_SUB_401_U49 = ~new_P3_SUB_401_U23;
  assign new_P3_SUB_401_U50 = ~new_P3_SUB_401_U49 | ~new_P3_SUB_401_U42;
  assign new_P3_SUB_401_U51 = ~new_P3_SUB_401_U23 | ~new_P3_SUB_401_U16;
  assign new_P3_SUB_401_U52 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_401_U14;
  assign new_P3_SUB_401_U53 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_401_U13;
  assign new_P3_SUB_401_U54 = ~new_P3_SUB_401_U24;
  assign new_P3_SUB_401_U55 = ~new_P3_SUB_401_U38 | ~new_P3_SUB_401_U54;
  assign new_P3_SUB_401_U56 = ~new_P3_SUB_401_U24 | ~new_P3_SUB_401_U27;
  assign new_P3_SUB_401_U57 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_401_U12;
  assign new_P3_SUB_401_U58 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_401_U11;
  assign new_P3_SUB_401_U59 = ~new_P3_SUB_401_U25;
  assign new_P3_SUB_401_U60 = ~new_P3_SUB_401_U34 | ~new_P3_SUB_401_U59;
  assign new_P3_SUB_401_U61 = ~new_P3_SUB_401_U25 | ~new_P3_SUB_401_U28;
  assign new_P3_SUB_401_U62 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_401_U10;
  assign new_P3_SUB_401_U63 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_401_U29;
  assign new_P3_SUB_401_U64 = ~new_P3_SUB_401_U26;
  assign new_P3_SUB_401_U65 = ~new_P3_SUB_401_U64 | ~new_P3_SUB_401_U30;
  assign new_P3_SUB_401_U66 = ~new_P3_SUB_401_U26 | ~new_P3_SUB_401_U9;
  assign new_P3_ADD_371_U4 = ~new_P3_U2621;
  assign new_P3_ADD_371_U5 = ~new_P3_ADD_371_U24 | ~new_P3_ADD_371_U32;
  assign new_P3_ADD_371_U6 = new_P3_ADD_371_U22 & new_P3_ADD_371_U30;
  assign new_P3_ADD_371_U7 = ~new_P3_U2622;
  assign new_P3_ADD_371_U8 = ~new_P3_U2624;
  assign new_P3_ADD_371_U9 = ~new_P3_U2624 | ~new_P3_ADD_371_U24;
  assign new_P3_ADD_371_U10 = ~new_P3_U2625;
  assign new_P3_ADD_371_U11 = ~new_P3_U2625 | ~new_P3_ADD_371_U28;
  assign new_P3_ADD_371_U12 = ~new_P3_U2626;
  assign new_P3_ADD_371_U13 = ~new_P3_U2626 | ~new_P3_ADD_371_U29;
  assign new_P3_ADD_371_U14 = ~new_P3_U2628;
  assign new_P3_ADD_371_U15 = ~new_P3_U2627;
  assign new_P3_ADD_371_U16 = ~new_P3_U2623;
  assign new_P3_ADD_371_U17 = ~new_P3_ADD_371_U34 | ~new_P3_ADD_371_U33;
  assign new_P3_ADD_371_U18 = ~new_P3_ADD_371_U36 | ~new_P3_ADD_371_U35;
  assign new_P3_ADD_371_U19 = ~new_P3_ADD_371_U38 | ~new_P3_ADD_371_U37;
  assign new_P3_ADD_371_U20 = ~new_P3_ADD_371_U40 | ~new_P3_ADD_371_U39;
  assign new_P3_ADD_371_U21 = ~new_P3_ADD_371_U44 | ~new_P3_ADD_371_U43;
  assign new_P3_ADD_371_U22 = new_P3_U2628 & new_P3_U2627;
  assign new_P3_ADD_371_U23 = ~new_P3_U2627 | ~new_P3_ADD_371_U30;
  assign new_P3_ADD_371_U24 = ~new_P3_ADD_371_U16 | ~new_P3_ADD_371_U26;
  assign new_P3_ADD_371_U25 = new_P3_ADD_371_U42 & new_P3_ADD_371_U41;
  assign new_P3_ADD_371_U26 = ~new_P3_U2622 | ~new_P3_U2621;
  assign new_P3_ADD_371_U27 = ~new_P3_ADD_371_U24;
  assign new_P3_ADD_371_U28 = ~new_P3_ADD_371_U9;
  assign new_P3_ADD_371_U29 = ~new_P3_ADD_371_U11;
  assign new_P3_ADD_371_U30 = ~new_P3_ADD_371_U13;
  assign new_P3_ADD_371_U31 = ~new_P3_ADD_371_U23;
  assign new_P3_ADD_371_U32 = ~new_P3_U2623 | ~new_P3_U2622 | ~new_P3_U2621;
  assign new_P3_ADD_371_U33 = ~new_P3_U2628 | ~new_P3_ADD_371_U23;
  assign new_P3_ADD_371_U34 = ~new_P3_ADD_371_U31 | ~new_P3_ADD_371_U14;
  assign new_P3_ADD_371_U35 = ~new_P3_U2627 | ~new_P3_ADD_371_U13;
  assign new_P3_ADD_371_U36 = ~new_P3_ADD_371_U30 | ~new_P3_ADD_371_U15;
  assign new_P3_ADD_371_U37 = ~new_P3_U2626 | ~new_P3_ADD_371_U11;
  assign new_P3_ADD_371_U38 = ~new_P3_ADD_371_U29 | ~new_P3_ADD_371_U12;
  assign new_P3_ADD_371_U39 = ~new_P3_U2625 | ~new_P3_ADD_371_U9;
  assign new_P3_ADD_371_U40 = ~new_P3_ADD_371_U28 | ~new_P3_ADD_371_U10;
  assign new_P3_ADD_371_U41 = ~new_P3_U2624 | ~new_P3_ADD_371_U24;
  assign new_P3_ADD_371_U42 = ~new_P3_ADD_371_U27 | ~new_P3_ADD_371_U8;
  assign new_P3_ADD_371_U43 = ~new_P3_U2622 | ~new_P3_ADD_371_U4;
  assign new_P3_ADD_371_U44 = ~new_P3_U2621 | ~new_P3_ADD_371_U7;
  assign new_P3_SUB_390_U6 = ~new_P3_SUB_390_U45 | ~new_P3_SUB_390_U44;
  assign new_P3_SUB_390_U7 = ~new_P3_SUB_390_U9 | ~new_P3_SUB_390_U46;
  assign new_P3_SUB_390_U8 = ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign new_P3_SUB_390_U9 = ~P3_INSTQUEUERD_ADDR_REG_0_ | ~new_P3_SUB_390_U18;
  assign new_P3_SUB_390_U10 = ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P3_SUB_390_U11 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_SUB_390_U12 = ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P3_SUB_390_U13 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_SUB_390_U14 = ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P3_SUB_390_U15 = ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P3_SUB_390_U16 = ~new_P3_SUB_390_U41 | ~new_P3_SUB_390_U40;
  assign new_P3_SUB_390_U17 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_SUB_390_U18 = ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P3_SUB_390_U19 = ~new_P3_SUB_390_U51 | ~new_P3_SUB_390_U50;
  assign new_P3_SUB_390_U20 = ~new_P3_SUB_390_U56 | ~new_P3_SUB_390_U55;
  assign new_P3_SUB_390_U21 = ~new_P3_SUB_390_U61 | ~new_P3_SUB_390_U60;
  assign new_P3_SUB_390_U22 = ~new_P3_SUB_390_U66 | ~new_P3_SUB_390_U65;
  assign new_P3_SUB_390_U23 = ~new_P3_SUB_390_U48 | ~new_P3_SUB_390_U47;
  assign new_P3_SUB_390_U24 = ~new_P3_SUB_390_U53 | ~new_P3_SUB_390_U52;
  assign new_P3_SUB_390_U25 = ~new_P3_SUB_390_U58 | ~new_P3_SUB_390_U57;
  assign new_P3_SUB_390_U26 = ~new_P3_SUB_390_U63 | ~new_P3_SUB_390_U62;
  assign new_P3_SUB_390_U27 = ~new_P3_SUB_390_U37 | ~new_P3_SUB_390_U36;
  assign new_P3_SUB_390_U28 = ~new_P3_SUB_390_U33 | ~new_P3_SUB_390_U32;
  assign new_P3_SUB_390_U29 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_SUB_390_U30 = ~new_P3_SUB_390_U9;
  assign new_P3_SUB_390_U31 = ~new_P3_SUB_390_U30 | ~new_P3_SUB_390_U10;
  assign new_P3_SUB_390_U32 = ~new_P3_SUB_390_U31 | ~new_P3_SUB_390_U29;
  assign new_P3_SUB_390_U33 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_390_U9;
  assign new_P3_SUB_390_U34 = ~new_P3_SUB_390_U28;
  assign new_P3_SUB_390_U35 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_390_U12;
  assign new_P3_SUB_390_U36 = ~new_P3_SUB_390_U35 | ~new_P3_SUB_390_U28;
  assign new_P3_SUB_390_U37 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_390_U11;
  assign new_P3_SUB_390_U38 = ~new_P3_SUB_390_U27;
  assign new_P3_SUB_390_U39 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_390_U14;
  assign new_P3_SUB_390_U40 = ~new_P3_SUB_390_U39 | ~new_P3_SUB_390_U27;
  assign new_P3_SUB_390_U41 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_390_U13;
  assign new_P3_SUB_390_U42 = ~new_P3_SUB_390_U16;
  assign new_P3_SUB_390_U43 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_390_U17;
  assign new_P3_SUB_390_U44 = ~new_P3_SUB_390_U42 | ~new_P3_SUB_390_U43;
  assign new_P3_SUB_390_U45 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_390_U15;
  assign new_P3_SUB_390_U46 = ~P3_INSTQUEUEWR_ADDR_REG_0_ | ~new_P3_SUB_390_U8;
  assign new_P3_SUB_390_U47 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_SUB_390_U15;
  assign new_P3_SUB_390_U48 = ~P3_INSTQUEUEWR_ADDR_REG_4_ | ~new_P3_SUB_390_U17;
  assign new_P3_SUB_390_U49 = ~new_P3_SUB_390_U23;
  assign new_P3_SUB_390_U50 = ~new_P3_SUB_390_U49 | ~new_P3_SUB_390_U42;
  assign new_P3_SUB_390_U51 = ~new_P3_SUB_390_U23 | ~new_P3_SUB_390_U16;
  assign new_P3_SUB_390_U52 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_SUB_390_U14;
  assign new_P3_SUB_390_U53 = ~P3_INSTQUEUEWR_ADDR_REG_3_ | ~new_P3_SUB_390_U13;
  assign new_P3_SUB_390_U54 = ~new_P3_SUB_390_U24;
  assign new_P3_SUB_390_U55 = ~new_P3_SUB_390_U38 | ~new_P3_SUB_390_U54;
  assign new_P3_SUB_390_U56 = ~new_P3_SUB_390_U24 | ~new_P3_SUB_390_U27;
  assign new_P3_SUB_390_U57 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_SUB_390_U12;
  assign new_P3_SUB_390_U58 = ~P3_INSTQUEUEWR_ADDR_REG_2_ | ~new_P3_SUB_390_U11;
  assign new_P3_SUB_390_U59 = ~new_P3_SUB_390_U25;
  assign new_P3_SUB_390_U60 = ~new_P3_SUB_390_U34 | ~new_P3_SUB_390_U59;
  assign new_P3_SUB_390_U61 = ~new_P3_SUB_390_U25 | ~new_P3_SUB_390_U28;
  assign new_P3_SUB_390_U62 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_SUB_390_U10;
  assign new_P3_SUB_390_U63 = ~P3_INSTQUEUEWR_ADDR_REG_1_ | ~new_P3_SUB_390_U29;
  assign new_P3_SUB_390_U64 = ~new_P3_SUB_390_U26;
  assign new_P3_SUB_390_U65 = ~new_P3_SUB_390_U64 | ~new_P3_SUB_390_U30;
  assign new_P3_SUB_390_U66 = ~new_P3_SUB_390_U26 | ~new_P3_SUB_390_U9;
  assign new_P3_SUB_357_U6 = ~new_P3_U2627;
  assign new_P3_SUB_357_U7 = ~new_P3_U2622;
  assign new_P3_SUB_357_U8 = ~new_P3_U2628;
  assign new_P3_SUB_357_U9 = ~new_P3_U2626;
  assign new_P3_SUB_357_U10 = ~new_P3_U2621;
  assign new_P3_SUB_357_U11 = ~new_P3_U2624;
  assign new_P3_SUB_357_U12 = ~new_P3_U2623;
  assign new_P3_SUB_357_U13 = ~new_P3_U2625;
  assign new_P3_ADD_495_U4 = ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_ADD_495_U5 = ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign new_P3_ADD_495_U6 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign new_P3_ADD_495_U7 = ~P3_INSTQUEUERD_ADDR_REG_3_;
  assign new_P3_ADD_495_U8 = ~new_P3_ADD_495_U16 | ~new_P3_ADD_495_U15;
  assign new_P3_ADD_495_U9 = ~new_P3_ADD_495_U18 | ~new_P3_ADD_495_U17;
  assign new_P3_ADD_495_U10 = ~new_P3_ADD_495_U20 | ~new_P3_ADD_495_U19;
  assign new_P3_ADD_495_U11 = ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign new_P3_ADD_495_U12 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_ADD_495_U13;
  assign new_P3_ADD_495_U13 = ~new_P3_ADD_495_U6;
  assign new_P3_ADD_495_U14 = ~new_P3_ADD_495_U12;
  assign new_P3_ADD_495_U15 = ~P3_INSTQUEUERD_ADDR_REG_4_ | ~new_P3_ADD_495_U12;
  assign new_P3_ADD_495_U16 = ~new_P3_ADD_495_U14 | ~new_P3_ADD_495_U11;
  assign new_P3_ADD_495_U17 = ~P3_INSTQUEUERD_ADDR_REG_3_ | ~new_P3_ADD_495_U6;
  assign new_P3_ADD_495_U18 = ~new_P3_ADD_495_U13 | ~new_P3_ADD_495_U7;
  assign new_P3_ADD_495_U19 = ~P3_INSTQUEUERD_ADDR_REG_2_ | ~new_P3_ADD_495_U4;
  assign new_P3_ADD_495_U20 = ~P3_INSTQUEUERD_ADDR_REG_1_ | ~new_P3_ADD_495_U5;
  assign new_P3_GTE_412_U6 = ~new_P3_SUB_412_U6 & ~new_P3_GTE_412_U7;
  assign new_P3_GTE_412_U7 = ~new_P3_SUB_412_U18 & ~new_P3_SUB_412_U19 & ~new_P3_SUB_412_U16 & ~new_P3_SUB_412_U17;
  assign new_P3_GTE_504_U6 = ~new_P3_SUB_504_U6 & ~new_P3_GTE_504_U7;
  assign new_P3_GTE_504_U7 = ~new_P3_SUB_504_U18 & ~new_P3_SUB_504_U19 & ~new_P3_SUB_504_U16 & ~new_P3_SUB_504_U17;
  assign new_P3_ADD_494_U4 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_494_U5 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_494_U6 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_494_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_494_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_494_U94;
  assign new_P3_ADD_494_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_494_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_494_U95;
  assign new_P3_ADD_494_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_494_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_494_U96;
  assign new_P3_ADD_494_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_494_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_494_U97;
  assign new_P3_ADD_494_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_494_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_494_U98;
  assign new_P3_ADD_494_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_494_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_494_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_494_U99;
  assign new_P3_ADD_494_U20 = ~new_P3_ADD_494_U100 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_494_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_494_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_494_U101;
  assign new_P3_ADD_494_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_494_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_494_U102;
  assign new_P3_ADD_494_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_494_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_494_U103;
  assign new_P3_ADD_494_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_494_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_494_U104;
  assign new_P3_ADD_494_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_494_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_494_U105;
  assign new_P3_ADD_494_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_494_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_494_U106;
  assign new_P3_ADD_494_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_494_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_494_U107;
  assign new_P3_ADD_494_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_494_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_494_U108;
  assign new_P3_ADD_494_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_494_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_494_U109;
  assign new_P3_ADD_494_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_494_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_494_U110;
  assign new_P3_ADD_494_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_494_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_494_U111;
  assign new_P3_ADD_494_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_494_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_494_U112;
  assign new_P3_ADD_494_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_494_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_494_U113;
  assign new_P3_ADD_494_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_494_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_494_U114;
  assign new_P3_ADD_494_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_494_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_494_U115;
  assign new_P3_ADD_494_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_494_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_494_U116;
  assign new_P3_ADD_494_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_494_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_494_U117;
  assign new_P3_ADD_494_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_494_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_494_U118;
  assign new_P3_ADD_494_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_494_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_494_U119;
  assign new_P3_ADD_494_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_494_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_494_U120;
  assign new_P3_ADD_494_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_494_U62 = ~new_P3_ADD_494_U124 | ~new_P3_ADD_494_U123;
  assign new_P3_ADD_494_U63 = ~new_P3_ADD_494_U126 | ~new_P3_ADD_494_U125;
  assign new_P3_ADD_494_U64 = ~new_P3_ADD_494_U128 | ~new_P3_ADD_494_U127;
  assign new_P3_ADD_494_U65 = ~new_P3_ADD_494_U130 | ~new_P3_ADD_494_U129;
  assign new_P3_ADD_494_U66 = ~new_P3_ADD_494_U132 | ~new_P3_ADD_494_U131;
  assign new_P3_ADD_494_U67 = ~new_P3_ADD_494_U134 | ~new_P3_ADD_494_U133;
  assign new_P3_ADD_494_U68 = ~new_P3_ADD_494_U136 | ~new_P3_ADD_494_U135;
  assign new_P3_ADD_494_U69 = ~new_P3_ADD_494_U138 | ~new_P3_ADD_494_U137;
  assign new_P3_ADD_494_U70 = ~new_P3_ADD_494_U140 | ~new_P3_ADD_494_U139;
  assign new_P3_ADD_494_U71 = ~new_P3_ADD_494_U142 | ~new_P3_ADD_494_U141;
  assign new_P3_ADD_494_U72 = ~new_P3_ADD_494_U144 | ~new_P3_ADD_494_U143;
  assign new_P3_ADD_494_U73 = ~new_P3_ADD_494_U146 | ~new_P3_ADD_494_U145;
  assign new_P3_ADD_494_U74 = ~new_P3_ADD_494_U148 | ~new_P3_ADD_494_U147;
  assign new_P3_ADD_494_U75 = ~new_P3_ADD_494_U150 | ~new_P3_ADD_494_U149;
  assign new_P3_ADD_494_U76 = ~new_P3_ADD_494_U152 | ~new_P3_ADD_494_U151;
  assign new_P3_ADD_494_U77 = ~new_P3_ADD_494_U154 | ~new_P3_ADD_494_U153;
  assign new_P3_ADD_494_U78 = ~new_P3_ADD_494_U156 | ~new_P3_ADD_494_U155;
  assign new_P3_ADD_494_U79 = ~new_P3_ADD_494_U158 | ~new_P3_ADD_494_U157;
  assign new_P3_ADD_494_U80 = ~new_P3_ADD_494_U160 | ~new_P3_ADD_494_U159;
  assign new_P3_ADD_494_U81 = ~new_P3_ADD_494_U162 | ~new_P3_ADD_494_U161;
  assign new_P3_ADD_494_U82 = ~new_P3_ADD_494_U164 | ~new_P3_ADD_494_U163;
  assign new_P3_ADD_494_U83 = ~new_P3_ADD_494_U166 | ~new_P3_ADD_494_U165;
  assign new_P3_ADD_494_U84 = ~new_P3_ADD_494_U168 | ~new_P3_ADD_494_U167;
  assign new_P3_ADD_494_U85 = ~new_P3_ADD_494_U170 | ~new_P3_ADD_494_U169;
  assign new_P3_ADD_494_U86 = ~new_P3_ADD_494_U172 | ~new_P3_ADD_494_U171;
  assign new_P3_ADD_494_U87 = ~new_P3_ADD_494_U174 | ~new_P3_ADD_494_U173;
  assign new_P3_ADD_494_U88 = ~new_P3_ADD_494_U176 | ~new_P3_ADD_494_U175;
  assign new_P3_ADD_494_U89 = ~new_P3_ADD_494_U178 | ~new_P3_ADD_494_U177;
  assign new_P3_ADD_494_U90 = ~new_P3_ADD_494_U180 | ~new_P3_ADD_494_U179;
  assign new_P3_ADD_494_U91 = ~new_P3_ADD_494_U182 | ~new_P3_ADD_494_U181;
  assign new_P3_ADD_494_U92 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_494_U93 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_494_U121;
  assign new_P3_ADD_494_U94 = ~new_P3_ADD_494_U6;
  assign new_P3_ADD_494_U95 = ~new_P3_ADD_494_U8;
  assign new_P3_ADD_494_U96 = ~new_P3_ADD_494_U10;
  assign new_P3_ADD_494_U97 = ~new_P3_ADD_494_U12;
  assign new_P3_ADD_494_U98 = ~new_P3_ADD_494_U14;
  assign new_P3_ADD_494_U99 = ~new_P3_ADD_494_U16;
  assign new_P3_ADD_494_U100 = ~new_P3_ADD_494_U19;
  assign new_P3_ADD_494_U101 = ~new_P3_ADD_494_U20;
  assign new_P3_ADD_494_U102 = ~new_P3_ADD_494_U22;
  assign new_P3_ADD_494_U103 = ~new_P3_ADD_494_U24;
  assign new_P3_ADD_494_U104 = ~new_P3_ADD_494_U26;
  assign new_P3_ADD_494_U105 = ~new_P3_ADD_494_U28;
  assign new_P3_ADD_494_U106 = ~new_P3_ADD_494_U30;
  assign new_P3_ADD_494_U107 = ~new_P3_ADD_494_U32;
  assign new_P3_ADD_494_U108 = ~new_P3_ADD_494_U34;
  assign new_P3_ADD_494_U109 = ~new_P3_ADD_494_U36;
  assign new_P3_ADD_494_U110 = ~new_P3_ADD_494_U38;
  assign new_P3_ADD_494_U111 = ~new_P3_ADD_494_U40;
  assign new_P3_ADD_494_U112 = ~new_P3_ADD_494_U42;
  assign new_P3_ADD_494_U113 = ~new_P3_ADD_494_U44;
  assign new_P3_ADD_494_U114 = ~new_P3_ADD_494_U46;
  assign new_P3_ADD_494_U115 = ~new_P3_ADD_494_U48;
  assign new_P3_ADD_494_U116 = ~new_P3_ADD_494_U50;
  assign new_P3_ADD_494_U117 = ~new_P3_ADD_494_U52;
  assign new_P3_ADD_494_U118 = ~new_P3_ADD_494_U54;
  assign new_P3_ADD_494_U119 = ~new_P3_ADD_494_U56;
  assign new_P3_ADD_494_U120 = ~new_P3_ADD_494_U58;
  assign new_P3_ADD_494_U121 = ~new_P3_ADD_494_U60;
  assign new_P3_ADD_494_U122 = ~new_P3_ADD_494_U93;
  assign new_P3_ADD_494_U123 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_494_U19;
  assign new_P3_ADD_494_U124 = ~new_P3_ADD_494_U100 | ~new_P3_ADD_494_U18;
  assign new_P3_ADD_494_U125 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_494_U16;
  assign new_P3_ADD_494_U126 = ~new_P3_ADD_494_U99 | ~new_P3_ADD_494_U17;
  assign new_P3_ADD_494_U127 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_494_U14;
  assign new_P3_ADD_494_U128 = ~new_P3_ADD_494_U98 | ~new_P3_ADD_494_U15;
  assign new_P3_ADD_494_U129 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_494_U12;
  assign new_P3_ADD_494_U130 = ~new_P3_ADD_494_U97 | ~new_P3_ADD_494_U13;
  assign new_P3_ADD_494_U131 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_494_U10;
  assign new_P3_ADD_494_U132 = ~new_P3_ADD_494_U96 | ~new_P3_ADD_494_U11;
  assign new_P3_ADD_494_U133 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_494_U8;
  assign new_P3_ADD_494_U134 = ~new_P3_ADD_494_U95 | ~new_P3_ADD_494_U9;
  assign new_P3_ADD_494_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_494_U6;
  assign new_P3_ADD_494_U136 = ~new_P3_ADD_494_U94 | ~new_P3_ADD_494_U7;
  assign new_P3_ADD_494_U137 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_494_U93;
  assign new_P3_ADD_494_U138 = ~new_P3_ADD_494_U122 | ~new_P3_ADD_494_U92;
  assign new_P3_ADD_494_U139 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_494_U60;
  assign new_P3_ADD_494_U140 = ~new_P3_ADD_494_U121 | ~new_P3_ADD_494_U61;
  assign new_P3_ADD_494_U141 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_494_U4;
  assign new_P3_ADD_494_U142 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_494_U5;
  assign new_P3_ADD_494_U143 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_494_U58;
  assign new_P3_ADD_494_U144 = ~new_P3_ADD_494_U120 | ~new_P3_ADD_494_U59;
  assign new_P3_ADD_494_U145 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_494_U56;
  assign new_P3_ADD_494_U146 = ~new_P3_ADD_494_U119 | ~new_P3_ADD_494_U57;
  assign new_P3_ADD_494_U147 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_494_U54;
  assign new_P3_ADD_494_U148 = ~new_P3_ADD_494_U118 | ~new_P3_ADD_494_U55;
  assign new_P3_ADD_494_U149 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_494_U52;
  assign new_P3_ADD_494_U150 = ~new_P3_ADD_494_U117 | ~new_P3_ADD_494_U53;
  assign new_P3_ADD_494_U151 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_494_U50;
  assign new_P3_ADD_494_U152 = ~new_P3_ADD_494_U116 | ~new_P3_ADD_494_U51;
  assign new_P3_ADD_494_U153 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_494_U48;
  assign new_P3_ADD_494_U154 = ~new_P3_ADD_494_U115 | ~new_P3_ADD_494_U49;
  assign new_P3_ADD_494_U155 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_494_U46;
  assign new_P3_ADD_494_U156 = ~new_P3_ADD_494_U114 | ~new_P3_ADD_494_U47;
  assign new_P3_ADD_494_U157 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_494_U44;
  assign new_P3_ADD_494_U158 = ~new_P3_ADD_494_U113 | ~new_P3_ADD_494_U45;
  assign new_P3_ADD_494_U159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_494_U42;
  assign new_P3_ADD_494_U160 = ~new_P3_ADD_494_U112 | ~new_P3_ADD_494_U43;
  assign new_P3_ADD_494_U161 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_494_U40;
  assign new_P3_ADD_494_U162 = ~new_P3_ADD_494_U111 | ~new_P3_ADD_494_U41;
  assign new_P3_ADD_494_U163 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_494_U38;
  assign new_P3_ADD_494_U164 = ~new_P3_ADD_494_U110 | ~new_P3_ADD_494_U39;
  assign new_P3_ADD_494_U165 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_494_U36;
  assign new_P3_ADD_494_U166 = ~new_P3_ADD_494_U109 | ~new_P3_ADD_494_U37;
  assign new_P3_ADD_494_U167 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_494_U34;
  assign new_P3_ADD_494_U168 = ~new_P3_ADD_494_U108 | ~new_P3_ADD_494_U35;
  assign new_P3_ADD_494_U169 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_494_U32;
  assign new_P3_ADD_494_U170 = ~new_P3_ADD_494_U107 | ~new_P3_ADD_494_U33;
  assign new_P3_ADD_494_U171 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_494_U30;
  assign new_P3_ADD_494_U172 = ~new_P3_ADD_494_U106 | ~new_P3_ADD_494_U31;
  assign new_P3_ADD_494_U173 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_494_U28;
  assign new_P3_ADD_494_U174 = ~new_P3_ADD_494_U105 | ~new_P3_ADD_494_U29;
  assign new_P3_ADD_494_U175 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_494_U26;
  assign new_P3_ADD_494_U176 = ~new_P3_ADD_494_U104 | ~new_P3_ADD_494_U27;
  assign new_P3_ADD_494_U177 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_494_U24;
  assign new_P3_ADD_494_U178 = ~new_P3_ADD_494_U103 | ~new_P3_ADD_494_U25;
  assign new_P3_ADD_494_U179 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_494_U22;
  assign new_P3_ADD_494_U180 = ~new_P3_ADD_494_U102 | ~new_P3_ADD_494_U23;
  assign new_P3_ADD_494_U181 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_494_U20;
  assign new_P3_ADD_494_U182 = ~new_P3_ADD_494_U101 | ~new_P3_ADD_494_U21;
  assign new_P3_ADD_536_U4 = ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_536_U5 = ~P3_INSTADDRPOINTER_REG_2_;
  assign new_P3_ADD_536_U6 = ~P3_INSTADDRPOINTER_REG_2_ | ~P3_INSTADDRPOINTER_REG_1_;
  assign new_P3_ADD_536_U7 = ~P3_INSTADDRPOINTER_REG_3_;
  assign new_P3_ADD_536_U8 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_536_U94;
  assign new_P3_ADD_536_U9 = ~P3_INSTADDRPOINTER_REG_4_;
  assign new_P3_ADD_536_U10 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_536_U95;
  assign new_P3_ADD_536_U11 = ~P3_INSTADDRPOINTER_REG_5_;
  assign new_P3_ADD_536_U12 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_536_U96;
  assign new_P3_ADD_536_U13 = ~P3_INSTADDRPOINTER_REG_6_;
  assign new_P3_ADD_536_U14 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_536_U97;
  assign new_P3_ADD_536_U15 = ~P3_INSTADDRPOINTER_REG_7_;
  assign new_P3_ADD_536_U16 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_536_U98;
  assign new_P3_ADD_536_U17 = ~P3_INSTADDRPOINTER_REG_8_;
  assign new_P3_ADD_536_U18 = ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_536_U19 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_536_U99;
  assign new_P3_ADD_536_U20 = ~new_P3_ADD_536_U100 | ~P3_INSTADDRPOINTER_REG_9_;
  assign new_P3_ADD_536_U21 = ~P3_INSTADDRPOINTER_REG_10_;
  assign new_P3_ADD_536_U22 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_536_U101;
  assign new_P3_ADD_536_U23 = ~P3_INSTADDRPOINTER_REG_11_;
  assign new_P3_ADD_536_U24 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_536_U102;
  assign new_P3_ADD_536_U25 = ~P3_INSTADDRPOINTER_REG_12_;
  assign new_P3_ADD_536_U26 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_536_U103;
  assign new_P3_ADD_536_U27 = ~P3_INSTADDRPOINTER_REG_13_;
  assign new_P3_ADD_536_U28 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_536_U104;
  assign new_P3_ADD_536_U29 = ~P3_INSTADDRPOINTER_REG_14_;
  assign new_P3_ADD_536_U30 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_536_U105;
  assign new_P3_ADD_536_U31 = ~P3_INSTADDRPOINTER_REG_15_;
  assign new_P3_ADD_536_U32 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_536_U106;
  assign new_P3_ADD_536_U33 = ~P3_INSTADDRPOINTER_REG_16_;
  assign new_P3_ADD_536_U34 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_536_U107;
  assign new_P3_ADD_536_U35 = ~P3_INSTADDRPOINTER_REG_17_;
  assign new_P3_ADD_536_U36 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_536_U108;
  assign new_P3_ADD_536_U37 = ~P3_INSTADDRPOINTER_REG_18_;
  assign new_P3_ADD_536_U38 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_536_U109;
  assign new_P3_ADD_536_U39 = ~P3_INSTADDRPOINTER_REG_19_;
  assign new_P3_ADD_536_U40 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_536_U110;
  assign new_P3_ADD_536_U41 = ~P3_INSTADDRPOINTER_REG_20_;
  assign new_P3_ADD_536_U42 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_536_U111;
  assign new_P3_ADD_536_U43 = ~P3_INSTADDRPOINTER_REG_21_;
  assign new_P3_ADD_536_U44 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_536_U112;
  assign new_P3_ADD_536_U45 = ~P3_INSTADDRPOINTER_REG_22_;
  assign new_P3_ADD_536_U46 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_536_U113;
  assign new_P3_ADD_536_U47 = ~P3_INSTADDRPOINTER_REG_23_;
  assign new_P3_ADD_536_U48 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_536_U114;
  assign new_P3_ADD_536_U49 = ~P3_INSTADDRPOINTER_REG_24_;
  assign new_P3_ADD_536_U50 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_536_U115;
  assign new_P3_ADD_536_U51 = ~P3_INSTADDRPOINTER_REG_25_;
  assign new_P3_ADD_536_U52 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_536_U116;
  assign new_P3_ADD_536_U53 = ~P3_INSTADDRPOINTER_REG_26_;
  assign new_P3_ADD_536_U54 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_536_U117;
  assign new_P3_ADD_536_U55 = ~P3_INSTADDRPOINTER_REG_27_;
  assign new_P3_ADD_536_U56 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_536_U118;
  assign new_P3_ADD_536_U57 = ~P3_INSTADDRPOINTER_REG_28_;
  assign new_P3_ADD_536_U58 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_536_U119;
  assign new_P3_ADD_536_U59 = ~P3_INSTADDRPOINTER_REG_29_;
  assign new_P3_ADD_536_U60 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_536_U120;
  assign new_P3_ADD_536_U61 = ~P3_INSTADDRPOINTER_REG_30_;
  assign new_P3_ADD_536_U62 = ~new_P3_ADD_536_U124 | ~new_P3_ADD_536_U123;
  assign new_P3_ADD_536_U63 = ~new_P3_ADD_536_U126 | ~new_P3_ADD_536_U125;
  assign new_P3_ADD_536_U64 = ~new_P3_ADD_536_U128 | ~new_P3_ADD_536_U127;
  assign new_P3_ADD_536_U65 = ~new_P3_ADD_536_U130 | ~new_P3_ADD_536_U129;
  assign new_P3_ADD_536_U66 = ~new_P3_ADD_536_U132 | ~new_P3_ADD_536_U131;
  assign new_P3_ADD_536_U67 = ~new_P3_ADD_536_U134 | ~new_P3_ADD_536_U133;
  assign new_P3_ADD_536_U68 = ~new_P3_ADD_536_U136 | ~new_P3_ADD_536_U135;
  assign new_P3_ADD_536_U69 = ~new_P3_ADD_536_U138 | ~new_P3_ADD_536_U137;
  assign new_P3_ADD_536_U70 = ~new_P3_ADD_536_U140 | ~new_P3_ADD_536_U139;
  assign new_P3_ADD_536_U71 = ~new_P3_ADD_536_U142 | ~new_P3_ADD_536_U141;
  assign new_P3_ADD_536_U72 = ~new_P3_ADD_536_U144 | ~new_P3_ADD_536_U143;
  assign new_P3_ADD_536_U73 = ~new_P3_ADD_536_U146 | ~new_P3_ADD_536_U145;
  assign new_P3_ADD_536_U74 = ~new_P3_ADD_536_U148 | ~new_P3_ADD_536_U147;
  assign new_P3_ADD_536_U75 = ~new_P3_ADD_536_U150 | ~new_P3_ADD_536_U149;
  assign new_P3_ADD_536_U76 = ~new_P3_ADD_536_U152 | ~new_P3_ADD_536_U151;
  assign new_P3_ADD_536_U77 = ~new_P3_ADD_536_U154 | ~new_P3_ADD_536_U153;
  assign new_P3_ADD_536_U78 = ~new_P3_ADD_536_U156 | ~new_P3_ADD_536_U155;
  assign new_P3_ADD_536_U79 = ~new_P3_ADD_536_U158 | ~new_P3_ADD_536_U157;
  assign new_P3_ADD_536_U80 = ~new_P3_ADD_536_U160 | ~new_P3_ADD_536_U159;
  assign new_P3_ADD_536_U81 = ~new_P3_ADD_536_U162 | ~new_P3_ADD_536_U161;
  assign new_P3_ADD_536_U82 = ~new_P3_ADD_536_U164 | ~new_P3_ADD_536_U163;
  assign new_P3_ADD_536_U83 = ~new_P3_ADD_536_U166 | ~new_P3_ADD_536_U165;
  assign new_P3_ADD_536_U84 = ~new_P3_ADD_536_U168 | ~new_P3_ADD_536_U167;
  assign new_P3_ADD_536_U85 = ~new_P3_ADD_536_U170 | ~new_P3_ADD_536_U169;
  assign new_P3_ADD_536_U86 = ~new_P3_ADD_536_U172 | ~new_P3_ADD_536_U171;
  assign new_P3_ADD_536_U87 = ~new_P3_ADD_536_U174 | ~new_P3_ADD_536_U173;
  assign new_P3_ADD_536_U88 = ~new_P3_ADD_536_U176 | ~new_P3_ADD_536_U175;
  assign new_P3_ADD_536_U89 = ~new_P3_ADD_536_U178 | ~new_P3_ADD_536_U177;
  assign new_P3_ADD_536_U90 = ~new_P3_ADD_536_U180 | ~new_P3_ADD_536_U179;
  assign new_P3_ADD_536_U91 = ~new_P3_ADD_536_U182 | ~new_P3_ADD_536_U181;
  assign new_P3_ADD_536_U92 = ~P3_INSTADDRPOINTER_REG_31_;
  assign new_P3_ADD_536_U93 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_536_U121;
  assign new_P3_ADD_536_U94 = ~new_P3_ADD_536_U6;
  assign new_P3_ADD_536_U95 = ~new_P3_ADD_536_U8;
  assign new_P3_ADD_536_U96 = ~new_P3_ADD_536_U10;
  assign new_P3_ADD_536_U97 = ~new_P3_ADD_536_U12;
  assign new_P3_ADD_536_U98 = ~new_P3_ADD_536_U14;
  assign new_P3_ADD_536_U99 = ~new_P3_ADD_536_U16;
  assign new_P3_ADD_536_U100 = ~new_P3_ADD_536_U19;
  assign new_P3_ADD_536_U101 = ~new_P3_ADD_536_U20;
  assign new_P3_ADD_536_U102 = ~new_P3_ADD_536_U22;
  assign new_P3_ADD_536_U103 = ~new_P3_ADD_536_U24;
  assign new_P3_ADD_536_U104 = ~new_P3_ADD_536_U26;
  assign new_P3_ADD_536_U105 = ~new_P3_ADD_536_U28;
  assign new_P3_ADD_536_U106 = ~new_P3_ADD_536_U30;
  assign new_P3_ADD_536_U107 = ~new_P3_ADD_536_U32;
  assign new_P3_ADD_536_U108 = ~new_P3_ADD_536_U34;
  assign new_P3_ADD_536_U109 = ~new_P3_ADD_536_U36;
  assign new_P3_ADD_536_U110 = ~new_P3_ADD_536_U38;
  assign new_P3_ADD_536_U111 = ~new_P3_ADD_536_U40;
  assign new_P3_ADD_536_U112 = ~new_P3_ADD_536_U42;
  assign new_P3_ADD_536_U113 = ~new_P3_ADD_536_U44;
  assign new_P3_ADD_536_U114 = ~new_P3_ADD_536_U46;
  assign new_P3_ADD_536_U115 = ~new_P3_ADD_536_U48;
  assign new_P3_ADD_536_U116 = ~new_P3_ADD_536_U50;
  assign new_P3_ADD_536_U117 = ~new_P3_ADD_536_U52;
  assign new_P3_ADD_536_U118 = ~new_P3_ADD_536_U54;
  assign new_P3_ADD_536_U119 = ~new_P3_ADD_536_U56;
  assign new_P3_ADD_536_U120 = ~new_P3_ADD_536_U58;
  assign new_P3_ADD_536_U121 = ~new_P3_ADD_536_U60;
  assign new_P3_ADD_536_U122 = ~new_P3_ADD_536_U93;
  assign new_P3_ADD_536_U123 = ~P3_INSTADDRPOINTER_REG_9_ | ~new_P3_ADD_536_U19;
  assign new_P3_ADD_536_U124 = ~new_P3_ADD_536_U100 | ~new_P3_ADD_536_U18;
  assign new_P3_ADD_536_U125 = ~P3_INSTADDRPOINTER_REG_8_ | ~new_P3_ADD_536_U16;
  assign new_P3_ADD_536_U126 = ~new_P3_ADD_536_U99 | ~new_P3_ADD_536_U17;
  assign new_P3_ADD_536_U127 = ~P3_INSTADDRPOINTER_REG_7_ | ~new_P3_ADD_536_U14;
  assign new_P3_ADD_536_U128 = ~new_P3_ADD_536_U98 | ~new_P3_ADD_536_U15;
  assign new_P3_ADD_536_U129 = ~P3_INSTADDRPOINTER_REG_6_ | ~new_P3_ADD_536_U12;
  assign new_P3_ADD_536_U130 = ~new_P3_ADD_536_U97 | ~new_P3_ADD_536_U13;
  assign new_P3_ADD_536_U131 = ~P3_INSTADDRPOINTER_REG_5_ | ~new_P3_ADD_536_U10;
  assign new_P3_ADD_536_U132 = ~new_P3_ADD_536_U96 | ~new_P3_ADD_536_U11;
  assign new_P3_ADD_536_U133 = ~P3_INSTADDRPOINTER_REG_4_ | ~new_P3_ADD_536_U8;
  assign new_P3_ADD_536_U134 = ~new_P3_ADD_536_U95 | ~new_P3_ADD_536_U9;
  assign new_P3_ADD_536_U135 = ~P3_INSTADDRPOINTER_REG_3_ | ~new_P3_ADD_536_U6;
  assign new_P3_ADD_536_U136 = ~new_P3_ADD_536_U94 | ~new_P3_ADD_536_U7;
  assign new_P3_ADD_536_U137 = ~P3_INSTADDRPOINTER_REG_31_ | ~new_P3_ADD_536_U93;
  assign new_P3_ADD_536_U138 = ~new_P3_ADD_536_U122 | ~new_P3_ADD_536_U92;
  assign new_P3_ADD_536_U139 = ~P3_INSTADDRPOINTER_REG_30_ | ~new_P3_ADD_536_U60;
  assign new_P3_ADD_536_U140 = ~new_P3_ADD_536_U121 | ~new_P3_ADD_536_U61;
  assign new_P3_ADD_536_U141 = ~P3_INSTADDRPOINTER_REG_2_ | ~new_P3_ADD_536_U4;
  assign new_P3_ADD_536_U142 = ~P3_INSTADDRPOINTER_REG_1_ | ~new_P3_ADD_536_U5;
  assign new_P3_ADD_536_U143 = ~P3_INSTADDRPOINTER_REG_29_ | ~new_P3_ADD_536_U58;
  assign new_P3_ADD_536_U144 = ~new_P3_ADD_536_U120 | ~new_P3_ADD_536_U59;
  assign new_P3_ADD_536_U145 = ~P3_INSTADDRPOINTER_REG_28_ | ~new_P3_ADD_536_U56;
  assign new_P3_ADD_536_U146 = ~new_P3_ADD_536_U119 | ~new_P3_ADD_536_U57;
  assign new_P3_ADD_536_U147 = ~P3_INSTADDRPOINTER_REG_27_ | ~new_P3_ADD_536_U54;
  assign new_P3_ADD_536_U148 = ~new_P3_ADD_536_U118 | ~new_P3_ADD_536_U55;
  assign new_P3_ADD_536_U149 = ~P3_INSTADDRPOINTER_REG_26_ | ~new_P3_ADD_536_U52;
  assign new_P3_ADD_536_U150 = ~new_P3_ADD_536_U117 | ~new_P3_ADD_536_U53;
  assign new_P3_ADD_536_U151 = ~P3_INSTADDRPOINTER_REG_25_ | ~new_P3_ADD_536_U50;
  assign new_P3_ADD_536_U152 = ~new_P3_ADD_536_U116 | ~new_P3_ADD_536_U51;
  assign new_P3_ADD_536_U153 = ~P3_INSTADDRPOINTER_REG_24_ | ~new_P3_ADD_536_U48;
  assign new_P3_ADD_536_U154 = ~new_P3_ADD_536_U115 | ~new_P3_ADD_536_U49;
  assign new_P3_ADD_536_U155 = ~P3_INSTADDRPOINTER_REG_23_ | ~new_P3_ADD_536_U46;
  assign new_P3_ADD_536_U156 = ~new_P3_ADD_536_U114 | ~new_P3_ADD_536_U47;
  assign new_P3_ADD_536_U157 = ~P3_INSTADDRPOINTER_REG_22_ | ~new_P3_ADD_536_U44;
  assign new_P3_ADD_536_U158 = ~new_P3_ADD_536_U113 | ~new_P3_ADD_536_U45;
  assign new_P3_ADD_536_U159 = ~P3_INSTADDRPOINTER_REG_21_ | ~new_P3_ADD_536_U42;
  assign new_P3_ADD_536_U160 = ~new_P3_ADD_536_U112 | ~new_P3_ADD_536_U43;
  assign new_P3_ADD_536_U161 = ~P3_INSTADDRPOINTER_REG_20_ | ~new_P3_ADD_536_U40;
  assign new_P3_ADD_536_U162 = ~new_P3_ADD_536_U111 | ~new_P3_ADD_536_U41;
  assign new_P3_ADD_536_U163 = ~P3_INSTADDRPOINTER_REG_19_ | ~new_P3_ADD_536_U38;
  assign new_P3_ADD_536_U164 = ~new_P3_ADD_536_U110 | ~new_P3_ADD_536_U39;
  assign new_P3_ADD_536_U165 = ~P3_INSTADDRPOINTER_REG_18_ | ~new_P3_ADD_536_U36;
  assign new_P3_ADD_536_U166 = ~new_P3_ADD_536_U109 | ~new_P3_ADD_536_U37;
  assign new_P3_ADD_536_U167 = ~P3_INSTADDRPOINTER_REG_17_ | ~new_P3_ADD_536_U34;
  assign new_P3_ADD_536_U168 = ~new_P3_ADD_536_U108 | ~new_P3_ADD_536_U35;
  assign new_P3_ADD_536_U169 = ~P3_INSTADDRPOINTER_REG_16_ | ~new_P3_ADD_536_U32;
  assign new_P3_ADD_536_U170 = ~new_P3_ADD_536_U107 | ~new_P3_ADD_536_U33;
  assign new_P3_ADD_536_U171 = ~P3_INSTADDRPOINTER_REG_15_ | ~new_P3_ADD_536_U30;
  assign new_P3_ADD_536_U172 = ~new_P3_ADD_536_U106 | ~new_P3_ADD_536_U31;
  assign new_P3_ADD_536_U173 = ~P3_INSTADDRPOINTER_REG_14_ | ~new_P3_ADD_536_U28;
  assign new_P3_ADD_536_U174 = ~new_P3_ADD_536_U105 | ~new_P3_ADD_536_U29;
  assign new_P3_ADD_536_U175 = ~P3_INSTADDRPOINTER_REG_13_ | ~new_P3_ADD_536_U26;
  assign new_P3_ADD_536_U176 = ~new_P3_ADD_536_U104 | ~new_P3_ADD_536_U27;
  assign new_P3_ADD_536_U177 = ~P3_INSTADDRPOINTER_REG_12_ | ~new_P3_ADD_536_U24;
  assign new_P3_ADD_536_U178 = ~new_P3_ADD_536_U103 | ~new_P3_ADD_536_U25;
  assign new_P3_ADD_536_U179 = ~P3_INSTADDRPOINTER_REG_11_ | ~new_P3_ADD_536_U22;
  assign new_P3_ADD_536_U180 = ~new_P3_ADD_536_U102 | ~new_P3_ADD_536_U23;
  assign new_P3_ADD_536_U181 = ~P3_INSTADDRPOINTER_REG_10_ | ~new_P3_ADD_536_U20;
  assign new_P3_ADD_536_U182 = ~new_P3_ADD_536_U101 | ~new_P3_ADD_536_U21;
  assign new_P3_ADD_402_1132_U4 = ~new_P3_U2613;
  assign new_P3_ADD_402_1132_U5 = ~new_P3_U3069;
  assign new_P3_ADD_402_1132_U6 = ~new_P3_U3069 | ~new_P3_U2613;
  assign new_P3_ADD_402_1132_U7 = ~new_P3_U2614;
  assign new_P3_ADD_402_1132_U8 = ~new_P3_U2614 | ~new_P3_ADD_402_1132_U28;
  assign new_P3_ADD_402_1132_U9 = ~new_P3_U2615;
  assign new_P3_ADD_402_1132_U10 = ~new_P3_U2615 | ~new_P3_ADD_402_1132_U29;
  assign new_P3_ADD_402_1132_U11 = ~new_P3_U2616;
  assign new_P3_ADD_402_1132_U12 = ~new_P3_U2616 | ~new_P3_ADD_402_1132_U30;
  assign new_P3_ADD_402_1132_U13 = ~new_P3_U2617;
  assign new_P3_ADD_402_1132_U14 = ~new_P3_U2617 | ~new_P3_ADD_402_1132_U31;
  assign new_P3_ADD_402_1132_U15 = ~new_P3_U2618;
  assign new_P3_ADD_402_1132_U16 = ~new_P3_U2618 | ~new_P3_ADD_402_1132_U32;
  assign new_P3_ADD_402_1132_U17 = ~new_P3_U2619;
  assign new_P3_ADD_402_1132_U18 = ~new_P3_ADD_402_1132_U36 | ~new_P3_ADD_402_1132_U35;
  assign new_P3_ADD_402_1132_U19 = ~new_P3_ADD_402_1132_U38 | ~new_P3_ADD_402_1132_U37;
  assign new_P3_ADD_402_1132_U20 = ~new_P3_ADD_402_1132_U40 | ~new_P3_ADD_402_1132_U39;
  assign new_P3_ADD_402_1132_U21 = ~new_P3_ADD_402_1132_U42 | ~new_P3_ADD_402_1132_U41;
  assign new_P3_ADD_402_1132_U22 = ~new_P3_ADD_402_1132_U44 | ~new_P3_ADD_402_1132_U43;
  assign new_P3_ADD_402_1132_U23 = ~new_P3_ADD_402_1132_U46 | ~new_P3_ADD_402_1132_U45;
  assign new_P3_ADD_402_1132_U24 = ~new_P3_ADD_402_1132_U48 | ~new_P3_ADD_402_1132_U47;
  assign new_P3_ADD_402_1132_U25 = ~new_P3_ADD_402_1132_U50 | ~new_P3_ADD_402_1132_U49;
  assign new_P3_ADD_402_1132_U26 = ~new_P3_U2620;
  assign new_P3_ADD_402_1132_U27 = ~new_P3_U2619 | ~new_P3_ADD_402_1132_U33;
  assign new_P3_ADD_402_1132_U28 = ~new_P3_ADD_402_1132_U6;
  assign new_P3_ADD_402_1132_U29 = ~new_P3_ADD_402_1132_U8;
  assign new_P3_ADD_402_1132_U30 = ~new_P3_ADD_402_1132_U10;
  assign new_P3_ADD_402_1132_U31 = ~new_P3_ADD_402_1132_U12;
  assign new_P3_ADD_402_1132_U32 = ~new_P3_ADD_402_1132_U14;
  assign new_P3_ADD_402_1132_U33 = ~new_P3_ADD_402_1132_U16;
  assign new_P3_ADD_402_1132_U34 = ~new_P3_ADD_402_1132_U27;
  assign new_P3_ADD_402_1132_U35 = ~new_P3_U2620 | ~new_P3_ADD_402_1132_U27;
  assign new_P3_ADD_402_1132_U36 = ~new_P3_ADD_402_1132_U34 | ~new_P3_ADD_402_1132_U26;
  assign new_P3_ADD_402_1132_U37 = ~new_P3_U2619 | ~new_P3_ADD_402_1132_U16;
  assign new_P3_ADD_402_1132_U38 = ~new_P3_ADD_402_1132_U33 | ~new_P3_ADD_402_1132_U17;
  assign new_P3_ADD_402_1132_U39 = ~new_P3_U2618 | ~new_P3_ADD_402_1132_U14;
  assign new_P3_ADD_402_1132_U40 = ~new_P3_ADD_402_1132_U32 | ~new_P3_ADD_402_1132_U15;
  assign new_P3_ADD_402_1132_U41 = ~new_P3_U2617 | ~new_P3_ADD_402_1132_U12;
  assign new_P3_ADD_402_1132_U42 = ~new_P3_ADD_402_1132_U31 | ~new_P3_ADD_402_1132_U13;
  assign new_P3_ADD_402_1132_U43 = ~new_P3_U2616 | ~new_P3_ADD_402_1132_U10;
  assign new_P3_ADD_402_1132_U44 = ~new_P3_ADD_402_1132_U30 | ~new_P3_ADD_402_1132_U11;
  assign new_P3_ADD_402_1132_U45 = ~new_P3_U2615 | ~new_P3_ADD_402_1132_U8;
  assign new_P3_ADD_402_1132_U46 = ~new_P3_ADD_402_1132_U29 | ~new_P3_ADD_402_1132_U9;
  assign new_P3_ADD_402_1132_U47 = ~new_P3_U2614 | ~new_P3_ADD_402_1132_U6;
  assign new_P3_ADD_402_1132_U48 = ~new_P3_ADD_402_1132_U28 | ~new_P3_ADD_402_1132_U7;
  assign new_P3_ADD_402_1132_U49 = ~new_P3_U3069 | ~new_P3_ADD_402_1132_U4;
  assign new_P3_ADD_402_1132_U50 = ~new_P3_U2613 | ~new_P3_ADD_402_1132_U5;
  assign new_P2_R2099_U5 = ~new_P2_R2099_U107 | ~new_P2_R2099_U148;
  assign new_P2_R2099_U6 = ~new_P2_U2747;
  assign new_P2_R2099_U7 = ~new_P2_U2751;
  assign new_P2_R2099_U8 = ~new_P2_U2750;
  assign new_P2_R2099_U9 = ~new_P2_U2746;
  assign new_P2_R2099_U10 = ~new_P2_U2749;
  assign new_P2_R2099_U11 = ~new_P2_U2745;
  assign new_P2_R2099_U12 = ~new_P2_U2748;
  assign new_P2_R2099_U13 = ~new_P2_U2744;
  assign new_P2_R2099_U14 = ~new_P2_U2743;
  assign new_P2_R2099_U15 = ~new_P2_U2743 | ~new_P2_R2099_U97;
  assign new_P2_R2099_U16 = ~new_P2_U2742;
  assign new_P2_R2099_U17 = ~new_P2_U2742 | ~new_P2_R2099_U120;
  assign new_P2_R2099_U18 = ~new_P2_U2741;
  assign new_P2_R2099_U19 = ~new_P2_U2741 | ~new_P2_R2099_U121;
  assign new_P2_R2099_U20 = ~new_P2_U2740;
  assign new_P2_R2099_U21 = ~new_P2_U2740 | ~new_P2_R2099_U122;
  assign new_P2_R2099_U22 = ~new_P2_U2739;
  assign new_P2_R2099_U23 = ~new_P2_U2738;
  assign new_P2_R2099_U24 = ~new_P2_U2739 | ~new_P2_R2099_U123;
  assign new_P2_R2099_U25 = ~new_P2_R2099_U124 | ~new_P2_U2738;
  assign new_P2_R2099_U26 = ~new_P2_U2737;
  assign new_P2_R2099_U27 = ~new_P2_U2737 | ~new_P2_R2099_U125;
  assign new_P2_R2099_U28 = ~new_P2_U2736;
  assign new_P2_R2099_U29 = ~new_P2_U2736 | ~new_P2_R2099_U126;
  assign new_P2_R2099_U30 = ~new_P2_U2735;
  assign new_P2_R2099_U31 = ~new_P2_U2735 | ~new_P2_R2099_U127;
  assign new_P2_R2099_U32 = ~new_P2_U2734;
  assign new_P2_R2099_U33 = ~new_P2_U2734 | ~new_P2_R2099_U128;
  assign new_P2_R2099_U34 = ~new_P2_U2733;
  assign new_P2_R2099_U35 = ~new_P2_U2733 | ~new_P2_R2099_U129;
  assign new_P2_R2099_U36 = ~new_P2_U2732;
  assign new_P2_R2099_U37 = ~new_P2_U2732 | ~new_P2_R2099_U130;
  assign new_P2_R2099_U38 = ~new_P2_U2731;
  assign new_P2_R2099_U39 = ~new_P2_U2731 | ~new_P2_R2099_U131;
  assign new_P2_R2099_U40 = ~new_P2_U2730;
  assign new_P2_R2099_U41 = ~new_P2_U2730 | ~new_P2_R2099_U132;
  assign new_P2_R2099_U42 = ~new_P2_U2729;
  assign new_P2_R2099_U43 = ~new_P2_U2729 | ~new_P2_R2099_U133;
  assign new_P2_R2099_U44 = ~new_P2_U2728;
  assign new_P2_R2099_U45 = ~new_P2_U2728 | ~new_P2_R2099_U134;
  assign new_P2_R2099_U46 = ~new_P2_U2727;
  assign new_P2_R2099_U47 = ~new_P2_U2727 | ~new_P2_R2099_U135;
  assign new_P2_R2099_U48 = ~new_P2_U2726;
  assign new_P2_R2099_U49 = ~new_P2_U2726 | ~new_P2_R2099_U136;
  assign new_P2_R2099_U50 = ~new_P2_U2725;
  assign new_P2_R2099_U51 = ~new_P2_U2725 | ~new_P2_R2099_U137;
  assign new_P2_R2099_U52 = ~new_P2_U2724;
  assign new_P2_R2099_U53 = ~new_P2_U2724 | ~new_P2_R2099_U138;
  assign new_P2_R2099_U54 = ~new_P2_U2723;
  assign new_P2_R2099_U55 = ~new_P2_U2723 | ~new_P2_R2099_U139;
  assign new_P2_R2099_U56 = ~new_P2_U2722;
  assign new_P2_R2099_U57 = ~new_P2_U2722 | ~new_P2_R2099_U140;
  assign new_P2_R2099_U58 = ~new_P2_U2721;
  assign new_P2_R2099_U59 = ~new_P2_U2721 | ~new_P2_R2099_U141;
  assign new_P2_R2099_U60 = ~new_P2_U2720;
  assign new_P2_R2099_U61 = ~new_P2_U2720 | ~new_P2_R2099_U142;
  assign new_P2_R2099_U62 = ~new_P2_U2719;
  assign new_P2_R2099_U63 = ~new_P2_U2719 | ~new_P2_R2099_U143;
  assign new_P2_R2099_U64 = ~new_P2_U2718;
  assign new_P2_R2099_U65 = ~new_P2_U2718 | ~new_P2_R2099_U144;
  assign new_P2_R2099_U66 = ~new_P2_U2717;
  assign new_P2_R2099_U67 = ~new_P2_R2099_U150 | ~new_P2_R2099_U149;
  assign new_P2_R2099_U68 = ~new_P2_R2099_U152 | ~new_P2_R2099_U151;
  assign new_P2_R2099_U69 = ~new_P2_R2099_U154 | ~new_P2_R2099_U153;
  assign new_P2_R2099_U70 = ~new_P2_R2099_U156 | ~new_P2_R2099_U155;
  assign new_P2_R2099_U71 = ~new_P2_R2099_U158 | ~new_P2_R2099_U157;
  assign new_P2_R2099_U72 = ~new_P2_R2099_U169 | ~new_P2_R2099_U168;
  assign new_P2_R2099_U73 = ~new_P2_R2099_U171 | ~new_P2_R2099_U170;
  assign new_P2_R2099_U74 = ~new_P2_R2099_U180 | ~new_P2_R2099_U179;
  assign new_P2_R2099_U75 = ~new_P2_R2099_U182 | ~new_P2_R2099_U181;
  assign new_P2_R2099_U76 = ~new_P2_R2099_U184 | ~new_P2_R2099_U183;
  assign new_P2_R2099_U77 = ~new_P2_R2099_U186 | ~new_P2_R2099_U185;
  assign new_P2_R2099_U78 = ~new_P2_R2099_U188 | ~new_P2_R2099_U187;
  assign new_P2_R2099_U79 = ~new_P2_R2099_U190 | ~new_P2_R2099_U189;
  assign new_P2_R2099_U80 = ~new_P2_R2099_U192 | ~new_P2_R2099_U191;
  assign new_P2_R2099_U81 = ~new_P2_R2099_U194 | ~new_P2_R2099_U193;
  assign new_P2_R2099_U82 = ~new_P2_R2099_U196 | ~new_P2_R2099_U195;
  assign new_P2_R2099_U83 = ~new_P2_R2099_U198 | ~new_P2_R2099_U197;
  assign new_P2_R2099_U84 = ~new_P2_R2099_U205 | ~new_P2_R2099_U204;
  assign new_P2_R2099_U85 = ~new_P2_R2099_U207 | ~new_P2_R2099_U206;
  assign new_P2_R2099_U86 = ~new_P2_R2099_U209 | ~new_P2_R2099_U208;
  assign new_P2_R2099_U87 = ~new_P2_R2099_U211 | ~new_P2_R2099_U210;
  assign new_P2_R2099_U88 = ~new_P2_R2099_U213 | ~new_P2_R2099_U212;
  assign new_P2_R2099_U89 = ~new_P2_R2099_U215 | ~new_P2_R2099_U214;
  assign new_P2_R2099_U90 = ~new_P2_R2099_U217 | ~new_P2_R2099_U216;
  assign new_P2_R2099_U91 = ~new_P2_R2099_U219 | ~new_P2_R2099_U218;
  assign new_P2_R2099_U92 = ~new_P2_R2099_U221 | ~new_P2_R2099_U220;
  assign new_P2_R2099_U93 = ~new_P2_R2099_U223 | ~new_P2_R2099_U222;
  assign new_P2_R2099_U94 = ~new_P2_R2099_U225 | ~new_P2_R2099_U224;
  assign new_P2_R2099_U95 = ~new_P2_R2099_U167 | ~new_P2_R2099_U166;
  assign new_P2_R2099_U96 = ~new_P2_R2099_U178 | ~new_P2_R2099_U177;
  assign new_P2_R2099_U97 = ~new_P2_R2099_U118 | ~new_P2_R2099_U117;
  assign new_P2_R2099_U98 = new_P2_R2099_U160 & new_P2_R2099_U159;
  assign new_P2_R2099_U99 = new_P2_R2099_U162 & new_P2_R2099_U161;
  assign new_P2_R2099_U100 = ~new_P2_R2099_U114 | ~new_P2_R2099_U113;
  assign new_P2_R2099_U101 = ~new_P2_U2716;
  assign new_P2_R2099_U102 = ~new_P2_U2717 | ~new_P2_R2099_U145;
  assign new_P2_R2099_U103 = new_P2_R2099_U173 & new_P2_R2099_U172;
  assign new_P2_R2099_U104 = ~new_P2_R2099_U106 | ~new_P2_R2099_U110;
  assign new_P2_R2099_U105 = ~new_P2_U2751 | ~new_P2_U2747;
  assign new_P2_R2099_U106 = ~new_P2_U2751 | ~new_P2_U2746 | ~new_P2_U2747;
  assign new_P2_R2099_U107 = new_P2_R2099_U203 & new_P2_R2099_U202;
  assign new_P2_R2099_U108 = ~new_P2_R2099_U106;
  assign new_P2_R2099_U109 = ~new_P2_R2099_U9 | ~new_P2_R2099_U105;
  assign new_P2_R2099_U110 = ~new_P2_U2750 | ~new_P2_R2099_U109;
  assign new_P2_R2099_U111 = ~new_P2_R2099_U104;
  assign new_P2_R2099_U112 = new_P2_U2749 | new_P2_U2745;
  assign new_P2_R2099_U113 = ~new_P2_R2099_U112 | ~new_P2_R2099_U104;
  assign new_P2_R2099_U114 = ~new_P2_U2745 | ~new_P2_U2749;
  assign new_P2_R2099_U115 = ~new_P2_R2099_U100;
  assign new_P2_R2099_U116 = new_P2_U2748 | new_P2_U2744;
  assign new_P2_R2099_U117 = ~new_P2_R2099_U116 | ~new_P2_R2099_U100;
  assign new_P2_R2099_U118 = ~new_P2_U2744 | ~new_P2_U2748;
  assign new_P2_R2099_U119 = ~new_P2_R2099_U97;
  assign new_P2_R2099_U120 = ~new_P2_R2099_U15;
  assign new_P2_R2099_U121 = ~new_P2_R2099_U17;
  assign new_P2_R2099_U122 = ~new_P2_R2099_U19;
  assign new_P2_R2099_U123 = ~new_P2_R2099_U21;
  assign new_P2_R2099_U124 = ~new_P2_R2099_U24;
  assign new_P2_R2099_U125 = ~new_P2_R2099_U25;
  assign new_P2_R2099_U126 = ~new_P2_R2099_U27;
  assign new_P2_R2099_U127 = ~new_P2_R2099_U29;
  assign new_P2_R2099_U128 = ~new_P2_R2099_U31;
  assign new_P2_R2099_U129 = ~new_P2_R2099_U33;
  assign new_P2_R2099_U130 = ~new_P2_R2099_U35;
  assign new_P2_R2099_U131 = ~new_P2_R2099_U37;
  assign new_P2_R2099_U132 = ~new_P2_R2099_U39;
  assign new_P2_R2099_U133 = ~new_P2_R2099_U41;
  assign new_P2_R2099_U134 = ~new_P2_R2099_U43;
  assign new_P2_R2099_U135 = ~new_P2_R2099_U45;
  assign new_P2_R2099_U136 = ~new_P2_R2099_U47;
  assign new_P2_R2099_U137 = ~new_P2_R2099_U49;
  assign new_P2_R2099_U138 = ~new_P2_R2099_U51;
  assign new_P2_R2099_U139 = ~new_P2_R2099_U53;
  assign new_P2_R2099_U140 = ~new_P2_R2099_U55;
  assign new_P2_R2099_U141 = ~new_P2_R2099_U57;
  assign new_P2_R2099_U142 = ~new_P2_R2099_U59;
  assign new_P2_R2099_U143 = ~new_P2_R2099_U61;
  assign new_P2_R2099_U144 = ~new_P2_R2099_U63;
  assign new_P2_R2099_U145 = ~new_P2_R2099_U65;
  assign new_P2_R2099_U146 = ~new_P2_R2099_U102;
  assign new_P2_R2099_U147 = ~new_P2_R2099_U105;
  assign new_P2_R2099_U148 = ~new_P2_R2099_U201 | ~new_P2_R2099_U9;
  assign new_P2_R2099_U149 = ~new_P2_U2738 | ~new_P2_R2099_U24;
  assign new_P2_R2099_U150 = ~new_P2_R2099_U124 | ~new_P2_R2099_U23;
  assign new_P2_R2099_U151 = ~new_P2_U2739 | ~new_P2_R2099_U21;
  assign new_P2_R2099_U152 = ~new_P2_R2099_U123 | ~new_P2_R2099_U22;
  assign new_P2_R2099_U153 = ~new_P2_U2740 | ~new_P2_R2099_U19;
  assign new_P2_R2099_U154 = ~new_P2_R2099_U122 | ~new_P2_R2099_U20;
  assign new_P2_R2099_U155 = ~new_P2_U2741 | ~new_P2_R2099_U17;
  assign new_P2_R2099_U156 = ~new_P2_R2099_U121 | ~new_P2_R2099_U18;
  assign new_P2_R2099_U157 = ~new_P2_U2742 | ~new_P2_R2099_U15;
  assign new_P2_R2099_U158 = ~new_P2_R2099_U120 | ~new_P2_R2099_U16;
  assign new_P2_R2099_U159 = ~new_P2_U2743 | ~new_P2_R2099_U97;
  assign new_P2_R2099_U160 = ~new_P2_R2099_U119 | ~new_P2_R2099_U14;
  assign new_P2_R2099_U161 = ~new_P2_U2744 | ~new_P2_R2099_U12;
  assign new_P2_R2099_U162 = ~new_P2_U2748 | ~new_P2_R2099_U13;
  assign new_P2_R2099_U163 = ~new_P2_U2744 | ~new_P2_R2099_U12;
  assign new_P2_R2099_U164 = ~new_P2_U2748 | ~new_P2_R2099_U13;
  assign new_P2_R2099_U165 = ~new_P2_R2099_U164 | ~new_P2_R2099_U163;
  assign new_P2_R2099_U166 = ~new_P2_R2099_U99 | ~new_P2_R2099_U100;
  assign new_P2_R2099_U167 = ~new_P2_R2099_U115 | ~new_P2_R2099_U165;
  assign new_P2_R2099_U168 = ~new_P2_U2716 | ~new_P2_R2099_U102;
  assign new_P2_R2099_U169 = ~new_P2_R2099_U146 | ~new_P2_R2099_U101;
  assign new_P2_R2099_U170 = ~new_P2_U2717 | ~new_P2_R2099_U65;
  assign new_P2_R2099_U171 = ~new_P2_R2099_U145 | ~new_P2_R2099_U66;
  assign new_P2_R2099_U172 = ~new_P2_U2745 | ~new_P2_R2099_U10;
  assign new_P2_R2099_U173 = ~new_P2_U2749 | ~new_P2_R2099_U11;
  assign new_P2_R2099_U174 = ~new_P2_U2745 | ~new_P2_R2099_U10;
  assign new_P2_R2099_U175 = ~new_P2_U2749 | ~new_P2_R2099_U11;
  assign new_P2_R2099_U176 = ~new_P2_R2099_U175 | ~new_P2_R2099_U174;
  assign new_P2_R2099_U177 = ~new_P2_R2099_U103 | ~new_P2_R2099_U104;
  assign new_P2_R2099_U178 = ~new_P2_R2099_U111 | ~new_P2_R2099_U176;
  assign new_P2_R2099_U179 = ~new_P2_U2718 | ~new_P2_R2099_U63;
  assign new_P2_R2099_U180 = ~new_P2_R2099_U144 | ~new_P2_R2099_U64;
  assign new_P2_R2099_U181 = ~new_P2_U2719 | ~new_P2_R2099_U61;
  assign new_P2_R2099_U182 = ~new_P2_R2099_U143 | ~new_P2_R2099_U62;
  assign new_P2_R2099_U183 = ~new_P2_U2720 | ~new_P2_R2099_U59;
  assign new_P2_R2099_U184 = ~new_P2_R2099_U142 | ~new_P2_R2099_U60;
  assign new_P2_R2099_U185 = ~new_P2_U2721 | ~new_P2_R2099_U57;
  assign new_P2_R2099_U186 = ~new_P2_R2099_U141 | ~new_P2_R2099_U58;
  assign new_P2_R2099_U187 = ~new_P2_U2722 | ~new_P2_R2099_U55;
  assign new_P2_R2099_U188 = ~new_P2_R2099_U140 | ~new_P2_R2099_U56;
  assign new_P2_R2099_U189 = ~new_P2_U2723 | ~new_P2_R2099_U53;
  assign new_P2_R2099_U190 = ~new_P2_R2099_U139 | ~new_P2_R2099_U54;
  assign new_P2_R2099_U191 = ~new_P2_U2724 | ~new_P2_R2099_U51;
  assign new_P2_R2099_U192 = ~new_P2_R2099_U138 | ~new_P2_R2099_U52;
  assign new_P2_R2099_U193 = ~new_P2_U2725 | ~new_P2_R2099_U49;
  assign new_P2_R2099_U194 = ~new_P2_R2099_U137 | ~new_P2_R2099_U50;
  assign new_P2_R2099_U195 = ~new_P2_U2726 | ~new_P2_R2099_U47;
  assign new_P2_R2099_U196 = ~new_P2_R2099_U136 | ~new_P2_R2099_U48;
  assign new_P2_R2099_U197 = ~new_P2_U2727 | ~new_P2_R2099_U45;
  assign new_P2_R2099_U198 = ~new_P2_R2099_U135 | ~new_P2_R2099_U46;
  assign new_P2_R2099_U199 = ~new_P2_U2750 | ~new_P2_R2099_U105;
  assign new_P2_R2099_U200 = ~new_P2_R2099_U147 | ~new_P2_R2099_U8;
  assign new_P2_R2099_U201 = ~new_P2_R2099_U200 | ~new_P2_R2099_U199;
  assign new_P2_R2099_U202 = ~new_P2_R2099_U8 | ~new_P2_U2746 | ~new_P2_R2099_U105;
  assign new_P2_R2099_U203 = ~new_P2_R2099_U108 | ~new_P2_U2750;
  assign new_P2_R2099_U204 = ~new_P2_U2728 | ~new_P2_R2099_U43;
  assign new_P2_R2099_U205 = ~new_P2_R2099_U134 | ~new_P2_R2099_U44;
  assign new_P2_R2099_U206 = ~new_P2_U2729 | ~new_P2_R2099_U41;
  assign new_P2_R2099_U207 = ~new_P2_R2099_U133 | ~new_P2_R2099_U42;
  assign new_P2_R2099_U208 = ~new_P2_U2730 | ~new_P2_R2099_U39;
  assign new_P2_R2099_U209 = ~new_P2_R2099_U132 | ~new_P2_R2099_U40;
  assign new_P2_R2099_U210 = ~new_P2_U2731 | ~new_P2_R2099_U37;
  assign new_P2_R2099_U211 = ~new_P2_R2099_U131 | ~new_P2_R2099_U38;
  assign new_P2_R2099_U212 = ~new_P2_U2732 | ~new_P2_R2099_U35;
  assign new_P2_R2099_U213 = ~new_P2_R2099_U130 | ~new_P2_R2099_U36;
  assign new_P2_R2099_U214 = ~new_P2_U2733 | ~new_P2_R2099_U33;
  assign new_P2_R2099_U215 = ~new_P2_R2099_U129 | ~new_P2_R2099_U34;
  assign new_P2_R2099_U216 = ~new_P2_U2734 | ~new_P2_R2099_U31;
  assign new_P2_R2099_U217 = ~new_P2_R2099_U128 | ~new_P2_R2099_U32;
  assign new_P2_R2099_U218 = ~new_P2_U2735 | ~new_P2_R2099_U29;
  assign new_P2_R2099_U219 = ~new_P2_R2099_U127 | ~new_P2_R2099_U30;
  assign new_P2_R2099_U220 = ~new_P2_U2736 | ~new_P2_R2099_U27;
  assign new_P2_R2099_U221 = ~new_P2_R2099_U126 | ~new_P2_R2099_U28;
  assign new_P2_R2099_U222 = ~new_P2_U2737 | ~new_P2_R2099_U25;
  assign new_P2_R2099_U223 = ~new_P2_R2099_U125 | ~new_P2_R2099_U26;
  assign new_P2_R2099_U224 = ~new_P2_U2751 | ~new_P2_R2099_U6;
  assign new_P2_R2099_U225 = ~new_P2_U2747 | ~new_P2_R2099_U7;
  assign new_P2_ADD_391_1196_U5 = new_P2_ADD_391_1196_U301 & new_P2_ADD_391_1196_U299;
  assign new_P2_ADD_391_1196_U6 = new_P2_ADD_391_1196_U296 & new_P2_ADD_391_1196_U294;
  assign new_P2_ADD_391_1196_U7 = new_P2_ADD_391_1196_U292 & new_P2_ADD_391_1196_U290;
  assign new_P2_ADD_391_1196_U8 = new_P2_ADD_391_1196_U287 & new_P2_ADD_391_1196_U283;
  assign new_P2_ADD_391_1196_U9 = new_P2_ADD_391_1196_U205 & new_P2_ADD_391_1196_U203;
  assign new_P2_ADD_391_1196_U10 = new_P2_ADD_391_1196_U201 & new_P2_ADD_391_1196_U199;
  assign new_P2_ADD_391_1196_U11 = new_P2_ADD_391_1196_U196 & new_P2_ADD_391_1196_U192;
  assign new_P2_ADD_391_1196_U12 = ~new_P2_ADD_391_1196_U144 | ~new_P2_ADD_391_1196_U306;
  assign new_P2_ADD_391_1196_U13 = ~new_P2_R2182_U72;
  assign new_P2_ADD_391_1196_U14 = ~new_P2_R2096_U71;
  assign new_P2_ADD_391_1196_U15 = ~new_P2_R2182_U73;
  assign new_P2_ADD_391_1196_U16 = ~new_P2_R2096_U72;
  assign new_P2_ADD_391_1196_U17 = ~new_P2_R2182_U74;
  assign new_P2_ADD_391_1196_U18 = ~new_P2_R2096_U73;
  assign new_P2_ADD_391_1196_U19 = ~new_P2_R2096_U68;
  assign new_P2_ADD_391_1196_U20 = ~new_P2_R2182_U69;
  assign new_P2_ADD_391_1196_U21 = ~new_P2_R2182_U68;
  assign new_P2_ADD_391_1196_U22 = ~new_P2_R2182_U69 | ~new_P2_R2096_U68;
  assign new_P2_ADD_391_1196_U23 = ~new_P2_R2096_U51;
  assign new_P2_ADD_391_1196_U24 = ~new_P2_R2182_U40;
  assign new_P2_ADD_391_1196_U25 = ~new_P2_R2096_U77;
  assign new_P2_ADD_391_1196_U26 = ~new_P2_R2182_U76;
  assign new_P2_ADD_391_1196_U27 = ~new_P2_R2096_U75;
  assign new_P2_ADD_391_1196_U28 = ~new_P2_R2182_U75;
  assign new_P2_ADD_391_1196_U29 = ~new_P2_R2096_U74;
  assign new_P2_ADD_391_1196_U30 = ~new_P2_ADD_391_1196_U39 | ~new_P2_ADD_391_1196_U180;
  assign new_P2_ADD_391_1196_U31 = ~new_P2_R2182_U71;
  assign new_P2_ADD_391_1196_U32 = ~new_P2_R2096_U70;
  assign new_P2_ADD_391_1196_U33 = ~new_P2_R2096_U69;
  assign new_P2_ADD_391_1196_U34 = ~new_P2_R2182_U70;
  assign new_P2_ADD_391_1196_U35 = ~new_P2_ADD_391_1196_U190 | ~new_P2_ADD_391_1196_U189;
  assign new_P2_ADD_391_1196_U36 = ~new_P2_ADD_391_1196_U35 | ~new_P2_ADD_391_1196_U193;
  assign new_P2_ADD_391_1196_U37 = ~new_P2_ADD_391_1196_U183 | ~new_P2_ADD_391_1196_U184 | ~new_P2_ADD_391_1196_U182;
  assign new_P2_ADD_391_1196_U38 = ~new_P2_ADD_391_1196_U176 | ~new_P2_ADD_391_1196_U175;
  assign new_P2_ADD_391_1196_U39 = ~new_P2_ADD_391_1196_U38 | ~new_P2_ADD_391_1196_U178;
  assign new_P2_ADD_391_1196_U40 = ~new_P2_R2182_U91;
  assign new_P2_ADD_391_1196_U41 = ~new_P2_R2096_U92;
  assign new_P2_ADD_391_1196_U42 = ~new_P2_R2182_U92;
  assign new_P2_ADD_391_1196_U43 = ~new_P2_R2096_U93;
  assign new_P2_ADD_391_1196_U44 = ~new_P2_R2182_U93;
  assign new_P2_ADD_391_1196_U45 = ~new_P2_R2096_U94;
  assign new_P2_ADD_391_1196_U46 = ~new_P2_R2182_U95;
  assign new_P2_ADD_391_1196_U47 = ~new_P2_R2096_U96;
  assign new_P2_ADD_391_1196_U48 = ~new_P2_R2182_U96;
  assign new_P2_ADD_391_1196_U49 = ~new_P2_R2096_U97;
  assign new_P2_ADD_391_1196_U50 = ~new_P2_ADD_391_1196_U36 | ~new_P2_ADD_391_1196_U206;
  assign new_P2_ADD_391_1196_U51 = ~new_P2_R2182_U94;
  assign new_P2_ADD_391_1196_U52 = ~new_P2_R2096_U95;
  assign new_P2_ADD_391_1196_U53 = ~new_P2_ADD_391_1196_U85 | ~new_P2_ADD_391_1196_U220;
  assign new_P2_ADD_391_1196_U54 = ~new_P2_R2182_U90;
  assign new_P2_ADD_391_1196_U55 = ~new_P2_R2096_U91;
  assign new_P2_ADD_391_1196_U56 = ~new_P2_R2182_U89;
  assign new_P2_ADD_391_1196_U57 = ~new_P2_R2096_U90;
  assign new_P2_ADD_391_1196_U58 = ~new_P2_R2182_U88;
  assign new_P2_ADD_391_1196_U59 = ~new_P2_R2096_U89;
  assign new_P2_ADD_391_1196_U60 = ~new_P2_R2182_U87;
  assign new_P2_ADD_391_1196_U61 = ~new_P2_R2096_U88;
  assign new_P2_ADD_391_1196_U62 = ~new_P2_R2182_U86;
  assign new_P2_ADD_391_1196_U63 = ~new_P2_R2096_U87;
  assign new_P2_ADD_391_1196_U64 = ~new_P2_R2182_U85;
  assign new_P2_ADD_391_1196_U65 = ~new_P2_R2096_U86;
  assign new_P2_ADD_391_1196_U66 = ~new_P2_R2182_U84;
  assign new_P2_ADD_391_1196_U67 = ~new_P2_R2096_U85;
  assign new_P2_ADD_391_1196_U68 = ~new_P2_R2182_U83;
  assign new_P2_ADD_391_1196_U69 = ~new_P2_R2096_U84;
  assign new_P2_ADD_391_1196_U70 = ~new_P2_R2182_U82;
  assign new_P2_ADD_391_1196_U71 = ~new_P2_R2096_U83;
  assign new_P2_ADD_391_1196_U72 = ~new_P2_R2182_U81;
  assign new_P2_ADD_391_1196_U73 = ~new_P2_R2096_U82;
  assign new_P2_ADD_391_1196_U74 = ~new_P2_R2182_U80;
  assign new_P2_ADD_391_1196_U75 = ~new_P2_R2096_U81;
  assign new_P2_ADD_391_1196_U76 = ~new_P2_R2182_U79;
  assign new_P2_ADD_391_1196_U77 = ~new_P2_R2096_U80;
  assign new_P2_ADD_391_1196_U78 = ~new_P2_R2096_U79;
  assign new_P2_ADD_391_1196_U79 = ~new_P2_R2182_U78;
  assign new_P2_ADD_391_1196_U80 = ~new_P2_R2096_U78;
  assign new_P2_ADD_391_1196_U81 = ~new_P2_R2182_U77;
  assign new_P2_ADD_391_1196_U82 = ~new_P2_ADD_391_1196_U278 | ~new_P2_ADD_391_1196_U277;
  assign new_P2_ADD_391_1196_U83 = ~new_P2_ADD_391_1196_U223 | ~new_P2_ADD_391_1196_U224 | ~new_P2_ADD_391_1196_U222;
  assign new_P2_ADD_391_1196_U84 = ~new_P2_ADD_391_1196_U216 | ~new_P2_ADD_391_1196_U215;
  assign new_P2_ADD_391_1196_U85 = ~new_P2_ADD_391_1196_U84 | ~new_P2_ADD_391_1196_U218;
  assign new_P2_ADD_391_1196_U86 = ~new_P2_ADD_391_1196_U209 | ~new_P2_ADD_391_1196_U210 | ~new_P2_ADD_391_1196_U208;
  assign new_P2_ADD_391_1196_U87 = ~new_P2_ADD_391_1196_U478 | ~new_P2_ADD_391_1196_U477;
  assign new_P2_ADD_391_1196_U88 = ~new_P2_ADD_391_1196_U315 | ~new_P2_ADD_391_1196_U314;
  assign new_P2_ADD_391_1196_U89 = ~new_P2_ADD_391_1196_U322 | ~new_P2_ADD_391_1196_U321;
  assign new_P2_ADD_391_1196_U90 = ~new_P2_ADD_391_1196_U331 | ~new_P2_ADD_391_1196_U330;
  assign new_P2_ADD_391_1196_U91 = ~new_P2_ADD_391_1196_U338 | ~new_P2_ADD_391_1196_U337;
  assign new_P2_ADD_391_1196_U92 = ~new_P2_ADD_391_1196_U350 | ~new_P2_ADD_391_1196_U349;
  assign new_P2_ADD_391_1196_U93 = ~new_P2_ADD_391_1196_U357 | ~new_P2_ADD_391_1196_U356;
  assign new_P2_ADD_391_1196_U94 = ~new_P2_ADD_391_1196_U364 | ~new_P2_ADD_391_1196_U363;
  assign new_P2_ADD_391_1196_U95 = ~new_P2_ADD_391_1196_U371 | ~new_P2_ADD_391_1196_U370;
  assign new_P2_ADD_391_1196_U96 = ~new_P2_ADD_391_1196_U378 | ~new_P2_ADD_391_1196_U377;
  assign new_P2_ADD_391_1196_U97 = ~new_P2_ADD_391_1196_U385 | ~new_P2_ADD_391_1196_U384;
  assign new_P2_ADD_391_1196_U98 = ~new_P2_ADD_391_1196_U392 | ~new_P2_ADD_391_1196_U391;
  assign new_P2_ADD_391_1196_U99 = ~new_P2_ADD_391_1196_U399 | ~new_P2_ADD_391_1196_U398;
  assign new_P2_ADD_391_1196_U100 = ~new_P2_ADD_391_1196_U406 | ~new_P2_ADD_391_1196_U405;
  assign new_P2_ADD_391_1196_U101 = ~new_P2_ADD_391_1196_U413 | ~new_P2_ADD_391_1196_U412;
  assign new_P2_ADD_391_1196_U102 = ~new_P2_ADD_391_1196_U420 | ~new_P2_ADD_391_1196_U419;
  assign new_P2_ADD_391_1196_U103 = ~new_P2_ADD_391_1196_U432 | ~new_P2_ADD_391_1196_U431;
  assign new_P2_ADD_391_1196_U104 = ~new_P2_ADD_391_1196_U439 | ~new_P2_ADD_391_1196_U438;
  assign new_P2_ADD_391_1196_U105 = ~new_P2_ADD_391_1196_U446 | ~new_P2_ADD_391_1196_U445;
  assign new_P2_ADD_391_1196_U106 = ~new_P2_ADD_391_1196_U453 | ~new_P2_ADD_391_1196_U452;
  assign new_P2_ADD_391_1196_U107 = ~new_P2_ADD_391_1196_U460 | ~new_P2_ADD_391_1196_U459;
  assign new_P2_ADD_391_1196_U108 = ~new_P2_ADD_391_1196_U469 | ~new_P2_ADD_391_1196_U468;
  assign new_P2_ADD_391_1196_U109 = ~new_P2_ADD_391_1196_U476 | ~new_P2_ADD_391_1196_U475;
  assign new_P2_ADD_391_1196_U110 = new_P2_ADD_391_1196_U308 & new_P2_ADD_391_1196_U307;
  assign new_P2_ADD_391_1196_U111 = new_P2_ADD_391_1196_U310 & new_P2_ADD_391_1196_U309;
  assign new_P2_ADD_391_1196_U112 = ~new_P2_ADD_391_1196_U37 | ~new_P2_ADD_391_1196_U186;
  assign new_P2_ADD_391_1196_U113 = new_P2_ADD_391_1196_U317 & new_P2_ADD_391_1196_U316;
  assign new_P2_ADD_391_1196_U114 = new_P2_ADD_391_1196_U324 & new_P2_ADD_391_1196_U323;
  assign new_P2_ADD_391_1196_U115 = new_P2_ADD_391_1196_U326 & new_P2_ADD_391_1196_U325;
  assign new_P2_ADD_391_1196_U116 = ~new_P2_ADD_391_1196_U172 | ~new_P2_ADD_391_1196_U171;
  assign new_P2_ADD_391_1196_U117 = new_P2_ADD_391_1196_U333 & new_P2_ADD_391_1196_U332;
  assign new_P2_ADD_391_1196_U118 = ~new_P2_ADD_391_1196_U168 | ~new_P2_ADD_391_1196_U167;
  assign new_P2_ADD_391_1196_U119 = ~new_P2_R2182_U41;
  assign new_P2_ADD_391_1196_U120 = ~new_P2_R2096_U76;
  assign new_P2_ADD_391_1196_U121 = new_P2_ADD_391_1196_U340 & new_P2_ADD_391_1196_U339;
  assign new_P2_ADD_391_1196_U122 = new_P2_ADD_391_1196_U345 & new_P2_ADD_391_1196_U344;
  assign new_P2_ADD_391_1196_U123 = ~new_P2_ADD_391_1196_U143 | ~new_P2_ADD_391_1196_U164;
  assign new_P2_ADD_391_1196_U124 = new_P2_ADD_391_1196_U352 & new_P2_ADD_391_1196_U351;
  assign new_P2_ADD_391_1196_U125 = new_P2_ADD_391_1196_U359 & new_P2_ADD_391_1196_U358;
  assign new_P2_ADD_391_1196_U126 = ~new_P2_ADD_391_1196_U274 | ~new_P2_ADD_391_1196_U273;
  assign new_P2_ADD_391_1196_U127 = new_P2_ADD_391_1196_U366 & new_P2_ADD_391_1196_U365;
  assign new_P2_ADD_391_1196_U128 = ~new_P2_ADD_391_1196_U270 | ~new_P2_ADD_391_1196_U269;
  assign new_P2_ADD_391_1196_U129 = new_P2_ADD_391_1196_U373 & new_P2_ADD_391_1196_U372;
  assign new_P2_ADD_391_1196_U130 = ~new_P2_ADD_391_1196_U266 | ~new_P2_ADD_391_1196_U265;
  assign new_P2_ADD_391_1196_U131 = new_P2_ADD_391_1196_U380 & new_P2_ADD_391_1196_U379;
  assign new_P2_ADD_391_1196_U132 = ~new_P2_ADD_391_1196_U262 | ~new_P2_ADD_391_1196_U261;
  assign new_P2_ADD_391_1196_U133 = new_P2_ADD_391_1196_U387 & new_P2_ADD_391_1196_U386;
  assign new_P2_ADD_391_1196_U134 = ~new_P2_ADD_391_1196_U258 | ~new_P2_ADD_391_1196_U257;
  assign new_P2_ADD_391_1196_U135 = new_P2_ADD_391_1196_U394 & new_P2_ADD_391_1196_U393;
  assign new_P2_ADD_391_1196_U136 = ~new_P2_ADD_391_1196_U254 | ~new_P2_ADD_391_1196_U253;
  assign new_P2_ADD_391_1196_U137 = new_P2_ADD_391_1196_U401 & new_P2_ADD_391_1196_U400;
  assign new_P2_ADD_391_1196_U138 = ~new_P2_ADD_391_1196_U250 | ~new_P2_ADD_391_1196_U249;
  assign new_P2_ADD_391_1196_U139 = new_P2_ADD_391_1196_U408 & new_P2_ADD_391_1196_U407;
  assign new_P2_ADD_391_1196_U140 = ~new_P2_ADD_391_1196_U246 | ~new_P2_ADD_391_1196_U245;
  assign new_P2_ADD_391_1196_U141 = new_P2_ADD_391_1196_U415 & new_P2_ADD_391_1196_U414;
  assign new_P2_ADD_391_1196_U142 = ~new_P2_ADD_391_1196_U242 | ~new_P2_ADD_391_1196_U241;
  assign new_P2_ADD_391_1196_U143 = ~new_P2_R2096_U51 | ~new_P2_ADD_391_1196_U162;
  assign new_P2_ADD_391_1196_U144 = new_P2_ADD_391_1196_U425 & new_P2_ADD_391_1196_U424;
  assign new_P2_ADD_391_1196_U145 = new_P2_ADD_391_1196_U427 & new_P2_ADD_391_1196_U426;
  assign new_P2_ADD_391_1196_U146 = ~new_P2_ADD_391_1196_U238 | ~new_P2_ADD_391_1196_U237;
  assign new_P2_ADD_391_1196_U147 = new_P2_ADD_391_1196_U434 & new_P2_ADD_391_1196_U433;
  assign new_P2_ADD_391_1196_U148 = ~new_P2_ADD_391_1196_U234 | ~new_P2_ADD_391_1196_U233;
  assign new_P2_ADD_391_1196_U149 = new_P2_ADD_391_1196_U441 & new_P2_ADD_391_1196_U440;
  assign new_P2_ADD_391_1196_U150 = ~new_P2_ADD_391_1196_U230 | ~new_P2_ADD_391_1196_U229;
  assign new_P2_ADD_391_1196_U151 = new_P2_ADD_391_1196_U448 & new_P2_ADD_391_1196_U447;
  assign new_P2_ADD_391_1196_U152 = ~new_P2_ADD_391_1196_U83 | ~new_P2_ADD_391_1196_U226;
  assign new_P2_ADD_391_1196_U153 = new_P2_ADD_391_1196_U455 & new_P2_ADD_391_1196_U454;
  assign new_P2_ADD_391_1196_U154 = new_P2_ADD_391_1196_U462 & new_P2_ADD_391_1196_U461;
  assign new_P2_ADD_391_1196_U155 = new_P2_ADD_391_1196_U464 & new_P2_ADD_391_1196_U463;
  assign new_P2_ADD_391_1196_U156 = ~new_P2_ADD_391_1196_U86 | ~new_P2_ADD_391_1196_U212;
  assign new_P2_ADD_391_1196_U157 = new_P2_ADD_391_1196_U471 & new_P2_ADD_391_1196_U470;
  assign new_P2_ADD_391_1196_U158 = ~new_P2_R2096_U97 | ~new_P2_R2182_U96;
  assign new_P2_ADD_391_1196_U159 = ~new_P2_R2096_U93 | ~new_P2_R2182_U92;
  assign new_P2_ADD_391_1196_U160 = ~new_P2_ADD_391_1196_U143;
  assign new_P2_ADD_391_1196_U161 = ~new_P2_R2096_U72 | ~new_P2_R2182_U73;
  assign new_P2_ADD_391_1196_U162 = ~new_P2_ADD_391_1196_U22;
  assign new_P2_ADD_391_1196_U163 = ~new_P2_ADD_391_1196_U23 | ~new_P2_ADD_391_1196_U22;
  assign new_P2_ADD_391_1196_U164 = ~new_P2_R2182_U68 | ~new_P2_ADD_391_1196_U163;
  assign new_P2_ADD_391_1196_U165 = ~new_P2_ADD_391_1196_U123;
  assign new_P2_ADD_391_1196_U166 = new_P2_R2182_U40 | new_P2_R2096_U77;
  assign new_P2_ADD_391_1196_U167 = ~new_P2_ADD_391_1196_U166 | ~new_P2_ADD_391_1196_U123;
  assign new_P2_ADD_391_1196_U168 = ~new_P2_R2096_U77 | ~new_P2_R2182_U40;
  assign new_P2_ADD_391_1196_U169 = ~new_P2_ADD_391_1196_U118;
  assign new_P2_ADD_391_1196_U170 = new_P2_R2182_U76 | new_P2_R2096_U75;
  assign new_P2_ADD_391_1196_U171 = ~new_P2_ADD_391_1196_U170 | ~new_P2_ADD_391_1196_U118;
  assign new_P2_ADD_391_1196_U172 = ~new_P2_R2096_U75 | ~new_P2_R2182_U76;
  assign new_P2_ADD_391_1196_U173 = ~new_P2_ADD_391_1196_U116;
  assign new_P2_ADD_391_1196_U174 = new_P2_R2182_U75 | new_P2_R2096_U74;
  assign new_P2_ADD_391_1196_U175 = ~new_P2_ADD_391_1196_U174 | ~new_P2_ADD_391_1196_U116;
  assign new_P2_ADD_391_1196_U176 = ~new_P2_R2096_U74 | ~new_P2_R2182_U75;
  assign new_P2_ADD_391_1196_U177 = ~new_P2_ADD_391_1196_U38;
  assign new_P2_ADD_391_1196_U178 = new_P2_R2096_U73 | new_P2_R2182_U74;
  assign new_P2_ADD_391_1196_U179 = ~new_P2_ADD_391_1196_U39;
  assign new_P2_ADD_391_1196_U180 = ~new_P2_R2096_U73 | ~new_P2_R2182_U74;
  assign new_P2_ADD_391_1196_U181 = ~new_P2_ADD_391_1196_U30;
  assign new_P2_ADD_391_1196_U182 = ~new_P2_ADD_391_1196_U181 | ~new_P2_ADD_391_1196_U161;
  assign new_P2_ADD_391_1196_U183 = new_P2_R2096_U71 | new_P2_R2182_U72;
  assign new_P2_ADD_391_1196_U184 = new_P2_R2096_U72 | new_P2_R2182_U73;
  assign new_P2_ADD_391_1196_U185 = ~new_P2_ADD_391_1196_U37;
  assign new_P2_ADD_391_1196_U186 = ~new_P2_R2096_U71 | ~new_P2_R2182_U72;
  assign new_P2_ADD_391_1196_U187 = ~new_P2_ADD_391_1196_U112;
  assign new_P2_ADD_391_1196_U188 = new_P2_R2182_U71 | new_P2_R2096_U70;
  assign new_P2_ADD_391_1196_U189 = ~new_P2_ADD_391_1196_U188 | ~new_P2_ADD_391_1196_U112;
  assign new_P2_ADD_391_1196_U190 = ~new_P2_R2096_U70 | ~new_P2_R2182_U71;
  assign new_P2_ADD_391_1196_U191 = ~new_P2_ADD_391_1196_U35;
  assign new_P2_ADD_391_1196_U192 = ~new_P2_ADD_391_1196_U110 | ~new_P2_ADD_391_1196_U191;
  assign new_P2_ADD_391_1196_U193 = new_P2_R2096_U69 | new_P2_R2182_U70;
  assign new_P2_ADD_391_1196_U194 = ~new_P2_ADD_391_1196_U36;
  assign new_P2_ADD_391_1196_U195 = ~new_P2_R2182_U70 | ~new_P2_R2096_U69;
  assign new_P2_ADD_391_1196_U196 = ~new_P2_ADD_391_1196_U194 | ~new_P2_ADD_391_1196_U195;
  assign new_P2_ADD_391_1196_U197 = new_P2_R2182_U73 | new_P2_R2096_U72;
  assign new_P2_ADD_391_1196_U198 = ~new_P2_ADD_391_1196_U197 | ~new_P2_ADD_391_1196_U30;
  assign new_P2_ADD_391_1196_U199 = ~new_P2_ADD_391_1196_U113 | ~new_P2_ADD_391_1196_U198 | ~new_P2_ADD_391_1196_U161;
  assign new_P2_ADD_391_1196_U200 = ~new_P2_R2096_U71 | ~new_P2_R2182_U72;
  assign new_P2_ADD_391_1196_U201 = ~new_P2_ADD_391_1196_U185 | ~new_P2_ADD_391_1196_U200;
  assign new_P2_ADD_391_1196_U202 = new_P2_R2096_U72 | new_P2_R2182_U73;
  assign new_P2_ADD_391_1196_U203 = ~new_P2_ADD_391_1196_U114 | ~new_P2_ADD_391_1196_U177;
  assign new_P2_ADD_391_1196_U204 = ~new_P2_R2096_U73 | ~new_P2_R2182_U74;
  assign new_P2_ADD_391_1196_U205 = ~new_P2_ADD_391_1196_U179 | ~new_P2_ADD_391_1196_U204;
  assign new_P2_ADD_391_1196_U206 = ~new_P2_R2182_U70 | ~new_P2_R2096_U69;
  assign new_P2_ADD_391_1196_U207 = ~new_P2_ADD_391_1196_U50;
  assign new_P2_ADD_391_1196_U208 = ~new_P2_ADD_391_1196_U207 | ~new_P2_ADD_391_1196_U158;
  assign new_P2_ADD_391_1196_U209 = new_P2_R2096_U96 | new_P2_R2182_U95;
  assign new_P2_ADD_391_1196_U210 = new_P2_R2096_U97 | new_P2_R2182_U96;
  assign new_P2_ADD_391_1196_U211 = ~new_P2_ADD_391_1196_U86;
  assign new_P2_ADD_391_1196_U212 = ~new_P2_R2096_U96 | ~new_P2_R2182_U95;
  assign new_P2_ADD_391_1196_U213 = ~new_P2_ADD_391_1196_U156;
  assign new_P2_ADD_391_1196_U214 = new_P2_R2182_U94 | new_P2_R2096_U95;
  assign new_P2_ADD_391_1196_U215 = ~new_P2_ADD_391_1196_U214 | ~new_P2_ADD_391_1196_U156;
  assign new_P2_ADD_391_1196_U216 = ~new_P2_R2096_U95 | ~new_P2_R2182_U94;
  assign new_P2_ADD_391_1196_U217 = ~new_P2_ADD_391_1196_U84;
  assign new_P2_ADD_391_1196_U218 = new_P2_R2096_U94 | new_P2_R2182_U93;
  assign new_P2_ADD_391_1196_U219 = ~new_P2_ADD_391_1196_U85;
  assign new_P2_ADD_391_1196_U220 = ~new_P2_R2096_U94 | ~new_P2_R2182_U93;
  assign new_P2_ADD_391_1196_U221 = ~new_P2_ADD_391_1196_U53;
  assign new_P2_ADD_391_1196_U222 = ~new_P2_ADD_391_1196_U221 | ~new_P2_ADD_391_1196_U159;
  assign new_P2_ADD_391_1196_U223 = new_P2_R2096_U92 | new_P2_R2182_U91;
  assign new_P2_ADD_391_1196_U224 = new_P2_R2096_U93 | new_P2_R2182_U92;
  assign new_P2_ADD_391_1196_U225 = ~new_P2_ADD_391_1196_U83;
  assign new_P2_ADD_391_1196_U226 = ~new_P2_R2096_U92 | ~new_P2_R2182_U91;
  assign new_P2_ADD_391_1196_U227 = ~new_P2_ADD_391_1196_U152;
  assign new_P2_ADD_391_1196_U228 = new_P2_R2182_U90 | new_P2_R2096_U91;
  assign new_P2_ADD_391_1196_U229 = ~new_P2_ADD_391_1196_U228 | ~new_P2_ADD_391_1196_U152;
  assign new_P2_ADD_391_1196_U230 = ~new_P2_R2096_U91 | ~new_P2_R2182_U90;
  assign new_P2_ADD_391_1196_U231 = ~new_P2_ADD_391_1196_U150;
  assign new_P2_ADD_391_1196_U232 = new_P2_R2182_U89 | new_P2_R2096_U90;
  assign new_P2_ADD_391_1196_U233 = ~new_P2_ADD_391_1196_U232 | ~new_P2_ADD_391_1196_U150;
  assign new_P2_ADD_391_1196_U234 = ~new_P2_R2096_U90 | ~new_P2_R2182_U89;
  assign new_P2_ADD_391_1196_U235 = ~new_P2_ADD_391_1196_U148;
  assign new_P2_ADD_391_1196_U236 = new_P2_R2182_U88 | new_P2_R2096_U89;
  assign new_P2_ADD_391_1196_U237 = ~new_P2_ADD_391_1196_U236 | ~new_P2_ADD_391_1196_U148;
  assign new_P2_ADD_391_1196_U238 = ~new_P2_R2096_U89 | ~new_P2_R2182_U88;
  assign new_P2_ADD_391_1196_U239 = ~new_P2_ADD_391_1196_U146;
  assign new_P2_ADD_391_1196_U240 = new_P2_R2182_U87 | new_P2_R2096_U88;
  assign new_P2_ADD_391_1196_U241 = ~new_P2_ADD_391_1196_U240 | ~new_P2_ADD_391_1196_U146;
  assign new_P2_ADD_391_1196_U242 = ~new_P2_R2096_U88 | ~new_P2_R2182_U87;
  assign new_P2_ADD_391_1196_U243 = ~new_P2_ADD_391_1196_U142;
  assign new_P2_ADD_391_1196_U244 = new_P2_R2182_U86 | new_P2_R2096_U87;
  assign new_P2_ADD_391_1196_U245 = ~new_P2_ADD_391_1196_U244 | ~new_P2_ADD_391_1196_U142;
  assign new_P2_ADD_391_1196_U246 = ~new_P2_R2096_U87 | ~new_P2_R2182_U86;
  assign new_P2_ADD_391_1196_U247 = ~new_P2_ADD_391_1196_U140;
  assign new_P2_ADD_391_1196_U248 = new_P2_R2182_U85 | new_P2_R2096_U86;
  assign new_P2_ADD_391_1196_U249 = ~new_P2_ADD_391_1196_U248 | ~new_P2_ADD_391_1196_U140;
  assign new_P2_ADD_391_1196_U250 = ~new_P2_R2096_U86 | ~new_P2_R2182_U85;
  assign new_P2_ADD_391_1196_U251 = ~new_P2_ADD_391_1196_U138;
  assign new_P2_ADD_391_1196_U252 = new_P2_R2182_U84 | new_P2_R2096_U85;
  assign new_P2_ADD_391_1196_U253 = ~new_P2_ADD_391_1196_U252 | ~new_P2_ADD_391_1196_U138;
  assign new_P2_ADD_391_1196_U254 = ~new_P2_R2096_U85 | ~new_P2_R2182_U84;
  assign new_P2_ADD_391_1196_U255 = ~new_P2_ADD_391_1196_U136;
  assign new_P2_ADD_391_1196_U256 = new_P2_R2182_U83 | new_P2_R2096_U84;
  assign new_P2_ADD_391_1196_U257 = ~new_P2_ADD_391_1196_U256 | ~new_P2_ADD_391_1196_U136;
  assign new_P2_ADD_391_1196_U258 = ~new_P2_R2096_U84 | ~new_P2_R2182_U83;
  assign new_P2_ADD_391_1196_U259 = ~new_P2_ADD_391_1196_U134;
  assign new_P2_ADD_391_1196_U260 = new_P2_R2182_U82 | new_P2_R2096_U83;
  assign new_P2_ADD_391_1196_U261 = ~new_P2_ADD_391_1196_U260 | ~new_P2_ADD_391_1196_U134;
  assign new_P2_ADD_391_1196_U262 = ~new_P2_R2096_U83 | ~new_P2_R2182_U82;
  assign new_P2_ADD_391_1196_U263 = ~new_P2_ADD_391_1196_U132;
  assign new_P2_ADD_391_1196_U264 = new_P2_R2182_U81 | new_P2_R2096_U82;
  assign new_P2_ADD_391_1196_U265 = ~new_P2_ADD_391_1196_U264 | ~new_P2_ADD_391_1196_U132;
  assign new_P2_ADD_391_1196_U266 = ~new_P2_R2096_U82 | ~new_P2_R2182_U81;
  assign new_P2_ADD_391_1196_U267 = ~new_P2_ADD_391_1196_U130;
  assign new_P2_ADD_391_1196_U268 = new_P2_R2182_U80 | new_P2_R2096_U81;
  assign new_P2_ADD_391_1196_U269 = ~new_P2_ADD_391_1196_U268 | ~new_P2_ADD_391_1196_U130;
  assign new_P2_ADD_391_1196_U270 = ~new_P2_R2096_U81 | ~new_P2_R2182_U80;
  assign new_P2_ADD_391_1196_U271 = ~new_P2_ADD_391_1196_U128;
  assign new_P2_ADD_391_1196_U272 = new_P2_R2182_U79 | new_P2_R2096_U80;
  assign new_P2_ADD_391_1196_U273 = ~new_P2_ADD_391_1196_U272 | ~new_P2_ADD_391_1196_U128;
  assign new_P2_ADD_391_1196_U274 = ~new_P2_R2096_U80 | ~new_P2_R2182_U79;
  assign new_P2_ADD_391_1196_U275 = ~new_P2_ADD_391_1196_U126;
  assign new_P2_ADD_391_1196_U276 = new_P2_R2096_U79 | new_P2_R2182_U78;
  assign new_P2_ADD_391_1196_U277 = ~new_P2_ADD_391_1196_U276 | ~new_P2_ADD_391_1196_U126;
  assign new_P2_ADD_391_1196_U278 = ~new_P2_R2182_U78 | ~new_P2_R2096_U79;
  assign new_P2_ADD_391_1196_U279 = ~new_P2_ADD_391_1196_U82;
  assign new_P2_ADD_391_1196_U280 = new_P2_R2096_U78 | new_P2_R2182_U77;
  assign new_P2_ADD_391_1196_U281 = ~new_P2_ADD_391_1196_U280 | ~new_P2_ADD_391_1196_U82;
  assign new_P2_ADD_391_1196_U282 = ~new_P2_R2182_U77 | ~new_P2_R2096_U78;
  assign new_P2_ADD_391_1196_U283 = ~new_P2_ADD_391_1196_U121 | ~new_P2_ADD_391_1196_U282 | ~new_P2_ADD_391_1196_U281;
  assign new_P2_ADD_391_1196_U284 = ~new_P2_R2182_U77 | ~new_P2_R2096_U78;
  assign new_P2_ADD_391_1196_U285 = ~new_P2_ADD_391_1196_U279 | ~new_P2_ADD_391_1196_U284;
  assign new_P2_ADD_391_1196_U286 = new_P2_R2182_U77 | new_P2_R2096_U78;
  assign new_P2_ADD_391_1196_U287 = ~new_P2_ADD_391_1196_U343 | ~new_P2_ADD_391_1196_U286 | ~new_P2_ADD_391_1196_U285;
  assign new_P2_ADD_391_1196_U288 = new_P2_R2182_U92 | new_P2_R2096_U93;
  assign new_P2_ADD_391_1196_U289 = ~new_P2_ADD_391_1196_U288 | ~new_P2_ADD_391_1196_U53;
  assign new_P2_ADD_391_1196_U290 = ~new_P2_ADD_391_1196_U153 | ~new_P2_ADD_391_1196_U289 | ~new_P2_ADD_391_1196_U159;
  assign new_P2_ADD_391_1196_U291 = ~new_P2_R2096_U92 | ~new_P2_R2182_U91;
  assign new_P2_ADD_391_1196_U292 = ~new_P2_ADD_391_1196_U225 | ~new_P2_ADD_391_1196_U291;
  assign new_P2_ADD_391_1196_U293 = new_P2_R2096_U93 | new_P2_R2182_U92;
  assign new_P2_ADD_391_1196_U294 = ~new_P2_ADD_391_1196_U154 | ~new_P2_ADD_391_1196_U217;
  assign new_P2_ADD_391_1196_U295 = ~new_P2_R2096_U94 | ~new_P2_R2182_U93;
  assign new_P2_ADD_391_1196_U296 = ~new_P2_ADD_391_1196_U219 | ~new_P2_ADD_391_1196_U295;
  assign new_P2_ADD_391_1196_U297 = new_P2_R2182_U96 | new_P2_R2096_U97;
  assign new_P2_ADD_391_1196_U298 = ~new_P2_ADD_391_1196_U297 | ~new_P2_ADD_391_1196_U50;
  assign new_P2_ADD_391_1196_U299 = ~new_P2_ADD_391_1196_U157 | ~new_P2_ADD_391_1196_U298 | ~new_P2_ADD_391_1196_U158;
  assign new_P2_ADD_391_1196_U300 = ~new_P2_R2096_U96 | ~new_P2_R2182_U95;
  assign new_P2_ADD_391_1196_U301 = ~new_P2_ADD_391_1196_U211 | ~new_P2_ADD_391_1196_U300;
  assign new_P2_ADD_391_1196_U302 = new_P2_R2096_U97 | new_P2_R2182_U96;
  assign new_P2_ADD_391_1196_U303 = ~new_P2_ADD_391_1196_U202 | ~new_P2_ADD_391_1196_U161;
  assign new_P2_ADD_391_1196_U304 = ~new_P2_ADD_391_1196_U293 | ~new_P2_ADD_391_1196_U159;
  assign new_P2_ADD_391_1196_U305 = ~new_P2_ADD_391_1196_U302 | ~new_P2_ADD_391_1196_U158;
  assign new_P2_ADD_391_1196_U306 = ~new_P2_ADD_391_1196_U423 | ~new_P2_ADD_391_1196_U23;
  assign new_P2_ADD_391_1196_U307 = ~new_P2_R2096_U69 | ~new_P2_ADD_391_1196_U34;
  assign new_P2_ADD_391_1196_U308 = ~new_P2_R2182_U70 | ~new_P2_ADD_391_1196_U33;
  assign new_P2_ADD_391_1196_U309 = ~new_P2_R2096_U70 | ~new_P2_ADD_391_1196_U31;
  assign new_P2_ADD_391_1196_U310 = ~new_P2_R2182_U71 | ~new_P2_ADD_391_1196_U32;
  assign new_P2_ADD_391_1196_U311 = ~new_P2_R2096_U70 | ~new_P2_ADD_391_1196_U31;
  assign new_P2_ADD_391_1196_U312 = ~new_P2_R2182_U71 | ~new_P2_ADD_391_1196_U32;
  assign new_P2_ADD_391_1196_U313 = ~new_P2_ADD_391_1196_U312 | ~new_P2_ADD_391_1196_U311;
  assign new_P2_ADD_391_1196_U314 = ~new_P2_ADD_391_1196_U111 | ~new_P2_ADD_391_1196_U112;
  assign new_P2_ADD_391_1196_U315 = ~new_P2_ADD_391_1196_U187 | ~new_P2_ADD_391_1196_U313;
  assign new_P2_ADD_391_1196_U316 = ~new_P2_R2096_U71 | ~new_P2_ADD_391_1196_U13;
  assign new_P2_ADD_391_1196_U317 = ~new_P2_R2182_U72 | ~new_P2_ADD_391_1196_U14;
  assign new_P2_ADD_391_1196_U318 = ~new_P2_R2096_U72 | ~new_P2_ADD_391_1196_U15;
  assign new_P2_ADD_391_1196_U319 = ~new_P2_R2182_U73 | ~new_P2_ADD_391_1196_U16;
  assign new_P2_ADD_391_1196_U320 = ~new_P2_ADD_391_1196_U319 | ~new_P2_ADD_391_1196_U318;
  assign new_P2_ADD_391_1196_U321 = ~new_P2_ADD_391_1196_U303 | ~new_P2_ADD_391_1196_U30;
  assign new_P2_ADD_391_1196_U322 = ~new_P2_ADD_391_1196_U320 | ~new_P2_ADD_391_1196_U181;
  assign new_P2_ADD_391_1196_U323 = ~new_P2_R2096_U73 | ~new_P2_ADD_391_1196_U17;
  assign new_P2_ADD_391_1196_U324 = ~new_P2_R2182_U74 | ~new_P2_ADD_391_1196_U18;
  assign new_P2_ADD_391_1196_U325 = ~new_P2_R2096_U74 | ~new_P2_ADD_391_1196_U28;
  assign new_P2_ADD_391_1196_U326 = ~new_P2_R2182_U75 | ~new_P2_ADD_391_1196_U29;
  assign new_P2_ADD_391_1196_U327 = ~new_P2_R2096_U74 | ~new_P2_ADD_391_1196_U28;
  assign new_P2_ADD_391_1196_U328 = ~new_P2_R2182_U75 | ~new_P2_ADD_391_1196_U29;
  assign new_P2_ADD_391_1196_U329 = ~new_P2_ADD_391_1196_U328 | ~new_P2_ADD_391_1196_U327;
  assign new_P2_ADD_391_1196_U330 = ~new_P2_ADD_391_1196_U115 | ~new_P2_ADD_391_1196_U116;
  assign new_P2_ADD_391_1196_U331 = ~new_P2_ADD_391_1196_U173 | ~new_P2_ADD_391_1196_U329;
  assign new_P2_ADD_391_1196_U332 = ~new_P2_R2096_U75 | ~new_P2_ADD_391_1196_U26;
  assign new_P2_ADD_391_1196_U333 = ~new_P2_R2182_U76 | ~new_P2_ADD_391_1196_U27;
  assign new_P2_ADD_391_1196_U334 = ~new_P2_R2096_U75 | ~new_P2_ADD_391_1196_U26;
  assign new_P2_ADD_391_1196_U335 = ~new_P2_R2182_U76 | ~new_P2_ADD_391_1196_U27;
  assign new_P2_ADD_391_1196_U336 = ~new_P2_ADD_391_1196_U335 | ~new_P2_ADD_391_1196_U334;
  assign new_P2_ADD_391_1196_U337 = ~new_P2_ADD_391_1196_U117 | ~new_P2_ADD_391_1196_U118;
  assign new_P2_ADD_391_1196_U338 = ~new_P2_ADD_391_1196_U169 | ~new_P2_ADD_391_1196_U336;
  assign new_P2_ADD_391_1196_U339 = ~new_P2_R2182_U41 | ~new_P2_ADD_391_1196_U120;
  assign new_P2_ADD_391_1196_U340 = ~new_P2_R2096_U76 | ~new_P2_ADD_391_1196_U119;
  assign new_P2_ADD_391_1196_U341 = ~new_P2_R2182_U41 | ~new_P2_ADD_391_1196_U120;
  assign new_P2_ADD_391_1196_U342 = ~new_P2_R2096_U76 | ~new_P2_ADD_391_1196_U119;
  assign new_P2_ADD_391_1196_U343 = ~new_P2_ADD_391_1196_U342 | ~new_P2_ADD_391_1196_U341;
  assign new_P2_ADD_391_1196_U344 = ~new_P2_R2096_U77 | ~new_P2_ADD_391_1196_U24;
  assign new_P2_ADD_391_1196_U345 = ~new_P2_R2182_U40 | ~new_P2_ADD_391_1196_U25;
  assign new_P2_ADD_391_1196_U346 = ~new_P2_R2096_U77 | ~new_P2_ADD_391_1196_U24;
  assign new_P2_ADD_391_1196_U347 = ~new_P2_R2182_U40 | ~new_P2_ADD_391_1196_U25;
  assign new_P2_ADD_391_1196_U348 = ~new_P2_ADD_391_1196_U347 | ~new_P2_ADD_391_1196_U346;
  assign new_P2_ADD_391_1196_U349 = ~new_P2_ADD_391_1196_U122 | ~new_P2_ADD_391_1196_U123;
  assign new_P2_ADD_391_1196_U350 = ~new_P2_ADD_391_1196_U165 | ~new_P2_ADD_391_1196_U348;
  assign new_P2_ADD_391_1196_U351 = ~new_P2_R2182_U77 | ~new_P2_ADD_391_1196_U80;
  assign new_P2_ADD_391_1196_U352 = ~new_P2_R2096_U78 | ~new_P2_ADD_391_1196_U81;
  assign new_P2_ADD_391_1196_U353 = ~new_P2_R2182_U77 | ~new_P2_ADD_391_1196_U80;
  assign new_P2_ADD_391_1196_U354 = ~new_P2_R2096_U78 | ~new_P2_ADD_391_1196_U81;
  assign new_P2_ADD_391_1196_U355 = ~new_P2_ADD_391_1196_U354 | ~new_P2_ADD_391_1196_U353;
  assign new_P2_ADD_391_1196_U356 = ~new_P2_ADD_391_1196_U124 | ~new_P2_ADD_391_1196_U82;
  assign new_P2_ADD_391_1196_U357 = ~new_P2_ADD_391_1196_U355 | ~new_P2_ADD_391_1196_U279;
  assign new_P2_ADD_391_1196_U358 = ~new_P2_R2182_U78 | ~new_P2_ADD_391_1196_U78;
  assign new_P2_ADD_391_1196_U359 = ~new_P2_R2096_U79 | ~new_P2_ADD_391_1196_U79;
  assign new_P2_ADD_391_1196_U360 = ~new_P2_R2182_U78 | ~new_P2_ADD_391_1196_U78;
  assign new_P2_ADD_391_1196_U361 = ~new_P2_R2096_U79 | ~new_P2_ADD_391_1196_U79;
  assign new_P2_ADD_391_1196_U362 = ~new_P2_ADD_391_1196_U361 | ~new_P2_ADD_391_1196_U360;
  assign new_P2_ADD_391_1196_U363 = ~new_P2_ADD_391_1196_U125 | ~new_P2_ADD_391_1196_U126;
  assign new_P2_ADD_391_1196_U364 = ~new_P2_ADD_391_1196_U275 | ~new_P2_ADD_391_1196_U362;
  assign new_P2_ADD_391_1196_U365 = ~new_P2_R2096_U80 | ~new_P2_ADD_391_1196_U76;
  assign new_P2_ADD_391_1196_U366 = ~new_P2_R2182_U79 | ~new_P2_ADD_391_1196_U77;
  assign new_P2_ADD_391_1196_U367 = ~new_P2_R2096_U80 | ~new_P2_ADD_391_1196_U76;
  assign new_P2_ADD_391_1196_U368 = ~new_P2_R2182_U79 | ~new_P2_ADD_391_1196_U77;
  assign new_P2_ADD_391_1196_U369 = ~new_P2_ADD_391_1196_U368 | ~new_P2_ADD_391_1196_U367;
  assign new_P2_ADD_391_1196_U370 = ~new_P2_ADD_391_1196_U127 | ~new_P2_ADD_391_1196_U128;
  assign new_P2_ADD_391_1196_U371 = ~new_P2_ADD_391_1196_U271 | ~new_P2_ADD_391_1196_U369;
  assign new_P2_ADD_391_1196_U372 = ~new_P2_R2096_U81 | ~new_P2_ADD_391_1196_U74;
  assign new_P2_ADD_391_1196_U373 = ~new_P2_R2182_U80 | ~new_P2_ADD_391_1196_U75;
  assign new_P2_ADD_391_1196_U374 = ~new_P2_R2096_U81 | ~new_P2_ADD_391_1196_U74;
  assign new_P2_ADD_391_1196_U375 = ~new_P2_R2182_U80 | ~new_P2_ADD_391_1196_U75;
  assign new_P2_ADD_391_1196_U376 = ~new_P2_ADD_391_1196_U375 | ~new_P2_ADD_391_1196_U374;
  assign new_P2_ADD_391_1196_U377 = ~new_P2_ADD_391_1196_U129 | ~new_P2_ADD_391_1196_U130;
  assign new_P2_ADD_391_1196_U378 = ~new_P2_ADD_391_1196_U267 | ~new_P2_ADD_391_1196_U376;
  assign new_P2_ADD_391_1196_U379 = ~new_P2_R2096_U82 | ~new_P2_ADD_391_1196_U72;
  assign new_P2_ADD_391_1196_U380 = ~new_P2_R2182_U81 | ~new_P2_ADD_391_1196_U73;
  assign new_P2_ADD_391_1196_U381 = ~new_P2_R2096_U82 | ~new_P2_ADD_391_1196_U72;
  assign new_P2_ADD_391_1196_U382 = ~new_P2_R2182_U81 | ~new_P2_ADD_391_1196_U73;
  assign new_P2_ADD_391_1196_U383 = ~new_P2_ADD_391_1196_U382 | ~new_P2_ADD_391_1196_U381;
  assign new_P2_ADD_391_1196_U384 = ~new_P2_ADD_391_1196_U131 | ~new_P2_ADD_391_1196_U132;
  assign new_P2_ADD_391_1196_U385 = ~new_P2_ADD_391_1196_U263 | ~new_P2_ADD_391_1196_U383;
  assign new_P2_ADD_391_1196_U386 = ~new_P2_R2096_U83 | ~new_P2_ADD_391_1196_U70;
  assign new_P2_ADD_391_1196_U387 = ~new_P2_R2182_U82 | ~new_P2_ADD_391_1196_U71;
  assign new_P2_ADD_391_1196_U388 = ~new_P2_R2096_U83 | ~new_P2_ADD_391_1196_U70;
  assign new_P2_ADD_391_1196_U389 = ~new_P2_R2182_U82 | ~new_P2_ADD_391_1196_U71;
  assign new_P2_ADD_391_1196_U390 = ~new_P2_ADD_391_1196_U389 | ~new_P2_ADD_391_1196_U388;
  assign new_P2_ADD_391_1196_U391 = ~new_P2_ADD_391_1196_U133 | ~new_P2_ADD_391_1196_U134;
  assign new_P2_ADD_391_1196_U392 = ~new_P2_ADD_391_1196_U259 | ~new_P2_ADD_391_1196_U390;
  assign new_P2_ADD_391_1196_U393 = ~new_P2_R2096_U84 | ~new_P2_ADD_391_1196_U68;
  assign new_P2_ADD_391_1196_U394 = ~new_P2_R2182_U83 | ~new_P2_ADD_391_1196_U69;
  assign new_P2_ADD_391_1196_U395 = ~new_P2_R2096_U84 | ~new_P2_ADD_391_1196_U68;
  assign new_P2_ADD_391_1196_U396 = ~new_P2_R2182_U83 | ~new_P2_ADD_391_1196_U69;
  assign new_P2_ADD_391_1196_U397 = ~new_P2_ADD_391_1196_U396 | ~new_P2_ADD_391_1196_U395;
  assign new_P2_ADD_391_1196_U398 = ~new_P2_ADD_391_1196_U135 | ~new_P2_ADD_391_1196_U136;
  assign new_P2_ADD_391_1196_U399 = ~new_P2_ADD_391_1196_U255 | ~new_P2_ADD_391_1196_U397;
  assign new_P2_ADD_391_1196_U400 = ~new_P2_R2096_U85 | ~new_P2_ADD_391_1196_U66;
  assign new_P2_ADD_391_1196_U401 = ~new_P2_R2182_U84 | ~new_P2_ADD_391_1196_U67;
  assign new_P2_ADD_391_1196_U402 = ~new_P2_R2096_U85 | ~new_P2_ADD_391_1196_U66;
  assign new_P2_ADD_391_1196_U403 = ~new_P2_R2182_U84 | ~new_P2_ADD_391_1196_U67;
  assign new_P2_ADD_391_1196_U404 = ~new_P2_ADD_391_1196_U403 | ~new_P2_ADD_391_1196_U402;
  assign new_P2_ADD_391_1196_U405 = ~new_P2_ADD_391_1196_U137 | ~new_P2_ADD_391_1196_U138;
  assign new_P2_ADD_391_1196_U406 = ~new_P2_ADD_391_1196_U251 | ~new_P2_ADD_391_1196_U404;
  assign new_P2_ADD_391_1196_U407 = ~new_P2_R2096_U86 | ~new_P2_ADD_391_1196_U64;
  assign new_P2_ADD_391_1196_U408 = ~new_P2_R2182_U85 | ~new_P2_ADD_391_1196_U65;
  assign new_P2_ADD_391_1196_U409 = ~new_P2_R2096_U86 | ~new_P2_ADD_391_1196_U64;
  assign new_P2_ADD_391_1196_U410 = ~new_P2_R2182_U85 | ~new_P2_ADD_391_1196_U65;
  assign new_P2_ADD_391_1196_U411 = ~new_P2_ADD_391_1196_U410 | ~new_P2_ADD_391_1196_U409;
  assign new_P2_ADD_391_1196_U412 = ~new_P2_ADD_391_1196_U139 | ~new_P2_ADD_391_1196_U140;
  assign new_P2_ADD_391_1196_U413 = ~new_P2_ADD_391_1196_U247 | ~new_P2_ADD_391_1196_U411;
  assign new_P2_ADD_391_1196_U414 = ~new_P2_R2096_U87 | ~new_P2_ADD_391_1196_U62;
  assign new_P2_ADD_391_1196_U415 = ~new_P2_R2182_U86 | ~new_P2_ADD_391_1196_U63;
  assign new_P2_ADD_391_1196_U416 = ~new_P2_R2096_U87 | ~new_P2_ADD_391_1196_U62;
  assign new_P2_ADD_391_1196_U417 = ~new_P2_R2182_U86 | ~new_P2_ADD_391_1196_U63;
  assign new_P2_ADD_391_1196_U418 = ~new_P2_ADD_391_1196_U417 | ~new_P2_ADD_391_1196_U416;
  assign new_P2_ADD_391_1196_U419 = ~new_P2_ADD_391_1196_U141 | ~new_P2_ADD_391_1196_U142;
  assign new_P2_ADD_391_1196_U420 = ~new_P2_ADD_391_1196_U243 | ~new_P2_ADD_391_1196_U418;
  assign new_P2_ADD_391_1196_U421 = ~new_P2_R2182_U68 | ~new_P2_ADD_391_1196_U22;
  assign new_P2_ADD_391_1196_U422 = ~new_P2_ADD_391_1196_U162 | ~new_P2_ADD_391_1196_U21;
  assign new_P2_ADD_391_1196_U423 = ~new_P2_ADD_391_1196_U422 | ~new_P2_ADD_391_1196_U421;
  assign new_P2_ADD_391_1196_U424 = ~new_P2_ADD_391_1196_U21 | ~new_P2_R2096_U51 | ~new_P2_ADD_391_1196_U22;
  assign new_P2_ADD_391_1196_U425 = ~new_P2_ADD_391_1196_U160 | ~new_P2_R2182_U68;
  assign new_P2_ADD_391_1196_U426 = ~new_P2_R2096_U88 | ~new_P2_ADD_391_1196_U60;
  assign new_P2_ADD_391_1196_U427 = ~new_P2_R2182_U87 | ~new_P2_ADD_391_1196_U61;
  assign new_P2_ADD_391_1196_U428 = ~new_P2_R2096_U88 | ~new_P2_ADD_391_1196_U60;
  assign new_P2_ADD_391_1196_U429 = ~new_P2_R2182_U87 | ~new_P2_ADD_391_1196_U61;
  assign new_P2_ADD_391_1196_U430 = ~new_P2_ADD_391_1196_U429 | ~new_P2_ADD_391_1196_U428;
  assign new_P2_ADD_391_1196_U431 = ~new_P2_ADD_391_1196_U145 | ~new_P2_ADD_391_1196_U146;
  assign new_P2_ADD_391_1196_U432 = ~new_P2_ADD_391_1196_U239 | ~new_P2_ADD_391_1196_U430;
  assign new_P2_ADD_391_1196_U433 = ~new_P2_R2096_U89 | ~new_P2_ADD_391_1196_U58;
  assign new_P2_ADD_391_1196_U434 = ~new_P2_R2182_U88 | ~new_P2_ADD_391_1196_U59;
  assign new_P2_ADD_391_1196_U435 = ~new_P2_R2096_U89 | ~new_P2_ADD_391_1196_U58;
  assign new_P2_ADD_391_1196_U436 = ~new_P2_R2182_U88 | ~new_P2_ADD_391_1196_U59;
  assign new_P2_ADD_391_1196_U437 = ~new_P2_ADD_391_1196_U436 | ~new_P2_ADD_391_1196_U435;
  assign new_P2_ADD_391_1196_U438 = ~new_P2_ADD_391_1196_U147 | ~new_P2_ADD_391_1196_U148;
  assign new_P2_ADD_391_1196_U439 = ~new_P2_ADD_391_1196_U235 | ~new_P2_ADD_391_1196_U437;
  assign new_P2_ADD_391_1196_U440 = ~new_P2_R2096_U90 | ~new_P2_ADD_391_1196_U56;
  assign new_P2_ADD_391_1196_U441 = ~new_P2_R2182_U89 | ~new_P2_ADD_391_1196_U57;
  assign new_P2_ADD_391_1196_U442 = ~new_P2_R2096_U90 | ~new_P2_ADD_391_1196_U56;
  assign new_P2_ADD_391_1196_U443 = ~new_P2_R2182_U89 | ~new_P2_ADD_391_1196_U57;
  assign new_P2_ADD_391_1196_U444 = ~new_P2_ADD_391_1196_U443 | ~new_P2_ADD_391_1196_U442;
  assign new_P2_ADD_391_1196_U445 = ~new_P2_ADD_391_1196_U149 | ~new_P2_ADD_391_1196_U150;
  assign new_P2_ADD_391_1196_U446 = ~new_P2_ADD_391_1196_U231 | ~new_P2_ADD_391_1196_U444;
  assign new_P2_ADD_391_1196_U447 = ~new_P2_R2096_U91 | ~new_P2_ADD_391_1196_U54;
  assign new_P2_ADD_391_1196_U448 = ~new_P2_R2182_U90 | ~new_P2_ADD_391_1196_U55;
  assign new_P2_ADD_391_1196_U449 = ~new_P2_R2096_U91 | ~new_P2_ADD_391_1196_U54;
  assign new_P2_ADD_391_1196_U450 = ~new_P2_R2182_U90 | ~new_P2_ADD_391_1196_U55;
  assign new_P2_ADD_391_1196_U451 = ~new_P2_ADD_391_1196_U450 | ~new_P2_ADD_391_1196_U449;
  assign new_P2_ADD_391_1196_U452 = ~new_P2_ADD_391_1196_U151 | ~new_P2_ADD_391_1196_U152;
  assign new_P2_ADD_391_1196_U453 = ~new_P2_ADD_391_1196_U227 | ~new_P2_ADD_391_1196_U451;
  assign new_P2_ADD_391_1196_U454 = ~new_P2_R2096_U92 | ~new_P2_ADD_391_1196_U40;
  assign new_P2_ADD_391_1196_U455 = ~new_P2_R2182_U91 | ~new_P2_ADD_391_1196_U41;
  assign new_P2_ADD_391_1196_U456 = ~new_P2_R2096_U93 | ~new_P2_ADD_391_1196_U42;
  assign new_P2_ADD_391_1196_U457 = ~new_P2_R2182_U92 | ~new_P2_ADD_391_1196_U43;
  assign new_P2_ADD_391_1196_U458 = ~new_P2_ADD_391_1196_U457 | ~new_P2_ADD_391_1196_U456;
  assign new_P2_ADD_391_1196_U459 = ~new_P2_ADD_391_1196_U304 | ~new_P2_ADD_391_1196_U53;
  assign new_P2_ADD_391_1196_U460 = ~new_P2_ADD_391_1196_U458 | ~new_P2_ADD_391_1196_U221;
  assign new_P2_ADD_391_1196_U461 = ~new_P2_R2096_U94 | ~new_P2_ADD_391_1196_U44;
  assign new_P2_ADD_391_1196_U462 = ~new_P2_R2182_U93 | ~new_P2_ADD_391_1196_U45;
  assign new_P2_ADD_391_1196_U463 = ~new_P2_R2096_U95 | ~new_P2_ADD_391_1196_U51;
  assign new_P2_ADD_391_1196_U464 = ~new_P2_R2182_U94 | ~new_P2_ADD_391_1196_U52;
  assign new_P2_ADD_391_1196_U465 = ~new_P2_R2096_U95 | ~new_P2_ADD_391_1196_U51;
  assign new_P2_ADD_391_1196_U466 = ~new_P2_R2182_U94 | ~new_P2_ADD_391_1196_U52;
  assign new_P2_ADD_391_1196_U467 = ~new_P2_ADD_391_1196_U466 | ~new_P2_ADD_391_1196_U465;
  assign new_P2_ADD_391_1196_U468 = ~new_P2_ADD_391_1196_U155 | ~new_P2_ADD_391_1196_U156;
  assign new_P2_ADD_391_1196_U469 = ~new_P2_ADD_391_1196_U213 | ~new_P2_ADD_391_1196_U467;
  assign new_P2_ADD_391_1196_U470 = ~new_P2_R2096_U96 | ~new_P2_ADD_391_1196_U46;
  assign new_P2_ADD_391_1196_U471 = ~new_P2_R2182_U95 | ~new_P2_ADD_391_1196_U47;
  assign new_P2_ADD_391_1196_U472 = ~new_P2_R2096_U97 | ~new_P2_ADD_391_1196_U48;
  assign new_P2_ADD_391_1196_U473 = ~new_P2_R2182_U96 | ~new_P2_ADD_391_1196_U49;
  assign new_P2_ADD_391_1196_U474 = ~new_P2_ADD_391_1196_U473 | ~new_P2_ADD_391_1196_U472;
  assign new_P2_ADD_391_1196_U475 = ~new_P2_ADD_391_1196_U305 | ~new_P2_ADD_391_1196_U50;
  assign new_P2_ADD_391_1196_U476 = ~new_P2_ADD_391_1196_U474 | ~new_P2_ADD_391_1196_U207;
  assign new_P2_ADD_391_1196_U477 = ~new_P2_R2182_U69 | ~new_P2_ADD_391_1196_U19;
  assign new_P2_ADD_391_1196_U478 = ~new_P2_R2096_U68 | ~new_P2_ADD_391_1196_U20;
  assign new_P2_ADD_402_1132_U4 = ~new_P2_U2606;
  assign new_P2_ADD_402_1132_U5 = ~new_P2_U2591;
  assign new_P2_ADD_402_1132_U6 = ~new_P2_U2591 | ~new_P2_U2606;
  assign new_P2_ADD_402_1132_U7 = ~new_P2_U2592;
  assign new_P2_ADD_402_1132_U8 = ~new_P2_U2592 | ~new_P2_ADD_402_1132_U28;
  assign new_P2_ADD_402_1132_U9 = ~new_P2_U2593;
  assign new_P2_ADD_402_1132_U10 = ~new_P2_U2593 | ~new_P2_ADD_402_1132_U29;
  assign new_P2_ADD_402_1132_U11 = ~new_P2_U2594;
  assign new_P2_ADD_402_1132_U12 = ~new_P2_U2594 | ~new_P2_ADD_402_1132_U30;
  assign new_P2_ADD_402_1132_U13 = ~new_P2_U2595;
  assign new_P2_ADD_402_1132_U14 = ~new_P2_U2595 | ~new_P2_ADD_402_1132_U31;
  assign new_P2_ADD_402_1132_U15 = ~new_P2_U2596;
  assign new_P2_ADD_402_1132_U16 = ~new_P2_U2596 | ~new_P2_ADD_402_1132_U32;
  assign new_P2_ADD_402_1132_U17 = ~new_P2_U2597;
  assign new_P2_ADD_402_1132_U18 = ~new_P2_ADD_402_1132_U36 | ~new_P2_ADD_402_1132_U35;
  assign new_P2_ADD_402_1132_U19 = ~new_P2_ADD_402_1132_U38 | ~new_P2_ADD_402_1132_U37;
  assign new_P2_ADD_402_1132_U20 = ~new_P2_ADD_402_1132_U40 | ~new_P2_ADD_402_1132_U39;
  assign new_P2_ADD_402_1132_U21 = ~new_P2_ADD_402_1132_U42 | ~new_P2_ADD_402_1132_U41;
  assign new_P2_ADD_402_1132_U22 = ~new_P2_ADD_402_1132_U44 | ~new_P2_ADD_402_1132_U43;
  assign new_P2_ADD_402_1132_U23 = ~new_P2_ADD_402_1132_U46 | ~new_P2_ADD_402_1132_U45;
  assign new_P2_ADD_402_1132_U24 = ~new_P2_ADD_402_1132_U48 | ~new_P2_ADD_402_1132_U47;
  assign new_P2_ADD_402_1132_U25 = ~new_P2_ADD_402_1132_U50 | ~new_P2_ADD_402_1132_U49;
  assign new_P2_ADD_402_1132_U26 = ~new_P2_U2598;
  assign new_P2_ADD_402_1132_U27 = ~new_P2_U2597 | ~new_P2_ADD_402_1132_U33;
  assign new_P2_ADD_402_1132_U28 = ~new_P2_ADD_402_1132_U6;
  assign new_P2_ADD_402_1132_U29 = ~new_P2_ADD_402_1132_U8;
  assign new_P2_ADD_402_1132_U30 = ~new_P2_ADD_402_1132_U10;
  assign new_P2_ADD_402_1132_U31 = ~new_P2_ADD_402_1132_U12;
  assign new_P2_ADD_402_1132_U32 = ~new_P2_ADD_402_1132_U14;
  assign new_P2_ADD_402_1132_U33 = ~new_P2_ADD_402_1132_U16;
  assign new_P2_ADD_402_1132_U34 = ~new_P2_ADD_402_1132_U27;
  assign new_P2_ADD_402_1132_U35 = ~new_P2_U2598 | ~new_P2_ADD_402_1132_U27;
  assign new_P2_ADD_402_1132_U36 = ~new_P2_ADD_402_1132_U34 | ~new_P2_ADD_402_1132_U26;
  assign new_P2_ADD_402_1132_U37 = ~new_P2_U2597 | ~new_P2_ADD_402_1132_U16;
  assign new_P2_ADD_402_1132_U38 = ~new_P2_ADD_402_1132_U33 | ~new_P2_ADD_402_1132_U17;
  assign new_P2_ADD_402_1132_U39 = ~new_P2_U2592 | ~new_P2_ADD_402_1132_U6;
  assign new_P2_ADD_402_1132_U40 = ~new_P2_ADD_402_1132_U28 | ~new_P2_ADD_402_1132_U7;
  assign new_P2_ADD_402_1132_U41 = ~new_P2_U2594 | ~new_P2_ADD_402_1132_U10;
  assign new_P2_ADD_402_1132_U42 = ~new_P2_ADD_402_1132_U30 | ~new_P2_ADD_402_1132_U11;
  assign new_P2_ADD_402_1132_U43 = ~new_P2_U2595 | ~new_P2_ADD_402_1132_U12;
  assign new_P2_ADD_402_1132_U44 = ~new_P2_ADD_402_1132_U31 | ~new_P2_ADD_402_1132_U13;
  assign new_P2_ADD_402_1132_U45 = ~new_P2_U2591 | ~new_P2_ADD_402_1132_U4;
  assign new_P2_ADD_402_1132_U46 = ~new_P2_U2606 | ~new_P2_ADD_402_1132_U5;
  assign new_P2_ADD_402_1132_U47 = ~new_P2_U2596 | ~new_P2_ADD_402_1132_U14;
  assign new_P2_ADD_402_1132_U48 = ~new_P2_ADD_402_1132_U32 | ~new_P2_ADD_402_1132_U15;
  assign new_P2_ADD_402_1132_U49 = ~new_P2_U2593 | ~new_P2_ADD_402_1132_U8;
  assign new_P2_ADD_402_1132_U50 = ~new_P2_ADD_402_1132_U29 | ~new_P2_ADD_402_1132_U9;
  assign new_P2_SUB_563_U6 = ~new_P2_U3618;
  assign new_P2_SUB_563_U7 = ~new_P2_U3619;
  assign new_P2_R2182_U4 = new_P2_U2671 & new_P2_R2182_U20;
  assign new_P2_R2182_U5 = new_P2_U2670 & new_P2_R2182_U4;
  assign new_P2_R2182_U6 = new_P2_U2669 & new_P2_R2182_U5;
  assign new_P2_R2182_U7 = new_P2_U2690 & new_P2_R2182_U8;
  assign new_P2_R2182_U8 = new_P2_U2691 & new_P2_R2182_U11;
  assign new_P2_R2182_U9 = new_P2_U2675 & new_P2_R2182_U21;
  assign new_P2_R2182_U10 = new_P2_U2674 & new_P2_R2182_U9;
  assign new_P2_R2182_U11 = new_P2_U2692 & new_P2_R2182_U13;
  assign new_P2_R2182_U12 = new_P2_U2694 & new_P2_R2182_U18;
  assign new_P2_R2182_U13 = new_P2_U2693 & new_P2_R2182_U12;
  assign new_P2_R2182_U14 = new_P2_U2668 & new_P2_R2182_U6;
  assign new_P2_R2182_U15 = new_P2_U2667 & new_P2_R2182_U14;
  assign new_P2_R2182_U16 = new_P2_U2666 & new_P2_R2182_U15;
  assign new_P2_R2182_U17 = new_P2_U2696 & new_P2_R2182_U16;
  assign new_P2_R2182_U18 = new_P2_U2695 & new_P2_R2182_U17;
  assign new_P2_R2182_U19 = new_P2_U2673 & new_P2_R2182_U10;
  assign new_P2_R2182_U20 = new_P2_U2672 & new_P2_R2182_U19;
  assign new_P2_R2182_U21 = new_P2_U2676 & new_P2_R2182_U102;
  assign new_P2_R2182_U22 = ~new_P2_U2675;
  assign new_P2_R2182_U23 = ~new_P2_U2671;
  assign new_P2_R2182_U24 = ~new_P2_U2676;
  assign new_P2_R2182_U25 = ~new_P2_U2666;
  assign new_P2_R2182_U26 = ~new_P2_U2667;
  assign new_P2_R2182_U27 = ~new_P2_U2696;
  assign new_P2_R2182_U28 = ~new_P2_U2695;
  assign new_P2_R2182_U29 = ~new_P2_U2694;
  assign new_P2_R2182_U30 = ~new_P2_U2693;
  assign new_P2_R2182_U31 = ~new_P2_U2692;
  assign new_P2_R2182_U32 = ~new_P2_U2691;
  assign new_P2_R2182_U33 = ~new_P2_U2670;
  assign new_P2_R2182_U34 = ~new_P2_U2672;
  assign new_P2_R2182_U35 = ~new_P2_U2674;
  assign new_P2_R2182_U36 = ~new_P2_U2673;
  assign new_P2_R2182_U37 = ~new_P2_U2690;
  assign new_P2_R2182_U38 = ~new_P2_U2668;
  assign new_P2_R2182_U39 = ~new_P2_U2669;
  assign new_P2_R2182_U40 = new_P2_R2182_U192 & new_P2_R2182_U190;
  assign new_P2_R2182_U41 = new_P2_R2182_U186 & new_P2_R2182_U182;
  assign new_P2_R2182_U42 = ~new_P2_U2700;
  assign new_P2_R2182_U43 = ~new_P2_U2679;
  assign new_P2_R2182_U44 = ~new_P2_U2702;
  assign new_P2_R2182_U45 = ~new_P2_U2681;
  assign new_P2_R2182_U46 = ~new_P2_U2681 | ~new_P2_U2702;
  assign new_P2_R2182_U47 = ~new_P2_U2680;
  assign new_P2_R2182_U48 = ~new_P2_U2699;
  assign new_P2_R2182_U49 = ~new_P2_U2678;
  assign new_P2_R2182_U50 = ~new_P2_U2698;
  assign new_P2_R2182_U51 = ~new_P2_U2677;
  assign new_P2_R2182_U52 = ~new_P2_U2689;
  assign new_P2_R2182_U53 = ~new_P2_U2665;
  assign new_P2_R2182_U54 = ~new_P2_U2688;
  assign new_P2_R2182_U55 = ~new_P2_U2664;
  assign new_P2_R2182_U56 = ~new_P2_U2687;
  assign new_P2_R2182_U57 = ~new_P2_U2663;
  assign new_P2_R2182_U58 = ~new_P2_U2686;
  assign new_P2_R2182_U59 = ~new_P2_U2662;
  assign new_P2_R2182_U60 = ~new_P2_U2685;
  assign new_P2_R2182_U61 = ~new_P2_U2661;
  assign new_P2_R2182_U62 = ~new_P2_U2684;
  assign new_P2_R2182_U63 = ~new_P2_U2660;
  assign new_P2_R2182_U64 = ~new_P2_U2683;
  assign new_P2_R2182_U65 = ~new_P2_U2659;
  assign new_P2_R2182_U66 = ~new_P2_R2182_U177 | ~new_P2_R2182_U176;
  assign new_P2_R2182_U67 = ~new_P2_U2701;
  assign new_P2_R2182_U68 = ~new_P2_R2182_U283 | ~new_P2_R2182_U282;
  assign new_P2_R2182_U69 = ~new_P2_R2182_U305 | ~new_P2_R2182_U304;
  assign new_P2_R2182_U70 = ~new_P2_R2182_U194 | ~new_P2_R2182_U193;
  assign new_P2_R2182_U71 = ~new_P2_R2182_U196 | ~new_P2_R2182_U195;
  assign new_P2_R2182_U72 = ~new_P2_R2182_U198 | ~new_P2_R2182_U197;
  assign new_P2_R2182_U73 = ~new_P2_R2182_U200 | ~new_P2_R2182_U199;
  assign new_P2_R2182_U74 = ~new_P2_R2182_U202 | ~new_P2_R2182_U201;
  assign new_P2_R2182_U75 = ~new_P2_R2182_U209 | ~new_P2_R2182_U208;
  assign new_P2_R2182_U76 = ~new_P2_R2182_U216 | ~new_P2_R2182_U215;
  assign new_P2_R2182_U77 = ~new_P2_R2182_U230 | ~new_P2_R2182_U229;
  assign new_P2_R2182_U78 = ~new_P2_R2182_U237 | ~new_P2_R2182_U236;
  assign new_P2_R2182_U79 = ~new_P2_R2182_U244 | ~new_P2_R2182_U243;
  assign new_P2_R2182_U80 = ~new_P2_R2182_U251 | ~new_P2_R2182_U250;
  assign new_P2_R2182_U81 = ~new_P2_R2182_U258 | ~new_P2_R2182_U257;
  assign new_P2_R2182_U82 = ~new_P2_R2182_U265 | ~new_P2_R2182_U264;
  assign new_P2_R2182_U83 = ~new_P2_R2182_U272 | ~new_P2_R2182_U271;
  assign new_P2_R2182_U84 = ~new_P2_R2182_U274 | ~new_P2_R2182_U273;
  assign new_P2_R2182_U85 = ~new_P2_R2182_U276 | ~new_P2_R2182_U275;
  assign new_P2_R2182_U86 = ~new_P2_R2182_U278 | ~new_P2_R2182_U277;
  assign new_P2_R2182_U87 = ~new_P2_R2182_U285 | ~new_P2_R2182_U284;
  assign new_P2_R2182_U88 = ~new_P2_R2182_U287 | ~new_P2_R2182_U286;
  assign new_P2_R2182_U89 = ~new_P2_R2182_U289 | ~new_P2_R2182_U288;
  assign new_P2_R2182_U90 = ~new_P2_R2182_U291 | ~new_P2_R2182_U290;
  assign new_P2_R2182_U91 = ~new_P2_R2182_U293 | ~new_P2_R2182_U292;
  assign new_P2_R2182_U92 = ~new_P2_R2182_U295 | ~new_P2_R2182_U294;
  assign new_P2_R2182_U93 = ~new_P2_R2182_U297 | ~new_P2_R2182_U296;
  assign new_P2_R2182_U94 = ~new_P2_R2182_U299 | ~new_P2_R2182_U298;
  assign new_P2_R2182_U95 = ~new_P2_R2182_U301 | ~new_P2_R2182_U300;
  assign new_P2_R2182_U96 = ~new_P2_R2182_U303 | ~new_P2_R2182_U302;
  assign new_P2_R2182_U97 = new_P2_R2182_U181 & new_P2_R2182_U218 & new_P2_R2182_U217;
  assign new_P2_R2182_U98 = new_P2_R2182_U185 & new_P2_R2182_U221;
  assign new_P2_R2182_U99 = new_P2_R2182_U189 & new_P2_R2182_U223 & new_P2_R2182_U222;
  assign new_P2_R2182_U100 = new_P2_R2182_U191 & new_P2_R2182_U125;
  assign new_P2_R2182_U101 = ~new_P2_R2182_U280 | ~new_P2_R2182_U279;
  assign new_P2_R2182_U102 = ~new_P2_R2182_U135 | ~new_P2_R2182_U134;
  assign new_P2_R2182_U103 = new_P2_R2182_U204 & new_P2_R2182_U203;
  assign new_P2_R2182_U104 = ~new_P2_R2182_U131 | ~new_P2_R2182_U130;
  assign new_P2_R2182_U105 = new_P2_R2182_U211 & new_P2_R2182_U210;
  assign new_P2_R2182_U106 = ~new_P2_R2182_U126 | ~new_P2_R2182_U127;
  assign new_P2_R2182_U107 = ~new_P2_U2658;
  assign new_P2_R2182_U108 = ~new_P2_U2682;
  assign new_P2_R2182_U109 = new_P2_R2182_U225 & new_P2_R2182_U224;
  assign new_P2_R2182_U110 = new_P2_R2182_U232 & new_P2_R2182_U231;
  assign new_P2_R2182_U111 = ~new_P2_R2182_U173 | ~new_P2_R2182_U172;
  assign new_P2_R2182_U112 = new_P2_R2182_U239 & new_P2_R2182_U238;
  assign new_P2_R2182_U113 = ~new_P2_R2182_U169 | ~new_P2_R2182_U168;
  assign new_P2_R2182_U114 = new_P2_R2182_U246 & new_P2_R2182_U245;
  assign new_P2_R2182_U115 = ~new_P2_R2182_U165 | ~new_P2_R2182_U164;
  assign new_P2_R2182_U116 = new_P2_R2182_U253 & new_P2_R2182_U252;
  assign new_P2_R2182_U117 = ~new_P2_R2182_U161 | ~new_P2_R2182_U160;
  assign new_P2_R2182_U118 = new_P2_R2182_U260 & new_P2_R2182_U259;
  assign new_P2_R2182_U119 = ~new_P2_R2182_U157 | ~new_P2_R2182_U156;
  assign new_P2_R2182_U120 = new_P2_R2182_U267 & new_P2_R2182_U266;
  assign new_P2_R2182_U121 = ~new_P2_R2182_U46;
  assign new_P2_R2182_U122 = ~new_P2_U2680 | ~new_P2_R2182_U121;
  assign new_P2_R2182_U123 = ~new_P2_R2182_U122 | ~new_P2_R2182_U67;
  assign new_P2_R2182_U124 = new_P2_U2679 | new_P2_U2700;
  assign new_P2_R2182_U125 = ~new_P2_R2182_U46 | ~new_P2_R2182_U47;
  assign new_P2_R2182_U126 = ~new_P2_R2182_U124 | ~new_P2_R2182_U125 | ~new_P2_R2182_U123;
  assign new_P2_R2182_U127 = ~new_P2_U2679 | ~new_P2_U2700;
  assign new_P2_R2182_U128 = ~new_P2_R2182_U106;
  assign new_P2_R2182_U129 = new_P2_U2699 | new_P2_U2678;
  assign new_P2_R2182_U130 = ~new_P2_R2182_U129 | ~new_P2_R2182_U106;
  assign new_P2_R2182_U131 = ~new_P2_U2678 | ~new_P2_U2699;
  assign new_P2_R2182_U132 = ~new_P2_R2182_U104;
  assign new_P2_R2182_U133 = new_P2_U2698 | new_P2_U2677;
  assign new_P2_R2182_U134 = ~new_P2_R2182_U133 | ~new_P2_R2182_U104;
  assign new_P2_R2182_U135 = ~new_P2_U2677 | ~new_P2_U2698;
  assign new_P2_R2182_U136 = ~new_P2_R2182_U102;
  assign new_P2_R2182_U137 = ~new_P2_R2182_U21;
  assign new_P2_R2182_U138 = ~new_P2_R2182_U9;
  assign new_P2_R2182_U139 = ~new_P2_R2182_U10;
  assign new_P2_R2182_U140 = ~new_P2_R2182_U19;
  assign new_P2_R2182_U141 = ~new_P2_R2182_U20;
  assign new_P2_R2182_U142 = ~new_P2_R2182_U4;
  assign new_P2_R2182_U143 = ~new_P2_R2182_U5;
  assign new_P2_R2182_U144 = ~new_P2_R2182_U6;
  assign new_P2_R2182_U145 = ~new_P2_R2182_U14;
  assign new_P2_R2182_U146 = ~new_P2_R2182_U15;
  assign new_P2_R2182_U147 = ~new_P2_R2182_U16;
  assign new_P2_R2182_U148 = ~new_P2_R2182_U17;
  assign new_P2_R2182_U149 = ~new_P2_R2182_U18;
  assign new_P2_R2182_U150 = ~new_P2_R2182_U12;
  assign new_P2_R2182_U151 = ~new_P2_R2182_U13;
  assign new_P2_R2182_U152 = ~new_P2_R2182_U11;
  assign new_P2_R2182_U153 = ~new_P2_R2182_U8;
  assign new_P2_R2182_U154 = ~new_P2_R2182_U7;
  assign new_P2_R2182_U155 = new_P2_U2689 | new_P2_U2665;
  assign new_P2_R2182_U156 = ~new_P2_R2182_U155 | ~new_P2_R2182_U7;
  assign new_P2_R2182_U157 = ~new_P2_U2665 | ~new_P2_U2689;
  assign new_P2_R2182_U158 = ~new_P2_R2182_U119;
  assign new_P2_R2182_U159 = new_P2_U2688 | new_P2_U2664;
  assign new_P2_R2182_U160 = ~new_P2_R2182_U159 | ~new_P2_R2182_U119;
  assign new_P2_R2182_U161 = ~new_P2_U2664 | ~new_P2_U2688;
  assign new_P2_R2182_U162 = ~new_P2_R2182_U117;
  assign new_P2_R2182_U163 = new_P2_U2687 | new_P2_U2663;
  assign new_P2_R2182_U164 = ~new_P2_R2182_U163 | ~new_P2_R2182_U117;
  assign new_P2_R2182_U165 = ~new_P2_U2663 | ~new_P2_U2687;
  assign new_P2_R2182_U166 = ~new_P2_R2182_U115;
  assign new_P2_R2182_U167 = new_P2_U2686 | new_P2_U2662;
  assign new_P2_R2182_U168 = ~new_P2_R2182_U167 | ~new_P2_R2182_U115;
  assign new_P2_R2182_U169 = ~new_P2_U2662 | ~new_P2_U2686;
  assign new_P2_R2182_U170 = ~new_P2_R2182_U113;
  assign new_P2_R2182_U171 = new_P2_U2685 | new_P2_U2661;
  assign new_P2_R2182_U172 = ~new_P2_R2182_U171 | ~new_P2_R2182_U113;
  assign new_P2_R2182_U173 = ~new_P2_U2661 | ~new_P2_U2685;
  assign new_P2_R2182_U174 = ~new_P2_R2182_U111;
  assign new_P2_R2182_U175 = new_P2_U2684 | new_P2_U2660;
  assign new_P2_R2182_U176 = ~new_P2_R2182_U175 | ~new_P2_R2182_U111;
  assign new_P2_R2182_U177 = ~new_P2_U2660 | ~new_P2_U2684;
  assign new_P2_R2182_U178 = ~new_P2_R2182_U66;
  assign new_P2_R2182_U179 = new_P2_U2683 | new_P2_U2659;
  assign new_P2_R2182_U180 = ~new_P2_R2182_U179 | ~new_P2_R2182_U66;
  assign new_P2_R2182_U181 = ~new_P2_U2659 | ~new_P2_U2683;
  assign new_P2_R2182_U182 = ~new_P2_R2182_U97 | ~new_P2_R2182_U180;
  assign new_P2_R2182_U183 = ~new_P2_U2659 | ~new_P2_U2683;
  assign new_P2_R2182_U184 = ~new_P2_R2182_U178 | ~new_P2_R2182_U183;
  assign new_P2_R2182_U185 = new_P2_U2659 | new_P2_U2683;
  assign new_P2_R2182_U186 = ~new_P2_R2182_U98 | ~new_P2_R2182_U184;
  assign new_P2_R2182_U187 = ~new_P2_R2182_U47 | ~new_P2_R2182_U46;
  assign new_P2_R2182_U188 = ~new_P2_U2701 | ~new_P2_R2182_U187;
  assign new_P2_R2182_U189 = ~new_P2_U2680 | ~new_P2_R2182_U121;
  assign new_P2_R2182_U190 = ~new_P2_R2182_U99 | ~new_P2_R2182_U188;
  assign new_P2_R2182_U191 = ~new_P2_U2679 | ~new_P2_U2700;
  assign new_P2_R2182_U192 = ~new_P2_R2182_U100 | ~new_P2_R2182_U124 | ~new_P2_R2182_U123;
  assign new_P2_R2182_U193 = ~new_P2_R2182_U34 | ~new_P2_R2182_U19;
  assign new_P2_R2182_U194 = ~new_P2_R2182_U140 | ~new_P2_U2672;
  assign new_P2_R2182_U195 = ~new_P2_R2182_U36 | ~new_P2_R2182_U10;
  assign new_P2_R2182_U196 = ~new_P2_R2182_U139 | ~new_P2_U2673;
  assign new_P2_R2182_U197 = ~new_P2_R2182_U35 | ~new_P2_R2182_U9;
  assign new_P2_R2182_U198 = ~new_P2_R2182_U138 | ~new_P2_U2674;
  assign new_P2_R2182_U199 = ~new_P2_R2182_U22 | ~new_P2_R2182_U21;
  assign new_P2_R2182_U200 = ~new_P2_R2182_U137 | ~new_P2_U2675;
  assign new_P2_R2182_U201 = ~new_P2_R2182_U24 | ~new_P2_R2182_U102;
  assign new_P2_R2182_U202 = ~new_P2_R2182_U136 | ~new_P2_U2676;
  assign new_P2_R2182_U203 = ~new_P2_U2677 | ~new_P2_R2182_U50;
  assign new_P2_R2182_U204 = ~new_P2_U2698 | ~new_P2_R2182_U51;
  assign new_P2_R2182_U205 = ~new_P2_U2677 | ~new_P2_R2182_U50;
  assign new_P2_R2182_U206 = ~new_P2_U2698 | ~new_P2_R2182_U51;
  assign new_P2_R2182_U207 = ~new_P2_R2182_U206 | ~new_P2_R2182_U205;
  assign new_P2_R2182_U208 = ~new_P2_R2182_U103 | ~new_P2_R2182_U104;
  assign new_P2_R2182_U209 = ~new_P2_R2182_U132 | ~new_P2_R2182_U207;
  assign new_P2_R2182_U210 = ~new_P2_U2678 | ~new_P2_R2182_U48;
  assign new_P2_R2182_U211 = ~new_P2_U2699 | ~new_P2_R2182_U49;
  assign new_P2_R2182_U212 = ~new_P2_U2678 | ~new_P2_R2182_U48;
  assign new_P2_R2182_U213 = ~new_P2_U2699 | ~new_P2_R2182_U49;
  assign new_P2_R2182_U214 = ~new_P2_R2182_U213 | ~new_P2_R2182_U212;
  assign new_P2_R2182_U215 = ~new_P2_R2182_U105 | ~new_P2_R2182_U106;
  assign new_P2_R2182_U216 = ~new_P2_R2182_U128 | ~new_P2_R2182_U214;
  assign new_P2_R2182_U217 = ~new_P2_U2658 | ~new_P2_R2182_U108;
  assign new_P2_R2182_U218 = ~new_P2_U2682 | ~new_P2_R2182_U107;
  assign new_P2_R2182_U219 = ~new_P2_U2658 | ~new_P2_R2182_U108;
  assign new_P2_R2182_U220 = ~new_P2_U2682 | ~new_P2_R2182_U107;
  assign new_P2_R2182_U221 = ~new_P2_R2182_U220 | ~new_P2_R2182_U219;
  assign new_P2_R2182_U222 = ~new_P2_U2679 | ~new_P2_R2182_U42;
  assign new_P2_R2182_U223 = ~new_P2_U2700 | ~new_P2_R2182_U43;
  assign new_P2_R2182_U224 = ~new_P2_U2659 | ~new_P2_R2182_U64;
  assign new_P2_R2182_U225 = ~new_P2_U2683 | ~new_P2_R2182_U65;
  assign new_P2_R2182_U226 = ~new_P2_U2659 | ~new_P2_R2182_U64;
  assign new_P2_R2182_U227 = ~new_P2_U2683 | ~new_P2_R2182_U65;
  assign new_P2_R2182_U228 = ~new_P2_R2182_U227 | ~new_P2_R2182_U226;
  assign new_P2_R2182_U229 = ~new_P2_R2182_U109 | ~new_P2_R2182_U66;
  assign new_P2_R2182_U230 = ~new_P2_R2182_U228 | ~new_P2_R2182_U178;
  assign new_P2_R2182_U231 = ~new_P2_U2660 | ~new_P2_R2182_U62;
  assign new_P2_R2182_U232 = ~new_P2_U2684 | ~new_P2_R2182_U63;
  assign new_P2_R2182_U233 = ~new_P2_U2660 | ~new_P2_R2182_U62;
  assign new_P2_R2182_U234 = ~new_P2_U2684 | ~new_P2_R2182_U63;
  assign new_P2_R2182_U235 = ~new_P2_R2182_U234 | ~new_P2_R2182_U233;
  assign new_P2_R2182_U236 = ~new_P2_R2182_U110 | ~new_P2_R2182_U111;
  assign new_P2_R2182_U237 = ~new_P2_R2182_U174 | ~new_P2_R2182_U235;
  assign new_P2_R2182_U238 = ~new_P2_U2661 | ~new_P2_R2182_U60;
  assign new_P2_R2182_U239 = ~new_P2_U2685 | ~new_P2_R2182_U61;
  assign new_P2_R2182_U240 = ~new_P2_U2661 | ~new_P2_R2182_U60;
  assign new_P2_R2182_U241 = ~new_P2_U2685 | ~new_P2_R2182_U61;
  assign new_P2_R2182_U242 = ~new_P2_R2182_U241 | ~new_P2_R2182_U240;
  assign new_P2_R2182_U243 = ~new_P2_R2182_U112 | ~new_P2_R2182_U113;
  assign new_P2_R2182_U244 = ~new_P2_R2182_U170 | ~new_P2_R2182_U242;
  assign new_P2_R2182_U245 = ~new_P2_U2662 | ~new_P2_R2182_U58;
  assign new_P2_R2182_U246 = ~new_P2_U2686 | ~new_P2_R2182_U59;
  assign new_P2_R2182_U247 = ~new_P2_U2662 | ~new_P2_R2182_U58;
  assign new_P2_R2182_U248 = ~new_P2_U2686 | ~new_P2_R2182_U59;
  assign new_P2_R2182_U249 = ~new_P2_R2182_U248 | ~new_P2_R2182_U247;
  assign new_P2_R2182_U250 = ~new_P2_R2182_U114 | ~new_P2_R2182_U115;
  assign new_P2_R2182_U251 = ~new_P2_R2182_U166 | ~new_P2_R2182_U249;
  assign new_P2_R2182_U252 = ~new_P2_U2663 | ~new_P2_R2182_U56;
  assign new_P2_R2182_U253 = ~new_P2_U2687 | ~new_P2_R2182_U57;
  assign new_P2_R2182_U254 = ~new_P2_U2663 | ~new_P2_R2182_U56;
  assign new_P2_R2182_U255 = ~new_P2_U2687 | ~new_P2_R2182_U57;
  assign new_P2_R2182_U256 = ~new_P2_R2182_U255 | ~new_P2_R2182_U254;
  assign new_P2_R2182_U257 = ~new_P2_R2182_U116 | ~new_P2_R2182_U117;
  assign new_P2_R2182_U258 = ~new_P2_R2182_U162 | ~new_P2_R2182_U256;
  assign new_P2_R2182_U259 = ~new_P2_U2664 | ~new_P2_R2182_U54;
  assign new_P2_R2182_U260 = ~new_P2_U2688 | ~new_P2_R2182_U55;
  assign new_P2_R2182_U261 = ~new_P2_U2664 | ~new_P2_R2182_U54;
  assign new_P2_R2182_U262 = ~new_P2_U2688 | ~new_P2_R2182_U55;
  assign new_P2_R2182_U263 = ~new_P2_R2182_U262 | ~new_P2_R2182_U261;
  assign new_P2_R2182_U264 = ~new_P2_R2182_U118 | ~new_P2_R2182_U119;
  assign new_P2_R2182_U265 = ~new_P2_R2182_U158 | ~new_P2_R2182_U263;
  assign new_P2_R2182_U266 = ~new_P2_U2665 | ~new_P2_R2182_U52;
  assign new_P2_R2182_U267 = ~new_P2_U2689 | ~new_P2_R2182_U53;
  assign new_P2_R2182_U268 = ~new_P2_U2665 | ~new_P2_R2182_U52;
  assign new_P2_R2182_U269 = ~new_P2_U2689 | ~new_P2_R2182_U53;
  assign new_P2_R2182_U270 = ~new_P2_R2182_U269 | ~new_P2_R2182_U268;
  assign new_P2_R2182_U271 = ~new_P2_R2182_U120 | ~new_P2_R2182_U7;
  assign new_P2_R2182_U272 = ~new_P2_R2182_U154 | ~new_P2_R2182_U270;
  assign new_P2_R2182_U273 = ~new_P2_R2182_U37 | ~new_P2_R2182_U8;
  assign new_P2_R2182_U274 = ~new_P2_R2182_U153 | ~new_P2_U2690;
  assign new_P2_R2182_U275 = ~new_P2_R2182_U32 | ~new_P2_R2182_U11;
  assign new_P2_R2182_U276 = ~new_P2_R2182_U152 | ~new_P2_U2691;
  assign new_P2_R2182_U277 = ~new_P2_R2182_U31 | ~new_P2_R2182_U13;
  assign new_P2_R2182_U278 = ~new_P2_R2182_U151 | ~new_P2_U2692;
  assign new_P2_R2182_U279 = ~new_P2_R2182_U121 | ~new_P2_R2182_U47;
  assign new_P2_R2182_U280 = ~new_P2_U2680 | ~new_P2_R2182_U46;
  assign new_P2_R2182_U281 = ~new_P2_R2182_U101;
  assign new_P2_R2182_U282 = ~new_P2_R2182_U281 | ~new_P2_U2701;
  assign new_P2_R2182_U283 = ~new_P2_R2182_U101 | ~new_P2_R2182_U67;
  assign new_P2_R2182_U284 = ~new_P2_R2182_U30 | ~new_P2_R2182_U12;
  assign new_P2_R2182_U285 = ~new_P2_R2182_U150 | ~new_P2_U2693;
  assign new_P2_R2182_U286 = ~new_P2_R2182_U29 | ~new_P2_R2182_U18;
  assign new_P2_R2182_U287 = ~new_P2_R2182_U149 | ~new_P2_U2694;
  assign new_P2_R2182_U288 = ~new_P2_R2182_U28 | ~new_P2_R2182_U17;
  assign new_P2_R2182_U289 = ~new_P2_R2182_U148 | ~new_P2_U2695;
  assign new_P2_R2182_U290 = ~new_P2_R2182_U27 | ~new_P2_R2182_U16;
  assign new_P2_R2182_U291 = ~new_P2_R2182_U147 | ~new_P2_U2696;
  assign new_P2_R2182_U292 = ~new_P2_R2182_U25 | ~new_P2_R2182_U15;
  assign new_P2_R2182_U293 = ~new_P2_R2182_U146 | ~new_P2_U2666;
  assign new_P2_R2182_U294 = ~new_P2_R2182_U26 | ~new_P2_R2182_U14;
  assign new_P2_R2182_U295 = ~new_P2_R2182_U145 | ~new_P2_U2667;
  assign new_P2_R2182_U296 = ~new_P2_R2182_U38 | ~new_P2_R2182_U6;
  assign new_P2_R2182_U297 = ~new_P2_R2182_U144 | ~new_P2_U2668;
  assign new_P2_R2182_U298 = ~new_P2_R2182_U39 | ~new_P2_R2182_U5;
  assign new_P2_R2182_U299 = ~new_P2_R2182_U143 | ~new_P2_U2669;
  assign new_P2_R2182_U300 = ~new_P2_R2182_U33 | ~new_P2_R2182_U4;
  assign new_P2_R2182_U301 = ~new_P2_R2182_U142 | ~new_P2_U2670;
  assign new_P2_R2182_U302 = ~new_P2_R2182_U23 | ~new_P2_R2182_U20;
  assign new_P2_R2182_U303 = ~new_P2_R2182_U141 | ~new_P2_U2671;
  assign new_P2_R2182_U304 = ~new_P2_U2681 | ~new_P2_R2182_U44;
  assign new_P2_R2182_U305 = ~new_P2_U2702 | ~new_P2_R2182_U45;
  assign new_P2_R2167_U6 = ~new_P2_R2167_U38 | ~new_P2_R2167_U42 | ~new_P2_R2167_U41;
  assign new_P2_R2167_U7 = ~new_P2_U2706;
  assign new_P2_R2167_U8 = ~new_P2_U2713;
  assign new_P2_R2167_U9 = ~new_P2_U2712;
  assign new_P2_R2167_U10 = ~new_P2_U2705;
  assign new_P2_R2167_U11 = ~new_P2_U2704;
  assign new_P2_R2167_U12 = ~new_P2_U2711;
  assign new_P2_R2167_U13 = ~new_P2_U2710;
  assign new_P2_R2167_U14 = ~new_P2_U2703;
  assign new_P2_R2167_U15 = ~new_P2_U2361;
  assign new_P2_R2167_U16 = ~new_P2_U2709;
  assign new_P2_R2167_U17 = ~P2_STATE2_REG_0_;
  assign new_P2_R2167_U18 = ~new_P2_U2708;
  assign new_P2_R2167_U19 = ~new_P2_U2714 | ~new_P2_U2715;
  assign new_P2_R2167_U20 = ~new_P2_U2707 | ~new_P2_R2167_U19;
  assign new_P2_R2167_U21 = new_P2_U2714 | new_P2_U2715;
  assign new_P2_R2167_U22 = ~new_P2_U2706 | ~new_P2_R2167_U8;
  assign new_P2_R2167_U23 = ~new_P2_R2167_U22 | ~new_P2_R2167_U21 | ~new_P2_R2167_U20;
  assign new_P2_R2167_U24 = ~new_P2_U2713 | ~new_P2_R2167_U7;
  assign new_P2_R2167_U25 = ~new_P2_U2712 | ~new_P2_R2167_U10;
  assign new_P2_R2167_U26 = ~new_P2_R2167_U23 | ~new_P2_R2167_U24 | ~new_P2_R2167_U25;
  assign new_P2_R2167_U27 = ~new_P2_U2705 | ~new_P2_R2167_U9;
  assign new_P2_R2167_U28 = ~new_P2_U2704 | ~new_P2_R2167_U12;
  assign new_P2_R2167_U29 = ~new_P2_R2167_U26 | ~new_P2_R2167_U27 | ~new_P2_R2167_U28;
  assign new_P2_R2167_U30 = ~new_P2_U2711 | ~new_P2_R2167_U11;
  assign new_P2_R2167_U31 = ~new_P2_U2710 | ~new_P2_R2167_U14;
  assign new_P2_R2167_U32 = ~new_P2_R2167_U31 | ~new_P2_R2167_U30 | ~new_P2_R2167_U29;
  assign new_P2_R2167_U33 = ~new_P2_U2703 | ~new_P2_R2167_U13;
  assign new_P2_R2167_U34 = ~new_P2_U2361 | ~new_P2_R2167_U16;
  assign new_P2_R2167_U35 = ~new_P2_R2167_U34 | ~new_P2_R2167_U33 | ~new_P2_R2167_U32;
  assign new_P2_R2167_U36 = ~new_P2_U2709 | ~new_P2_R2167_U15;
  assign new_P2_R2167_U37 = ~new_P2_R2167_U36 | ~new_P2_R2167_U35;
  assign new_P2_R2167_U38 = ~new_P2_R2167_U37 | ~new_P2_R2167_U40 | ~new_P2_R2167_U39;
  assign new_P2_R2167_U39 = ~new_P2_U2361 | ~new_P2_R2167_U18;
  assign new_P2_R2167_U40 = ~new_P2_U2708 | ~new_P2_R2167_U15;
  assign new_P2_R2167_U41 = ~new_P2_R2167_U18 | ~P2_STATE2_REG_0_ | ~new_P2_U2361;
  assign new_P2_R2167_U42 = ~new_P2_U2708 | ~new_P2_R2167_U17 | ~new_P2_R2167_U15;
  assign new_P2_R2027_U5 = ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_R2027_U6 = ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_R2027_U7 = ~P2_INSTADDRPOINTER_REG_1_ | ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_R2027_U8 = ~P2_INSTADDRPOINTER_REG_2_;
  assign new_P2_R2027_U9 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_R2027_U98;
  assign new_P2_R2027_U10 = ~P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_R2027_U11 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_R2027_U99;
  assign new_P2_R2027_U12 = ~P2_INSTADDRPOINTER_REG_4_;
  assign new_P2_R2027_U13 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_R2027_U100;
  assign new_P2_R2027_U14 = ~P2_INSTADDRPOINTER_REG_5_;
  assign new_P2_R2027_U15 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_R2027_U101;
  assign new_P2_R2027_U16 = ~P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_R2027_U17 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_R2027_U102;
  assign new_P2_R2027_U18 = ~P2_INSTADDRPOINTER_REG_7_;
  assign new_P2_R2027_U19 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_R2027_U103;
  assign new_P2_R2027_U20 = ~P2_INSTADDRPOINTER_REG_8_;
  assign new_P2_R2027_U21 = ~P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_R2027_U22 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_R2027_U104;
  assign new_P2_R2027_U23 = ~new_P2_R2027_U105 | ~P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_R2027_U24 = ~P2_INSTADDRPOINTER_REG_10_;
  assign new_P2_R2027_U25 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_R2027_U106;
  assign new_P2_R2027_U26 = ~P2_INSTADDRPOINTER_REG_11_;
  assign new_P2_R2027_U27 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_R2027_U107;
  assign new_P2_R2027_U28 = ~P2_INSTADDRPOINTER_REG_12_;
  assign new_P2_R2027_U29 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_R2027_U108;
  assign new_P2_R2027_U30 = ~P2_INSTADDRPOINTER_REG_13_;
  assign new_P2_R2027_U31 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_R2027_U109;
  assign new_P2_R2027_U32 = ~P2_INSTADDRPOINTER_REG_14_;
  assign new_P2_R2027_U33 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_R2027_U110;
  assign new_P2_R2027_U34 = ~P2_INSTADDRPOINTER_REG_15_;
  assign new_P2_R2027_U35 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_R2027_U111;
  assign new_P2_R2027_U36 = ~P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_R2027_U37 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_R2027_U112;
  assign new_P2_R2027_U38 = ~P2_INSTADDRPOINTER_REG_17_;
  assign new_P2_R2027_U39 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_R2027_U113;
  assign new_P2_R2027_U40 = ~P2_INSTADDRPOINTER_REG_18_;
  assign new_P2_R2027_U41 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_R2027_U114;
  assign new_P2_R2027_U42 = ~P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_R2027_U43 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_R2027_U115;
  assign new_P2_R2027_U44 = ~P2_INSTADDRPOINTER_REG_20_;
  assign new_P2_R2027_U45 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_R2027_U116;
  assign new_P2_R2027_U46 = ~P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_R2027_U47 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_R2027_U117;
  assign new_P2_R2027_U48 = ~P2_INSTADDRPOINTER_REG_22_;
  assign new_P2_R2027_U49 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_R2027_U118;
  assign new_P2_R2027_U50 = ~P2_INSTADDRPOINTER_REG_23_;
  assign new_P2_R2027_U51 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_R2027_U119;
  assign new_P2_R2027_U52 = ~P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_R2027_U53 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_R2027_U120;
  assign new_P2_R2027_U54 = ~P2_INSTADDRPOINTER_REG_25_;
  assign new_P2_R2027_U55 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_R2027_U121;
  assign new_P2_R2027_U56 = ~P2_INSTADDRPOINTER_REG_26_;
  assign new_P2_R2027_U57 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_R2027_U122;
  assign new_P2_R2027_U58 = ~P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_R2027_U59 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_R2027_U123;
  assign new_P2_R2027_U60 = ~P2_INSTADDRPOINTER_REG_28_;
  assign new_P2_R2027_U61 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_R2027_U124;
  assign new_P2_R2027_U62 = ~P2_INSTADDRPOINTER_REG_29_;
  assign new_P2_R2027_U63 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_R2027_U125;
  assign new_P2_R2027_U64 = ~P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_R2027_U65 = ~new_P2_R2027_U129 | ~new_P2_R2027_U128;
  assign new_P2_R2027_U66 = ~new_P2_R2027_U131 | ~new_P2_R2027_U130;
  assign new_P2_R2027_U67 = ~new_P2_R2027_U133 | ~new_P2_R2027_U132;
  assign new_P2_R2027_U68 = ~new_P2_R2027_U135 | ~new_P2_R2027_U134;
  assign new_P2_R2027_U69 = ~new_P2_R2027_U137 | ~new_P2_R2027_U136;
  assign new_P2_R2027_U70 = ~new_P2_R2027_U139 | ~new_P2_R2027_U138;
  assign new_P2_R2027_U71 = ~new_P2_R2027_U141 | ~new_P2_R2027_U140;
  assign new_P2_R2027_U72 = ~new_P2_R2027_U143 | ~new_P2_R2027_U142;
  assign new_P2_R2027_U73 = ~new_P2_R2027_U145 | ~new_P2_R2027_U144;
  assign new_P2_R2027_U74 = ~new_P2_R2027_U147 | ~new_P2_R2027_U146;
  assign new_P2_R2027_U75 = ~new_P2_R2027_U149 | ~new_P2_R2027_U148;
  assign new_P2_R2027_U76 = ~new_P2_R2027_U151 | ~new_P2_R2027_U150;
  assign new_P2_R2027_U77 = ~new_P2_R2027_U153 | ~new_P2_R2027_U152;
  assign new_P2_R2027_U78 = ~new_P2_R2027_U155 | ~new_P2_R2027_U154;
  assign new_P2_R2027_U79 = ~new_P2_R2027_U157 | ~new_P2_R2027_U156;
  assign new_P2_R2027_U80 = ~new_P2_R2027_U159 | ~new_P2_R2027_U158;
  assign new_P2_R2027_U81 = ~new_P2_R2027_U161 | ~new_P2_R2027_U160;
  assign new_P2_R2027_U82 = ~new_P2_R2027_U163 | ~new_P2_R2027_U162;
  assign new_P2_R2027_U83 = ~new_P2_R2027_U165 | ~new_P2_R2027_U164;
  assign new_P2_R2027_U84 = ~new_P2_R2027_U167 | ~new_P2_R2027_U166;
  assign new_P2_R2027_U85 = ~new_P2_R2027_U169 | ~new_P2_R2027_U168;
  assign new_P2_R2027_U86 = ~new_P2_R2027_U171 | ~new_P2_R2027_U170;
  assign new_P2_R2027_U87 = ~new_P2_R2027_U173 | ~new_P2_R2027_U172;
  assign new_P2_R2027_U88 = ~new_P2_R2027_U175 | ~new_P2_R2027_U174;
  assign new_P2_R2027_U89 = ~new_P2_R2027_U177 | ~new_P2_R2027_U176;
  assign new_P2_R2027_U90 = ~new_P2_R2027_U179 | ~new_P2_R2027_U178;
  assign new_P2_R2027_U91 = ~new_P2_R2027_U181 | ~new_P2_R2027_U180;
  assign new_P2_R2027_U92 = ~new_P2_R2027_U183 | ~new_P2_R2027_U182;
  assign new_P2_R2027_U93 = ~new_P2_R2027_U185 | ~new_P2_R2027_U184;
  assign new_P2_R2027_U94 = ~new_P2_R2027_U187 | ~new_P2_R2027_U186;
  assign new_P2_R2027_U95 = ~new_P2_R2027_U189 | ~new_P2_R2027_U188;
  assign new_P2_R2027_U96 = ~P2_INSTADDRPOINTER_REG_31_;
  assign new_P2_R2027_U97 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_R2027_U126;
  assign new_P2_R2027_U98 = ~new_P2_R2027_U7;
  assign new_P2_R2027_U99 = ~new_P2_R2027_U9;
  assign new_P2_R2027_U100 = ~new_P2_R2027_U11;
  assign new_P2_R2027_U101 = ~new_P2_R2027_U13;
  assign new_P2_R2027_U102 = ~new_P2_R2027_U15;
  assign new_P2_R2027_U103 = ~new_P2_R2027_U17;
  assign new_P2_R2027_U104 = ~new_P2_R2027_U19;
  assign new_P2_R2027_U105 = ~new_P2_R2027_U22;
  assign new_P2_R2027_U106 = ~new_P2_R2027_U23;
  assign new_P2_R2027_U107 = ~new_P2_R2027_U25;
  assign new_P2_R2027_U108 = ~new_P2_R2027_U27;
  assign new_P2_R2027_U109 = ~new_P2_R2027_U29;
  assign new_P2_R2027_U110 = ~new_P2_R2027_U31;
  assign new_P2_R2027_U111 = ~new_P2_R2027_U33;
  assign new_P2_R2027_U112 = ~new_P2_R2027_U35;
  assign new_P2_R2027_U113 = ~new_P2_R2027_U37;
  assign new_P2_R2027_U114 = ~new_P2_R2027_U39;
  assign new_P2_R2027_U115 = ~new_P2_R2027_U41;
  assign new_P2_R2027_U116 = ~new_P2_R2027_U43;
  assign new_P2_R2027_U117 = ~new_P2_R2027_U45;
  assign new_P2_R2027_U118 = ~new_P2_R2027_U47;
  assign new_P2_R2027_U119 = ~new_P2_R2027_U49;
  assign new_P2_R2027_U120 = ~new_P2_R2027_U51;
  assign new_P2_R2027_U121 = ~new_P2_R2027_U53;
  assign new_P2_R2027_U122 = ~new_P2_R2027_U55;
  assign new_P2_R2027_U123 = ~new_P2_R2027_U57;
  assign new_P2_R2027_U124 = ~new_P2_R2027_U59;
  assign new_P2_R2027_U125 = ~new_P2_R2027_U61;
  assign new_P2_R2027_U126 = ~new_P2_R2027_U63;
  assign new_P2_R2027_U127 = ~new_P2_R2027_U97;
  assign new_P2_R2027_U128 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_R2027_U22;
  assign new_P2_R2027_U129 = ~new_P2_R2027_U105 | ~new_P2_R2027_U21;
  assign new_P2_R2027_U130 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_R2027_U19;
  assign new_P2_R2027_U131 = ~new_P2_R2027_U104 | ~new_P2_R2027_U20;
  assign new_P2_R2027_U132 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_R2027_U17;
  assign new_P2_R2027_U133 = ~new_P2_R2027_U103 | ~new_P2_R2027_U18;
  assign new_P2_R2027_U134 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_R2027_U15;
  assign new_P2_R2027_U135 = ~new_P2_R2027_U102 | ~new_P2_R2027_U16;
  assign new_P2_R2027_U136 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_R2027_U13;
  assign new_P2_R2027_U137 = ~new_P2_R2027_U101 | ~new_P2_R2027_U14;
  assign new_P2_R2027_U138 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_R2027_U11;
  assign new_P2_R2027_U139 = ~new_P2_R2027_U100 | ~new_P2_R2027_U12;
  assign new_P2_R2027_U140 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_R2027_U9;
  assign new_P2_R2027_U141 = ~new_P2_R2027_U99 | ~new_P2_R2027_U10;
  assign new_P2_R2027_U142 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_R2027_U97;
  assign new_P2_R2027_U143 = ~new_P2_R2027_U127 | ~new_P2_R2027_U96;
  assign new_P2_R2027_U144 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_R2027_U63;
  assign new_P2_R2027_U145 = ~new_P2_R2027_U126 | ~new_P2_R2027_U64;
  assign new_P2_R2027_U146 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_R2027_U7;
  assign new_P2_R2027_U147 = ~new_P2_R2027_U98 | ~new_P2_R2027_U8;
  assign new_P2_R2027_U148 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_R2027_U61;
  assign new_P2_R2027_U149 = ~new_P2_R2027_U125 | ~new_P2_R2027_U62;
  assign new_P2_R2027_U150 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_R2027_U59;
  assign new_P2_R2027_U151 = ~new_P2_R2027_U124 | ~new_P2_R2027_U60;
  assign new_P2_R2027_U152 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_R2027_U57;
  assign new_P2_R2027_U153 = ~new_P2_R2027_U123 | ~new_P2_R2027_U58;
  assign new_P2_R2027_U154 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_R2027_U55;
  assign new_P2_R2027_U155 = ~new_P2_R2027_U122 | ~new_P2_R2027_U56;
  assign new_P2_R2027_U156 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_R2027_U53;
  assign new_P2_R2027_U157 = ~new_P2_R2027_U121 | ~new_P2_R2027_U54;
  assign new_P2_R2027_U158 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_R2027_U51;
  assign new_P2_R2027_U159 = ~new_P2_R2027_U120 | ~new_P2_R2027_U52;
  assign new_P2_R2027_U160 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_R2027_U49;
  assign new_P2_R2027_U161 = ~new_P2_R2027_U119 | ~new_P2_R2027_U50;
  assign new_P2_R2027_U162 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_R2027_U47;
  assign new_P2_R2027_U163 = ~new_P2_R2027_U118 | ~new_P2_R2027_U48;
  assign new_P2_R2027_U164 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_R2027_U45;
  assign new_P2_R2027_U165 = ~new_P2_R2027_U117 | ~new_P2_R2027_U46;
  assign new_P2_R2027_U166 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_R2027_U43;
  assign new_P2_R2027_U167 = ~new_P2_R2027_U116 | ~new_P2_R2027_U44;
  assign new_P2_R2027_U168 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_R2027_U5;
  assign new_P2_R2027_U169 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_R2027_U6;
  assign new_P2_R2027_U170 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_R2027_U41;
  assign new_P2_R2027_U171 = ~new_P2_R2027_U115 | ~new_P2_R2027_U42;
  assign new_P2_R2027_U172 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_R2027_U39;
  assign new_P2_R2027_U173 = ~new_P2_R2027_U114 | ~new_P2_R2027_U40;
  assign new_P2_R2027_U174 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_R2027_U37;
  assign new_P2_R2027_U175 = ~new_P2_R2027_U113 | ~new_P2_R2027_U38;
  assign new_P2_R2027_U176 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_R2027_U35;
  assign new_P2_R2027_U177 = ~new_P2_R2027_U112 | ~new_P2_R2027_U36;
  assign new_P2_R2027_U178 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_R2027_U33;
  assign new_P2_R2027_U179 = ~new_P2_R2027_U111 | ~new_P2_R2027_U34;
  assign new_P2_R2027_U180 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_R2027_U31;
  assign new_P2_R2027_U181 = ~new_P2_R2027_U110 | ~new_P2_R2027_U32;
  assign new_P2_R2027_U182 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_R2027_U29;
  assign new_P2_R2027_U183 = ~new_P2_R2027_U109 | ~new_P2_R2027_U30;
  assign new_P2_R2027_U184 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_R2027_U27;
  assign new_P2_R2027_U185 = ~new_P2_R2027_U108 | ~new_P2_R2027_U28;
  assign new_P2_R2027_U186 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_R2027_U25;
  assign new_P2_R2027_U187 = ~new_P2_R2027_U107 | ~new_P2_R2027_U26;
  assign new_P2_R2027_U188 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_R2027_U23;
  assign new_P2_R2027_U189 = ~new_P2_R2027_U106 | ~new_P2_R2027_U24;
  assign new_P2_LT_563_1260_U6 = new_P2_LT_563_1260_U7 | new_P2_U3617;
  assign new_P2_LT_563_1260_U7 = ~new_P2_SUB_563_U6 & ~new_P2_SUB_563_U7;
  assign new_P2_R2337_U4 = ~P2_PHYADDRPOINTER_REG_1_;
  assign new_P2_R2337_U5 = ~P2_PHYADDRPOINTER_REG_3_;
  assign new_P2_R2337_U6 = ~P2_PHYADDRPOINTER_REG_2_;
  assign new_P2_R2337_U7 = ~P2_PHYADDRPOINTER_REG_2_ | ~P2_PHYADDRPOINTER_REG_3_ | ~P2_PHYADDRPOINTER_REG_1_;
  assign new_P2_R2337_U8 = ~P2_PHYADDRPOINTER_REG_4_;
  assign new_P2_R2337_U9 = ~P2_PHYADDRPOINTER_REG_4_ | ~new_P2_R2337_U95;
  assign new_P2_R2337_U10 = ~P2_PHYADDRPOINTER_REG_5_;
  assign new_P2_R2337_U11 = ~P2_PHYADDRPOINTER_REG_5_ | ~new_P2_R2337_U96;
  assign new_P2_R2337_U12 = ~P2_PHYADDRPOINTER_REG_6_;
  assign new_P2_R2337_U13 = ~P2_PHYADDRPOINTER_REG_6_ | ~new_P2_R2337_U97;
  assign new_P2_R2337_U14 = ~P2_PHYADDRPOINTER_REG_7_;
  assign new_P2_R2337_U15 = ~P2_PHYADDRPOINTER_REG_7_ | ~new_P2_R2337_U98;
  assign new_P2_R2337_U16 = ~P2_PHYADDRPOINTER_REG_8_;
  assign new_P2_R2337_U17 = ~P2_PHYADDRPOINTER_REG_9_;
  assign new_P2_R2337_U18 = ~P2_PHYADDRPOINTER_REG_8_ | ~new_P2_R2337_U99;
  assign new_P2_R2337_U19 = ~new_P2_R2337_U100 | ~P2_PHYADDRPOINTER_REG_9_;
  assign new_P2_R2337_U20 = ~P2_PHYADDRPOINTER_REG_10_;
  assign new_P2_R2337_U21 = ~P2_PHYADDRPOINTER_REG_10_ | ~new_P2_R2337_U101;
  assign new_P2_R2337_U22 = ~P2_PHYADDRPOINTER_REG_11_;
  assign new_P2_R2337_U23 = ~P2_PHYADDRPOINTER_REG_11_ | ~new_P2_R2337_U102;
  assign new_P2_R2337_U24 = ~P2_PHYADDRPOINTER_REG_12_;
  assign new_P2_R2337_U25 = ~P2_PHYADDRPOINTER_REG_12_ | ~new_P2_R2337_U103;
  assign new_P2_R2337_U26 = ~P2_PHYADDRPOINTER_REG_13_;
  assign new_P2_R2337_U27 = ~P2_PHYADDRPOINTER_REG_13_ | ~new_P2_R2337_U104;
  assign new_P2_R2337_U28 = ~P2_PHYADDRPOINTER_REG_14_;
  assign new_P2_R2337_U29 = ~P2_PHYADDRPOINTER_REG_14_ | ~new_P2_R2337_U105;
  assign new_P2_R2337_U30 = ~P2_PHYADDRPOINTER_REG_15_;
  assign new_P2_R2337_U31 = ~P2_PHYADDRPOINTER_REG_15_ | ~new_P2_R2337_U106;
  assign new_P2_R2337_U32 = ~P2_PHYADDRPOINTER_REG_16_;
  assign new_P2_R2337_U33 = ~P2_PHYADDRPOINTER_REG_16_ | ~new_P2_R2337_U107;
  assign new_P2_R2337_U34 = ~P2_PHYADDRPOINTER_REG_17_;
  assign new_P2_R2337_U35 = ~P2_PHYADDRPOINTER_REG_17_ | ~new_P2_R2337_U108;
  assign new_P2_R2337_U36 = ~P2_PHYADDRPOINTER_REG_18_;
  assign new_P2_R2337_U37 = ~P2_PHYADDRPOINTER_REG_18_ | ~new_P2_R2337_U109;
  assign new_P2_R2337_U38 = ~P2_PHYADDRPOINTER_REG_19_;
  assign new_P2_R2337_U39 = ~P2_PHYADDRPOINTER_REG_19_ | ~new_P2_R2337_U110;
  assign new_P2_R2337_U40 = ~P2_PHYADDRPOINTER_REG_20_;
  assign new_P2_R2337_U41 = ~P2_PHYADDRPOINTER_REG_20_ | ~new_P2_R2337_U111;
  assign new_P2_R2337_U42 = ~P2_PHYADDRPOINTER_REG_21_;
  assign new_P2_R2337_U43 = ~P2_PHYADDRPOINTER_REG_21_ | ~new_P2_R2337_U112;
  assign new_P2_R2337_U44 = ~P2_PHYADDRPOINTER_REG_22_;
  assign new_P2_R2337_U45 = ~P2_PHYADDRPOINTER_REG_22_ | ~new_P2_R2337_U113;
  assign new_P2_R2337_U46 = ~P2_PHYADDRPOINTER_REG_23_;
  assign new_P2_R2337_U47 = ~P2_PHYADDRPOINTER_REG_23_ | ~new_P2_R2337_U114;
  assign new_P2_R2337_U48 = ~P2_PHYADDRPOINTER_REG_24_;
  assign new_P2_R2337_U49 = ~P2_PHYADDRPOINTER_REG_24_ | ~new_P2_R2337_U115;
  assign new_P2_R2337_U50 = ~P2_PHYADDRPOINTER_REG_25_;
  assign new_P2_R2337_U51 = ~P2_PHYADDRPOINTER_REG_25_ | ~new_P2_R2337_U116;
  assign new_P2_R2337_U52 = ~P2_PHYADDRPOINTER_REG_26_;
  assign new_P2_R2337_U53 = ~P2_PHYADDRPOINTER_REG_26_ | ~new_P2_R2337_U117;
  assign new_P2_R2337_U54 = ~P2_PHYADDRPOINTER_REG_27_;
  assign new_P2_R2337_U55 = ~P2_PHYADDRPOINTER_REG_27_ | ~new_P2_R2337_U118;
  assign new_P2_R2337_U56 = ~P2_PHYADDRPOINTER_REG_28_;
  assign new_P2_R2337_U57 = ~P2_PHYADDRPOINTER_REG_28_ | ~new_P2_R2337_U119;
  assign new_P2_R2337_U58 = ~P2_PHYADDRPOINTER_REG_29_;
  assign new_P2_R2337_U59 = ~P2_PHYADDRPOINTER_REG_29_ | ~new_P2_R2337_U120;
  assign new_P2_R2337_U60 = ~P2_PHYADDRPOINTER_REG_30_;
  assign new_P2_R2337_U61 = ~new_P2_R2337_U124 | ~new_P2_R2337_U123;
  assign new_P2_R2337_U62 = ~new_P2_R2337_U126 | ~new_P2_R2337_U125;
  assign new_P2_R2337_U63 = ~new_P2_R2337_U128 | ~new_P2_R2337_U127;
  assign new_P2_R2337_U64 = ~new_P2_R2337_U130 | ~new_P2_R2337_U129;
  assign new_P2_R2337_U65 = ~new_P2_R2337_U132 | ~new_P2_R2337_U131;
  assign new_P2_R2337_U66 = ~new_P2_R2337_U134 | ~new_P2_R2337_U133;
  assign new_P2_R2337_U67 = ~new_P2_R2337_U136 | ~new_P2_R2337_U135;
  assign new_P2_R2337_U68 = ~new_P2_R2337_U138 | ~new_P2_R2337_U137;
  assign new_P2_R2337_U69 = ~new_P2_R2337_U140 | ~new_P2_R2337_U139;
  assign new_P2_R2337_U70 = ~new_P2_R2337_U142 | ~new_P2_R2337_U141;
  assign new_P2_R2337_U71 = ~new_P2_R2337_U144 | ~new_P2_R2337_U143;
  assign new_P2_R2337_U72 = ~new_P2_R2337_U146 | ~new_P2_R2337_U145;
  assign new_P2_R2337_U73 = ~new_P2_R2337_U148 | ~new_P2_R2337_U147;
  assign new_P2_R2337_U74 = ~new_P2_R2337_U150 | ~new_P2_R2337_U149;
  assign new_P2_R2337_U75 = ~new_P2_R2337_U152 | ~new_P2_R2337_U151;
  assign new_P2_R2337_U76 = ~new_P2_R2337_U154 | ~new_P2_R2337_U153;
  assign new_P2_R2337_U77 = ~new_P2_R2337_U156 | ~new_P2_R2337_U155;
  assign new_P2_R2337_U78 = ~new_P2_R2337_U158 | ~new_P2_R2337_U157;
  assign new_P2_R2337_U79 = ~new_P2_R2337_U160 | ~new_P2_R2337_U159;
  assign new_P2_R2337_U80 = ~new_P2_R2337_U162 | ~new_P2_R2337_U161;
  assign new_P2_R2337_U81 = ~new_P2_R2337_U164 | ~new_P2_R2337_U163;
  assign new_P2_R2337_U82 = ~new_P2_R2337_U166 | ~new_P2_R2337_U165;
  assign new_P2_R2337_U83 = ~new_P2_R2337_U168 | ~new_P2_R2337_U167;
  assign new_P2_R2337_U84 = ~new_P2_R2337_U170 | ~new_P2_R2337_U169;
  assign new_P2_R2337_U85 = ~new_P2_R2337_U172 | ~new_P2_R2337_U171;
  assign new_P2_R2337_U86 = ~new_P2_R2337_U174 | ~new_P2_R2337_U173;
  assign new_P2_R2337_U87 = ~new_P2_R2337_U176 | ~new_P2_R2337_U175;
  assign new_P2_R2337_U88 = ~new_P2_R2337_U178 | ~new_P2_R2337_U177;
  assign new_P2_R2337_U89 = ~new_P2_R2337_U180 | ~new_P2_R2337_U179;
  assign new_P2_R2337_U90 = ~new_P2_R2337_U182 | ~new_P2_R2337_U181;
  assign new_P2_R2337_U91 = ~P2_PHYADDRPOINTER_REG_2_ | ~P2_PHYADDRPOINTER_REG_1_;
  assign new_P2_R2337_U92 = ~P2_PHYADDRPOINTER_REG_31_;
  assign new_P2_R2337_U93 = ~P2_PHYADDRPOINTER_REG_30_ | ~new_P2_R2337_U121;
  assign new_P2_R2337_U94 = ~new_P2_R2337_U91;
  assign new_P2_R2337_U95 = ~new_P2_R2337_U7;
  assign new_P2_R2337_U96 = ~new_P2_R2337_U9;
  assign new_P2_R2337_U97 = ~new_P2_R2337_U11;
  assign new_P2_R2337_U98 = ~new_P2_R2337_U13;
  assign new_P2_R2337_U99 = ~new_P2_R2337_U15;
  assign new_P2_R2337_U100 = ~new_P2_R2337_U18;
  assign new_P2_R2337_U101 = ~new_P2_R2337_U19;
  assign new_P2_R2337_U102 = ~new_P2_R2337_U21;
  assign new_P2_R2337_U103 = ~new_P2_R2337_U23;
  assign new_P2_R2337_U104 = ~new_P2_R2337_U25;
  assign new_P2_R2337_U105 = ~new_P2_R2337_U27;
  assign new_P2_R2337_U106 = ~new_P2_R2337_U29;
  assign new_P2_R2337_U107 = ~new_P2_R2337_U31;
  assign new_P2_R2337_U108 = ~new_P2_R2337_U33;
  assign new_P2_R2337_U109 = ~new_P2_R2337_U35;
  assign new_P2_R2337_U110 = ~new_P2_R2337_U37;
  assign new_P2_R2337_U111 = ~new_P2_R2337_U39;
  assign new_P2_R2337_U112 = ~new_P2_R2337_U41;
  assign new_P2_R2337_U113 = ~new_P2_R2337_U43;
  assign new_P2_R2337_U114 = ~new_P2_R2337_U45;
  assign new_P2_R2337_U115 = ~new_P2_R2337_U47;
  assign new_P2_R2337_U116 = ~new_P2_R2337_U49;
  assign new_P2_R2337_U117 = ~new_P2_R2337_U51;
  assign new_P2_R2337_U118 = ~new_P2_R2337_U53;
  assign new_P2_R2337_U119 = ~new_P2_R2337_U55;
  assign new_P2_R2337_U120 = ~new_P2_R2337_U57;
  assign new_P2_R2337_U121 = ~new_P2_R2337_U59;
  assign new_P2_R2337_U122 = ~new_P2_R2337_U93;
  assign new_P2_R2337_U123 = ~P2_PHYADDRPOINTER_REG_9_ | ~new_P2_R2337_U18;
  assign new_P2_R2337_U124 = ~new_P2_R2337_U100 | ~new_P2_R2337_U17;
  assign new_P2_R2337_U125 = ~P2_PHYADDRPOINTER_REG_8_ | ~new_P2_R2337_U15;
  assign new_P2_R2337_U126 = ~new_P2_R2337_U99 | ~new_P2_R2337_U16;
  assign new_P2_R2337_U127 = ~P2_PHYADDRPOINTER_REG_7_ | ~new_P2_R2337_U13;
  assign new_P2_R2337_U128 = ~new_P2_R2337_U98 | ~new_P2_R2337_U14;
  assign new_P2_R2337_U129 = ~P2_PHYADDRPOINTER_REG_6_ | ~new_P2_R2337_U11;
  assign new_P2_R2337_U130 = ~new_P2_R2337_U97 | ~new_P2_R2337_U12;
  assign new_P2_R2337_U131 = ~P2_PHYADDRPOINTER_REG_5_ | ~new_P2_R2337_U9;
  assign new_P2_R2337_U132 = ~new_P2_R2337_U96 | ~new_P2_R2337_U10;
  assign new_P2_R2337_U133 = ~P2_PHYADDRPOINTER_REG_4_ | ~new_P2_R2337_U7;
  assign new_P2_R2337_U134 = ~new_P2_R2337_U95 | ~new_P2_R2337_U8;
  assign new_P2_R2337_U135 = ~P2_PHYADDRPOINTER_REG_3_ | ~new_P2_R2337_U91;
  assign new_P2_R2337_U136 = ~new_P2_R2337_U94 | ~new_P2_R2337_U5;
  assign new_P2_R2337_U137 = ~P2_PHYADDRPOINTER_REG_31_ | ~new_P2_R2337_U93;
  assign new_P2_R2337_U138 = ~new_P2_R2337_U122 | ~new_P2_R2337_U92;
  assign new_P2_R2337_U139 = ~P2_PHYADDRPOINTER_REG_30_ | ~new_P2_R2337_U59;
  assign new_P2_R2337_U140 = ~new_P2_R2337_U121 | ~new_P2_R2337_U60;
  assign new_P2_R2337_U141 = ~P2_PHYADDRPOINTER_REG_2_ | ~new_P2_R2337_U4;
  assign new_P2_R2337_U142 = ~P2_PHYADDRPOINTER_REG_1_ | ~new_P2_R2337_U6;
  assign new_P2_R2337_U143 = ~P2_PHYADDRPOINTER_REG_29_ | ~new_P2_R2337_U57;
  assign new_P2_R2337_U144 = ~new_P2_R2337_U120 | ~new_P2_R2337_U58;
  assign new_P2_R2337_U145 = ~P2_PHYADDRPOINTER_REG_28_ | ~new_P2_R2337_U55;
  assign new_P2_R2337_U146 = ~new_P2_R2337_U119 | ~new_P2_R2337_U56;
  assign new_P2_R2337_U147 = ~P2_PHYADDRPOINTER_REG_27_ | ~new_P2_R2337_U53;
  assign new_P2_R2337_U148 = ~new_P2_R2337_U118 | ~new_P2_R2337_U54;
  assign new_P2_R2337_U149 = ~P2_PHYADDRPOINTER_REG_26_ | ~new_P2_R2337_U51;
  assign new_P2_R2337_U150 = ~new_P2_R2337_U117 | ~new_P2_R2337_U52;
  assign new_P2_R2337_U151 = ~P2_PHYADDRPOINTER_REG_25_ | ~new_P2_R2337_U49;
  assign new_P2_R2337_U152 = ~new_P2_R2337_U116 | ~new_P2_R2337_U50;
  assign new_P2_R2337_U153 = ~P2_PHYADDRPOINTER_REG_24_ | ~new_P2_R2337_U47;
  assign new_P2_R2337_U154 = ~new_P2_R2337_U115 | ~new_P2_R2337_U48;
  assign new_P2_R2337_U155 = ~P2_PHYADDRPOINTER_REG_23_ | ~new_P2_R2337_U45;
  assign new_P2_R2337_U156 = ~new_P2_R2337_U114 | ~new_P2_R2337_U46;
  assign new_P2_R2337_U157 = ~P2_PHYADDRPOINTER_REG_22_ | ~new_P2_R2337_U43;
  assign new_P2_R2337_U158 = ~new_P2_R2337_U113 | ~new_P2_R2337_U44;
  assign new_P2_R2337_U159 = ~P2_PHYADDRPOINTER_REG_21_ | ~new_P2_R2337_U41;
  assign new_P2_R2337_U160 = ~new_P2_R2337_U112 | ~new_P2_R2337_U42;
  assign new_P2_R2337_U161 = ~P2_PHYADDRPOINTER_REG_20_ | ~new_P2_R2337_U39;
  assign new_P2_R2337_U162 = ~new_P2_R2337_U111 | ~new_P2_R2337_U40;
  assign new_P2_R2337_U163 = ~P2_PHYADDRPOINTER_REG_19_ | ~new_P2_R2337_U37;
  assign new_P2_R2337_U164 = ~new_P2_R2337_U110 | ~new_P2_R2337_U38;
  assign new_P2_R2337_U165 = ~P2_PHYADDRPOINTER_REG_18_ | ~new_P2_R2337_U35;
  assign new_P2_R2337_U166 = ~new_P2_R2337_U109 | ~new_P2_R2337_U36;
  assign new_P2_R2337_U167 = ~P2_PHYADDRPOINTER_REG_17_ | ~new_P2_R2337_U33;
  assign new_P2_R2337_U168 = ~new_P2_R2337_U108 | ~new_P2_R2337_U34;
  assign new_P2_R2337_U169 = ~P2_PHYADDRPOINTER_REG_16_ | ~new_P2_R2337_U31;
  assign new_P2_R2337_U170 = ~new_P2_R2337_U107 | ~new_P2_R2337_U32;
  assign new_P2_R2337_U171 = ~P2_PHYADDRPOINTER_REG_15_ | ~new_P2_R2337_U29;
  assign new_P2_R2337_U172 = ~new_P2_R2337_U106 | ~new_P2_R2337_U30;
  assign new_P2_R2337_U173 = ~P2_PHYADDRPOINTER_REG_14_ | ~new_P2_R2337_U27;
  assign new_P2_R2337_U174 = ~new_P2_R2337_U105 | ~new_P2_R2337_U28;
  assign new_P2_R2337_U175 = ~P2_PHYADDRPOINTER_REG_13_ | ~new_P2_R2337_U25;
  assign new_P2_R2337_U176 = ~new_P2_R2337_U104 | ~new_P2_R2337_U26;
  assign new_P2_R2337_U177 = ~P2_PHYADDRPOINTER_REG_12_ | ~new_P2_R2337_U23;
  assign new_P2_R2337_U178 = ~new_P2_R2337_U103 | ~new_P2_R2337_U24;
  assign new_P2_R2337_U179 = ~P2_PHYADDRPOINTER_REG_11_ | ~new_P2_R2337_U21;
  assign new_P2_R2337_U180 = ~new_P2_R2337_U102 | ~new_P2_R2337_U22;
  assign new_P2_R2337_U181 = ~P2_PHYADDRPOINTER_REG_10_ | ~new_P2_R2337_U19;
  assign new_P2_R2337_U182 = ~new_P2_R2337_U101 | ~new_P2_R2337_U20;
  assign new_P2_R2147_U4 = ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_R2147_U5 = ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign new_P2_R2147_U6 = ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign new_P2_R2147_U7 = ~new_P2_R2147_U16 | ~new_P2_R2147_U15;
  assign new_P2_R2147_U8 = ~new_P2_R2147_U18 | ~new_P2_R2147_U17;
  assign new_P2_R2147_U9 = ~new_P2_R2147_U20 | ~new_P2_R2147_U19;
  assign new_P2_R2147_U10 = ~new_P2_U2752;
  assign new_P2_R2147_U11 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~P2_INSTQUEUERD_ADDR_REG_3_ | ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_R2147_U12 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_R2147_U13 = ~new_P2_R2147_U11;
  assign new_P2_R2147_U14 = ~new_P2_R2147_U12;
  assign new_P2_R2147_U15 = ~new_P2_U2752 | ~new_P2_R2147_U11;
  assign new_P2_R2147_U16 = ~new_P2_R2147_U13 | ~new_P2_R2147_U10;
  assign new_P2_R2147_U17 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_R2147_U12;
  assign new_P2_R2147_U18 = ~new_P2_R2147_U14 | ~new_P2_R2147_U5;
  assign new_P2_R2147_U19 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_R2147_U4;
  assign new_P2_R2147_U20 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_R2147_U6;
  assign new_P2_R2219_U6 = new_P2_R2219_U52 & new_P2_R2219_U48;
  assign new_P2_R2219_U7 = new_P2_R2219_U68 & new_P2_R2219_U66;
  assign new_P2_R2219_U8 = ~new_P2_R2219_U45 | ~new_P2_R2219_U69;
  assign new_P2_R2219_U9 = ~new_P2_U4428;
  assign new_P2_R2219_U10 = ~new_P2_U2753;
  assign new_P2_R2219_U11 = ~new_P2_U2761;
  assign new_P2_R2219_U12 = ~new_P2_U2763;
  assign new_P2_R2219_U13 = ~new_P2_U2762;
  assign new_P2_R2219_U14 = ~new_P2_U2756;
  assign new_P2_R2219_U15 = ~new_P2_U2765;
  assign new_P2_R2219_U16 = ~new_P2_U2764;
  assign new_P2_R2219_U17 = ~new_P2_U2755;
  assign new_P2_R2219_U18 = ~new_P2_U2754;
  assign new_P2_R2219_U19 = ~new_P2_R2219_U72 | ~new_P2_R2219_U76;
  assign new_P2_R2219_U20 = ~new_P2_U2760;
  assign new_P2_R2219_U21 = ~new_P2_U2759;
  assign new_P2_R2219_U22 = ~new_P2_U2758;
  assign new_P2_R2219_U23 = ~new_P2_U2757;
  assign new_P2_R2219_U24 = ~new_P2_R2219_U86 | ~new_P2_R2219_U85;
  assign new_P2_R2219_U25 = ~new_P2_R2219_U91 | ~new_P2_R2219_U90;
  assign new_P2_R2219_U26 = ~new_P2_R2219_U96 | ~new_P2_R2219_U95;
  assign new_P2_R2219_U27 = ~new_P2_R2219_U101 | ~new_P2_R2219_U100;
  assign new_P2_R2219_U28 = ~new_P2_R2219_U106 | ~new_P2_R2219_U105;
  assign new_P2_R2219_U29 = ~new_P2_R2219_U111 | ~new_P2_R2219_U110;
  assign new_P2_R2219_U30 = ~new_P2_R2219_U116 | ~new_P2_R2219_U115;
  assign new_P2_R2219_U31 = new_P2_R2219_U6 & new_P2_R2219_U55;
  assign new_P2_R2219_U32 = ~new_P2_R2219_U83 | ~new_P2_R2219_U82;
  assign new_P2_R2219_U33 = ~new_P2_R2219_U88 | ~new_P2_R2219_U87;
  assign new_P2_R2219_U34 = ~new_P2_R2219_U93 | ~new_P2_R2219_U92;
  assign new_P2_R2219_U35 = ~new_P2_R2219_U98 | ~new_P2_R2219_U97;
  assign new_P2_R2219_U36 = ~new_P2_R2219_U103 | ~new_P2_R2219_U102;
  assign new_P2_R2219_U37 = ~new_P2_R2219_U108 | ~new_P2_R2219_U107;
  assign new_P2_R2219_U38 = ~new_P2_R2219_U113 | ~new_P2_R2219_U112;
  assign new_P2_R2219_U39 = ~new_P2_R2219_U64 | ~new_P2_R2219_U63;
  assign new_P2_R2219_U40 = ~new_P2_R2219_U60 | ~new_P2_R2219_U59;
  assign new_P2_R2219_U41 = ~new_P2_R2219_U74 | ~new_P2_R2219_U75 | ~new_P2_R2219_U56;
  assign new_P2_R2219_U42 = ~new_P2_R2219_U19 | ~new_P2_R2219_U71;
  assign new_P2_R2219_U43 = ~new_P2_R2219_U50 | ~new_P2_R2219_U49;
  assign new_P2_R2219_U44 = ~new_P2_R2219_U78 | ~new_P2_R2219_U70;
  assign new_P2_R2219_U45 = ~new_P2_U2765 | ~new_P2_R2219_U23;
  assign new_P2_R2219_U46 = ~new_P2_R2219_U45;
  assign new_P2_R2219_U47 = ~new_P2_U2764 | ~new_P2_R2219_U14;
  assign new_P2_R2219_U48 = ~new_P2_U2763 | ~new_P2_R2219_U17;
  assign new_P2_R2219_U49 = ~new_P2_R2219_U48 | ~new_P2_R2219_U81;
  assign new_P2_R2219_U50 = ~new_P2_U2755 | ~new_P2_R2219_U12;
  assign new_P2_R2219_U51 = ~new_P2_R2219_U43;
  assign new_P2_R2219_U52 = ~new_P2_U2762 | ~new_P2_R2219_U18;
  assign new_P2_R2219_U53 = ~new_P2_U2754 | ~new_P2_R2219_U13;
  assign new_P2_R2219_U54 = ~new_P2_R2219_U42;
  assign new_P2_R2219_U55 = ~new_P2_U2761 | ~new_P2_R2219_U10;
  assign new_P2_R2219_U56 = ~new_P2_U2753 | ~new_P2_R2219_U11;
  assign new_P2_R2219_U57 = ~new_P2_R2219_U41;
  assign new_P2_R2219_U58 = ~new_P2_U2760 | ~new_P2_R2219_U9;
  assign new_P2_R2219_U59 = ~new_P2_R2219_U58 | ~new_P2_R2219_U41;
  assign new_P2_R2219_U60 = ~new_P2_U4428 | ~new_P2_R2219_U20;
  assign new_P2_R2219_U61 = ~new_P2_R2219_U40;
  assign new_P2_R2219_U62 = ~new_P2_U2759 | ~new_P2_R2219_U9;
  assign new_P2_R2219_U63 = ~new_P2_R2219_U62 | ~new_P2_R2219_U40;
  assign new_P2_R2219_U64 = ~new_P2_U4428 | ~new_P2_R2219_U21;
  assign new_P2_R2219_U65 = ~new_P2_R2219_U39;
  assign new_P2_R2219_U66 = ~new_P2_U4428 | ~new_P2_R2219_U22;
  assign new_P2_R2219_U67 = ~new_P2_U2758 | ~new_P2_R2219_U9;
  assign new_P2_R2219_U68 = ~new_P2_R2219_U67 | ~new_P2_R2219_U39;
  assign new_P2_R2219_U69 = ~new_P2_U2757 | ~new_P2_R2219_U15;
  assign new_P2_R2219_U70 = ~new_P2_U2756 | ~new_P2_R2219_U16;
  assign new_P2_R2219_U71 = ~new_P2_R2219_U6 | ~new_P2_R2219_U44;
  assign new_P2_R2219_U72 = ~new_P2_R2219_U53 | ~new_P2_R2219_U50;
  assign new_P2_R2219_U73 = ~new_P2_R2219_U19;
  assign new_P2_R2219_U74 = ~new_P2_R2219_U31 | ~new_P2_R2219_U44;
  assign new_P2_R2219_U75 = ~new_P2_R2219_U73 | ~new_P2_R2219_U55;
  assign new_P2_R2219_U76 = ~new_P2_U2762 | ~new_P2_R2219_U18;
  assign new_P2_R2219_U77 = ~new_P2_U2764 | ~new_P2_R2219_U14;
  assign new_P2_R2219_U78 = ~new_P2_R2219_U47 | ~new_P2_R2219_U45;
  assign new_P2_R2219_U79 = ~new_P2_R2219_U44;
  assign new_P2_R2219_U80 = ~new_P2_R2219_U77 | ~new_P2_R2219_U45;
  assign new_P2_R2219_U81 = ~new_P2_R2219_U80 | ~new_P2_R2219_U70;
  assign new_P2_R2219_U82 = ~new_P2_U2758 | ~new_P2_R2219_U9;
  assign new_P2_R2219_U83 = ~new_P2_U4428 | ~new_P2_R2219_U22;
  assign new_P2_R2219_U84 = ~new_P2_R2219_U32;
  assign new_P2_R2219_U85 = ~new_P2_R2219_U65 | ~new_P2_R2219_U84;
  assign new_P2_R2219_U86 = ~new_P2_R2219_U32 | ~new_P2_R2219_U39;
  assign new_P2_R2219_U87 = ~new_P2_U2759 | ~new_P2_R2219_U9;
  assign new_P2_R2219_U88 = ~new_P2_U4428 | ~new_P2_R2219_U21;
  assign new_P2_R2219_U89 = ~new_P2_R2219_U33;
  assign new_P2_R2219_U90 = ~new_P2_R2219_U61 | ~new_P2_R2219_U89;
  assign new_P2_R2219_U91 = ~new_P2_R2219_U33 | ~new_P2_R2219_U40;
  assign new_P2_R2219_U92 = ~new_P2_U2760 | ~new_P2_R2219_U9;
  assign new_P2_R2219_U93 = ~new_P2_U4428 | ~new_P2_R2219_U20;
  assign new_P2_R2219_U94 = ~new_P2_R2219_U34;
  assign new_P2_R2219_U95 = ~new_P2_R2219_U57 | ~new_P2_R2219_U94;
  assign new_P2_R2219_U96 = ~new_P2_R2219_U34 | ~new_P2_R2219_U41;
  assign new_P2_R2219_U97 = ~new_P2_U2761 | ~new_P2_R2219_U10;
  assign new_P2_R2219_U98 = ~new_P2_U2753 | ~new_P2_R2219_U11;
  assign new_P2_R2219_U99 = ~new_P2_R2219_U35;
  assign new_P2_R2219_U100 = ~new_P2_R2219_U54 | ~new_P2_R2219_U99;
  assign new_P2_R2219_U101 = ~new_P2_R2219_U35 | ~new_P2_R2219_U42;
  assign new_P2_R2219_U102 = ~new_P2_U2762 | ~new_P2_R2219_U18;
  assign new_P2_R2219_U103 = ~new_P2_U2754 | ~new_P2_R2219_U13;
  assign new_P2_R2219_U104 = ~new_P2_R2219_U36;
  assign new_P2_R2219_U105 = ~new_P2_R2219_U51 | ~new_P2_R2219_U104;
  assign new_P2_R2219_U106 = ~new_P2_R2219_U36 | ~new_P2_R2219_U43;
  assign new_P2_R2219_U107 = ~new_P2_U2763 | ~new_P2_R2219_U17;
  assign new_P2_R2219_U108 = ~new_P2_U2755 | ~new_P2_R2219_U12;
  assign new_P2_R2219_U109 = ~new_P2_R2219_U37;
  assign new_P2_R2219_U110 = ~new_P2_R2219_U79 | ~new_P2_R2219_U109;
  assign new_P2_R2219_U111 = ~new_P2_R2219_U37 | ~new_P2_R2219_U44;
  assign new_P2_R2219_U112 = ~new_P2_U2764 | ~new_P2_R2219_U14;
  assign new_P2_R2219_U113 = ~new_P2_U2756 | ~new_P2_R2219_U16;
  assign new_P2_R2219_U114 = ~new_P2_R2219_U38;
  assign new_P2_R2219_U115 = ~new_P2_R2219_U46 | ~new_P2_R2219_U114;
  assign new_P2_R2219_U116 = ~new_P2_R2219_U38 | ~new_P2_R2219_U45;
  assign new_P2_R2243_U6 = ~new_P2_U3687 & ~new_P2_U3684 & ~new_P2_U3686 & ~new_P2_U3685;
  assign new_P2_R2243_U7 = ~new_P2_U3684 & ~new_P2_R2243_U9;
  assign new_P2_R2243_U8 = ~new_P2_R2243_U7 | ~new_P2_R2243_U11;
  assign new_P2_R2243_U9 = ~new_P2_U3685 & ~new_P2_U3686 & ~new_P2_U3684 & ~new_P2_U3689 & ~new_P2_U3687;
  assign new_P2_R2243_U10 = ~new_P2_U3688;
  assign new_P2_R2243_U11 = ~new_P2_R2243_U6 | ~new_P2_R2243_U10;
  assign new_P2_SUB_589_U6 = ~new_P2_U3614;
  assign new_P2_SUB_589_U7 = ~new_P2_U3615;
  assign new_P2_SUB_589_U8 = ~new_P2_U2813;
  assign new_P2_SUB_589_U9 = ~new_P2_U3613;
  assign new_P2_R2096_U4 = new_P2_U2640 & new_P2_R2096_U23;
  assign new_P2_R2096_U5 = new_P2_U2633 & new_P2_R2096_U18;
  assign new_P2_R2096_U6 = new_P2_U2631 & new_P2_R2096_U25;
  assign new_P2_R2096_U7 = new_P2_U2629 & new_P2_R2096_U16;
  assign new_P2_R2096_U8 = new_P2_U2628 & new_P2_R2096_U7;
  assign new_P2_R2096_U9 = new_P2_U2627 & new_P2_R2096_U8;
  assign new_P2_R2096_U10 = new_P2_U2626 & new_P2_R2096_U9;
  assign new_P2_R2096_U11 = new_P2_U2625 & new_P2_R2096_U10;
  assign new_P2_R2096_U12 = new_P2_U2624 & new_P2_R2096_U11;
  assign new_P2_R2096_U13 = new_P2_U2622 & new_P2_R2096_U15;
  assign new_P2_R2096_U14 = new_P2_U2621 & new_P2_R2096_U13;
  assign new_P2_R2096_U15 = new_P2_U2623 & new_P2_R2096_U12;
  assign new_P2_R2096_U16 = new_P2_U2630 & new_P2_R2096_U6;
  assign new_P2_R2096_U17 = new_P2_U2635 & new_P2_R2096_U21;
  assign new_P2_R2096_U18 = new_P2_U2634 & new_P2_R2096_U17;
  assign new_P2_R2096_U19 = new_P2_U2638 & new_P2_R2096_U24;
  assign new_P2_R2096_U20 = new_P2_U2637 & new_P2_R2096_U19;
  assign new_P2_R2096_U21 = new_P2_U2636 & new_P2_R2096_U20;
  assign new_P2_R2096_U22 = new_P2_U2620 & new_P2_R2096_U14;
  assign new_P2_R2096_U23 = new_P2_U2641 & new_P2_R2096_U99;
  assign new_P2_R2096_U24 = new_P2_U2639 & new_P2_R2096_U4;
  assign new_P2_R2096_U25 = new_P2_U2632 & new_P2_R2096_U5;
  assign new_P2_R2096_U26 = ~new_P2_U2631;
  assign new_P2_R2096_U27 = ~new_P2_U2638;
  assign new_P2_R2096_U28 = ~new_P2_U2640;
  assign new_P2_R2096_U29 = ~new_P2_U2618;
  assign new_P2_R2096_U30 = ~new_P2_U2619;
  assign new_P2_R2096_U31 = ~new_P2_U2635;
  assign new_P2_R2096_U32 = ~new_P2_U2636;
  assign new_P2_R2096_U33 = ~new_P2_U2637;
  assign new_P2_R2096_U34 = ~new_P2_U2633;
  assign new_P2_R2096_U35 = ~new_P2_U2634;
  assign new_P2_R2096_U36 = ~new_P2_U2629;
  assign new_P2_R2096_U37 = ~new_P2_U2641;
  assign new_P2_R2096_U38 = ~new_P2_U2622;
  assign new_P2_R2096_U39 = ~new_P2_U2627;
  assign new_P2_R2096_U40 = ~new_P2_U2620;
  assign new_P2_R2096_U41 = ~new_P2_U2621;
  assign new_P2_R2096_U42 = ~new_P2_U2623;
  assign new_P2_R2096_U43 = ~new_P2_U2624;
  assign new_P2_R2096_U44 = ~new_P2_U2625;
  assign new_P2_R2096_U45 = ~new_P2_U2626;
  assign new_P2_R2096_U46 = ~new_P2_U2628;
  assign new_P2_R2096_U47 = ~new_P2_U2630;
  assign new_P2_R2096_U48 = ~new_P2_U2632;
  assign new_P2_R2096_U49 = ~new_P2_U2639;
  assign new_P2_R2096_U50 = new_P2_R2096_U168 & new_P2_R2096_U167;
  assign new_P2_R2096_U51 = ~new_P2_R2096_U114 | ~new_P2_R2096_U170;
  assign new_P2_R2096_U52 = ~new_P2_U2657;
  assign new_P2_R2096_U53 = ~new_P2_U2649;
  assign new_P2_R2096_U54 = ~new_P2_U2648;
  assign new_P2_R2096_U55 = ~new_P2_U2656;
  assign new_P2_R2096_U56 = ~new_P2_U2655;
  assign new_P2_R2096_U57 = ~new_P2_U2647;
  assign new_P2_R2096_U58 = ~new_P2_U2654;
  assign new_P2_R2096_U59 = ~new_P2_U2646;
  assign new_P2_R2096_U60 = ~new_P2_U2653;
  assign new_P2_R2096_U61 = ~new_P2_U2645;
  assign new_P2_R2096_U62 = ~new_P2_U2652;
  assign new_P2_R2096_U63 = ~new_P2_U2644;
  assign new_P2_R2096_U64 = ~new_P2_U2651;
  assign new_P2_R2096_U65 = ~new_P2_U2643;
  assign new_P2_R2096_U66 = ~new_P2_U2650;
  assign new_P2_R2096_U67 = ~new_P2_U2642;
  assign new_P2_R2096_U68 = ~new_P2_R2096_U265 | ~new_P2_R2096_U264;
  assign new_P2_R2096_U69 = ~new_P2_R2096_U172 | ~new_P2_R2096_U171;
  assign new_P2_R2096_U70 = ~new_P2_R2096_U174 | ~new_P2_R2096_U173;
  assign new_P2_R2096_U71 = ~new_P2_R2096_U181 | ~new_P2_R2096_U180;
  assign new_P2_R2096_U72 = ~new_P2_R2096_U188 | ~new_P2_R2096_U187;
  assign new_P2_R2096_U73 = ~new_P2_R2096_U195 | ~new_P2_R2096_U194;
  assign new_P2_R2096_U74 = ~new_P2_R2096_U202 | ~new_P2_R2096_U201;
  assign new_P2_R2096_U75 = ~new_P2_R2096_U209 | ~new_P2_R2096_U208;
  assign new_P2_R2096_U76 = ~new_P2_R2096_U211 | ~new_P2_R2096_U210;
  assign new_P2_R2096_U77 = ~new_P2_R2096_U218 | ~new_P2_R2096_U217;
  assign new_P2_R2096_U78 = ~new_P2_R2096_U220 | ~new_P2_R2096_U219;
  assign new_P2_R2096_U79 = ~new_P2_R2096_U222 | ~new_P2_R2096_U221;
  assign new_P2_R2096_U80 = ~new_P2_R2096_U224 | ~new_P2_R2096_U223;
  assign new_P2_R2096_U81 = ~new_P2_R2096_U226 | ~new_P2_R2096_U225;
  assign new_P2_R2096_U82 = ~new_P2_R2096_U228 | ~new_P2_R2096_U227;
  assign new_P2_R2096_U83 = ~new_P2_R2096_U230 | ~new_P2_R2096_U229;
  assign new_P2_R2096_U84 = ~new_P2_R2096_U232 | ~new_P2_R2096_U231;
  assign new_P2_R2096_U85 = ~new_P2_R2096_U234 | ~new_P2_R2096_U233;
  assign new_P2_R2096_U86 = ~new_P2_R2096_U236 | ~new_P2_R2096_U235;
  assign new_P2_R2096_U87 = ~new_P2_R2096_U238 | ~new_P2_R2096_U237;
  assign new_P2_R2096_U88 = ~new_P2_R2096_U245 | ~new_P2_R2096_U244;
  assign new_P2_R2096_U89 = ~new_P2_R2096_U247 | ~new_P2_R2096_U246;
  assign new_P2_R2096_U90 = ~new_P2_R2096_U249 | ~new_P2_R2096_U248;
  assign new_P2_R2096_U91 = ~new_P2_R2096_U251 | ~new_P2_R2096_U250;
  assign new_P2_R2096_U92 = ~new_P2_R2096_U253 | ~new_P2_R2096_U252;
  assign new_P2_R2096_U93 = ~new_P2_R2096_U255 | ~new_P2_R2096_U254;
  assign new_P2_R2096_U94 = ~new_P2_R2096_U257 | ~new_P2_R2096_U256;
  assign new_P2_R2096_U95 = ~new_P2_R2096_U259 | ~new_P2_R2096_U258;
  assign new_P2_R2096_U96 = ~new_P2_R2096_U261 | ~new_P2_R2096_U260;
  assign new_P2_R2096_U97 = ~new_P2_R2096_U263 | ~new_P2_R2096_U262;
  assign new_P2_R2096_U98 = new_P2_U2619 & new_P2_U2618;
  assign new_P2_R2096_U99 = ~new_P2_R2096_U142 | ~new_P2_R2096_U141;
  assign new_P2_R2096_U100 = new_P2_R2096_U176 & new_P2_R2096_U175;
  assign new_P2_R2096_U101 = ~new_P2_R2096_U138 | ~new_P2_R2096_U137;
  assign new_P2_R2096_U102 = new_P2_R2096_U183 & new_P2_R2096_U182;
  assign new_P2_R2096_U103 = ~new_P2_R2096_U134 | ~new_P2_R2096_U133;
  assign new_P2_R2096_U104 = new_P2_R2096_U190 & new_P2_R2096_U189;
  assign new_P2_R2096_U105 = ~new_P2_R2096_U130 | ~new_P2_R2096_U129;
  assign new_P2_R2096_U106 = new_P2_R2096_U197 & new_P2_R2096_U196;
  assign new_P2_R2096_U107 = ~new_P2_R2096_U126 | ~new_P2_R2096_U125;
  assign new_P2_R2096_U108 = new_P2_R2096_U204 & new_P2_R2096_U203;
  assign new_P2_R2096_U109 = ~new_P2_R2096_U122 | ~new_P2_R2096_U121;
  assign new_P2_R2096_U110 = new_P2_R2096_U213 & new_P2_R2096_U212;
  assign new_P2_R2096_U111 = ~new_P2_R2096_U113 | ~new_P2_R2096_U118;
  assign new_P2_R2096_U112 = ~new_P2_U2649 | ~new_P2_U2657;
  assign new_P2_R2096_U113 = ~new_P2_U2656 | ~new_P2_U2649 | ~new_P2_U2657;
  assign new_P2_R2096_U114 = new_P2_R2096_U243 & new_P2_R2096_U242;
  assign new_P2_R2096_U115 = ~new_P2_R2096_U113;
  assign new_P2_R2096_U116 = ~new_P2_U2649 | ~new_P2_U2657;
  assign new_P2_R2096_U117 = ~new_P2_R2096_U55 | ~new_P2_R2096_U116;
  assign new_P2_R2096_U118 = ~new_P2_U2648 | ~new_P2_R2096_U117;
  assign new_P2_R2096_U119 = ~new_P2_R2096_U111;
  assign new_P2_R2096_U120 = new_P2_U2655 | new_P2_U2647;
  assign new_P2_R2096_U121 = ~new_P2_R2096_U120 | ~new_P2_R2096_U111;
  assign new_P2_R2096_U122 = ~new_P2_U2647 | ~new_P2_U2655;
  assign new_P2_R2096_U123 = ~new_P2_R2096_U109;
  assign new_P2_R2096_U124 = new_P2_U2654 | new_P2_U2646;
  assign new_P2_R2096_U125 = ~new_P2_R2096_U124 | ~new_P2_R2096_U109;
  assign new_P2_R2096_U126 = ~new_P2_U2646 | ~new_P2_U2654;
  assign new_P2_R2096_U127 = ~new_P2_R2096_U107;
  assign new_P2_R2096_U128 = new_P2_U2653 | new_P2_U2645;
  assign new_P2_R2096_U129 = ~new_P2_R2096_U128 | ~new_P2_R2096_U107;
  assign new_P2_R2096_U130 = ~new_P2_U2645 | ~new_P2_U2653;
  assign new_P2_R2096_U131 = ~new_P2_R2096_U105;
  assign new_P2_R2096_U132 = new_P2_U2652 | new_P2_U2644;
  assign new_P2_R2096_U133 = ~new_P2_R2096_U132 | ~new_P2_R2096_U105;
  assign new_P2_R2096_U134 = ~new_P2_U2644 | ~new_P2_U2652;
  assign new_P2_R2096_U135 = ~new_P2_R2096_U103;
  assign new_P2_R2096_U136 = new_P2_U2651 | new_P2_U2643;
  assign new_P2_R2096_U137 = ~new_P2_R2096_U136 | ~new_P2_R2096_U103;
  assign new_P2_R2096_U138 = ~new_P2_U2643 | ~new_P2_U2651;
  assign new_P2_R2096_U139 = ~new_P2_R2096_U101;
  assign new_P2_R2096_U140 = new_P2_U2650 | new_P2_U2642;
  assign new_P2_R2096_U141 = ~new_P2_R2096_U140 | ~new_P2_R2096_U101;
  assign new_P2_R2096_U142 = ~new_P2_U2642 | ~new_P2_U2650;
  assign new_P2_R2096_U143 = ~new_P2_R2096_U99;
  assign new_P2_R2096_U144 = ~new_P2_R2096_U23;
  assign new_P2_R2096_U145 = ~new_P2_R2096_U4;
  assign new_P2_R2096_U146 = ~new_P2_R2096_U24;
  assign new_P2_R2096_U147 = ~new_P2_R2096_U19;
  assign new_P2_R2096_U148 = ~new_P2_R2096_U20;
  assign new_P2_R2096_U149 = ~new_P2_R2096_U21;
  assign new_P2_R2096_U150 = ~new_P2_R2096_U17;
  assign new_P2_R2096_U151 = ~new_P2_R2096_U18;
  assign new_P2_R2096_U152 = ~new_P2_R2096_U5;
  assign new_P2_R2096_U153 = ~new_P2_R2096_U25;
  assign new_P2_R2096_U154 = ~new_P2_R2096_U6;
  assign new_P2_R2096_U155 = ~new_P2_R2096_U16;
  assign new_P2_R2096_U156 = ~new_P2_R2096_U7;
  assign new_P2_R2096_U157 = ~new_P2_R2096_U8;
  assign new_P2_R2096_U158 = ~new_P2_R2096_U9;
  assign new_P2_R2096_U159 = ~new_P2_R2096_U10;
  assign new_P2_R2096_U160 = ~new_P2_R2096_U11;
  assign new_P2_R2096_U161 = ~new_P2_R2096_U12;
  assign new_P2_R2096_U162 = ~new_P2_R2096_U15;
  assign new_P2_R2096_U163 = ~new_P2_R2096_U13;
  assign new_P2_R2096_U164 = ~new_P2_R2096_U14;
  assign new_P2_R2096_U165 = ~new_P2_R2096_U22;
  assign new_P2_R2096_U166 = ~new_P2_U2619 | ~new_P2_R2096_U22;
  assign new_P2_R2096_U167 = ~new_P2_R2096_U29 | ~new_P2_R2096_U166;
  assign new_P2_R2096_U168 = ~new_P2_R2096_U98 | ~new_P2_R2096_U22;
  assign new_P2_R2096_U169 = ~new_P2_R2096_U112;
  assign new_P2_R2096_U170 = ~new_P2_R2096_U241 | ~new_P2_R2096_U55;
  assign new_P2_R2096_U171 = ~new_P2_R2096_U28 | ~new_P2_R2096_U23;
  assign new_P2_R2096_U172 = ~new_P2_R2096_U144 | ~new_P2_U2640;
  assign new_P2_R2096_U173 = ~new_P2_R2096_U37 | ~new_P2_R2096_U99;
  assign new_P2_R2096_U174 = ~new_P2_R2096_U143 | ~new_P2_U2641;
  assign new_P2_R2096_U175 = ~new_P2_U2642 | ~new_P2_R2096_U66;
  assign new_P2_R2096_U176 = ~new_P2_U2650 | ~new_P2_R2096_U67;
  assign new_P2_R2096_U177 = ~new_P2_U2642 | ~new_P2_R2096_U66;
  assign new_P2_R2096_U178 = ~new_P2_U2650 | ~new_P2_R2096_U67;
  assign new_P2_R2096_U179 = ~new_P2_R2096_U178 | ~new_P2_R2096_U177;
  assign new_P2_R2096_U180 = ~new_P2_R2096_U100 | ~new_P2_R2096_U101;
  assign new_P2_R2096_U181 = ~new_P2_R2096_U139 | ~new_P2_R2096_U179;
  assign new_P2_R2096_U182 = ~new_P2_U2643 | ~new_P2_R2096_U64;
  assign new_P2_R2096_U183 = ~new_P2_U2651 | ~new_P2_R2096_U65;
  assign new_P2_R2096_U184 = ~new_P2_U2643 | ~new_P2_R2096_U64;
  assign new_P2_R2096_U185 = ~new_P2_U2651 | ~new_P2_R2096_U65;
  assign new_P2_R2096_U186 = ~new_P2_R2096_U185 | ~new_P2_R2096_U184;
  assign new_P2_R2096_U187 = ~new_P2_R2096_U102 | ~new_P2_R2096_U103;
  assign new_P2_R2096_U188 = ~new_P2_R2096_U135 | ~new_P2_R2096_U186;
  assign new_P2_R2096_U189 = ~new_P2_U2644 | ~new_P2_R2096_U62;
  assign new_P2_R2096_U190 = ~new_P2_U2652 | ~new_P2_R2096_U63;
  assign new_P2_R2096_U191 = ~new_P2_U2644 | ~new_P2_R2096_U62;
  assign new_P2_R2096_U192 = ~new_P2_U2652 | ~new_P2_R2096_U63;
  assign new_P2_R2096_U193 = ~new_P2_R2096_U192 | ~new_P2_R2096_U191;
  assign new_P2_R2096_U194 = ~new_P2_R2096_U104 | ~new_P2_R2096_U105;
  assign new_P2_R2096_U195 = ~new_P2_R2096_U131 | ~new_P2_R2096_U193;
  assign new_P2_R2096_U196 = ~new_P2_U2645 | ~new_P2_R2096_U60;
  assign new_P2_R2096_U197 = ~new_P2_U2653 | ~new_P2_R2096_U61;
  assign new_P2_R2096_U198 = ~new_P2_U2645 | ~new_P2_R2096_U60;
  assign new_P2_R2096_U199 = ~new_P2_U2653 | ~new_P2_R2096_U61;
  assign new_P2_R2096_U200 = ~new_P2_R2096_U199 | ~new_P2_R2096_U198;
  assign new_P2_R2096_U201 = ~new_P2_R2096_U106 | ~new_P2_R2096_U107;
  assign new_P2_R2096_U202 = ~new_P2_R2096_U127 | ~new_P2_R2096_U200;
  assign new_P2_R2096_U203 = ~new_P2_U2646 | ~new_P2_R2096_U58;
  assign new_P2_R2096_U204 = ~new_P2_U2654 | ~new_P2_R2096_U59;
  assign new_P2_R2096_U205 = ~new_P2_U2646 | ~new_P2_R2096_U58;
  assign new_P2_R2096_U206 = ~new_P2_U2654 | ~new_P2_R2096_U59;
  assign new_P2_R2096_U207 = ~new_P2_R2096_U206 | ~new_P2_R2096_U205;
  assign new_P2_R2096_U208 = ~new_P2_R2096_U108 | ~new_P2_R2096_U109;
  assign new_P2_R2096_U209 = ~new_P2_R2096_U123 | ~new_P2_R2096_U207;
  assign new_P2_R2096_U210 = ~new_P2_R2096_U30 | ~new_P2_R2096_U22;
  assign new_P2_R2096_U211 = ~new_P2_U2619 | ~new_P2_R2096_U165;
  assign new_P2_R2096_U212 = ~new_P2_U2647 | ~new_P2_R2096_U56;
  assign new_P2_R2096_U213 = ~new_P2_U2655 | ~new_P2_R2096_U57;
  assign new_P2_R2096_U214 = ~new_P2_U2647 | ~new_P2_R2096_U56;
  assign new_P2_R2096_U215 = ~new_P2_U2655 | ~new_P2_R2096_U57;
  assign new_P2_R2096_U216 = ~new_P2_R2096_U215 | ~new_P2_R2096_U214;
  assign new_P2_R2096_U217 = ~new_P2_R2096_U110 | ~new_P2_R2096_U111;
  assign new_P2_R2096_U218 = ~new_P2_R2096_U119 | ~new_P2_R2096_U216;
  assign new_P2_R2096_U219 = ~new_P2_R2096_U40 | ~new_P2_R2096_U14;
  assign new_P2_R2096_U220 = ~new_P2_R2096_U164 | ~new_P2_U2620;
  assign new_P2_R2096_U221 = ~new_P2_R2096_U41 | ~new_P2_R2096_U13;
  assign new_P2_R2096_U222 = ~new_P2_R2096_U163 | ~new_P2_U2621;
  assign new_P2_R2096_U223 = ~new_P2_R2096_U38 | ~new_P2_R2096_U15;
  assign new_P2_R2096_U224 = ~new_P2_R2096_U162 | ~new_P2_U2622;
  assign new_P2_R2096_U225 = ~new_P2_R2096_U42 | ~new_P2_R2096_U12;
  assign new_P2_R2096_U226 = ~new_P2_R2096_U161 | ~new_P2_U2623;
  assign new_P2_R2096_U227 = ~new_P2_R2096_U43 | ~new_P2_R2096_U11;
  assign new_P2_R2096_U228 = ~new_P2_R2096_U160 | ~new_P2_U2624;
  assign new_P2_R2096_U229 = ~new_P2_R2096_U44 | ~new_P2_R2096_U10;
  assign new_P2_R2096_U230 = ~new_P2_R2096_U159 | ~new_P2_U2625;
  assign new_P2_R2096_U231 = ~new_P2_R2096_U45 | ~new_P2_R2096_U9;
  assign new_P2_R2096_U232 = ~new_P2_R2096_U158 | ~new_P2_U2626;
  assign new_P2_R2096_U233 = ~new_P2_R2096_U39 | ~new_P2_R2096_U8;
  assign new_P2_R2096_U234 = ~new_P2_R2096_U157 | ~new_P2_U2627;
  assign new_P2_R2096_U235 = ~new_P2_R2096_U46 | ~new_P2_R2096_U7;
  assign new_P2_R2096_U236 = ~new_P2_R2096_U156 | ~new_P2_U2628;
  assign new_P2_R2096_U237 = ~new_P2_R2096_U36 | ~new_P2_R2096_U16;
  assign new_P2_R2096_U238 = ~new_P2_R2096_U155 | ~new_P2_U2629;
  assign new_P2_R2096_U239 = ~new_P2_U2648 | ~new_P2_R2096_U112;
  assign new_P2_R2096_U240 = ~new_P2_R2096_U169 | ~new_P2_R2096_U54;
  assign new_P2_R2096_U241 = ~new_P2_R2096_U240 | ~new_P2_R2096_U239;
  assign new_P2_R2096_U242 = ~new_P2_R2096_U54 | ~new_P2_U2656 | ~new_P2_R2096_U116;
  assign new_P2_R2096_U243 = ~new_P2_R2096_U115 | ~new_P2_U2648;
  assign new_P2_R2096_U244 = ~new_P2_R2096_U47 | ~new_P2_R2096_U6;
  assign new_P2_R2096_U245 = ~new_P2_R2096_U154 | ~new_P2_U2630;
  assign new_P2_R2096_U246 = ~new_P2_R2096_U26 | ~new_P2_R2096_U25;
  assign new_P2_R2096_U247 = ~new_P2_R2096_U153 | ~new_P2_U2631;
  assign new_P2_R2096_U248 = ~new_P2_R2096_U48 | ~new_P2_R2096_U5;
  assign new_P2_R2096_U249 = ~new_P2_R2096_U152 | ~new_P2_U2632;
  assign new_P2_R2096_U250 = ~new_P2_R2096_U34 | ~new_P2_R2096_U18;
  assign new_P2_R2096_U251 = ~new_P2_R2096_U151 | ~new_P2_U2633;
  assign new_P2_R2096_U252 = ~new_P2_R2096_U35 | ~new_P2_R2096_U17;
  assign new_P2_R2096_U253 = ~new_P2_R2096_U150 | ~new_P2_U2634;
  assign new_P2_R2096_U254 = ~new_P2_R2096_U31 | ~new_P2_R2096_U21;
  assign new_P2_R2096_U255 = ~new_P2_R2096_U149 | ~new_P2_U2635;
  assign new_P2_R2096_U256 = ~new_P2_R2096_U32 | ~new_P2_R2096_U20;
  assign new_P2_R2096_U257 = ~new_P2_R2096_U148 | ~new_P2_U2636;
  assign new_P2_R2096_U258 = ~new_P2_R2096_U33 | ~new_P2_R2096_U19;
  assign new_P2_R2096_U259 = ~new_P2_R2096_U147 | ~new_P2_U2637;
  assign new_P2_R2096_U260 = ~new_P2_R2096_U27 | ~new_P2_R2096_U24;
  assign new_P2_R2096_U261 = ~new_P2_R2096_U146 | ~new_P2_U2638;
  assign new_P2_R2096_U262 = ~new_P2_R2096_U49 | ~new_P2_R2096_U4;
  assign new_P2_R2096_U263 = ~new_P2_R2096_U145 | ~new_P2_U2639;
  assign new_P2_R2096_U264 = ~new_P2_U2649 | ~new_P2_R2096_U52;
  assign new_P2_R2096_U265 = ~new_P2_U2657 | ~new_P2_R2096_U53;
  assign new_P2_GTE_370_U6 = ~new_P2_R2219_U25 & ~new_P2_GTE_370_U8;
  assign new_P2_GTE_370_U7 = new_P2_R2219_U29 & new_P2_GTE_370_U9;
  assign new_P2_GTE_370_U8 = ~new_P2_GTE_370_U7 & ~new_P2_R2219_U28 & ~new_P2_R2219_U26 & ~new_P2_R2219_U27;
  assign new_P2_GTE_370_U9 = new_P2_R2219_U8 | new_P2_R2219_U30;
  assign new_P2_LT_563_U6 = new_P2_LT_563_U27 & new_P2_LT_563_U26;
  assign new_P2_LT_563_U7 = ~new_P2_U3620;
  assign new_P2_LT_563_U8 = ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_LT_563_U9 = ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P2_LT_563_U10 = ~new_P2_U3619;
  assign new_P2_LT_563_U11 = ~new_P2_U3618;
  assign new_P2_LT_563_U12 = ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_LT_563_U13 = ~P2_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P2_LT_563_U14 = ~new_P2_U3617;
  assign new_P2_LT_563_U15 = ~new_P2_U3621;
  assign new_P2_LT_563_U16 = ~new_P2_U3620 | ~new_P2_LT_563_U8;
  assign new_P2_LT_563_U17 = ~new_P2_LT_563_U16 | ~P2_INSTQUEUEWR_ADDR_REG_0_ | ~new_P2_LT_563_U15;
  assign new_P2_LT_563_U18 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_LT_563_U7;
  assign new_P2_LT_563_U19 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_LT_563_U10;
  assign new_P2_LT_563_U20 = ~new_P2_LT_563_U17 | ~new_P2_LT_563_U18 | ~new_P2_LT_563_U19;
  assign new_P2_LT_563_U21 = ~new_P2_U3619 | ~new_P2_LT_563_U9;
  assign new_P2_LT_563_U22 = ~new_P2_U3618 | ~new_P2_LT_563_U12;
  assign new_P2_LT_563_U23 = ~new_P2_LT_563_U20 | ~new_P2_LT_563_U21 | ~new_P2_LT_563_U22;
  assign new_P2_LT_563_U24 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_LT_563_U11;
  assign new_P2_LT_563_U25 = ~P2_INSTQUEUEWR_ADDR_REG_4_ | ~new_P2_LT_563_U14;
  assign new_P2_LT_563_U26 = ~new_P2_LT_563_U23 | ~new_P2_LT_563_U24 | ~new_P2_LT_563_U25;
  assign new_P2_LT_563_U27 = ~new_P2_U3617 | ~new_P2_LT_563_U13;
  assign new_P2_R2256_U4 = ~new_P2_R2256_U31 | ~new_P2_R2256_U46;
  assign new_P2_R2256_U5 = new_P2_R2256_U23 & new_P2_R2256_U43;
  assign new_P2_R2256_U6 = ~new_P2_U3629;
  assign new_P2_R2256_U7 = ~new_P2_U3628;
  assign new_P2_R2256_U8 = ~new_P2_U3627;
  assign new_P2_R2256_U9 = ~new_P2_U3626;
  assign new_P2_R2256_U10 = ~new_P2_U3626 | ~new_P2_R2256_U25;
  assign new_P2_R2256_U11 = ~new_P2_U3625;
  assign new_P2_R2256_U12 = ~new_P2_U3625 | ~new_P2_R2256_U41;
  assign new_P2_R2256_U13 = ~new_P2_U3624;
  assign new_P2_R2256_U14 = ~new_P2_U3624 | ~new_P2_R2256_U42;
  assign new_P2_R2256_U15 = ~new_P2_U3622;
  assign new_P2_R2256_U16 = ~new_P2_U3623;
  assign new_P2_R2256_U17 = ~new_P2_R2256_U48 | ~new_P2_R2256_U47;
  assign new_P2_R2256_U18 = ~new_P2_R2256_U50 | ~new_P2_R2256_U49;
  assign new_P2_R2256_U19 = ~new_P2_R2256_U52 | ~new_P2_R2256_U51;
  assign new_P2_R2256_U20 = ~new_P2_R2256_U54 | ~new_P2_R2256_U53;
  assign new_P2_R2256_U21 = ~new_P2_R2256_U70 | ~new_P2_R2256_U69;
  assign new_P2_R2256_U22 = ~new_P2_R2256_U63 | ~new_P2_R2256_U62;
  assign new_P2_R2256_U23 = new_P2_U3622 & new_P2_U3623;
  assign new_P2_R2256_U24 = ~new_P2_U3623 | ~new_P2_R2256_U43;
  assign new_P2_R2256_U25 = ~new_P2_R2256_U39 | ~new_P2_R2256_U38;
  assign new_P2_R2256_U26 = new_P2_R2256_U56 & new_P2_R2256_U55;
  assign new_P2_R2256_U27 = new_P2_R2256_U58 & new_P2_R2256_U57;
  assign new_P2_R2256_U28 = ~new_P2_R2256_U30 | ~new_P2_R2256_U35;
  assign new_P2_R2256_U29 = ~new_P2_U7873 | ~new_P2_U3629;
  assign new_P2_R2256_U30 = ~new_P2_U3628 | ~new_P2_U7873 | ~new_P2_U3629;
  assign new_P2_R2256_U31 = new_P2_R2256_U68 & new_P2_R2256_U67;
  assign new_P2_R2256_U32 = ~new_P2_R2256_U30;
  assign new_P2_R2256_U33 = ~new_P2_U7873 | ~new_P2_U3629;
  assign new_P2_R2256_U34 = ~new_P2_R2256_U7 | ~new_P2_R2256_U33;
  assign new_P2_R2256_U35 = ~new_P2_U2616 | ~new_P2_R2256_U34;
  assign new_P2_R2256_U36 = ~new_P2_R2256_U28;
  assign new_P2_R2256_U37 = new_P2_U3627 | new_P2_U7873;
  assign new_P2_R2256_U38 = ~new_P2_R2256_U37 | ~new_P2_R2256_U28;
  assign new_P2_R2256_U39 = ~new_P2_U7873 | ~new_P2_U3627;
  assign new_P2_R2256_U40 = ~new_P2_R2256_U25;
  assign new_P2_R2256_U41 = ~new_P2_R2256_U10;
  assign new_P2_R2256_U42 = ~new_P2_R2256_U12;
  assign new_P2_R2256_U43 = ~new_P2_R2256_U14;
  assign new_P2_R2256_U44 = ~new_P2_R2256_U24;
  assign new_P2_R2256_U45 = ~new_P2_R2256_U29;
  assign new_P2_R2256_U46 = ~new_P2_R2256_U66 | ~new_P2_R2256_U7;
  assign new_P2_R2256_U47 = ~new_P2_U3622 | ~new_P2_R2256_U24;
  assign new_P2_R2256_U48 = ~new_P2_R2256_U44 | ~new_P2_R2256_U15;
  assign new_P2_R2256_U49 = ~new_P2_U3623 | ~new_P2_R2256_U14;
  assign new_P2_R2256_U50 = ~new_P2_R2256_U43 | ~new_P2_R2256_U16;
  assign new_P2_R2256_U51 = ~new_P2_U3624 | ~new_P2_R2256_U12;
  assign new_P2_R2256_U52 = ~new_P2_R2256_U42 | ~new_P2_R2256_U13;
  assign new_P2_R2256_U53 = ~new_P2_U3625 | ~new_P2_R2256_U10;
  assign new_P2_R2256_U54 = ~new_P2_R2256_U41 | ~new_P2_R2256_U11;
  assign new_P2_R2256_U55 = ~new_P2_U3626 | ~new_P2_R2256_U25;
  assign new_P2_R2256_U56 = ~new_P2_R2256_U40 | ~new_P2_R2256_U9;
  assign new_P2_R2256_U57 = ~new_P2_U7873 | ~new_P2_R2256_U8;
  assign new_P2_R2256_U58 = ~new_P2_U3627 | ~new_P2_U2616;
  assign new_P2_R2256_U59 = ~new_P2_U7873 | ~new_P2_R2256_U8;
  assign new_P2_R2256_U60 = ~new_P2_U3627 | ~new_P2_U2616;
  assign new_P2_R2256_U61 = ~new_P2_R2256_U60 | ~new_P2_R2256_U59;
  assign new_P2_R2256_U62 = ~new_P2_R2256_U27 | ~new_P2_R2256_U28;
  assign new_P2_R2256_U63 = ~new_P2_R2256_U36 | ~new_P2_R2256_U61;
  assign new_P2_R2256_U64 = ~new_P2_U2616 | ~new_P2_R2256_U29;
  assign new_P2_R2256_U65 = ~new_P2_R2256_U45 | ~new_P2_U7873;
  assign new_P2_R2256_U66 = ~new_P2_R2256_U65 | ~new_P2_R2256_U64;
  assign new_P2_R2256_U67 = ~new_P2_U7873 | ~new_P2_U3628 | ~new_P2_R2256_U33;
  assign new_P2_R2256_U68 = ~new_P2_R2256_U32 | ~new_P2_U2616;
  assign new_P2_R2256_U69 = ~new_P2_U7873 | ~new_P2_R2256_U6;
  assign new_P2_R2256_U70 = ~new_P2_U3629 | ~new_P2_U2616;
  assign new_P2_R2238_U6 = ~new_P2_R2238_U45 | ~new_P2_R2238_U44;
  assign new_P2_R2238_U7 = ~new_P2_R2238_U9 | ~new_P2_R2238_U46;
  assign new_P2_R2238_U8 = ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign new_P2_R2238_U9 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_R2238_U18;
  assign new_P2_R2238_U10 = ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_R2238_U11 = ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign new_P2_R2238_U12 = ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P2_R2238_U13 = ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign new_P2_R2238_U14 = ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_R2238_U15 = ~P2_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P2_R2238_U16 = ~new_P2_R2238_U41 | ~new_P2_R2238_U40;
  assign new_P2_R2238_U17 = ~P2_INSTQUEUERD_ADDR_REG_4_;
  assign new_P2_R2238_U18 = ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P2_R2238_U19 = ~new_P2_R2238_U51 | ~new_P2_R2238_U50;
  assign new_P2_R2238_U20 = ~new_P2_R2238_U56 | ~new_P2_R2238_U55;
  assign new_P2_R2238_U21 = ~new_P2_R2238_U61 | ~new_P2_R2238_U60;
  assign new_P2_R2238_U22 = ~new_P2_R2238_U66 | ~new_P2_R2238_U65;
  assign new_P2_R2238_U23 = ~new_P2_R2238_U48 | ~new_P2_R2238_U47;
  assign new_P2_R2238_U24 = ~new_P2_R2238_U53 | ~new_P2_R2238_U52;
  assign new_P2_R2238_U25 = ~new_P2_R2238_U58 | ~new_P2_R2238_U57;
  assign new_P2_R2238_U26 = ~new_P2_R2238_U63 | ~new_P2_R2238_U62;
  assign new_P2_R2238_U27 = ~new_P2_R2238_U37 | ~new_P2_R2238_U36;
  assign new_P2_R2238_U28 = ~new_P2_R2238_U33 | ~new_P2_R2238_U32;
  assign new_P2_R2238_U29 = ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_R2238_U30 = ~new_P2_R2238_U9;
  assign new_P2_R2238_U31 = ~new_P2_R2238_U30 | ~new_P2_R2238_U10;
  assign new_P2_R2238_U32 = ~new_P2_R2238_U31 | ~new_P2_R2238_U29;
  assign new_P2_R2238_U33 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_R2238_U9;
  assign new_P2_R2238_U34 = ~new_P2_R2238_U28;
  assign new_P2_R2238_U35 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_R2238_U12;
  assign new_P2_R2238_U36 = ~new_P2_R2238_U35 | ~new_P2_R2238_U28;
  assign new_P2_R2238_U37 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_R2238_U11;
  assign new_P2_R2238_U38 = ~new_P2_R2238_U27;
  assign new_P2_R2238_U39 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_R2238_U14;
  assign new_P2_R2238_U40 = ~new_P2_R2238_U39 | ~new_P2_R2238_U27;
  assign new_P2_R2238_U41 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_R2238_U13;
  assign new_P2_R2238_U42 = ~new_P2_R2238_U16;
  assign new_P2_R2238_U43 = ~P2_INSTQUEUEWR_ADDR_REG_4_ | ~new_P2_R2238_U17;
  assign new_P2_R2238_U44 = ~new_P2_R2238_U42 | ~new_P2_R2238_U43;
  assign new_P2_R2238_U45 = ~P2_INSTQUEUERD_ADDR_REG_4_ | ~new_P2_R2238_U15;
  assign new_P2_R2238_U46 = ~P2_INSTQUEUEWR_ADDR_REG_0_ | ~new_P2_R2238_U8;
  assign new_P2_R2238_U47 = ~P2_INSTQUEUERD_ADDR_REG_4_ | ~new_P2_R2238_U15;
  assign new_P2_R2238_U48 = ~P2_INSTQUEUEWR_ADDR_REG_4_ | ~new_P2_R2238_U17;
  assign new_P2_R2238_U49 = ~new_P2_R2238_U23;
  assign new_P2_R2238_U50 = ~new_P2_R2238_U49 | ~new_P2_R2238_U42;
  assign new_P2_R2238_U51 = ~new_P2_R2238_U23 | ~new_P2_R2238_U16;
  assign new_P2_R2238_U52 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_R2238_U14;
  assign new_P2_R2238_U53 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_R2238_U13;
  assign new_P2_R2238_U54 = ~new_P2_R2238_U24;
  assign new_P2_R2238_U55 = ~new_P2_R2238_U38 | ~new_P2_R2238_U54;
  assign new_P2_R2238_U56 = ~new_P2_R2238_U24 | ~new_P2_R2238_U27;
  assign new_P2_R2238_U57 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_R2238_U12;
  assign new_P2_R2238_U58 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_R2238_U11;
  assign new_P2_R2238_U59 = ~new_P2_R2238_U25;
  assign new_P2_R2238_U60 = ~new_P2_R2238_U34 | ~new_P2_R2238_U59;
  assign new_P2_R2238_U61 = ~new_P2_R2238_U25 | ~new_P2_R2238_U28;
  assign new_P2_R2238_U62 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_R2238_U10;
  assign new_P2_R2238_U63 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_R2238_U29;
  assign new_P2_R2238_U64 = ~new_P2_R2238_U26;
  assign new_P2_R2238_U65 = ~new_P2_R2238_U64 | ~new_P2_R2238_U30;
  assign new_P2_R2238_U66 = ~new_P2_R2238_U26 | ~new_P2_R2238_U9;
  assign new_P2_R1957_U6 = new_P2_R1957_U126 & new_P2_R1957_U27;
  assign new_P2_R1957_U7 = new_P2_R1957_U124 & new_P2_R1957_U28;
  assign new_P2_R1957_U8 = new_P2_R1957_U122 & new_P2_R1957_U29;
  assign new_P2_R1957_U9 = new_P2_R1957_U120 & new_P2_R1957_U30;
  assign new_P2_R1957_U10 = new_P2_R1957_U118 & new_P2_R1957_U31;
  assign new_P2_R1957_U11 = new_P2_R1957_U116 & new_P2_R1957_U32;
  assign new_P2_R1957_U12 = new_P2_R1957_U114 & new_P2_R1957_U33;
  assign new_P2_R1957_U13 = new_P2_R1957_U112 & new_P2_R1957_U34;
  assign new_P2_R1957_U14 = new_P2_R1957_U110 & new_P2_R1957_U35;
  assign new_P2_R1957_U15 = new_P2_R1957_U108 & new_P2_R1957_U36;
  assign new_P2_R1957_U16 = new_P2_R1957_U106 & new_P2_R1957_U37;
  assign new_P2_R1957_U17 = new_P2_R1957_U105 & new_P2_R1957_U21;
  assign new_P2_R1957_U18 = new_P2_R1957_U92 & new_P2_R1957_U22;
  assign new_P2_R1957_U19 = new_P2_R1957_U90 & new_P2_R1957_U23;
  assign new_P2_R1957_U20 = new_P2_R1957_U88 & new_P2_R1957_U24;
  assign new_P2_R1957_U21 = new_P2_U3671 | new_P2_U3682 | new_P2_U3683;
  assign new_P2_R1957_U22 = ~new_P2_R1957_U51 | ~new_P2_R1957_U83;
  assign new_P2_R1957_U23 = ~new_P2_R1957_U26 | ~new_P2_R1957_U84 | ~new_P2_R1957_U56;
  assign new_P2_R1957_U24 = ~new_P2_R1957_U25 | ~new_P2_R1957_U85 | ~new_P2_R1957_U54;
  assign new_P2_R1957_U25 = ~new_P2_U3654;
  assign new_P2_R1957_U26 = ~new_P2_U3656;
  assign new_P2_R1957_U27 = ~new_P2_R1957_U48 | ~new_P2_R1957_U52 | ~new_P2_R1957_U86;
  assign new_P2_R1957_U28 = ~new_P2_R1957_U47 | ~new_P2_R1957_U93 | ~new_P2_R1957_U81;
  assign new_P2_R1957_U29 = ~new_P2_R1957_U46 | ~new_P2_R1957_U94 | ~new_P2_R1957_U79;
  assign new_P2_R1957_U30 = ~new_P2_R1957_U45 | ~new_P2_R1957_U95 | ~new_P2_R1957_U77;
  assign new_P2_R1957_U31 = ~new_P2_R1957_U44 | ~new_P2_R1957_U96 | ~new_P2_R1957_U75;
  assign new_P2_R1957_U32 = ~new_P2_R1957_U43 | ~new_P2_R1957_U97 | ~new_P2_R1957_U73;
  assign new_P2_R1957_U33 = ~new_P2_R1957_U42 | ~new_P2_R1957_U98 | ~new_P2_R1957_U69;
  assign new_P2_R1957_U34 = ~new_P2_R1957_U41 | ~new_P2_R1957_U99 | ~new_P2_R1957_U67;
  assign new_P2_R1957_U35 = ~new_P2_R1957_U40 | ~new_P2_R1957_U100 | ~new_P2_R1957_U65;
  assign new_P2_R1957_U36 = ~new_P2_R1957_U39 | ~new_P2_R1957_U101 | ~new_P2_R1957_U63;
  assign new_P2_R1957_U37 = ~new_P2_R1957_U102 | ~new_P2_R1957_U38;
  assign new_P2_R1957_U38 = ~new_P2_U3661;
  assign new_P2_R1957_U39 = ~new_P2_U3662;
  assign new_P2_R1957_U40 = ~new_P2_U3664;
  assign new_P2_R1957_U41 = ~new_P2_U3666;
  assign new_P2_R1957_U42 = ~new_P2_U3668;
  assign new_P2_R1957_U43 = ~new_P2_U3670;
  assign new_P2_R1957_U44 = ~new_P2_U3673;
  assign new_P2_R1957_U45 = ~new_P2_U3675;
  assign new_P2_R1957_U46 = ~new_P2_U3677;
  assign new_P2_R1957_U47 = ~new_P2_U3679;
  assign new_P2_R1957_U48 = ~new_P2_U3681;
  assign new_P2_R1957_U49 = ~new_P2_R1957_U149 | ~new_P2_R1957_U148;
  assign new_P2_R1957_U50 = ~new_P2_R1957_U137 | ~new_P2_R1957_U136;
  assign new_P2_R1957_U51 = ~new_P2_U3660 & ~new_P2_U3658;
  assign new_P2_R1957_U52 = ~new_P2_U3653;
  assign new_P2_R1957_U53 = new_P2_R1957_U129 & new_P2_R1957_U128;
  assign new_P2_R1957_U54 = ~new_P2_U3655;
  assign new_P2_R1957_U55 = new_P2_R1957_U131 & new_P2_R1957_U130;
  assign new_P2_R1957_U56 = ~new_P2_U3657;
  assign new_P2_R1957_U57 = new_P2_R1957_U133 & new_P2_R1957_U132;
  assign new_P2_R1957_U58 = ~new_P2_U3660;
  assign new_P2_R1957_U59 = new_P2_R1957_U135 & new_P2_R1957_U134;
  assign new_P2_R1957_U60 = ~new_P2_U3647;
  assign new_P2_R1957_U61 = ~new_P2_U3659;
  assign new_P2_R1957_U62 = new_P2_R1957_U139 & new_P2_R1957_U138;
  assign new_P2_R1957_U63 = ~new_P2_U3663;
  assign new_P2_R1957_U64 = new_P2_R1957_U141 & new_P2_R1957_U140;
  assign new_P2_R1957_U65 = ~new_P2_U3665;
  assign new_P2_R1957_U66 = new_P2_R1957_U143 & new_P2_R1957_U142;
  assign new_P2_R1957_U67 = ~new_P2_U3667;
  assign new_P2_R1957_U68 = new_P2_R1957_U145 & new_P2_R1957_U144;
  assign new_P2_R1957_U69 = ~new_P2_U3669;
  assign new_P2_R1957_U70 = new_P2_R1957_U147 & new_P2_R1957_U146;
  assign new_P2_R1957_U71 = ~new_P2_U3682;
  assign new_P2_R1957_U72 = ~new_P2_U3683;
  assign new_P2_R1957_U73 = ~new_P2_U3672;
  assign new_P2_R1957_U74 = new_P2_R1957_U151 & new_P2_R1957_U150;
  assign new_P2_R1957_U75 = ~new_P2_U3674;
  assign new_P2_R1957_U76 = new_P2_R1957_U153 & new_P2_R1957_U152;
  assign new_P2_R1957_U77 = ~new_P2_U3676;
  assign new_P2_R1957_U78 = new_P2_R1957_U155 & new_P2_R1957_U154;
  assign new_P2_R1957_U79 = ~new_P2_U3678;
  assign new_P2_R1957_U80 = new_P2_R1957_U157 & new_P2_R1957_U156;
  assign new_P2_R1957_U81 = ~new_P2_U3680;
  assign new_P2_R1957_U82 = new_P2_R1957_U159 & new_P2_R1957_U158;
  assign new_P2_R1957_U83 = ~new_P2_R1957_U21;
  assign new_P2_R1957_U84 = ~new_P2_R1957_U22;
  assign new_P2_R1957_U85 = ~new_P2_R1957_U23;
  assign new_P2_R1957_U86 = ~new_P2_R1957_U24;
  assign new_P2_R1957_U87 = ~new_P2_R1957_U85 | ~new_P2_R1957_U54;
  assign new_P2_R1957_U88 = ~new_P2_U3654 | ~new_P2_R1957_U87;
  assign new_P2_R1957_U89 = ~new_P2_R1957_U84 | ~new_P2_R1957_U56;
  assign new_P2_R1957_U90 = ~new_P2_U3656 | ~new_P2_R1957_U89;
  assign new_P2_R1957_U91 = ~new_P2_R1957_U83 | ~new_P2_R1957_U58;
  assign new_P2_R1957_U92 = ~new_P2_U3658 | ~new_P2_R1957_U91;
  assign new_P2_R1957_U93 = ~new_P2_R1957_U27;
  assign new_P2_R1957_U94 = ~new_P2_R1957_U28;
  assign new_P2_R1957_U95 = ~new_P2_R1957_U29;
  assign new_P2_R1957_U96 = ~new_P2_R1957_U30;
  assign new_P2_R1957_U97 = ~new_P2_R1957_U31;
  assign new_P2_R1957_U98 = ~new_P2_R1957_U32;
  assign new_P2_R1957_U99 = ~new_P2_R1957_U33;
  assign new_P2_R1957_U100 = ~new_P2_R1957_U34;
  assign new_P2_R1957_U101 = ~new_P2_R1957_U35;
  assign new_P2_R1957_U102 = ~new_P2_R1957_U36;
  assign new_P2_R1957_U103 = ~new_P2_R1957_U37;
  assign new_P2_R1957_U104 = new_P2_U3682 | new_P2_U3683;
  assign new_P2_R1957_U105 = ~new_P2_U3671 | ~new_P2_R1957_U104;
  assign new_P2_R1957_U106 = ~new_P2_U3661 | ~new_P2_R1957_U36;
  assign new_P2_R1957_U107 = ~new_P2_R1957_U101 | ~new_P2_R1957_U63;
  assign new_P2_R1957_U108 = ~new_P2_U3662 | ~new_P2_R1957_U107;
  assign new_P2_R1957_U109 = ~new_P2_R1957_U100 | ~new_P2_R1957_U65;
  assign new_P2_R1957_U110 = ~new_P2_U3664 | ~new_P2_R1957_U109;
  assign new_P2_R1957_U111 = ~new_P2_R1957_U99 | ~new_P2_R1957_U67;
  assign new_P2_R1957_U112 = ~new_P2_U3666 | ~new_P2_R1957_U111;
  assign new_P2_R1957_U113 = ~new_P2_R1957_U98 | ~new_P2_R1957_U69;
  assign new_P2_R1957_U114 = ~new_P2_U3668 | ~new_P2_R1957_U113;
  assign new_P2_R1957_U115 = ~new_P2_R1957_U97 | ~new_P2_R1957_U73;
  assign new_P2_R1957_U116 = ~new_P2_U3670 | ~new_P2_R1957_U115;
  assign new_P2_R1957_U117 = ~new_P2_R1957_U96 | ~new_P2_R1957_U75;
  assign new_P2_R1957_U118 = ~new_P2_U3673 | ~new_P2_R1957_U117;
  assign new_P2_R1957_U119 = ~new_P2_R1957_U95 | ~new_P2_R1957_U77;
  assign new_P2_R1957_U120 = ~new_P2_U3675 | ~new_P2_R1957_U119;
  assign new_P2_R1957_U121 = ~new_P2_R1957_U94 | ~new_P2_R1957_U79;
  assign new_P2_R1957_U122 = ~new_P2_U3677 | ~new_P2_R1957_U121;
  assign new_P2_R1957_U123 = ~new_P2_R1957_U93 | ~new_P2_R1957_U81;
  assign new_P2_R1957_U124 = ~new_P2_U3679 | ~new_P2_R1957_U123;
  assign new_P2_R1957_U125 = ~new_P2_R1957_U86 | ~new_P2_R1957_U52;
  assign new_P2_R1957_U126 = ~new_P2_U3681 | ~new_P2_R1957_U125;
  assign new_P2_R1957_U127 = ~new_P2_R1957_U103 | ~new_P2_R1957_U61;
  assign new_P2_R1957_U128 = ~new_P2_U3653 | ~new_P2_R1957_U24;
  assign new_P2_R1957_U129 = ~new_P2_R1957_U86 | ~new_P2_R1957_U52;
  assign new_P2_R1957_U130 = ~new_P2_U3655 | ~new_P2_R1957_U23;
  assign new_P2_R1957_U131 = ~new_P2_R1957_U85 | ~new_P2_R1957_U54;
  assign new_P2_R1957_U132 = ~new_P2_U3657 | ~new_P2_R1957_U22;
  assign new_P2_R1957_U133 = ~new_P2_R1957_U84 | ~new_P2_R1957_U56;
  assign new_P2_R1957_U134 = ~new_P2_U3660 | ~new_P2_R1957_U21;
  assign new_P2_R1957_U135 = ~new_P2_R1957_U83 | ~new_P2_R1957_U58;
  assign new_P2_R1957_U136 = ~new_P2_R1957_U127 | ~new_P2_R1957_U60;
  assign new_P2_R1957_U137 = ~new_P2_U3647 | ~new_P2_R1957_U103 | ~new_P2_R1957_U61;
  assign new_P2_R1957_U138 = ~new_P2_U3659 | ~new_P2_R1957_U37;
  assign new_P2_R1957_U139 = ~new_P2_R1957_U103 | ~new_P2_R1957_U61;
  assign new_P2_R1957_U140 = ~new_P2_U3663 | ~new_P2_R1957_U35;
  assign new_P2_R1957_U141 = ~new_P2_R1957_U101 | ~new_P2_R1957_U63;
  assign new_P2_R1957_U142 = ~new_P2_U3665 | ~new_P2_R1957_U34;
  assign new_P2_R1957_U143 = ~new_P2_R1957_U100 | ~new_P2_R1957_U65;
  assign new_P2_R1957_U144 = ~new_P2_U3667 | ~new_P2_R1957_U33;
  assign new_P2_R1957_U145 = ~new_P2_R1957_U99 | ~new_P2_R1957_U67;
  assign new_P2_R1957_U146 = ~new_P2_U3669 | ~new_P2_R1957_U32;
  assign new_P2_R1957_U147 = ~new_P2_R1957_U98 | ~new_P2_R1957_U69;
  assign new_P2_R1957_U148 = ~new_P2_U3682 | ~new_P2_R1957_U72;
  assign new_P2_R1957_U149 = ~new_P2_U3683 | ~new_P2_R1957_U71;
  assign new_P2_R1957_U150 = ~new_P2_U3672 | ~new_P2_R1957_U31;
  assign new_P2_R1957_U151 = ~new_P2_R1957_U97 | ~new_P2_R1957_U73;
  assign new_P2_R1957_U152 = ~new_P2_U3674 | ~new_P2_R1957_U30;
  assign new_P2_R1957_U153 = ~new_P2_R1957_U96 | ~new_P2_R1957_U75;
  assign new_P2_R1957_U154 = ~new_P2_U3676 | ~new_P2_R1957_U29;
  assign new_P2_R1957_U155 = ~new_P2_R1957_U95 | ~new_P2_R1957_U77;
  assign new_P2_R1957_U156 = ~new_P2_U3678 | ~new_P2_R1957_U28;
  assign new_P2_R1957_U157 = ~new_P2_R1957_U94 | ~new_P2_R1957_U79;
  assign new_P2_R1957_U158 = ~new_P2_U3680 | ~new_P2_R1957_U27;
  assign new_P2_R1957_U159 = ~new_P2_R1957_U93 | ~new_P2_R1957_U81;
  assign new_P2_R2278_U4 = new_P2_R2278_U399 & new_P2_R2278_U398;
  assign new_P2_R2278_U5 = new_P2_R2278_U206 & new_P2_R2278_U161 & new_P2_R2278_U309;
  assign new_P2_R2278_U6 = ~new_P2_R2278_U345 | ~new_P2_R2278_U490 | ~new_P2_R2278_U489;
  assign new_P2_R2278_U7 = ~new_P2_U3631;
  assign new_P2_R2278_U8 = ~P2_INSTADDRPOINTER_REG_7_;
  assign new_P2_R2278_U9 = ~new_P2_U3633;
  assign new_P2_R2278_U10 = ~P2_INSTADDRPOINTER_REG_5_;
  assign new_P2_R2278_U11 = ~new_P2_U3635;
  assign new_P2_R2278_U12 = ~P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_R2278_U13 = ~new_P2_U3638;
  assign new_P2_R2278_U14 = ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_R2278_U15 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_U3638;
  assign new_P2_R2278_U16 = ~new_P2_U3637;
  assign new_P2_R2278_U17 = ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_R2278_U18 = ~new_P2_U3636;
  assign new_P2_R2278_U19 = ~P2_INSTADDRPOINTER_REG_2_;
  assign new_P2_R2278_U20 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_U3636;
  assign new_P2_R2278_U21 = ~new_P2_U3634;
  assign new_P2_R2278_U22 = ~P2_INSTADDRPOINTER_REG_4_;
  assign new_P2_R2278_U23 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_U3634;
  assign new_P2_R2278_U24 = ~new_P2_U3632;
  assign new_P2_R2278_U25 = ~P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_R2278_U26 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_U3632;
  assign new_P2_R2278_U27 = ~new_P2_U3630;
  assign new_P2_R2278_U28 = ~P2_INSTADDRPOINTER_REG_8_;
  assign new_P2_R2278_U29 = ~P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_R2278_U30 = ~new_P2_U2812;
  assign new_P2_R2278_U31 = ~new_P2_U2793;
  assign new_P2_R2278_U32 = ~P2_INSTADDRPOINTER_REG_28_;
  assign new_P2_R2278_U33 = ~new_P2_U2792;
  assign new_P2_R2278_U34 = ~P2_INSTADDRPOINTER_REG_29_;
  assign new_P2_R2278_U35 = ~new_P2_U2797;
  assign new_P2_R2278_U36 = ~P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_R2278_U37 = ~new_P2_U2799;
  assign new_P2_R2278_U38 = ~P2_INSTADDRPOINTER_REG_22_;
  assign new_P2_R2278_U39 = ~new_P2_U2801;
  assign new_P2_R2278_U40 = ~P2_INSTADDRPOINTER_REG_20_;
  assign new_P2_R2278_U41 = ~new_P2_U2804;
  assign new_P2_R2278_U42 = ~P2_INSTADDRPOINTER_REG_17_;
  assign new_P2_R2278_U43 = ~new_P2_U2806;
  assign new_P2_R2278_U44 = ~P2_INSTADDRPOINTER_REG_15_;
  assign new_P2_R2278_U45 = ~new_P2_U2808;
  assign new_P2_R2278_U46 = ~P2_INSTADDRPOINTER_REG_13_;
  assign new_P2_R2278_U47 = ~new_P2_U2810;
  assign new_P2_R2278_U48 = ~P2_INSTADDRPOINTER_REG_11_;
  assign new_P2_R2278_U49 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_U3630;
  assign new_P2_R2278_U50 = ~new_P2_U2811;
  assign new_P2_R2278_U51 = ~P2_INSTADDRPOINTER_REG_10_;
  assign new_P2_R2278_U52 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_U2811;
  assign new_P2_R2278_U53 = ~new_P2_U2809;
  assign new_P2_R2278_U54 = ~P2_INSTADDRPOINTER_REG_12_;
  assign new_P2_R2278_U55 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_U2809;
  assign new_P2_R2278_U56 = ~new_P2_U2807;
  assign new_P2_R2278_U57 = ~P2_INSTADDRPOINTER_REG_14_;
  assign new_P2_R2278_U58 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_U2807;
  assign new_P2_R2278_U59 = ~new_P2_U2805;
  assign new_P2_R2278_U60 = ~P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_R2278_U61 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_U2805;
  assign new_P2_R2278_U62 = ~new_P2_U2802;
  assign new_P2_R2278_U63 = ~P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_R2278_U64 = ~new_P2_U2803;
  assign new_P2_R2278_U65 = ~P2_INSTADDRPOINTER_REG_18_;
  assign new_P2_R2278_U66 = ~new_P2_U2800;
  assign new_P2_R2278_U67 = ~P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_R2278_U68 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_U2800;
  assign new_P2_R2278_U69 = ~new_P2_U2798;
  assign new_P2_R2278_U70 = ~P2_INSTADDRPOINTER_REG_23_;
  assign new_P2_R2278_U71 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_U2798;
  assign new_P2_R2278_U72 = ~new_P2_U2796;
  assign new_P2_R2278_U73 = ~P2_INSTADDRPOINTER_REG_25_;
  assign new_P2_R2278_U74 = ~new_P2_U2794;
  assign new_P2_R2278_U75 = ~P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_R2278_U76 = ~new_P2_U2795;
  assign new_P2_R2278_U77 = ~P2_INSTADDRPOINTER_REG_26_;
  assign new_P2_R2278_U78 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_U2795;
  assign new_P2_R2278_U79 = ~new_P2_U2791;
  assign new_P2_R2278_U80 = ~P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_R2278_U81 = ~new_P2_R2278_U340 | ~new_P2_R2278_U297;
  assign new_P2_R2278_U82 = ~new_P2_U3637 | ~new_P2_R2278_U208;
  assign new_P2_R2278_U83 = ~new_P2_R2278_U562 | ~new_P2_R2278_U561;
  assign new_P2_R2278_U84 = ~new_P2_R2278_U352 | ~new_P2_R2278_U351;
  assign new_P2_R2278_U85 = ~new_P2_R2278_U359 | ~new_P2_R2278_U358;
  assign new_P2_R2278_U86 = ~new_P2_R2278_U366 | ~new_P2_R2278_U365;
  assign new_P2_R2278_U87 = ~new_P2_R2278_U373 | ~new_P2_R2278_U372;
  assign new_P2_R2278_U88 = ~new_P2_R2278_U380 | ~new_P2_R2278_U379;
  assign new_P2_R2278_U89 = ~new_P2_R2278_U387 | ~new_P2_R2278_U386;
  assign new_P2_R2278_U90 = ~new_P2_R2278_U394 | ~new_P2_R2278_U393;
  assign new_P2_R2278_U91 = ~new_P2_R2278_U408 | ~new_P2_R2278_U407;
  assign new_P2_R2278_U92 = ~new_P2_R2278_U415 | ~new_P2_R2278_U414;
  assign new_P2_R2278_U93 = ~new_P2_R2278_U422 | ~new_P2_R2278_U421;
  assign new_P2_R2278_U94 = ~new_P2_R2278_U429 | ~new_P2_R2278_U428;
  assign new_P2_R2278_U95 = ~new_P2_R2278_U436 | ~new_P2_R2278_U435;
  assign new_P2_R2278_U96 = ~new_P2_R2278_U443 | ~new_P2_R2278_U442;
  assign new_P2_R2278_U97 = ~new_P2_R2278_U450 | ~new_P2_R2278_U449;
  assign new_P2_R2278_U98 = ~new_P2_R2278_U457 | ~new_P2_R2278_U456;
  assign new_P2_R2278_U99 = ~new_P2_R2278_U464 | ~new_P2_R2278_U463;
  assign new_P2_R2278_U100 = ~new_P2_R2278_U471 | ~new_P2_R2278_U470;
  assign new_P2_R2278_U101 = ~new_P2_R2278_U478 | ~new_P2_R2278_U477;
  assign new_P2_R2278_U102 = ~new_P2_R2278_U485 | ~new_P2_R2278_U484;
  assign new_P2_R2278_U103 = ~new_P2_R2278_U497 | ~new_P2_R2278_U496;
  assign new_P2_R2278_U104 = ~new_P2_R2278_U504 | ~new_P2_R2278_U503;
  assign new_P2_R2278_U105 = ~new_P2_R2278_U511 | ~new_P2_R2278_U510;
  assign new_P2_R2278_U106 = ~new_P2_R2278_U518 | ~new_P2_R2278_U517;
  assign new_P2_R2278_U107 = ~new_P2_R2278_U525 | ~new_P2_R2278_U524;
  assign new_P2_R2278_U108 = ~new_P2_R2278_U532 | ~new_P2_R2278_U531;
  assign new_P2_R2278_U109 = ~new_P2_R2278_U539 | ~new_P2_R2278_U538;
  assign new_P2_R2278_U110 = ~new_P2_R2278_U546 | ~new_P2_R2278_U545;
  assign new_P2_R2278_U111 = ~new_P2_R2278_U553 | ~new_P2_R2278_U552;
  assign new_P2_R2278_U112 = ~new_P2_R2278_U560 | ~new_P2_R2278_U559;
  assign new_P2_R2278_U113 = new_P2_R2278_U210 & new_P2_R2278_U314;
  assign new_P2_R2278_U114 = new_P2_R2278_U313 & new_P2_R2278_U215;
  assign new_P2_R2278_U115 = new_P2_R2278_U217 & new_P2_R2278_U221;
  assign new_P2_R2278_U116 = new_P2_R2278_U316 & new_P2_R2278_U222;
  assign new_P2_R2278_U117 = new_P2_R2278_U224 & new_P2_R2278_U228;
  assign new_P2_R2278_U118 = new_P2_R2278_U318 & new_P2_R2278_U229;
  assign new_P2_R2278_U119 = new_P2_R2278_U231 & new_P2_R2278_U235;
  assign new_P2_R2278_U120 = new_P2_R2278_U320 & new_P2_R2278_U236;
  assign new_P2_R2278_U121 = new_P2_R2278_U238 & new_P2_R2278_U242;
  assign new_P2_R2278_U122 = new_P2_R2278_U322 & new_P2_R2278_U243;
  assign new_P2_R2278_U123 = new_P2_R2278_U245 & new_P2_R2278_U249;
  assign new_P2_R2278_U124 = new_P2_R2278_U324 & new_P2_R2278_U250;
  assign new_P2_R2278_U125 = new_P2_R2278_U252 & new_P2_R2278_U256;
  assign new_P2_R2278_U126 = new_P2_R2278_U326 & new_P2_R2278_U257;
  assign new_P2_R2278_U127 = new_P2_R2278_U259 & new_P2_R2278_U263;
  assign new_P2_R2278_U128 = new_P2_R2278_U328 & new_P2_R2278_U264;
  assign new_P2_R2278_U129 = new_P2_R2278_U273 & new_P2_R2278_U270;
  assign new_P2_R2278_U130 = new_P2_R2278_U331 & new_P2_R2278_U273;
  assign new_P2_R2278_U131 = new_P2_R2278_U334 & new_P2_R2278_U274;
  assign new_P2_R2278_U132 = new_P2_R2278_U276 & new_P2_R2278_U280;
  assign new_P2_R2278_U133 = new_P2_R2278_U336 & new_P2_R2278_U281;
  assign new_P2_R2278_U134 = new_P2_R2278_U283 & new_P2_R2278_U287;
  assign new_P2_R2278_U135 = new_P2_R2278_U338 & new_P2_R2278_U288;
  assign new_P2_R2278_U136 = new_P2_R2278_U292 & new_P2_R2278_U299 & new_P2_R2278_U296;
  assign new_P2_R2278_U137 = new_P2_R2278_U304 & new_P2_R2278_U300;
  assign new_P2_R2278_U138 = new_P2_R2278_U307 & new_P2_R2278_U302;
  assign new_P2_R2278_U139 = new_P2_R2278_U397 & new_P2_R2278_U138;
  assign new_P2_R2278_U140 = new_P2_R2278_U343 & new_P2_R2278_U300;
  assign new_P2_R2278_U141 = new_P2_R2278_U4 & new_P2_R2278_U142;
  assign new_P2_R2278_U142 = new_P2_R2278_U304 & new_P2_R2278_U306;
  assign new_P2_R2278_U143 = new_P2_R2278_U292 & new_P2_R2278_U296;
  assign new_P2_R2278_U144 = new_P2_R2278_U266 & new_P2_R2278_U270;
  assign new_P2_R2278_U145 = new_P2_R2278_U347 & new_P2_R2278_U346;
  assign new_P2_R2278_U146 = ~new_P2_R2278_U49 | ~new_P2_R2278_U232;
  assign new_P2_R2278_U147 = new_P2_R2278_U354 & new_P2_R2278_U353;
  assign new_P2_R2278_U148 = ~new_P2_R2278_U118 | ~new_P2_R2278_U317;
  assign new_P2_R2278_U149 = new_P2_R2278_U361 & new_P2_R2278_U360;
  assign new_P2_R2278_U150 = ~new_P2_R2278_U26 | ~new_P2_R2278_U225;
  assign new_P2_R2278_U151 = new_P2_R2278_U368 & new_P2_R2278_U367;
  assign new_P2_R2278_U152 = ~new_P2_R2278_U116 | ~new_P2_R2278_U315;
  assign new_P2_R2278_U153 = new_P2_R2278_U375 & new_P2_R2278_U374;
  assign new_P2_R2278_U154 = ~new_P2_R2278_U23 | ~new_P2_R2278_U218;
  assign new_P2_R2278_U155 = new_P2_R2278_U382 & new_P2_R2278_U381;
  assign new_P2_R2278_U156 = ~new_P2_R2278_U114 | ~new_P2_R2278_U312;
  assign new_P2_R2278_U157 = new_P2_R2278_U389 & new_P2_R2278_U388;
  assign new_P2_R2278_U158 = ~new_P2_R2278_U20 | ~new_P2_R2278_U211;
  assign new_P2_R2278_U159 = ~P2_INSTADDRPOINTER_REG_31_;
  assign new_P2_R2278_U160 = ~new_P2_U2790;
  assign new_P2_R2278_U161 = new_P2_R2278_U401 & new_P2_R2278_U400;
  assign new_P2_R2278_U162 = new_P2_R2278_U403 & new_P2_R2278_U402;
  assign new_P2_R2278_U163 = ~new_P2_R2278_U304 | ~new_P2_R2278_U303;
  assign new_P2_R2278_U164 = new_P2_R2278_U410 & new_P2_R2278_U409;
  assign new_P2_R2278_U165 = ~new_P2_R2278_U311 | ~new_P2_R2278_U310 | ~new_P2_R2278_U82;
  assign new_P2_R2278_U166 = new_P2_R2278_U417 & new_P2_R2278_U416;
  assign new_P2_R2278_U167 = ~new_P2_R2278_U140 | ~new_P2_R2278_U342;
  assign new_P2_R2278_U168 = new_P2_R2278_U424 & new_P2_R2278_U423;
  assign new_P2_R2278_U169 = ~new_P2_R2278_U341 | ~new_P2_R2278_U339;
  assign new_P2_R2278_U170 = new_P2_R2278_U431 & new_P2_R2278_U430;
  assign new_P2_R2278_U171 = ~new_P2_R2278_U78 | ~new_P2_R2278_U293;
  assign new_P2_R2278_U172 = new_P2_R2278_U438 & new_P2_R2278_U437;
  assign new_P2_R2278_U173 = ~new_P2_R2278_U308 | ~new_P2_R2278_U290 | ~new_P2_R2278_U205;
  assign new_P2_R2278_U174 = ~new_P2_R2278_U135 | ~new_P2_R2278_U337;
  assign new_P2_R2278_U175 = new_P2_R2278_U452 & new_P2_R2278_U451;
  assign new_P2_R2278_U176 = ~new_P2_R2278_U71 | ~new_P2_R2278_U284;
  assign new_P2_R2278_U177 = new_P2_R2278_U459 & new_P2_R2278_U458;
  assign new_P2_R2278_U178 = ~new_P2_R2278_U133 | ~new_P2_R2278_U335;
  assign new_P2_R2278_U179 = new_P2_R2278_U466 & new_P2_R2278_U465;
  assign new_P2_R2278_U180 = ~new_P2_R2278_U68 | ~new_P2_R2278_U277;
  assign new_P2_R2278_U181 = new_P2_R2278_U473 & new_P2_R2278_U472;
  assign new_P2_R2278_U182 = ~new_P2_R2278_U131 | ~new_P2_R2278_U333;
  assign new_P2_R2278_U183 = new_P2_R2278_U480 & new_P2_R2278_U479;
  assign new_P2_R2278_U184 = ~new_P2_R2278_U330 | ~new_P2_R2278_U329;
  assign new_P2_R2278_U185 = new_P2_R2278_U492 & new_P2_R2278_U491;
  assign new_P2_R2278_U186 = ~new_P2_R2278_U268 | ~new_P2_R2278_U267;
  assign new_P2_R2278_U187 = new_P2_R2278_U499 & new_P2_R2278_U498;
  assign new_P2_R2278_U188 = ~new_P2_R2278_U128 | ~new_P2_R2278_U327;
  assign new_P2_R2278_U189 = new_P2_R2278_U506 & new_P2_R2278_U505;
  assign new_P2_R2278_U190 = ~new_P2_R2278_U61 | ~new_P2_R2278_U260;
  assign new_P2_R2278_U191 = new_P2_R2278_U513 & new_P2_R2278_U512;
  assign new_P2_R2278_U192 = ~new_P2_R2278_U126 | ~new_P2_R2278_U325;
  assign new_P2_R2278_U193 = new_P2_R2278_U520 & new_P2_R2278_U519;
  assign new_P2_R2278_U194 = ~new_P2_R2278_U58 | ~new_P2_R2278_U253;
  assign new_P2_R2278_U195 = new_P2_R2278_U527 & new_P2_R2278_U526;
  assign new_P2_R2278_U196 = ~new_P2_R2278_U124 | ~new_P2_R2278_U323;
  assign new_P2_R2278_U197 = new_P2_R2278_U534 & new_P2_R2278_U533;
  assign new_P2_R2278_U198 = ~new_P2_R2278_U55 | ~new_P2_R2278_U246;
  assign new_P2_R2278_U199 = new_P2_R2278_U541 & new_P2_R2278_U540;
  assign new_P2_R2278_U200 = ~new_P2_R2278_U122 | ~new_P2_R2278_U321;
  assign new_P2_R2278_U201 = new_P2_R2278_U548 & new_P2_R2278_U547;
  assign new_P2_R2278_U202 = ~new_P2_R2278_U52 | ~new_P2_R2278_U239;
  assign new_P2_R2278_U203 = new_P2_R2278_U555 & new_P2_R2278_U554;
  assign new_P2_R2278_U204 = ~new_P2_R2278_U120 | ~new_P2_R2278_U319;
  assign new_P2_R2278_U205 = ~new_P2_U2796 | ~new_P2_R2278_U174;
  assign new_P2_R2278_U206 = ~new_P2_R2278_U139 | ~new_P2_R2278_U344;
  assign new_P2_R2278_U207 = ~new_P2_R2278_U82;
  assign new_P2_R2278_U208 = ~new_P2_R2278_U15;
  assign new_P2_R2278_U209 = ~new_P2_R2278_U165;
  assign new_P2_R2278_U210 = new_P2_U3636 | P2_INSTADDRPOINTER_REG_2_;
  assign new_P2_R2278_U211 = ~new_P2_R2278_U210 | ~new_P2_R2278_U165;
  assign new_P2_R2278_U212 = ~new_P2_R2278_U20;
  assign new_P2_R2278_U213 = ~new_P2_R2278_U158;
  assign new_P2_R2278_U214 = new_P2_U3635 | P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_R2278_U215 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_U3635;
  assign new_P2_R2278_U216 = ~new_P2_R2278_U156;
  assign new_P2_R2278_U217 = new_P2_U3634 | P2_INSTADDRPOINTER_REG_4_;
  assign new_P2_R2278_U218 = ~new_P2_R2278_U217 | ~new_P2_R2278_U156;
  assign new_P2_R2278_U219 = ~new_P2_R2278_U23;
  assign new_P2_R2278_U220 = ~new_P2_R2278_U154;
  assign new_P2_R2278_U221 = new_P2_U3633 | P2_INSTADDRPOINTER_REG_5_;
  assign new_P2_R2278_U222 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_U3633;
  assign new_P2_R2278_U223 = ~new_P2_R2278_U152;
  assign new_P2_R2278_U224 = new_P2_U3632 | P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_R2278_U225 = ~new_P2_R2278_U224 | ~new_P2_R2278_U152;
  assign new_P2_R2278_U226 = ~new_P2_R2278_U26;
  assign new_P2_R2278_U227 = ~new_P2_R2278_U150;
  assign new_P2_R2278_U228 = new_P2_U3631 | P2_INSTADDRPOINTER_REG_7_;
  assign new_P2_R2278_U229 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_U3631;
  assign new_P2_R2278_U230 = ~new_P2_R2278_U148;
  assign new_P2_R2278_U231 = new_P2_U3630 | P2_INSTADDRPOINTER_REG_8_;
  assign new_P2_R2278_U232 = ~new_P2_R2278_U231 | ~new_P2_R2278_U148;
  assign new_P2_R2278_U233 = ~new_P2_R2278_U49;
  assign new_P2_R2278_U234 = ~new_P2_R2278_U146;
  assign new_P2_R2278_U235 = new_P2_U2812 | P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_R2278_U236 = ~new_P2_U2812 | ~P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_R2278_U237 = ~new_P2_R2278_U204;
  assign new_P2_R2278_U238 = new_P2_U2811 | P2_INSTADDRPOINTER_REG_10_;
  assign new_P2_R2278_U239 = ~new_P2_R2278_U238 | ~new_P2_R2278_U204;
  assign new_P2_R2278_U240 = ~new_P2_R2278_U52;
  assign new_P2_R2278_U241 = ~new_P2_R2278_U202;
  assign new_P2_R2278_U242 = new_P2_U2810 | P2_INSTADDRPOINTER_REG_11_;
  assign new_P2_R2278_U243 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_U2810;
  assign new_P2_R2278_U244 = ~new_P2_R2278_U200;
  assign new_P2_R2278_U245 = new_P2_U2809 | P2_INSTADDRPOINTER_REG_12_;
  assign new_P2_R2278_U246 = ~new_P2_R2278_U245 | ~new_P2_R2278_U200;
  assign new_P2_R2278_U247 = ~new_P2_R2278_U55;
  assign new_P2_R2278_U248 = ~new_P2_R2278_U198;
  assign new_P2_R2278_U249 = new_P2_U2808 | P2_INSTADDRPOINTER_REG_13_;
  assign new_P2_R2278_U250 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_U2808;
  assign new_P2_R2278_U251 = ~new_P2_R2278_U196;
  assign new_P2_R2278_U252 = new_P2_U2807 | P2_INSTADDRPOINTER_REG_14_;
  assign new_P2_R2278_U253 = ~new_P2_R2278_U252 | ~new_P2_R2278_U196;
  assign new_P2_R2278_U254 = ~new_P2_R2278_U58;
  assign new_P2_R2278_U255 = ~new_P2_R2278_U194;
  assign new_P2_R2278_U256 = new_P2_U2806 | P2_INSTADDRPOINTER_REG_15_;
  assign new_P2_R2278_U257 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_U2806;
  assign new_P2_R2278_U258 = ~new_P2_R2278_U192;
  assign new_P2_R2278_U259 = new_P2_U2805 | P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_R2278_U260 = ~new_P2_R2278_U259 | ~new_P2_R2278_U192;
  assign new_P2_R2278_U261 = ~new_P2_R2278_U61;
  assign new_P2_R2278_U262 = ~new_P2_R2278_U190;
  assign new_P2_R2278_U263 = new_P2_U2804 | P2_INSTADDRPOINTER_REG_17_;
  assign new_P2_R2278_U264 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_U2804;
  assign new_P2_R2278_U265 = ~new_P2_R2278_U188;
  assign new_P2_R2278_U266 = new_P2_U2803 | P2_INSTADDRPOINTER_REG_18_;
  assign new_P2_R2278_U267 = ~new_P2_R2278_U266 | ~new_P2_R2278_U188;
  assign new_P2_R2278_U268 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_U2803;
  assign new_P2_R2278_U269 = ~new_P2_R2278_U186;
  assign new_P2_R2278_U270 = new_P2_U2802 | P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_R2278_U271 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_U2802;
  assign new_P2_R2278_U272 = ~new_P2_R2278_U184;
  assign new_P2_R2278_U273 = new_P2_U2801 | P2_INSTADDRPOINTER_REG_20_;
  assign new_P2_R2278_U274 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_U2801;
  assign new_P2_R2278_U275 = ~new_P2_R2278_U182;
  assign new_P2_R2278_U276 = new_P2_U2800 | P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_R2278_U277 = ~new_P2_R2278_U276 | ~new_P2_R2278_U182;
  assign new_P2_R2278_U278 = ~new_P2_R2278_U68;
  assign new_P2_R2278_U279 = ~new_P2_R2278_U180;
  assign new_P2_R2278_U280 = new_P2_U2799 | P2_INSTADDRPOINTER_REG_22_;
  assign new_P2_R2278_U281 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_U2799;
  assign new_P2_R2278_U282 = ~new_P2_R2278_U178;
  assign new_P2_R2278_U283 = new_P2_U2798 | P2_INSTADDRPOINTER_REG_23_;
  assign new_P2_R2278_U284 = ~new_P2_R2278_U283 | ~new_P2_R2278_U178;
  assign new_P2_R2278_U285 = ~new_P2_R2278_U71;
  assign new_P2_R2278_U286 = ~new_P2_R2278_U176;
  assign new_P2_R2278_U287 = new_P2_U2797 | P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_R2278_U288 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_U2797;
  assign new_P2_R2278_U289 = ~new_P2_R2278_U174;
  assign new_P2_R2278_U290 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_R2278_U174;
  assign new_P2_R2278_U291 = ~new_P2_R2278_U173;
  assign new_P2_R2278_U292 = new_P2_U2795 | P2_INSTADDRPOINTER_REG_26_;
  assign new_P2_R2278_U293 = ~new_P2_R2278_U292 | ~new_P2_R2278_U173;
  assign new_P2_R2278_U294 = ~new_P2_R2278_U78;
  assign new_P2_R2278_U295 = ~new_P2_R2278_U171;
  assign new_P2_R2278_U296 = new_P2_U2794 | P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_R2278_U297 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_U2794;
  assign new_P2_R2278_U298 = ~new_P2_R2278_U169;
  assign new_P2_R2278_U299 = new_P2_U2793 | P2_INSTADDRPOINTER_REG_28_;
  assign new_P2_R2278_U300 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_U2793;
  assign new_P2_R2278_U301 = ~new_P2_R2278_U167;
  assign new_P2_R2278_U302 = new_P2_U2792 | P2_INSTADDRPOINTER_REG_29_;
  assign new_P2_R2278_U303 = ~new_P2_R2278_U302 | ~new_P2_R2278_U167;
  assign new_P2_R2278_U304 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_U2792;
  assign new_P2_R2278_U305 = ~new_P2_R2278_U163;
  assign new_P2_R2278_U306 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_U2791;
  assign new_P2_R2278_U307 = P2_INSTADDRPOINTER_REG_30_ | new_P2_U2791;
  assign new_P2_R2278_U308 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_U2796;
  assign new_P2_R2278_U309 = ~new_P2_R2278_U303 | ~new_P2_R2278_U141;
  assign new_P2_R2278_U310 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_R2278_U208;
  assign new_P2_R2278_U311 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_U3637;
  assign new_P2_R2278_U312 = ~new_P2_R2278_U113 | ~new_P2_R2278_U165;
  assign new_P2_R2278_U313 = ~new_P2_R2278_U212 | ~new_P2_R2278_U214;
  assign new_P2_R2278_U314 = new_P2_U3635 | P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_R2278_U315 = ~new_P2_R2278_U115 | ~new_P2_R2278_U156;
  assign new_P2_R2278_U316 = ~new_P2_R2278_U219 | ~new_P2_R2278_U221;
  assign new_P2_R2278_U317 = ~new_P2_R2278_U117 | ~new_P2_R2278_U152;
  assign new_P2_R2278_U318 = ~new_P2_R2278_U226 | ~new_P2_R2278_U228;
  assign new_P2_R2278_U319 = ~new_P2_R2278_U119 | ~new_P2_R2278_U148;
  assign new_P2_R2278_U320 = ~new_P2_R2278_U233 | ~new_P2_R2278_U235;
  assign new_P2_R2278_U321 = ~new_P2_R2278_U121 | ~new_P2_R2278_U204;
  assign new_P2_R2278_U322 = ~new_P2_R2278_U240 | ~new_P2_R2278_U242;
  assign new_P2_R2278_U323 = ~new_P2_R2278_U123 | ~new_P2_R2278_U200;
  assign new_P2_R2278_U324 = ~new_P2_R2278_U247 | ~new_P2_R2278_U249;
  assign new_P2_R2278_U325 = ~new_P2_R2278_U125 | ~new_P2_R2278_U196;
  assign new_P2_R2278_U326 = ~new_P2_R2278_U254 | ~new_P2_R2278_U256;
  assign new_P2_R2278_U327 = ~new_P2_R2278_U127 | ~new_P2_R2278_U192;
  assign new_P2_R2278_U328 = ~new_P2_R2278_U261 | ~new_P2_R2278_U263;
  assign new_P2_R2278_U329 = ~new_P2_R2278_U144 | ~new_P2_R2278_U188;
  assign new_P2_R2278_U330 = ~new_P2_R2278_U331 | ~new_P2_R2278_U332;
  assign new_P2_R2278_U331 = new_P2_U2802 | P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_R2278_U332 = ~new_P2_R2278_U268 | ~new_P2_R2278_U271;
  assign new_P2_R2278_U333 = ~new_P2_R2278_U129 | ~new_P2_R2278_U266 | ~new_P2_R2278_U188;
  assign new_P2_R2278_U334 = ~new_P2_R2278_U130 | ~new_P2_R2278_U332;
  assign new_P2_R2278_U335 = ~new_P2_R2278_U132 | ~new_P2_R2278_U182;
  assign new_P2_R2278_U336 = ~new_P2_R2278_U278 | ~new_P2_R2278_U280;
  assign new_P2_R2278_U337 = ~new_P2_R2278_U134 | ~new_P2_R2278_U178;
  assign new_P2_R2278_U338 = ~new_P2_R2278_U285 | ~new_P2_R2278_U287;
  assign new_P2_R2278_U339 = ~new_P2_R2278_U143 | ~new_P2_R2278_U173;
  assign new_P2_R2278_U340 = ~new_P2_R2278_U294 | ~new_P2_R2278_U296;
  assign new_P2_R2278_U341 = ~new_P2_R2278_U81;
  assign new_P2_R2278_U342 = ~new_P2_R2278_U173 | ~new_P2_R2278_U136;
  assign new_P2_R2278_U343 = ~new_P2_R2278_U81 | ~new_P2_R2278_U299;
  assign new_P2_R2278_U344 = ~new_P2_R2278_U137 | ~new_P2_R2278_U343 | ~new_P2_R2278_U342;
  assign new_P2_R2278_U345 = ~new_P2_R2278_U207 | ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_R2278_U346 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_R2278_U30;
  assign new_P2_R2278_U347 = ~new_P2_U2812 | ~new_P2_R2278_U29;
  assign new_P2_R2278_U348 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_R2278_U30;
  assign new_P2_R2278_U349 = ~new_P2_U2812 | ~new_P2_R2278_U29;
  assign new_P2_R2278_U350 = ~new_P2_R2278_U349 | ~new_P2_R2278_U348;
  assign new_P2_R2278_U351 = ~new_P2_R2278_U145 | ~new_P2_R2278_U146;
  assign new_P2_R2278_U352 = ~new_P2_R2278_U234 | ~new_P2_R2278_U350;
  assign new_P2_R2278_U353 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_R2278_U27;
  assign new_P2_R2278_U354 = ~new_P2_U3630 | ~new_P2_R2278_U28;
  assign new_P2_R2278_U355 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_R2278_U27;
  assign new_P2_R2278_U356 = ~new_P2_U3630 | ~new_P2_R2278_U28;
  assign new_P2_R2278_U357 = ~new_P2_R2278_U356 | ~new_P2_R2278_U355;
  assign new_P2_R2278_U358 = ~new_P2_R2278_U147 | ~new_P2_R2278_U148;
  assign new_P2_R2278_U359 = ~new_P2_R2278_U230 | ~new_P2_R2278_U357;
  assign new_P2_R2278_U360 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_R2278_U7;
  assign new_P2_R2278_U361 = ~new_P2_U3631 | ~new_P2_R2278_U8;
  assign new_P2_R2278_U362 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_R2278_U7;
  assign new_P2_R2278_U363 = ~new_P2_U3631 | ~new_P2_R2278_U8;
  assign new_P2_R2278_U364 = ~new_P2_R2278_U363 | ~new_P2_R2278_U362;
  assign new_P2_R2278_U365 = ~new_P2_R2278_U149 | ~new_P2_R2278_U150;
  assign new_P2_R2278_U366 = ~new_P2_R2278_U227 | ~new_P2_R2278_U364;
  assign new_P2_R2278_U367 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_R2278_U24;
  assign new_P2_R2278_U368 = ~new_P2_U3632 | ~new_P2_R2278_U25;
  assign new_P2_R2278_U369 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_R2278_U24;
  assign new_P2_R2278_U370 = ~new_P2_U3632 | ~new_P2_R2278_U25;
  assign new_P2_R2278_U371 = ~new_P2_R2278_U370 | ~new_P2_R2278_U369;
  assign new_P2_R2278_U372 = ~new_P2_R2278_U151 | ~new_P2_R2278_U152;
  assign new_P2_R2278_U373 = ~new_P2_R2278_U223 | ~new_P2_R2278_U371;
  assign new_P2_R2278_U374 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_R2278_U9;
  assign new_P2_R2278_U375 = ~new_P2_U3633 | ~new_P2_R2278_U10;
  assign new_P2_R2278_U376 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_R2278_U9;
  assign new_P2_R2278_U377 = ~new_P2_U3633 | ~new_P2_R2278_U10;
  assign new_P2_R2278_U378 = ~new_P2_R2278_U377 | ~new_P2_R2278_U376;
  assign new_P2_R2278_U379 = ~new_P2_R2278_U153 | ~new_P2_R2278_U154;
  assign new_P2_R2278_U380 = ~new_P2_R2278_U220 | ~new_P2_R2278_U378;
  assign new_P2_R2278_U381 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_R2278_U21;
  assign new_P2_R2278_U382 = ~new_P2_U3634 | ~new_P2_R2278_U22;
  assign new_P2_R2278_U383 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_R2278_U21;
  assign new_P2_R2278_U384 = ~new_P2_U3634 | ~new_P2_R2278_U22;
  assign new_P2_R2278_U385 = ~new_P2_R2278_U384 | ~new_P2_R2278_U383;
  assign new_P2_R2278_U386 = ~new_P2_R2278_U155 | ~new_P2_R2278_U156;
  assign new_P2_R2278_U387 = ~new_P2_R2278_U216 | ~new_P2_R2278_U385;
  assign new_P2_R2278_U388 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_R2278_U11;
  assign new_P2_R2278_U389 = ~new_P2_U3635 | ~new_P2_R2278_U12;
  assign new_P2_R2278_U390 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_R2278_U11;
  assign new_P2_R2278_U391 = ~new_P2_U3635 | ~new_P2_R2278_U12;
  assign new_P2_R2278_U392 = ~new_P2_R2278_U391 | ~new_P2_R2278_U390;
  assign new_P2_R2278_U393 = ~new_P2_R2278_U157 | ~new_P2_R2278_U158;
  assign new_P2_R2278_U394 = ~new_P2_R2278_U213 | ~new_P2_R2278_U392;
  assign new_P2_R2278_U395 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_R2278_U160;
  assign new_P2_R2278_U396 = ~new_P2_U2790 | ~new_P2_R2278_U159;
  assign new_P2_R2278_U397 = ~new_P2_R2278_U396 | ~new_P2_R2278_U395;
  assign new_P2_R2278_U398 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_R2278_U160;
  assign new_P2_R2278_U399 = ~new_P2_U2790 | ~new_P2_R2278_U159;
  assign new_P2_R2278_U400 = ~new_P2_R2278_U80 | ~new_P2_R2278_U4 | ~new_P2_R2278_U79;
  assign new_P2_R2278_U401 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_U2791 | ~new_P2_R2278_U397;
  assign new_P2_R2278_U402 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_R2278_U79;
  assign new_P2_R2278_U403 = ~new_P2_U2791 | ~new_P2_R2278_U80;
  assign new_P2_R2278_U404 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_R2278_U79;
  assign new_P2_R2278_U405 = ~new_P2_U2791 | ~new_P2_R2278_U80;
  assign new_P2_R2278_U406 = ~new_P2_R2278_U405 | ~new_P2_R2278_U404;
  assign new_P2_R2278_U407 = ~new_P2_R2278_U162 | ~new_P2_R2278_U163;
  assign new_P2_R2278_U408 = ~new_P2_R2278_U305 | ~new_P2_R2278_U406;
  assign new_P2_R2278_U409 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_R2278_U18;
  assign new_P2_R2278_U410 = ~new_P2_U3636 | ~new_P2_R2278_U19;
  assign new_P2_R2278_U411 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_R2278_U18;
  assign new_P2_R2278_U412 = ~new_P2_U3636 | ~new_P2_R2278_U19;
  assign new_P2_R2278_U413 = ~new_P2_R2278_U412 | ~new_P2_R2278_U411;
  assign new_P2_R2278_U414 = ~new_P2_R2278_U164 | ~new_P2_R2278_U165;
  assign new_P2_R2278_U415 = ~new_P2_R2278_U209 | ~new_P2_R2278_U413;
  assign new_P2_R2278_U416 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_R2278_U33;
  assign new_P2_R2278_U417 = ~new_P2_U2792 | ~new_P2_R2278_U34;
  assign new_P2_R2278_U418 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_R2278_U33;
  assign new_P2_R2278_U419 = ~new_P2_U2792 | ~new_P2_R2278_U34;
  assign new_P2_R2278_U420 = ~new_P2_R2278_U419 | ~new_P2_R2278_U418;
  assign new_P2_R2278_U421 = ~new_P2_R2278_U166 | ~new_P2_R2278_U167;
  assign new_P2_R2278_U422 = ~new_P2_R2278_U301 | ~new_P2_R2278_U420;
  assign new_P2_R2278_U423 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_R2278_U31;
  assign new_P2_R2278_U424 = ~new_P2_U2793 | ~new_P2_R2278_U32;
  assign new_P2_R2278_U425 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_R2278_U31;
  assign new_P2_R2278_U426 = ~new_P2_U2793 | ~new_P2_R2278_U32;
  assign new_P2_R2278_U427 = ~new_P2_R2278_U426 | ~new_P2_R2278_U425;
  assign new_P2_R2278_U428 = ~new_P2_R2278_U168 | ~new_P2_R2278_U169;
  assign new_P2_R2278_U429 = ~new_P2_R2278_U298 | ~new_P2_R2278_U427;
  assign new_P2_R2278_U430 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_R2278_U74;
  assign new_P2_R2278_U431 = ~new_P2_U2794 | ~new_P2_R2278_U75;
  assign new_P2_R2278_U432 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_R2278_U74;
  assign new_P2_R2278_U433 = ~new_P2_U2794 | ~new_P2_R2278_U75;
  assign new_P2_R2278_U434 = ~new_P2_R2278_U433 | ~new_P2_R2278_U432;
  assign new_P2_R2278_U435 = ~new_P2_R2278_U170 | ~new_P2_R2278_U171;
  assign new_P2_R2278_U436 = ~new_P2_R2278_U295 | ~new_P2_R2278_U434;
  assign new_P2_R2278_U437 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_R2278_U76;
  assign new_P2_R2278_U438 = ~new_P2_U2795 | ~new_P2_R2278_U77;
  assign new_P2_R2278_U439 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_R2278_U76;
  assign new_P2_R2278_U440 = ~new_P2_U2795 | ~new_P2_R2278_U77;
  assign new_P2_R2278_U441 = ~new_P2_R2278_U440 | ~new_P2_R2278_U439;
  assign new_P2_R2278_U442 = ~new_P2_R2278_U172 | ~new_P2_R2278_U173;
  assign new_P2_R2278_U443 = ~new_P2_R2278_U291 | ~new_P2_R2278_U441;
  assign new_P2_R2278_U444 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_R2278_U174;
  assign new_P2_R2278_U445 = ~new_P2_R2278_U289 | ~new_P2_R2278_U73;
  assign new_P2_R2278_U446 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_R2278_U174;
  assign new_P2_R2278_U447 = ~new_P2_R2278_U289 | ~new_P2_R2278_U73;
  assign new_P2_R2278_U448 = ~new_P2_R2278_U447 | ~new_P2_R2278_U446;
  assign new_P2_R2278_U449 = ~new_P2_R2278_U72 | ~new_P2_R2278_U445 | ~new_P2_R2278_U444;
  assign new_P2_R2278_U450 = ~new_P2_R2278_U448 | ~new_P2_U2796;
  assign new_P2_R2278_U451 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_R2278_U35;
  assign new_P2_R2278_U452 = ~new_P2_U2797 | ~new_P2_R2278_U36;
  assign new_P2_R2278_U453 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_R2278_U35;
  assign new_P2_R2278_U454 = ~new_P2_U2797 | ~new_P2_R2278_U36;
  assign new_P2_R2278_U455 = ~new_P2_R2278_U454 | ~new_P2_R2278_U453;
  assign new_P2_R2278_U456 = ~new_P2_R2278_U175 | ~new_P2_R2278_U176;
  assign new_P2_R2278_U457 = ~new_P2_R2278_U286 | ~new_P2_R2278_U455;
  assign new_P2_R2278_U458 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_R2278_U69;
  assign new_P2_R2278_U459 = ~new_P2_U2798 | ~new_P2_R2278_U70;
  assign new_P2_R2278_U460 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_R2278_U69;
  assign new_P2_R2278_U461 = ~new_P2_U2798 | ~new_P2_R2278_U70;
  assign new_P2_R2278_U462 = ~new_P2_R2278_U461 | ~new_P2_R2278_U460;
  assign new_P2_R2278_U463 = ~new_P2_R2278_U177 | ~new_P2_R2278_U178;
  assign new_P2_R2278_U464 = ~new_P2_R2278_U282 | ~new_P2_R2278_U462;
  assign new_P2_R2278_U465 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_R2278_U37;
  assign new_P2_R2278_U466 = ~new_P2_U2799 | ~new_P2_R2278_U38;
  assign new_P2_R2278_U467 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_R2278_U37;
  assign new_P2_R2278_U468 = ~new_P2_U2799 | ~new_P2_R2278_U38;
  assign new_P2_R2278_U469 = ~new_P2_R2278_U468 | ~new_P2_R2278_U467;
  assign new_P2_R2278_U470 = ~new_P2_R2278_U179 | ~new_P2_R2278_U180;
  assign new_P2_R2278_U471 = ~new_P2_R2278_U279 | ~new_P2_R2278_U469;
  assign new_P2_R2278_U472 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_R2278_U66;
  assign new_P2_R2278_U473 = ~new_P2_U2800 | ~new_P2_R2278_U67;
  assign new_P2_R2278_U474 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_R2278_U66;
  assign new_P2_R2278_U475 = ~new_P2_U2800 | ~new_P2_R2278_U67;
  assign new_P2_R2278_U476 = ~new_P2_R2278_U475 | ~new_P2_R2278_U474;
  assign new_P2_R2278_U477 = ~new_P2_R2278_U181 | ~new_P2_R2278_U182;
  assign new_P2_R2278_U478 = ~new_P2_R2278_U275 | ~new_P2_R2278_U476;
  assign new_P2_R2278_U479 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_R2278_U39;
  assign new_P2_R2278_U480 = ~new_P2_U2801 | ~new_P2_R2278_U40;
  assign new_P2_R2278_U481 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_R2278_U39;
  assign new_P2_R2278_U482 = ~new_P2_U2801 | ~new_P2_R2278_U40;
  assign new_P2_R2278_U483 = ~new_P2_R2278_U482 | ~new_P2_R2278_U481;
  assign new_P2_R2278_U484 = ~new_P2_R2278_U183 | ~new_P2_R2278_U184;
  assign new_P2_R2278_U485 = ~new_P2_R2278_U272 | ~new_P2_R2278_U483;
  assign new_P2_R2278_U486 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_R2278_U15;
  assign new_P2_R2278_U487 = ~new_P2_R2278_U208 | ~new_P2_R2278_U17;
  assign new_P2_R2278_U488 = ~new_P2_R2278_U487 | ~new_P2_R2278_U486;
  assign new_P2_R2278_U489 = ~new_P2_U3637 | ~new_P2_R2278_U15 | ~new_P2_R2278_U17;
  assign new_P2_R2278_U490 = ~new_P2_R2278_U488 | ~new_P2_R2278_U16;
  assign new_P2_R2278_U491 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_R2278_U62;
  assign new_P2_R2278_U492 = ~new_P2_U2802 | ~new_P2_R2278_U63;
  assign new_P2_R2278_U493 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_R2278_U62;
  assign new_P2_R2278_U494 = ~new_P2_U2802 | ~new_P2_R2278_U63;
  assign new_P2_R2278_U495 = ~new_P2_R2278_U494 | ~new_P2_R2278_U493;
  assign new_P2_R2278_U496 = ~new_P2_R2278_U185 | ~new_P2_R2278_U186;
  assign new_P2_R2278_U497 = ~new_P2_R2278_U269 | ~new_P2_R2278_U495;
  assign new_P2_R2278_U498 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_R2278_U64;
  assign new_P2_R2278_U499 = ~new_P2_U2803 | ~new_P2_R2278_U65;
  assign new_P2_R2278_U500 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_R2278_U64;
  assign new_P2_R2278_U501 = ~new_P2_U2803 | ~new_P2_R2278_U65;
  assign new_P2_R2278_U502 = ~new_P2_R2278_U501 | ~new_P2_R2278_U500;
  assign new_P2_R2278_U503 = ~new_P2_R2278_U187 | ~new_P2_R2278_U188;
  assign new_P2_R2278_U504 = ~new_P2_R2278_U265 | ~new_P2_R2278_U502;
  assign new_P2_R2278_U505 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_R2278_U41;
  assign new_P2_R2278_U506 = ~new_P2_U2804 | ~new_P2_R2278_U42;
  assign new_P2_R2278_U507 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_R2278_U41;
  assign new_P2_R2278_U508 = ~new_P2_U2804 | ~new_P2_R2278_U42;
  assign new_P2_R2278_U509 = ~new_P2_R2278_U508 | ~new_P2_R2278_U507;
  assign new_P2_R2278_U510 = ~new_P2_R2278_U189 | ~new_P2_R2278_U190;
  assign new_P2_R2278_U511 = ~new_P2_R2278_U262 | ~new_P2_R2278_U509;
  assign new_P2_R2278_U512 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_R2278_U59;
  assign new_P2_R2278_U513 = ~new_P2_U2805 | ~new_P2_R2278_U60;
  assign new_P2_R2278_U514 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_R2278_U59;
  assign new_P2_R2278_U515 = ~new_P2_U2805 | ~new_P2_R2278_U60;
  assign new_P2_R2278_U516 = ~new_P2_R2278_U515 | ~new_P2_R2278_U514;
  assign new_P2_R2278_U517 = ~new_P2_R2278_U191 | ~new_P2_R2278_U192;
  assign new_P2_R2278_U518 = ~new_P2_R2278_U258 | ~new_P2_R2278_U516;
  assign new_P2_R2278_U519 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_R2278_U43;
  assign new_P2_R2278_U520 = ~new_P2_U2806 | ~new_P2_R2278_U44;
  assign new_P2_R2278_U521 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_R2278_U43;
  assign new_P2_R2278_U522 = ~new_P2_U2806 | ~new_P2_R2278_U44;
  assign new_P2_R2278_U523 = ~new_P2_R2278_U522 | ~new_P2_R2278_U521;
  assign new_P2_R2278_U524 = ~new_P2_R2278_U193 | ~new_P2_R2278_U194;
  assign new_P2_R2278_U525 = ~new_P2_R2278_U255 | ~new_P2_R2278_U523;
  assign new_P2_R2278_U526 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_R2278_U56;
  assign new_P2_R2278_U527 = ~new_P2_U2807 | ~new_P2_R2278_U57;
  assign new_P2_R2278_U528 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_R2278_U56;
  assign new_P2_R2278_U529 = ~new_P2_U2807 | ~new_P2_R2278_U57;
  assign new_P2_R2278_U530 = ~new_P2_R2278_U529 | ~new_P2_R2278_U528;
  assign new_P2_R2278_U531 = ~new_P2_R2278_U195 | ~new_P2_R2278_U196;
  assign new_P2_R2278_U532 = ~new_P2_R2278_U251 | ~new_P2_R2278_U530;
  assign new_P2_R2278_U533 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_R2278_U45;
  assign new_P2_R2278_U534 = ~new_P2_U2808 | ~new_P2_R2278_U46;
  assign new_P2_R2278_U535 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_R2278_U45;
  assign new_P2_R2278_U536 = ~new_P2_U2808 | ~new_P2_R2278_U46;
  assign new_P2_R2278_U537 = ~new_P2_R2278_U536 | ~new_P2_R2278_U535;
  assign new_P2_R2278_U538 = ~new_P2_R2278_U197 | ~new_P2_R2278_U198;
  assign new_P2_R2278_U539 = ~new_P2_R2278_U248 | ~new_P2_R2278_U537;
  assign new_P2_R2278_U540 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_R2278_U53;
  assign new_P2_R2278_U541 = ~new_P2_U2809 | ~new_P2_R2278_U54;
  assign new_P2_R2278_U542 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_R2278_U53;
  assign new_P2_R2278_U543 = ~new_P2_U2809 | ~new_P2_R2278_U54;
  assign new_P2_R2278_U544 = ~new_P2_R2278_U543 | ~new_P2_R2278_U542;
  assign new_P2_R2278_U545 = ~new_P2_R2278_U199 | ~new_P2_R2278_U200;
  assign new_P2_R2278_U546 = ~new_P2_R2278_U244 | ~new_P2_R2278_U544;
  assign new_P2_R2278_U547 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_R2278_U47;
  assign new_P2_R2278_U548 = ~new_P2_U2810 | ~new_P2_R2278_U48;
  assign new_P2_R2278_U549 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_R2278_U47;
  assign new_P2_R2278_U550 = ~new_P2_U2810 | ~new_P2_R2278_U48;
  assign new_P2_R2278_U551 = ~new_P2_R2278_U550 | ~new_P2_R2278_U549;
  assign new_P2_R2278_U552 = ~new_P2_R2278_U201 | ~new_P2_R2278_U202;
  assign new_P2_R2278_U553 = ~new_P2_R2278_U241 | ~new_P2_R2278_U551;
  assign new_P2_R2278_U554 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_R2278_U50;
  assign new_P2_R2278_U555 = ~new_P2_U2811 | ~new_P2_R2278_U51;
  assign new_P2_R2278_U556 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_R2278_U50;
  assign new_P2_R2278_U557 = ~new_P2_U2811 | ~new_P2_R2278_U51;
  assign new_P2_R2278_U558 = ~new_P2_R2278_U557 | ~new_P2_R2278_U556;
  assign new_P2_R2278_U559 = ~new_P2_R2278_U203 | ~new_P2_R2278_U204;
  assign new_P2_R2278_U560 = ~new_P2_R2278_U237 | ~new_P2_R2278_U558;
  assign new_P2_R2278_U561 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_R2278_U13;
  assign new_P2_R2278_U562 = ~new_P2_U3638 | ~new_P2_R2278_U14;
  assign new_P2_SUB_450_U6 = ~new_P2_SUB_450_U43 | ~new_P2_SUB_450_U42;
  assign new_P2_SUB_450_U7 = ~P2_INSTQUEUERD_ADDR_REG_0_ | ~new_P2_SUB_450_U16;
  assign new_P2_SUB_450_U8 = ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P2_SUB_450_U9 = ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign new_P2_SUB_450_U10 = ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P2_SUB_450_U11 = ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign new_P2_SUB_450_U12 = ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P2_SUB_450_U13 = ~P2_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P2_SUB_450_U14 = ~new_P2_SUB_450_U39 | ~new_P2_SUB_450_U38;
  assign new_P2_SUB_450_U15 = ~P2_INSTQUEUERD_ADDR_REG_4_;
  assign new_P2_SUB_450_U16 = ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P2_SUB_450_U17 = ~new_P2_SUB_450_U48 | ~new_P2_SUB_450_U47;
  assign new_P2_SUB_450_U18 = ~new_P2_SUB_450_U53 | ~new_P2_SUB_450_U52;
  assign new_P2_SUB_450_U19 = ~new_P2_SUB_450_U58 | ~new_P2_SUB_450_U57;
  assign new_P2_SUB_450_U20 = ~new_P2_SUB_450_U63 | ~new_P2_SUB_450_U62;
  assign new_P2_SUB_450_U21 = ~new_P2_SUB_450_U45 | ~new_P2_SUB_450_U44;
  assign new_P2_SUB_450_U22 = ~new_P2_SUB_450_U50 | ~new_P2_SUB_450_U49;
  assign new_P2_SUB_450_U23 = ~new_P2_SUB_450_U55 | ~new_P2_SUB_450_U54;
  assign new_P2_SUB_450_U24 = ~new_P2_SUB_450_U60 | ~new_P2_SUB_450_U59;
  assign new_P2_SUB_450_U25 = ~new_P2_SUB_450_U35 | ~new_P2_SUB_450_U34;
  assign new_P2_SUB_450_U26 = ~new_P2_SUB_450_U31 | ~new_P2_SUB_450_U30;
  assign new_P2_SUB_450_U27 = ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign new_P2_SUB_450_U28 = ~new_P2_SUB_450_U7;
  assign new_P2_SUB_450_U29 = ~new_P2_SUB_450_U28 | ~new_P2_SUB_450_U8;
  assign new_P2_SUB_450_U30 = ~new_P2_SUB_450_U29 | ~new_P2_SUB_450_U27;
  assign new_P2_SUB_450_U31 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_SUB_450_U7;
  assign new_P2_SUB_450_U32 = ~new_P2_SUB_450_U26;
  assign new_P2_SUB_450_U33 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_SUB_450_U10;
  assign new_P2_SUB_450_U34 = ~new_P2_SUB_450_U33 | ~new_P2_SUB_450_U26;
  assign new_P2_SUB_450_U35 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_SUB_450_U9;
  assign new_P2_SUB_450_U36 = ~new_P2_SUB_450_U25;
  assign new_P2_SUB_450_U37 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_SUB_450_U12;
  assign new_P2_SUB_450_U38 = ~new_P2_SUB_450_U37 | ~new_P2_SUB_450_U25;
  assign new_P2_SUB_450_U39 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_SUB_450_U11;
  assign new_P2_SUB_450_U40 = ~new_P2_SUB_450_U14;
  assign new_P2_SUB_450_U41 = ~P2_INSTQUEUEWR_ADDR_REG_4_ | ~new_P2_SUB_450_U15;
  assign new_P2_SUB_450_U42 = ~new_P2_SUB_450_U40 | ~new_P2_SUB_450_U41;
  assign new_P2_SUB_450_U43 = ~P2_INSTQUEUERD_ADDR_REG_4_ | ~new_P2_SUB_450_U13;
  assign new_P2_SUB_450_U44 = ~P2_INSTQUEUERD_ADDR_REG_4_ | ~new_P2_SUB_450_U13;
  assign new_P2_SUB_450_U45 = ~P2_INSTQUEUEWR_ADDR_REG_4_ | ~new_P2_SUB_450_U15;
  assign new_P2_SUB_450_U46 = ~new_P2_SUB_450_U21;
  assign new_P2_SUB_450_U47 = ~new_P2_SUB_450_U46 | ~new_P2_SUB_450_U40;
  assign new_P2_SUB_450_U48 = ~new_P2_SUB_450_U21 | ~new_P2_SUB_450_U14;
  assign new_P2_SUB_450_U49 = ~P2_INSTQUEUERD_ADDR_REG_3_ | ~new_P2_SUB_450_U12;
  assign new_P2_SUB_450_U50 = ~P2_INSTQUEUEWR_ADDR_REG_3_ | ~new_P2_SUB_450_U11;
  assign new_P2_SUB_450_U51 = ~new_P2_SUB_450_U22;
  assign new_P2_SUB_450_U52 = ~new_P2_SUB_450_U36 | ~new_P2_SUB_450_U51;
  assign new_P2_SUB_450_U53 = ~new_P2_SUB_450_U22 | ~new_P2_SUB_450_U25;
  assign new_P2_SUB_450_U54 = ~P2_INSTQUEUERD_ADDR_REG_2_ | ~new_P2_SUB_450_U10;
  assign new_P2_SUB_450_U55 = ~P2_INSTQUEUEWR_ADDR_REG_2_ | ~new_P2_SUB_450_U9;
  assign new_P2_SUB_450_U56 = ~new_P2_SUB_450_U23;
  assign new_P2_SUB_450_U57 = ~new_P2_SUB_450_U32 | ~new_P2_SUB_450_U56;
  assign new_P2_SUB_450_U58 = ~new_P2_SUB_450_U23 | ~new_P2_SUB_450_U26;
  assign new_P2_SUB_450_U59 = ~P2_INSTQUEUERD_ADDR_REG_1_ | ~new_P2_SUB_450_U8;
  assign new_P2_SUB_450_U60 = ~P2_INSTQUEUEWR_ADDR_REG_1_ | ~new_P2_SUB_450_U27;
  assign new_P2_SUB_450_U61 = ~new_P2_SUB_450_U24;
  assign new_P2_SUB_450_U62 = ~new_P2_SUB_450_U61 | ~new_P2_SUB_450_U28;
  assign new_P2_SUB_450_U63 = ~new_P2_SUB_450_U24 | ~new_P2_SUB_450_U7;
  assign new_P2_R2088_U6 = ~new_P2_U3648 & ~new_P2_R2088_U7;
  assign new_P2_R2088_U7 = ~new_P2_U3651 & ~new_P2_U3652 & ~new_P2_U3650 & ~new_P2_U3648 & ~new_P2_U3649;
  assign new_P2_ADD_394_U4 = ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_ADD_394_U5 = ~new_P2_ADD_394_U94 | ~new_P2_ADD_394_U125;
  assign new_P2_ADD_394_U6 = ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_ADD_394_U7 = ~P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_ADD_394_U8 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_ADD_394_U94;
  assign new_P2_ADD_394_U9 = ~P2_INSTADDRPOINTER_REG_4_;
  assign new_P2_ADD_394_U10 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_ADD_394_U98;
  assign new_P2_ADD_394_U11 = ~P2_INSTADDRPOINTER_REG_5_;
  assign new_P2_ADD_394_U12 = ~P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_ADD_394_U13 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_ADD_394_U99;
  assign new_P2_ADD_394_U14 = ~new_P2_ADD_394_U100 | ~P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_ADD_394_U15 = ~P2_INSTADDRPOINTER_REG_7_;
  assign new_P2_ADD_394_U16 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_ADD_394_U101;
  assign new_P2_ADD_394_U17 = ~P2_INSTADDRPOINTER_REG_8_;
  assign new_P2_ADD_394_U18 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_ADD_394_U102;
  assign new_P2_ADD_394_U19 = ~P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_ADD_394_U20 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_ADD_394_U103;
  assign new_P2_ADD_394_U21 = ~P2_INSTADDRPOINTER_REG_10_;
  assign new_P2_ADD_394_U22 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_ADD_394_U104;
  assign new_P2_ADD_394_U23 = ~P2_INSTADDRPOINTER_REG_11_;
  assign new_P2_ADD_394_U24 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_ADD_394_U105;
  assign new_P2_ADD_394_U25 = ~P2_INSTADDRPOINTER_REG_12_;
  assign new_P2_ADD_394_U26 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_ADD_394_U106;
  assign new_P2_ADD_394_U27 = ~P2_INSTADDRPOINTER_REG_13_;
  assign new_P2_ADD_394_U28 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_ADD_394_U107;
  assign new_P2_ADD_394_U29 = ~P2_INSTADDRPOINTER_REG_14_;
  assign new_P2_ADD_394_U30 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_ADD_394_U108;
  assign new_P2_ADD_394_U31 = ~P2_INSTADDRPOINTER_REG_15_;
  assign new_P2_ADD_394_U32 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_ADD_394_U109;
  assign new_P2_ADD_394_U33 = ~P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_ADD_394_U34 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_ADD_394_U110;
  assign new_P2_ADD_394_U35 = ~P2_INSTADDRPOINTER_REG_17_;
  assign new_P2_ADD_394_U36 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_ADD_394_U111;
  assign new_P2_ADD_394_U37 = ~P2_INSTADDRPOINTER_REG_18_;
  assign new_P2_ADD_394_U38 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_ADD_394_U112;
  assign new_P2_ADD_394_U39 = ~P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_ADD_394_U40 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_ADD_394_U113;
  assign new_P2_ADD_394_U41 = ~P2_INSTADDRPOINTER_REG_20_;
  assign new_P2_ADD_394_U42 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_ADD_394_U114;
  assign new_P2_ADD_394_U43 = ~P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_ADD_394_U44 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_ADD_394_U115;
  assign new_P2_ADD_394_U45 = ~P2_INSTADDRPOINTER_REG_22_;
  assign new_P2_ADD_394_U46 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_ADD_394_U116;
  assign new_P2_ADD_394_U47 = ~P2_INSTADDRPOINTER_REG_23_;
  assign new_P2_ADD_394_U48 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_ADD_394_U117;
  assign new_P2_ADD_394_U49 = ~P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_ADD_394_U50 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_ADD_394_U118;
  assign new_P2_ADD_394_U51 = ~P2_INSTADDRPOINTER_REG_25_;
  assign new_P2_ADD_394_U52 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_ADD_394_U119;
  assign new_P2_ADD_394_U53 = ~P2_INSTADDRPOINTER_REG_26_;
  assign new_P2_ADD_394_U54 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_ADD_394_U120;
  assign new_P2_ADD_394_U55 = ~P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_ADD_394_U56 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_ADD_394_U121;
  assign new_P2_ADD_394_U57 = ~P2_INSTADDRPOINTER_REG_28_;
  assign new_P2_ADD_394_U58 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_ADD_394_U122;
  assign new_P2_ADD_394_U59 = ~P2_INSTADDRPOINTER_REG_29_;
  assign new_P2_ADD_394_U60 = ~P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_ADD_394_U61 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_ADD_394_U123;
  assign new_P2_ADD_394_U62 = ~P2_INSTADDRPOINTER_REG_2_;
  assign new_P2_ADD_394_U63 = ~new_P2_ADD_394_U128 | ~new_P2_ADD_394_U127;
  assign new_P2_ADD_394_U64 = ~new_P2_ADD_394_U130 | ~new_P2_ADD_394_U129;
  assign new_P2_ADD_394_U65 = ~new_P2_ADD_394_U132 | ~new_P2_ADD_394_U131;
  assign new_P2_ADD_394_U66 = ~new_P2_ADD_394_U134 | ~new_P2_ADD_394_U133;
  assign new_P2_ADD_394_U67 = ~new_P2_ADD_394_U136 | ~new_P2_ADD_394_U135;
  assign new_P2_ADD_394_U68 = ~new_P2_ADD_394_U138 | ~new_P2_ADD_394_U137;
  assign new_P2_ADD_394_U69 = ~new_P2_ADD_394_U140 | ~new_P2_ADD_394_U139;
  assign new_P2_ADD_394_U70 = ~new_P2_ADD_394_U142 | ~new_P2_ADD_394_U141;
  assign new_P2_ADD_394_U71 = ~new_P2_ADD_394_U144 | ~new_P2_ADD_394_U143;
  assign new_P2_ADD_394_U72 = ~new_P2_ADD_394_U146 | ~new_P2_ADD_394_U145;
  assign new_P2_ADD_394_U73 = ~new_P2_ADD_394_U148 | ~new_P2_ADD_394_U147;
  assign new_P2_ADD_394_U74 = ~new_P2_ADD_394_U150 | ~new_P2_ADD_394_U149;
  assign new_P2_ADD_394_U75 = ~new_P2_ADD_394_U152 | ~new_P2_ADD_394_U151;
  assign new_P2_ADD_394_U76 = ~new_P2_ADD_394_U154 | ~new_P2_ADD_394_U153;
  assign new_P2_ADD_394_U77 = ~new_P2_ADD_394_U156 | ~new_P2_ADD_394_U155;
  assign new_P2_ADD_394_U78 = ~new_P2_ADD_394_U158 | ~new_P2_ADD_394_U157;
  assign new_P2_ADD_394_U79 = ~new_P2_ADD_394_U160 | ~new_P2_ADD_394_U159;
  assign new_P2_ADD_394_U80 = ~new_P2_ADD_394_U162 | ~new_P2_ADD_394_U161;
  assign new_P2_ADD_394_U81 = ~new_P2_ADD_394_U164 | ~new_P2_ADD_394_U163;
  assign new_P2_ADD_394_U82 = ~new_P2_ADD_394_U166 | ~new_P2_ADD_394_U165;
  assign new_P2_ADD_394_U83 = ~new_P2_ADD_394_U168 | ~new_P2_ADD_394_U167;
  assign new_P2_ADD_394_U84 = ~new_P2_ADD_394_U170 | ~new_P2_ADD_394_U169;
  assign new_P2_ADD_394_U85 = ~new_P2_ADD_394_U174 | ~new_P2_ADD_394_U173;
  assign new_P2_ADD_394_U86 = ~new_P2_ADD_394_U176 | ~new_P2_ADD_394_U175;
  assign new_P2_ADD_394_U87 = ~new_P2_ADD_394_U178 | ~new_P2_ADD_394_U177;
  assign new_P2_ADD_394_U88 = ~new_P2_ADD_394_U180 | ~new_P2_ADD_394_U179;
  assign new_P2_ADD_394_U89 = ~new_P2_ADD_394_U182 | ~new_P2_ADD_394_U181;
  assign new_P2_ADD_394_U90 = ~new_P2_ADD_394_U184 | ~new_P2_ADD_394_U183;
  assign new_P2_ADD_394_U91 = ~new_P2_ADD_394_U186 | ~new_P2_ADD_394_U185;
  assign new_P2_ADD_394_U92 = ~P2_INSTADDRPOINTER_REG_31_;
  assign new_P2_ADD_394_U93 = ~new_P2_ADD_394_U124 | ~P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_ADD_394_U94 = ~new_P2_ADD_394_U62 | ~new_P2_ADD_394_U96;
  assign new_P2_ADD_394_U95 = new_P2_ADD_394_U172 & new_P2_ADD_394_U171;
  assign new_P2_ADD_394_U96 = ~P2_INSTADDRPOINTER_REG_1_ | ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_ADD_394_U97 = ~new_P2_ADD_394_U94;
  assign new_P2_ADD_394_U98 = ~new_P2_ADD_394_U8;
  assign new_P2_ADD_394_U99 = ~new_P2_ADD_394_U10;
  assign new_P2_ADD_394_U100 = ~new_P2_ADD_394_U13;
  assign new_P2_ADD_394_U101 = ~new_P2_ADD_394_U14;
  assign new_P2_ADD_394_U102 = ~new_P2_ADD_394_U16;
  assign new_P2_ADD_394_U103 = ~new_P2_ADD_394_U18;
  assign new_P2_ADD_394_U104 = ~new_P2_ADD_394_U20;
  assign new_P2_ADD_394_U105 = ~new_P2_ADD_394_U22;
  assign new_P2_ADD_394_U106 = ~new_P2_ADD_394_U24;
  assign new_P2_ADD_394_U107 = ~new_P2_ADD_394_U26;
  assign new_P2_ADD_394_U108 = ~new_P2_ADD_394_U28;
  assign new_P2_ADD_394_U109 = ~new_P2_ADD_394_U30;
  assign new_P2_ADD_394_U110 = ~new_P2_ADD_394_U32;
  assign new_P2_ADD_394_U111 = ~new_P2_ADD_394_U34;
  assign new_P2_ADD_394_U112 = ~new_P2_ADD_394_U36;
  assign new_P2_ADD_394_U113 = ~new_P2_ADD_394_U38;
  assign new_P2_ADD_394_U114 = ~new_P2_ADD_394_U40;
  assign new_P2_ADD_394_U115 = ~new_P2_ADD_394_U42;
  assign new_P2_ADD_394_U116 = ~new_P2_ADD_394_U44;
  assign new_P2_ADD_394_U117 = ~new_P2_ADD_394_U46;
  assign new_P2_ADD_394_U118 = ~new_P2_ADD_394_U48;
  assign new_P2_ADD_394_U119 = ~new_P2_ADD_394_U50;
  assign new_P2_ADD_394_U120 = ~new_P2_ADD_394_U52;
  assign new_P2_ADD_394_U121 = ~new_P2_ADD_394_U54;
  assign new_P2_ADD_394_U122 = ~new_P2_ADD_394_U56;
  assign new_P2_ADD_394_U123 = ~new_P2_ADD_394_U58;
  assign new_P2_ADD_394_U124 = ~new_P2_ADD_394_U61;
  assign new_P2_ADD_394_U125 = ~P2_INSTADDRPOINTER_REG_2_ | ~P2_INSTADDRPOINTER_REG_1_ | ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_ADD_394_U126 = ~new_P2_ADD_394_U93;
  assign new_P2_ADD_394_U127 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_ADD_394_U13;
  assign new_P2_ADD_394_U128 = ~new_P2_ADD_394_U100 | ~new_P2_ADD_394_U12;
  assign new_P2_ADD_394_U129 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_ADD_394_U61;
  assign new_P2_ADD_394_U130 = ~new_P2_ADD_394_U124 | ~new_P2_ADD_394_U60;
  assign new_P2_ADD_394_U131 = ~P2_INSTADDRPOINTER_REG_29_ | ~new_P2_ADD_394_U58;
  assign new_P2_ADD_394_U132 = ~new_P2_ADD_394_U123 | ~new_P2_ADD_394_U59;
  assign new_P2_ADD_394_U133 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_ADD_394_U48;
  assign new_P2_ADD_394_U134 = ~new_P2_ADD_394_U118 | ~new_P2_ADD_394_U49;
  assign new_P2_ADD_394_U135 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_ADD_394_U34;
  assign new_P2_ADD_394_U136 = ~new_P2_ADD_394_U111 | ~new_P2_ADD_394_U35;
  assign new_P2_ADD_394_U137 = ~P2_INSTADDRPOINTER_REG_20_ | ~new_P2_ADD_394_U40;
  assign new_P2_ADD_394_U138 = ~new_P2_ADD_394_U114 | ~new_P2_ADD_394_U41;
  assign new_P2_ADD_394_U139 = ~P2_INSTADDRPOINTER_REG_13_ | ~new_P2_ADD_394_U26;
  assign new_P2_ADD_394_U140 = ~new_P2_ADD_394_U107 | ~new_P2_ADD_394_U27;
  assign new_P2_ADD_394_U141 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_ADD_394_U18;
  assign new_P2_ADD_394_U142 = ~new_P2_ADD_394_U103 | ~new_P2_ADD_394_U19;
  assign new_P2_ADD_394_U143 = ~P2_INSTADDRPOINTER_REG_22_ | ~new_P2_ADD_394_U44;
  assign new_P2_ADD_394_U144 = ~new_P2_ADD_394_U116 | ~new_P2_ADD_394_U45;
  assign new_P2_ADD_394_U145 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_ADD_394_U36;
  assign new_P2_ADD_394_U146 = ~new_P2_ADD_394_U112 | ~new_P2_ADD_394_U37;
  assign new_P2_ADD_394_U147 = ~P2_INSTADDRPOINTER_REG_11_ | ~new_P2_ADD_394_U22;
  assign new_P2_ADD_394_U148 = ~new_P2_ADD_394_U105 | ~new_P2_ADD_394_U23;
  assign new_P2_ADD_394_U149 = ~P2_INSTADDRPOINTER_REG_26_ | ~new_P2_ADD_394_U52;
  assign new_P2_ADD_394_U150 = ~new_P2_ADD_394_U120 | ~new_P2_ADD_394_U53;
  assign new_P2_ADD_394_U151 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_ADD_394_U30;
  assign new_P2_ADD_394_U152 = ~new_P2_ADD_394_U109 | ~new_P2_ADD_394_U31;
  assign new_P2_ADD_394_U153 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_ADD_394_U8;
  assign new_P2_ADD_394_U154 = ~new_P2_ADD_394_U98 | ~new_P2_ADD_394_U9;
  assign new_P2_ADD_394_U155 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_ADD_394_U54;
  assign new_P2_ADD_394_U156 = ~new_P2_ADD_394_U121 | ~new_P2_ADD_394_U55;
  assign new_P2_ADD_394_U157 = ~P2_INSTADDRPOINTER_REG_14_ | ~new_P2_ADD_394_U28;
  assign new_P2_ADD_394_U158 = ~new_P2_ADD_394_U108 | ~new_P2_ADD_394_U29;
  assign new_P2_ADD_394_U159 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_ADD_394_U10;
  assign new_P2_ADD_394_U160 = ~new_P2_ADD_394_U99 | ~new_P2_ADD_394_U11;
  assign new_P2_ADD_394_U161 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_ADD_394_U16;
  assign new_P2_ADD_394_U162 = ~new_P2_ADD_394_U102 | ~new_P2_ADD_394_U17;
  assign new_P2_ADD_394_U163 = ~P2_INSTADDRPOINTER_REG_23_ | ~new_P2_ADD_394_U46;
  assign new_P2_ADD_394_U164 = ~new_P2_ADD_394_U117 | ~new_P2_ADD_394_U47;
  assign new_P2_ADD_394_U165 = ~P2_INSTADDRPOINTER_REG_19_ | ~new_P2_ADD_394_U38;
  assign new_P2_ADD_394_U166 = ~new_P2_ADD_394_U113 | ~new_P2_ADD_394_U39;
  assign new_P2_ADD_394_U167 = ~P2_INSTADDRPOINTER_REG_10_ | ~new_P2_ADD_394_U20;
  assign new_P2_ADD_394_U168 = ~new_P2_ADD_394_U104 | ~new_P2_ADD_394_U21;
  assign new_P2_ADD_394_U169 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_ADD_394_U93;
  assign new_P2_ADD_394_U170 = ~new_P2_ADD_394_U126 | ~new_P2_ADD_394_U92;
  assign new_P2_ADD_394_U171 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_ADD_394_U94;
  assign new_P2_ADD_394_U172 = ~new_P2_ADD_394_U97 | ~new_P2_ADD_394_U7;
  assign new_P2_ADD_394_U173 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_ADD_394_U4;
  assign new_P2_ADD_394_U174 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_ADD_394_U6;
  assign new_P2_ADD_394_U175 = ~P2_INSTADDRPOINTER_REG_28_ | ~new_P2_ADD_394_U56;
  assign new_P2_ADD_394_U176 = ~new_P2_ADD_394_U122 | ~new_P2_ADD_394_U57;
  assign new_P2_ADD_394_U177 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_ADD_394_U42;
  assign new_P2_ADD_394_U178 = ~new_P2_ADD_394_U115 | ~new_P2_ADD_394_U43;
  assign new_P2_ADD_394_U179 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_ADD_394_U24;
  assign new_P2_ADD_394_U180 = ~new_P2_ADD_394_U106 | ~new_P2_ADD_394_U25;
  assign new_P2_ADD_394_U181 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_ADD_394_U14;
  assign new_P2_ADD_394_U182 = ~new_P2_ADD_394_U101 | ~new_P2_ADD_394_U15;
  assign new_P2_ADD_394_U183 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_ADD_394_U50;
  assign new_P2_ADD_394_U184 = ~new_P2_ADD_394_U119 | ~new_P2_ADD_394_U51;
  assign new_P2_ADD_394_U185 = ~P2_INSTADDRPOINTER_REG_16_ | ~new_P2_ADD_394_U32;
  assign new_P2_ADD_394_U186 = ~new_P2_ADD_394_U110 | ~new_P2_ADD_394_U33;
  assign new_P2_R2267_U6 = new_P2_R2267_U133 & new_P2_R2267_U31;
  assign new_P2_R2267_U7 = new_P2_R2267_U131 & new_P2_R2267_U32;
  assign new_P2_R2267_U8 = new_P2_R2267_U129 & new_P2_R2267_U33;
  assign new_P2_R2267_U9 = new_P2_R2267_U127 & new_P2_R2267_U34;
  assign new_P2_R2267_U10 = new_P2_R2267_U125 & new_P2_R2267_U35;
  assign new_P2_R2267_U11 = new_P2_R2267_U123 & new_P2_R2267_U36;
  assign new_P2_R2267_U12 = new_P2_R2267_U121 & new_P2_R2267_U37;
  assign new_P2_R2267_U13 = new_P2_R2267_U119 & new_P2_R2267_U38;
  assign new_P2_R2267_U14 = new_P2_R2267_U117 & new_P2_R2267_U39;
  assign new_P2_R2267_U15 = new_P2_R2267_U115 & new_P2_R2267_U40;
  assign new_P2_R2267_U16 = new_P2_R2267_U113 & new_P2_R2267_U62;
  assign new_P2_R2267_U17 = new_P2_R2267_U101 & new_P2_R2267_U24;
  assign new_P2_R2267_U18 = new_P2_R2267_U99 & new_P2_R2267_U25;
  assign new_P2_R2267_U19 = new_P2_R2267_U97 & new_P2_R2267_U26;
  assign new_P2_R2267_U20 = new_P2_R2267_U95 & new_P2_R2267_U30;
  assign new_P2_R2267_U21 = ~new_P2_R2267_U77 | ~new_P2_R2267_U134;
  assign new_P2_R2267_U22 = ~new_P2_U3646;
  assign new_P2_R2267_U23 = ~new_P2_R2267_U76 | ~new_P2_R2267_U77;
  assign new_P2_R2267_U24 = ~new_P2_R2267_U29 | ~new_P2_R2267_U89 | ~new_P2_R2267_U64;
  assign new_P2_R2267_U25 = ~new_P2_R2267_U28 | ~new_P2_R2267_U90 | ~new_P2_R2267_U59;
  assign new_P2_R2267_U26 = ~new_P2_R2267_U27 | ~new_P2_R2267_U91 | ~new_P2_R2267_U57;
  assign new_P2_R2267_U27 = ~new_P2_U3639;
  assign new_P2_R2267_U28 = ~new_P2_U3641;
  assign new_P2_R2267_U29 = ~new_P2_U3643;
  assign new_P2_R2267_U30 = ~new_P2_R2267_U44 | ~new_P2_R2267_U92;
  assign new_P2_R2267_U31 = ~new_P2_R2267_U45 | ~new_P2_R2267_U93;
  assign new_P2_R2267_U32 = ~new_P2_R2267_U46 | ~new_P2_R2267_U102;
  assign new_P2_R2267_U33 = ~new_P2_R2267_U47 | ~new_P2_R2267_U103;
  assign new_P2_R2267_U34 = ~new_P2_R2267_U48 | ~new_P2_R2267_U104;
  assign new_P2_R2267_U35 = ~new_P2_R2267_U49 | ~new_P2_R2267_U105;
  assign new_P2_R2267_U36 = ~new_P2_R2267_U50 | ~new_P2_R2267_U106;
  assign new_P2_R2267_U37 = ~new_P2_R2267_U51 | ~new_P2_R2267_U107;
  assign new_P2_R2267_U38 = ~new_P2_R2267_U52 | ~new_P2_R2267_U108;
  assign new_P2_R2267_U39 = ~new_P2_R2267_U53 | ~new_P2_R2267_U109;
  assign new_P2_R2267_U40 = ~new_P2_R2267_U54 | ~new_P2_R2267_U110;
  assign new_P2_R2267_U41 = ~new_P2_U2767;
  assign new_P2_R2267_U42 = ~new_P2_U2617;
  assign new_P2_R2267_U43 = ~new_P2_R2267_U156 | ~new_P2_R2267_U155;
  assign new_P2_R2267_U44 = ~new_P2_U2789 & ~new_P2_U2788;
  assign new_P2_R2267_U45 = ~new_P2_U2787 & ~new_P2_U2786;
  assign new_P2_R2267_U46 = ~new_P2_U2785 & ~new_P2_U2784;
  assign new_P2_R2267_U47 = ~new_P2_U2783 & ~new_P2_U2782;
  assign new_P2_R2267_U48 = ~new_P2_U2781 & ~new_P2_U2780;
  assign new_P2_R2267_U49 = ~new_P2_U2779 & ~new_P2_U2778;
  assign new_P2_R2267_U50 = ~new_P2_U2777 & ~new_P2_U2776;
  assign new_P2_R2267_U51 = ~new_P2_U2775 & ~new_P2_U2774;
  assign new_P2_R2267_U52 = ~new_P2_U2773 & ~new_P2_U2772;
  assign new_P2_R2267_U53 = ~new_P2_U2771 & ~new_P2_U2770;
  assign new_P2_R2267_U54 = ~new_P2_U2769 & ~new_P2_U2768;
  assign new_P2_R2267_U55 = ~new_P2_U2789;
  assign new_P2_R2267_U56 = new_P2_R2267_U136 & new_P2_R2267_U135;
  assign new_P2_R2267_U57 = ~new_P2_U3640;
  assign new_P2_R2267_U58 = new_P2_R2267_U138 & new_P2_R2267_U137;
  assign new_P2_R2267_U59 = ~new_P2_U3642;
  assign new_P2_R2267_U60 = new_P2_R2267_U140 & new_P2_R2267_U139;
  assign new_P2_R2267_U61 = ~new_P2_U2766;
  assign new_P2_R2267_U62 = ~new_P2_R2267_U111 | ~new_P2_R2267_U41;
  assign new_P2_R2267_U63 = new_P2_R2267_U142 & new_P2_R2267_U141;
  assign new_P2_R2267_U64 = ~new_P2_U3644;
  assign new_P2_R2267_U65 = new_P2_R2267_U144 & new_P2_R2267_U143;
  assign new_P2_R2267_U66 = ~new_P2_U2769;
  assign new_P2_R2267_U67 = new_P2_R2267_U146 & new_P2_R2267_U145;
  assign new_P2_R2267_U68 = ~new_P2_U2771;
  assign new_P2_R2267_U69 = new_P2_R2267_U148 & new_P2_R2267_U147;
  assign new_P2_R2267_U70 = ~new_P2_U2773;
  assign new_P2_R2267_U71 = new_P2_R2267_U150 & new_P2_R2267_U149;
  assign new_P2_R2267_U72 = ~new_P2_U2775;
  assign new_P2_R2267_U73 = new_P2_R2267_U152 & new_P2_R2267_U151;
  assign new_P2_R2267_U74 = ~new_P2_U2777;
  assign new_P2_R2267_U75 = new_P2_R2267_U154 & new_P2_R2267_U153;
  assign new_P2_R2267_U76 = ~new_P2_U3645;
  assign new_P2_R2267_U77 = ~new_P2_U3646 | ~new_P2_R2267_U42;
  assign new_P2_R2267_U78 = ~new_P2_U2779;
  assign new_P2_R2267_U79 = new_P2_R2267_U158 & new_P2_R2267_U157;
  assign new_P2_R2267_U80 = ~new_P2_U2781;
  assign new_P2_R2267_U81 = new_P2_R2267_U160 & new_P2_R2267_U159;
  assign new_P2_R2267_U82 = ~new_P2_U2783;
  assign new_P2_R2267_U83 = new_P2_R2267_U162 & new_P2_R2267_U161;
  assign new_P2_R2267_U84 = ~new_P2_U2785;
  assign new_P2_R2267_U85 = new_P2_R2267_U164 & new_P2_R2267_U163;
  assign new_P2_R2267_U86 = ~new_P2_U2787;
  assign new_P2_R2267_U87 = new_P2_R2267_U166 & new_P2_R2267_U165;
  assign new_P2_R2267_U88 = ~new_P2_R2267_U77;
  assign new_P2_R2267_U89 = ~new_P2_R2267_U23;
  assign new_P2_R2267_U90 = ~new_P2_R2267_U24;
  assign new_P2_R2267_U91 = ~new_P2_R2267_U25;
  assign new_P2_R2267_U92 = ~new_P2_R2267_U26;
  assign new_P2_R2267_U93 = ~new_P2_R2267_U30;
  assign new_P2_R2267_U94 = ~new_P2_R2267_U92 | ~new_P2_R2267_U55;
  assign new_P2_R2267_U95 = ~new_P2_U2788 | ~new_P2_R2267_U94;
  assign new_P2_R2267_U96 = ~new_P2_R2267_U91 | ~new_P2_R2267_U57;
  assign new_P2_R2267_U97 = ~new_P2_U3639 | ~new_P2_R2267_U96;
  assign new_P2_R2267_U98 = ~new_P2_R2267_U90 | ~new_P2_R2267_U59;
  assign new_P2_R2267_U99 = ~new_P2_U3641 | ~new_P2_R2267_U98;
  assign new_P2_R2267_U100 = ~new_P2_R2267_U89 | ~new_P2_R2267_U64;
  assign new_P2_R2267_U101 = ~new_P2_U3643 | ~new_P2_R2267_U100;
  assign new_P2_R2267_U102 = ~new_P2_R2267_U31;
  assign new_P2_R2267_U103 = ~new_P2_R2267_U32;
  assign new_P2_R2267_U104 = ~new_P2_R2267_U33;
  assign new_P2_R2267_U105 = ~new_P2_R2267_U34;
  assign new_P2_R2267_U106 = ~new_P2_R2267_U35;
  assign new_P2_R2267_U107 = ~new_P2_R2267_U36;
  assign new_P2_R2267_U108 = ~new_P2_R2267_U37;
  assign new_P2_R2267_U109 = ~new_P2_R2267_U38;
  assign new_P2_R2267_U110 = ~new_P2_R2267_U39;
  assign new_P2_R2267_U111 = ~new_P2_R2267_U40;
  assign new_P2_R2267_U112 = ~new_P2_R2267_U62;
  assign new_P2_R2267_U113 = ~new_P2_U2767 | ~new_P2_R2267_U40;
  assign new_P2_R2267_U114 = ~new_P2_R2267_U110 | ~new_P2_R2267_U66;
  assign new_P2_R2267_U115 = ~new_P2_U2768 | ~new_P2_R2267_U114;
  assign new_P2_R2267_U116 = ~new_P2_R2267_U109 | ~new_P2_R2267_U68;
  assign new_P2_R2267_U117 = ~new_P2_U2770 | ~new_P2_R2267_U116;
  assign new_P2_R2267_U118 = ~new_P2_R2267_U108 | ~new_P2_R2267_U70;
  assign new_P2_R2267_U119 = ~new_P2_U2772 | ~new_P2_R2267_U118;
  assign new_P2_R2267_U120 = ~new_P2_R2267_U107 | ~new_P2_R2267_U72;
  assign new_P2_R2267_U121 = ~new_P2_U2774 | ~new_P2_R2267_U120;
  assign new_P2_R2267_U122 = ~new_P2_R2267_U106 | ~new_P2_R2267_U74;
  assign new_P2_R2267_U123 = ~new_P2_U2776 | ~new_P2_R2267_U122;
  assign new_P2_R2267_U124 = ~new_P2_R2267_U105 | ~new_P2_R2267_U78;
  assign new_P2_R2267_U125 = ~new_P2_U2778 | ~new_P2_R2267_U124;
  assign new_P2_R2267_U126 = ~new_P2_R2267_U104 | ~new_P2_R2267_U80;
  assign new_P2_R2267_U127 = ~new_P2_U2780 | ~new_P2_R2267_U126;
  assign new_P2_R2267_U128 = ~new_P2_R2267_U103 | ~new_P2_R2267_U82;
  assign new_P2_R2267_U129 = ~new_P2_U2782 | ~new_P2_R2267_U128;
  assign new_P2_R2267_U130 = ~new_P2_R2267_U102 | ~new_P2_R2267_U84;
  assign new_P2_R2267_U131 = ~new_P2_U2784 | ~new_P2_R2267_U130;
  assign new_P2_R2267_U132 = ~new_P2_R2267_U93 | ~new_P2_R2267_U86;
  assign new_P2_R2267_U133 = ~new_P2_U2786 | ~new_P2_R2267_U132;
  assign new_P2_R2267_U134 = ~new_P2_U2617 | ~new_P2_R2267_U22;
  assign new_P2_R2267_U135 = ~new_P2_U2789 | ~new_P2_R2267_U26;
  assign new_P2_R2267_U136 = ~new_P2_R2267_U92 | ~new_P2_R2267_U55;
  assign new_P2_R2267_U137 = ~new_P2_U3640 | ~new_P2_R2267_U25;
  assign new_P2_R2267_U138 = ~new_P2_R2267_U91 | ~new_P2_R2267_U57;
  assign new_P2_R2267_U139 = ~new_P2_U3642 | ~new_P2_R2267_U24;
  assign new_P2_R2267_U140 = ~new_P2_R2267_U90 | ~new_P2_R2267_U59;
  assign new_P2_R2267_U141 = ~new_P2_U2766 | ~new_P2_R2267_U62;
  assign new_P2_R2267_U142 = ~new_P2_R2267_U112 | ~new_P2_R2267_U61;
  assign new_P2_R2267_U143 = ~new_P2_U3644 | ~new_P2_R2267_U23;
  assign new_P2_R2267_U144 = ~new_P2_R2267_U89 | ~new_P2_R2267_U64;
  assign new_P2_R2267_U145 = ~new_P2_U2769 | ~new_P2_R2267_U39;
  assign new_P2_R2267_U146 = ~new_P2_R2267_U110 | ~new_P2_R2267_U66;
  assign new_P2_R2267_U147 = ~new_P2_U2771 | ~new_P2_R2267_U38;
  assign new_P2_R2267_U148 = ~new_P2_R2267_U109 | ~new_P2_R2267_U68;
  assign new_P2_R2267_U149 = ~new_P2_U2773 | ~new_P2_R2267_U37;
  assign new_P2_R2267_U150 = ~new_P2_R2267_U108 | ~new_P2_R2267_U70;
  assign new_P2_R2267_U151 = ~new_P2_U2775 | ~new_P2_R2267_U36;
  assign new_P2_R2267_U152 = ~new_P2_R2267_U107 | ~new_P2_R2267_U72;
  assign new_P2_R2267_U153 = ~new_P2_U2777 | ~new_P2_R2267_U35;
  assign new_P2_R2267_U154 = ~new_P2_R2267_U106 | ~new_P2_R2267_U74;
  assign new_P2_R2267_U155 = ~new_P2_U3645 | ~new_P2_R2267_U77;
  assign new_P2_R2267_U156 = ~new_P2_R2267_U88 | ~new_P2_R2267_U76;
  assign new_P2_R2267_U157 = ~new_P2_U2779 | ~new_P2_R2267_U34;
  assign new_P2_R2267_U158 = ~new_P2_R2267_U105 | ~new_P2_R2267_U78;
  assign new_P2_R2267_U159 = ~new_P2_U2781 | ~new_P2_R2267_U33;
  assign new_P2_R2267_U160 = ~new_P2_R2267_U104 | ~new_P2_R2267_U80;
  assign new_P2_R2267_U161 = ~new_P2_U2783 | ~new_P2_R2267_U32;
  assign new_P2_R2267_U162 = ~new_P2_R2267_U103 | ~new_P2_R2267_U82;
  assign new_P2_R2267_U163 = ~new_P2_U2785 | ~new_P2_R2267_U31;
  assign new_P2_R2267_U164 = ~new_P2_R2267_U102 | ~new_P2_R2267_U84;
  assign new_P2_R2267_U165 = ~new_P2_U2787 | ~new_P2_R2267_U30;
  assign new_P2_R2267_U166 = ~new_P2_R2267_U93 | ~new_P2_R2267_U86;
  assign new_P2_ADD_371_1212_U4 = P2_INSTADDRPOINTER_REG_13_ & new_P2_ADD_371_1212_U10;
  assign new_P2_ADD_371_1212_U5 = P2_INSTADDRPOINTER_REG_10_ & P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_ADD_371_1212_U6 = new_P2_ADD_371_1212_U89 & new_P2_ADD_371_1212_U11;
  assign new_P2_ADD_371_1212_U7 = new_P2_ADD_371_1212_U10 & new_P2_ADD_371_1212_U87;
  assign new_P2_ADD_371_1212_U8 = new_P2_ADD_371_1212_U9 & new_P2_ADD_371_1212_U91;
  assign new_P2_ADD_371_1212_U9 = new_P2_ADD_371_1212_U6 & new_P2_ADD_371_1212_U90;
  assign new_P2_ADD_371_1212_U10 = P2_INSTADDRPOINTER_REG_9_ & P2_INSTADDRPOINTER_REG_10_ & P2_INSTADDRPOINTER_REG_12_ & P2_INSTADDRPOINTER_REG_11_;
  assign new_P2_ADD_371_1212_U11 = new_P2_ADD_371_1212_U7 & new_P2_ADD_371_1212_U88;
  assign new_P2_ADD_371_1212_U12 = new_P2_ADD_371_1212_U8 & new_P2_ADD_371_1212_U92;
  assign new_P2_ADD_371_1212_U13 = new_P2_ADD_371_1212_U196 & new_P2_ADD_371_1212_U168;
  assign new_P2_ADD_371_1212_U14 = new_P2_ADD_371_1212_U188 & new_P2_ADD_371_1212_U132;
  assign new_P2_ADD_371_1212_U15 = new_P2_ADD_371_1212_U185 & new_P2_ADD_371_1212_U170;
  assign new_P2_ADD_371_1212_U16 = new_P2_ADD_371_1212_U191 & new_P2_ADD_371_1212_U120;
  assign new_P2_ADD_371_1212_U17 = new_P2_ADD_371_1212_U200 & new_P2_ADD_371_1212_U114;
  assign new_P2_ADD_371_1212_U18 = new_P2_ADD_371_1212_U194 & new_P2_ADD_371_1212_U174;
  assign new_P2_ADD_371_1212_U19 = new_P2_ADD_371_1212_U183 & new_P2_ADD_371_1212_U131;
  assign new_P2_ADD_371_1212_U20 = new_P2_ADD_371_1212_U187 & new_P2_ADD_371_1212_U176;
  assign new_P2_ADD_371_1212_U21 = new_P2_ADD_371_1212_U192 & new_P2_ADD_371_1212_U113;
  assign new_P2_ADD_371_1212_U22 = new_P2_ADD_371_1212_U190 & new_P2_ADD_371_1212_U123;
  assign new_P2_ADD_371_1212_U23 = new_P2_ADD_371_1212_U198 & new_P2_ADD_371_1212_U180;
  assign new_P2_ADD_371_1212_U24 = new_P2_ADD_371_1212_U182 & new_P2_ADD_371_1212_U112;
  assign new_P2_ADD_371_1212_U25 = ~new_P2_ADD_371_1212_U204 | ~new_P2_ADD_371_1212_U269 | ~new_P2_ADD_371_1212_U268;
  assign new_P2_ADD_371_1212_U26 = ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_ADD_371_1212_U27 = ~new_P2_R2256_U21;
  assign new_P2_ADD_371_1212_U28 = ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_ADD_371_1212_U29 = ~new_P2_R2256_U21 | ~P2_INSTADDRPOINTER_REG_0_;
  assign new_P2_ADD_371_1212_U30 = ~new_P2_R2256_U4;
  assign new_P2_ADD_371_1212_U31 = ~new_P2_R2256_U22;
  assign new_P2_ADD_371_1212_U32 = ~P2_INSTADDRPOINTER_REG_2_;
  assign new_P2_ADD_371_1212_U33 = ~new_P2_R2256_U26;
  assign new_P2_ADD_371_1212_U34 = ~P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_ADD_371_1212_U35 = ~new_P2_R2256_U20;
  assign new_P2_ADD_371_1212_U36 = ~P2_INSTADDRPOINTER_REG_4_;
  assign new_P2_ADD_371_1212_U37 = ~new_P2_R2256_U19;
  assign new_P2_ADD_371_1212_U38 = ~P2_INSTADDRPOINTER_REG_5_;
  assign new_P2_ADD_371_1212_U39 = ~P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_ADD_371_1212_U40 = ~new_P2_R2256_U18;
  assign new_P2_ADD_371_1212_U41 = ~new_P2_R2256_U5;
  assign new_P2_ADD_371_1212_U42 = ~P2_INSTADDRPOINTER_REG_8_;
  assign new_P2_ADD_371_1212_U43 = ~new_P2_R2256_U17;
  assign new_P2_ADD_371_1212_U44 = ~P2_INSTADDRPOINTER_REG_7_;
  assign new_P2_ADD_371_1212_U45 = ~P2_INSTADDRPOINTER_REG_9_;
  assign new_P2_ADD_371_1212_U46 = ~P2_INSTADDRPOINTER_REG_10_;
  assign new_P2_ADD_371_1212_U47 = ~P2_INSTADDRPOINTER_REG_11_;
  assign new_P2_ADD_371_1212_U48 = ~P2_INSTADDRPOINTER_REG_12_;
  assign new_P2_ADD_371_1212_U49 = ~P2_INSTADDRPOINTER_REG_13_;
  assign new_P2_ADD_371_1212_U50 = ~P2_INSTADDRPOINTER_REG_14_;
  assign new_P2_ADD_371_1212_U51 = ~P2_INSTADDRPOINTER_REG_15_;
  assign new_P2_ADD_371_1212_U52 = ~P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_ADD_371_1212_U53 = ~P2_INSTADDRPOINTER_REG_18_;
  assign new_P2_ADD_371_1212_U54 = ~P2_INSTADDRPOINTER_REG_17_;
  assign new_P2_ADD_371_1212_U55 = ~P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_ADD_371_1212_U56 = ~P2_INSTADDRPOINTER_REG_20_;
  assign new_P2_ADD_371_1212_U57 = ~P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_ADD_371_1212_U58 = ~P2_INSTADDRPOINTER_REG_22_;
  assign new_P2_ADD_371_1212_U59 = ~P2_INSTADDRPOINTER_REG_23_;
  assign new_P2_ADD_371_1212_U60 = ~P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_ADD_371_1212_U61 = ~P2_INSTADDRPOINTER_REG_26_;
  assign new_P2_ADD_371_1212_U62 = ~P2_INSTADDRPOINTER_REG_25_;
  assign new_P2_ADD_371_1212_U63 = ~P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_ADD_371_1212_U64 = ~P2_INSTADDRPOINTER_REG_28_;
  assign new_P2_ADD_371_1212_U65 = ~P2_INSTADDRPOINTER_REG_29_;
  assign new_P2_ADD_371_1212_U66 = ~P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_ADD_371_1212_U67 = ~new_P2_R2256_U4 | ~new_P2_ADD_371_1212_U137;
  assign new_P2_ADD_371_1212_U68 = ~new_P2_ADD_371_1212_U206 | ~new_P2_ADD_371_1212_U205;
  assign new_P2_ADD_371_1212_U69 = ~new_P2_ADD_371_1212_U215 | ~new_P2_ADD_371_1212_U214;
  assign new_P2_ADD_371_1212_U70 = ~new_P2_ADD_371_1212_U217 | ~new_P2_ADD_371_1212_U216;
  assign new_P2_ADD_371_1212_U71 = ~new_P2_ADD_371_1212_U219 | ~new_P2_ADD_371_1212_U218;
  assign new_P2_ADD_371_1212_U72 = ~new_P2_ADD_371_1212_U230 | ~new_P2_ADD_371_1212_U229;
  assign new_P2_ADD_371_1212_U73 = ~new_P2_ADD_371_1212_U232 | ~new_P2_ADD_371_1212_U231;
  assign new_P2_ADD_371_1212_U74 = ~new_P2_ADD_371_1212_U241 | ~new_P2_ADD_371_1212_U240;
  assign new_P2_ADD_371_1212_U75 = ~new_P2_ADD_371_1212_U271 | ~new_P2_ADD_371_1212_U270;
  assign new_P2_ADD_371_1212_U76 = ~new_P2_ADD_371_1212_U273 | ~new_P2_ADD_371_1212_U272;
  assign new_P2_ADD_371_1212_U77 = ~new_P2_ADD_371_1212_U282 | ~new_P2_ADD_371_1212_U281;
  assign new_P2_ADD_371_1212_U78 = ~new_P2_ADD_371_1212_U213 | ~new_P2_ADD_371_1212_U212;
  assign new_P2_ADD_371_1212_U79 = ~new_P2_ADD_371_1212_U226 | ~new_P2_ADD_371_1212_U225;
  assign new_P2_ADD_371_1212_U80 = ~new_P2_ADD_371_1212_U239 | ~new_P2_ADD_371_1212_U238;
  assign new_P2_ADD_371_1212_U81 = ~new_P2_ADD_371_1212_U248 | ~new_P2_ADD_371_1212_U247;
  assign new_P2_ADD_371_1212_U82 = ~new_P2_ADD_371_1212_U255 | ~new_P2_ADD_371_1212_U254;
  assign new_P2_ADD_371_1212_U83 = ~new_P2_ADD_371_1212_U257 | ~new_P2_ADD_371_1212_U256;
  assign new_P2_ADD_371_1212_U84 = ~new_P2_ADD_371_1212_U264 | ~new_P2_ADD_371_1212_U263;
  assign new_P2_ADD_371_1212_U85 = ~new_P2_ADD_371_1212_U280 | ~new_P2_ADD_371_1212_U279;
  assign new_P2_ADD_371_1212_U86 = new_P2_ADD_371_1212_U203 & new_P2_ADD_371_1212_U166;
  assign new_P2_ADD_371_1212_U87 = P2_INSTADDRPOINTER_REG_13_ & P2_INSTADDRPOINTER_REG_15_ & P2_INSTADDRPOINTER_REG_14_;
  assign new_P2_ADD_371_1212_U88 = P2_INSTADDRPOINTER_REG_16_ & P2_INSTADDRPOINTER_REG_17_ & P2_INSTADDRPOINTER_REG_18_;
  assign new_P2_ADD_371_1212_U89 = P2_INSTADDRPOINTER_REG_19_ & P2_INSTADDRPOINTER_REG_20_;
  assign new_P2_ADD_371_1212_U90 = P2_INSTADDRPOINTER_REG_21_ & P2_INSTADDRPOINTER_REG_23_ & P2_INSTADDRPOINTER_REG_22_;
  assign new_P2_ADD_371_1212_U91 = P2_INSTADDRPOINTER_REG_24_ & P2_INSTADDRPOINTER_REG_25_ & P2_INSTADDRPOINTER_REG_26_;
  assign new_P2_ADD_371_1212_U92 = P2_INSTADDRPOINTER_REG_27_ & P2_INSTADDRPOINTER_REG_29_ & P2_INSTADDRPOINTER_REG_28_;
  assign new_P2_ADD_371_1212_U93 = new_P2_ADD_371_1212_U8 & new_P2_ADD_371_1212_U94;
  assign new_P2_ADD_371_1212_U94 = P2_INSTADDRPOINTER_REG_28_ & P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_ADD_371_1212_U95 = new_P2_ADD_371_1212_U7 & P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_ADD_371_1212_U96 = new_P2_ADD_371_1212_U11 & P2_INSTADDRPOINTER_REG_19_;
  assign new_P2_ADD_371_1212_U97 = new_P2_ADD_371_1212_U6 & new_P2_ADD_371_1212_U98;
  assign new_P2_ADD_371_1212_U98 = P2_INSTADDRPOINTER_REG_22_ & P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_ADD_371_1212_U99 = new_P2_ADD_371_1212_U6 & P2_INSTADDRPOINTER_REG_21_;
  assign new_P2_ADD_371_1212_U100 = new_P2_ADD_371_1212_U7 & new_P2_ADD_371_1212_U101;
  assign new_P2_ADD_371_1212_U101 = P2_INSTADDRPOINTER_REG_17_ & P2_INSTADDRPOINTER_REG_16_;
  assign new_P2_ADD_371_1212_U102 = P2_INSTADDRPOINTER_REG_11_ & new_P2_ADD_371_1212_U5;
  assign new_P2_ADD_371_1212_U103 = new_P2_ADD_371_1212_U9 & new_P2_ADD_371_1212_U104;
  assign new_P2_ADD_371_1212_U104 = P2_INSTADDRPOINTER_REG_25_ & P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_ADD_371_1212_U105 = P2_INSTADDRPOINTER_REG_14_ & new_P2_ADD_371_1212_U4;
  assign new_P2_ADD_371_1212_U106 = new_P2_ADD_371_1212_U12 & P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_ADD_371_1212_U107 = new_P2_ADD_371_1212_U12 & P2_INSTADDRPOINTER_REG_30_;
  assign new_P2_ADD_371_1212_U108 = new_P2_ADD_371_1212_U8 & P2_INSTADDRPOINTER_REG_27_;
  assign new_P2_ADD_371_1212_U109 = new_P2_ADD_371_1212_U9 & P2_INSTADDRPOINTER_REG_24_;
  assign new_P2_ADD_371_1212_U110 = new_P2_ADD_371_1212_U208 & new_P2_ADD_371_1212_U207;
  assign new_P2_ADD_371_1212_U111 = ~new_P2_ADD_371_1212_U155 | ~new_P2_ADD_371_1212_U154;
  assign new_P2_ADD_371_1212_U112 = ~new_P2_ADD_371_1212_U12 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U113 = ~new_P2_ADD_371_1212_U9 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U114 = ~new_P2_ADD_371_1212_U95 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U115 = new_P2_ADD_371_1212_U221 & new_P2_ADD_371_1212_U220;
  assign new_P2_ADD_371_1212_U116 = ~new_P2_ADD_371_1212_U67 | ~new_P2_ADD_371_1212_U139;
  assign new_P2_ADD_371_1212_U117 = ~new_P2_ADD_371_1212_U86 | ~new_P2_ADD_371_1212_U202;
  assign new_P2_ADD_371_1212_U118 = new_P2_ADD_371_1212_U228 & new_P2_ADD_371_1212_U227;
  assign new_P2_ADD_371_1212_U119 = ~new_P2_ADD_371_1212_U117 | ~new_P2_ADD_371_1212_U100;
  assign new_P2_ADD_371_1212_U120 = ~new_P2_ADD_371_1212_U105 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U121 = new_P2_ADD_371_1212_U234 & new_P2_ADD_371_1212_U233;
  assign new_P2_ADD_371_1212_U122 = ~new_P2_ADD_371_1212_U147 | ~new_P2_ADD_371_1212_U146;
  assign new_P2_ADD_371_1212_U123 = ~new_P2_ADD_371_1212_U8 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U124 = new_P2_ADD_371_1212_U243 & new_P2_ADD_371_1212_U242;
  assign new_P2_ADD_371_1212_U125 = ~new_P2_ADD_371_1212_U151 | ~new_P2_ADD_371_1212_U150;
  assign new_P2_ADD_371_1212_U126 = new_P2_ADD_371_1212_U250 & new_P2_ADD_371_1212_U249;
  assign new_P2_ADD_371_1212_U127 = ~new_P2_ADD_371_1212_U163 | ~new_P2_ADD_371_1212_U162;
  assign new_P2_ADD_371_1212_U128 = ~P2_INSTADDRPOINTER_REG_31_;
  assign new_P2_ADD_371_1212_U129 = new_P2_ADD_371_1212_U259 & new_P2_ADD_371_1212_U258;
  assign new_P2_ADD_371_1212_U130 = ~new_P2_ADD_371_1212_U143 | ~new_P2_ADD_371_1212_U142;
  assign new_P2_ADD_371_1212_U131 = ~new_P2_ADD_371_1212_U6 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U132 = ~new_P2_ADD_371_1212_U102 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U133 = new_P2_ADD_371_1212_U275 & new_P2_ADD_371_1212_U274;
  assign new_P2_ADD_371_1212_U134 = ~new_P2_ADD_371_1212_U159 | ~new_P2_ADD_371_1212_U158;
  assign new_P2_ADD_371_1212_U135 = ~new_P2_ADD_371_1212_U109 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U136 = ~new_P2_ADD_371_1212_U67;
  assign new_P2_ADD_371_1212_U137 = ~new_P2_ADD_371_1212_U29;
  assign new_P2_ADD_371_1212_U138 = ~new_P2_ADD_371_1212_U30 | ~new_P2_ADD_371_1212_U29;
  assign new_P2_ADD_371_1212_U139 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_ADD_371_1212_U138;
  assign new_P2_ADD_371_1212_U140 = ~new_P2_ADD_371_1212_U116;
  assign new_P2_ADD_371_1212_U141 = new_P2_R2256_U22 | P2_INSTADDRPOINTER_REG_2_;
  assign new_P2_ADD_371_1212_U142 = ~new_P2_ADD_371_1212_U141 | ~new_P2_ADD_371_1212_U116;
  assign new_P2_ADD_371_1212_U143 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_R2256_U22;
  assign new_P2_ADD_371_1212_U144 = ~new_P2_ADD_371_1212_U130;
  assign new_P2_ADD_371_1212_U145 = new_P2_R2256_U26 | P2_INSTADDRPOINTER_REG_3_;
  assign new_P2_ADD_371_1212_U146 = ~new_P2_ADD_371_1212_U145 | ~new_P2_ADD_371_1212_U130;
  assign new_P2_ADD_371_1212_U147 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_R2256_U26;
  assign new_P2_ADD_371_1212_U148 = ~new_P2_ADD_371_1212_U122;
  assign new_P2_ADD_371_1212_U149 = new_P2_R2256_U20 | P2_INSTADDRPOINTER_REG_4_;
  assign new_P2_ADD_371_1212_U150 = ~new_P2_ADD_371_1212_U149 | ~new_P2_ADD_371_1212_U122;
  assign new_P2_ADD_371_1212_U151 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_R2256_U20;
  assign new_P2_ADD_371_1212_U152 = ~new_P2_ADD_371_1212_U125;
  assign new_P2_ADD_371_1212_U153 = new_P2_R2256_U19 | P2_INSTADDRPOINTER_REG_5_;
  assign new_P2_ADD_371_1212_U154 = ~new_P2_ADD_371_1212_U153 | ~new_P2_ADD_371_1212_U125;
  assign new_P2_ADD_371_1212_U155 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_R2256_U19;
  assign new_P2_ADD_371_1212_U156 = ~new_P2_ADD_371_1212_U111;
  assign new_P2_ADD_371_1212_U157 = new_P2_R2256_U18 | P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_ADD_371_1212_U158 = ~new_P2_ADD_371_1212_U157 | ~new_P2_ADD_371_1212_U111;
  assign new_P2_ADD_371_1212_U159 = ~new_P2_R2256_U18 | ~P2_INSTADDRPOINTER_REG_6_;
  assign new_P2_ADD_371_1212_U160 = ~new_P2_ADD_371_1212_U134;
  assign new_P2_ADD_371_1212_U161 = new_P2_R2256_U17 | P2_INSTADDRPOINTER_REG_7_;
  assign new_P2_ADD_371_1212_U162 = ~new_P2_ADD_371_1212_U161 | ~new_P2_ADD_371_1212_U134;
  assign new_P2_ADD_371_1212_U163 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_R2256_U17;
  assign new_P2_ADD_371_1212_U164 = ~new_P2_ADD_371_1212_U127;
  assign new_P2_ADD_371_1212_U165 = new_P2_R2256_U5 | P2_INSTADDRPOINTER_REG_8_;
  assign new_P2_ADD_371_1212_U166 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_R2256_U5;
  assign new_P2_ADD_371_1212_U167 = ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U168 = ~new_P2_ADD_371_1212_U5 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U169 = ~new_P2_ADD_371_1212_U132;
  assign new_P2_ADD_371_1212_U170 = ~new_P2_ADD_371_1212_U4 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U171 = ~new_P2_ADD_371_1212_U120;
  assign new_P2_ADD_371_1212_U172 = ~new_P2_ADD_371_1212_U114;
  assign new_P2_ADD_371_1212_U173 = ~new_P2_ADD_371_1212_U119;
  assign new_P2_ADD_371_1212_U174 = ~new_P2_ADD_371_1212_U96 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U175 = ~new_P2_ADD_371_1212_U131;
  assign new_P2_ADD_371_1212_U176 = ~new_P2_ADD_371_1212_U117 | ~new_P2_ADD_371_1212_U97;
  assign new_P2_ADD_371_1212_U177 = ~new_P2_ADD_371_1212_U113;
  assign new_P2_ADD_371_1212_U178 = ~new_P2_ADD_371_1212_U135;
  assign new_P2_ADD_371_1212_U179 = ~new_P2_ADD_371_1212_U123;
  assign new_P2_ADD_371_1212_U180 = ~new_P2_ADD_371_1212_U117 | ~new_P2_ADD_371_1212_U93;
  assign new_P2_ADD_371_1212_U181 = ~new_P2_ADD_371_1212_U112;
  assign new_P2_ADD_371_1212_U182 = ~new_P2_ADD_371_1212_U65 | ~new_P2_ADD_371_1212_U180;
  assign new_P2_ADD_371_1212_U183 = ~new_P2_ADD_371_1212_U56 | ~new_P2_ADD_371_1212_U174;
  assign new_P2_ADD_371_1212_U184 = ~new_P2_ADD_371_1212_U10 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U185 = ~new_P2_ADD_371_1212_U49 | ~new_P2_ADD_371_1212_U184;
  assign new_P2_ADD_371_1212_U186 = ~new_P2_ADD_371_1212_U99 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U187 = ~new_P2_ADD_371_1212_U58 | ~new_P2_ADD_371_1212_U186;
  assign new_P2_ADD_371_1212_U188 = ~new_P2_ADD_371_1212_U47 | ~new_P2_ADD_371_1212_U168;
  assign new_P2_ADD_371_1212_U189 = ~new_P2_ADD_371_1212_U117 | ~new_P2_ADD_371_1212_U103;
  assign new_P2_ADD_371_1212_U190 = ~new_P2_ADD_371_1212_U61 | ~new_P2_ADD_371_1212_U189;
  assign new_P2_ADD_371_1212_U191 = ~new_P2_ADD_371_1212_U50 | ~new_P2_ADD_371_1212_U170;
  assign new_P2_ADD_371_1212_U192 = ~new_P2_ADD_371_1212_U59 | ~new_P2_ADD_371_1212_U176;
  assign new_P2_ADD_371_1212_U193 = ~new_P2_ADD_371_1212_U11 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U194 = ~new_P2_ADD_371_1212_U55 | ~new_P2_ADD_371_1212_U193;
  assign new_P2_ADD_371_1212_U195 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U196 = ~new_P2_ADD_371_1212_U46 | ~new_P2_ADD_371_1212_U195;
  assign new_P2_ADD_371_1212_U197 = ~new_P2_ADD_371_1212_U108 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U198 = ~new_P2_ADD_371_1212_U64 | ~new_P2_ADD_371_1212_U197;
  assign new_P2_ADD_371_1212_U199 = ~new_P2_ADD_371_1212_U7 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U200 = ~new_P2_ADD_371_1212_U52 | ~new_P2_ADD_371_1212_U199;
  assign new_P2_ADD_371_1212_U201 = ~new_P2_ADD_371_1212_U107 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U202 = ~new_P2_ADD_371_1212_U161 | ~new_P2_ADD_371_1212_U165 | ~new_P2_ADD_371_1212_U134;
  assign new_P2_ADD_371_1212_U203 = ~new_P2_R2256_U17 | ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_ADD_371_1212_U165;
  assign new_P2_ADD_371_1212_U204 = ~new_P2_ADD_371_1212_U136 | ~P2_INSTADDRPOINTER_REG_1_;
  assign new_P2_ADD_371_1212_U205 = ~P2_INSTADDRPOINTER_REG_0_ | ~new_P2_ADD_371_1212_U27;
  assign new_P2_ADD_371_1212_U206 = ~new_P2_R2256_U21 | ~new_P2_ADD_371_1212_U26;
  assign new_P2_ADD_371_1212_U207 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_ADD_371_1212_U40;
  assign new_P2_ADD_371_1212_U208 = ~new_P2_R2256_U18 | ~new_P2_ADD_371_1212_U39;
  assign new_P2_ADD_371_1212_U209 = ~P2_INSTADDRPOINTER_REG_6_ | ~new_P2_ADD_371_1212_U40;
  assign new_P2_ADD_371_1212_U210 = ~new_P2_R2256_U18 | ~new_P2_ADD_371_1212_U39;
  assign new_P2_ADD_371_1212_U211 = ~new_P2_ADD_371_1212_U210 | ~new_P2_ADD_371_1212_U209;
  assign new_P2_ADD_371_1212_U212 = ~new_P2_ADD_371_1212_U110 | ~new_P2_ADD_371_1212_U111;
  assign new_P2_ADD_371_1212_U213 = ~new_P2_ADD_371_1212_U156 | ~new_P2_ADD_371_1212_U211;
  assign new_P2_ADD_371_1212_U214 = ~P2_INSTADDRPOINTER_REG_30_ | ~new_P2_ADD_371_1212_U112;
  assign new_P2_ADD_371_1212_U215 = ~new_P2_ADD_371_1212_U181 | ~new_P2_ADD_371_1212_U66;
  assign new_P2_ADD_371_1212_U216 = ~P2_INSTADDRPOINTER_REG_24_ | ~new_P2_ADD_371_1212_U113;
  assign new_P2_ADD_371_1212_U217 = ~new_P2_ADD_371_1212_U177 | ~new_P2_ADD_371_1212_U60;
  assign new_P2_ADD_371_1212_U218 = ~P2_INSTADDRPOINTER_REG_17_ | ~new_P2_ADD_371_1212_U114;
  assign new_P2_ADD_371_1212_U219 = ~new_P2_ADD_371_1212_U172 | ~new_P2_ADD_371_1212_U54;
  assign new_P2_ADD_371_1212_U220 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_ADD_371_1212_U31;
  assign new_P2_ADD_371_1212_U221 = ~new_P2_R2256_U22 | ~new_P2_ADD_371_1212_U32;
  assign new_P2_ADD_371_1212_U222 = ~P2_INSTADDRPOINTER_REG_2_ | ~new_P2_ADD_371_1212_U31;
  assign new_P2_ADD_371_1212_U223 = ~new_P2_R2256_U22 | ~new_P2_ADD_371_1212_U32;
  assign new_P2_ADD_371_1212_U224 = ~new_P2_ADD_371_1212_U223 | ~new_P2_ADD_371_1212_U222;
  assign new_P2_ADD_371_1212_U225 = ~new_P2_ADD_371_1212_U115 | ~new_P2_ADD_371_1212_U116;
  assign new_P2_ADD_371_1212_U226 = ~new_P2_ADD_371_1212_U140 | ~new_P2_ADD_371_1212_U224;
  assign new_P2_ADD_371_1212_U227 = ~P2_INSTADDRPOINTER_REG_9_ | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U228 = ~new_P2_ADD_371_1212_U167 | ~new_P2_ADD_371_1212_U45;
  assign new_P2_ADD_371_1212_U229 = ~P2_INSTADDRPOINTER_REG_18_ | ~new_P2_ADD_371_1212_U119;
  assign new_P2_ADD_371_1212_U230 = ~new_P2_ADD_371_1212_U173 | ~new_P2_ADD_371_1212_U53;
  assign new_P2_ADD_371_1212_U231 = ~P2_INSTADDRPOINTER_REG_15_ | ~new_P2_ADD_371_1212_U120;
  assign new_P2_ADD_371_1212_U232 = ~new_P2_ADD_371_1212_U171 | ~new_P2_ADD_371_1212_U51;
  assign new_P2_ADD_371_1212_U233 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_ADD_371_1212_U35;
  assign new_P2_ADD_371_1212_U234 = ~new_P2_R2256_U20 | ~new_P2_ADD_371_1212_U36;
  assign new_P2_ADD_371_1212_U235 = ~P2_INSTADDRPOINTER_REG_4_ | ~new_P2_ADD_371_1212_U35;
  assign new_P2_ADD_371_1212_U236 = ~new_P2_R2256_U20 | ~new_P2_ADD_371_1212_U36;
  assign new_P2_ADD_371_1212_U237 = ~new_P2_ADD_371_1212_U236 | ~new_P2_ADD_371_1212_U235;
  assign new_P2_ADD_371_1212_U238 = ~new_P2_ADD_371_1212_U121 | ~new_P2_ADD_371_1212_U122;
  assign new_P2_ADD_371_1212_U239 = ~new_P2_ADD_371_1212_U148 | ~new_P2_ADD_371_1212_U237;
  assign new_P2_ADD_371_1212_U240 = ~P2_INSTADDRPOINTER_REG_27_ | ~new_P2_ADD_371_1212_U123;
  assign new_P2_ADD_371_1212_U241 = ~new_P2_ADD_371_1212_U179 | ~new_P2_ADD_371_1212_U63;
  assign new_P2_ADD_371_1212_U242 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_ADD_371_1212_U37;
  assign new_P2_ADD_371_1212_U243 = ~new_P2_R2256_U19 | ~new_P2_ADD_371_1212_U38;
  assign new_P2_ADD_371_1212_U244 = ~P2_INSTADDRPOINTER_REG_5_ | ~new_P2_ADD_371_1212_U37;
  assign new_P2_ADD_371_1212_U245 = ~new_P2_R2256_U19 | ~new_P2_ADD_371_1212_U38;
  assign new_P2_ADD_371_1212_U246 = ~new_P2_ADD_371_1212_U245 | ~new_P2_ADD_371_1212_U244;
  assign new_P2_ADD_371_1212_U247 = ~new_P2_ADD_371_1212_U124 | ~new_P2_ADD_371_1212_U125;
  assign new_P2_ADD_371_1212_U248 = ~new_P2_ADD_371_1212_U152 | ~new_P2_ADD_371_1212_U246;
  assign new_P2_ADD_371_1212_U249 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_ADD_371_1212_U41;
  assign new_P2_ADD_371_1212_U250 = ~new_P2_R2256_U5 | ~new_P2_ADD_371_1212_U42;
  assign new_P2_ADD_371_1212_U251 = ~P2_INSTADDRPOINTER_REG_8_ | ~new_P2_ADD_371_1212_U41;
  assign new_P2_ADD_371_1212_U252 = ~new_P2_R2256_U5 | ~new_P2_ADD_371_1212_U42;
  assign new_P2_ADD_371_1212_U253 = ~new_P2_ADD_371_1212_U252 | ~new_P2_ADD_371_1212_U251;
  assign new_P2_ADD_371_1212_U254 = ~new_P2_ADD_371_1212_U126 | ~new_P2_ADD_371_1212_U127;
  assign new_P2_ADD_371_1212_U255 = ~new_P2_ADD_371_1212_U164 | ~new_P2_ADD_371_1212_U253;
  assign new_P2_ADD_371_1212_U256 = ~P2_INSTADDRPOINTER_REG_31_ | ~new_P2_ADD_371_1212_U201;
  assign new_P2_ADD_371_1212_U257 = ~new_P2_ADD_371_1212_U128 | ~new_P2_ADD_371_1212_U106 | ~new_P2_ADD_371_1212_U117;
  assign new_P2_ADD_371_1212_U258 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_ADD_371_1212_U33;
  assign new_P2_ADD_371_1212_U259 = ~new_P2_R2256_U26 | ~new_P2_ADD_371_1212_U34;
  assign new_P2_ADD_371_1212_U260 = ~P2_INSTADDRPOINTER_REG_3_ | ~new_P2_ADD_371_1212_U33;
  assign new_P2_ADD_371_1212_U261 = ~new_P2_R2256_U26 | ~new_P2_ADD_371_1212_U34;
  assign new_P2_ADD_371_1212_U262 = ~new_P2_ADD_371_1212_U261 | ~new_P2_ADD_371_1212_U260;
  assign new_P2_ADD_371_1212_U263 = ~new_P2_ADD_371_1212_U129 | ~new_P2_ADD_371_1212_U130;
  assign new_P2_ADD_371_1212_U264 = ~new_P2_ADD_371_1212_U144 | ~new_P2_ADD_371_1212_U262;
  assign new_P2_ADD_371_1212_U265 = ~P2_INSTADDRPOINTER_REG_1_ | ~new_P2_ADD_371_1212_U29;
  assign new_P2_ADD_371_1212_U266 = ~new_P2_ADD_371_1212_U137 | ~new_P2_ADD_371_1212_U28;
  assign new_P2_ADD_371_1212_U267 = ~new_P2_ADD_371_1212_U266 | ~new_P2_ADD_371_1212_U265;
  assign new_P2_ADD_371_1212_U268 = ~new_P2_R2256_U4 | ~new_P2_ADD_371_1212_U29 | ~new_P2_ADD_371_1212_U28;
  assign new_P2_ADD_371_1212_U269 = ~new_P2_ADD_371_1212_U267 | ~new_P2_ADD_371_1212_U30;
  assign new_P2_ADD_371_1212_U270 = ~P2_INSTADDRPOINTER_REG_21_ | ~new_P2_ADD_371_1212_U131;
  assign new_P2_ADD_371_1212_U271 = ~new_P2_ADD_371_1212_U175 | ~new_P2_ADD_371_1212_U57;
  assign new_P2_ADD_371_1212_U272 = ~P2_INSTADDRPOINTER_REG_12_ | ~new_P2_ADD_371_1212_U132;
  assign new_P2_ADD_371_1212_U273 = ~new_P2_ADD_371_1212_U169 | ~new_P2_ADD_371_1212_U48;
  assign new_P2_ADD_371_1212_U274 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_ADD_371_1212_U43;
  assign new_P2_ADD_371_1212_U275 = ~new_P2_R2256_U17 | ~new_P2_ADD_371_1212_U44;
  assign new_P2_ADD_371_1212_U276 = ~P2_INSTADDRPOINTER_REG_7_ | ~new_P2_ADD_371_1212_U43;
  assign new_P2_ADD_371_1212_U277 = ~new_P2_R2256_U17 | ~new_P2_ADD_371_1212_U44;
  assign new_P2_ADD_371_1212_U278 = ~new_P2_ADD_371_1212_U277 | ~new_P2_ADD_371_1212_U276;
  assign new_P2_ADD_371_1212_U279 = ~new_P2_ADD_371_1212_U133 | ~new_P2_ADD_371_1212_U134;
  assign new_P2_ADD_371_1212_U280 = ~new_P2_ADD_371_1212_U160 | ~new_P2_ADD_371_1212_U278;
  assign new_P2_ADD_371_1212_U281 = ~P2_INSTADDRPOINTER_REG_25_ | ~new_P2_ADD_371_1212_U135;
  assign new_P2_ADD_371_1212_U282 = ~new_P2_ADD_371_1212_U178 | ~new_P2_ADD_371_1212_U62;
  assign new_P1_R2027_U5 = ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_R2027_U6 = ~P1_INSTADDRPOINTER_REG_2_;
  assign new_P1_R2027_U7 = ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_R2027_U8 = ~P1_INSTADDRPOINTER_REG_4_;
  assign new_P1_R2027_U9 = ~P1_INSTADDRPOINTER_REG_3_;
  assign new_P1_R2027_U10 = ~P1_INSTADDRPOINTER_REG_1_ | ~P1_INSTADDRPOINTER_REG_2_ | ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_R2027_U11 = ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_R2027_U12 = ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_R2027_U13 = ~new_P1_R2027_U82 | ~new_P1_R2027_U111;
  assign new_P1_R2027_U14 = ~P1_INSTADDRPOINTER_REG_8_;
  assign new_P1_R2027_U15 = ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_R2027_U16 = ~new_P1_R2027_U83 | ~new_P1_R2027_U112;
  assign new_P1_R2027_U17 = ~new_P1_R2027_U84 | ~new_P1_R2027_U118;
  assign new_P1_R2027_U18 = ~P1_INSTADDRPOINTER_REG_9_;
  assign new_P1_R2027_U19 = ~P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_R2027_U20 = ~P1_INSTADDRPOINTER_REG_12_;
  assign new_P1_R2027_U21 = ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_R2027_U22 = ~new_P1_R2027_U85 | ~new_P1_R2027_U120;
  assign new_P1_R2027_U23 = ~P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_R2027_U24 = ~P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_R2027_U25 = ~new_P1_R2027_U86 | ~new_P1_R2027_U113;
  assign new_P1_R2027_U26 = ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_R2027_U27 = ~new_P1_R2027_U87 | ~new_P1_R2027_U119;
  assign new_P1_R2027_U28 = ~P1_INSTADDRPOINTER_REG_16_;
  assign new_P1_R2027_U29 = ~P1_INSTADDRPOINTER_REG_18_;
  assign new_P1_R2027_U30 = ~P1_INSTADDRPOINTER_REG_17_;
  assign new_P1_R2027_U31 = ~new_P1_R2027_U88 | ~new_P1_R2027_U124;
  assign new_P1_R2027_U32 = ~P1_INSTADDRPOINTER_REG_20_;
  assign new_P1_R2027_U33 = ~P1_INSTADDRPOINTER_REG_19_;
  assign new_P1_R2027_U34 = ~new_P1_R2027_U89 | ~new_P1_R2027_U117;
  assign new_P1_R2027_U35 = ~P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_R2027_U36 = ~new_P1_R2027_U90 | ~new_P1_R2027_U114;
  assign new_P1_R2027_U37 = ~P1_INSTADDRPOINTER_REG_22_;
  assign new_P1_R2027_U38 = ~P1_INSTADDRPOINTER_REG_24_;
  assign new_P1_R2027_U39 = ~P1_INSTADDRPOINTER_REG_23_;
  assign new_P1_R2027_U40 = ~new_P1_R2027_U91 | ~new_P1_R2027_U121;
  assign new_P1_R2027_U41 = ~P1_INSTADDRPOINTER_REG_26_;
  assign new_P1_R2027_U42 = ~P1_INSTADDRPOINTER_REG_25_;
  assign new_P1_R2027_U43 = ~new_P1_R2027_U92 | ~new_P1_R2027_U115;
  assign new_P1_R2027_U44 = ~P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_R2027_U45 = ~P1_INSTADDRPOINTER_REG_28_;
  assign new_P1_R2027_U46 = ~new_P1_R2027_U93 | ~new_P1_R2027_U116;
  assign new_P1_R2027_U47 = ~P1_INSTADDRPOINTER_REG_29_;
  assign new_P1_R2027_U48 = ~new_P1_R2027_U94 | ~new_P1_R2027_U122;
  assign new_P1_R2027_U49 = ~new_P1_R2027_U123 | ~P1_INSTADDRPOINTER_REG_29_;
  assign new_P1_R2027_U50 = ~P1_INSTADDRPOINTER_REG_30_;
  assign new_P1_R2027_U51 = ~new_P1_R2027_U142 | ~new_P1_R2027_U141;
  assign new_P1_R2027_U52 = ~new_P1_R2027_U144 | ~new_P1_R2027_U143;
  assign new_P1_R2027_U53 = ~new_P1_R2027_U146 | ~new_P1_R2027_U145;
  assign new_P1_R2027_U54 = ~new_P1_R2027_U148 | ~new_P1_R2027_U147;
  assign new_P1_R2027_U55 = ~new_P1_R2027_U150 | ~new_P1_R2027_U149;
  assign new_P1_R2027_U56 = ~new_P1_R2027_U152 | ~new_P1_R2027_U151;
  assign new_P1_R2027_U57 = ~new_P1_R2027_U154 | ~new_P1_R2027_U153;
  assign new_P1_R2027_U58 = ~new_P1_R2027_U156 | ~new_P1_R2027_U155;
  assign new_P1_R2027_U59 = ~new_P1_R2027_U158 | ~new_P1_R2027_U157;
  assign new_P1_R2027_U60 = ~new_P1_R2027_U160 | ~new_P1_R2027_U159;
  assign new_P1_R2027_U61 = ~new_P1_R2027_U162 | ~new_P1_R2027_U161;
  assign new_P1_R2027_U62 = ~new_P1_R2027_U164 | ~new_P1_R2027_U163;
  assign new_P1_R2027_U63 = ~new_P1_R2027_U166 | ~new_P1_R2027_U165;
  assign new_P1_R2027_U64 = ~new_P1_R2027_U168 | ~new_P1_R2027_U167;
  assign new_P1_R2027_U65 = ~new_P1_R2027_U170 | ~new_P1_R2027_U169;
  assign new_P1_R2027_U66 = ~new_P1_R2027_U172 | ~new_P1_R2027_U171;
  assign new_P1_R2027_U67 = ~new_P1_R2027_U174 | ~new_P1_R2027_U173;
  assign new_P1_R2027_U68 = ~new_P1_R2027_U176 | ~new_P1_R2027_U175;
  assign new_P1_R2027_U69 = ~new_P1_R2027_U178 | ~new_P1_R2027_U177;
  assign new_P1_R2027_U70 = ~new_P1_R2027_U180 | ~new_P1_R2027_U179;
  assign new_P1_R2027_U71 = ~new_P1_R2027_U182 | ~new_P1_R2027_U181;
  assign new_P1_R2027_U72 = ~new_P1_R2027_U184 | ~new_P1_R2027_U183;
  assign new_P1_R2027_U73 = ~new_P1_R2027_U186 | ~new_P1_R2027_U185;
  assign new_P1_R2027_U74 = ~new_P1_R2027_U188 | ~new_P1_R2027_U187;
  assign new_P1_R2027_U75 = ~new_P1_R2027_U190 | ~new_P1_R2027_U189;
  assign new_P1_R2027_U76 = ~new_P1_R2027_U192 | ~new_P1_R2027_U191;
  assign new_P1_R2027_U77 = ~new_P1_R2027_U194 | ~new_P1_R2027_U193;
  assign new_P1_R2027_U78 = ~new_P1_R2027_U196 | ~new_P1_R2027_U195;
  assign new_P1_R2027_U79 = ~new_P1_R2027_U198 | ~new_P1_R2027_U197;
  assign new_P1_R2027_U80 = ~new_P1_R2027_U200 | ~new_P1_R2027_U199;
  assign new_P1_R2027_U81 = ~new_P1_R2027_U202 | ~new_P1_R2027_U201;
  assign new_P1_R2027_U82 = P1_INSTADDRPOINTER_REG_3_ & P1_INSTADDRPOINTER_REG_4_;
  assign new_P1_R2027_U83 = P1_INSTADDRPOINTER_REG_5_ & P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_R2027_U84 = P1_INSTADDRPOINTER_REG_7_ & P1_INSTADDRPOINTER_REG_8_;
  assign new_P1_R2027_U85 = P1_INSTADDRPOINTER_REG_9_ & P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_R2027_U86 = P1_INSTADDRPOINTER_REG_11_ & P1_INSTADDRPOINTER_REG_12_;
  assign new_P1_R2027_U87 = P1_INSTADDRPOINTER_REG_13_ & P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_R2027_U88 = P1_INSTADDRPOINTER_REG_16_ & P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_R2027_U89 = P1_INSTADDRPOINTER_REG_17_ & P1_INSTADDRPOINTER_REG_18_;
  assign new_P1_R2027_U90 = P1_INSTADDRPOINTER_REG_19_ & P1_INSTADDRPOINTER_REG_20_;
  assign new_P1_R2027_U91 = P1_INSTADDRPOINTER_REG_22_ & P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_R2027_U92 = P1_INSTADDRPOINTER_REG_23_ & P1_INSTADDRPOINTER_REG_24_;
  assign new_P1_R2027_U93 = P1_INSTADDRPOINTER_REG_25_ & P1_INSTADDRPOINTER_REG_26_;
  assign new_P1_R2027_U94 = P1_INSTADDRPOINTER_REG_28_ & P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_R2027_U95 = ~new_P1_R2027_U118 | ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_R2027_U96 = ~new_P1_R2027_U112 | ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_R2027_U97 = ~new_P1_R2027_U111 | ~P1_INSTADDRPOINTER_REG_3_;
  assign new_P1_R2027_U98 = ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_R2027_U99 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_R2027_U128;
  assign new_P1_R2027_U100 = ~P1_INSTADDRPOINTER_REG_1_ | ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_R2027_U101 = ~new_P1_R2027_U122 | ~P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_R2027_U102 = ~new_P1_R2027_U116 | ~P1_INSTADDRPOINTER_REG_25_;
  assign new_P1_R2027_U103 = ~new_P1_R2027_U115 | ~P1_INSTADDRPOINTER_REG_23_;
  assign new_P1_R2027_U104 = ~new_P1_R2027_U121 | ~P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_R2027_U105 = ~new_P1_R2027_U114 | ~P1_INSTADDRPOINTER_REG_19_;
  assign new_P1_R2027_U106 = ~new_P1_R2027_U117 | ~P1_INSTADDRPOINTER_REG_17_;
  assign new_P1_R2027_U107 = ~new_P1_R2027_U124 | ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_R2027_U108 = ~new_P1_R2027_U119 | ~P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_R2027_U109 = ~new_P1_R2027_U113 | ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_R2027_U110 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_R2027_U120;
  assign new_P1_R2027_U111 = ~new_P1_R2027_U10;
  assign new_P1_R2027_U112 = ~new_P1_R2027_U13;
  assign new_P1_R2027_U113 = ~new_P1_R2027_U22;
  assign new_P1_R2027_U114 = ~new_P1_R2027_U34;
  assign new_P1_R2027_U115 = ~new_P1_R2027_U40;
  assign new_P1_R2027_U116 = ~new_P1_R2027_U43;
  assign new_P1_R2027_U117 = ~new_P1_R2027_U31;
  assign new_P1_R2027_U118 = ~new_P1_R2027_U16;
  assign new_P1_R2027_U119 = ~new_P1_R2027_U25;
  assign new_P1_R2027_U120 = ~new_P1_R2027_U17;
  assign new_P1_R2027_U121 = ~new_P1_R2027_U36;
  assign new_P1_R2027_U122 = ~new_P1_R2027_U46;
  assign new_P1_R2027_U123 = ~new_P1_R2027_U48;
  assign new_P1_R2027_U124 = ~new_P1_R2027_U27;
  assign new_P1_R2027_U125 = ~new_P1_R2027_U95;
  assign new_P1_R2027_U126 = ~new_P1_R2027_U96;
  assign new_P1_R2027_U127 = ~new_P1_R2027_U97;
  assign new_P1_R2027_U128 = ~new_P1_R2027_U49;
  assign new_P1_R2027_U129 = ~new_P1_R2027_U99;
  assign new_P1_R2027_U130 = ~new_P1_R2027_U100;
  assign new_P1_R2027_U131 = ~new_P1_R2027_U101;
  assign new_P1_R2027_U132 = ~new_P1_R2027_U102;
  assign new_P1_R2027_U133 = ~new_P1_R2027_U103;
  assign new_P1_R2027_U134 = ~new_P1_R2027_U104;
  assign new_P1_R2027_U135 = ~new_P1_R2027_U105;
  assign new_P1_R2027_U136 = ~new_P1_R2027_U106;
  assign new_P1_R2027_U137 = ~new_P1_R2027_U107;
  assign new_P1_R2027_U138 = ~new_P1_R2027_U108;
  assign new_P1_R2027_U139 = ~new_P1_R2027_U109;
  assign new_P1_R2027_U140 = ~new_P1_R2027_U110;
  assign new_P1_R2027_U141 = ~new_P1_R2027_U120 | ~new_P1_R2027_U18;
  assign new_P1_R2027_U142 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_R2027_U17;
  assign new_P1_R2027_U143 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_R2027_U95;
  assign new_P1_R2027_U144 = ~new_P1_R2027_U125 | ~new_P1_R2027_U14;
  assign new_P1_R2027_U145 = ~new_P1_R2027_U118 | ~new_P1_R2027_U15;
  assign new_P1_R2027_U146 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_R2027_U16;
  assign new_P1_R2027_U147 = ~P1_INSTADDRPOINTER_REG_6_ | ~new_P1_R2027_U96;
  assign new_P1_R2027_U148 = ~new_P1_R2027_U126 | ~new_P1_R2027_U11;
  assign new_P1_R2027_U149 = ~new_P1_R2027_U112 | ~new_P1_R2027_U12;
  assign new_P1_R2027_U150 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_R2027_U13;
  assign new_P1_R2027_U151 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_R2027_U97;
  assign new_P1_R2027_U152 = ~new_P1_R2027_U127 | ~new_P1_R2027_U8;
  assign new_P1_R2027_U153 = ~new_P1_R2027_U111 | ~new_P1_R2027_U9;
  assign new_P1_R2027_U154 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_R2027_U10;
  assign new_P1_R2027_U155 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_R2027_U99;
  assign new_P1_R2027_U156 = ~new_P1_R2027_U129 | ~new_P1_R2027_U98;
  assign new_P1_R2027_U157 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_R2027_U49;
  assign new_P1_R2027_U158 = ~new_P1_R2027_U128 | ~new_P1_R2027_U50;
  assign new_P1_R2027_U159 = ~P1_INSTADDRPOINTER_REG_2_ | ~new_P1_R2027_U100;
  assign new_P1_R2027_U160 = ~new_P1_R2027_U130 | ~new_P1_R2027_U6;
  assign new_P1_R2027_U161 = ~new_P1_R2027_U123 | ~new_P1_R2027_U47;
  assign new_P1_R2027_U162 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_R2027_U48;
  assign new_P1_R2027_U163 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_R2027_U101;
  assign new_P1_R2027_U164 = ~new_P1_R2027_U131 | ~new_P1_R2027_U45;
  assign new_P1_R2027_U165 = ~new_P1_R2027_U122 | ~new_P1_R2027_U44;
  assign new_P1_R2027_U166 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_R2027_U46;
  assign new_P1_R2027_U167 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_R2027_U102;
  assign new_P1_R2027_U168 = ~new_P1_R2027_U132 | ~new_P1_R2027_U41;
  assign new_P1_R2027_U169 = ~new_P1_R2027_U116 | ~new_P1_R2027_U42;
  assign new_P1_R2027_U170 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_R2027_U43;
  assign new_P1_R2027_U171 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_R2027_U103;
  assign new_P1_R2027_U172 = ~new_P1_R2027_U133 | ~new_P1_R2027_U38;
  assign new_P1_R2027_U173 = ~new_P1_R2027_U115 | ~new_P1_R2027_U39;
  assign new_P1_R2027_U174 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_R2027_U40;
  assign new_P1_R2027_U175 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_R2027_U104;
  assign new_P1_R2027_U176 = ~new_P1_R2027_U134 | ~new_P1_R2027_U37;
  assign new_P1_R2027_U177 = ~new_P1_R2027_U121 | ~new_P1_R2027_U35;
  assign new_P1_R2027_U178 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_R2027_U36;
  assign new_P1_R2027_U179 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_R2027_U105;
  assign new_P1_R2027_U180 = ~new_P1_R2027_U135 | ~new_P1_R2027_U32;
  assign new_P1_R2027_U181 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_R2027_U7;
  assign new_P1_R2027_U182 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_R2027_U5;
  assign new_P1_R2027_U183 = ~new_P1_R2027_U114 | ~new_P1_R2027_U33;
  assign new_P1_R2027_U184 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_R2027_U34;
  assign new_P1_R2027_U185 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_R2027_U106;
  assign new_P1_R2027_U186 = ~new_P1_R2027_U136 | ~new_P1_R2027_U29;
  assign new_P1_R2027_U187 = ~new_P1_R2027_U117 | ~new_P1_R2027_U30;
  assign new_P1_R2027_U188 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_R2027_U31;
  assign new_P1_R2027_U189 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_R2027_U107;
  assign new_P1_R2027_U190 = ~new_P1_R2027_U137 | ~new_P1_R2027_U28;
  assign new_P1_R2027_U191 = ~new_P1_R2027_U124 | ~new_P1_R2027_U26;
  assign new_P1_R2027_U192 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_R2027_U27;
  assign new_P1_R2027_U193 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_R2027_U108;
  assign new_P1_R2027_U194 = ~new_P1_R2027_U138 | ~new_P1_R2027_U23;
  assign new_P1_R2027_U195 = ~new_P1_R2027_U119 | ~new_P1_R2027_U24;
  assign new_P1_R2027_U196 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_R2027_U25;
  assign new_P1_R2027_U197 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_R2027_U109;
  assign new_P1_R2027_U198 = ~new_P1_R2027_U139 | ~new_P1_R2027_U20;
  assign new_P1_R2027_U199 = ~new_P1_R2027_U113 | ~new_P1_R2027_U21;
  assign new_P1_R2027_U200 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_R2027_U22;
  assign new_P1_R2027_U201 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_R2027_U110;
  assign new_P1_R2027_U202 = ~new_P1_R2027_U140 | ~new_P1_R2027_U19;
  assign new_P1_R2182_U5 = new_P1_R2182_U47 & new_P1_U2740;
  assign new_P1_R2182_U6 = new_P1_R2182_U60 & new_P1_R2182_U16;
  assign new_P1_R2182_U7 = ~new_P1_U2744;
  assign new_P1_R2182_U8 = ~new_P1_U3246;
  assign new_P1_R2182_U9 = ~new_P1_U3246 | ~new_P1_U2744;
  assign new_P1_R2182_U10 = ~new_P1_U2742;
  assign new_P1_R2182_U11 = ~new_P1_U2741;
  assign new_P1_R2182_U12 = ~new_P1_U2740;
  assign new_P1_R2182_U13 = ~new_P1_R2182_U35 | ~new_P1_R2182_U41;
  assign new_P1_R2182_U14 = ~new_P1_U2737;
  assign new_P1_R2182_U15 = ~new_P1_U2738;
  assign new_P1_R2182_U16 = ~new_P1_U2723 | ~new_P1_U2739;
  assign new_P1_R2182_U17 = ~new_P1_U2736;
  assign new_P1_R2182_U18 = ~new_P1_U2735;
  assign new_P1_R2182_U19 = ~new_P1_R2182_U36 | ~new_P1_R2182_U49;
  assign new_P1_R2182_U20 = ~new_P1_U2734;
  assign new_P1_R2182_U21 = ~new_P1_R2182_U37 | ~new_P1_R2182_U46;
  assign new_P1_R2182_U22 = ~new_P1_R2182_U48 | ~new_P1_U2734;
  assign new_P1_R2182_U23 = ~new_P1_U2733;
  assign new_P1_R2182_U24 = ~new_P1_R2182_U64 | ~new_P1_R2182_U63;
  assign new_P1_R2182_U25 = ~new_P1_R2182_U66 | ~new_P1_R2182_U65;
  assign new_P1_R2182_U26 = ~new_P1_R2182_U68 | ~new_P1_R2182_U67;
  assign new_P1_R2182_U27 = ~new_P1_R2182_U72 | ~new_P1_R2182_U71;
  assign new_P1_R2182_U28 = ~new_P1_R2182_U74 | ~new_P1_R2182_U73;
  assign new_P1_R2182_U29 = ~new_P1_R2182_U76 | ~new_P1_R2182_U75;
  assign new_P1_R2182_U30 = ~new_P1_R2182_U78 | ~new_P1_R2182_U77;
  assign new_P1_R2182_U31 = ~new_P1_R2182_U80 | ~new_P1_R2182_U79;
  assign new_P1_R2182_U32 = ~new_P1_R2182_U82 | ~new_P1_R2182_U81;
  assign new_P1_R2182_U33 = ~new_P1_R2182_U84 | ~new_P1_R2182_U83;
  assign new_P1_R2182_U34 = ~new_P1_R2182_U86 | ~new_P1_R2182_U85;
  assign new_P1_R2182_U35 = new_P1_U2742 & new_P1_U2741;
  assign new_P1_R2182_U36 = new_P1_U2738 & new_P1_U2737;
  assign new_P1_R2182_U37 = new_P1_U2735 & new_P1_U2736;
  assign new_P1_R2182_U38 = ~new_P1_U2742 | ~new_P1_R2182_U41;
  assign new_P1_R2182_U39 = ~new_P1_U2732;
  assign new_P1_R2182_U40 = ~new_P1_U2733 | ~new_P1_R2182_U56;
  assign new_P1_R2182_U41 = ~new_P1_R2182_U52 | ~new_P1_R2182_U53;
  assign new_P1_R2182_U42 = new_P1_R2182_U70 & new_P1_R2182_U69;
  assign new_P1_R2182_U43 = ~new_P1_R2182_U46 | ~new_P1_U2736;
  assign new_P1_R2182_U44 = ~new_P1_R2182_U49 | ~new_P1_U2738;
  assign new_P1_R2182_U45 = ~new_P1_R2182_U51 | ~new_P1_R2182_U62;
  assign new_P1_R2182_U46 = ~new_P1_R2182_U19;
  assign new_P1_R2182_U47 = ~new_P1_R2182_U13;
  assign new_P1_R2182_U48 = ~new_P1_R2182_U21;
  assign new_P1_R2182_U49 = ~new_P1_R2182_U16;
  assign new_P1_R2182_U50 = ~new_P1_R2182_U9;
  assign new_P1_R2182_U51 = new_P1_U2743 | new_P1_U2731;
  assign new_P1_R2182_U52 = ~new_P1_U2731 | ~new_P1_U2743;
  assign new_P1_R2182_U53 = ~new_P1_R2182_U50 | ~new_P1_R2182_U51;
  assign new_P1_R2182_U54 = ~new_P1_R2182_U41;
  assign new_P1_R2182_U55 = ~new_P1_R2182_U38;
  assign new_P1_R2182_U56 = ~new_P1_R2182_U22;
  assign new_P1_R2182_U57 = ~new_P1_R2182_U40;
  assign new_P1_R2182_U58 = ~new_P1_R2182_U43;
  assign new_P1_R2182_U59 = ~new_P1_R2182_U44;
  assign new_P1_R2182_U60 = new_P1_U2739 | new_P1_U2723;
  assign new_P1_R2182_U61 = ~new_P1_R2182_U45;
  assign new_P1_R2182_U62 = ~new_P1_U2731 | ~new_P1_U2743;
  assign new_P1_R2182_U63 = ~new_P1_R2182_U47 | ~new_P1_R2182_U12;
  assign new_P1_R2182_U64 = ~new_P1_U2740 | ~new_P1_R2182_U13;
  assign new_P1_R2182_U65 = ~new_P1_U2741 | ~new_P1_R2182_U38;
  assign new_P1_R2182_U66 = ~new_P1_R2182_U55 | ~new_P1_R2182_U11;
  assign new_P1_R2182_U67 = ~new_P1_U2732 | ~new_P1_R2182_U40;
  assign new_P1_R2182_U68 = ~new_P1_R2182_U57 | ~new_P1_R2182_U39;
  assign new_P1_R2182_U69 = ~new_P1_U2742 | ~new_P1_R2182_U41;
  assign new_P1_R2182_U70 = ~new_P1_R2182_U54 | ~new_P1_R2182_U10;
  assign new_P1_R2182_U71 = ~new_P1_U2733 | ~new_P1_R2182_U22;
  assign new_P1_R2182_U72 = ~new_P1_R2182_U56 | ~new_P1_R2182_U23;
  assign new_P1_R2182_U73 = ~new_P1_R2182_U48 | ~new_P1_R2182_U20;
  assign new_P1_R2182_U74 = ~new_P1_U2734 | ~new_P1_R2182_U21;
  assign new_P1_R2182_U75 = ~new_P1_U2735 | ~new_P1_R2182_U43;
  assign new_P1_R2182_U76 = ~new_P1_R2182_U58 | ~new_P1_R2182_U18;
  assign new_P1_R2182_U77 = ~new_P1_R2182_U46 | ~new_P1_R2182_U17;
  assign new_P1_R2182_U78 = ~new_P1_U2736 | ~new_P1_R2182_U19;
  assign new_P1_R2182_U79 = ~new_P1_U2737 | ~new_P1_R2182_U44;
  assign new_P1_R2182_U80 = ~new_P1_R2182_U59 | ~new_P1_R2182_U14;
  assign new_P1_R2182_U81 = ~new_P1_R2182_U49 | ~new_P1_R2182_U15;
  assign new_P1_R2182_U82 = ~new_P1_U2738 | ~new_P1_R2182_U16;
  assign new_P1_R2182_U83 = ~new_P1_R2182_U50 | ~new_P1_R2182_U45;
  assign new_P1_R2182_U84 = ~new_P1_R2182_U61 | ~new_P1_R2182_U9;
  assign new_P1_R2182_U85 = ~new_P1_U3246 | ~new_P1_R2182_U7;
  assign new_P1_R2182_U86 = ~new_P1_U2744 | ~new_P1_R2182_U8;
  assign new_P1_R2144_U5 = new_P1_R2144_U104 & new_P1_R2144_U103;
  assign new_P1_R2144_U6 = new_P1_R2144_U29 & new_P1_R2144_U27 & new_P1_R2144_U36 & new_P1_R2144_U35;
  assign new_P1_R2144_U7 = new_P1_R2144_U104 & new_P1_R2144_U81;
  assign new_P1_R2144_U8 = new_P1_R2144_U138 & new_P1_R2144_U136;
  assign new_P1_R2144_U9 = new_P1_R2144_U128 & new_P1_R2144_U127;
  assign new_P1_R2144_U10 = new_P1_R2144_U82 & new_P1_R2144_U213 & new_P1_R2144_U212;
  assign new_P1_R2144_U11 = ~new_P1_R2144_U144 | ~new_P1_R2144_U146;
  assign new_P1_R2144_U12 = ~new_P1_U2355;
  assign new_P1_R2144_U13 = ~new_P1_U2750;
  assign new_P1_R2144_U14 = ~new_P1_U2751;
  assign new_P1_R2144_U15 = ~new_P1_U2752;
  assign new_P1_R2144_U16 = ~new_P1_U2749;
  assign new_P1_R2144_U17 = ~new_P1_U2745;
  assign new_P1_R2144_U18 = ~new_P1_U2748;
  assign new_P1_R2144_U19 = ~new_P1_U2748 | ~new_P1_R2144_U178;
  assign new_P1_R2144_U20 = ~new_P1_U2747;
  assign new_P1_R2144_U21 = ~new_P1_U2747 | ~new_P1_R2144_U170;
  assign new_P1_R2144_U22 = ~new_P1_U2746;
  assign new_P1_R2144_U23 = ~new_P1_U2746 | ~new_P1_R2144_U173;
  assign new_P1_R2144_U24 = ~new_P1_R2144_U79 | ~new_P1_R2144_U63;
  assign new_P1_R2144_U25 = ~new_P1_R2144_U6 | ~new_P1_R2144_U79;
  assign new_P1_R2144_U26 = ~new_P1_R2144_U65 | ~new_P1_R2144_U141;
  assign new_P1_R2144_U27 = ~new_P1_R2144_U206 | ~new_P1_R2144_U205;
  assign new_P1_R2144_U28 = ~new_P1_R2144_U186 | ~new_P1_R2144_U185;
  assign new_P1_R2144_U29 = ~new_P1_R2144_U203 | ~new_P1_R2144_U202;
  assign new_P1_R2144_U30 = ~new_P1_R2144_U209 | ~new_P1_R2144_U208;
  assign new_P1_R2144_U31 = ~new_P1_R2144_U224 | ~new_P1_R2144_U223;
  assign new_P1_R2144_U32 = ~new_P1_R2144_U221 | ~new_P1_R2144_U220;
  assign new_P1_R2144_U33 = ~new_P1_R2144_U227 | ~new_P1_R2144_U226;
  assign new_P1_R2144_U34 = ~new_P1_R2144_U230 | ~new_P1_R2144_U229;
  assign new_P1_R2144_U35 = ~new_P1_R2144_U233 | ~new_P1_R2144_U232;
  assign new_P1_R2144_U36 = ~new_P1_R2144_U236 | ~new_P1_R2144_U235;
  assign new_P1_R2144_U37 = ~new_P1_R2144_U248 | ~new_P1_R2144_U247;
  assign new_P1_R2144_U38 = ~new_P1_R2144_U250 | ~new_P1_R2144_U249;
  assign new_P1_R2144_U39 = ~new_P1_R2144_U252 | ~new_P1_R2144_U251;
  assign new_P1_R2144_U40 = ~new_P1_R2144_U254 | ~new_P1_R2144_U253;
  assign new_P1_R2144_U41 = ~new_P1_R2144_U256 | ~new_P1_R2144_U255;
  assign new_P1_R2144_U42 = ~new_P1_R2144_U258 | ~new_P1_R2144_U257;
  assign new_P1_R2144_U43 = ~new_P1_R2144_U260 | ~new_P1_R2144_U259;
  assign new_P1_R2144_U44 = new_P1_R2144_U21 & new_P1_R2144_U105;
  assign new_P1_R2144_U45 = ~new_P1_R2144_U217 | ~new_P1_R2144_U216;
  assign new_P1_R2144_U46 = new_P1_R2144_U19 & new_P1_R2144_U106;
  assign new_P1_R2144_U47 = ~new_P1_R2144_U219 | ~new_P1_R2144_U218;
  assign new_P1_R2144_U48 = new_P1_R2144_U162 & new_P1_R2144_U109;
  assign new_P1_R2144_U49 = ~new_P1_R2144_U239 | ~new_P1_R2144_U238;
  assign new_P1_R2144_U50 = ~new_P1_R2144_U246 | ~new_P1_R2144_U245;
  assign new_P1_R2144_U51 = new_P1_R2144_U110 & new_P1_R2144_U109;
  assign new_P1_R2144_U52 = new_P1_R2144_U106 & new_P1_R2144_U105;
  assign new_P1_R2144_U53 = new_P1_R2144_U7 & new_P1_R2144_U52;
  assign new_P1_R2144_U54 = new_P1_R2144_U152 & new_P1_R2144_U153 & new_P1_R2144_U103 & new_P1_R2144_U151;
  assign new_P1_R2144_U55 = new_P1_R2144_U109 & new_P1_R2144_U106;
  assign new_P1_R2144_U56 = new_P1_R2144_U159 & new_P1_R2144_U19;
  assign new_P1_R2144_U57 = new_P1_R2144_U156 & new_P1_R2144_U21;
  assign new_P1_R2144_U58 = new_P1_R2144_U159 & new_P1_R2144_U19 & new_P1_R2144_U21;
  assign new_P1_R2144_U59 = new_P1_R2144_U5 & new_P1_R2144_U105;
  assign new_P1_R2144_U60 = new_P1_R2144_U126 & new_P1_R2144_U21;
  assign new_P1_R2144_U61 = new_P1_R2144_U23 & new_P1_R2144_U81;
  assign new_P1_R2144_U62 = new_P1_R2144_U111 & new_P1_R2144_U110;
  assign new_P1_R2144_U63 = new_P1_R2144_U6 & new_P1_R2144_U64;
  assign new_P1_R2144_U64 = new_P1_R2144_U32 & new_P1_R2144_U31 & new_P1_R2144_U34 & new_P1_R2144_U33;
  assign new_P1_R2144_U65 = new_P1_R2144_U34 & new_P1_R2144_U33;
  assign new_P1_R2144_U66 = new_P1_R2144_U29 & new_P1_R2144_U36 & new_P1_R2144_U27;
  assign new_P1_R2144_U67 = new_P1_R2144_U29 & new_P1_R2144_U27;
  assign new_P1_R2144_U68 = ~new_P1_U2762;
  assign new_P1_R2144_U69 = ~new_P1_U2761;
  assign new_P1_R2144_U70 = ~new_P1_U2763;
  assign new_P1_R2144_U71 = ~new_P1_U2764;
  assign new_P1_R2144_U72 = ~new_P1_U2766;
  assign new_P1_R2144_U73 = ~new_P1_U2767;
  assign new_P1_R2144_U74 = ~new_P1_U2768;
  assign new_P1_R2144_U75 = ~new_P1_U2765;
  assign new_P1_R2144_U76 = ~new_P1_U2760;
  assign new_P1_R2144_U77 = ~new_P1_U2759;
  assign new_P1_R2144_U78 = ~new_P1_R2144_U29 | ~new_P1_R2144_U79;
  assign new_P1_R2144_U79 = ~new_P1_R2144_U99 | ~new_P1_R2144_U54;
  assign new_P1_R2144_U80 = new_P1_R2144_U211 & new_P1_R2144_U210;
  assign new_P1_R2144_U81 = ~new_P1_R2144_U22 | ~new_P1_R2144_U165 | ~new_P1_R2144_U164;
  assign new_P1_R2144_U82 = new_P1_R2144_U215 & new_P1_R2144_U214;
  assign new_P1_R2144_U83 = ~new_P1_R2144_U56 | ~new_P1_R2144_U158;
  assign new_P1_R2144_U84 = ~new_P1_R2144_U111 | ~new_P1_R2144_U118;
  assign new_P1_R2144_U85 = ~new_P1_U2754;
  assign new_P1_R2144_U86 = ~new_P1_U2753;
  assign new_P1_R2144_U87 = ~new_P1_U2755;
  assign new_P1_R2144_U88 = ~new_P1_U2756;
  assign new_P1_R2144_U89 = ~new_P1_U2757;
  assign new_P1_R2144_U90 = ~new_P1_U2758;
  assign new_P1_R2144_U91 = ~new_P1_R2144_U100 | ~new_P1_R2144_U132;
  assign new_P1_R2144_U92 = new_P1_R2144_U241 & new_P1_R2144_U240;
  assign new_P1_R2144_U93 = ~new_P1_R2144_U129 | ~new_P1_R2144_U113;
  assign new_P1_R2144_U94 = ~new_P1_R2144_U143 | ~new_P1_R2144_U32;
  assign new_P1_R2144_U95 = ~new_P1_R2144_U141 | ~new_P1_R2144_U34;
  assign new_P1_R2144_U96 = ~new_P1_R2144_U79 | ~new_P1_R2144_U66;
  assign new_P1_R2144_U97 = ~new_P1_R2144_U67 | ~new_P1_R2144_U79;
  assign new_P1_R2144_U98 = ~new_P1_R2144_U113 | ~new_P1_R2144_U112;
  assign new_P1_R2144_U99 = ~new_P1_R2144_U53 | ~new_P1_R2144_U84;
  assign new_P1_R2144_U100 = ~new_P1_U2751 | ~new_P1_R2144_U28;
  assign new_P1_R2144_U101 = ~new_P1_R2144_U24;
  assign new_P1_R2144_U102 = ~new_P1_R2144_U81;
  assign new_P1_R2144_U103 = ~new_P1_U2745 | ~new_P1_R2144_U181;
  assign new_P1_R2144_U104 = ~new_P1_R2144_U17 | ~new_P1_R2144_U167 | ~new_P1_R2144_U166;
  assign new_P1_R2144_U105 = ~new_P1_R2144_U20 | ~new_P1_R2144_U175 | ~new_P1_R2144_U174;
  assign new_P1_R2144_U106 = ~new_P1_R2144_U18 | ~new_P1_R2144_U201 | ~new_P1_R2144_U200;
  assign new_P1_R2144_U107 = ~new_P1_R2144_U21;
  assign new_P1_R2144_U108 = ~new_P1_R2144_U23;
  assign new_P1_R2144_U109 = ~new_P1_R2144_U13 | ~new_P1_R2144_U194 | ~new_P1_R2144_U193;
  assign new_P1_R2144_U110 = ~new_P1_R2144_U16 | ~new_P1_R2144_U196 | ~new_P1_R2144_U195;
  assign new_P1_R2144_U111 = ~new_P1_U2749 | ~new_P1_R2144_U199;
  assign new_P1_R2144_U112 = ~new_P1_R2144_U15 | ~new_P1_R2144_U189 | ~new_P1_R2144_U188;
  assign new_P1_R2144_U113 = ~new_P1_U2752 | ~new_P1_R2144_U192;
  assign new_P1_R2144_U114 = ~new_P1_R2144_U187 | ~new_P1_R2144_U14;
  assign new_P1_R2144_U115 = ~new_P1_U2355 | ~new_P1_R2144_U112;
  assign new_P1_R2144_U116 = ~new_P1_U2750 | ~new_P1_R2144_U184;
  assign new_P1_R2144_U117 = ~new_P1_R2144_U155 | ~new_P1_R2144_U157;
  assign new_P1_R2144_U118 = ~new_P1_R2144_U51 | ~new_P1_R2144_U117;
  assign new_P1_R2144_U119 = ~new_P1_R2144_U84;
  assign new_P1_R2144_U120 = ~new_P1_R2144_U19;
  assign new_P1_R2144_U121 = ~new_P1_R2144_U79;
  assign new_P1_R2144_U122 = ~new_P1_R2144_U78;
  assign new_P1_R2144_U123 = ~new_P1_R2144_U83;
  assign new_P1_R2144_U124 = ~new_P1_R2144_U83 | ~new_P1_R2144_U105;
  assign new_P1_R2144_U125 = ~new_P1_R2144_U21 | ~new_P1_R2144_U124;
  assign new_P1_R2144_U126 = ~new_P1_R2144_U23 | ~new_P1_R2144_U81;
  assign new_P1_R2144_U127 = ~new_P1_R2144_U60 | ~new_P1_R2144_U124;
  assign new_P1_R2144_U128 = ~new_P1_R2144_U61 | ~new_P1_R2144_U125;
  assign new_P1_R2144_U129 = ~new_P1_U2355 | ~new_P1_R2144_U112;
  assign new_P1_R2144_U130 = ~new_P1_R2144_U93;
  assign new_P1_R2144_U131 = ~new_P1_R2144_U187 | ~new_P1_R2144_U14;
  assign new_P1_R2144_U132 = ~new_P1_R2144_U131 | ~new_P1_R2144_U93;
  assign new_P1_R2144_U133 = ~new_P1_R2144_U91;
  assign new_P1_R2144_U134 = ~new_P1_R2144_U91 | ~new_P1_R2144_U109;
  assign new_P1_R2144_U135 = ~new_P1_R2144_U134 | ~new_P1_R2144_U116;
  assign new_P1_R2144_U136 = ~new_P1_R2144_U62 | ~new_P1_R2144_U135;
  assign new_P1_R2144_U137 = ~new_P1_R2144_U161 | ~new_P1_R2144_U110;
  assign new_P1_R2144_U138 = ~new_P1_R2144_U137 | ~new_P1_R2144_U134 | ~new_P1_R2144_U116;
  assign new_P1_R2144_U139 = ~new_P1_R2144_U97;
  assign new_P1_R2144_U140 = ~new_P1_R2144_U96;
  assign new_P1_R2144_U141 = ~new_P1_R2144_U25;
  assign new_P1_R2144_U142 = ~new_P1_R2144_U95;
  assign new_P1_R2144_U143 = ~new_P1_R2144_U26;
  assign new_P1_R2144_U144 = ~new_P1_U2355 | ~new_P1_R2144_U24;
  assign new_P1_R2144_U145 = ~new_P1_R2144_U144;
  assign new_P1_R2144_U146 = ~new_P1_R2144_U101 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U147 = ~new_P1_R2144_U94;
  assign new_P1_R2144_U148 = ~new_P1_R2144_U98;
  assign new_P1_R2144_U149 = ~new_P1_R2144_U21 | ~new_P1_R2144_U105;
  assign new_P1_R2144_U150 = ~new_P1_R2144_U19 | ~new_P1_R2144_U106;
  assign new_P1_R2144_U151 = ~new_P1_R2144_U7 | ~new_P1_R2144_U120 | ~new_P1_R2144_U105;
  assign new_P1_R2144_U152 = ~new_P1_R2144_U107 | ~new_P1_R2144_U7;
  assign new_P1_R2144_U153 = ~new_P1_R2144_U108 | ~new_P1_R2144_U7;
  assign new_P1_R2144_U154 = ~new_P1_R2144_U100 | ~new_P1_R2144_U113 | ~new_P1_R2144_U115;
  assign new_P1_R2144_U155 = ~new_P1_R2144_U154 | ~new_P1_R2144_U114;
  assign new_P1_R2144_U156 = ~new_P1_R2144_U104 | ~new_P1_R2144_U103;
  assign new_P1_R2144_U157 = ~new_P1_U2750 | ~new_P1_R2144_U184;
  assign new_P1_R2144_U158 = ~new_P1_R2144_U55 | ~new_P1_R2144_U117 | ~new_P1_R2144_U110;
  assign new_P1_R2144_U159 = ~new_P1_R2144_U199 | ~new_P1_U2749 | ~new_P1_R2144_U106;
  assign new_P1_R2144_U160 = ~new_P1_R2144_U58 | ~new_P1_R2144_U158;
  assign new_P1_R2144_U161 = ~new_P1_U2749 | ~new_P1_R2144_U199;
  assign new_P1_R2144_U162 = ~new_P1_U2750 | ~new_P1_R2144_U184;
  assign new_P1_R2144_U163 = ~new_P1_R2144_U116 | ~new_P1_R2144_U109;
  assign new_P1_R2144_U164 = ~new_P1_U2355 | ~new_P1_R2144_U68;
  assign new_P1_R2144_U165 = ~new_P1_U2762 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U166 = ~new_P1_U2355 | ~new_P1_R2144_U69;
  assign new_P1_R2144_U167 = ~new_P1_U2761 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U168 = ~new_P1_U2355 | ~new_P1_R2144_U70;
  assign new_P1_R2144_U169 = ~new_P1_U2763 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U170 = ~new_P1_R2144_U169 | ~new_P1_R2144_U168;
  assign new_P1_R2144_U171 = ~new_P1_U2355 | ~new_P1_R2144_U68;
  assign new_P1_R2144_U172 = ~new_P1_U2762 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U173 = ~new_P1_R2144_U172 | ~new_P1_R2144_U171;
  assign new_P1_R2144_U174 = ~new_P1_U2355 | ~new_P1_R2144_U70;
  assign new_P1_R2144_U175 = ~new_P1_U2763 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U176 = ~new_P1_U2355 | ~new_P1_R2144_U71;
  assign new_P1_R2144_U177 = ~new_P1_U2764 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U178 = ~new_P1_R2144_U177 | ~new_P1_R2144_U176;
  assign new_P1_R2144_U179 = ~new_P1_U2355 | ~new_P1_R2144_U69;
  assign new_P1_R2144_U180 = ~new_P1_U2761 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U181 = ~new_P1_R2144_U180 | ~new_P1_R2144_U179;
  assign new_P1_R2144_U182 = ~new_P1_U2355 | ~new_P1_R2144_U72;
  assign new_P1_R2144_U183 = ~new_P1_U2766 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U184 = ~new_P1_R2144_U183 | ~new_P1_R2144_U182;
  assign new_P1_R2144_U185 = ~new_P1_U2355 | ~new_P1_R2144_U73;
  assign new_P1_R2144_U186 = ~new_P1_U2767 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U187 = ~new_P1_R2144_U28;
  assign new_P1_R2144_U188 = ~new_P1_U2355 | ~new_P1_R2144_U74;
  assign new_P1_R2144_U189 = ~new_P1_U2768 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U190 = ~new_P1_U2355 | ~new_P1_R2144_U74;
  assign new_P1_R2144_U191 = ~new_P1_U2768 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U192 = ~new_P1_R2144_U191 | ~new_P1_R2144_U190;
  assign new_P1_R2144_U193 = ~new_P1_U2355 | ~new_P1_R2144_U72;
  assign new_P1_R2144_U194 = ~new_P1_U2766 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U195 = ~new_P1_U2355 | ~new_P1_R2144_U75;
  assign new_P1_R2144_U196 = ~new_P1_U2765 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U197 = ~new_P1_U2355 | ~new_P1_R2144_U75;
  assign new_P1_R2144_U198 = ~new_P1_U2765 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U199 = ~new_P1_R2144_U198 | ~new_P1_R2144_U197;
  assign new_P1_R2144_U200 = ~new_P1_U2355 | ~new_P1_R2144_U71;
  assign new_P1_R2144_U201 = ~new_P1_U2764 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U202 = ~new_P1_U2355 | ~new_P1_R2144_U76;
  assign new_P1_R2144_U203 = ~new_P1_U2760 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U204 = ~new_P1_R2144_U29;
  assign new_P1_R2144_U205 = ~new_P1_U2355 | ~new_P1_R2144_U77;
  assign new_P1_R2144_U206 = ~new_P1_U2759 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U207 = ~new_P1_R2144_U27;
  assign new_P1_R2144_U208 = ~new_P1_R2144_U122 | ~new_P1_R2144_U207;
  assign new_P1_R2144_U209 = ~new_P1_R2144_U27 | ~new_P1_R2144_U78;
  assign new_P1_R2144_U210 = ~new_P1_R2144_U121 | ~new_P1_R2144_U204;
  assign new_P1_R2144_U211 = ~new_P1_R2144_U29 | ~new_P1_R2144_U79;
  assign new_P1_R2144_U212 = ~new_P1_R2144_U23 | ~new_P1_R2144_U57 | ~new_P1_R2144_U124;
  assign new_P1_R2144_U213 = ~new_P1_R2144_U5 | ~new_P1_R2144_U108;
  assign new_P1_R2144_U214 = ~new_P1_R2144_U102 | ~new_P1_R2144_U156;
  assign new_P1_R2144_U215 = ~new_P1_R2144_U81 | ~new_P1_R2144_U59 | ~new_P1_R2144_U160;
  assign new_P1_R2144_U216 = ~new_P1_R2144_U149 | ~new_P1_R2144_U83;
  assign new_P1_R2144_U217 = ~new_P1_R2144_U44 | ~new_P1_R2144_U123;
  assign new_P1_R2144_U218 = ~new_P1_R2144_U150 | ~new_P1_R2144_U84;
  assign new_P1_R2144_U219 = ~new_P1_R2144_U46 | ~new_P1_R2144_U119;
  assign new_P1_R2144_U220 = ~new_P1_U2355 | ~new_P1_R2144_U85;
  assign new_P1_R2144_U221 = ~new_P1_U2754 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U222 = ~new_P1_R2144_U32;
  assign new_P1_R2144_U223 = ~new_P1_U2355 | ~new_P1_R2144_U86;
  assign new_P1_R2144_U224 = ~new_P1_U2753 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U225 = ~new_P1_R2144_U31;
  assign new_P1_R2144_U226 = ~new_P1_U2355 | ~new_P1_R2144_U87;
  assign new_P1_R2144_U227 = ~new_P1_U2755 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U228 = ~new_P1_R2144_U33;
  assign new_P1_R2144_U229 = ~new_P1_U2355 | ~new_P1_R2144_U88;
  assign new_P1_R2144_U230 = ~new_P1_U2756 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U231 = ~new_P1_R2144_U34;
  assign new_P1_R2144_U232 = ~new_P1_U2355 | ~new_P1_R2144_U89;
  assign new_P1_R2144_U233 = ~new_P1_U2757 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U234 = ~new_P1_R2144_U35;
  assign new_P1_R2144_U235 = ~new_P1_U2355 | ~new_P1_R2144_U90;
  assign new_P1_R2144_U236 = ~new_P1_U2758 | ~new_P1_R2144_U12;
  assign new_P1_R2144_U237 = ~new_P1_R2144_U36;
  assign new_P1_R2144_U238 = ~new_P1_R2144_U163 | ~new_P1_R2144_U91;
  assign new_P1_R2144_U239 = ~new_P1_R2144_U48 | ~new_P1_R2144_U133;
  assign new_P1_R2144_U240 = ~new_P1_R2144_U187 | ~new_P1_U2751;
  assign new_P1_R2144_U241 = ~new_P1_R2144_U28 | ~new_P1_R2144_U14;
  assign new_P1_R2144_U242 = ~new_P1_R2144_U187 | ~new_P1_U2751;
  assign new_P1_R2144_U243 = ~new_P1_R2144_U28 | ~new_P1_R2144_U14;
  assign new_P1_R2144_U244 = ~new_P1_R2144_U243 | ~new_P1_R2144_U242;
  assign new_P1_R2144_U245 = ~new_P1_R2144_U92 | ~new_P1_R2144_U93;
  assign new_P1_R2144_U246 = ~new_P1_R2144_U130 | ~new_P1_R2144_U244;
  assign new_P1_R2144_U247 = ~new_P1_R2144_U147 | ~new_P1_R2144_U225;
  assign new_P1_R2144_U248 = ~new_P1_R2144_U31 | ~new_P1_R2144_U94;
  assign new_P1_R2144_U249 = ~new_P1_R2144_U222 | ~new_P1_R2144_U143;
  assign new_P1_R2144_U250 = ~new_P1_R2144_U32 | ~new_P1_R2144_U26;
  assign new_P1_R2144_U251 = ~new_P1_R2144_U142 | ~new_P1_R2144_U228;
  assign new_P1_R2144_U252 = ~new_P1_R2144_U33 | ~new_P1_R2144_U95;
  assign new_P1_R2144_U253 = ~new_P1_R2144_U231 | ~new_P1_R2144_U141;
  assign new_P1_R2144_U254 = ~new_P1_R2144_U34 | ~new_P1_R2144_U25;
  assign new_P1_R2144_U255 = ~new_P1_R2144_U140 | ~new_P1_R2144_U234;
  assign new_P1_R2144_U256 = ~new_P1_R2144_U35 | ~new_P1_R2144_U96;
  assign new_P1_R2144_U257 = ~new_P1_R2144_U139 | ~new_P1_R2144_U237;
  assign new_P1_R2144_U258 = ~new_P1_R2144_U36 | ~new_P1_R2144_U97;
  assign new_P1_R2144_U259 = ~new_P1_U2355 | ~new_P1_R2144_U98;
  assign new_P1_R2144_U260 = ~new_P1_R2144_U148 | ~new_P1_R2144_U12;
  assign new_P1_R2278_U5 = new_P1_R2278_U466 & new_P1_R2278_U327;
  assign new_P1_R2278_U6 = new_P1_R2278_U292 & new_P1_R2278_U288;
  assign new_P1_R2278_U7 = new_P1_R2278_U6 & new_P1_R2278_U295;
  assign new_P1_R2278_U8 = new_P1_R2278_U305 & new_P1_R2278_U302 & new_P1_R2278_U298;
  assign new_P1_R2278_U9 = new_P1_R2278_U8 & new_P1_R2278_U308;
  assign new_P1_R2278_U10 = new_P1_R2278_U315 & new_P1_R2278_U313 & new_P1_R2278_U311;
  assign new_P1_R2278_U11 = new_P1_R2278_U134 & new_P1_R2278_U10;
  assign new_P1_R2278_U12 = new_P1_R2278_U295 & new_P1_R2278_U292;
  assign new_P1_R2278_U13 = new_P1_R2278_U9 & new_P1_R2278_U321;
  assign new_P1_R2278_U14 = new_P1_R2278_U463 & new_P1_R2278_U462;
  assign new_P1_R2278_U15 = new_P1_R2278_U344 & new_P1_R2278_U342;
  assign new_P1_R2278_U16 = new_P1_R2278_U467 & new_P1_R2278_U468 & new_P1_R2278_U188 & new_P1_R2278_U375;
  assign new_P1_R2278_U17 = new_P1_R2278_U272 & new_P1_R2278_U270;
  assign new_P1_R2278_U18 = new_P1_R2278_U268 & new_P1_R2278_U266;
  assign new_P1_R2278_U19 = ~new_P1_R2278_U214 | ~new_P1_R2278_U429;
  assign new_P1_R2278_U20 = new_P1_R2278_U414 & new_P1_R2278_U335;
  assign new_P1_R2278_U21 = ~P1_INSTADDRPOINTER_REG_8_;
  assign new_P1_R2278_U22 = ~new_P1_U2792;
  assign new_P1_R2278_U23 = ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_R2278_U24 = ~new_P1_U2793;
  assign new_P1_R2278_U25 = ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_R2278_U26 = ~new_P1_U2794;
  assign new_P1_R2278_U27 = ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_R2278_U28 = ~new_P1_U2795;
  assign new_P1_R2278_U29 = ~new_P1_U2800;
  assign new_P1_R2278_U30 = ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_R2278_U31 = ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_R2278_U32 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_U2800;
  assign new_P1_R2278_U33 = ~new_P1_U2799;
  assign new_P1_R2278_U34 = ~P1_INSTADDRPOINTER_REG_2_;
  assign new_P1_R2278_U35 = ~new_P1_U2798;
  assign new_P1_R2278_U36 = ~P1_INSTADDRPOINTER_REG_3_;
  assign new_P1_R2278_U37 = ~new_P1_U2797;
  assign new_P1_R2278_U38 = ~P1_INSTADDRPOINTER_REG_4_;
  assign new_P1_R2278_U39 = ~new_P1_U2796;
  assign new_P1_R2278_U40 = ~new_P1_R2278_U43 | ~new_P1_R2278_U250;
  assign new_P1_R2278_U41 = ~new_P1_R2278_U253 | ~new_P1_R2278_U254 | ~new_P1_R2278_U252;
  assign new_P1_R2278_U42 = ~new_P1_R2278_U246 | ~new_P1_R2278_U245;
  assign new_P1_R2278_U43 = ~new_P1_R2278_U42 | ~new_P1_R2278_U248;
  assign new_P1_R2278_U44 = ~P1_INSTADDRPOINTER_REG_25_;
  assign new_P1_R2278_U45 = ~new_P1_U2775;
  assign new_P1_R2278_U46 = ~P1_INSTADDRPOINTER_REG_26_;
  assign new_P1_R2278_U47 = ~new_P1_U2774;
  assign new_P1_R2278_U48 = ~P1_INSTADDRPOINTER_REG_24_;
  assign new_P1_R2278_U49 = ~new_P1_U2776;
  assign new_P1_R2278_U50 = ~P1_INSTADDRPOINTER_REG_23_;
  assign new_P1_R2278_U51 = ~new_P1_U2777;
  assign new_P1_R2278_U52 = ~P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_R2278_U53 = ~new_P1_U2779;
  assign new_P1_R2278_U54 = ~P1_INSTADDRPOINTER_REG_20_;
  assign new_P1_R2278_U55 = ~new_P1_U2780;
  assign new_P1_R2278_U56 = ~P1_INSTADDRPOINTER_REG_19_;
  assign new_P1_R2278_U57 = ~new_P1_U2781;
  assign new_P1_R2278_U58 = ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_R2278_U59 = ~new_P1_U2789;
  assign new_P1_R2278_U60 = ~P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_R2278_U61 = ~new_P1_U2790;
  assign new_P1_R2278_U62 = ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_R2278_U63 = ~new_P1_U2785;
  assign new_P1_R2278_U64 = ~P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_R2278_U65 = ~new_P1_U2787;
  assign new_P1_R2278_U66 = ~P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_R2278_U67 = ~new_P1_U2786;
  assign new_P1_R2278_U68 = ~new_P1_U2788 | ~P1_INSTADDRPOINTER_REG_12_;
  assign new_P1_R2278_U69 = ~P1_INSTADDRPOINTER_REG_16_;
  assign new_P1_R2278_U70 = ~new_P1_U2784;
  assign new_P1_R2278_U71 = ~P1_INSTADDRPOINTER_REG_17_;
  assign new_P1_R2278_U72 = ~new_P1_U2783;
  assign new_P1_R2278_U73 = ~new_P1_R2278_U308 | ~new_P1_R2278_U359 | ~new_P1_R2278_U12 | ~new_P1_R2278_U8;
  assign new_P1_R2278_U74 = ~P1_INSTADDRPOINTER_REG_22_;
  assign new_P1_R2278_U75 = ~new_P1_U2778;
  assign new_P1_R2278_U76 = ~new_P1_U2778 | ~P1_INSTADDRPOINTER_REG_22_;
  assign new_P1_R2278_U77 = ~P1_INSTADDRPOINTER_REG_18_;
  assign new_P1_R2278_U78 = ~new_P1_U2782;
  assign new_P1_R2278_U79 = ~new_P1_U2782 | ~P1_INSTADDRPOINTER_REG_18_;
  assign new_P1_R2278_U80 = ~new_P1_R2278_U144 | ~new_P1_R2278_U8;
  assign new_P1_R2278_U81 = ~new_P1_U2772;
  assign new_P1_R2278_U82 = ~P1_INSTADDRPOINTER_REG_28_;
  assign new_P1_R2278_U83 = ~P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_R2278_U84 = ~new_P1_U2773;
  assign new_P1_R2278_U85 = ~new_P1_U2773 | ~P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_R2278_U86 = ~new_P1_R2278_U379 | ~new_P1_R2278_U322;
  assign new_P1_R2278_U87 = ~new_P1_R2278_U93 | ~new_P1_R2278_U392 | ~new_P1_R2278_U92;
  assign new_P1_R2278_U88 = ~new_P1_U2770;
  assign new_P1_R2278_U89 = ~P1_INSTADDRPOINTER_REG_30_;
  assign new_P1_R2278_U90 = ~new_P1_U2771;
  assign new_P1_R2278_U91 = ~P1_INSTADDRPOINTER_REG_29_;
  assign new_P1_R2278_U92 = ~new_P1_R2278_U143 | ~new_P1_R2278_U11;
  assign new_P1_R2278_U93 = ~new_P1_R2278_U377 | ~new_P1_R2278_U11 | ~new_P1_R2278_U321;
  assign new_P1_R2278_U94 = ~new_P1_R2278_U132 | ~new_P1_R2278_U372;
  assign new_P1_R2278_U95 = ~new_P1_R2278_U136 | ~new_P1_R2278_U368;
  assign new_P1_R2278_U96 = ~new_P1_R2278_U378 | ~new_P1_R2278_U11 | ~new_P1_R2278_U321;
  assign new_P1_R2278_U97 = ~new_P1_R2278_U229 | ~new_P1_R2278_U331;
  assign new_P1_R2278_U98 = ~new_P1_R2278_U138 | ~new_P1_R2278_U354;
  assign new_P1_R2278_U99 = ~new_P1_R2278_U610 | ~new_P1_R2278_U609;
  assign new_P1_R2278_U100 = new_P1_R2278_U262 & new_P1_R2278_U261;
  assign new_P1_R2278_U101 = ~new_P1_R2278_U431 | ~new_P1_R2278_U430;
  assign new_P1_R2278_U102 = ~new_P1_R2278_U438 | ~new_P1_R2278_U437;
  assign new_P1_R2278_U103 = ~new_P1_R2278_U445 | ~new_P1_R2278_U444;
  assign new_P1_R2278_U104 = ~new_P1_R2278_U454 | ~new_P1_R2278_U453;
  assign new_P1_R2278_U105 = ~new_P1_R2278_U461 | ~new_P1_R2278_U460;
  assign new_P1_R2278_U106 = ~new_P1_R2278_U477 | ~new_P1_R2278_U476;
  assign new_P1_R2278_U107 = ~new_P1_R2278_U484 | ~new_P1_R2278_U483;
  assign new_P1_R2278_U108 = ~new_P1_R2278_U491 | ~new_P1_R2278_U490;
  assign new_P1_R2278_U109 = ~new_P1_R2278_U498 | ~new_P1_R2278_U497;
  assign new_P1_R2278_U110 = ~new_P1_R2278_U505 | ~new_P1_R2278_U504;
  assign new_P1_R2278_U111 = ~new_P1_R2278_U512 | ~new_P1_R2278_U511;
  assign new_P1_R2278_U112 = ~new_P1_R2278_U519 | ~new_P1_R2278_U518;
  assign new_P1_R2278_U113 = ~new_P1_R2278_U526 | ~new_P1_R2278_U525;
  assign new_P1_R2278_U114 = ~new_P1_R2278_U533 | ~new_P1_R2278_U532;
  assign new_P1_R2278_U115 = ~new_P1_R2278_U540 | ~new_P1_R2278_U539;
  assign new_P1_R2278_U116 = ~new_P1_R2278_U547 | ~new_P1_R2278_U546;
  assign new_P1_R2278_U117 = ~new_P1_R2278_U554 | ~new_P1_R2278_U553;
  assign new_P1_R2278_U118 = ~new_P1_R2278_U566 | ~new_P1_R2278_U565;
  assign new_P1_R2278_U119 = ~new_P1_R2278_U573 | ~new_P1_R2278_U572;
  assign new_P1_R2278_U120 = ~new_P1_R2278_U580 | ~new_P1_R2278_U579;
  assign new_P1_R2278_U121 = ~new_P1_R2278_U587 | ~new_P1_R2278_U586;
  assign new_P1_R2278_U122 = ~new_P1_R2278_U594 | ~new_P1_R2278_U593;
  assign new_P1_R2278_U123 = ~new_P1_R2278_U599 | ~new_P1_R2278_U598;
  assign new_P1_R2278_U124 = new_P1_R2278_U68 & new_P1_R2278_U281;
  assign new_P1_R2278_U125 = ~new_P1_R2278_U601 | ~new_P1_R2278_U600;
  assign new_P1_R2278_U126 = ~new_P1_R2278_U608 | ~new_P1_R2278_U607;
  assign new_P1_R2278_U127 = P1_INSTADDRPOINTER_REG_7_ & new_P1_U2793;
  assign new_P1_R2278_U128 = new_P1_R2278_U258 & new_P1_R2278_U254;
  assign new_P1_R2278_U129 = new_P1_R2278_U352 & new_P1_R2278_U259;
  assign new_P1_R2278_U130 = P1_INSTADDRPOINTER_REG_23_ & new_P1_U2777;
  assign new_P1_R2278_U131 = new_P1_R2278_U318 & new_P1_R2278_U316;
  assign new_P1_R2278_U132 = new_P1_R2278_U321 & new_P1_R2278_U319 & new_P1_R2278_U317;
  assign new_P1_R2278_U133 = P1_INSTADDRPOINTER_REG_19_ & new_P1_U2781;
  assign new_P1_R2278_U134 = new_P1_R2278_U319 & new_P1_R2278_U317;
  assign new_P1_R2278_U135 = new_P1_R2278_U321 & new_P1_R2278_U308;
  assign new_P1_R2278_U136 = new_P1_R2278_U11 & new_P1_R2278_U135;
  assign new_P1_R2278_U137 = new_P1_R2278_U273 & new_P1_R2278_U259 & new_P1_R2278_U228;
  assign new_P1_R2278_U138 = new_P1_R2278_U389 & new_P1_R2278_U276;
  assign new_P1_R2278_U139 = new_P1_R2278_U357 & new_P1_R2278_U140;
  assign new_P1_R2278_U140 = new_P1_R2278_U284 & new_P1_R2278_U281 & new_P1_R2278_U283;
  assign new_P1_R2278_U141 = new_P1_R2278_U286 & new_P1_R2278_U410;
  assign new_P1_R2278_U142 = new_P1_R2278_U7 & new_P1_R2278_U13;
  assign new_P1_R2278_U143 = new_P1_R2278_U309 & new_P1_R2278_U321;
  assign new_P1_R2278_U144 = new_P1_R2278_U296 & new_P1_R2278_U308;
  assign new_P1_R2278_U145 = new_P1_R2278_U95 & new_P1_R2278_U94;
  assign new_P1_R2278_U146 = new_P1_R2278_U401 & new_P1_R2278_U96;
  assign new_P1_R2278_U147 = new_P1_R2278_U324 & new_P1_R2278_U5;
  assign new_P1_R2278_U148 = new_P1_R2278_U317 & new_P1_R2278_U319 & new_P1_R2278_U324 & new_P1_R2278_U321;
  assign new_P1_R2278_U149 = new_P1_R2278_U324 & new_P1_R2278_U321 & new_P1_R2278_U308;
  assign new_P1_R2278_U150 = new_P1_R2278_U11 & new_P1_R2278_U149;
  assign new_P1_R2278_U151 = new_P1_R2278_U286 & new_P1_R2278_U412;
  assign new_P1_R2278_U152 = new_P1_R2278_U11 & new_P1_R2278_U324;
  assign new_P1_R2278_U153 = new_P1_R2278_U7 & new_P1_R2278_U13;
  assign new_P1_R2278_U154 = new_P1_R2278_U324 & new_P1_R2278_U321;
  assign new_P1_R2278_U155 = new_P1_R2278_U156 & new_P1_R2278_U398 & new_P1_R2278_U395 & new_P1_R2278_U394 & new_P1_R2278_U393;
  assign new_P1_R2278_U156 = new_P1_R2278_U399 & new_P1_R2278_U14 & new_P1_R2278_U400;
  assign new_P1_R2278_U157 = new_P1_R2278_U11 & new_P1_R2278_U324;
  assign new_P1_R2278_U158 = new_P1_R2278_U7 & new_P1_R2278_U13;
  assign new_P1_R2278_U159 = new_P1_R2278_U404 & new_P1_R2278_U403 & new_P1_R2278_U187;
  assign new_P1_R2278_U160 = new_P1_R2278_U286 & new_P1_R2278_U417;
  assign new_P1_R2278_U161 = new_P1_R2278_U9 & new_P1_R2278_U7;
  assign new_P1_R2278_U162 = new_P1_R2278_U369 & new_P1_R2278_U76;
  assign new_P1_R2278_U163 = new_P1_R2278_U73 & new_P1_R2278_U80;
  assign new_P1_R2278_U164 = new_P1_R2278_U317 & new_P1_R2278_U10;
  assign new_P1_R2278_U165 = new_P1_R2278_U371 & new_P1_R2278_U316;
  assign new_P1_R2278_U166 = new_P1_R2278_U311 & new_P1_R2278_U313;
  assign new_P1_R2278_U167 = new_P1_R2278_U370 & new_P1_R2278_U314;
  assign new_P1_R2278_U168 = new_P1_R2278_U286 & new_P1_R2278_U415;
  assign new_P1_R2278_U169 = new_P1_R2278_U362 & new_P1_R2278_U79;
  assign new_P1_R2278_U170 = new_P1_R2278_U367 & new_P1_R2278_U306;
  assign new_P1_R2278_U171 = new_P1_R2278_U298 & new_P1_R2278_U302;
  assign new_P1_R2278_U172 = new_P1_R2278_U364 & new_P1_R2278_U303;
  assign new_P1_R2278_U173 = new_P1_R2278_U285 & new_P1_R2278_U589 & new_P1_R2278_U588;
  assign new_P1_R2278_U174 = new_P1_R2278_U337 & new_P1_R2278_U227;
  assign new_P1_R2278_U175 = new_P1_R2278_U228 & new_P1_R2278_U603 & new_P1_R2278_U602;
  assign new_P1_R2278_U176 = ~new_P1_R2278_U129 | ~new_P1_R2278_U353;
  assign new_P1_R2278_U177 = new_P1_R2278_U433 & new_P1_R2278_U432;
  assign new_P1_R2278_U178 = ~new_P1_R2278_U41 | ~new_P1_R2278_U256;
  assign new_P1_R2278_U179 = new_P1_R2278_U440 & new_P1_R2278_U439;
  assign new_P1_R2278_U180 = new_P1_R2278_U447 & new_P1_R2278_U446;
  assign new_P1_R2278_U181 = new_P1_R2278_U449 & new_P1_R2278_U448;
  assign new_P1_R2278_U182 = ~new_P1_R2278_U242 | ~new_P1_R2278_U241;
  assign new_P1_R2278_U183 = new_P1_R2278_U456 & new_P1_R2278_U455;
  assign new_P1_R2278_U184 = ~new_P1_R2278_U238 | ~new_P1_R2278_U237;
  assign new_P1_R2278_U185 = ~P1_INSTADDRPOINTER_REG_31_;
  assign new_P1_R2278_U186 = ~new_P1_U2769;
  assign new_P1_R2278_U187 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_U2771;
  assign new_P1_R2278_U188 = new_P1_R2278_U470 & new_P1_R2278_U469;
  assign new_P1_R2278_U189 = new_P1_R2278_U472 & new_P1_R2278_U471;
  assign new_P1_R2278_U190 = ~new_P1_R2278_U159 | ~new_P1_R2278_U407 | ~new_P1_R2278_U406 | ~new_P1_R2278_U405;
  assign new_P1_R2278_U191 = new_P1_R2278_U479 & new_P1_R2278_U478;
  assign new_P1_R2278_U192 = ~new_P1_R2278_U213 | ~new_P1_R2278_U234;
  assign new_P1_R2278_U193 = new_P1_R2278_U486 & new_P1_R2278_U485;
  assign new_P1_R2278_U194 = ~new_P1_R2278_U146 | ~new_P1_R2278_U145 | ~new_P1_R2278_U385;
  assign new_P1_R2278_U195 = new_P1_R2278_U493 & new_P1_R2278_U492;
  assign new_P1_R2278_U196 = ~new_P1_R2278_U419 | ~new_P1_R2278_U409;
  assign new_P1_R2278_U197 = new_P1_R2278_U500 & new_P1_R2278_U499;
  assign new_P1_R2278_U198 = ~new_P1_R2278_U425 | ~new_P1_R2278_U373;
  assign new_P1_R2278_U199 = new_P1_R2278_U507 & new_P1_R2278_U506;
  assign new_P1_R2278_U200 = ~new_P1_R2278_U165 | ~new_P1_R2278_U423;
  assign new_P1_R2278_U201 = new_P1_R2278_U514 & new_P1_R2278_U513;
  assign new_P1_R2278_U202 = ~new_P1_R2278_U167 | ~new_P1_R2278_U427;
  assign new_P1_R2278_U203 = new_P1_R2278_U521 & new_P1_R2278_U520;
  assign new_P1_R2278_U204 = ~new_P1_R2278_U421 | ~new_P1_R2278_U312;
  assign new_P1_R2278_U205 = new_P1_R2278_U528 & new_P1_R2278_U527;
  assign new_P1_R2278_U206 = ~new_P1_R2278_U162 | ~new_P1_R2278_U163 | ~new_P1_R2278_U376;
  assign new_P1_R2278_U207 = new_P1_R2278_U535 & new_P1_R2278_U534;
  assign new_P1_R2278_U208 = ~new_P1_R2278_U170 | ~new_P1_R2278_U365;
  assign new_P1_R2278_U209 = new_P1_R2278_U542 & new_P1_R2278_U541;
  assign new_P1_R2278_U210 = ~new_P1_R2278_U172 | ~new_P1_R2278_U363;
  assign new_P1_R2278_U211 = new_P1_R2278_U549 & new_P1_R2278_U548;
  assign new_P1_R2278_U212 = ~new_P1_R2278_U300 | ~new_P1_R2278_U299;
  assign new_P1_R2278_U213 = ~new_P1_U2799 | ~new_P1_R2278_U232;
  assign new_P1_R2278_U214 = new_P1_R2278_U559 & new_P1_R2278_U558;
  assign new_P1_R2278_U215 = new_P1_R2278_U561 & new_P1_R2278_U560;
  assign new_P1_R2278_U216 = ~new_P1_R2278_U169 | ~new_P1_R2278_U361;
  assign new_P1_R2278_U217 = new_P1_R2278_U568 & new_P1_R2278_U567;
  assign new_P1_R2278_U218 = ~new_P1_R2278_U360 | ~new_P1_R2278_U358;
  assign new_P1_R2278_U219 = new_P1_R2278_U575 & new_P1_R2278_U574;
  assign new_P1_R2278_U220 = ~new_P1_R2278_U290 | ~new_P1_R2278_U289;
  assign new_P1_R2278_U221 = new_P1_R2278_U582 & new_P1_R2278_U581;
  assign new_P1_R2278_U222 = ~new_P1_R2278_U168 | ~new_P1_R2278_U226;
  assign new_P1_R2278_U223 = ~new_P1_R2278_U68 | ~new_P1_R2278_U328;
  assign new_P1_R2278_U224 = ~new_P1_R2278_U98 | ~new_P1_R2278_U279;
  assign new_P1_R2278_U225 = ~new_P1_R2278_U274 | ~new_P1_R2278_U273;
  assign new_P1_R2278_U226 = ~new_P1_R2278_U224 | ~new_P1_R2278_U139;
  assign new_P1_R2278_U227 = ~new_P1_R2278_U356 | ~new_P1_R2278_U355;
  assign new_P1_R2278_U228 = ~new_P1_U2790 | ~P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_R2278_U229 = ~new_P1_U2787 | ~P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_R2278_U230 = ~new_P1_R2278_U213;
  assign new_P1_R2278_U231 = ~new_P1_U2794 | ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_R2278_U232 = ~new_P1_R2278_U32;
  assign new_P1_R2278_U233 = ~new_P1_R2278_U33 | ~new_P1_R2278_U32;
  assign new_P1_R2278_U234 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_R2278_U233;
  assign new_P1_R2278_U235 = ~new_P1_R2278_U192;
  assign new_P1_R2278_U236 = P1_INSTADDRPOINTER_REG_2_ | new_P1_U2798;
  assign new_P1_R2278_U237 = ~new_P1_R2278_U236 | ~new_P1_R2278_U192;
  assign new_P1_R2278_U238 = ~new_P1_U2798 | ~P1_INSTADDRPOINTER_REG_2_;
  assign new_P1_R2278_U239 = ~new_P1_R2278_U184;
  assign new_P1_R2278_U240 = P1_INSTADDRPOINTER_REG_3_ | new_P1_U2797;
  assign new_P1_R2278_U241 = ~new_P1_R2278_U240 | ~new_P1_R2278_U184;
  assign new_P1_R2278_U242 = ~new_P1_U2797 | ~P1_INSTADDRPOINTER_REG_3_;
  assign new_P1_R2278_U243 = ~new_P1_R2278_U182;
  assign new_P1_R2278_U244 = P1_INSTADDRPOINTER_REG_4_ | new_P1_U2796;
  assign new_P1_R2278_U245 = ~new_P1_R2278_U244 | ~new_P1_R2278_U182;
  assign new_P1_R2278_U246 = ~new_P1_U2796 | ~P1_INSTADDRPOINTER_REG_4_;
  assign new_P1_R2278_U247 = ~new_P1_R2278_U42;
  assign new_P1_R2278_U248 = new_P1_U2795 | P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_R2278_U249 = ~new_P1_R2278_U43;
  assign new_P1_R2278_U250 = ~new_P1_U2795 | ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_R2278_U251 = ~new_P1_R2278_U40;
  assign new_P1_R2278_U252 = ~new_P1_R2278_U251 | ~new_P1_R2278_U231;
  assign new_P1_R2278_U253 = new_P1_U2793 | P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_R2278_U254 = new_P1_U2794 | P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_R2278_U255 = ~new_P1_R2278_U41;
  assign new_P1_R2278_U256 = ~new_P1_U2793 | ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_R2278_U257 = ~new_P1_R2278_U178;
  assign new_P1_R2278_U258 = P1_INSTADDRPOINTER_REG_8_ | new_P1_U2792;
  assign new_P1_R2278_U259 = ~new_P1_U2792 | ~P1_INSTADDRPOINTER_REG_8_;
  assign new_P1_R2278_U260 = ~new_P1_R2278_U176;
  assign new_P1_R2278_U261 = P1_INSTADDRPOINTER_REG_9_ | new_P1_U2791;
  assign new_P1_R2278_U262 = ~new_P1_U2791 | ~P1_INSTADDRPOINTER_REG_9_;
  assign new_P1_R2278_U263 = ~new_P1_U2791 | ~P1_INSTADDRPOINTER_REG_9_;
  assign new_P1_R2278_U264 = P1_INSTADDRPOINTER_REG_6_ | new_P1_U2794;
  assign new_P1_R2278_U265 = ~new_P1_R2278_U264 | ~new_P1_R2278_U40;
  assign new_P1_R2278_U266 = ~new_P1_R2278_U179 | ~new_P1_R2278_U265 | ~new_P1_R2278_U231;
  assign new_P1_R2278_U267 = ~new_P1_U2793 | ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_R2278_U268 = ~new_P1_R2278_U255 | ~new_P1_R2278_U267;
  assign new_P1_R2278_U269 = new_P1_U2794 | P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_R2278_U270 = ~new_P1_R2278_U180 | ~new_P1_R2278_U247;
  assign new_P1_R2278_U271 = ~new_P1_U2795 | ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_R2278_U272 = ~new_P1_R2278_U249 | ~new_P1_R2278_U271;
  assign new_P1_R2278_U273 = ~new_P1_U2791 | ~P1_INSTADDRPOINTER_REG_9_;
  assign new_P1_R2278_U274 = ~new_P1_R2278_U261 | ~new_P1_R2278_U176;
  assign new_P1_R2278_U275 = ~new_P1_R2278_U225;
  assign new_P1_R2278_U276 = new_P1_U2789 | P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_R2278_U277 = new_P1_U2790 | P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_R2278_U278 = ~new_P1_R2278_U98;
  assign new_P1_R2278_U279 = ~new_P1_U2789 | ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_R2278_U280 = ~new_P1_R2278_U224;
  assign new_P1_R2278_U281 = P1_INSTADDRPOINTER_REG_12_ | new_P1_U2788;
  assign new_P1_R2278_U282 = ~new_P1_R2278_U68;
  assign new_P1_R2278_U283 = new_P1_U2787 | P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_R2278_U284 = new_P1_U2786 | P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_R2278_U285 = ~new_P1_U2786 | ~P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_R2278_U286 = ~new_P1_U2785 | ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_R2278_U287 = ~new_P1_R2278_U285 | ~new_P1_R2278_U391 | ~new_P1_R2278_U229;
  assign new_P1_R2278_U288 = P1_INSTADDRPOINTER_REG_16_ | new_P1_U2784;
  assign new_P1_R2278_U289 = ~new_P1_R2278_U288 | ~new_P1_R2278_U222;
  assign new_P1_R2278_U290 = ~new_P1_U2784 | ~P1_INSTADDRPOINTER_REG_16_;
  assign new_P1_R2278_U291 = ~new_P1_R2278_U220;
  assign new_P1_R2278_U292 = P1_INSTADDRPOINTER_REG_17_ | new_P1_U2783;
  assign new_P1_R2278_U293 = ~new_P1_U2783 | ~P1_INSTADDRPOINTER_REG_17_;
  assign new_P1_R2278_U294 = ~new_P1_R2278_U218;
  assign new_P1_R2278_U295 = P1_INSTADDRPOINTER_REG_18_ | new_P1_U2782;
  assign new_P1_R2278_U296 = ~new_P1_R2278_U79;
  assign new_P1_R2278_U297 = ~new_P1_R2278_U216;
  assign new_P1_R2278_U298 = P1_INSTADDRPOINTER_REG_19_ | new_P1_U2781;
  assign new_P1_R2278_U299 = ~new_P1_R2278_U298 | ~new_P1_R2278_U216;
  assign new_P1_R2278_U300 = ~new_P1_U2781 | ~P1_INSTADDRPOINTER_REG_19_;
  assign new_P1_R2278_U301 = ~new_P1_R2278_U212;
  assign new_P1_R2278_U302 = P1_INSTADDRPOINTER_REG_20_ | new_P1_U2780;
  assign new_P1_R2278_U303 = ~new_P1_U2780 | ~P1_INSTADDRPOINTER_REG_20_;
  assign new_P1_R2278_U304 = ~new_P1_R2278_U210;
  assign new_P1_R2278_U305 = P1_INSTADDRPOINTER_REG_21_ | new_P1_U2779;
  assign new_P1_R2278_U306 = ~new_P1_U2779 | ~P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_R2278_U307 = ~new_P1_R2278_U208;
  assign new_P1_R2278_U308 = P1_INSTADDRPOINTER_REG_22_ | new_P1_U2778;
  assign new_P1_R2278_U309 = ~new_P1_R2278_U76;
  assign new_P1_R2278_U310 = ~new_P1_R2278_U206;
  assign new_P1_R2278_U311 = P1_INSTADDRPOINTER_REG_23_ | new_P1_U2777;
  assign new_P1_R2278_U312 = ~new_P1_U2777 | ~P1_INSTADDRPOINTER_REG_23_;
  assign new_P1_R2278_U313 = P1_INSTADDRPOINTER_REG_24_ | new_P1_U2776;
  assign new_P1_R2278_U314 = ~new_P1_U2776 | ~P1_INSTADDRPOINTER_REG_24_;
  assign new_P1_R2278_U315 = P1_INSTADDRPOINTER_REG_25_ | new_P1_U2775;
  assign new_P1_R2278_U316 = ~new_P1_U2775 | ~P1_INSTADDRPOINTER_REG_25_;
  assign new_P1_R2278_U317 = P1_INSTADDRPOINTER_REG_26_ | new_P1_U2774;
  assign new_P1_R2278_U318 = ~new_P1_U2774 | ~P1_INSTADDRPOINTER_REG_26_;
  assign new_P1_R2278_U319 = P1_INSTADDRPOINTER_REG_27_ | new_P1_U2773;
  assign new_P1_R2278_U320 = ~new_P1_R2278_U85;
  assign new_P1_R2278_U321 = new_P1_U2772 | P1_INSTADDRPOINTER_REG_28_;
  assign new_P1_R2278_U322 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_U2772;
  assign new_P1_R2278_U323 = ~new_P1_R2278_U194;
  assign new_P1_R2278_U324 = new_P1_U2771 | P1_INSTADDRPOINTER_REG_29_;
  assign new_P1_R2278_U325 = ~new_P1_R2278_U187;
  assign new_P1_R2278_U326 = ~new_P1_R2278_U190;
  assign new_P1_R2278_U327 = P1_INSTADDRPOINTER_REG_30_ | new_P1_U2770;
  assign new_P1_R2278_U328 = ~new_P1_R2278_U281 | ~new_P1_R2278_U224;
  assign new_P1_R2278_U329 = ~new_P1_R2278_U223;
  assign new_P1_R2278_U330 = P1_INSTADDRPOINTER_REG_13_ | new_P1_U2787;
  assign new_P1_R2278_U331 = ~new_P1_R2278_U330 | ~new_P1_R2278_U223;
  assign new_P1_R2278_U332 = ~new_P1_R2278_U97;
  assign new_P1_R2278_U333 = P1_INSTADDRPOINTER_REG_14_ | new_P1_U2786;
  assign new_P1_R2278_U334 = ~new_P1_R2278_U333 | ~new_P1_R2278_U97;
  assign new_P1_R2278_U335 = ~new_P1_R2278_U173 | ~new_P1_R2278_U334;
  assign new_P1_R2278_U336 = ~new_P1_R2278_U332 | ~new_P1_R2278_U285;
  assign new_P1_R2278_U337 = ~new_P1_U2785 | ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_R2278_U338 = new_P1_U2786 | P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_R2278_U339 = new_P1_U2787 | P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_R2278_U340 = P1_INSTADDRPOINTER_REG_10_ | new_P1_U2790;
  assign new_P1_R2278_U341 = ~new_P1_R2278_U340 | ~new_P1_R2278_U225;
  assign new_P1_R2278_U342 = ~new_P1_R2278_U175 | ~new_P1_R2278_U341;
  assign new_P1_R2278_U343 = ~new_P1_U2789 | ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_R2278_U344 = ~new_P1_R2278_U278 | ~new_P1_R2278_U343;
  assign new_P1_R2278_U345 = new_P1_U2790 | P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_R2278_U346 = ~new_P1_R2278_U263 | ~new_P1_R2278_U261;
  assign new_P1_R2278_U347 = ~new_P1_R2278_U269 | ~new_P1_R2278_U231;
  assign new_P1_R2278_U348 = ~new_P1_R2278_U338 | ~new_P1_R2278_U285;
  assign new_P1_R2278_U349 = ~new_P1_R2278_U339 | ~new_P1_R2278_U229;
  assign new_P1_R2278_U350 = ~new_P1_R2278_U68 | ~new_P1_R2278_U281;
  assign new_P1_R2278_U351 = ~new_P1_R2278_U345 | ~new_P1_R2278_U228;
  assign new_P1_R2278_U352 = ~new_P1_R2278_U127 | ~new_P1_R2278_U258;
  assign new_P1_R2278_U353 = ~new_P1_R2278_U128 | ~new_P1_R2278_U253 | ~new_P1_R2278_U252;
  assign new_P1_R2278_U354 = ~new_P1_R2278_U137 | ~new_P1_R2278_U353 | ~new_P1_R2278_U352;
  assign new_P1_R2278_U355 = ~new_P1_U2785 | ~new_P1_R2278_U284;
  assign new_P1_R2278_U356 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_R2278_U284;
  assign new_P1_R2278_U357 = ~new_P1_R2278_U356 | ~new_P1_R2278_U63;
  assign new_P1_R2278_U358 = ~new_P1_R2278_U6 | ~new_P1_R2278_U222;
  assign new_P1_R2278_U359 = ~new_P1_R2278_U293 | ~new_P1_R2278_U290;
  assign new_P1_R2278_U360 = ~new_P1_R2278_U359 | ~new_P1_R2278_U292;
  assign new_P1_R2278_U361 = ~new_P1_R2278_U7 | ~new_P1_R2278_U222;
  assign new_P1_R2278_U362 = ~new_P1_R2278_U12 | ~new_P1_R2278_U359;
  assign new_P1_R2278_U363 = ~new_P1_R2278_U171 | ~new_P1_R2278_U216;
  assign new_P1_R2278_U364 = ~new_P1_R2278_U133 | ~new_P1_R2278_U302;
  assign new_P1_R2278_U365 = ~new_P1_R2278_U8 | ~new_P1_R2278_U216;
  assign new_P1_R2278_U366 = ~new_P1_R2278_U364 | ~new_P1_R2278_U303;
  assign new_P1_R2278_U367 = ~new_P1_R2278_U366 | ~new_P1_R2278_U305;
  assign new_P1_R2278_U368 = ~new_P1_R2278_U367 | ~new_P1_R2278_U306;
  assign new_P1_R2278_U369 = ~new_P1_R2278_U368 | ~new_P1_R2278_U308;
  assign new_P1_R2278_U370 = ~new_P1_R2278_U130 | ~new_P1_R2278_U313;
  assign new_P1_R2278_U371 = ~new_P1_R2278_U381 | ~new_P1_R2278_U315;
  assign new_P1_R2278_U372 = ~new_P1_R2278_U131 | ~new_P1_R2278_U371;
  assign new_P1_R2278_U373 = ~new_P1_R2278_U372 | ~new_P1_R2278_U317;
  assign new_P1_R2278_U374 = ~new_P1_R2278_U372 | ~new_P1_R2278_U317;
  assign new_P1_R2278_U375 = ~new_P1_R2278_U147 | ~new_P1_R2278_U194;
  assign new_P1_R2278_U376 = ~new_P1_R2278_U161 | ~new_P1_R2278_U418;
  assign new_P1_R2278_U377 = ~new_P1_R2278_U80;
  assign new_P1_R2278_U378 = ~new_P1_R2278_U73;
  assign new_P1_R2278_U379 = ~new_P1_R2278_U320 | ~new_P1_R2278_U321;
  assign new_P1_R2278_U380 = ~new_P1_R2278_U94;
  assign new_P1_R2278_U381 = ~new_P1_R2278_U370 | ~new_P1_R2278_U314;
  assign new_P1_R2278_U382 = ~new_P1_R2278_U285 | ~new_P1_R2278_U391 | ~new_P1_R2278_U229;
  assign new_P1_R2278_U383 = ~new_P1_R2278_U92;
  assign new_P1_R2278_U384 = ~new_P1_R2278_U95;
  assign new_P1_R2278_U385 = ~new_P1_R2278_U142 | ~new_P1_R2278_U11 | ~new_P1_R2278_U411;
  assign new_P1_R2278_U386 = ~new_P1_R2278_U93;
  assign new_P1_R2278_U387 = ~new_P1_R2278_U96;
  assign new_P1_R2278_U388 = ~new_P1_R2278_U277 | ~new_P1_R2278_U261;
  assign new_P1_R2278_U389 = ~new_P1_R2278_U388 | ~new_P1_R2278_U228;
  assign new_P1_R2278_U390 = ~new_P1_R2278_U285 | ~new_P1_R2278_U391 | ~new_P1_R2278_U229;
  assign new_P1_R2278_U391 = ~new_P1_R2278_U282 | ~new_P1_R2278_U283;
  assign new_P1_R2278_U392 = ~new_P1_R2278_U86;
  assign new_P1_R2278_U393 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_U2770;
  assign new_P1_R2278_U394 = ~new_P1_R2278_U148 | ~new_P1_R2278_U372;
  assign new_P1_R2278_U395 = ~new_P1_R2278_U383 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U396 = ~new_P1_R2278_U150 | ~new_P1_R2278_U368;
  assign new_P1_R2278_U397 = ~new_P1_R2278_U153 | ~new_P1_R2278_U152 | ~new_P1_R2278_U413;
  assign new_P1_R2278_U398 = ~new_P1_R2278_U386 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U399 = ~new_P1_R2278_U378 | ~new_P1_R2278_U154 | ~new_P1_R2278_U11;
  assign new_P1_R2278_U400 = ~new_P1_R2278_U86 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U401 = ~new_P1_R2278_U87;
  assign new_P1_R2278_U402 = ~new_P1_R2278_U285 | ~new_P1_R2278_U391 | ~new_P1_R2278_U229;
  assign new_P1_R2278_U403 = ~new_P1_R2278_U380 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U404 = ~new_P1_R2278_U384 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U405 = ~new_P1_R2278_U158 | ~new_P1_R2278_U157 | ~new_P1_R2278_U411;
  assign new_P1_R2278_U406 = ~new_P1_R2278_U387 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U407 = ~new_P1_R2278_U87 | ~new_P1_R2278_U324;
  assign new_P1_R2278_U408 = ~new_P1_R2278_U374 | ~new_P1_R2278_U85;
  assign new_P1_R2278_U409 = ~new_P1_R2278_U408 | ~new_P1_R2278_U319;
  assign new_P1_R2278_U410 = ~new_P1_R2278_U402 | ~new_P1_R2278_U227;
  assign new_P1_R2278_U411 = ~new_P1_R2278_U141 | ~new_P1_R2278_U226;
  assign new_P1_R2278_U412 = ~new_P1_R2278_U390 | ~new_P1_R2278_U227;
  assign new_P1_R2278_U413 = ~new_P1_R2278_U151 | ~new_P1_R2278_U226;
  assign new_P1_R2278_U414 = ~new_P1_R2278_U174 | ~new_P1_R2278_U336;
  assign new_P1_R2278_U415 = ~new_P1_R2278_U287 | ~new_P1_R2278_U227;
  assign new_P1_R2278_U416 = ~new_P1_R2278_U222;
  assign new_P1_R2278_U417 = ~new_P1_R2278_U382 | ~new_P1_R2278_U227;
  assign new_P1_R2278_U418 = ~new_P1_R2278_U160 | ~new_P1_R2278_U226;
  assign new_P1_R2278_U419 = ~new_P1_R2278_U11 | ~new_P1_R2278_U206;
  assign new_P1_R2278_U420 = ~new_P1_R2278_U196;
  assign new_P1_R2278_U421 = ~new_P1_R2278_U311 | ~new_P1_R2278_U206;
  assign new_P1_R2278_U422 = ~new_P1_R2278_U204;
  assign new_P1_R2278_U423 = ~new_P1_R2278_U10 | ~new_P1_R2278_U206;
  assign new_P1_R2278_U424 = ~new_P1_R2278_U200;
  assign new_P1_R2278_U425 = ~new_P1_R2278_U164 | ~new_P1_R2278_U206;
  assign new_P1_R2278_U426 = ~new_P1_R2278_U198;
  assign new_P1_R2278_U427 = ~new_P1_R2278_U166 | ~new_P1_R2278_U206;
  assign new_P1_R2278_U428 = ~new_P1_R2278_U202;
  assign new_P1_R2278_U429 = ~new_P1_R2278_U557 | ~new_P1_R2278_U33;
  assign new_P1_R2278_U430 = ~new_P1_R2278_U346 | ~new_P1_R2278_U176;
  assign new_P1_R2278_U431 = ~new_P1_R2278_U100 | ~new_P1_R2278_U260;
  assign new_P1_R2278_U432 = ~new_P1_U2792 | ~new_P1_R2278_U21;
  assign new_P1_R2278_U433 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_R2278_U22;
  assign new_P1_R2278_U434 = ~new_P1_U2792 | ~new_P1_R2278_U21;
  assign new_P1_R2278_U435 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_R2278_U22;
  assign new_P1_R2278_U436 = ~new_P1_R2278_U435 | ~new_P1_R2278_U434;
  assign new_P1_R2278_U437 = ~new_P1_R2278_U177 | ~new_P1_R2278_U178;
  assign new_P1_R2278_U438 = ~new_P1_R2278_U257 | ~new_P1_R2278_U436;
  assign new_P1_R2278_U439 = ~new_P1_U2793 | ~new_P1_R2278_U23;
  assign new_P1_R2278_U440 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_R2278_U24;
  assign new_P1_R2278_U441 = ~new_P1_U2794 | ~new_P1_R2278_U25;
  assign new_P1_R2278_U442 = ~P1_INSTADDRPOINTER_REG_6_ | ~new_P1_R2278_U26;
  assign new_P1_R2278_U443 = ~new_P1_R2278_U442 | ~new_P1_R2278_U441;
  assign new_P1_R2278_U444 = ~new_P1_R2278_U347 | ~new_P1_R2278_U40;
  assign new_P1_R2278_U445 = ~new_P1_R2278_U443 | ~new_P1_R2278_U251;
  assign new_P1_R2278_U446 = ~new_P1_U2795 | ~new_P1_R2278_U27;
  assign new_P1_R2278_U447 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_R2278_U28;
  assign new_P1_R2278_U448 = ~new_P1_U2796 | ~new_P1_R2278_U38;
  assign new_P1_R2278_U449 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_R2278_U39;
  assign new_P1_R2278_U450 = ~new_P1_U2796 | ~new_P1_R2278_U38;
  assign new_P1_R2278_U451 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_R2278_U39;
  assign new_P1_R2278_U452 = ~new_P1_R2278_U451 | ~new_P1_R2278_U450;
  assign new_P1_R2278_U453 = ~new_P1_R2278_U181 | ~new_P1_R2278_U182;
  assign new_P1_R2278_U454 = ~new_P1_R2278_U243 | ~new_P1_R2278_U452;
  assign new_P1_R2278_U455 = ~new_P1_U2797 | ~new_P1_R2278_U36;
  assign new_P1_R2278_U456 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_R2278_U37;
  assign new_P1_R2278_U457 = ~new_P1_U2797 | ~new_P1_R2278_U36;
  assign new_P1_R2278_U458 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_R2278_U37;
  assign new_P1_R2278_U459 = ~new_P1_R2278_U458 | ~new_P1_R2278_U457;
  assign new_P1_R2278_U460 = ~new_P1_R2278_U183 | ~new_P1_R2278_U184;
  assign new_P1_R2278_U461 = ~new_P1_R2278_U239 | ~new_P1_R2278_U459;
  assign new_P1_R2278_U462 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_R2278_U186;
  assign new_P1_R2278_U463 = ~new_P1_U2769 | ~new_P1_R2278_U185;
  assign new_P1_R2278_U464 = ~P1_INSTADDRPOINTER_REG_31_ | ~new_P1_R2278_U186;
  assign new_P1_R2278_U465 = ~new_P1_U2769 | ~new_P1_R2278_U185;
  assign new_P1_R2278_U466 = ~new_P1_R2278_U465 | ~new_P1_R2278_U464;
  assign new_P1_R2278_U467 = ~new_P1_R2278_U187 | ~new_P1_R2278_U155 | ~new_P1_R2278_U397 | ~new_P1_R2278_U396;
  assign new_P1_R2278_U468 = ~new_P1_R2278_U325 | ~new_P1_R2278_U5;
  assign new_P1_R2278_U469 = ~new_P1_R2278_U89 | ~new_P1_R2278_U14 | ~new_P1_R2278_U88;
  assign new_P1_R2278_U470 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_U2770 | ~new_P1_R2278_U466;
  assign new_P1_R2278_U471 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_R2278_U88;
  assign new_P1_R2278_U472 = ~new_P1_U2770 | ~new_P1_R2278_U89;
  assign new_P1_R2278_U473 = ~P1_INSTADDRPOINTER_REG_30_ | ~new_P1_R2278_U88;
  assign new_P1_R2278_U474 = ~new_P1_U2770 | ~new_P1_R2278_U89;
  assign new_P1_R2278_U475 = ~new_P1_R2278_U474 | ~new_P1_R2278_U473;
  assign new_P1_R2278_U476 = ~new_P1_R2278_U189 | ~new_P1_R2278_U190;
  assign new_P1_R2278_U477 = ~new_P1_R2278_U326 | ~new_P1_R2278_U475;
  assign new_P1_R2278_U478 = ~new_P1_U2798 | ~new_P1_R2278_U34;
  assign new_P1_R2278_U479 = ~P1_INSTADDRPOINTER_REG_2_ | ~new_P1_R2278_U35;
  assign new_P1_R2278_U480 = ~new_P1_U2798 | ~new_P1_R2278_U34;
  assign new_P1_R2278_U481 = ~P1_INSTADDRPOINTER_REG_2_ | ~new_P1_R2278_U35;
  assign new_P1_R2278_U482 = ~new_P1_R2278_U481 | ~new_P1_R2278_U480;
  assign new_P1_R2278_U483 = ~new_P1_R2278_U191 | ~new_P1_R2278_U192;
  assign new_P1_R2278_U484 = ~new_P1_R2278_U235 | ~new_P1_R2278_U482;
  assign new_P1_R2278_U485 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_R2278_U90;
  assign new_P1_R2278_U486 = ~new_P1_U2771 | ~new_P1_R2278_U91;
  assign new_P1_R2278_U487 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_R2278_U90;
  assign new_P1_R2278_U488 = ~new_P1_U2771 | ~new_P1_R2278_U91;
  assign new_P1_R2278_U489 = ~new_P1_R2278_U488 | ~new_P1_R2278_U487;
  assign new_P1_R2278_U490 = ~new_P1_R2278_U193 | ~new_P1_R2278_U194;
  assign new_P1_R2278_U491 = ~new_P1_R2278_U323 | ~new_P1_R2278_U489;
  assign new_P1_R2278_U492 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_R2278_U81;
  assign new_P1_R2278_U493 = ~new_P1_U2772 | ~new_P1_R2278_U82;
  assign new_P1_R2278_U494 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_R2278_U81;
  assign new_P1_R2278_U495 = ~new_P1_U2772 | ~new_P1_R2278_U82;
  assign new_P1_R2278_U496 = ~new_P1_R2278_U495 | ~new_P1_R2278_U494;
  assign new_P1_R2278_U497 = ~new_P1_R2278_U195 | ~new_P1_R2278_U196;
  assign new_P1_R2278_U498 = ~new_P1_R2278_U420 | ~new_P1_R2278_U496;
  assign new_P1_R2278_U499 = ~new_P1_U2773 | ~new_P1_R2278_U83;
  assign new_P1_R2278_U500 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_R2278_U84;
  assign new_P1_R2278_U501 = ~new_P1_U2773 | ~new_P1_R2278_U83;
  assign new_P1_R2278_U502 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_R2278_U84;
  assign new_P1_R2278_U503 = ~new_P1_R2278_U502 | ~new_P1_R2278_U501;
  assign new_P1_R2278_U504 = ~new_P1_R2278_U197 | ~new_P1_R2278_U198;
  assign new_P1_R2278_U505 = ~new_P1_R2278_U426 | ~new_P1_R2278_U503;
  assign new_P1_R2278_U506 = ~new_P1_U2774 | ~new_P1_R2278_U46;
  assign new_P1_R2278_U507 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_R2278_U47;
  assign new_P1_R2278_U508 = ~new_P1_U2774 | ~new_P1_R2278_U46;
  assign new_P1_R2278_U509 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_R2278_U47;
  assign new_P1_R2278_U510 = ~new_P1_R2278_U509 | ~new_P1_R2278_U508;
  assign new_P1_R2278_U511 = ~new_P1_R2278_U199 | ~new_P1_R2278_U200;
  assign new_P1_R2278_U512 = ~new_P1_R2278_U424 | ~new_P1_R2278_U510;
  assign new_P1_R2278_U513 = ~new_P1_U2775 | ~new_P1_R2278_U44;
  assign new_P1_R2278_U514 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_R2278_U45;
  assign new_P1_R2278_U515 = ~new_P1_U2775 | ~new_P1_R2278_U44;
  assign new_P1_R2278_U516 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_R2278_U45;
  assign new_P1_R2278_U517 = ~new_P1_R2278_U516 | ~new_P1_R2278_U515;
  assign new_P1_R2278_U518 = ~new_P1_R2278_U201 | ~new_P1_R2278_U202;
  assign new_P1_R2278_U519 = ~new_P1_R2278_U428 | ~new_P1_R2278_U517;
  assign new_P1_R2278_U520 = ~new_P1_U2776 | ~new_P1_R2278_U48;
  assign new_P1_R2278_U521 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_R2278_U49;
  assign new_P1_R2278_U522 = ~new_P1_U2776 | ~new_P1_R2278_U48;
  assign new_P1_R2278_U523 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_R2278_U49;
  assign new_P1_R2278_U524 = ~new_P1_R2278_U523 | ~new_P1_R2278_U522;
  assign new_P1_R2278_U525 = ~new_P1_R2278_U203 | ~new_P1_R2278_U204;
  assign new_P1_R2278_U526 = ~new_P1_R2278_U422 | ~new_P1_R2278_U524;
  assign new_P1_R2278_U527 = ~new_P1_U2777 | ~new_P1_R2278_U50;
  assign new_P1_R2278_U528 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_R2278_U51;
  assign new_P1_R2278_U529 = ~new_P1_U2777 | ~new_P1_R2278_U50;
  assign new_P1_R2278_U530 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_R2278_U51;
  assign new_P1_R2278_U531 = ~new_P1_R2278_U530 | ~new_P1_R2278_U529;
  assign new_P1_R2278_U532 = ~new_P1_R2278_U205 | ~new_P1_R2278_U206;
  assign new_P1_R2278_U533 = ~new_P1_R2278_U310 | ~new_P1_R2278_U531;
  assign new_P1_R2278_U534 = ~new_P1_U2778 | ~new_P1_R2278_U74;
  assign new_P1_R2278_U535 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_R2278_U75;
  assign new_P1_R2278_U536 = ~new_P1_U2778 | ~new_P1_R2278_U74;
  assign new_P1_R2278_U537 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_R2278_U75;
  assign new_P1_R2278_U538 = ~new_P1_R2278_U537 | ~new_P1_R2278_U536;
  assign new_P1_R2278_U539 = ~new_P1_R2278_U207 | ~new_P1_R2278_U208;
  assign new_P1_R2278_U540 = ~new_P1_R2278_U307 | ~new_P1_R2278_U538;
  assign new_P1_R2278_U541 = ~new_P1_U2779 | ~new_P1_R2278_U52;
  assign new_P1_R2278_U542 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_R2278_U53;
  assign new_P1_R2278_U543 = ~new_P1_U2779 | ~new_P1_R2278_U52;
  assign new_P1_R2278_U544 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_R2278_U53;
  assign new_P1_R2278_U545 = ~new_P1_R2278_U544 | ~new_P1_R2278_U543;
  assign new_P1_R2278_U546 = ~new_P1_R2278_U209 | ~new_P1_R2278_U210;
  assign new_P1_R2278_U547 = ~new_P1_R2278_U304 | ~new_P1_R2278_U545;
  assign new_P1_R2278_U548 = ~new_P1_U2780 | ~new_P1_R2278_U54;
  assign new_P1_R2278_U549 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_R2278_U55;
  assign new_P1_R2278_U550 = ~new_P1_U2780 | ~new_P1_R2278_U54;
  assign new_P1_R2278_U551 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_R2278_U55;
  assign new_P1_R2278_U552 = ~new_P1_R2278_U551 | ~new_P1_R2278_U550;
  assign new_P1_R2278_U553 = ~new_P1_R2278_U211 | ~new_P1_R2278_U212;
  assign new_P1_R2278_U554 = ~new_P1_R2278_U301 | ~new_P1_R2278_U552;
  assign new_P1_R2278_U555 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_R2278_U32;
  assign new_P1_R2278_U556 = ~new_P1_R2278_U232 | ~new_P1_R2278_U31;
  assign new_P1_R2278_U557 = ~new_P1_R2278_U556 | ~new_P1_R2278_U555;
  assign new_P1_R2278_U558 = ~new_P1_R2278_U31 | ~new_P1_U2799 | ~new_P1_R2278_U32;
  assign new_P1_R2278_U559 = ~new_P1_R2278_U230 | ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_R2278_U560 = ~new_P1_U2781 | ~new_P1_R2278_U56;
  assign new_P1_R2278_U561 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_R2278_U57;
  assign new_P1_R2278_U562 = ~new_P1_U2781 | ~new_P1_R2278_U56;
  assign new_P1_R2278_U563 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_R2278_U57;
  assign new_P1_R2278_U564 = ~new_P1_R2278_U563 | ~new_P1_R2278_U562;
  assign new_P1_R2278_U565 = ~new_P1_R2278_U215 | ~new_P1_R2278_U216;
  assign new_P1_R2278_U566 = ~new_P1_R2278_U297 | ~new_P1_R2278_U564;
  assign new_P1_R2278_U567 = ~new_P1_U2782 | ~new_P1_R2278_U77;
  assign new_P1_R2278_U568 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_R2278_U78;
  assign new_P1_R2278_U569 = ~new_P1_U2782 | ~new_P1_R2278_U77;
  assign new_P1_R2278_U570 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_R2278_U78;
  assign new_P1_R2278_U571 = ~new_P1_R2278_U570 | ~new_P1_R2278_U569;
  assign new_P1_R2278_U572 = ~new_P1_R2278_U217 | ~new_P1_R2278_U218;
  assign new_P1_R2278_U573 = ~new_P1_R2278_U294 | ~new_P1_R2278_U571;
  assign new_P1_R2278_U574 = ~new_P1_U2783 | ~new_P1_R2278_U71;
  assign new_P1_R2278_U575 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_R2278_U72;
  assign new_P1_R2278_U576 = ~new_P1_U2783 | ~new_P1_R2278_U71;
  assign new_P1_R2278_U577 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_R2278_U72;
  assign new_P1_R2278_U578 = ~new_P1_R2278_U577 | ~new_P1_R2278_U576;
  assign new_P1_R2278_U579 = ~new_P1_R2278_U219 | ~new_P1_R2278_U220;
  assign new_P1_R2278_U580 = ~new_P1_R2278_U291 | ~new_P1_R2278_U578;
  assign new_P1_R2278_U581 = ~new_P1_U2784 | ~new_P1_R2278_U69;
  assign new_P1_R2278_U582 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_R2278_U70;
  assign new_P1_R2278_U583 = ~new_P1_U2784 | ~new_P1_R2278_U69;
  assign new_P1_R2278_U584 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_R2278_U70;
  assign new_P1_R2278_U585 = ~new_P1_R2278_U584 | ~new_P1_R2278_U583;
  assign new_P1_R2278_U586 = ~new_P1_R2278_U221 | ~new_P1_R2278_U222;
  assign new_P1_R2278_U587 = ~new_P1_R2278_U416 | ~new_P1_R2278_U585;
  assign new_P1_R2278_U588 = ~new_P1_U2785 | ~new_P1_R2278_U62;
  assign new_P1_R2278_U589 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_R2278_U63;
  assign new_P1_R2278_U590 = ~new_P1_U2786 | ~new_P1_R2278_U66;
  assign new_P1_R2278_U591 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_R2278_U67;
  assign new_P1_R2278_U592 = ~new_P1_R2278_U591 | ~new_P1_R2278_U590;
  assign new_P1_R2278_U593 = ~new_P1_R2278_U348 | ~new_P1_R2278_U97;
  assign new_P1_R2278_U594 = ~new_P1_R2278_U592 | ~new_P1_R2278_U332;
  assign new_P1_R2278_U595 = ~new_P1_U2787 | ~new_P1_R2278_U64;
  assign new_P1_R2278_U596 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_R2278_U65;
  assign new_P1_R2278_U597 = ~new_P1_R2278_U596 | ~new_P1_R2278_U595;
  assign new_P1_R2278_U598 = ~new_P1_R2278_U349 | ~new_P1_R2278_U223;
  assign new_P1_R2278_U599 = ~new_P1_R2278_U329 | ~new_P1_R2278_U597;
  assign new_P1_R2278_U600 = ~new_P1_R2278_U350 | ~new_P1_R2278_U224;
  assign new_P1_R2278_U601 = ~new_P1_R2278_U124 | ~new_P1_R2278_U280;
  assign new_P1_R2278_U602 = ~new_P1_U2789 | ~new_P1_R2278_U58;
  assign new_P1_R2278_U603 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_R2278_U59;
  assign new_P1_R2278_U604 = ~new_P1_U2790 | ~new_P1_R2278_U60;
  assign new_P1_R2278_U605 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_R2278_U61;
  assign new_P1_R2278_U606 = ~new_P1_R2278_U605 | ~new_P1_R2278_U604;
  assign new_P1_R2278_U607 = ~new_P1_R2278_U351 | ~new_P1_R2278_U225;
  assign new_P1_R2278_U608 = ~new_P1_R2278_U275 | ~new_P1_R2278_U606;
  assign new_P1_R2278_U609 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_R2278_U29;
  assign new_P1_R2278_U610 = ~new_P1_U2800 | ~new_P1_R2278_U30;
  assign new_P1_R2358_U5 = new_P1_R2358_U274 & new_P1_R2358_U272;
  assign new_P1_R2358_U6 = new_P1_R2358_U280 & new_P1_R2358_U278;
  assign new_P1_R2358_U7 = new_P1_R2358_U6 & new_P1_R2358_U282;
  assign new_P1_R2358_U8 = new_P1_R2358_U288 & new_P1_R2358_U286;
  assign new_P1_R2358_U9 = new_P1_R2358_U8 & new_P1_R2358_U290;
  assign new_P1_R2358_U10 = new_P1_R2358_U9 & new_P1_R2358_U292;
  assign new_P1_R2358_U11 = new_P1_R2358_U458 & new_P1_R2358_U457;
  assign new_P1_R2358_U12 = new_P1_R2358_U481 & new_P1_R2358_U480;
  assign new_P1_R2358_U13 = new_P1_R2358_U555 & new_P1_R2358_U554;
  assign new_P1_R2358_U14 = new_P1_R2358_U330 & new_P1_R2358_U329;
  assign new_P1_R2358_U15 = new_P1_R2358_U327 & new_P1_R2358_U325;
  assign new_P1_R2358_U16 = new_P1_R2358_U320 & new_P1_R2358_U319;
  assign new_P1_R2358_U17 = new_P1_R2358_U317 & new_P1_R2358_U315;
  assign new_P1_R2358_U18 = new_P1_R2358_U308 & new_P1_R2358_U307;
  assign new_P1_R2358_U19 = new_P1_R2358_U254 & new_P1_R2358_U252;
  assign new_P1_R2358_U20 = new_P1_R2358_U245 & new_P1_R2358_U244;
  assign new_P1_R2358_U21 = new_P1_R2358_U242 & new_P1_R2358_U240;
  assign new_P1_R2358_U22 = new_P1_R2358_U136 & new_P1_R2358_U566 & new_P1_R2358_U565;
  assign new_P1_R2358_U23 = ~new_P1_U2352;
  assign new_P1_R2358_U24 = ~new_P1_U2643;
  assign new_P1_R2358_U25 = ~new_P1_U2644;
  assign new_P1_R2358_U26 = ~new_P1_U2645;
  assign new_P1_R2358_U27 = ~new_P1_U2646;
  assign new_P1_R2358_U28 = ~new_P1_U2646 | ~new_P1_R2358_U413;
  assign new_P1_R2358_U29 = ~new_P1_U2649;
  assign new_P1_R2358_U30 = ~new_P1_U2648;
  assign new_P1_R2358_U31 = ~new_P1_U2650;
  assign new_P1_R2358_U32 = ~new_P1_U2647;
  assign new_P1_R2358_U33 = ~new_P1_U2642;
  assign new_P1_R2358_U34 = ~new_P1_U2641;
  assign new_P1_R2358_U35 = ~new_P1_R2358_U236 | ~new_P1_R2358_U220;
  assign new_P1_R2358_U36 = ~new_P1_R2358_U35 | ~new_P1_R2358_U218;
  assign new_P1_R2358_U37 = ~new_P1_U2623;
  assign new_P1_R2358_U38 = ~new_P1_U2624;
  assign new_P1_R2358_U39 = ~new_P1_U2625;
  assign new_P1_R2358_U40 = ~new_P1_U2626;
  assign new_P1_R2358_U41 = ~new_P1_U2627;
  assign new_P1_R2358_U42 = ~new_P1_U2627 | ~new_P1_R2358_U546;
  assign new_P1_R2358_U43 = ~new_P1_U2628;
  assign new_P1_R2358_U44 = ~new_P1_U2629;
  assign new_P1_R2358_U45 = ~new_P1_U2630;
  assign new_P1_R2358_U46 = ~new_P1_U2631;
  assign new_P1_R2358_U47 = ~new_P1_U2631 | ~new_P1_R2358_U521;
  assign new_P1_R2358_U48 = ~new_P1_U2632;
  assign new_P1_R2358_U49 = ~new_P1_U2633;
  assign new_P1_R2358_U50 = ~new_P1_U2634;
  assign new_P1_R2358_U51 = ~new_P1_U2634 | ~new_P1_R2358_U501;
  assign new_P1_R2358_U52 = ~new_P1_U2639;
  assign new_P1_R2358_U53 = ~new_P1_U2640;
  assign new_P1_R2358_U54 = ~new_P1_R2358_U34 | ~new_P1_R2358_U400 | ~new_P1_R2358_U399;
  assign new_P1_R2358_U55 = ~new_P1_U2635;
  assign new_P1_R2358_U56 = ~new_P1_U2638;
  assign new_P1_R2358_U57 = ~new_P1_U2638 | ~new_P1_R2358_U471;
  assign new_P1_R2358_U58 = ~new_P1_U2637;
  assign new_P1_R2358_U59 = ~new_P1_U2637 | ~new_P1_R2358_U463;
  assign new_P1_R2358_U60 = ~new_P1_U2636;
  assign new_P1_R2358_U61 = ~new_P1_U2636 | ~new_P1_R2358_U466;
  assign new_P1_R2358_U62 = ~new_P1_U2622;
  assign new_P1_R2358_U63 = ~new_P1_U2620;
  assign new_P1_R2358_U64 = ~new_P1_U2621;
  assign new_P1_R2358_U65 = ~new_P1_R2358_U206 | ~new_P1_R2358_U248;
  assign new_P1_R2358_U66 = ~new_P1_R2358_U65 | ~new_P1_R2358_U202;
  assign new_P1_R2358_U67 = ~new_P1_R2358_U371 | ~new_P1_R2358_U293;
  assign new_P1_R2358_U68 = ~new_P1_R2358_U369 | ~new_P1_R2358_U291;
  assign new_P1_R2358_U69 = ~new_P1_R2358_U364 | ~new_P1_R2358_U283;
  assign new_P1_R2358_U70 = ~new_P1_R2358_U358 | ~new_P1_R2358_U275;
  assign new_P1_R2358_U71 = ~new_P1_R2358_U59 | ~new_P1_R2358_U311;
  assign new_P1_R2358_U72 = ~new_P1_R2358_U71 | ~new_P1_R2358_U255;
  assign new_P1_R2358_U73 = ~new_P1_R2358_U233 | ~new_P1_R2358_U321;
  assign new_P1_R2358_U74 = ~new_P1_R2358_U73 | ~new_P1_R2358_U262;
  assign new_P1_R2358_U75 = ~new_P1_R2358_U557 | ~new_P1_R2358_U556;
  assign new_P1_R2358_U76 = ~new_P1_R2358_U611 | ~new_P1_R2358_U610;
  assign new_P1_R2358_U77 = new_P1_R2358_U233 & new_P1_R2358_U54;
  assign new_P1_R2358_U78 = ~new_P1_R2358_U450 | ~new_P1_R2358_U449;
  assign new_P1_R2358_U79 = new_P1_R2358_U229 & new_P1_R2358_U228;
  assign new_P1_R2358_U80 = ~new_P1_R2358_U452 | ~new_P1_R2358_U451;
  assign new_P1_R2358_U81 = new_P1_R2358_U220 & new_P1_R2358_U219;
  assign new_P1_R2358_U82 = ~new_P1_R2358_U454 | ~new_P1_R2358_U453;
  assign new_P1_R2358_U83 = new_P1_R2358_U225 & new_P1_R2358_U28;
  assign new_P1_R2358_U84 = ~new_P1_R2358_U456 | ~new_P1_R2358_U455;
  assign new_P1_R2358_U85 = ~new_P1_R2358_U575 | ~new_P1_R2358_U574;
  assign new_P1_R2358_U86 = new_P1_R2358_U179 & new_P1_R2358_U300;
  assign new_P1_R2358_U87 = ~new_P1_R2358_U577 | ~new_P1_R2358_U576;
  assign new_P1_R2358_U88 = new_P1_R2358_U297 & new_P1_R2358_U296;
  assign new_P1_R2358_U89 = ~new_P1_R2358_U579 | ~new_P1_R2358_U578;
  assign new_P1_R2358_U90 = new_P1_R2358_U295 & new_P1_R2358_U294;
  assign new_P1_R2358_U91 = ~new_P1_R2358_U581 | ~new_P1_R2358_U580;
  assign new_P1_R2358_U92 = new_P1_R2358_U293 & new_P1_R2358_U292;
  assign new_P1_R2358_U93 = ~new_P1_R2358_U583 | ~new_P1_R2358_U582;
  assign new_P1_R2358_U94 = new_P1_R2358_U291 & new_P1_R2358_U290;
  assign new_P1_R2358_U95 = ~new_P1_R2358_U585 | ~new_P1_R2358_U584;
  assign new_P1_R2358_U96 = new_P1_R2358_U289 & new_P1_R2358_U288;
  assign new_P1_R2358_U97 = ~new_P1_R2358_U587 | ~new_P1_R2358_U586;
  assign new_P1_R2358_U98 = new_P1_R2358_U42 & new_P1_R2358_U286;
  assign new_P1_R2358_U99 = ~new_P1_R2358_U589 | ~new_P1_R2358_U588;
  assign new_P1_R2358_U100 = new_P1_R2358_U285 & new_P1_R2358_U284;
  assign new_P1_R2358_U101 = ~new_P1_R2358_U591 | ~new_P1_R2358_U590;
  assign new_P1_R2358_U102 = new_P1_R2358_U283 & new_P1_R2358_U282;
  assign new_P1_R2358_U103 = ~new_P1_R2358_U593 | ~new_P1_R2358_U592;
  assign new_P1_R2358_U104 = new_P1_R2358_U281 & new_P1_R2358_U280;
  assign new_P1_R2358_U105 = ~new_P1_R2358_U595 | ~new_P1_R2358_U594;
  assign new_P1_R2358_U106 = new_P1_R2358_U206 & new_P1_R2358_U205;
  assign new_P1_R2358_U107 = ~new_P1_R2358_U597 | ~new_P1_R2358_U596;
  assign new_P1_R2358_U108 = new_P1_R2358_U47 & new_P1_R2358_U278;
  assign new_P1_R2358_U109 = ~new_P1_R2358_U599 | ~new_P1_R2358_U598;
  assign new_P1_R2358_U110 = new_P1_R2358_U277 & new_P1_R2358_U276;
  assign new_P1_R2358_U111 = ~new_P1_R2358_U601 | ~new_P1_R2358_U600;
  assign new_P1_R2358_U112 = new_P1_R2358_U275 & new_P1_R2358_U274;
  assign new_P1_R2358_U113 = ~new_P1_R2358_U603 | ~new_P1_R2358_U602;
  assign new_P1_R2358_U114 = new_P1_R2358_U51 & new_P1_R2358_U272;
  assign new_P1_R2358_U115 = ~new_P1_R2358_U605 | ~new_P1_R2358_U604;
  assign new_P1_R2358_U116 = new_P1_R2358_U59 & new_P1_R2358_U258;
  assign new_P1_R2358_U117 = ~new_P1_R2358_U607 | ~new_P1_R2358_U606;
  assign new_P1_R2358_U118 = new_P1_R2358_U57 & new_P1_R2358_U259;
  assign new_P1_R2358_U119 = ~new_P1_R2358_U609 | ~new_P1_R2358_U608;
  assign new_P1_R2358_U120 = new_P1_R2358_U208 & new_P1_R2358_U205;
  assign new_P1_R2358_U121 = new_P1_R2358_U204 & new_P1_R2358_U202;
  assign new_P1_R2358_U122 = new_P1_R2358_U217 & new_P1_R2358_U216;
  assign new_P1_R2358_U123 = new_P1_R2358_U204 & new_P1_R2358_U203;
  assign new_P1_R2358_U124 = new_P1_R2358_U229 & new_P1_R2358_U54;
  assign new_P1_R2358_U125 = new_P1_R2358_U265 & new_P1_R2358_U262;
  assign new_P1_R2358_U126 = new_P1_R2358_U356 & new_P1_R2358_U255 & new_P1_R2358_U258 & new_P1_R2358_U259;
  assign new_P1_R2358_U127 = new_P1_R2358_U354 & new_P1_R2358_U355 & new_P1_R2358_U256 & new_P1_R2358_U353;
  assign new_P1_R2358_U128 = new_P1_R2358_U276 & new_P1_R2358_U5;
  assign new_P1_R2358_U129 = new_P1_R2358_U361 & new_P1_R2358_U277;
  assign new_P1_R2358_U130 = new_P1_R2358_U7 & new_P1_R2358_U284;
  assign new_P1_R2358_U131 = new_P1_R2358_U366 & new_P1_R2358_U285;
  assign new_P1_R2358_U132 = new_P1_R2358_U10 & new_P1_R2358_U294;
  assign new_P1_R2358_U133 = new_P1_R2358_U373 & new_P1_R2358_U295;
  assign new_P1_R2358_U134 = new_P1_R2358_U561 & new_P1_R2358_U305;
  assign new_P1_R2358_U135 = new_P1_R2358_U304 & new_P1_R2358_U13;
  assign new_P1_R2358_U136 = new_P1_R2358_U180 & new_P1_R2358_U374;
  assign new_P1_R2358_U137 = new_P1_R2358_U367 & new_P1_R2358_U289;
  assign new_P1_R2358_U138 = new_P1_R2358_U362 & new_P1_R2358_U281;
  assign new_P1_R2358_U139 = new_P1_R2358_U257 & new_P1_R2358_U256;
  assign new_P1_R2358_U140 = new_P1_R2358_U316 & new_P1_R2358_U61;
  assign new_P1_R2358_U141 = new_P1_R2358_U265 & new_P1_R2358_U264;
  assign new_P1_R2358_U142 = new_P1_R2358_U326 & new_P1_R2358_U263;
  assign new_P1_R2358_U143 = ~new_P1_U2618;
  assign new_P1_R2358_U144 = ~new_P1_U2615;
  assign new_P1_R2358_U145 = ~new_P1_U2614;
  assign new_P1_R2358_U146 = ~new_P1_U2667;
  assign new_P1_R2358_U147 = ~new_P1_U2668;
  assign new_P1_R2358_U148 = ~new_P1_U2670;
  assign new_P1_R2358_U149 = ~new_P1_U2671;
  assign new_P1_R2358_U150 = ~new_P1_U2672;
  assign new_P1_R2358_U151 = ~new_P1_U2669;
  assign new_P1_R2358_U152 = ~new_P1_U2617;
  assign new_P1_R2358_U153 = ~new_P1_R2358_U228 | ~new_P1_R2358_U230;
  assign new_P1_R2358_U154 = ~new_P1_R2358_U224 | ~new_P1_R2358_U226 | ~new_P1_R2358_U216;
  assign new_P1_R2358_U155 = ~new_P1_R2358_U28 | ~new_P1_R2358_U234;
  assign new_P1_R2358_U156 = ~new_P1_R2358_U203 | ~new_P1_R2358_U213;
  assign new_P1_R2358_U157 = ~new_P1_U2611;
  assign new_P1_R2358_U158 = ~new_P1_U2612;
  assign new_P1_R2358_U159 = ~new_P1_U2613;
  assign new_P1_R2358_U160 = ~new_P1_U2616;
  assign new_P1_R2358_U161 = ~new_P1_U2610;
  assign new_P1_R2358_U162 = ~new_P1_U2609;
  assign new_P1_R2358_U163 = ~new_P1_U2666;
  assign new_P1_R2358_U164 = ~new_P1_U2665;
  assign new_P1_R2358_U165 = ~new_P1_U2664;
  assign new_P1_R2358_U166 = ~new_P1_U2660;
  assign new_P1_R2358_U167 = ~new_P1_U2661;
  assign new_P1_R2358_U168 = ~new_P1_U2663;
  assign new_P1_R2358_U169 = ~new_P1_U2662;
  assign new_P1_R2358_U170 = ~new_P1_U2655;
  assign new_P1_R2358_U171 = ~new_P1_U2656;
  assign new_P1_R2358_U172 = ~new_P1_U2657;
  assign new_P1_R2358_U173 = ~new_P1_U2659;
  assign new_P1_R2358_U174 = ~new_P1_U2658;
  assign new_P1_R2358_U175 = ~new_P1_U2654;
  assign new_P1_R2358_U176 = ~new_P1_U2653;
  assign new_P1_R2358_U177 = ~new_P1_U2651;
  assign new_P1_R2358_U178 = ~new_P1_U2652;
  assign new_P1_R2358_U179 = ~new_P1_U2621 | ~new_P1_R2358_U564;
  assign new_P1_R2358_U180 = new_P1_R2358_U568 & new_P1_R2358_U567;
  assign new_P1_R2358_U181 = new_P1_R2358_U570 & new_P1_R2358_U569;
  assign new_P1_R2358_U182 = ~new_P1_R2358_U179 | ~new_P1_R2358_U302;
  assign new_P1_R2358_U183 = ~new_P1_R2358_U297 | ~new_P1_R2358_U298;
  assign new_P1_R2358_U184 = ~new_P1_R2358_U133 | ~new_P1_R2358_U383;
  assign new_P1_R2358_U185 = ~new_P1_R2358_U372 | ~new_P1_R2358_U381;
  assign new_P1_R2358_U186 = ~new_P1_R2358_U370 | ~new_P1_R2358_U379;
  assign new_P1_R2358_U187 = ~new_P1_R2358_U137 | ~new_P1_R2358_U377;
  assign new_P1_R2358_U188 = ~new_P1_R2358_U375 | ~new_P1_R2358_U42;
  assign new_P1_R2358_U189 = ~new_P1_R2358_U131 | ~new_P1_R2358_U385;
  assign new_P1_R2358_U190 = ~new_P1_R2358_U365 | ~new_P1_R2358_U387;
  assign new_P1_R2358_U191 = ~new_P1_R2358_U138 | ~new_P1_R2358_U389;
  assign new_P1_R2358_U192 = ~new_P1_R2358_U391 | ~new_P1_R2358_U47;
  assign new_P1_R2358_U193 = ~new_P1_R2358_U209 | ~new_P1_R2358_U246;
  assign new_P1_R2358_U194 = ~new_P1_R2358_U129 | ~new_P1_R2358_U393;
  assign new_P1_R2358_U195 = ~new_P1_R2358_U359 | ~new_P1_R2358_U395;
  assign new_P1_R2358_U196 = ~new_P1_R2358_U397 | ~new_P1_R2358_U51;
  assign new_P1_R2358_U197 = ~new_P1_R2358_U201 | ~new_P1_R2358_U127;
  assign new_P1_R2358_U198 = ~new_P1_R2358_U57 | ~new_P1_R2358_U309;
  assign new_P1_R2358_U199 = ~new_P1_R2358_U267 | ~new_P1_R2358_U268 | ~new_P1_R2358_U264;
  assign new_P1_R2358_U200 = ~new_P1_R2358_U209 | ~new_P1_R2358_U208;
  assign new_P1_R2358_U201 = ~new_P1_R2358_U126 | ~new_P1_R2358_U199;
  assign new_P1_R2358_U202 = ~new_P1_R2358_U30 | ~new_P1_R2358_U436 | ~new_P1_R2358_U435;
  assign new_P1_R2358_U203 = ~new_P1_U2647 | ~new_P1_R2358_U441;
  assign new_P1_R2358_U204 = ~new_P1_R2358_U32 | ~new_P1_R2358_U438 | ~new_P1_R2358_U437;
  assign new_P1_R2358_U205 = ~new_P1_R2358_U29 | ~new_P1_R2358_U432 | ~new_P1_R2358_U431;
  assign new_P1_R2358_U206 = ~new_P1_U2649 | ~new_P1_R2358_U427;
  assign new_P1_R2358_U207 = ~new_P1_U2648 | ~new_P1_R2358_U424;
  assign new_P1_R2358_U208 = ~new_P1_R2358_U31 | ~new_P1_R2358_U434 | ~new_P1_R2358_U433;
  assign new_P1_R2358_U209 = ~new_P1_U2650 | ~new_P1_R2358_U430;
  assign new_P1_R2358_U210 = ~new_P1_R2358_U209 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U211 = ~new_P1_R2358_U120 | ~new_P1_R2358_U210;
  assign new_P1_R2358_U212 = ~new_P1_R2358_U207 | ~new_P1_R2358_U211 | ~new_P1_R2358_U206;
  assign new_P1_R2358_U213 = ~new_P1_R2358_U121 | ~new_P1_R2358_U212;
  assign new_P1_R2358_U214 = ~new_P1_R2358_U156;
  assign new_P1_R2358_U215 = ~new_P1_U2644 | ~new_P1_R2358_U408;
  assign new_P1_R2358_U216 = ~new_P1_U2643 | ~new_P1_R2358_U421;
  assign new_P1_R2358_U217 = ~new_P1_R2358_U24 | ~new_P1_R2358_U405 | ~new_P1_R2358_U404;
  assign new_P1_R2358_U218 = ~new_P1_R2358_U25 | ~new_P1_R2358_U418 | ~new_P1_R2358_U417;
  assign new_P1_R2358_U219 = ~new_P1_R2358_U26 | ~new_P1_R2358_U410 | ~new_P1_R2358_U409;
  assign new_P1_R2358_U220 = ~new_P1_U2645 | ~new_P1_R2358_U416;
  assign new_P1_R2358_U221 = ~new_P1_R2358_U28;
  assign new_P1_R2358_U222 = ~new_P1_R2358_U221 | ~new_P1_R2358_U219;
  assign new_P1_R2358_U223 = ~new_P1_R2358_U215 | ~new_P1_R2358_U220 | ~new_P1_R2358_U222;
  assign new_P1_R2358_U224 = ~new_P1_R2358_U217 | ~new_P1_R2358_U218 | ~new_P1_R2358_U223;
  assign new_P1_R2358_U225 = ~new_P1_R2358_U27 | ~new_P1_R2358_U443 | ~new_P1_R2358_U442;
  assign new_P1_R2358_U226 = ~new_P1_R2358_U217 | ~new_P1_R2358_U218 | ~new_P1_R2358_U219 | ~new_P1_R2358_U225 | ~new_P1_R2358_U156;
  assign new_P1_R2358_U227 = ~new_P1_R2358_U154;
  assign new_P1_R2358_U228 = ~new_P1_U2642 | ~new_P1_R2358_U448;
  assign new_P1_R2358_U229 = ~new_P1_R2358_U33 | ~new_P1_R2358_U445 | ~new_P1_R2358_U444;
  assign new_P1_R2358_U230 = ~new_P1_R2358_U229 | ~new_P1_R2358_U154;
  assign new_P1_R2358_U231 = ~new_P1_R2358_U153;
  assign new_P1_R2358_U232 = ~new_P1_R2358_U54;
  assign new_P1_R2358_U233 = ~new_P1_U2641 | ~new_P1_R2358_U403;
  assign new_P1_R2358_U234 = ~new_P1_R2358_U225 | ~new_P1_R2358_U156;
  assign new_P1_R2358_U235 = ~new_P1_R2358_U155;
  assign new_P1_R2358_U236 = ~new_P1_R2358_U155 | ~new_P1_R2358_U219;
  assign new_P1_R2358_U237 = ~new_P1_R2358_U35;
  assign new_P1_R2358_U238 = ~new_P1_R2358_U36;
  assign new_P1_R2358_U239 = ~new_P1_R2358_U36 | ~new_P1_R2358_U215;
  assign new_P1_R2358_U240 = ~new_P1_R2358_U122 | ~new_P1_R2358_U239;
  assign new_P1_R2358_U241 = ~new_P1_R2358_U217 | ~new_P1_R2358_U216;
  assign new_P1_R2358_U242 = ~new_P1_R2358_U241 | ~new_P1_R2358_U36 | ~new_P1_R2358_U215;
  assign new_P1_R2358_U243 = ~new_P1_R2358_U218 | ~new_P1_R2358_U215;
  assign new_P1_R2358_U244 = ~new_P1_R2358_U237 | ~new_P1_R2358_U243;
  assign new_P1_R2358_U245 = ~new_P1_R2358_U238 | ~new_P1_R2358_U215;
  assign new_P1_R2358_U246 = ~new_P1_U2352 | ~new_P1_R2358_U208;
  assign new_P1_R2358_U247 = ~new_P1_R2358_U193;
  assign new_P1_R2358_U248 = ~new_P1_R2358_U193 | ~new_P1_R2358_U205;
  assign new_P1_R2358_U249 = ~new_P1_R2358_U65;
  assign new_P1_R2358_U250 = ~new_P1_R2358_U66;
  assign new_P1_R2358_U251 = ~new_P1_R2358_U66 | ~new_P1_R2358_U207;
  assign new_P1_R2358_U252 = ~new_P1_R2358_U123 | ~new_P1_R2358_U251;
  assign new_P1_R2358_U253 = ~new_P1_R2358_U204 | ~new_P1_R2358_U203;
  assign new_P1_R2358_U254 = ~new_P1_R2358_U253 | ~new_P1_R2358_U66 | ~new_P1_R2358_U207;
  assign new_P1_R2358_U255 = ~new_P1_R2358_U60 | ~new_P1_R2358_U460 | ~new_P1_R2358_U459;
  assign new_P1_R2358_U256 = ~new_P1_U2635 | ~new_P1_R2358_U474;
  assign new_P1_R2358_U257 = ~new_P1_R2358_U11 | ~new_P1_R2358_U55;
  assign new_P1_R2358_U258 = ~new_P1_R2358_U58 | ~new_P1_R2358_U468 | ~new_P1_R2358_U467;
  assign new_P1_R2358_U259 = ~new_P1_R2358_U56 | ~new_P1_R2358_U486 | ~new_P1_R2358_U485;
  assign new_P1_R2358_U260 = ~new_P1_R2358_U59;
  assign new_P1_R2358_U261 = ~new_P1_R2358_U61;
  assign new_P1_R2358_U262 = ~new_P1_R2358_U53 | ~new_P1_R2358_U476 | ~new_P1_R2358_U475;
  assign new_P1_R2358_U263 = ~new_P1_U2640 | ~new_P1_R2358_U479;
  assign new_P1_R2358_U264 = ~new_P1_U2639 | ~new_P1_R2358_U484;
  assign new_P1_R2358_U265 = ~new_P1_R2358_U12 | ~new_P1_R2358_U52;
  assign new_P1_R2358_U266 = ~new_P1_R2358_U263 | ~new_P1_R2358_U233 | ~new_P1_R2358_U228;
  assign new_P1_R2358_U267 = ~new_P1_R2358_U262 | ~new_P1_R2358_U266 | ~new_P1_R2358_U360 | ~new_P1_R2358_U357;
  assign new_P1_R2358_U268 = ~new_P1_R2358_U125 | ~new_P1_R2358_U124 | ~new_P1_R2358_U154;
  assign new_P1_R2358_U269 = ~new_P1_R2358_U199;
  assign new_P1_R2358_U270 = ~new_P1_R2358_U57;
  assign new_P1_R2358_U271 = ~new_P1_R2358_U197;
  assign new_P1_R2358_U272 = ~new_P1_R2358_U50 | ~new_P1_R2358_U488 | ~new_P1_R2358_U487;
  assign new_P1_R2358_U273 = ~new_P1_R2358_U51;
  assign new_P1_R2358_U274 = ~new_P1_R2358_U49 | ~new_P1_R2358_U490 | ~new_P1_R2358_U489;
  assign new_P1_R2358_U275 = ~new_P1_U2633 | ~new_P1_R2358_U498;
  assign new_P1_R2358_U276 = ~new_P1_R2358_U48 | ~new_P1_R2358_U492 | ~new_P1_R2358_U491;
  assign new_P1_R2358_U277 = ~new_P1_U2632 | ~new_P1_R2358_U495;
  assign new_P1_R2358_U278 = ~new_P1_R2358_U46 | ~new_P1_R2358_U507 | ~new_P1_R2358_U506;
  assign new_P1_R2358_U279 = ~new_P1_R2358_U47;
  assign new_P1_R2358_U280 = ~new_P1_R2358_U45 | ~new_P1_R2358_U509 | ~new_P1_R2358_U508;
  assign new_P1_R2358_U281 = ~new_P1_U2630 | ~new_P1_R2358_U518;
  assign new_P1_R2358_U282 = ~new_P1_R2358_U44 | ~new_P1_R2358_U505 | ~new_P1_R2358_U504;
  assign new_P1_R2358_U283 = ~new_P1_U2629 | ~new_P1_R2358_U515;
  assign new_P1_R2358_U284 = ~new_P1_R2358_U43 | ~new_P1_R2358_U503 | ~new_P1_R2358_U502;
  assign new_P1_R2358_U285 = ~new_P1_U2628 | ~new_P1_R2358_U512;
  assign new_P1_R2358_U286 = ~new_P1_R2358_U41 | ~new_P1_R2358_U529 | ~new_P1_R2358_U528;
  assign new_P1_R2358_U287 = ~new_P1_R2358_U42;
  assign new_P1_R2358_U288 = ~new_P1_R2358_U40 | ~new_P1_R2358_U531 | ~new_P1_R2358_U530;
  assign new_P1_R2358_U289 = ~new_P1_U2626 | ~new_P1_R2358_U543;
  assign new_P1_R2358_U290 = ~new_P1_R2358_U39 | ~new_P1_R2358_U527 | ~new_P1_R2358_U526;
  assign new_P1_R2358_U291 = ~new_P1_U2625 | ~new_P1_R2358_U540;
  assign new_P1_R2358_U292 = ~new_P1_R2358_U38 | ~new_P1_R2358_U525 | ~new_P1_R2358_U524;
  assign new_P1_R2358_U293 = ~new_P1_U2624 | ~new_P1_R2358_U537;
  assign new_P1_R2358_U294 = ~new_P1_R2358_U37 | ~new_P1_R2358_U523 | ~new_P1_R2358_U522;
  assign new_P1_R2358_U295 = ~new_P1_U2623 | ~new_P1_R2358_U534;
  assign new_P1_R2358_U296 = ~new_P1_R2358_U62 | ~new_P1_R2358_U548 | ~new_P1_R2358_U547;
  assign new_P1_R2358_U297 = ~new_P1_U2622 | ~new_P1_R2358_U551;
  assign new_P1_R2358_U298 = ~new_P1_R2358_U296 | ~new_P1_R2358_U184;
  assign new_P1_R2358_U299 = ~new_P1_R2358_U183;
  assign new_P1_R2358_U300 = ~new_P1_R2358_U64 | ~new_P1_R2358_U553 | ~new_P1_R2358_U552;
  assign new_P1_R2358_U301 = ~new_P1_R2358_U179;
  assign new_P1_R2358_U302 = ~new_P1_R2358_U300 | ~new_P1_R2358_U183;
  assign new_P1_R2358_U303 = ~new_P1_R2358_U182;
  assign new_P1_R2358_U304 = ~new_P1_U2620 | ~new_P1_R2358_U75;
  assign new_P1_R2358_U305 = ~new_P1_R2358_U558 | ~new_P1_R2358_U63;
  assign new_P1_R2358_U306 = ~new_P1_R2358_U207 | ~new_P1_R2358_U202;
  assign new_P1_R2358_U307 = ~new_P1_R2358_U249 | ~new_P1_R2358_U306;
  assign new_P1_R2358_U308 = ~new_P1_R2358_U250 | ~new_P1_R2358_U207;
  assign new_P1_R2358_U309 = ~new_P1_R2358_U199 | ~new_P1_R2358_U259;
  assign new_P1_R2358_U310 = ~new_P1_R2358_U198;
  assign new_P1_R2358_U311 = ~new_P1_R2358_U198 | ~new_P1_R2358_U258;
  assign new_P1_R2358_U312 = ~new_P1_R2358_U71;
  assign new_P1_R2358_U313 = ~new_P1_R2358_U72;
  assign new_P1_R2358_U314 = ~new_P1_R2358_U72 | ~new_P1_R2358_U61;
  assign new_P1_R2358_U315 = ~new_P1_R2358_U139 | ~new_P1_R2358_U314;
  assign new_P1_R2358_U316 = ~new_P1_R2358_U257 | ~new_P1_R2358_U256;
  assign new_P1_R2358_U317 = ~new_P1_R2358_U140 | ~new_P1_R2358_U72;
  assign new_P1_R2358_U318 = ~new_P1_R2358_U61 | ~new_P1_R2358_U255;
  assign new_P1_R2358_U319 = ~new_P1_R2358_U312 | ~new_P1_R2358_U318;
  assign new_P1_R2358_U320 = ~new_P1_R2358_U313 | ~new_P1_R2358_U61;
  assign new_P1_R2358_U321 = ~new_P1_R2358_U54 | ~new_P1_R2358_U153;
  assign new_P1_R2358_U322 = ~new_P1_R2358_U73;
  assign new_P1_R2358_U323 = ~new_P1_R2358_U74;
  assign new_P1_R2358_U324 = ~new_P1_R2358_U74 | ~new_P1_R2358_U263;
  assign new_P1_R2358_U325 = ~new_P1_R2358_U141 | ~new_P1_R2358_U324;
  assign new_P1_R2358_U326 = ~new_P1_R2358_U265 | ~new_P1_R2358_U264;
  assign new_P1_R2358_U327 = ~new_P1_R2358_U142 | ~new_P1_R2358_U74;
  assign new_P1_R2358_U328 = ~new_P1_R2358_U263 | ~new_P1_R2358_U262;
  assign new_P1_R2358_U329 = ~new_P1_R2358_U322 | ~new_P1_R2358_U328;
  assign new_P1_R2358_U330 = ~new_P1_R2358_U323 | ~new_P1_R2358_U263;
  assign new_P1_R2358_U331 = ~new_P1_R2358_U200;
  assign new_P1_R2358_U332 = ~new_P1_R2358_U233 | ~new_P1_R2358_U54;
  assign new_P1_R2358_U333 = ~new_P1_R2358_U229 | ~new_P1_R2358_U228;
  assign new_P1_R2358_U334 = ~new_P1_R2358_U220 | ~new_P1_R2358_U219;
  assign new_P1_R2358_U335 = ~new_P1_R2358_U225 | ~new_P1_R2358_U28;
  assign new_P1_R2358_U336 = ~new_P1_R2358_U179 | ~new_P1_R2358_U300;
  assign new_P1_R2358_U337 = ~new_P1_R2358_U297 | ~new_P1_R2358_U296;
  assign new_P1_R2358_U338 = ~new_P1_R2358_U295 | ~new_P1_R2358_U294;
  assign new_P1_R2358_U339 = ~new_P1_R2358_U293 | ~new_P1_R2358_U292;
  assign new_P1_R2358_U340 = ~new_P1_R2358_U291 | ~new_P1_R2358_U290;
  assign new_P1_R2358_U341 = ~new_P1_R2358_U289 | ~new_P1_R2358_U288;
  assign new_P1_R2358_U342 = ~new_P1_R2358_U42 | ~new_P1_R2358_U286;
  assign new_P1_R2358_U343 = ~new_P1_R2358_U285 | ~new_P1_R2358_U284;
  assign new_P1_R2358_U344 = ~new_P1_R2358_U283 | ~new_P1_R2358_U282;
  assign new_P1_R2358_U345 = ~new_P1_R2358_U281 | ~new_P1_R2358_U280;
  assign new_P1_R2358_U346 = ~new_P1_R2358_U206 | ~new_P1_R2358_U205;
  assign new_P1_R2358_U347 = ~new_P1_R2358_U47 | ~new_P1_R2358_U278;
  assign new_P1_R2358_U348 = ~new_P1_R2358_U277 | ~new_P1_R2358_U276;
  assign new_P1_R2358_U349 = ~new_P1_R2358_U275 | ~new_P1_R2358_U274;
  assign new_P1_R2358_U350 = ~new_P1_R2358_U51 | ~new_P1_R2358_U272;
  assign new_P1_R2358_U351 = ~new_P1_R2358_U59 | ~new_P1_R2358_U258;
  assign new_P1_R2358_U352 = ~new_P1_R2358_U57 | ~new_P1_R2358_U259;
  assign new_P1_R2358_U353 = ~new_P1_R2358_U257 | ~new_P1_R2358_U255 | ~new_P1_R2358_U270 | ~new_P1_R2358_U258;
  assign new_P1_R2358_U354 = ~new_P1_R2358_U257 | ~new_P1_R2358_U260 | ~new_P1_R2358_U255;
  assign new_P1_R2358_U355 = ~new_P1_R2358_U261 | ~new_P1_R2358_U257;
  assign new_P1_R2358_U356 = ~new_P1_R2358_U11 | ~new_P1_R2358_U55;
  assign new_P1_R2358_U357 = ~new_P1_R2358_U232 | ~new_P1_R2358_U263;
  assign new_P1_R2358_U358 = ~new_P1_R2358_U273 | ~new_P1_R2358_U274;
  assign new_P1_R2358_U359 = ~new_P1_R2358_U70;
  assign new_P1_R2358_U360 = ~new_P1_R2358_U12 | ~new_P1_R2358_U52;
  assign new_P1_R2358_U361 = ~new_P1_R2358_U70 | ~new_P1_R2358_U276;
  assign new_P1_R2358_U362 = ~new_P1_R2358_U279 | ~new_P1_R2358_U280;
  assign new_P1_R2358_U363 = ~new_P1_R2358_U362 | ~new_P1_R2358_U281;
  assign new_P1_R2358_U364 = ~new_P1_R2358_U363 | ~new_P1_R2358_U282;
  assign new_P1_R2358_U365 = ~new_P1_R2358_U69;
  assign new_P1_R2358_U366 = ~new_P1_R2358_U69 | ~new_P1_R2358_U284;
  assign new_P1_R2358_U367 = ~new_P1_R2358_U287 | ~new_P1_R2358_U288;
  assign new_P1_R2358_U368 = ~new_P1_R2358_U367 | ~new_P1_R2358_U289;
  assign new_P1_R2358_U369 = ~new_P1_R2358_U368 | ~new_P1_R2358_U290;
  assign new_P1_R2358_U370 = ~new_P1_R2358_U68;
  assign new_P1_R2358_U371 = ~new_P1_R2358_U68 | ~new_P1_R2358_U292;
  assign new_P1_R2358_U372 = ~new_P1_R2358_U67;
  assign new_P1_R2358_U373 = ~new_P1_R2358_U67 | ~new_P1_R2358_U294;
  assign new_P1_R2358_U374 = ~new_P1_R2358_U134 | ~new_P1_R2358_U300 | ~new_P1_R2358_U183;
  assign new_P1_R2358_U375 = ~new_P1_R2358_U286 | ~new_P1_R2358_U189;
  assign new_P1_R2358_U376 = ~new_P1_R2358_U188;
  assign new_P1_R2358_U377 = ~new_P1_R2358_U8 | ~new_P1_R2358_U189;
  assign new_P1_R2358_U378 = ~new_P1_R2358_U187;
  assign new_P1_R2358_U379 = ~new_P1_R2358_U9 | ~new_P1_R2358_U189;
  assign new_P1_R2358_U380 = ~new_P1_R2358_U186;
  assign new_P1_R2358_U381 = ~new_P1_R2358_U10 | ~new_P1_R2358_U189;
  assign new_P1_R2358_U382 = ~new_P1_R2358_U185;
  assign new_P1_R2358_U383 = ~new_P1_R2358_U132 | ~new_P1_R2358_U189;
  assign new_P1_R2358_U384 = ~new_P1_R2358_U184;
  assign new_P1_R2358_U385 = ~new_P1_R2358_U130 | ~new_P1_R2358_U194;
  assign new_P1_R2358_U386 = ~new_P1_R2358_U189;
  assign new_P1_R2358_U387 = ~new_P1_R2358_U7 | ~new_P1_R2358_U194;
  assign new_P1_R2358_U388 = ~new_P1_R2358_U190;
  assign new_P1_R2358_U389 = ~new_P1_R2358_U6 | ~new_P1_R2358_U194;
  assign new_P1_R2358_U390 = ~new_P1_R2358_U191;
  assign new_P1_R2358_U391 = ~new_P1_R2358_U278 | ~new_P1_R2358_U194;
  assign new_P1_R2358_U392 = ~new_P1_R2358_U192;
  assign new_P1_R2358_U393 = ~new_P1_R2358_U128 | ~new_P1_R2358_U197;
  assign new_P1_R2358_U394 = ~new_P1_R2358_U194;
  assign new_P1_R2358_U395 = ~new_P1_R2358_U5 | ~new_P1_R2358_U197;
  assign new_P1_R2358_U396 = ~new_P1_R2358_U195;
  assign new_P1_R2358_U397 = ~new_P1_R2358_U272 | ~new_P1_R2358_U197;
  assign new_P1_R2358_U398 = ~new_P1_R2358_U196;
  assign new_P1_R2358_U399 = ~new_P1_U2352 | ~new_P1_R2358_U143;
  assign new_P1_R2358_U400 = ~new_P1_U2618 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U401 = ~new_P1_U2352 | ~new_P1_R2358_U143;
  assign new_P1_R2358_U402 = ~new_P1_U2618 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U403 = ~new_P1_R2358_U402 | ~new_P1_R2358_U401;
  assign new_P1_R2358_U404 = ~new_P1_U2352 | ~new_P1_R2358_U144;
  assign new_P1_R2358_U405 = ~new_P1_U2615 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U406 = ~new_P1_U2352 | ~new_P1_R2358_U145;
  assign new_P1_R2358_U407 = ~new_P1_U2614 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U408 = ~new_P1_R2358_U407 | ~new_P1_R2358_U406;
  assign new_P1_R2358_U409 = ~new_P1_U2352 | ~new_P1_R2358_U146;
  assign new_P1_R2358_U410 = ~new_P1_U2667 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U411 = ~new_P1_U2352 | ~new_P1_R2358_U147;
  assign new_P1_R2358_U412 = ~new_P1_U2668 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U413 = ~new_P1_R2358_U412 | ~new_P1_R2358_U411;
  assign new_P1_R2358_U414 = ~new_P1_U2352 | ~new_P1_R2358_U146;
  assign new_P1_R2358_U415 = ~new_P1_U2667 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U416 = ~new_P1_R2358_U415 | ~new_P1_R2358_U414;
  assign new_P1_R2358_U417 = ~new_P1_U2352 | ~new_P1_R2358_U145;
  assign new_P1_R2358_U418 = ~new_P1_U2614 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U419 = ~new_P1_U2352 | ~new_P1_R2358_U144;
  assign new_P1_R2358_U420 = ~new_P1_U2615 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U421 = ~new_P1_R2358_U420 | ~new_P1_R2358_U419;
  assign new_P1_R2358_U422 = ~new_P1_U2352 | ~new_P1_R2358_U148;
  assign new_P1_R2358_U423 = ~new_P1_U2670 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U424 = ~new_P1_R2358_U423 | ~new_P1_R2358_U422;
  assign new_P1_R2358_U425 = ~new_P1_U2352 | ~new_P1_R2358_U149;
  assign new_P1_R2358_U426 = ~new_P1_U2671 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U427 = ~new_P1_R2358_U426 | ~new_P1_R2358_U425;
  assign new_P1_R2358_U428 = ~new_P1_U2352 | ~new_P1_R2358_U150;
  assign new_P1_R2358_U429 = ~new_P1_U2672 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U430 = ~new_P1_R2358_U429 | ~new_P1_R2358_U428;
  assign new_P1_R2358_U431 = ~new_P1_U2352 | ~new_P1_R2358_U149;
  assign new_P1_R2358_U432 = ~new_P1_U2671 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U433 = ~new_P1_U2352 | ~new_P1_R2358_U150;
  assign new_P1_R2358_U434 = ~new_P1_U2672 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U435 = ~new_P1_U2352 | ~new_P1_R2358_U148;
  assign new_P1_R2358_U436 = ~new_P1_U2670 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U437 = ~new_P1_U2352 | ~new_P1_R2358_U151;
  assign new_P1_R2358_U438 = ~new_P1_U2669 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U439 = ~new_P1_U2352 | ~new_P1_R2358_U151;
  assign new_P1_R2358_U440 = ~new_P1_U2669 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U441 = ~new_P1_R2358_U440 | ~new_P1_R2358_U439;
  assign new_P1_R2358_U442 = ~new_P1_U2352 | ~new_P1_R2358_U147;
  assign new_P1_R2358_U443 = ~new_P1_U2668 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U444 = ~new_P1_U2352 | ~new_P1_R2358_U152;
  assign new_P1_R2358_U445 = ~new_P1_U2617 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U446 = ~new_P1_U2352 | ~new_P1_R2358_U152;
  assign new_P1_R2358_U447 = ~new_P1_U2617 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U448 = ~new_P1_R2358_U447 | ~new_P1_R2358_U446;
  assign new_P1_R2358_U449 = ~new_P1_R2358_U332 | ~new_P1_R2358_U153;
  assign new_P1_R2358_U450 = ~new_P1_R2358_U77 | ~new_P1_R2358_U231;
  assign new_P1_R2358_U451 = ~new_P1_R2358_U333 | ~new_P1_R2358_U154;
  assign new_P1_R2358_U452 = ~new_P1_R2358_U79 | ~new_P1_R2358_U227;
  assign new_P1_R2358_U453 = ~new_P1_R2358_U334 | ~new_P1_R2358_U155;
  assign new_P1_R2358_U454 = ~new_P1_R2358_U81 | ~new_P1_R2358_U235;
  assign new_P1_R2358_U455 = ~new_P1_R2358_U335 | ~new_P1_R2358_U156;
  assign new_P1_R2358_U456 = ~new_P1_R2358_U83 | ~new_P1_R2358_U214;
  assign new_P1_R2358_U457 = ~new_P1_U2352 | ~new_P1_R2358_U157;
  assign new_P1_R2358_U458 = ~new_P1_U2611 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U459 = ~new_P1_U2352 | ~new_P1_R2358_U158;
  assign new_P1_R2358_U460 = ~new_P1_U2612 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U461 = ~new_P1_U2352 | ~new_P1_R2358_U159;
  assign new_P1_R2358_U462 = ~new_P1_U2613 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U463 = ~new_P1_R2358_U462 | ~new_P1_R2358_U461;
  assign new_P1_R2358_U464 = ~new_P1_U2352 | ~new_P1_R2358_U158;
  assign new_P1_R2358_U465 = ~new_P1_U2612 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U466 = ~new_P1_R2358_U465 | ~new_P1_R2358_U464;
  assign new_P1_R2358_U467 = ~new_P1_U2352 | ~new_P1_R2358_U159;
  assign new_P1_R2358_U468 = ~new_P1_U2613 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U469 = ~new_P1_U2352 | ~new_P1_R2358_U160;
  assign new_P1_R2358_U470 = ~new_P1_U2616 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U471 = ~new_P1_R2358_U470 | ~new_P1_R2358_U469;
  assign new_P1_R2358_U472 = ~new_P1_U2352 | ~new_P1_R2358_U157;
  assign new_P1_R2358_U473 = ~new_P1_U2611 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U474 = ~new_P1_R2358_U473 | ~new_P1_R2358_U472;
  assign new_P1_R2358_U475 = ~new_P1_U2352 | ~new_P1_R2358_U161;
  assign new_P1_R2358_U476 = ~new_P1_U2610 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U477 = ~new_P1_U2352 | ~new_P1_R2358_U161;
  assign new_P1_R2358_U478 = ~new_P1_U2610 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U479 = ~new_P1_R2358_U478 | ~new_P1_R2358_U477;
  assign new_P1_R2358_U480 = ~new_P1_U2352 | ~new_P1_R2358_U162;
  assign new_P1_R2358_U481 = ~new_P1_U2609 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U482 = ~new_P1_U2352 | ~new_P1_R2358_U162;
  assign new_P1_R2358_U483 = ~new_P1_U2609 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U484 = ~new_P1_R2358_U483 | ~new_P1_R2358_U482;
  assign new_P1_R2358_U485 = ~new_P1_U2352 | ~new_P1_R2358_U160;
  assign new_P1_R2358_U486 = ~new_P1_U2616 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U487 = ~new_P1_U2352 | ~new_P1_R2358_U163;
  assign new_P1_R2358_U488 = ~new_P1_U2666 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U489 = ~new_P1_U2352 | ~new_P1_R2358_U164;
  assign new_P1_R2358_U490 = ~new_P1_U2665 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U491 = ~new_P1_U2352 | ~new_P1_R2358_U165;
  assign new_P1_R2358_U492 = ~new_P1_U2664 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U493 = ~new_P1_U2352 | ~new_P1_R2358_U165;
  assign new_P1_R2358_U494 = ~new_P1_U2664 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U495 = ~new_P1_R2358_U494 | ~new_P1_R2358_U493;
  assign new_P1_R2358_U496 = ~new_P1_U2352 | ~new_P1_R2358_U164;
  assign new_P1_R2358_U497 = ~new_P1_U2665 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U498 = ~new_P1_R2358_U497 | ~new_P1_R2358_U496;
  assign new_P1_R2358_U499 = ~new_P1_U2352 | ~new_P1_R2358_U163;
  assign new_P1_R2358_U500 = ~new_P1_U2666 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U501 = ~new_P1_R2358_U500 | ~new_P1_R2358_U499;
  assign new_P1_R2358_U502 = ~new_P1_U2352 | ~new_P1_R2358_U166;
  assign new_P1_R2358_U503 = ~new_P1_U2660 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U504 = ~new_P1_U2352 | ~new_P1_R2358_U167;
  assign new_P1_R2358_U505 = ~new_P1_U2661 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U506 = ~new_P1_U2352 | ~new_P1_R2358_U168;
  assign new_P1_R2358_U507 = ~new_P1_U2663 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U508 = ~new_P1_U2352 | ~new_P1_R2358_U169;
  assign new_P1_R2358_U509 = ~new_P1_U2662 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U510 = ~new_P1_U2352 | ~new_P1_R2358_U166;
  assign new_P1_R2358_U511 = ~new_P1_U2660 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U512 = ~new_P1_R2358_U511 | ~new_P1_R2358_U510;
  assign new_P1_R2358_U513 = ~new_P1_U2352 | ~new_P1_R2358_U167;
  assign new_P1_R2358_U514 = ~new_P1_U2661 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U515 = ~new_P1_R2358_U514 | ~new_P1_R2358_U513;
  assign new_P1_R2358_U516 = ~new_P1_U2352 | ~new_P1_R2358_U169;
  assign new_P1_R2358_U517 = ~new_P1_U2662 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U518 = ~new_P1_R2358_U517 | ~new_P1_R2358_U516;
  assign new_P1_R2358_U519 = ~new_P1_U2352 | ~new_P1_R2358_U168;
  assign new_P1_R2358_U520 = ~new_P1_U2663 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U521 = ~new_P1_R2358_U520 | ~new_P1_R2358_U519;
  assign new_P1_R2358_U522 = ~new_P1_U2352 | ~new_P1_R2358_U170;
  assign new_P1_R2358_U523 = ~new_P1_U2655 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U524 = ~new_P1_U2352 | ~new_P1_R2358_U171;
  assign new_P1_R2358_U525 = ~new_P1_U2656 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U526 = ~new_P1_U2352 | ~new_P1_R2358_U172;
  assign new_P1_R2358_U527 = ~new_P1_U2657 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U528 = ~new_P1_U2352 | ~new_P1_R2358_U173;
  assign new_P1_R2358_U529 = ~new_P1_U2659 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U530 = ~new_P1_U2352 | ~new_P1_R2358_U174;
  assign new_P1_R2358_U531 = ~new_P1_U2658 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U532 = ~new_P1_U2352 | ~new_P1_R2358_U170;
  assign new_P1_R2358_U533 = ~new_P1_U2655 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U534 = ~new_P1_R2358_U533 | ~new_P1_R2358_U532;
  assign new_P1_R2358_U535 = ~new_P1_U2352 | ~new_P1_R2358_U171;
  assign new_P1_R2358_U536 = ~new_P1_U2656 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U537 = ~new_P1_R2358_U536 | ~new_P1_R2358_U535;
  assign new_P1_R2358_U538 = ~new_P1_U2352 | ~new_P1_R2358_U172;
  assign new_P1_R2358_U539 = ~new_P1_U2657 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U540 = ~new_P1_R2358_U539 | ~new_P1_R2358_U538;
  assign new_P1_R2358_U541 = ~new_P1_U2352 | ~new_P1_R2358_U174;
  assign new_P1_R2358_U542 = ~new_P1_U2658 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U543 = ~new_P1_R2358_U542 | ~new_P1_R2358_U541;
  assign new_P1_R2358_U544 = ~new_P1_U2352 | ~new_P1_R2358_U173;
  assign new_P1_R2358_U545 = ~new_P1_U2659 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U546 = ~new_P1_R2358_U545 | ~new_P1_R2358_U544;
  assign new_P1_R2358_U547 = ~new_P1_U2352 | ~new_P1_R2358_U175;
  assign new_P1_R2358_U548 = ~new_P1_U2654 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U549 = ~new_P1_U2352 | ~new_P1_R2358_U175;
  assign new_P1_R2358_U550 = ~new_P1_U2654 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U551 = ~new_P1_R2358_U550 | ~new_P1_R2358_U549;
  assign new_P1_R2358_U552 = ~new_P1_U2352 | ~new_P1_R2358_U176;
  assign new_P1_R2358_U553 = ~new_P1_U2653 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U554 = ~new_P1_U2352 | ~new_P1_R2358_U177;
  assign new_P1_R2358_U555 = ~new_P1_U2651 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U556 = ~new_P1_U2352 | ~new_P1_R2358_U178;
  assign new_P1_R2358_U557 = ~new_P1_U2652 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U558 = ~new_P1_R2358_U75;
  assign new_P1_R2358_U559 = ~new_P1_U2352 | ~new_P1_R2358_U177;
  assign new_P1_R2358_U560 = ~new_P1_U2651 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U561 = ~new_P1_R2358_U560 | ~new_P1_R2358_U559;
  assign new_P1_R2358_U562 = ~new_P1_U2352 | ~new_P1_R2358_U176;
  assign new_P1_R2358_U563 = ~new_P1_U2653 | ~new_P1_R2358_U23;
  assign new_P1_R2358_U564 = ~new_P1_R2358_U563 | ~new_P1_R2358_U562;
  assign new_P1_R2358_U565 = ~new_P1_R2358_U179 | ~new_P1_R2358_U135 | ~new_P1_R2358_U302;
  assign new_P1_R2358_U566 = ~new_P1_R2358_U301 | ~new_P1_R2358_U561 | ~new_P1_R2358_U305;
  assign new_P1_R2358_U567 = ~new_P1_R2358_U63 | ~new_P1_R2358_U13 | ~new_P1_R2358_U558;
  assign new_P1_R2358_U568 = ~new_P1_U2620 | ~new_P1_R2358_U561 | ~new_P1_R2358_U75;
  assign new_P1_R2358_U569 = ~new_P1_R2358_U558 | ~new_P1_U2620;
  assign new_P1_R2358_U570 = ~new_P1_R2358_U75 | ~new_P1_R2358_U63;
  assign new_P1_R2358_U571 = ~new_P1_R2358_U558 | ~new_P1_U2620;
  assign new_P1_R2358_U572 = ~new_P1_R2358_U75 | ~new_P1_R2358_U63;
  assign new_P1_R2358_U573 = ~new_P1_R2358_U572 | ~new_P1_R2358_U571;
  assign new_P1_R2358_U574 = ~new_P1_R2358_U181 | ~new_P1_R2358_U182;
  assign new_P1_R2358_U575 = ~new_P1_R2358_U303 | ~new_P1_R2358_U573;
  assign new_P1_R2358_U576 = ~new_P1_R2358_U336 | ~new_P1_R2358_U183;
  assign new_P1_R2358_U577 = ~new_P1_R2358_U86 | ~new_P1_R2358_U299;
  assign new_P1_R2358_U578 = ~new_P1_R2358_U184 | ~new_P1_R2358_U337;
  assign new_P1_R2358_U579 = ~new_P1_R2358_U88 | ~new_P1_R2358_U384;
  assign new_P1_R2358_U580 = ~new_P1_R2358_U185 | ~new_P1_R2358_U338;
  assign new_P1_R2358_U581 = ~new_P1_R2358_U90 | ~new_P1_R2358_U382;
  assign new_P1_R2358_U582 = ~new_P1_R2358_U186 | ~new_P1_R2358_U339;
  assign new_P1_R2358_U583 = ~new_P1_R2358_U92 | ~new_P1_R2358_U380;
  assign new_P1_R2358_U584 = ~new_P1_R2358_U187 | ~new_P1_R2358_U340;
  assign new_P1_R2358_U585 = ~new_P1_R2358_U94 | ~new_P1_R2358_U378;
  assign new_P1_R2358_U586 = ~new_P1_R2358_U188 | ~new_P1_R2358_U341;
  assign new_P1_R2358_U587 = ~new_P1_R2358_U96 | ~new_P1_R2358_U376;
  assign new_P1_R2358_U588 = ~new_P1_R2358_U189 | ~new_P1_R2358_U342;
  assign new_P1_R2358_U589 = ~new_P1_R2358_U98 | ~new_P1_R2358_U386;
  assign new_P1_R2358_U590 = ~new_P1_R2358_U190 | ~new_P1_R2358_U343;
  assign new_P1_R2358_U591 = ~new_P1_R2358_U100 | ~new_P1_R2358_U388;
  assign new_P1_R2358_U592 = ~new_P1_R2358_U191 | ~new_P1_R2358_U344;
  assign new_P1_R2358_U593 = ~new_P1_R2358_U102 | ~new_P1_R2358_U390;
  assign new_P1_R2358_U594 = ~new_P1_R2358_U192 | ~new_P1_R2358_U345;
  assign new_P1_R2358_U595 = ~new_P1_R2358_U104 | ~new_P1_R2358_U392;
  assign new_P1_R2358_U596 = ~new_P1_R2358_U346 | ~new_P1_R2358_U193;
  assign new_P1_R2358_U597 = ~new_P1_R2358_U106 | ~new_P1_R2358_U247;
  assign new_P1_R2358_U598 = ~new_P1_R2358_U194 | ~new_P1_R2358_U347;
  assign new_P1_R2358_U599 = ~new_P1_R2358_U108 | ~new_P1_R2358_U394;
  assign new_P1_R2358_U600 = ~new_P1_R2358_U195 | ~new_P1_R2358_U348;
  assign new_P1_R2358_U601 = ~new_P1_R2358_U110 | ~new_P1_R2358_U396;
  assign new_P1_R2358_U602 = ~new_P1_R2358_U196 | ~new_P1_R2358_U349;
  assign new_P1_R2358_U603 = ~new_P1_R2358_U112 | ~new_P1_R2358_U398;
  assign new_P1_R2358_U604 = ~new_P1_R2358_U350 | ~new_P1_R2358_U197;
  assign new_P1_R2358_U605 = ~new_P1_R2358_U114 | ~new_P1_R2358_U271;
  assign new_P1_R2358_U606 = ~new_P1_R2358_U351 | ~new_P1_R2358_U198;
  assign new_P1_R2358_U607 = ~new_P1_R2358_U116 | ~new_P1_R2358_U310;
  assign new_P1_R2358_U608 = ~new_P1_R2358_U352 | ~new_P1_R2358_U199;
  assign new_P1_R2358_U609 = ~new_P1_R2358_U118 | ~new_P1_R2358_U269;
  assign new_P1_R2358_U610 = ~new_P1_U2352 | ~new_P1_R2358_U200;
  assign new_P1_R2358_U611 = ~new_P1_R2358_U331 | ~new_P1_R2358_U23;
  assign new_P1_LT_589_U6 = new_P1_LT_589_U8 | new_P1_U2673;
  assign new_P1_LT_589_U7 = new_P1_R584_U7 & new_P1_R584_U6;
  assign new_P1_LT_589_U8 = ~new_P1_R584_U8 & ~new_P1_LT_589_U7 & ~new_P1_R584_U9;
  assign new_P1_R584_U6 = ~new_P1_U2676;
  assign new_P1_R584_U7 = ~new_P1_U2677;
  assign new_P1_R584_U8 = ~new_P1_U2674;
  assign new_P1_R584_U9 = ~new_P1_U2675;
  assign new_P1_R2099_U4 = ~new_P1_U4190;
  assign new_P1_R2099_U5 = ~new_P1_U4189;
  assign new_P1_R2099_U6 = ~new_P1_U2678;
  assign new_P1_R2099_U7 = ~new_P1_R2099_U88 | ~new_P1_R2099_U137;
  assign new_P1_R2099_U8 = ~new_P1_R2099_U89 | ~new_P1_R2099_U155;
  assign new_P1_R2099_U9 = ~new_P1_R2099_U90 | ~new_P1_R2099_U157;
  assign new_P1_R2099_U10 = ~new_P1_R2099_U91 | ~new_P1_R2099_U159;
  assign new_P1_R2099_U11 = ~new_P1_R2099_U92 | ~new_P1_R2099_U161;
  assign new_P1_R2099_U12 = ~new_P1_R2099_U93 | ~new_P1_R2099_U163;
  assign new_P1_R2099_U13 = ~new_P1_R2099_U94 | ~new_P1_R2099_U165;
  assign new_P1_R2099_U14 = ~new_P1_R2099_U95 | ~new_P1_R2099_U167;
  assign new_P1_R2099_U15 = ~new_P1_R2099_U169 | ~new_P1_R2099_U55;
  assign new_P1_R2099_U16 = ~new_P1_R2099_U170 | ~new_P1_R2099_U54;
  assign new_P1_R2099_U17 = ~new_P1_R2099_U171 | ~new_P1_R2099_U53;
  assign new_P1_R2099_U18 = ~new_P1_R2099_U172 | ~new_P1_R2099_U52;
  assign new_P1_R2099_U19 = ~new_P1_R2099_U173 | ~new_P1_R2099_U51;
  assign new_P1_R2099_U20 = ~new_P1_R2099_U174 | ~new_P1_R2099_U50;
  assign new_P1_R2099_U21 = ~new_P1_R2099_U175 | ~new_P1_R2099_U49;
  assign new_P1_R2099_U22 = ~new_P1_R2099_U176 | ~new_P1_R2099_U48;
  assign new_P1_R2099_U23 = ~new_P1_R2099_U177 | ~new_P1_R2099_U47;
  assign new_P1_R2099_U24 = ~new_P1_R2099_U178 | ~new_P1_R2099_U46;
  assign new_P1_R2099_U25 = ~new_P1_R2099_U179 | ~new_P1_R2099_U45;
  assign new_P1_R2099_U26 = ~new_P1_R2099_U210 | ~new_P1_R2099_U209;
  assign new_P1_R2099_U27 = ~new_P1_R2099_U183 | ~new_P1_R2099_U182;
  assign new_P1_R2099_U28 = ~new_P1_R2099_U204 | ~new_P1_R2099_U203;
  assign new_P1_R2099_U29 = ~new_P1_R2099_U207 | ~new_P1_R2099_U206;
  assign new_P1_R2099_U30 = ~new_P1_R2099_U198 | ~new_P1_R2099_U197;
  assign new_P1_R2099_U31 = ~new_P1_R2099_U201 | ~new_P1_R2099_U200;
  assign new_P1_R2099_U32 = ~new_P1_R2099_U186 | ~new_P1_R2099_U185;
  assign new_P1_R2099_U33 = ~new_P1_R2099_U189 | ~new_P1_R2099_U188;
  assign new_P1_R2099_U34 = ~new_P1_R2099_U195 | ~new_P1_R2099_U194;
  assign new_P1_R2099_U35 = ~new_P1_R2099_U192 | ~new_P1_R2099_U191;
  assign new_P1_R2099_U36 = ~new_P1_R2099_U213 | ~new_P1_R2099_U212;
  assign new_P1_R2099_U37 = ~new_P1_R2099_U215 | ~new_P1_R2099_U214;
  assign new_P1_R2099_U38 = ~new_P1_R2099_U217 | ~new_P1_R2099_U216;
  assign new_P1_R2099_U39 = ~new_P1_R2099_U219 | ~new_P1_R2099_U218;
  assign new_P1_R2099_U40 = ~new_P1_R2099_U221 | ~new_P1_R2099_U220;
  assign new_P1_R2099_U41 = ~new_P1_R2099_U223 | ~new_P1_R2099_U222;
  assign new_P1_R2099_U42 = ~new_P1_R2099_U225 | ~new_P1_R2099_U224;
  assign new_P1_R2099_U43 = ~new_P1_R2099_U284 | ~new_P1_R2099_U283;
  assign new_P1_R2099_U44 = ~new_P1_R2099_U287 | ~new_P1_R2099_U286;
  assign new_P1_R2099_U45 = ~new_P1_R2099_U227 | ~new_P1_R2099_U226;
  assign new_P1_R2099_U46 = ~new_P1_R2099_U230 | ~new_P1_R2099_U229;
  assign new_P1_R2099_U47 = ~new_P1_R2099_U233 | ~new_P1_R2099_U232;
  assign new_P1_R2099_U48 = ~new_P1_R2099_U236 | ~new_P1_R2099_U235;
  assign new_P1_R2099_U49 = ~new_P1_R2099_U239 | ~new_P1_R2099_U238;
  assign new_P1_R2099_U50 = ~new_P1_R2099_U242 | ~new_P1_R2099_U241;
  assign new_P1_R2099_U51 = ~new_P1_R2099_U245 | ~new_P1_R2099_U244;
  assign new_P1_R2099_U52 = ~new_P1_R2099_U248 | ~new_P1_R2099_U247;
  assign new_P1_R2099_U53 = ~new_P1_R2099_U251 | ~new_P1_R2099_U250;
  assign new_P1_R2099_U54 = ~new_P1_R2099_U254 | ~new_P1_R2099_U253;
  assign new_P1_R2099_U55 = ~new_P1_R2099_U257 | ~new_P1_R2099_U256;
  assign new_P1_R2099_U56 = ~new_P1_R2099_U278 | ~new_P1_R2099_U277;
  assign new_P1_R2099_U57 = ~new_P1_R2099_U281 | ~new_P1_R2099_U280;
  assign new_P1_R2099_U58 = ~new_P1_R2099_U272 | ~new_P1_R2099_U271;
  assign new_P1_R2099_U59 = ~new_P1_R2099_U275 | ~new_P1_R2099_U274;
  assign new_P1_R2099_U60 = ~new_P1_R2099_U266 | ~new_P1_R2099_U265;
  assign new_P1_R2099_U61 = ~new_P1_R2099_U269 | ~new_P1_R2099_U268;
  assign new_P1_R2099_U62 = ~new_P1_R2099_U260 | ~new_P1_R2099_U259;
  assign new_P1_R2099_U63 = ~new_P1_R2099_U263 | ~new_P1_R2099_U262;
  assign new_P1_R2099_U64 = ~new_P1_R2099_U293 | ~new_P1_R2099_U292;
  assign new_P1_R2099_U65 = ~new_P1_R2099_U295 | ~new_P1_R2099_U294;
  assign new_P1_R2099_U66 = ~new_P1_R2099_U299 | ~new_P1_R2099_U298;
  assign new_P1_R2099_U67 = ~new_P1_R2099_U301 | ~new_P1_R2099_U300;
  assign new_P1_R2099_U68 = ~new_P1_R2099_U303 | ~new_P1_R2099_U302;
  assign new_P1_R2099_U69 = ~new_P1_R2099_U305 | ~new_P1_R2099_U304;
  assign new_P1_R2099_U70 = ~new_P1_R2099_U307 | ~new_P1_R2099_U306;
  assign new_P1_R2099_U71 = ~new_P1_R2099_U309 | ~new_P1_R2099_U308;
  assign new_P1_R2099_U72 = ~new_P1_R2099_U311 | ~new_P1_R2099_U310;
  assign new_P1_R2099_U73 = ~new_P1_R2099_U313 | ~new_P1_R2099_U312;
  assign new_P1_R2099_U74 = ~new_P1_R2099_U315 | ~new_P1_R2099_U314;
  assign new_P1_R2099_U75 = ~new_P1_R2099_U317 | ~new_P1_R2099_U316;
  assign new_P1_R2099_U76 = ~new_P1_R2099_U326 | ~new_P1_R2099_U325;
  assign new_P1_R2099_U77 = ~new_P1_R2099_U328 | ~new_P1_R2099_U327;
  assign new_P1_R2099_U78 = ~new_P1_R2099_U330 | ~new_P1_R2099_U329;
  assign new_P1_R2099_U79 = ~new_P1_R2099_U332 | ~new_P1_R2099_U331;
  assign new_P1_R2099_U80 = ~new_P1_R2099_U334 | ~new_P1_R2099_U333;
  assign new_P1_R2099_U81 = ~new_P1_R2099_U336 | ~new_P1_R2099_U335;
  assign new_P1_R2099_U82 = ~new_P1_R2099_U338 | ~new_P1_R2099_U337;
  assign new_P1_R2099_U83 = ~new_P1_R2099_U340 | ~new_P1_R2099_U339;
  assign new_P1_R2099_U84 = ~new_P1_R2099_U342 | ~new_P1_R2099_U341;
  assign new_P1_R2099_U85 = ~new_P1_R2099_U344 | ~new_P1_R2099_U343;
  assign new_P1_R2099_U86 = ~new_P1_R2099_U349 | ~new_P1_R2099_U348;
  assign new_P1_R2099_U87 = ~new_P1_R2099_U324 | ~new_P1_R2099_U323;
  assign new_P1_R2099_U88 = new_P1_R2099_U34 & new_P1_R2099_U35;
  assign new_P1_R2099_U89 = new_P1_R2099_U31 & new_P1_R2099_U30;
  assign new_P1_R2099_U90 = new_P1_R2099_U29 & new_P1_R2099_U28;
  assign new_P1_R2099_U91 = new_P1_R2099_U26 & new_P1_R2099_U27;
  assign new_P1_R2099_U92 = new_P1_R2099_U63 & new_P1_R2099_U62;
  assign new_P1_R2099_U93 = new_P1_R2099_U61 & new_P1_R2099_U60;
  assign new_P1_R2099_U94 = new_P1_R2099_U59 & new_P1_R2099_U58;
  assign new_P1_R2099_U95 = new_P1_R2099_U57 & new_P1_R2099_U56;
  assign new_P1_R2099_U96 = new_P1_R2099_U44 & new_P1_R2099_U43;
  assign new_P1_R2099_U97 = ~new_P1_R2099_U290 | ~new_P1_R2099_U289;
  assign new_P1_R2099_U98 = ~new_P1_R2099_U346 | ~new_P1_R2099_U345;
  assign new_P1_R2099_U99 = ~new_P1_U2702;
  assign new_P1_R2099_U100 = ~new_P1_U2710;
  assign new_P1_R2099_U101 = ~new_P1_U2709;
  assign new_P1_R2099_U102 = ~new_P1_U2708;
  assign new_P1_R2099_U103 = ~new_P1_U2707;
  assign new_P1_R2099_U104 = ~new_P1_U2706;
  assign new_P1_R2099_U105 = ~new_P1_U2705;
  assign new_P1_R2099_U106 = ~new_P1_U2704;
  assign new_P1_R2099_U107 = ~new_P1_U2703;
  assign new_P1_R2099_U108 = ~new_P1_U2701;
  assign new_P1_R2099_U109 = ~new_P1_R2099_U159 | ~new_P1_R2099_U27;
  assign new_P1_R2099_U110 = ~new_P1_R2099_U157 | ~new_P1_R2099_U28;
  assign new_P1_R2099_U111 = ~new_P1_R2099_U155 | ~new_P1_R2099_U30;
  assign new_P1_R2099_U112 = ~new_P1_R2099_U35 | ~new_P1_R2099_U137;
  assign new_P1_R2099_U113 = ~new_P1_U2682;
  assign new_P1_R2099_U114 = ~new_P1_U2683;
  assign new_P1_R2099_U115 = ~new_P1_U2684;
  assign new_P1_R2099_U116 = ~new_P1_U2685;
  assign new_P1_R2099_U117 = ~new_P1_U2686;
  assign new_P1_R2099_U118 = ~new_P1_U2687;
  assign new_P1_R2099_U119 = ~new_P1_U2688;
  assign new_P1_R2099_U120 = ~new_P1_U2689;
  assign new_P1_R2099_U121 = ~new_P1_U2690;
  assign new_P1_R2099_U122 = ~new_P1_U2691;
  assign new_P1_R2099_U123 = ~new_P1_U2692;
  assign new_P1_R2099_U124 = ~new_P1_U2700;
  assign new_P1_R2099_U125 = ~new_P1_U2699;
  assign new_P1_R2099_U126 = ~new_P1_U2698;
  assign new_P1_R2099_U127 = ~new_P1_U2697;
  assign new_P1_R2099_U128 = ~new_P1_U2696;
  assign new_P1_R2099_U129 = ~new_P1_U2695;
  assign new_P1_R2099_U130 = ~new_P1_U2694;
  assign new_P1_R2099_U131 = ~new_P1_U2693;
  assign new_P1_R2099_U132 = ~new_P1_U2680;
  assign new_P1_R2099_U133 = ~new_P1_U2681;
  assign new_P1_R2099_U134 = ~new_P1_U2679;
  assign new_P1_R2099_U135 = ~new_P1_R2099_U96 | ~new_P1_R2099_U180;
  assign new_P1_R2099_U136 = ~new_P1_R2099_U180 | ~new_P1_R2099_U44;
  assign new_P1_R2099_U137 = ~new_P1_R2099_U152 | ~new_P1_R2099_U151;
  assign new_P1_R2099_U138 = new_P1_R2099_U297 & new_P1_R2099_U296;
  assign new_P1_R2099_U139 = new_P1_R2099_U319 & new_P1_R2099_U318;
  assign new_P1_R2099_U140 = ~new_P1_R2099_U148 | ~new_P1_R2099_U147;
  assign new_P1_R2099_U141 = ~new_P1_R2099_U167 | ~new_P1_R2099_U56;
  assign new_P1_R2099_U142 = ~new_P1_R2099_U165 | ~new_P1_R2099_U58;
  assign new_P1_R2099_U143 = ~new_P1_R2099_U163 | ~new_P1_R2099_U60;
  assign new_P1_R2099_U144 = ~new_P1_R2099_U161 | ~new_P1_R2099_U62;
  assign new_P1_R2099_U145 = ~new_P1_R2099_U135;
  assign new_P1_R2099_U146 = new_P1_U4190 | new_P1_U4189;
  assign new_P1_R2099_U147 = ~new_P1_R2099_U32 | ~new_P1_R2099_U146;
  assign new_P1_R2099_U148 = ~new_P1_U4189 | ~new_P1_U4190;
  assign new_P1_R2099_U149 = ~new_P1_R2099_U140;
  assign new_P1_R2099_U150 = ~new_P1_R2099_U190 | ~new_P1_R2099_U6;
  assign new_P1_R2099_U151 = ~new_P1_R2099_U150 | ~new_P1_R2099_U140;
  assign new_P1_R2099_U152 = ~new_P1_U2678 | ~new_P1_R2099_U33;
  assign new_P1_R2099_U153 = ~new_P1_R2099_U137;
  assign new_P1_R2099_U154 = ~new_P1_R2099_U112;
  assign new_P1_R2099_U155 = ~new_P1_R2099_U7;
  assign new_P1_R2099_U156 = ~new_P1_R2099_U111;
  assign new_P1_R2099_U157 = ~new_P1_R2099_U8;
  assign new_P1_R2099_U158 = ~new_P1_R2099_U110;
  assign new_P1_R2099_U159 = ~new_P1_R2099_U9;
  assign new_P1_R2099_U160 = ~new_P1_R2099_U109;
  assign new_P1_R2099_U161 = ~new_P1_R2099_U10;
  assign new_P1_R2099_U162 = ~new_P1_R2099_U144;
  assign new_P1_R2099_U163 = ~new_P1_R2099_U11;
  assign new_P1_R2099_U164 = ~new_P1_R2099_U143;
  assign new_P1_R2099_U165 = ~new_P1_R2099_U12;
  assign new_P1_R2099_U166 = ~new_P1_R2099_U142;
  assign new_P1_R2099_U167 = ~new_P1_R2099_U13;
  assign new_P1_R2099_U168 = ~new_P1_R2099_U141;
  assign new_P1_R2099_U169 = ~new_P1_R2099_U14;
  assign new_P1_R2099_U170 = ~new_P1_R2099_U15;
  assign new_P1_R2099_U171 = ~new_P1_R2099_U16;
  assign new_P1_R2099_U172 = ~new_P1_R2099_U17;
  assign new_P1_R2099_U173 = ~new_P1_R2099_U18;
  assign new_P1_R2099_U174 = ~new_P1_R2099_U19;
  assign new_P1_R2099_U175 = ~new_P1_R2099_U20;
  assign new_P1_R2099_U176 = ~new_P1_R2099_U21;
  assign new_P1_R2099_U177 = ~new_P1_R2099_U22;
  assign new_P1_R2099_U178 = ~new_P1_R2099_U23;
  assign new_P1_R2099_U179 = ~new_P1_R2099_U24;
  assign new_P1_R2099_U180 = ~new_P1_R2099_U25;
  assign new_P1_R2099_U181 = ~new_P1_R2099_U136;
  assign new_P1_R2099_U182 = ~new_P1_U4190 | ~new_P1_R2099_U99;
  assign new_P1_R2099_U183 = ~new_P1_U2702 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U184 = ~new_P1_R2099_U27;
  assign new_P1_R2099_U185 = ~new_P1_U4190 | ~new_P1_R2099_U100;
  assign new_P1_R2099_U186 = ~new_P1_U2710 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U187 = ~new_P1_R2099_U32;
  assign new_P1_R2099_U188 = ~new_P1_U4190 | ~new_P1_R2099_U101;
  assign new_P1_R2099_U189 = ~new_P1_U2709 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U190 = ~new_P1_R2099_U33;
  assign new_P1_R2099_U191 = ~new_P1_U4190 | ~new_P1_R2099_U102;
  assign new_P1_R2099_U192 = ~new_P1_U2708 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U193 = ~new_P1_R2099_U35;
  assign new_P1_R2099_U194 = ~new_P1_U4190 | ~new_P1_R2099_U103;
  assign new_P1_R2099_U195 = ~new_P1_U2707 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U196 = ~new_P1_R2099_U34;
  assign new_P1_R2099_U197 = ~new_P1_U4190 | ~new_P1_R2099_U104;
  assign new_P1_R2099_U198 = ~new_P1_U2706 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U199 = ~new_P1_R2099_U30;
  assign new_P1_R2099_U200 = ~new_P1_U4190 | ~new_P1_R2099_U105;
  assign new_P1_R2099_U201 = ~new_P1_U2705 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U202 = ~new_P1_R2099_U31;
  assign new_P1_R2099_U203 = ~new_P1_U4190 | ~new_P1_R2099_U106;
  assign new_P1_R2099_U204 = ~new_P1_U2704 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U205 = ~new_P1_R2099_U28;
  assign new_P1_R2099_U206 = ~new_P1_U4190 | ~new_P1_R2099_U107;
  assign new_P1_R2099_U207 = ~new_P1_U2703 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U208 = ~new_P1_R2099_U29;
  assign new_P1_R2099_U209 = ~new_P1_U4190 | ~new_P1_R2099_U108;
  assign new_P1_R2099_U210 = ~new_P1_U2701 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U211 = ~new_P1_R2099_U26;
  assign new_P1_R2099_U212 = ~new_P1_R2099_U160 | ~new_P1_R2099_U211;
  assign new_P1_R2099_U213 = ~new_P1_R2099_U26 | ~new_P1_R2099_U109;
  assign new_P1_R2099_U214 = ~new_P1_R2099_U184 | ~new_P1_R2099_U159;
  assign new_P1_R2099_U215 = ~new_P1_R2099_U27 | ~new_P1_R2099_U9;
  assign new_P1_R2099_U216 = ~new_P1_R2099_U158 | ~new_P1_R2099_U208;
  assign new_P1_R2099_U217 = ~new_P1_R2099_U29 | ~new_P1_R2099_U110;
  assign new_P1_R2099_U218 = ~new_P1_R2099_U205 | ~new_P1_R2099_U157;
  assign new_P1_R2099_U219 = ~new_P1_R2099_U28 | ~new_P1_R2099_U8;
  assign new_P1_R2099_U220 = ~new_P1_R2099_U156 | ~new_P1_R2099_U202;
  assign new_P1_R2099_U221 = ~new_P1_R2099_U31 | ~new_P1_R2099_U111;
  assign new_P1_R2099_U222 = ~new_P1_R2099_U199 | ~new_P1_R2099_U155;
  assign new_P1_R2099_U223 = ~new_P1_R2099_U30 | ~new_P1_R2099_U7;
  assign new_P1_R2099_U224 = ~new_P1_R2099_U154 | ~new_P1_R2099_U196;
  assign new_P1_R2099_U225 = ~new_P1_R2099_U34 | ~new_P1_R2099_U112;
  assign new_P1_R2099_U226 = ~new_P1_U4190 | ~new_P1_R2099_U113;
  assign new_P1_R2099_U227 = ~new_P1_U2682 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U228 = ~new_P1_R2099_U45;
  assign new_P1_R2099_U229 = ~new_P1_U4190 | ~new_P1_R2099_U114;
  assign new_P1_R2099_U230 = ~new_P1_U2683 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U231 = ~new_P1_R2099_U46;
  assign new_P1_R2099_U232 = ~new_P1_U4190 | ~new_P1_R2099_U115;
  assign new_P1_R2099_U233 = ~new_P1_U2684 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U234 = ~new_P1_R2099_U47;
  assign new_P1_R2099_U235 = ~new_P1_U4190 | ~new_P1_R2099_U116;
  assign new_P1_R2099_U236 = ~new_P1_U2685 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U237 = ~new_P1_R2099_U48;
  assign new_P1_R2099_U238 = ~new_P1_U4190 | ~new_P1_R2099_U117;
  assign new_P1_R2099_U239 = ~new_P1_U2686 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U240 = ~new_P1_R2099_U49;
  assign new_P1_R2099_U241 = ~new_P1_U4190 | ~new_P1_R2099_U118;
  assign new_P1_R2099_U242 = ~new_P1_U2687 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U243 = ~new_P1_R2099_U50;
  assign new_P1_R2099_U244 = ~new_P1_U4190 | ~new_P1_R2099_U119;
  assign new_P1_R2099_U245 = ~new_P1_U2688 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U246 = ~new_P1_R2099_U51;
  assign new_P1_R2099_U247 = ~new_P1_U4190 | ~new_P1_R2099_U120;
  assign new_P1_R2099_U248 = ~new_P1_U2689 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U249 = ~new_P1_R2099_U52;
  assign new_P1_R2099_U250 = ~new_P1_U4190 | ~new_P1_R2099_U121;
  assign new_P1_R2099_U251 = ~new_P1_U2690 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U252 = ~new_P1_R2099_U53;
  assign new_P1_R2099_U253 = ~new_P1_U4190 | ~new_P1_R2099_U122;
  assign new_P1_R2099_U254 = ~new_P1_U2691 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U255 = ~new_P1_R2099_U54;
  assign new_P1_R2099_U256 = ~new_P1_U4190 | ~new_P1_R2099_U123;
  assign new_P1_R2099_U257 = ~new_P1_U2692 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U258 = ~new_P1_R2099_U55;
  assign new_P1_R2099_U259 = ~new_P1_U4190 | ~new_P1_R2099_U124;
  assign new_P1_R2099_U260 = ~new_P1_U2700 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U261 = ~new_P1_R2099_U62;
  assign new_P1_R2099_U262 = ~new_P1_U4190 | ~new_P1_R2099_U125;
  assign new_P1_R2099_U263 = ~new_P1_U2699 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U264 = ~new_P1_R2099_U63;
  assign new_P1_R2099_U265 = ~new_P1_U4190 | ~new_P1_R2099_U126;
  assign new_P1_R2099_U266 = ~new_P1_U2698 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U267 = ~new_P1_R2099_U60;
  assign new_P1_R2099_U268 = ~new_P1_U4190 | ~new_P1_R2099_U127;
  assign new_P1_R2099_U269 = ~new_P1_U2697 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U270 = ~new_P1_R2099_U61;
  assign new_P1_R2099_U271 = ~new_P1_U4190 | ~new_P1_R2099_U128;
  assign new_P1_R2099_U272 = ~new_P1_U2696 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U273 = ~new_P1_R2099_U58;
  assign new_P1_R2099_U274 = ~new_P1_U4190 | ~new_P1_R2099_U129;
  assign new_P1_R2099_U275 = ~new_P1_U2695 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U276 = ~new_P1_R2099_U59;
  assign new_P1_R2099_U277 = ~new_P1_U4190 | ~new_P1_R2099_U130;
  assign new_P1_R2099_U278 = ~new_P1_U2694 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U279 = ~new_P1_R2099_U56;
  assign new_P1_R2099_U280 = ~new_P1_U4190 | ~new_P1_R2099_U131;
  assign new_P1_R2099_U281 = ~new_P1_U2693 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U282 = ~new_P1_R2099_U57;
  assign new_P1_R2099_U283 = ~new_P1_U4190 | ~new_P1_R2099_U132;
  assign new_P1_R2099_U284 = ~new_P1_U2680 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U285 = ~new_P1_R2099_U43;
  assign new_P1_R2099_U286 = ~new_P1_U4190 | ~new_P1_R2099_U133;
  assign new_P1_R2099_U287 = ~new_P1_U2681 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U288 = ~new_P1_R2099_U44;
  assign new_P1_R2099_U289 = ~new_P1_U4190 | ~new_P1_R2099_U134;
  assign new_P1_R2099_U290 = ~new_P1_U2679 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U291 = ~new_P1_R2099_U97;
  assign new_P1_R2099_U292 = ~new_P1_R2099_U145 | ~new_P1_R2099_U291;
  assign new_P1_R2099_U293 = ~new_P1_R2099_U97 | ~new_P1_R2099_U135;
  assign new_P1_R2099_U294 = ~new_P1_R2099_U181 | ~new_P1_R2099_U285;
  assign new_P1_R2099_U295 = ~new_P1_R2099_U43 | ~new_P1_R2099_U136;
  assign new_P1_R2099_U296 = ~new_P1_R2099_U153 | ~new_P1_R2099_U193;
  assign new_P1_R2099_U297 = ~new_P1_R2099_U35 | ~new_P1_R2099_U137;
  assign new_P1_R2099_U298 = ~new_P1_R2099_U288 | ~new_P1_R2099_U180;
  assign new_P1_R2099_U299 = ~new_P1_R2099_U44 | ~new_P1_R2099_U25;
  assign new_P1_R2099_U300 = ~new_P1_R2099_U228 | ~new_P1_R2099_U179;
  assign new_P1_R2099_U301 = ~new_P1_R2099_U45 | ~new_P1_R2099_U24;
  assign new_P1_R2099_U302 = ~new_P1_R2099_U231 | ~new_P1_R2099_U178;
  assign new_P1_R2099_U303 = ~new_P1_R2099_U46 | ~new_P1_R2099_U23;
  assign new_P1_R2099_U304 = ~new_P1_R2099_U234 | ~new_P1_R2099_U177;
  assign new_P1_R2099_U305 = ~new_P1_R2099_U47 | ~new_P1_R2099_U22;
  assign new_P1_R2099_U306 = ~new_P1_R2099_U237 | ~new_P1_R2099_U176;
  assign new_P1_R2099_U307 = ~new_P1_R2099_U48 | ~new_P1_R2099_U21;
  assign new_P1_R2099_U308 = ~new_P1_R2099_U240 | ~new_P1_R2099_U175;
  assign new_P1_R2099_U309 = ~new_P1_R2099_U49 | ~new_P1_R2099_U20;
  assign new_P1_R2099_U310 = ~new_P1_R2099_U243 | ~new_P1_R2099_U174;
  assign new_P1_R2099_U311 = ~new_P1_R2099_U50 | ~new_P1_R2099_U19;
  assign new_P1_R2099_U312 = ~new_P1_R2099_U246 | ~new_P1_R2099_U173;
  assign new_P1_R2099_U313 = ~new_P1_R2099_U51 | ~new_P1_R2099_U18;
  assign new_P1_R2099_U314 = ~new_P1_R2099_U249 | ~new_P1_R2099_U172;
  assign new_P1_R2099_U315 = ~new_P1_R2099_U52 | ~new_P1_R2099_U17;
  assign new_P1_R2099_U316 = ~new_P1_R2099_U252 | ~new_P1_R2099_U171;
  assign new_P1_R2099_U317 = ~new_P1_R2099_U53 | ~new_P1_R2099_U16;
  assign new_P1_R2099_U318 = ~new_P1_R2099_U190 | ~new_P1_U2678;
  assign new_P1_R2099_U319 = ~new_P1_R2099_U33 | ~new_P1_R2099_U6;
  assign new_P1_R2099_U320 = ~new_P1_R2099_U190 | ~new_P1_U2678;
  assign new_P1_R2099_U321 = ~new_P1_R2099_U33 | ~new_P1_R2099_U6;
  assign new_P1_R2099_U322 = ~new_P1_R2099_U321 | ~new_P1_R2099_U320;
  assign new_P1_R2099_U323 = ~new_P1_R2099_U139 | ~new_P1_R2099_U140;
  assign new_P1_R2099_U324 = ~new_P1_R2099_U149 | ~new_P1_R2099_U322;
  assign new_P1_R2099_U325 = ~new_P1_R2099_U255 | ~new_P1_R2099_U170;
  assign new_P1_R2099_U326 = ~new_P1_R2099_U54 | ~new_P1_R2099_U15;
  assign new_P1_R2099_U327 = ~new_P1_R2099_U258 | ~new_P1_R2099_U169;
  assign new_P1_R2099_U328 = ~new_P1_R2099_U55 | ~new_P1_R2099_U14;
  assign new_P1_R2099_U329 = ~new_P1_R2099_U168 | ~new_P1_R2099_U282;
  assign new_P1_R2099_U330 = ~new_P1_R2099_U57 | ~new_P1_R2099_U141;
  assign new_P1_R2099_U331 = ~new_P1_R2099_U279 | ~new_P1_R2099_U167;
  assign new_P1_R2099_U332 = ~new_P1_R2099_U56 | ~new_P1_R2099_U13;
  assign new_P1_R2099_U333 = ~new_P1_R2099_U166 | ~new_P1_R2099_U276;
  assign new_P1_R2099_U334 = ~new_P1_R2099_U59 | ~new_P1_R2099_U142;
  assign new_P1_R2099_U335 = ~new_P1_R2099_U273 | ~new_P1_R2099_U165;
  assign new_P1_R2099_U336 = ~new_P1_R2099_U58 | ~new_P1_R2099_U12;
  assign new_P1_R2099_U337 = ~new_P1_R2099_U164 | ~new_P1_R2099_U270;
  assign new_P1_R2099_U338 = ~new_P1_R2099_U61 | ~new_P1_R2099_U143;
  assign new_P1_R2099_U339 = ~new_P1_R2099_U267 | ~new_P1_R2099_U163;
  assign new_P1_R2099_U340 = ~new_P1_R2099_U60 | ~new_P1_R2099_U11;
  assign new_P1_R2099_U341 = ~new_P1_R2099_U162 | ~new_P1_R2099_U264;
  assign new_P1_R2099_U342 = ~new_P1_R2099_U63 | ~new_P1_R2099_U144;
  assign new_P1_R2099_U343 = ~new_P1_R2099_U261 | ~new_P1_R2099_U161;
  assign new_P1_R2099_U344 = ~new_P1_R2099_U62 | ~new_P1_R2099_U10;
  assign new_P1_R2099_U345 = ~new_P1_U4189 | ~new_P1_R2099_U4;
  assign new_P1_R2099_U346 = ~new_P1_U4190 | ~new_P1_R2099_U5;
  assign new_P1_R2099_U347 = ~new_P1_R2099_U98;
  assign new_P1_R2099_U348 = ~new_P1_R2099_U32 | ~new_P1_R2099_U347;
  assign new_P1_R2099_U349 = ~new_P1_R2099_U98 | ~new_P1_R2099_U187;
  assign new_P1_R2167_U6 = ~new_P1_U2716;
  assign new_P1_R2167_U7 = ~new_P1_U2714;
  assign new_P1_R2167_U8 = ~new_P1_U2720;
  assign new_P1_R2167_U9 = ~new_P1_U2719;
  assign new_P1_R2167_U10 = ~new_P1_U2713;
  assign new_P1_R2167_U11 = ~new_P1_U2712;
  assign new_P1_R2167_U12 = ~new_P1_U2718;
  assign new_P1_R2167_U13 = ~new_P1_U2717;
  assign new_P1_R2167_U14 = ~new_P1_U2711;
  assign new_P1_R2167_U15 = ~new_P1_U2356;
  assign new_P1_R2167_U16 = ~P1_STATE2_REG_0_;
  assign new_P1_R2167_U17 = ~new_P1_R2167_U50 | ~new_P1_R2167_U49;
  assign new_P1_R2167_U18 = new_P1_R2167_U29 & new_P1_R2167_U30;
  assign new_P1_R2167_U19 = new_P1_R2167_U32 & new_P1_R2167_U33;
  assign new_P1_R2167_U20 = new_P1_R2167_U35 & new_P1_R2167_U36;
  assign new_P1_R2167_U21 = new_P1_R2167_U38 & new_P1_R2167_U39;
  assign new_P1_R2167_U22 = ~new_P1_U2721;
  assign new_P1_R2167_U23 = ~new_P1_U2722;
  assign new_P1_R2167_U24 = ~new_P1_U2715 | ~new_P1_R2167_U23;
  assign new_P1_R2167_U25 = ~new_P1_U2715 | ~new_P1_R2167_U22;
  assign new_P1_R2167_U26 = new_P1_U2721 | new_P1_U2722;
  assign new_P1_R2167_U27 = ~new_P1_U2714 | ~new_P1_R2167_U8;
  assign new_P1_R2167_U28 = ~new_P1_R2167_U24 | ~new_P1_R2167_U25 | ~new_P1_R2167_U27 | ~new_P1_R2167_U26;
  assign new_P1_R2167_U29 = ~new_P1_U2720 | ~new_P1_R2167_U7;
  assign new_P1_R2167_U30 = ~new_P1_U2719 | ~new_P1_R2167_U10;
  assign new_P1_R2167_U31 = ~new_P1_R2167_U18 | ~new_P1_R2167_U28;
  assign new_P1_R2167_U32 = ~new_P1_U2713 | ~new_P1_R2167_U9;
  assign new_P1_R2167_U33 = ~new_P1_U2712 | ~new_P1_R2167_U12;
  assign new_P1_R2167_U34 = ~new_P1_R2167_U19 | ~new_P1_R2167_U31;
  assign new_P1_R2167_U35 = ~new_P1_U2718 | ~new_P1_R2167_U11;
  assign new_P1_R2167_U36 = ~new_P1_U2717 | ~new_P1_R2167_U14;
  assign new_P1_R2167_U37 = ~new_P1_R2167_U20 | ~new_P1_R2167_U34;
  assign new_P1_R2167_U38 = ~new_P1_U2711 | ~new_P1_R2167_U13;
  assign new_P1_R2167_U39 = ~new_P1_U2356 | ~new_P1_R2167_U6;
  assign new_P1_R2167_U40 = ~new_P1_R2167_U21 | ~new_P1_R2167_U37;
  assign new_P1_R2167_U41 = ~new_P1_U2716 | ~new_P1_R2167_U15;
  assign new_P1_R2167_U42 = ~new_P1_R2167_U40 | ~new_P1_R2167_U41;
  assign new_P1_R2167_U43 = ~new_P1_U2716 | ~new_P1_R2167_U16;
  assign new_P1_R2167_U44 = ~new_P1_R2167_U42 | ~new_P1_R2167_U6;
  assign new_P1_R2167_U45 = ~new_P1_R2167_U44 | ~new_P1_R2167_U43;
  assign new_P1_R2167_U46 = ~P1_STATE2_REG_0_ | ~new_P1_R2167_U6;
  assign new_P1_R2167_U47 = ~new_P1_U2716 | ~new_P1_R2167_U42;
  assign new_P1_R2167_U48 = ~new_P1_R2167_U47 | ~new_P1_R2167_U46;
  assign new_P1_R2167_U49 = ~new_P1_R2167_U45 | ~new_P1_R2167_U15;
  assign new_P1_R2167_U50 = ~new_P1_U2356 | ~new_P1_R2167_U48;
  assign new_P1_R2337_U4 = ~P1_PHYADDRPOINTER_REG_1_;
  assign new_P1_R2337_U5 = ~P1_PHYADDRPOINTER_REG_2_;
  assign new_P1_R2337_U6 = ~P1_PHYADDRPOINTER_REG_2_ | ~P1_PHYADDRPOINTER_REG_1_;
  assign new_P1_R2337_U7 = ~P1_PHYADDRPOINTER_REG_3_;
  assign new_P1_R2337_U8 = ~P1_PHYADDRPOINTER_REG_3_ | ~new_P1_R2337_U94;
  assign new_P1_R2337_U9 = ~P1_PHYADDRPOINTER_REG_4_;
  assign new_P1_R2337_U10 = ~P1_PHYADDRPOINTER_REG_4_ | ~new_P1_R2337_U95;
  assign new_P1_R2337_U11 = ~P1_PHYADDRPOINTER_REG_5_;
  assign new_P1_R2337_U12 = ~P1_PHYADDRPOINTER_REG_5_ | ~new_P1_R2337_U96;
  assign new_P1_R2337_U13 = ~P1_PHYADDRPOINTER_REG_6_;
  assign new_P1_R2337_U14 = ~P1_PHYADDRPOINTER_REG_6_ | ~new_P1_R2337_U97;
  assign new_P1_R2337_U15 = ~P1_PHYADDRPOINTER_REG_7_;
  assign new_P1_R2337_U16 = ~P1_PHYADDRPOINTER_REG_7_ | ~new_P1_R2337_U98;
  assign new_P1_R2337_U17 = ~P1_PHYADDRPOINTER_REG_8_;
  assign new_P1_R2337_U18 = ~P1_PHYADDRPOINTER_REG_9_;
  assign new_P1_R2337_U19 = ~P1_PHYADDRPOINTER_REG_8_ | ~new_P1_R2337_U99;
  assign new_P1_R2337_U20 = ~new_P1_R2337_U100 | ~P1_PHYADDRPOINTER_REG_9_;
  assign new_P1_R2337_U21 = ~P1_PHYADDRPOINTER_REG_10_;
  assign new_P1_R2337_U22 = ~P1_PHYADDRPOINTER_REG_10_ | ~new_P1_R2337_U101;
  assign new_P1_R2337_U23 = ~P1_PHYADDRPOINTER_REG_11_;
  assign new_P1_R2337_U24 = ~P1_PHYADDRPOINTER_REG_11_ | ~new_P1_R2337_U102;
  assign new_P1_R2337_U25 = ~P1_PHYADDRPOINTER_REG_12_;
  assign new_P1_R2337_U26 = ~P1_PHYADDRPOINTER_REG_12_ | ~new_P1_R2337_U103;
  assign new_P1_R2337_U27 = ~P1_PHYADDRPOINTER_REG_13_;
  assign new_P1_R2337_U28 = ~P1_PHYADDRPOINTER_REG_13_ | ~new_P1_R2337_U104;
  assign new_P1_R2337_U29 = ~P1_PHYADDRPOINTER_REG_14_;
  assign new_P1_R2337_U30 = ~P1_PHYADDRPOINTER_REG_14_ | ~new_P1_R2337_U105;
  assign new_P1_R2337_U31 = ~P1_PHYADDRPOINTER_REG_15_;
  assign new_P1_R2337_U32 = ~P1_PHYADDRPOINTER_REG_15_ | ~new_P1_R2337_U106;
  assign new_P1_R2337_U33 = ~P1_PHYADDRPOINTER_REG_16_;
  assign new_P1_R2337_U34 = ~P1_PHYADDRPOINTER_REG_16_ | ~new_P1_R2337_U107;
  assign new_P1_R2337_U35 = ~P1_PHYADDRPOINTER_REG_17_;
  assign new_P1_R2337_U36 = ~P1_PHYADDRPOINTER_REG_17_ | ~new_P1_R2337_U108;
  assign new_P1_R2337_U37 = ~P1_PHYADDRPOINTER_REG_18_;
  assign new_P1_R2337_U38 = ~P1_PHYADDRPOINTER_REG_18_ | ~new_P1_R2337_U109;
  assign new_P1_R2337_U39 = ~P1_PHYADDRPOINTER_REG_19_;
  assign new_P1_R2337_U40 = ~P1_PHYADDRPOINTER_REG_19_ | ~new_P1_R2337_U110;
  assign new_P1_R2337_U41 = ~P1_PHYADDRPOINTER_REG_20_;
  assign new_P1_R2337_U42 = ~P1_PHYADDRPOINTER_REG_20_ | ~new_P1_R2337_U111;
  assign new_P1_R2337_U43 = ~P1_PHYADDRPOINTER_REG_21_;
  assign new_P1_R2337_U44 = ~P1_PHYADDRPOINTER_REG_21_ | ~new_P1_R2337_U112;
  assign new_P1_R2337_U45 = ~P1_PHYADDRPOINTER_REG_22_;
  assign new_P1_R2337_U46 = ~P1_PHYADDRPOINTER_REG_22_ | ~new_P1_R2337_U113;
  assign new_P1_R2337_U47 = ~P1_PHYADDRPOINTER_REG_23_;
  assign new_P1_R2337_U48 = ~P1_PHYADDRPOINTER_REG_23_ | ~new_P1_R2337_U114;
  assign new_P1_R2337_U49 = ~P1_PHYADDRPOINTER_REG_24_;
  assign new_P1_R2337_U50 = ~P1_PHYADDRPOINTER_REG_24_ | ~new_P1_R2337_U115;
  assign new_P1_R2337_U51 = ~P1_PHYADDRPOINTER_REG_25_;
  assign new_P1_R2337_U52 = ~P1_PHYADDRPOINTER_REG_25_ | ~new_P1_R2337_U116;
  assign new_P1_R2337_U53 = ~P1_PHYADDRPOINTER_REG_26_;
  assign new_P1_R2337_U54 = ~P1_PHYADDRPOINTER_REG_26_ | ~new_P1_R2337_U117;
  assign new_P1_R2337_U55 = ~P1_PHYADDRPOINTER_REG_27_;
  assign new_P1_R2337_U56 = ~P1_PHYADDRPOINTER_REG_27_ | ~new_P1_R2337_U118;
  assign new_P1_R2337_U57 = ~P1_PHYADDRPOINTER_REG_28_;
  assign new_P1_R2337_U58 = ~P1_PHYADDRPOINTER_REG_28_ | ~new_P1_R2337_U119;
  assign new_P1_R2337_U59 = ~P1_PHYADDRPOINTER_REG_29_;
  assign new_P1_R2337_U60 = ~P1_PHYADDRPOINTER_REG_29_ | ~new_P1_R2337_U120;
  assign new_P1_R2337_U61 = ~P1_PHYADDRPOINTER_REG_30_;
  assign new_P1_R2337_U62 = ~new_P1_R2337_U124 | ~new_P1_R2337_U123;
  assign new_P1_R2337_U63 = ~new_P1_R2337_U126 | ~new_P1_R2337_U125;
  assign new_P1_R2337_U64 = ~new_P1_R2337_U128 | ~new_P1_R2337_U127;
  assign new_P1_R2337_U65 = ~new_P1_R2337_U130 | ~new_P1_R2337_U129;
  assign new_P1_R2337_U66 = ~new_P1_R2337_U132 | ~new_P1_R2337_U131;
  assign new_P1_R2337_U67 = ~new_P1_R2337_U134 | ~new_P1_R2337_U133;
  assign new_P1_R2337_U68 = ~new_P1_R2337_U136 | ~new_P1_R2337_U135;
  assign new_P1_R2337_U69 = ~new_P1_R2337_U138 | ~new_P1_R2337_U137;
  assign new_P1_R2337_U70 = ~new_P1_R2337_U140 | ~new_P1_R2337_U139;
  assign new_P1_R2337_U71 = ~new_P1_R2337_U142 | ~new_P1_R2337_U141;
  assign new_P1_R2337_U72 = ~new_P1_R2337_U144 | ~new_P1_R2337_U143;
  assign new_P1_R2337_U73 = ~new_P1_R2337_U146 | ~new_P1_R2337_U145;
  assign new_P1_R2337_U74 = ~new_P1_R2337_U148 | ~new_P1_R2337_U147;
  assign new_P1_R2337_U75 = ~new_P1_R2337_U150 | ~new_P1_R2337_U149;
  assign new_P1_R2337_U76 = ~new_P1_R2337_U152 | ~new_P1_R2337_U151;
  assign new_P1_R2337_U77 = ~new_P1_R2337_U154 | ~new_P1_R2337_U153;
  assign new_P1_R2337_U78 = ~new_P1_R2337_U156 | ~new_P1_R2337_U155;
  assign new_P1_R2337_U79 = ~new_P1_R2337_U158 | ~new_P1_R2337_U157;
  assign new_P1_R2337_U80 = ~new_P1_R2337_U160 | ~new_P1_R2337_U159;
  assign new_P1_R2337_U81 = ~new_P1_R2337_U162 | ~new_P1_R2337_U161;
  assign new_P1_R2337_U82 = ~new_P1_R2337_U164 | ~new_P1_R2337_U163;
  assign new_P1_R2337_U83 = ~new_P1_R2337_U166 | ~new_P1_R2337_U165;
  assign new_P1_R2337_U84 = ~new_P1_R2337_U168 | ~new_P1_R2337_U167;
  assign new_P1_R2337_U85 = ~new_P1_R2337_U170 | ~new_P1_R2337_U169;
  assign new_P1_R2337_U86 = ~new_P1_R2337_U172 | ~new_P1_R2337_U171;
  assign new_P1_R2337_U87 = ~new_P1_R2337_U174 | ~new_P1_R2337_U173;
  assign new_P1_R2337_U88 = ~new_P1_R2337_U176 | ~new_P1_R2337_U175;
  assign new_P1_R2337_U89 = ~new_P1_R2337_U178 | ~new_P1_R2337_U177;
  assign new_P1_R2337_U90 = ~new_P1_R2337_U180 | ~new_P1_R2337_U179;
  assign new_P1_R2337_U91 = ~new_P1_R2337_U182 | ~new_P1_R2337_U181;
  assign new_P1_R2337_U92 = ~P1_PHYADDRPOINTER_REG_31_;
  assign new_P1_R2337_U93 = ~P1_PHYADDRPOINTER_REG_30_ | ~new_P1_R2337_U121;
  assign new_P1_R2337_U94 = ~new_P1_R2337_U6;
  assign new_P1_R2337_U95 = ~new_P1_R2337_U8;
  assign new_P1_R2337_U96 = ~new_P1_R2337_U10;
  assign new_P1_R2337_U97 = ~new_P1_R2337_U12;
  assign new_P1_R2337_U98 = ~new_P1_R2337_U14;
  assign new_P1_R2337_U99 = ~new_P1_R2337_U16;
  assign new_P1_R2337_U100 = ~new_P1_R2337_U19;
  assign new_P1_R2337_U101 = ~new_P1_R2337_U20;
  assign new_P1_R2337_U102 = ~new_P1_R2337_U22;
  assign new_P1_R2337_U103 = ~new_P1_R2337_U24;
  assign new_P1_R2337_U104 = ~new_P1_R2337_U26;
  assign new_P1_R2337_U105 = ~new_P1_R2337_U28;
  assign new_P1_R2337_U106 = ~new_P1_R2337_U30;
  assign new_P1_R2337_U107 = ~new_P1_R2337_U32;
  assign new_P1_R2337_U108 = ~new_P1_R2337_U34;
  assign new_P1_R2337_U109 = ~new_P1_R2337_U36;
  assign new_P1_R2337_U110 = ~new_P1_R2337_U38;
  assign new_P1_R2337_U111 = ~new_P1_R2337_U40;
  assign new_P1_R2337_U112 = ~new_P1_R2337_U42;
  assign new_P1_R2337_U113 = ~new_P1_R2337_U44;
  assign new_P1_R2337_U114 = ~new_P1_R2337_U46;
  assign new_P1_R2337_U115 = ~new_P1_R2337_U48;
  assign new_P1_R2337_U116 = ~new_P1_R2337_U50;
  assign new_P1_R2337_U117 = ~new_P1_R2337_U52;
  assign new_P1_R2337_U118 = ~new_P1_R2337_U54;
  assign new_P1_R2337_U119 = ~new_P1_R2337_U56;
  assign new_P1_R2337_U120 = ~new_P1_R2337_U58;
  assign new_P1_R2337_U121 = ~new_P1_R2337_U60;
  assign new_P1_R2337_U122 = ~new_P1_R2337_U93;
  assign new_P1_R2337_U123 = ~P1_PHYADDRPOINTER_REG_9_ | ~new_P1_R2337_U19;
  assign new_P1_R2337_U124 = ~new_P1_R2337_U100 | ~new_P1_R2337_U18;
  assign new_P1_R2337_U125 = ~P1_PHYADDRPOINTER_REG_8_ | ~new_P1_R2337_U16;
  assign new_P1_R2337_U126 = ~new_P1_R2337_U99 | ~new_P1_R2337_U17;
  assign new_P1_R2337_U127 = ~P1_PHYADDRPOINTER_REG_7_ | ~new_P1_R2337_U14;
  assign new_P1_R2337_U128 = ~new_P1_R2337_U98 | ~new_P1_R2337_U15;
  assign new_P1_R2337_U129 = ~P1_PHYADDRPOINTER_REG_6_ | ~new_P1_R2337_U12;
  assign new_P1_R2337_U130 = ~new_P1_R2337_U97 | ~new_P1_R2337_U13;
  assign new_P1_R2337_U131 = ~P1_PHYADDRPOINTER_REG_5_ | ~new_P1_R2337_U10;
  assign new_P1_R2337_U132 = ~new_P1_R2337_U96 | ~new_P1_R2337_U11;
  assign new_P1_R2337_U133 = ~P1_PHYADDRPOINTER_REG_4_ | ~new_P1_R2337_U8;
  assign new_P1_R2337_U134 = ~new_P1_R2337_U95 | ~new_P1_R2337_U9;
  assign new_P1_R2337_U135 = ~P1_PHYADDRPOINTER_REG_3_ | ~new_P1_R2337_U6;
  assign new_P1_R2337_U136 = ~new_P1_R2337_U94 | ~new_P1_R2337_U7;
  assign new_P1_R2337_U137 = ~P1_PHYADDRPOINTER_REG_31_ | ~new_P1_R2337_U93;
  assign new_P1_R2337_U138 = ~new_P1_R2337_U122 | ~new_P1_R2337_U92;
  assign new_P1_R2337_U139 = ~P1_PHYADDRPOINTER_REG_30_ | ~new_P1_R2337_U60;
  assign new_P1_R2337_U140 = ~new_P1_R2337_U121 | ~new_P1_R2337_U61;
  assign new_P1_R2337_U141 = ~P1_PHYADDRPOINTER_REG_2_ | ~new_P1_R2337_U4;
  assign new_P1_R2337_U142 = ~P1_PHYADDRPOINTER_REG_1_ | ~new_P1_R2337_U5;
  assign new_P1_R2337_U143 = ~P1_PHYADDRPOINTER_REG_29_ | ~new_P1_R2337_U58;
  assign new_P1_R2337_U144 = ~new_P1_R2337_U120 | ~new_P1_R2337_U59;
  assign new_P1_R2337_U145 = ~P1_PHYADDRPOINTER_REG_28_ | ~new_P1_R2337_U56;
  assign new_P1_R2337_U146 = ~new_P1_R2337_U119 | ~new_P1_R2337_U57;
  assign new_P1_R2337_U147 = ~P1_PHYADDRPOINTER_REG_27_ | ~new_P1_R2337_U54;
  assign new_P1_R2337_U148 = ~new_P1_R2337_U118 | ~new_P1_R2337_U55;
  assign new_P1_R2337_U149 = ~P1_PHYADDRPOINTER_REG_26_ | ~new_P1_R2337_U52;
  assign new_P1_R2337_U150 = ~new_P1_R2337_U117 | ~new_P1_R2337_U53;
  assign new_P1_R2337_U151 = ~P1_PHYADDRPOINTER_REG_25_ | ~new_P1_R2337_U50;
  assign new_P1_R2337_U152 = ~new_P1_R2337_U116 | ~new_P1_R2337_U51;
  assign new_P1_R2337_U153 = ~P1_PHYADDRPOINTER_REG_24_ | ~new_P1_R2337_U48;
  assign new_P1_R2337_U154 = ~new_P1_R2337_U115 | ~new_P1_R2337_U49;
  assign new_P1_R2337_U155 = ~P1_PHYADDRPOINTER_REG_23_ | ~new_P1_R2337_U46;
  assign new_P1_R2337_U156 = ~new_P1_R2337_U114 | ~new_P1_R2337_U47;
  assign new_P1_R2337_U157 = ~P1_PHYADDRPOINTER_REG_22_ | ~new_P1_R2337_U44;
  assign new_P1_R2337_U158 = ~new_P1_R2337_U113 | ~new_P1_R2337_U45;
  assign new_P1_R2337_U159 = ~P1_PHYADDRPOINTER_REG_21_ | ~new_P1_R2337_U42;
  assign new_P1_R2337_U160 = ~new_P1_R2337_U112 | ~new_P1_R2337_U43;
  assign new_P1_R2337_U161 = ~P1_PHYADDRPOINTER_REG_20_ | ~new_P1_R2337_U40;
  assign new_P1_R2337_U162 = ~new_P1_R2337_U111 | ~new_P1_R2337_U41;
  assign new_P1_R2337_U163 = ~P1_PHYADDRPOINTER_REG_19_ | ~new_P1_R2337_U38;
  assign new_P1_R2337_U164 = ~new_P1_R2337_U110 | ~new_P1_R2337_U39;
  assign new_P1_R2337_U165 = ~P1_PHYADDRPOINTER_REG_18_ | ~new_P1_R2337_U36;
  assign new_P1_R2337_U166 = ~new_P1_R2337_U109 | ~new_P1_R2337_U37;
  assign new_P1_R2337_U167 = ~P1_PHYADDRPOINTER_REG_17_ | ~new_P1_R2337_U34;
  assign new_P1_R2337_U168 = ~new_P1_R2337_U108 | ~new_P1_R2337_U35;
  assign new_P1_R2337_U169 = ~P1_PHYADDRPOINTER_REG_16_ | ~new_P1_R2337_U32;
  assign new_P1_R2337_U170 = ~new_P1_R2337_U107 | ~new_P1_R2337_U33;
  assign new_P1_R2337_U171 = ~P1_PHYADDRPOINTER_REG_15_ | ~new_P1_R2337_U30;
  assign new_P1_R2337_U172 = ~new_P1_R2337_U106 | ~new_P1_R2337_U31;
  assign new_P1_R2337_U173 = ~P1_PHYADDRPOINTER_REG_14_ | ~new_P1_R2337_U28;
  assign new_P1_R2337_U174 = ~new_P1_R2337_U105 | ~new_P1_R2337_U29;
  assign new_P1_R2337_U175 = ~P1_PHYADDRPOINTER_REG_13_ | ~new_P1_R2337_U26;
  assign new_P1_R2337_U176 = ~new_P1_R2337_U104 | ~new_P1_R2337_U27;
  assign new_P1_R2337_U177 = ~P1_PHYADDRPOINTER_REG_12_ | ~new_P1_R2337_U24;
  assign new_P1_R2337_U178 = ~new_P1_R2337_U103 | ~new_P1_R2337_U25;
  assign new_P1_R2337_U179 = ~P1_PHYADDRPOINTER_REG_11_ | ~new_P1_R2337_U22;
  assign new_P1_R2337_U180 = ~new_P1_R2337_U102 | ~new_P1_R2337_U23;
  assign new_P1_R2337_U181 = ~P1_PHYADDRPOINTER_REG_10_ | ~new_P1_R2337_U20;
  assign new_P1_R2337_U182 = ~new_P1_R2337_U101 | ~new_P1_R2337_U21;
  assign new_P1_SUB_357_U6 = ~new_P1_U3233;
  assign new_P1_SUB_357_U7 = ~new_P1_U3228;
  assign new_P1_SUB_357_U8 = ~new_P1_U3234;
  assign new_P1_SUB_357_U9 = ~new_P1_U3232;
  assign new_P1_SUB_357_U10 = ~new_P1_U3227;
  assign new_P1_SUB_357_U11 = ~new_P1_U3230;
  assign new_P1_SUB_357_U12 = ~new_P1_U3229;
  assign new_P1_SUB_357_U13 = ~new_P1_U3231;
  assign new_P1_LT_563_1260_U6 = new_P1_LT_563_1260_U9 & new_P1_LT_563_1260_U8;
  assign new_P1_LT_563_1260_U7 = ~new_P1_U2673;
  assign new_P1_LT_563_1260_U8 = ~new_P1_R584_U8 | ~new_P1_LT_563_1260_U7;
  assign new_P1_LT_563_1260_U9 = ~new_P1_R584_U9 | ~new_P1_LT_563_1260_U7;
  assign new_P1_SUB_580_U6 = ~new_P1_SUB_580_U10 | ~new_P1_SUB_580_U9;
  assign new_P1_SUB_580_U7 = ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_SUB_580_U8 = ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_SUB_580_U9 = ~P1_INSTADDRPOINTER_REG_1_ | ~new_P1_SUB_580_U8;
  assign new_P1_SUB_580_U10 = ~P1_INSTADDRPOINTER_REG_0_ | ~new_P1_SUB_580_U7;
  assign new_P1_R2096_U4 = ~P1_REIP_REG_1_;
  assign new_P1_R2096_U5 = ~P1_REIP_REG_2_;
  assign new_P1_R2096_U6 = ~P1_REIP_REG_2_ | ~P1_REIP_REG_1_;
  assign new_P1_R2096_U7 = ~P1_REIP_REG_3_;
  assign new_P1_R2096_U8 = ~P1_REIP_REG_3_ | ~new_P1_R2096_U94;
  assign new_P1_R2096_U9 = ~P1_REIP_REG_4_;
  assign new_P1_R2096_U10 = ~P1_REIP_REG_4_ | ~new_P1_R2096_U95;
  assign new_P1_R2096_U11 = ~P1_REIP_REG_5_;
  assign new_P1_R2096_U12 = ~P1_REIP_REG_5_ | ~new_P1_R2096_U96;
  assign new_P1_R2096_U13 = ~P1_REIP_REG_6_;
  assign new_P1_R2096_U14 = ~P1_REIP_REG_6_ | ~new_P1_R2096_U97;
  assign new_P1_R2096_U15 = ~P1_REIP_REG_7_;
  assign new_P1_R2096_U16 = ~P1_REIP_REG_7_ | ~new_P1_R2096_U98;
  assign new_P1_R2096_U17 = ~P1_REIP_REG_8_;
  assign new_P1_R2096_U18 = ~P1_REIP_REG_9_;
  assign new_P1_R2096_U19 = ~P1_REIP_REG_8_ | ~new_P1_R2096_U99;
  assign new_P1_R2096_U20 = ~new_P1_R2096_U100 | ~P1_REIP_REG_9_;
  assign new_P1_R2096_U21 = ~P1_REIP_REG_10_;
  assign new_P1_R2096_U22 = ~P1_REIP_REG_10_ | ~new_P1_R2096_U101;
  assign new_P1_R2096_U23 = ~P1_REIP_REG_11_;
  assign new_P1_R2096_U24 = ~P1_REIP_REG_11_ | ~new_P1_R2096_U102;
  assign new_P1_R2096_U25 = ~P1_REIP_REG_12_;
  assign new_P1_R2096_U26 = ~P1_REIP_REG_12_ | ~new_P1_R2096_U103;
  assign new_P1_R2096_U27 = ~P1_REIP_REG_13_;
  assign new_P1_R2096_U28 = ~P1_REIP_REG_13_ | ~new_P1_R2096_U104;
  assign new_P1_R2096_U29 = ~P1_REIP_REG_14_;
  assign new_P1_R2096_U30 = ~P1_REIP_REG_14_ | ~new_P1_R2096_U105;
  assign new_P1_R2096_U31 = ~P1_REIP_REG_15_;
  assign new_P1_R2096_U32 = ~P1_REIP_REG_15_ | ~new_P1_R2096_U106;
  assign new_P1_R2096_U33 = ~P1_REIP_REG_16_;
  assign new_P1_R2096_U34 = ~P1_REIP_REG_16_ | ~new_P1_R2096_U107;
  assign new_P1_R2096_U35 = ~P1_REIP_REG_17_;
  assign new_P1_R2096_U36 = ~P1_REIP_REG_17_ | ~new_P1_R2096_U108;
  assign new_P1_R2096_U37 = ~P1_REIP_REG_18_;
  assign new_P1_R2096_U38 = ~P1_REIP_REG_18_ | ~new_P1_R2096_U109;
  assign new_P1_R2096_U39 = ~P1_REIP_REG_19_;
  assign new_P1_R2096_U40 = ~P1_REIP_REG_19_ | ~new_P1_R2096_U110;
  assign new_P1_R2096_U41 = ~P1_REIP_REG_20_;
  assign new_P1_R2096_U42 = ~P1_REIP_REG_20_ | ~new_P1_R2096_U111;
  assign new_P1_R2096_U43 = ~P1_REIP_REG_21_;
  assign new_P1_R2096_U44 = ~P1_REIP_REG_21_ | ~new_P1_R2096_U112;
  assign new_P1_R2096_U45 = ~P1_REIP_REG_22_;
  assign new_P1_R2096_U46 = ~P1_REIP_REG_22_ | ~new_P1_R2096_U113;
  assign new_P1_R2096_U47 = ~P1_REIP_REG_23_;
  assign new_P1_R2096_U48 = ~P1_REIP_REG_23_ | ~new_P1_R2096_U114;
  assign new_P1_R2096_U49 = ~P1_REIP_REG_24_;
  assign new_P1_R2096_U50 = ~P1_REIP_REG_24_ | ~new_P1_R2096_U115;
  assign new_P1_R2096_U51 = ~P1_REIP_REG_25_;
  assign new_P1_R2096_U52 = ~P1_REIP_REG_25_ | ~new_P1_R2096_U116;
  assign new_P1_R2096_U53 = ~P1_REIP_REG_26_;
  assign new_P1_R2096_U54 = ~P1_REIP_REG_26_ | ~new_P1_R2096_U117;
  assign new_P1_R2096_U55 = ~P1_REIP_REG_27_;
  assign new_P1_R2096_U56 = ~P1_REIP_REG_27_ | ~new_P1_R2096_U118;
  assign new_P1_R2096_U57 = ~P1_REIP_REG_28_;
  assign new_P1_R2096_U58 = ~P1_REIP_REG_28_ | ~new_P1_R2096_U119;
  assign new_P1_R2096_U59 = ~P1_REIP_REG_29_;
  assign new_P1_R2096_U60 = ~P1_REIP_REG_29_ | ~new_P1_R2096_U120;
  assign new_P1_R2096_U61 = ~P1_REIP_REG_30_;
  assign new_P1_R2096_U62 = ~new_P1_R2096_U124 | ~new_P1_R2096_U123;
  assign new_P1_R2096_U63 = ~new_P1_R2096_U126 | ~new_P1_R2096_U125;
  assign new_P1_R2096_U64 = ~new_P1_R2096_U128 | ~new_P1_R2096_U127;
  assign new_P1_R2096_U65 = ~new_P1_R2096_U130 | ~new_P1_R2096_U129;
  assign new_P1_R2096_U66 = ~new_P1_R2096_U132 | ~new_P1_R2096_U131;
  assign new_P1_R2096_U67 = ~new_P1_R2096_U134 | ~new_P1_R2096_U133;
  assign new_P1_R2096_U68 = ~new_P1_R2096_U136 | ~new_P1_R2096_U135;
  assign new_P1_R2096_U69 = ~new_P1_R2096_U138 | ~new_P1_R2096_U137;
  assign new_P1_R2096_U70 = ~new_P1_R2096_U140 | ~new_P1_R2096_U139;
  assign new_P1_R2096_U71 = ~new_P1_R2096_U142 | ~new_P1_R2096_U141;
  assign new_P1_R2096_U72 = ~new_P1_R2096_U144 | ~new_P1_R2096_U143;
  assign new_P1_R2096_U73 = ~new_P1_R2096_U146 | ~new_P1_R2096_U145;
  assign new_P1_R2096_U74 = ~new_P1_R2096_U148 | ~new_P1_R2096_U147;
  assign new_P1_R2096_U75 = ~new_P1_R2096_U150 | ~new_P1_R2096_U149;
  assign new_P1_R2096_U76 = ~new_P1_R2096_U152 | ~new_P1_R2096_U151;
  assign new_P1_R2096_U77 = ~new_P1_R2096_U154 | ~new_P1_R2096_U153;
  assign new_P1_R2096_U78 = ~new_P1_R2096_U156 | ~new_P1_R2096_U155;
  assign new_P1_R2096_U79 = ~new_P1_R2096_U158 | ~new_P1_R2096_U157;
  assign new_P1_R2096_U80 = ~new_P1_R2096_U160 | ~new_P1_R2096_U159;
  assign new_P1_R2096_U81 = ~new_P1_R2096_U162 | ~new_P1_R2096_U161;
  assign new_P1_R2096_U82 = ~new_P1_R2096_U164 | ~new_P1_R2096_U163;
  assign new_P1_R2096_U83 = ~new_P1_R2096_U166 | ~new_P1_R2096_U165;
  assign new_P1_R2096_U84 = ~new_P1_R2096_U168 | ~new_P1_R2096_U167;
  assign new_P1_R2096_U85 = ~new_P1_R2096_U170 | ~new_P1_R2096_U169;
  assign new_P1_R2096_U86 = ~new_P1_R2096_U172 | ~new_P1_R2096_U171;
  assign new_P1_R2096_U87 = ~new_P1_R2096_U174 | ~new_P1_R2096_U173;
  assign new_P1_R2096_U88 = ~new_P1_R2096_U176 | ~new_P1_R2096_U175;
  assign new_P1_R2096_U89 = ~new_P1_R2096_U178 | ~new_P1_R2096_U177;
  assign new_P1_R2096_U90 = ~new_P1_R2096_U180 | ~new_P1_R2096_U179;
  assign new_P1_R2096_U91 = ~new_P1_R2096_U182 | ~new_P1_R2096_U181;
  assign new_P1_R2096_U92 = ~P1_REIP_REG_31_;
  assign new_P1_R2096_U93 = ~P1_REIP_REG_30_ | ~new_P1_R2096_U121;
  assign new_P1_R2096_U94 = ~new_P1_R2096_U6;
  assign new_P1_R2096_U95 = ~new_P1_R2096_U8;
  assign new_P1_R2096_U96 = ~new_P1_R2096_U10;
  assign new_P1_R2096_U97 = ~new_P1_R2096_U12;
  assign new_P1_R2096_U98 = ~new_P1_R2096_U14;
  assign new_P1_R2096_U99 = ~new_P1_R2096_U16;
  assign new_P1_R2096_U100 = ~new_P1_R2096_U19;
  assign new_P1_R2096_U101 = ~new_P1_R2096_U20;
  assign new_P1_R2096_U102 = ~new_P1_R2096_U22;
  assign new_P1_R2096_U103 = ~new_P1_R2096_U24;
  assign new_P1_R2096_U104 = ~new_P1_R2096_U26;
  assign new_P1_R2096_U105 = ~new_P1_R2096_U28;
  assign new_P1_R2096_U106 = ~new_P1_R2096_U30;
  assign new_P1_R2096_U107 = ~new_P1_R2096_U32;
  assign new_P1_R2096_U108 = ~new_P1_R2096_U34;
  assign new_P1_R2096_U109 = ~new_P1_R2096_U36;
  assign new_P1_R2096_U110 = ~new_P1_R2096_U38;
  assign new_P1_R2096_U111 = ~new_P1_R2096_U40;
  assign new_P1_R2096_U112 = ~new_P1_R2096_U42;
  assign new_P1_R2096_U113 = ~new_P1_R2096_U44;
  assign new_P1_R2096_U114 = ~new_P1_R2096_U46;
  assign new_P1_R2096_U115 = ~new_P1_R2096_U48;
  assign new_P1_R2096_U116 = ~new_P1_R2096_U50;
  assign new_P1_R2096_U117 = ~new_P1_R2096_U52;
  assign new_P1_R2096_U118 = ~new_P1_R2096_U54;
  assign new_P1_R2096_U119 = ~new_P1_R2096_U56;
  assign new_P1_R2096_U120 = ~new_P1_R2096_U58;
  assign new_P1_R2096_U121 = ~new_P1_R2096_U60;
  assign new_P1_R2096_U122 = ~new_P1_R2096_U93;
  assign new_P1_R2096_U123 = ~P1_REIP_REG_9_ | ~new_P1_R2096_U19;
  assign new_P1_R2096_U124 = ~new_P1_R2096_U100 | ~new_P1_R2096_U18;
  assign new_P1_R2096_U125 = ~P1_REIP_REG_8_ | ~new_P1_R2096_U16;
  assign new_P1_R2096_U126 = ~new_P1_R2096_U99 | ~new_P1_R2096_U17;
  assign new_P1_R2096_U127 = ~P1_REIP_REG_7_ | ~new_P1_R2096_U14;
  assign new_P1_R2096_U128 = ~new_P1_R2096_U98 | ~new_P1_R2096_U15;
  assign new_P1_R2096_U129 = ~P1_REIP_REG_6_ | ~new_P1_R2096_U12;
  assign new_P1_R2096_U130 = ~new_P1_R2096_U97 | ~new_P1_R2096_U13;
  assign new_P1_R2096_U131 = ~P1_REIP_REG_5_ | ~new_P1_R2096_U10;
  assign new_P1_R2096_U132 = ~new_P1_R2096_U96 | ~new_P1_R2096_U11;
  assign new_P1_R2096_U133 = ~P1_REIP_REG_4_ | ~new_P1_R2096_U8;
  assign new_P1_R2096_U134 = ~new_P1_R2096_U95 | ~new_P1_R2096_U9;
  assign new_P1_R2096_U135 = ~P1_REIP_REG_3_ | ~new_P1_R2096_U6;
  assign new_P1_R2096_U136 = ~new_P1_R2096_U94 | ~new_P1_R2096_U7;
  assign new_P1_R2096_U137 = ~P1_REIP_REG_31_ | ~new_P1_R2096_U93;
  assign new_P1_R2096_U138 = ~new_P1_R2096_U122 | ~new_P1_R2096_U92;
  assign new_P1_R2096_U139 = ~P1_REIP_REG_30_ | ~new_P1_R2096_U60;
  assign new_P1_R2096_U140 = ~new_P1_R2096_U121 | ~new_P1_R2096_U61;
  assign new_P1_R2096_U141 = ~P1_REIP_REG_2_ | ~new_P1_R2096_U4;
  assign new_P1_R2096_U142 = ~P1_REIP_REG_1_ | ~new_P1_R2096_U5;
  assign new_P1_R2096_U143 = ~P1_REIP_REG_29_ | ~new_P1_R2096_U58;
  assign new_P1_R2096_U144 = ~new_P1_R2096_U120 | ~new_P1_R2096_U59;
  assign new_P1_R2096_U145 = ~P1_REIP_REG_28_ | ~new_P1_R2096_U56;
  assign new_P1_R2096_U146 = ~new_P1_R2096_U119 | ~new_P1_R2096_U57;
  assign new_P1_R2096_U147 = ~P1_REIP_REG_27_ | ~new_P1_R2096_U54;
  assign new_P1_R2096_U148 = ~new_P1_R2096_U118 | ~new_P1_R2096_U55;
  assign new_P1_R2096_U149 = ~P1_REIP_REG_26_ | ~new_P1_R2096_U52;
  assign new_P1_R2096_U150 = ~new_P1_R2096_U117 | ~new_P1_R2096_U53;
  assign new_P1_R2096_U151 = ~P1_REIP_REG_25_ | ~new_P1_R2096_U50;
  assign new_P1_R2096_U152 = ~new_P1_R2096_U116 | ~new_P1_R2096_U51;
  assign new_P1_R2096_U153 = ~P1_REIP_REG_24_ | ~new_P1_R2096_U48;
  assign new_P1_R2096_U154 = ~new_P1_R2096_U115 | ~new_P1_R2096_U49;
  assign new_P1_R2096_U155 = ~P1_REIP_REG_23_ | ~new_P1_R2096_U46;
  assign new_P1_R2096_U156 = ~new_P1_R2096_U114 | ~new_P1_R2096_U47;
  assign new_P1_R2096_U157 = ~P1_REIP_REG_22_ | ~new_P1_R2096_U44;
  assign new_P1_R2096_U158 = ~new_P1_R2096_U113 | ~new_P1_R2096_U45;
  assign new_P1_R2096_U159 = ~P1_REIP_REG_21_ | ~new_P1_R2096_U42;
  assign new_P1_R2096_U160 = ~new_P1_R2096_U112 | ~new_P1_R2096_U43;
  assign new_P1_R2096_U161 = ~P1_REIP_REG_20_ | ~new_P1_R2096_U40;
  assign new_P1_R2096_U162 = ~new_P1_R2096_U111 | ~new_P1_R2096_U41;
  assign new_P1_R2096_U163 = ~P1_REIP_REG_19_ | ~new_P1_R2096_U38;
  assign new_P1_R2096_U164 = ~new_P1_R2096_U110 | ~new_P1_R2096_U39;
  assign new_P1_R2096_U165 = ~P1_REIP_REG_18_ | ~new_P1_R2096_U36;
  assign new_P1_R2096_U166 = ~new_P1_R2096_U109 | ~new_P1_R2096_U37;
  assign new_P1_R2096_U167 = ~P1_REIP_REG_17_ | ~new_P1_R2096_U34;
  assign new_P1_R2096_U168 = ~new_P1_R2096_U108 | ~new_P1_R2096_U35;
  assign new_P1_R2096_U169 = ~P1_REIP_REG_16_ | ~new_P1_R2096_U32;
  assign new_P1_R2096_U170 = ~new_P1_R2096_U107 | ~new_P1_R2096_U33;
  assign new_P1_R2096_U171 = ~P1_REIP_REG_15_ | ~new_P1_R2096_U30;
  assign new_P1_R2096_U172 = ~new_P1_R2096_U106 | ~new_P1_R2096_U31;
  assign new_P1_R2096_U173 = ~P1_REIP_REG_14_ | ~new_P1_R2096_U28;
  assign new_P1_R2096_U174 = ~new_P1_R2096_U105 | ~new_P1_R2096_U29;
  assign new_P1_R2096_U175 = ~P1_REIP_REG_13_ | ~new_P1_R2096_U26;
  assign new_P1_R2096_U176 = ~new_P1_R2096_U104 | ~new_P1_R2096_U27;
  assign new_P1_R2096_U177 = ~P1_REIP_REG_12_ | ~new_P1_R2096_U24;
  assign new_P1_R2096_U178 = ~new_P1_R2096_U103 | ~new_P1_R2096_U25;
  assign new_P1_R2096_U179 = ~P1_REIP_REG_11_ | ~new_P1_R2096_U22;
  assign new_P1_R2096_U180 = ~new_P1_R2096_U102 | ~new_P1_R2096_U23;
  assign new_P1_R2096_U181 = ~P1_REIP_REG_10_ | ~new_P1_R2096_U20;
  assign new_P1_R2096_U182 = ~new_P1_R2096_U101 | ~new_P1_R2096_U21;
  assign new_P1_LT_563_U6 = new_P1_LT_563_U27 & new_P1_LT_563_U26;
  assign new_P1_LT_563_U7 = ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P1_LT_563_U8 = ~new_P1_U3491;
  assign new_P1_LT_563_U9 = ~new_P1_U3490;
  assign new_P1_LT_563_U10 = ~P1_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P1_LT_563_U11 = ~P1_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P1_LT_563_U12 = ~new_P1_U3489;
  assign new_P1_LT_563_U13 = new_P1_LT_563_U21 & new_P1_LT_563_U22;
  assign new_P1_LT_563_U14 = new_P1_LT_563_U24 & new_P1_LT_563_U25;
  assign new_P1_LT_563_U15 = ~new_P1_U3492;
  assign new_P1_LT_563_U16 = ~new_P1_U3493;
  assign new_P1_LT_563_U17 = ~P1_INSTQUEUEWR_ADDR_REG_0_ | ~new_P1_LT_563_U16 | ~new_P1_LT_563_U15;
  assign new_P1_LT_563_U18 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_LT_563_U15;
  assign new_P1_LT_563_U19 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_LT_563_U8;
  assign new_P1_LT_563_U20 = ~new_P1_LT_563_U17 | ~new_P1_LT_563_U18 | ~new_P1_LT_563_U28 | ~new_P1_LT_563_U19;
  assign new_P1_LT_563_U21 = ~new_P1_U3491 | ~new_P1_LT_563_U7;
  assign new_P1_LT_563_U22 = ~new_P1_U3490 | ~new_P1_LT_563_U10;
  assign new_P1_LT_563_U23 = ~new_P1_LT_563_U13 | ~new_P1_LT_563_U20;
  assign new_P1_LT_563_U24 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_LT_563_U9;
  assign new_P1_LT_563_U25 = ~P1_INSTQUEUEWR_ADDR_REG_4_ | ~new_P1_LT_563_U12;
  assign new_P1_LT_563_U26 = ~new_P1_LT_563_U14 | ~new_P1_LT_563_U23;
  assign new_P1_LT_563_U27 = ~new_P1_U3489 | ~new_P1_LT_563_U11;
  assign new_P1_LT_563_U28 = ~new_P1_LT_563_U16 | ~P1_INSTQUEUEWR_ADDR_REG_0_ | ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P1_R2238_U6 = ~new_P1_R2238_U45 | ~new_P1_R2238_U44;
  assign new_P1_R2238_U7 = ~new_P1_R2238_U9 | ~new_P1_R2238_U46;
  assign new_P1_R2238_U8 = ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_R2238_U9 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~new_P1_R2238_U18;
  assign new_P1_R2238_U10 = ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P1_R2238_U11 = ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_R2238_U12 = ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P1_R2238_U13 = ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_R2238_U14 = ~P1_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P1_R2238_U15 = ~P1_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P1_R2238_U16 = ~new_P1_R2238_U41 | ~new_P1_R2238_U40;
  assign new_P1_R2238_U17 = ~P1_INSTQUEUERD_ADDR_REG_4_;
  assign new_P1_R2238_U18 = ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P1_R2238_U19 = ~new_P1_R2238_U51 | ~new_P1_R2238_U50;
  assign new_P1_R2238_U20 = ~new_P1_R2238_U56 | ~new_P1_R2238_U55;
  assign new_P1_R2238_U21 = ~new_P1_R2238_U61 | ~new_P1_R2238_U60;
  assign new_P1_R2238_U22 = ~new_P1_R2238_U66 | ~new_P1_R2238_U65;
  assign new_P1_R2238_U23 = ~new_P1_R2238_U48 | ~new_P1_R2238_U47;
  assign new_P1_R2238_U24 = ~new_P1_R2238_U53 | ~new_P1_R2238_U52;
  assign new_P1_R2238_U25 = ~new_P1_R2238_U58 | ~new_P1_R2238_U57;
  assign new_P1_R2238_U26 = ~new_P1_R2238_U63 | ~new_P1_R2238_U62;
  assign new_P1_R2238_U27 = ~new_P1_R2238_U37 | ~new_P1_R2238_U36;
  assign new_P1_R2238_U28 = ~new_P1_R2238_U33 | ~new_P1_R2238_U32;
  assign new_P1_R2238_U29 = ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_R2238_U30 = ~new_P1_R2238_U9;
  assign new_P1_R2238_U31 = ~new_P1_R2238_U30 | ~new_P1_R2238_U10;
  assign new_P1_R2238_U32 = ~new_P1_R2238_U31 | ~new_P1_R2238_U29;
  assign new_P1_R2238_U33 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_R2238_U9;
  assign new_P1_R2238_U34 = ~new_P1_R2238_U28;
  assign new_P1_R2238_U35 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_R2238_U12;
  assign new_P1_R2238_U36 = ~new_P1_R2238_U35 | ~new_P1_R2238_U28;
  assign new_P1_R2238_U37 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_R2238_U11;
  assign new_P1_R2238_U38 = ~new_P1_R2238_U27;
  assign new_P1_R2238_U39 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_R2238_U14;
  assign new_P1_R2238_U40 = ~new_P1_R2238_U39 | ~new_P1_R2238_U27;
  assign new_P1_R2238_U41 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_R2238_U13;
  assign new_P1_R2238_U42 = ~new_P1_R2238_U16;
  assign new_P1_R2238_U43 = ~P1_INSTQUEUEWR_ADDR_REG_4_ | ~new_P1_R2238_U17;
  assign new_P1_R2238_U44 = ~new_P1_R2238_U42 | ~new_P1_R2238_U43;
  assign new_P1_R2238_U45 = ~P1_INSTQUEUERD_ADDR_REG_4_ | ~new_P1_R2238_U15;
  assign new_P1_R2238_U46 = ~P1_INSTQUEUEWR_ADDR_REG_0_ | ~new_P1_R2238_U8;
  assign new_P1_R2238_U47 = ~P1_INSTQUEUERD_ADDR_REG_4_ | ~new_P1_R2238_U15;
  assign new_P1_R2238_U48 = ~P1_INSTQUEUEWR_ADDR_REG_4_ | ~new_P1_R2238_U17;
  assign new_P1_R2238_U49 = ~new_P1_R2238_U23;
  assign new_P1_R2238_U50 = ~new_P1_R2238_U49 | ~new_P1_R2238_U42;
  assign new_P1_R2238_U51 = ~new_P1_R2238_U23 | ~new_P1_R2238_U16;
  assign new_P1_R2238_U52 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_R2238_U14;
  assign new_P1_R2238_U53 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_R2238_U13;
  assign new_P1_R2238_U54 = ~new_P1_R2238_U24;
  assign new_P1_R2238_U55 = ~new_P1_R2238_U38 | ~new_P1_R2238_U54;
  assign new_P1_R2238_U56 = ~new_P1_R2238_U24 | ~new_P1_R2238_U27;
  assign new_P1_R2238_U57 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_R2238_U12;
  assign new_P1_R2238_U58 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_R2238_U11;
  assign new_P1_R2238_U59 = ~new_P1_R2238_U25;
  assign new_P1_R2238_U60 = ~new_P1_R2238_U34 | ~new_P1_R2238_U59;
  assign new_P1_R2238_U61 = ~new_P1_R2238_U25 | ~new_P1_R2238_U28;
  assign new_P1_R2238_U62 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_R2238_U10;
  assign new_P1_R2238_U63 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_R2238_U29;
  assign new_P1_R2238_U64 = ~new_P1_R2238_U26;
  assign new_P1_R2238_U65 = ~new_P1_R2238_U64 | ~new_P1_R2238_U30;
  assign new_P1_R2238_U66 = ~new_P1_R2238_U26 | ~new_P1_R2238_U9;
  assign new_P1_SUB_450_U6 = ~new_P1_SUB_450_U45 | ~new_P1_SUB_450_U44;
  assign new_P1_SUB_450_U7 = ~new_P1_SUB_450_U9 | ~new_P1_SUB_450_U46;
  assign new_P1_SUB_450_U8 = ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign new_P1_SUB_450_U9 = ~P1_INSTQUEUERD_ADDR_REG_0_ | ~new_P1_SUB_450_U18;
  assign new_P1_SUB_450_U10 = ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign new_P1_SUB_450_U11 = ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign new_P1_SUB_450_U12 = ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign new_P1_SUB_450_U13 = ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign new_P1_SUB_450_U14 = ~P1_INSTQUEUEWR_ADDR_REG_3_;
  assign new_P1_SUB_450_U15 = ~P1_INSTQUEUEWR_ADDR_REG_4_;
  assign new_P1_SUB_450_U16 = ~new_P1_SUB_450_U41 | ~new_P1_SUB_450_U40;
  assign new_P1_SUB_450_U17 = ~P1_INSTQUEUERD_ADDR_REG_4_;
  assign new_P1_SUB_450_U18 = ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign new_P1_SUB_450_U19 = ~new_P1_SUB_450_U51 | ~new_P1_SUB_450_U50;
  assign new_P1_SUB_450_U20 = ~new_P1_SUB_450_U56 | ~new_P1_SUB_450_U55;
  assign new_P1_SUB_450_U21 = ~new_P1_SUB_450_U61 | ~new_P1_SUB_450_U60;
  assign new_P1_SUB_450_U22 = ~new_P1_SUB_450_U66 | ~new_P1_SUB_450_U65;
  assign new_P1_SUB_450_U23 = ~new_P1_SUB_450_U48 | ~new_P1_SUB_450_U47;
  assign new_P1_SUB_450_U24 = ~new_P1_SUB_450_U53 | ~new_P1_SUB_450_U52;
  assign new_P1_SUB_450_U25 = ~new_P1_SUB_450_U58 | ~new_P1_SUB_450_U57;
  assign new_P1_SUB_450_U26 = ~new_P1_SUB_450_U63 | ~new_P1_SUB_450_U62;
  assign new_P1_SUB_450_U27 = ~new_P1_SUB_450_U37 | ~new_P1_SUB_450_U36;
  assign new_P1_SUB_450_U28 = ~new_P1_SUB_450_U33 | ~new_P1_SUB_450_U32;
  assign new_P1_SUB_450_U29 = ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign new_P1_SUB_450_U30 = ~new_P1_SUB_450_U9;
  assign new_P1_SUB_450_U31 = ~new_P1_SUB_450_U30 | ~new_P1_SUB_450_U10;
  assign new_P1_SUB_450_U32 = ~new_P1_SUB_450_U31 | ~new_P1_SUB_450_U29;
  assign new_P1_SUB_450_U33 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_SUB_450_U9;
  assign new_P1_SUB_450_U34 = ~new_P1_SUB_450_U28;
  assign new_P1_SUB_450_U35 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_SUB_450_U12;
  assign new_P1_SUB_450_U36 = ~new_P1_SUB_450_U35 | ~new_P1_SUB_450_U28;
  assign new_P1_SUB_450_U37 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_SUB_450_U11;
  assign new_P1_SUB_450_U38 = ~new_P1_SUB_450_U27;
  assign new_P1_SUB_450_U39 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_SUB_450_U14;
  assign new_P1_SUB_450_U40 = ~new_P1_SUB_450_U39 | ~new_P1_SUB_450_U27;
  assign new_P1_SUB_450_U41 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_SUB_450_U13;
  assign new_P1_SUB_450_U42 = ~new_P1_SUB_450_U16;
  assign new_P1_SUB_450_U43 = ~P1_INSTQUEUEWR_ADDR_REG_4_ | ~new_P1_SUB_450_U17;
  assign new_P1_SUB_450_U44 = ~new_P1_SUB_450_U42 | ~new_P1_SUB_450_U43;
  assign new_P1_SUB_450_U45 = ~P1_INSTQUEUERD_ADDR_REG_4_ | ~new_P1_SUB_450_U15;
  assign new_P1_SUB_450_U46 = ~P1_INSTQUEUEWR_ADDR_REG_0_ | ~new_P1_SUB_450_U8;
  assign new_P1_SUB_450_U47 = ~P1_INSTQUEUERD_ADDR_REG_4_ | ~new_P1_SUB_450_U15;
  assign new_P1_SUB_450_U48 = ~P1_INSTQUEUEWR_ADDR_REG_4_ | ~new_P1_SUB_450_U17;
  assign new_P1_SUB_450_U49 = ~new_P1_SUB_450_U23;
  assign new_P1_SUB_450_U50 = ~new_P1_SUB_450_U49 | ~new_P1_SUB_450_U42;
  assign new_P1_SUB_450_U51 = ~new_P1_SUB_450_U23 | ~new_P1_SUB_450_U16;
  assign new_P1_SUB_450_U52 = ~P1_INSTQUEUERD_ADDR_REG_3_ | ~new_P1_SUB_450_U14;
  assign new_P1_SUB_450_U53 = ~P1_INSTQUEUEWR_ADDR_REG_3_ | ~new_P1_SUB_450_U13;
  assign new_P1_SUB_450_U54 = ~new_P1_SUB_450_U24;
  assign new_P1_SUB_450_U55 = ~new_P1_SUB_450_U38 | ~new_P1_SUB_450_U54;
  assign new_P1_SUB_450_U56 = ~new_P1_SUB_450_U24 | ~new_P1_SUB_450_U27;
  assign new_P1_SUB_450_U57 = ~P1_INSTQUEUERD_ADDR_REG_2_ | ~new_P1_SUB_450_U12;
  assign new_P1_SUB_450_U58 = ~P1_INSTQUEUEWR_ADDR_REG_2_ | ~new_P1_SUB_450_U11;
  assign new_P1_SUB_450_U59 = ~new_P1_SUB_450_U25;
  assign new_P1_SUB_450_U60 = ~new_P1_SUB_450_U34 | ~new_P1_SUB_450_U59;
  assign new_P1_SUB_450_U61 = ~new_P1_SUB_450_U25 | ~new_P1_SUB_450_U28;
  assign new_P1_SUB_450_U62 = ~P1_INSTQUEUERD_ADDR_REG_1_ | ~new_P1_SUB_450_U10;
  assign new_P1_SUB_450_U63 = ~P1_INSTQUEUEWR_ADDR_REG_1_ | ~new_P1_SUB_450_U29;
  assign new_P1_SUB_450_U64 = ~new_P1_SUB_450_U26;
  assign new_P1_SUB_450_U65 = ~new_P1_SUB_450_U64 | ~new_P1_SUB_450_U30;
  assign new_P1_SUB_450_U66 = ~new_P1_SUB_450_U26 | ~new_P1_SUB_450_U9;
  assign new_P1_ADD_371_U4 = ~new_P1_U3227;
  assign new_P1_ADD_371_U5 = ~new_P1_ADD_371_U23 | ~new_P1_ADD_371_U31;
  assign new_P1_ADD_371_U6 = new_P1_ADD_371_U22 & new_P1_ADD_371_U30;
  assign new_P1_ADD_371_U7 = ~new_P1_U3228;
  assign new_P1_ADD_371_U8 = ~new_P1_U3230;
  assign new_P1_ADD_371_U9 = ~new_P1_U3230 | ~new_P1_ADD_371_U23;
  assign new_P1_ADD_371_U10 = ~new_P1_U3231;
  assign new_P1_ADD_371_U11 = ~new_P1_U3231 | ~new_P1_ADD_371_U28;
  assign new_P1_ADD_371_U12 = ~new_P1_U3232;
  assign new_P1_ADD_371_U13 = ~new_P1_U3233;
  assign new_P1_ADD_371_U14 = ~new_P1_U3232 | ~new_P1_ADD_371_U29;
  assign new_P1_ADD_371_U15 = ~new_P1_U3229;
  assign new_P1_ADD_371_U16 = ~new_P1_U3234;
  assign new_P1_ADD_371_U17 = ~new_P1_ADD_371_U34 | ~new_P1_ADD_371_U33;
  assign new_P1_ADD_371_U18 = ~new_P1_ADD_371_U36 | ~new_P1_ADD_371_U35;
  assign new_P1_ADD_371_U19 = ~new_P1_ADD_371_U38 | ~new_P1_ADD_371_U37;
  assign new_P1_ADD_371_U20 = ~new_P1_ADD_371_U42 | ~new_P1_ADD_371_U41;
  assign new_P1_ADD_371_U21 = ~new_P1_ADD_371_U44 | ~new_P1_ADD_371_U43;
  assign new_P1_ADD_371_U22 = new_P1_U3234 & new_P1_U3233;
  assign new_P1_ADD_371_U23 = ~new_P1_ADD_371_U15 | ~new_P1_ADD_371_U26;
  assign new_P1_ADD_371_U24 = new_P1_ADD_371_U40 & new_P1_ADD_371_U39;
  assign new_P1_ADD_371_U25 = ~new_P1_ADD_371_U30 | ~new_P1_U3233;
  assign new_P1_ADD_371_U26 = ~new_P1_U3228 | ~new_P1_U3227;
  assign new_P1_ADD_371_U27 = ~new_P1_ADD_371_U23;
  assign new_P1_ADD_371_U28 = ~new_P1_ADD_371_U9;
  assign new_P1_ADD_371_U29 = ~new_P1_ADD_371_U11;
  assign new_P1_ADD_371_U30 = ~new_P1_ADD_371_U14;
  assign new_P1_ADD_371_U31 = ~new_P1_U3229 | ~new_P1_U3228 | ~new_P1_U3227;
  assign new_P1_ADD_371_U32 = ~new_P1_ADD_371_U25;
  assign new_P1_ADD_371_U33 = ~new_P1_U3233 | ~new_P1_ADD_371_U14;
  assign new_P1_ADD_371_U34 = ~new_P1_ADD_371_U30 | ~new_P1_ADD_371_U13;
  assign new_P1_ADD_371_U35 = ~new_P1_U3231 | ~new_P1_ADD_371_U9;
  assign new_P1_ADD_371_U36 = ~new_P1_ADD_371_U28 | ~new_P1_ADD_371_U10;
  assign new_P1_ADD_371_U37 = ~new_P1_U3232 | ~new_P1_ADD_371_U11;
  assign new_P1_ADD_371_U38 = ~new_P1_ADD_371_U29 | ~new_P1_ADD_371_U12;
  assign new_P1_ADD_371_U39 = ~new_P1_U3230 | ~new_P1_ADD_371_U23;
  assign new_P1_ADD_371_U40 = ~new_P1_ADD_371_U27 | ~new_P1_ADD_371_U8;
  assign new_P1_ADD_371_U41 = ~new_P1_U3228 | ~new_P1_ADD_371_U4;
  assign new_P1_ADD_371_U42 = ~new_P1_U3227 | ~new_P1_ADD_371_U7;
  assign new_P1_ADD_371_U43 = ~new_P1_U3234 | ~new_P1_ADD_371_U25;
  assign new_P1_ADD_371_U44 = ~new_P1_ADD_371_U32 | ~new_P1_ADD_371_U16;
  assign new_P1_ADD_405_U4 = ~P1_INSTADDRPOINTER_REG_0_;
  assign new_P1_ADD_405_U5 = ~new_P1_ADD_405_U94 | ~new_P1_ADD_405_U125;
  assign new_P1_ADD_405_U6 = ~P1_INSTADDRPOINTER_REG_1_;
  assign new_P1_ADD_405_U7 = ~P1_INSTADDRPOINTER_REG_3_;
  assign new_P1_ADD_405_U8 = ~P1_INSTADDRPOINTER_REG_3_ | ~new_P1_ADD_405_U94;
  assign new_P1_ADD_405_U9 = ~P1_INSTADDRPOINTER_REG_4_;
  assign new_P1_ADD_405_U10 = ~P1_INSTADDRPOINTER_REG_4_ | ~new_P1_ADD_405_U98;
  assign new_P1_ADD_405_U11 = ~P1_INSTADDRPOINTER_REG_5_;
  assign new_P1_ADD_405_U12 = ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_ADD_405_U13 = ~P1_INSTADDRPOINTER_REG_5_ | ~new_P1_ADD_405_U99;
  assign new_P1_ADD_405_U14 = ~new_P1_ADD_405_U100 | ~P1_INSTADDRPOINTER_REG_6_;
  assign new_P1_ADD_405_U15 = ~P1_INSTADDRPOINTER_REG_7_;
  assign new_P1_ADD_405_U16 = ~P1_INSTADDRPOINTER_REG_7_ | ~new_P1_ADD_405_U101;
  assign new_P1_ADD_405_U17 = ~P1_INSTADDRPOINTER_REG_8_;
  assign new_P1_ADD_405_U18 = ~P1_INSTADDRPOINTER_REG_8_ | ~new_P1_ADD_405_U102;
  assign new_P1_ADD_405_U19 = ~P1_INSTADDRPOINTER_REG_9_;
  assign new_P1_ADD_405_U20 = ~P1_INSTADDRPOINTER_REG_9_ | ~new_P1_ADD_405_U103;
  assign new_P1_ADD_405_U21 = ~P1_INSTADDRPOINTER_REG_10_;
  assign new_P1_ADD_405_U22 = ~P1_INSTADDRPOINTER_REG_10_ | ~new_P1_ADD_405_U104;
  assign new_P1_ADD_405_U23 = ~P1_INSTADDRPOINTER_REG_11_;
  assign new_P1_ADD_405_U24 = ~P1_INSTADDRPOINTER_REG_11_ | ~new_P1_ADD_405_U105;
  assign new_P1_ADD_405_U25 = ~P1_INSTADDRPOINTER_REG_12_;
  assign new_P1_ADD_405_U26 = ~P1_INSTADDRPOINTER_REG_12_ | ~new_P1_ADD_405_U106;
  assign new_P1_ADD_405_U27 = ~P1_INSTADDRPOINTER_REG_13_;
  assign new_P1_ADD_405_U28 = ~P1_INSTADDRPOINTER_REG_13_ | ~new_P1_ADD_405_U107;
  assign new_P1_ADD_405_U29 = ~P1_INSTADDRPOINTER_REG_14_;
  assign new_P1_ADD_405_U30 = ~P1_INSTADDRPOINTER_REG_14_ | ~new_P1_ADD_405_U108;
  assign new_P1_ADD_405_U31 = ~P1_INSTADDRPOINTER_REG_15_;
  assign new_P1_ADD_405_U32 = ~P1_INSTADDRPOINTER_REG_15_ | ~new_P1_ADD_405_U109;
  assign new_P1_ADD_405_U33 = ~P1_INSTADDRPOINTER_REG_16_;
  assign new_P1_ADD_405_U34 = ~P1_INSTADDRPOINTER_REG_16_ | ~new_P1_ADD_405_U110;
  assign new_P1_ADD_405_U35 = ~P1_INSTADDRPOINTER_REG_17_;
  assign new_P1_ADD_405_U36 = ~P1_INSTADDRPOINTER_REG_17_ | ~new_P1_ADD_405_U111;
  assign new_P1_ADD_405_U37 = ~P1_INSTADDRPOINTER_REG_18_;
  assign new_P1_ADD_405_U38 = ~P1_INSTADDRPOINTER_REG_18_ | ~new_P1_ADD_405_U112;
  assign new_P1_ADD_405_U39 = ~P1_INSTADDRPOINTER_REG_19_;
  assign new_P1_ADD_405_U40 = ~P1_INSTADDRPOINTER_REG_19_ | ~new_P1_ADD_405_U113;
  assign new_P1_ADD_405_U41 = ~P1_INSTADDRPOINTER_REG_20_;
  assign new_P1_ADD_405_U42 = ~P1_INSTADDRPOINTER_REG_20_ | ~new_P1_ADD_405_U114;
  assign new_P1_ADD_405_U43 = ~P1_INSTADDRPOINTER_REG_21_;
  assign new_P1_ADD_405_U44 = ~P1_INSTADDRPOINTER_REG_21_ | ~new_P1_ADD_405_U115;
  assign new_P1_ADD_405_U45 = ~P1_INSTADDRPOINTER_REG_22_;
  assign new_P1_ADD_405_U46 = ~P1_INSTADDRPOINTER_REG_22_ | ~new_P1_ADD_405_U116;
  assign new_P1_ADD_405_U47 = ~P1_INSTADDRPOINTER_REG_23_;
  assign new_P1_ADD_405_U48 = ~P1_INSTADDRPOINTER_REG_23_ | ~new_P1_ADD_405_U117;
  assign new_P1_ADD_405_U49 = ~P1_INSTADDRPOINTER_REG_24_;
  assign new_P1_ADD_405_U50 = ~P1_INSTADDRPOINTER_REG_24_ | ~new_P1_ADD_405_U118;
  assign new_P1_ADD_405_U51 = ~P1_INSTADDRPOINTER_REG_25_;
  assign new_P1_ADD_405_U52 = ~P1_INSTADDRPOINTER_REG_25_ | ~new_P1_ADD_405_U119;
  assign new_P1_ADD_405_U53 = ~P1_INSTADDRPOINTER_REG_26_;
  assign new_P1_ADD_405_U54 = ~P1_INSTADDRPOINTER_REG_26_ | ~new_P1_ADD_405_U120;
  assign new_P1_ADD_405_U55 = ~P1_INSTADDRPOINTER_REG_27_;
  assign new_P1_ADD_405_U56 = ~P1_INSTADDRPOINTER_REG_27_ | ~new_P1_ADD_405_U121;
  assign new_P1_ADD_405_U57 = ~P1_INSTADDRPOINTER_REG_28_;
  assign new_P1_ADD_405_U58 = ~P1_INSTADDRPOINTER_REG_28_ | ~new_P1_ADD_405_U122;
  assign new_P1_ADD_405_U59 = ~P1_INSTADDRPOINTER_REG_29_;
  assign new_P1_ADD_405_U60 = ~P1_INSTADDRPOINTER_REG_30_;
  assign new_P1_ADD_405_U61 = ~P1_INSTADDRPOINTER_REG_29_ | ~new_P1_ADD_405_U123;
  assign new_P1_ADD_405_U62 = ~P1_INSTADDRPOINTER_REG_2_;
  assign new_P1_ADD_405_U63 = ~new_P1_ADD_405_U128 | ~new_P1_ADD_405_U127;
  assign new_P1_ADD_405_U64 = ~new_P1_ADD_405_U130 | ~new_P1_ADD_405_U129;
  assign new_P1_ADD_405_U65 = ~new_P1_ADD_405_U132 | ~new_P1_ADD_405_U131;
  assign new_P1_ADD_405_U66 = ~new_P1_ADD_405_U134 | ~new_P1_ADD_405_U133;
  assign new_P1_ADD_405_U67 = ~new_P1_ADD_405_U136 | ~new_P1_ADD_405_U135;
  assign new_P1_ADD_405_U68 = ~new_P1_ADD_405_U138 | ~new_P1_ADD_405_U137;
  assign new_P1_ADD_405_U69 = ~new_P1_ADD_405_U140 | ~new_P1_ADD_405_U139;
  assign new_P1_ADD_405_U70 = ~new_P1_ADD_405_U142 | ~new_P1_ADD_405_U141;
  assign new_P1_ADD_405_U71 = ~new_P1_ADD_405_U144 | ~new_P1_ADD_405_U143;
  assign new_P1_ADD_405_U72 = ~new_P1_ADD_405_U146 | ~new_P1_ADD_405_U145;
  assign new_P1_ADD_405_U73 = ~new_P1_ADD_405_U148 | ~new_P1_ADD_405_U147;
  assign new_P1_ADD_405_U74 = ~new_P1_ADD_405_U150 | ~new_P1_ADD_405_U149;
  assign new_P1_ADD_405_U75 = ~new_P1_ADD_405_U152 | ~new_P1_ADD_405_U151;
  assign new_P1_ADD_405_U76 = ~new_P1_ADD_405_U154 | ~new_P1_ADD_405_U153;
  assign new_P1_ADD_405_U77 = ~new_P1_ADD_405_U156 | ~new_P1_ADD_405_U155;
  assign new_P1_ADD_405_U78 = ~new_P1_ADD_405_U158 | ~new_P1_ADD_405_U157;
  assign new_P1_ADD_405_U79 = ~new_P1_ADD_405_U160 | ~new_P1_ADD_405_U159;
  assign new_P1_ADD_405_U80 = ~new_P1_ADD_405_U162 | ~new_P1_ADD_405_U161;
  assign new_P1_ADD_405_U81 = ~new_P1_ADD_405_U164 | ~new_P1_ADD_405_U163;
  assign new_P1_ADD_405_U82 = ~new_P1_ADD_405_U166 | ~new_P1_ADD_405_U165;
  assign new_P1_ADD_405_U83 = ~new_P1_ADD_405_U168 | ~new_P1_ADD_405_U167;
  assign new_P1_ADD_405_U84 = ~new_P1_ADD_405_U170 | ~new_P1_ADD_405_U169;
  assign new_P1_ADD_405_U85 = ~new_P1_ADD_405_U174 | ~new_P1_ADD_405_U173;
  assign new_P1_ADD_405_U86 = ~new_P1_ADD_405_U176 | ~new_P1_ADD_405_U175;
  assign new_not_keyinput0 = ~keyinput0;
  assign new_not_keyinput1 = ~keyinput1;
  assign new_not_keyinput2 = ~keyinput2;
  assign new_not_keyinput3 = ~keyinput3;
  assign new_not_keyinput4 = ~keyinput4;
  assign new_not_0 = ~Q_1;
  assign new_and_1 = new_not_0 & Q_3;
  assign new_not_2 = ~Q_2;
  assign new_and_3 = new_not_2 & Q_3;
  assign new_not_4 = ~Q_0;
  assign new_and_5 = new_not_4 & Q_3;
  assign new_not_6 = ~Q_3;
  assign new_and_7 = new_not_6 & Q_2 & Q_0 & Q_1;
  assign n67464 = new_and_7 | new_and_5 | new_and_1 | new_and_3;
  assign new_not_9 = ~Q_2;
  assign new_and_10 = new_not_9 & Q_0 & Q_1;
  assign new_not_11 = ~Q_0;
  assign new_and_12 = new_not_11 & Q_2;
  assign new_not_13 = ~Q_1;
  assign new_and_14 = new_not_13 & Q_2;
  assign n67461 = new_and_14 | new_and_10 | new_and_12;
  assign new_not_16 = ~Q_1;
  assign new_and_17 = Q_0 & new_not_16;
  assign new_not_18 = ~Q_0;
  assign new_and_19 = new_not_18 & Q_1;
  assign n67458 = new_and_17 | new_and_19;
  assign n67455 = ~Q_0;
  assign new_not_Q_0 = ~Q_0;
  assign new_not_Q_1 = ~Q_1;
  assign new_not_Q_2 = ~Q_2;
  assign new_not_Q_3 = ~Q_3;
  assign new_count_state_1 = Q_0 & new_not_Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_2 = new_not_Q_0 & Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_3 = Q_0 & Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_4 = new_not_Q_0 & new_not_Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_5 = Q_0 & new_not_Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_6 = new_not_Q_0 & Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_7 = Q_0 & Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_8 = new_not_Q_0 & new_not_Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_9 = Q_0 & new_not_Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_10 = new_not_Q_0 & Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_11 = Q_0 & Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_12 = new_not_Q_0 & new_not_Q_1 & Q_3 & Q_2;
  assign new_count_state_13 = Q_0 & new_not_Q_1 & Q_3 & Q_2;
  assign new_count_state_14 = new_not_Q_0 & Q_1 & Q_3 & Q_2;
  assign new_count_state_15 = Q_0 & Q_1 & Q_3 & Q_2;
  assign new_y_mux_key0_and_0 = n290 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key0_and_1 = new_U247 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0 = new_y_mux_key0_and_0 | new_y_mux_key0_and_1;
  assign new_y_mux_key1_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_1 = new_U247 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1 = new_y_mux_key1_and_0 | new_y_mux_key1_and_1;
  assign new_y_mux_key2_and_0 = n290 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_1 = new_U247 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2 = new_y_mux_key2_and_0 | new_y_mux_key2_and_1;
  assign new_y_mux_key3_and_0 = n290 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key3_and_1 = new_U247 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3 = new_y_mux_key3_and_0 | new_y_mux_key3_and_1;
  assign new_y_mux_key4_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key4_and_1 = new_U247 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4 = new_y_mux_key4_and_0 | new_y_mux_key4_and_1;
  assign new_y_mux_key5_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key5_and_1 = new_U247 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5 = new_y_mux_key5_and_0 | new_y_mux_key5_and_1;
  assign new_y_mux_key6_and_0 = n290 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6_and_1 = new_U247 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6 = new_y_mux_key6_and_0 | new_y_mux_key6_and_1;
  assign new_y_mux_key7_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_1 = new_U247 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7 = new_y_mux_key7_and_0 | new_y_mux_key7_and_1;
  assign new_y_mux_key8_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key8_and_1 = new_U247 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8 = new_y_mux_key8_and_0 | new_y_mux_key8_and_1;
  assign new_y_mux_key9_and_0 = n290 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_1 = new_U247 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9 = new_y_mux_key9_and_0 | new_y_mux_key9_and_1;
  assign new_y_mux_key10_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key10_and_1 = new_U247 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10 = new_y_mux_key10_and_0 | new_y_mux_key10_and_1;
  assign new_y_mux_key11_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11_and_1 = new_U247 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11 = new_y_mux_key11_and_0 | new_y_mux_key11_and_1;
  assign new_y_mux_key12_and_0 = n290 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key12_and_1 = new_U247 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12 = new_y_mux_key12_and_0 | new_y_mux_key12_and_1;
  assign new_y_mux_key13_and_0 = n290 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key13_and_1 = new_U247 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key13 = new_y_mux_key13_and_0 | new_y_mux_key13_and_1;
  assign new_y_mux_key14_and_0 = n290 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14_and_1 = new_U247 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14 = new_y_mux_key14_and_0 | new_y_mux_key14_and_1;
  assign new_y_mux_key15_and_0 = n290 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key15_and_1 = new_U247 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15 = new_y_mux_key15_and_0 | new_y_mux_key15_and_1;
  assign new__state_1 = new_count_state_1;
  assign new__state_2 = new_count_state_2;
  assign new__state_3 = new_count_state_3;
  assign new__state_4 = new_count_state_4;
  assign new__state_5 = new_count_state_5;
  assign new__state_6 = new_count_state_6;
  assign new__state_7 = new_count_state_7;
  assign new__state_8 = new_count_state_8;
  assign new__state_9 = new_count_state_9;
  assign new__state_10 = new_count_state_10;
  assign new__state_11 = new_count_state_11;
  assign new__state_12 = new_count_state_12;
  assign new__state_13 = new_count_state_13;
  assign new__state_14 = new_count_state_14;
  assign new__state_15 = new_count_state_15;
  assign new__state_17 = new__state_2 | new__state_3;
  assign new__state_18 = new__state_4 | new__state_5;
  assign new__state_19 = new__state_6 | new__state_7;
  assign new__state_20 = new__state_8 | new__state_9;
  assign new__state_21 = new__state_10 | new__state_11;
  assign new__state_22 = new__state_12 | new__state_13;
  assign new__state_23 = new__state_14 | new__state_15;
  assign new__state_25 = new__state_18 | new__state_19;
  assign new__state_26 = new__state_20 | new__state_21;
  assign new__state_27 = new__state_22 | new__state_23;
  assign new__state_29 = new__state_26 | new__state_27;
  assign new_s__state_1 = new__state_1;
  assign new_not_s__state_1 = ~new_s__state_1;
  assign new_I0__state_1 = new_y_mux_key0;
  assign new_I1__state_1 = new_y_mux_key1;
  assign new_and_mux__state_1 = new_not_s__state_1 & new_I0__state_1;
  assign new_and_mux__state_1_2 = new_s__state_1 & new_I1__state_1;
  assign new_y_mux_16 = new_and_mux__state_1 | new_and_mux__state_1_2;
  assign new_s__state_3 = new__state_3;
  assign new_not_s__state_3 = ~new_s__state_3;
  assign new_I0__state_3 = new_y_mux_key2;
  assign new_I1__state_3 = new_y_mux_key3;
  assign new_and_mux__state_3 = new_not_s__state_3 & new_I0__state_3;
  assign new_and_mux__state_3_2 = new_s__state_3 & new_I1__state_3;
  assign new_y_mux_17 = new_and_mux__state_3 | new_and_mux__state_3_2;
  assign new_s__state_5 = new__state_5;
  assign new_not_s__state_5 = ~new_s__state_5;
  assign new_I0__state_5 = new_y_mux_key4;
  assign new_I1__state_5 = new_y_mux_key5;
  assign new_and_mux__state_5 = new_not_s__state_5 & new_I0__state_5;
  assign new_and_mux__state_5_2 = new_s__state_5 & new_I1__state_5;
  assign new_y_mux_18 = new_and_mux__state_5 | new_and_mux__state_5_2;
  assign new_s__state_7 = new__state_7;
  assign new_not_s__state_7 = ~new_s__state_7;
  assign new_I0__state_7 = new_y_mux_key6;
  assign new_I1__state_7 = new_y_mux_key7;
  assign new_and_mux__state_7 = new_not_s__state_7 & new_I0__state_7;
  assign new_and_mux__state_7_2 = new_s__state_7 & new_I1__state_7;
  assign new_y_mux_19 = new_and_mux__state_7 | new_and_mux__state_7_2;
  assign new_s__state_9 = new__state_9;
  assign new_not_s__state_9 = ~new_s__state_9;
  assign new_I0__state_9 = new_y_mux_key8;
  assign new_I1__state_9 = new_y_mux_key9;
  assign new_and_mux__state_9 = new_not_s__state_9 & new_I0__state_9;
  assign new_and_mux__state_9_2 = new_s__state_9 & new_I1__state_9;
  assign new_y_mux_20 = new_and_mux__state_9 | new_and_mux__state_9_2;
  assign new_s__state_11 = new__state_11;
  assign new_not_s__state_11 = ~new_s__state_11;
  assign new_I0__state_11 = new_y_mux_key10;
  assign new_I1__state_11 = new_y_mux_key11;
  assign new_and_mux__state_11 = new_not_s__state_11 & new_I0__state_11;
  assign new_and_mux__state_11_2 = new_s__state_11 & new_I1__state_11;
  assign new_y_mux_21 = new_and_mux__state_11 | new_and_mux__state_11_2;
  assign new_s__state_13 = new__state_13;
  assign new_not_s__state_13 = ~new_s__state_13;
  assign new_I0__state_13 = new_y_mux_key12;
  assign new_I1__state_13 = new_y_mux_key13;
  assign new_and_mux__state_13 = new_not_s__state_13 & new_I0__state_13;
  assign new_and_mux__state_13_2 = new_s__state_13 & new_I1__state_13;
  assign new_y_mux_22 = new_and_mux__state_13 | new_and_mux__state_13_2;
  assign new_s__state_15 = new__state_15;
  assign new_not_s__state_15 = ~new_s__state_15;
  assign new_I0__state_15 = new_y_mux_key14;
  assign new_I1__state_15 = new_y_mux_key15;
  assign new_and_mux__state_15 = new_not_s__state_15 & new_I0__state_15;
  assign new_and_mux__state_15_2 = new_s__state_15 & new_I1__state_15;
  assign new_y_mux_23 = new_and_mux__state_15 | new_and_mux__state_15_2;
  assign new_s__state_17 = new__state_17;
  assign new_not_s__state_17 = ~new_s__state_17;
  assign new_I0__state_17 = new_y_mux_16;
  assign new_I1__state_17 = new_y_mux_17;
  assign new_and_mux__state_17 = new_not_s__state_17 & new_I0__state_17;
  assign new_and_mux__state_17_2 = new_s__state_17 & new_I1__state_17;
  assign new_y_mux_24 = new_and_mux__state_17 | new_and_mux__state_17_2;
  assign new_s__state_19 = new__state_19;
  assign new_not_s__state_19 = ~new_s__state_19;
  assign new_I0__state_19 = new_y_mux_18;
  assign new_I1__state_19 = new_y_mux_19;
  assign new_and_mux__state_19 = new_not_s__state_19 & new_I0__state_19;
  assign new_and_mux__state_19_2 = new_s__state_19 & new_I1__state_19;
  assign new_y_mux_25 = new_and_mux__state_19 | new_and_mux__state_19_2;
  assign new_s__state_21 = new__state_21;
  assign new_not_s__state_21 = ~new_s__state_21;
  assign new_I0__state_21 = new_y_mux_20;
  assign new_I1__state_21 = new_y_mux_21;
  assign new_and_mux__state_21 = new_not_s__state_21 & new_I0__state_21;
  assign new_and_mux__state_21_2 = new_s__state_21 & new_I1__state_21;
  assign new_y_mux_26 = new_and_mux__state_21 | new_and_mux__state_21_2;
  assign new_s__state_23 = new__state_23;
  assign new_not_s__state_23 = ~new_s__state_23;
  assign new_I0__state_23 = new_y_mux_22;
  assign new_I1__state_23 = new_y_mux_23;
  assign new_and_mux__state_23 = new_not_s__state_23 & new_I0__state_23;
  assign new_and_mux__state_23_2 = new_s__state_23 & new_I1__state_23;
  assign new_y_mux_27 = new_and_mux__state_23 | new_and_mux__state_23_2;
  assign new_s__state_25 = new__state_25;
  assign new_not_s__state_25 = ~new_s__state_25;
  assign new_I0__state_25 = new_y_mux_24;
  assign new_I1__state_25 = new_y_mux_25;
  assign new_and_mux__state_25 = new_not_s__state_25 & new_I0__state_25;
  assign new_and_mux__state_25_2 = new_s__state_25 & new_I1__state_25;
  assign new_y_mux_28 = new_and_mux__state_25 | new_and_mux__state_25_2;
  assign new_s__state_27 = new__state_27;
  assign new_not_s__state_27 = ~new_s__state_27;
  assign new_I0__state_27 = new_y_mux_26;
  assign new_I1__state_27 = new_y_mux_27;
  assign new_and_mux__state_27 = new_not_s__state_27 & new_I0__state_27;
  assign new_and_mux__state_27_2 = new_s__state_27 & new_I1__state_27;
  assign new_y_mux_29 = new_and_mux__state_27 | new_and_mux__state_27_2;
  assign new_s__state_29 = new__state_29;
  assign new_not_s__state_29 = ~new_s__state_29;
  assign new_I0__state_29 = new_y_mux_28;
  assign new_I1__state_29 = new_y_mux_29;
  assign new_and_mux__state_29 = new_not_s__state_29 & new_I0__state_29;
  assign new_and_mux__state_29_2 = new_s__state_29 & new_I1__state_29;
  assign n280 = new_and_mux__state_29 | new_and_mux__state_29_2;
  always @ (posedge clock) begin
    BUF1_REG_0_ <= n280;
    BUF1_REG_1_ <= n285;
    BUF1_REG_2_ <= n290;
    BUF1_REG_3_ <= n295;
    BUF1_REG_4_ <= n300;
    BUF1_REG_5_ <= n305;
    BUF1_REG_6_ <= n310;
    BUF1_REG_7_ <= n315;
    BUF1_REG_8_ <= n320;
    BUF1_REG_9_ <= n325;
    BUF1_REG_10_ <= n330;
    BUF1_REG_11_ <= n335;
    BUF1_REG_12_ <= n340;
    BUF1_REG_13_ <= n345;
    BUF1_REG_14_ <= n350;
    BUF1_REG_15_ <= n355;
    BUF1_REG_16_ <= n360;
    BUF1_REG_17_ <= n365;
    BUF1_REG_18_ <= n370;
    BUF1_REG_19_ <= n375;
    BUF1_REG_20_ <= n380;
    BUF1_REG_21_ <= n385;
    BUF1_REG_22_ <= n390;
    BUF1_REG_23_ <= n395;
    BUF1_REG_24_ <= n400;
    BUF1_REG_25_ <= n405;
    BUF1_REG_26_ <= n410;
    BUF1_REG_27_ <= n415;
    BUF1_REG_28_ <= n420;
    BUF1_REG_29_ <= n425;
    BUF1_REG_30_ <= n430;
    BUF1_REG_31_ <= n435;
    BUF2_REG_0_ <= n440;
    BUF2_REG_1_ <= n445;
    BUF2_REG_2_ <= n450;
    BUF2_REG_3_ <= n455;
    BUF2_REG_4_ <= n460;
    BUF2_REG_5_ <= n465;
    BUF2_REG_6_ <= n470;
    BUF2_REG_7_ <= n475;
    BUF2_REG_8_ <= n480;
    BUF2_REG_9_ <= n485;
    BUF2_REG_10_ <= n490;
    BUF2_REG_11_ <= n495;
    BUF2_REG_12_ <= n500;
    BUF2_REG_13_ <= n505;
    BUF2_REG_14_ <= n510;
    BUF2_REG_15_ <= n515;
    BUF2_REG_16_ <= n520;
    BUF2_REG_17_ <= n525;
    BUF2_REG_18_ <= n530;
    BUF2_REG_19_ <= n535;
    BUF2_REG_20_ <= n540;
    BUF2_REG_21_ <= n545;
    BUF2_REG_22_ <= n550;
    BUF2_REG_23_ <= n555;
    BUF2_REG_24_ <= n560;
    BUF2_REG_25_ <= n565;
    BUF2_REG_26_ <= n570;
    BUF2_REG_27_ <= n575;
    BUF2_REG_28_ <= n580;
    BUF2_REG_29_ <= n585;
    BUF2_REG_30_ <= n590;
    BUF2_REG_31_ <= n595;
    READY12_REG <= n600;
    READY21_REG <= n605;
    READY22_REG <= n610;
    READY11_REG <= n615;
    P3_BE_N_REG_3_ <= n620;
    P3_BE_N_REG_2_ <= n625;
    P3_BE_N_REG_1_ <= n630;
    P3_BE_N_REG_0_ <= n635;
    P3_ADDRESS_REG_29_ <= n640;
    P3_ADDRESS_REG_28_ <= n645;
    P3_ADDRESS_REG_27_ <= n650;
    P3_ADDRESS_REG_26_ <= n655;
    P3_ADDRESS_REG_25_ <= n660;
    P3_ADDRESS_REG_24_ <= n665;
    P3_ADDRESS_REG_23_ <= n670;
    P3_ADDRESS_REG_22_ <= n675;
    P3_ADDRESS_REG_21_ <= n680;
    P3_ADDRESS_REG_20_ <= n685;
    P3_ADDRESS_REG_19_ <= n690;
    P3_ADDRESS_REG_18_ <= n695;
    P3_ADDRESS_REG_17_ <= n700;
    P3_ADDRESS_REG_16_ <= n705;
    P3_ADDRESS_REG_15_ <= n710;
    P3_ADDRESS_REG_14_ <= n715;
    P3_ADDRESS_REG_13_ <= n720;
    P3_ADDRESS_REG_12_ <= n725;
    P3_ADDRESS_REG_11_ <= n730;
    P3_ADDRESS_REG_10_ <= n735;
    P3_ADDRESS_REG_9_ <= n740;
    P3_ADDRESS_REG_8_ <= n745;
    P3_ADDRESS_REG_7_ <= n750;
    P3_ADDRESS_REG_6_ <= n755;
    P3_ADDRESS_REG_5_ <= n760;
    P3_ADDRESS_REG_4_ <= n765;
    P3_ADDRESS_REG_3_ <= n770;
    P3_ADDRESS_REG_2_ <= n775;
    P3_ADDRESS_REG_1_ <= n780;
    P3_ADDRESS_REG_0_ <= n785;
    P3_STATE_REG_2_ <= n790;
    P3_STATE_REG_1_ <= n795;
    P3_STATE_REG_0_ <= n800;
    P3_DATAWIDTH_REG_0_ <= n805;
    P3_DATAWIDTH_REG_1_ <= n810;
    P3_DATAWIDTH_REG_2_ <= n815;
    P3_DATAWIDTH_REG_3_ <= n820;
    P3_DATAWIDTH_REG_4_ <= n825;
    P3_DATAWIDTH_REG_5_ <= n830;
    P3_DATAWIDTH_REG_6_ <= n835;
    P3_DATAWIDTH_REG_7_ <= n840;
    P3_DATAWIDTH_REG_8_ <= n845;
    P3_DATAWIDTH_REG_9_ <= n850;
    P3_DATAWIDTH_REG_10_ <= n855;
    P3_DATAWIDTH_REG_11_ <= n860;
    P3_DATAWIDTH_REG_12_ <= n865;
    P3_DATAWIDTH_REG_13_ <= n870;
    P3_DATAWIDTH_REG_14_ <= n875;
    P3_DATAWIDTH_REG_15_ <= n880;
    P3_DATAWIDTH_REG_16_ <= n885;
    P3_DATAWIDTH_REG_17_ <= n890;
    P3_DATAWIDTH_REG_18_ <= n895;
    P3_DATAWIDTH_REG_19_ <= n900;
    P3_DATAWIDTH_REG_20_ <= n905;
    P3_DATAWIDTH_REG_21_ <= n910;
    P3_DATAWIDTH_REG_22_ <= n915;
    P3_DATAWIDTH_REG_23_ <= n920;
    P3_DATAWIDTH_REG_24_ <= n925;
    P3_DATAWIDTH_REG_25_ <= n930;
    P3_DATAWIDTH_REG_26_ <= n935;
    P3_DATAWIDTH_REG_27_ <= n940;
    P3_DATAWIDTH_REG_28_ <= n945;
    P3_DATAWIDTH_REG_29_ <= n950;
    P3_DATAWIDTH_REG_30_ <= n955;
    P3_DATAWIDTH_REG_31_ <= n960;
    P3_STATE2_REG_3_ <= n965;
    P3_STATE2_REG_2_ <= n970;
    P3_STATE2_REG_1_ <= n975;
    P3_STATE2_REG_0_ <= n980;
    P3_INSTQUEUE_REG_15__7_ <= n985;
    P3_INSTQUEUE_REG_15__6_ <= n990;
    P3_INSTQUEUE_REG_15__5_ <= n995;
    P3_INSTQUEUE_REG_15__4_ <= n1000;
    P3_INSTQUEUE_REG_15__3_ <= n1005;
    P3_INSTQUEUE_REG_15__2_ <= n1010;
    P3_INSTQUEUE_REG_15__1_ <= n1015;
    P3_INSTQUEUE_REG_15__0_ <= n1020;
    P3_INSTQUEUE_REG_14__7_ <= n1025;
    P3_INSTQUEUE_REG_14__6_ <= n1030;
    P3_INSTQUEUE_REG_14__5_ <= n1035;
    P3_INSTQUEUE_REG_14__4_ <= n1040;
    P3_INSTQUEUE_REG_14__3_ <= n1045;
    P3_INSTQUEUE_REG_14__2_ <= n1050;
    P3_INSTQUEUE_REG_14__1_ <= n1055;
    P3_INSTQUEUE_REG_14__0_ <= n1060;
    P3_INSTQUEUE_REG_13__7_ <= n1065;
    P3_INSTQUEUE_REG_13__6_ <= n1070;
    P3_INSTQUEUE_REG_13__5_ <= n1075;
    P3_INSTQUEUE_REG_13__4_ <= n1080;
    P3_INSTQUEUE_REG_13__3_ <= n1085;
    P3_INSTQUEUE_REG_13__2_ <= n1090;
    P3_INSTQUEUE_REG_13__1_ <= n1095;
    P3_INSTQUEUE_REG_13__0_ <= n1100;
    P3_INSTQUEUE_REG_12__7_ <= n1105;
    P3_INSTQUEUE_REG_12__6_ <= n1110;
    P3_INSTQUEUE_REG_12__5_ <= n1115;
    P3_INSTQUEUE_REG_12__4_ <= n1120;
    P3_INSTQUEUE_REG_12__3_ <= n1125;
    P3_INSTQUEUE_REG_12__2_ <= n1130;
    P3_INSTQUEUE_REG_12__1_ <= n1135;
    P3_INSTQUEUE_REG_12__0_ <= n1140;
    P3_INSTQUEUE_REG_11__7_ <= n1145;
    P3_INSTQUEUE_REG_11__6_ <= n1150;
    P3_INSTQUEUE_REG_11__5_ <= n1155;
    P3_INSTQUEUE_REG_11__4_ <= n1160;
    P3_INSTQUEUE_REG_11__3_ <= n1165;
    P3_INSTQUEUE_REG_11__2_ <= n1170;
    P3_INSTQUEUE_REG_11__1_ <= n1175;
    P3_INSTQUEUE_REG_11__0_ <= n1180;
    P3_INSTQUEUE_REG_10__7_ <= n1185;
    P3_INSTQUEUE_REG_10__6_ <= n1190;
    P3_INSTQUEUE_REG_10__5_ <= n1195;
    P3_INSTQUEUE_REG_10__4_ <= n1200;
    P3_INSTQUEUE_REG_10__3_ <= n1205;
    P3_INSTQUEUE_REG_10__2_ <= n1210;
    P3_INSTQUEUE_REG_10__1_ <= n1215;
    P3_INSTQUEUE_REG_10__0_ <= n1220;
    P3_INSTQUEUE_REG_9__7_ <= n1225;
    P3_INSTQUEUE_REG_9__6_ <= n1230;
    P3_INSTQUEUE_REG_9__5_ <= n1235;
    P3_INSTQUEUE_REG_9__4_ <= n1240;
    P3_INSTQUEUE_REG_9__3_ <= n1245;
    P3_INSTQUEUE_REG_9__2_ <= n1250;
    P3_INSTQUEUE_REG_9__1_ <= n1255;
    P3_INSTQUEUE_REG_9__0_ <= n1260;
    P3_INSTQUEUE_REG_8__7_ <= n1265;
    P3_INSTQUEUE_REG_8__6_ <= n1270;
    P3_INSTQUEUE_REG_8__5_ <= n1275;
    P3_INSTQUEUE_REG_8__4_ <= n1280;
    P3_INSTQUEUE_REG_8__3_ <= n1285;
    P3_INSTQUEUE_REG_8__2_ <= n1290;
    P3_INSTQUEUE_REG_8__1_ <= n1295;
    P3_INSTQUEUE_REG_8__0_ <= n1300;
    P3_INSTQUEUE_REG_7__7_ <= n1305;
    P3_INSTQUEUE_REG_7__6_ <= n1310;
    P3_INSTQUEUE_REG_7__5_ <= n1315;
    P3_INSTQUEUE_REG_7__4_ <= n1320;
    P3_INSTQUEUE_REG_7__3_ <= n1325;
    P3_INSTQUEUE_REG_7__2_ <= n1330;
    P3_INSTQUEUE_REG_7__1_ <= n1335;
    P3_INSTQUEUE_REG_7__0_ <= n1340;
    P3_INSTQUEUE_REG_6__7_ <= n1345;
    P3_INSTQUEUE_REG_6__6_ <= n1350;
    P3_INSTQUEUE_REG_6__5_ <= n1355;
    P3_INSTQUEUE_REG_6__4_ <= n1360;
    P3_INSTQUEUE_REG_6__3_ <= n1365;
    P3_INSTQUEUE_REG_6__2_ <= n1370;
    P3_INSTQUEUE_REG_6__1_ <= n1375;
    P3_INSTQUEUE_REG_6__0_ <= n1380;
    P3_INSTQUEUE_REG_5__7_ <= n1385;
    P3_INSTQUEUE_REG_5__6_ <= n1390;
    P3_INSTQUEUE_REG_5__5_ <= n1395;
    P3_INSTQUEUE_REG_5__4_ <= n1400;
    P3_INSTQUEUE_REG_5__3_ <= n1405;
    P3_INSTQUEUE_REG_5__2_ <= n1410;
    P3_INSTQUEUE_REG_5__1_ <= n1415;
    P3_INSTQUEUE_REG_5__0_ <= n1420;
    P3_INSTQUEUE_REG_4__7_ <= n1425;
    P3_INSTQUEUE_REG_4__6_ <= n1430;
    P3_INSTQUEUE_REG_4__5_ <= n1435;
    P3_INSTQUEUE_REG_4__4_ <= n1440;
    P3_INSTQUEUE_REG_4__3_ <= n1445;
    P3_INSTQUEUE_REG_4__2_ <= n1450;
    P3_INSTQUEUE_REG_4__1_ <= n1455;
    P3_INSTQUEUE_REG_4__0_ <= n1460;
    P3_INSTQUEUE_REG_3__7_ <= n1465;
    P3_INSTQUEUE_REG_3__6_ <= n1470;
    P3_INSTQUEUE_REG_3__5_ <= n1475;
    P3_INSTQUEUE_REG_3__4_ <= n1480;
    P3_INSTQUEUE_REG_3__3_ <= n1485;
    P3_INSTQUEUE_REG_3__2_ <= n1490;
    P3_INSTQUEUE_REG_3__1_ <= n1495;
    P3_INSTQUEUE_REG_3__0_ <= n1500;
    P3_INSTQUEUE_REG_2__7_ <= n1505;
    P3_INSTQUEUE_REG_2__6_ <= n1510;
    P3_INSTQUEUE_REG_2__5_ <= n1515;
    P3_INSTQUEUE_REG_2__4_ <= n1520;
    P3_INSTQUEUE_REG_2__3_ <= n1525;
    P3_INSTQUEUE_REG_2__2_ <= n1530;
    P3_INSTQUEUE_REG_2__1_ <= n1535;
    P3_INSTQUEUE_REG_2__0_ <= n1540;
    P3_INSTQUEUE_REG_1__7_ <= n1545;
    P3_INSTQUEUE_REG_1__6_ <= n1550;
    P3_INSTQUEUE_REG_1__5_ <= n1555;
    P3_INSTQUEUE_REG_1__4_ <= n1560;
    P3_INSTQUEUE_REG_1__3_ <= n1565;
    P3_INSTQUEUE_REG_1__2_ <= n1570;
    P3_INSTQUEUE_REG_1__1_ <= n1575;
    P3_INSTQUEUE_REG_1__0_ <= n1580;
    P3_INSTQUEUE_REG_0__7_ <= n1585;
    P3_INSTQUEUE_REG_0__6_ <= n1590;
    P3_INSTQUEUE_REG_0__5_ <= n1595;
    P3_INSTQUEUE_REG_0__4_ <= n1600;
    P3_INSTQUEUE_REG_0__3_ <= n1605;
    P3_INSTQUEUE_REG_0__2_ <= n1610;
    P3_INSTQUEUE_REG_0__1_ <= n1615;
    P3_INSTQUEUE_REG_0__0_ <= n1620;
    P3_INSTQUEUERD_ADDR_REG_4_ <= n1625;
    P3_INSTQUEUERD_ADDR_REG_3_ <= n1630;
    P3_INSTQUEUERD_ADDR_REG_2_ <= n1635;
    P3_INSTQUEUERD_ADDR_REG_1_ <= n1640;
    P3_INSTQUEUERD_ADDR_REG_0_ <= n1645;
    P3_INSTQUEUEWR_ADDR_REG_4_ <= n1650;
    P3_INSTQUEUEWR_ADDR_REG_3_ <= n1655;
    P3_INSTQUEUEWR_ADDR_REG_2_ <= n1660;
    P3_INSTQUEUEWR_ADDR_REG_1_ <= n1665;
    P3_INSTQUEUEWR_ADDR_REG_0_ <= n1670;
    P3_INSTADDRPOINTER_REG_0_ <= n1675;
    P3_INSTADDRPOINTER_REG_1_ <= n1680;
    P3_INSTADDRPOINTER_REG_2_ <= n1685;
    P3_INSTADDRPOINTER_REG_3_ <= n1690;
    P3_INSTADDRPOINTER_REG_4_ <= n1695;
    P3_INSTADDRPOINTER_REG_5_ <= n1700;
    P3_INSTADDRPOINTER_REG_6_ <= n1705;
    P3_INSTADDRPOINTER_REG_7_ <= n1710;
    P3_INSTADDRPOINTER_REG_8_ <= n1715;
    P3_INSTADDRPOINTER_REG_9_ <= n1720;
    P3_INSTADDRPOINTER_REG_10_ <= n1725;
    P3_INSTADDRPOINTER_REG_11_ <= n1730;
    P3_INSTADDRPOINTER_REG_12_ <= n1735;
    P3_INSTADDRPOINTER_REG_13_ <= n1740;
    P3_INSTADDRPOINTER_REG_14_ <= n1745;
    P3_INSTADDRPOINTER_REG_15_ <= n1750;
    P3_INSTADDRPOINTER_REG_16_ <= n1755;
    P3_INSTADDRPOINTER_REG_17_ <= n1760;
    P3_INSTADDRPOINTER_REG_18_ <= n1765;
    P3_INSTADDRPOINTER_REG_19_ <= n1770;
    P3_INSTADDRPOINTER_REG_20_ <= n1775;
    P3_INSTADDRPOINTER_REG_21_ <= n1780;
    P3_INSTADDRPOINTER_REG_22_ <= n1785;
    P3_INSTADDRPOINTER_REG_23_ <= n1790;
    P3_INSTADDRPOINTER_REG_24_ <= n1795;
    P3_INSTADDRPOINTER_REG_25_ <= n1800;
    P3_INSTADDRPOINTER_REG_26_ <= n1805;
    P3_INSTADDRPOINTER_REG_27_ <= n1810;
    P3_INSTADDRPOINTER_REG_28_ <= n1815;
    P3_INSTADDRPOINTER_REG_29_ <= n1820;
    P3_INSTADDRPOINTER_REG_30_ <= n1825;
    P3_INSTADDRPOINTER_REG_31_ <= n1830;
    P3_PHYADDRPOINTER_REG_0_ <= n1835;
    P3_PHYADDRPOINTER_REG_1_ <= n1840;
    P3_PHYADDRPOINTER_REG_2_ <= n1845;
    P3_PHYADDRPOINTER_REG_3_ <= n1850;
    P3_PHYADDRPOINTER_REG_4_ <= n1855;
    P3_PHYADDRPOINTER_REG_5_ <= n1860;
    P3_PHYADDRPOINTER_REG_6_ <= n1865;
    P3_PHYADDRPOINTER_REG_7_ <= n1870;
    P3_PHYADDRPOINTER_REG_8_ <= n1875;
    P3_PHYADDRPOINTER_REG_9_ <= n1880;
    P3_PHYADDRPOINTER_REG_10_ <= n1885;
    P3_PHYADDRPOINTER_REG_11_ <= n1890;
    P3_PHYADDRPOINTER_REG_12_ <= n1895;
    P3_PHYADDRPOINTER_REG_13_ <= n1900;
    P3_PHYADDRPOINTER_REG_14_ <= n1905;
    P3_PHYADDRPOINTER_REG_15_ <= n1910;
    P3_PHYADDRPOINTER_REG_16_ <= n1915;
    P3_PHYADDRPOINTER_REG_17_ <= n1920;
    P3_PHYADDRPOINTER_REG_18_ <= n1925;
    P3_PHYADDRPOINTER_REG_19_ <= n1930;
    P3_PHYADDRPOINTER_REG_20_ <= n1935;
    P3_PHYADDRPOINTER_REG_21_ <= n1940;
    P3_PHYADDRPOINTER_REG_22_ <= n1945;
    P3_PHYADDRPOINTER_REG_23_ <= n1950;
    P3_PHYADDRPOINTER_REG_24_ <= n1955;
    P3_PHYADDRPOINTER_REG_25_ <= n1960;
    P3_PHYADDRPOINTER_REG_26_ <= n1965;
    P3_PHYADDRPOINTER_REG_27_ <= n1970;
    P3_PHYADDRPOINTER_REG_28_ <= n1975;
    P3_PHYADDRPOINTER_REG_29_ <= n1980;
    P3_PHYADDRPOINTER_REG_30_ <= n1985;
    P3_PHYADDRPOINTER_REG_31_ <= n1990;
    P3_LWORD_REG_15_ <= n1995;
    P3_LWORD_REG_14_ <= n2000;
    P3_LWORD_REG_13_ <= n2005;
    P3_LWORD_REG_12_ <= n2010;
    P3_LWORD_REG_11_ <= n2015;
    P3_LWORD_REG_10_ <= n2020;
    P3_LWORD_REG_9_ <= n2025;
    P3_LWORD_REG_8_ <= n2030;
    P3_LWORD_REG_7_ <= n2035;
    P3_LWORD_REG_6_ <= n2040;
    P3_LWORD_REG_5_ <= n2045;
    P3_LWORD_REG_4_ <= n2050;
    P3_LWORD_REG_3_ <= n2055;
    P3_LWORD_REG_2_ <= n2060;
    P3_LWORD_REG_1_ <= n2065;
    P3_LWORD_REG_0_ <= n2070;
    P3_UWORD_REG_14_ <= n2075;
    P3_UWORD_REG_13_ <= n2080;
    P3_UWORD_REG_12_ <= n2085;
    P3_UWORD_REG_11_ <= n2090;
    P3_UWORD_REG_10_ <= n2095;
    P3_UWORD_REG_9_ <= n2100;
    P3_UWORD_REG_8_ <= n2105;
    P3_UWORD_REG_7_ <= n2110;
    P3_UWORD_REG_6_ <= n2115;
    P3_UWORD_REG_5_ <= n2120;
    P3_UWORD_REG_4_ <= n2125;
    P3_UWORD_REG_3_ <= n2130;
    P3_UWORD_REG_2_ <= n2135;
    P3_UWORD_REG_1_ <= n2140;
    P3_UWORD_REG_0_ <= n2145;
    P3_DATAO_REG_0_ <= n2150;
    P3_DATAO_REG_1_ <= n2154;
    P3_DATAO_REG_2_ <= n2158;
    P3_DATAO_REG_3_ <= n2162;
    P3_DATAO_REG_4_ <= n2166;
    P3_DATAO_REG_5_ <= n2170;
    P3_DATAO_REG_6_ <= n2174;
    P3_DATAO_REG_7_ <= n2178;
    P3_DATAO_REG_8_ <= n2182;
    P3_DATAO_REG_9_ <= n2186;
    P3_DATAO_REG_10_ <= n2190;
    P3_DATAO_REG_11_ <= n2194;
    P3_DATAO_REG_12_ <= n2198;
    P3_DATAO_REG_13_ <= n2202;
    P3_DATAO_REG_14_ <= n2206;
    P3_DATAO_REG_15_ <= n2210;
    P3_DATAO_REG_16_ <= n2214;
    P3_DATAO_REG_17_ <= n2218;
    P3_DATAO_REG_18_ <= n2222;
    P3_DATAO_REG_19_ <= n2226;
    P3_DATAO_REG_20_ <= n2230;
    P3_DATAO_REG_21_ <= n2234;
    P3_DATAO_REG_22_ <= n2238;
    P3_DATAO_REG_23_ <= n2242;
    P3_DATAO_REG_24_ <= n2246;
    P3_DATAO_REG_25_ <= n2250;
    P3_DATAO_REG_26_ <= n2254;
    P3_DATAO_REG_27_ <= n2258;
    P3_DATAO_REG_28_ <= n2262;
    P3_DATAO_REG_29_ <= n2266;
    P3_DATAO_REG_30_ <= n2270;
    P3_DATAO_REG_31_ <= n2274;
    P3_EAX_REG_0_ <= n2278;
    P3_EAX_REG_1_ <= n2283;
    P3_EAX_REG_2_ <= n2288;
    P3_EAX_REG_3_ <= n2293;
    P3_EAX_REG_4_ <= n2298;
    P3_EAX_REG_5_ <= n2303;
    P3_EAX_REG_6_ <= n2308;
    P3_EAX_REG_7_ <= n2313;
    P3_EAX_REG_8_ <= n2318;
    P3_EAX_REG_9_ <= n2323;
    P3_EAX_REG_10_ <= n2328;
    P3_EAX_REG_11_ <= n2333;
    P3_EAX_REG_12_ <= n2338;
    P3_EAX_REG_13_ <= n2343;
    P3_EAX_REG_14_ <= n2348;
    P3_EAX_REG_15_ <= n2353;
    P3_EAX_REG_16_ <= n2358;
    P3_EAX_REG_17_ <= n2363;
    P3_EAX_REG_18_ <= n2368;
    P3_EAX_REG_19_ <= n2373;
    P3_EAX_REG_20_ <= n2378;
    P3_EAX_REG_21_ <= n2383;
    P3_EAX_REG_22_ <= n2388;
    P3_EAX_REG_23_ <= n2393;
    P3_EAX_REG_24_ <= n2398;
    P3_EAX_REG_25_ <= n2403;
    P3_EAX_REG_26_ <= n2408;
    P3_EAX_REG_27_ <= n2413;
    P3_EAX_REG_28_ <= n2418;
    P3_EAX_REG_29_ <= n2423;
    P3_EAX_REG_30_ <= n2428;
    P3_EAX_REG_31_ <= n2433;
    P3_EBX_REG_0_ <= n2438;
    P3_EBX_REG_1_ <= n2443;
    P3_EBX_REG_2_ <= n2448;
    P3_EBX_REG_3_ <= n2453;
    P3_EBX_REG_4_ <= n2458;
    P3_EBX_REG_5_ <= n2463;
    P3_EBX_REG_6_ <= n2468;
    P3_EBX_REG_7_ <= n2473;
    P3_EBX_REG_8_ <= n2478;
    P3_EBX_REG_9_ <= n2483;
    P3_EBX_REG_10_ <= n2488;
    P3_EBX_REG_11_ <= n2493;
    P3_EBX_REG_12_ <= n2498;
    P3_EBX_REG_13_ <= n2503;
    P3_EBX_REG_14_ <= n2508;
    P3_EBX_REG_15_ <= n2513;
    P3_EBX_REG_16_ <= n2518;
    P3_EBX_REG_17_ <= n2523;
    P3_EBX_REG_18_ <= n2528;
    P3_EBX_REG_19_ <= n2533;
    P3_EBX_REG_20_ <= n2538;
    P3_EBX_REG_21_ <= n2543;
    P3_EBX_REG_22_ <= n2548;
    P3_EBX_REG_23_ <= n2553;
    P3_EBX_REG_24_ <= n2558;
    P3_EBX_REG_25_ <= n2563;
    P3_EBX_REG_26_ <= n2568;
    P3_EBX_REG_27_ <= n2573;
    P3_EBX_REG_28_ <= n2578;
    P3_EBX_REG_29_ <= n2583;
    P3_EBX_REG_30_ <= n2588;
    P3_EBX_REG_31_ <= n2593;
    P3_REIP_REG_0_ <= n2598;
    P3_REIP_REG_1_ <= n2603;
    P3_REIP_REG_2_ <= n2608;
    P3_REIP_REG_3_ <= n2613;
    P3_REIP_REG_4_ <= n2618;
    P3_REIP_REG_5_ <= n2623;
    P3_REIP_REG_6_ <= n2628;
    P3_REIP_REG_7_ <= n2633;
    P3_REIP_REG_8_ <= n2638;
    P3_REIP_REG_9_ <= n2643;
    P3_REIP_REG_10_ <= n2648;
    P3_REIP_REG_11_ <= n2653;
    P3_REIP_REG_12_ <= n2658;
    P3_REIP_REG_13_ <= n2663;
    P3_REIP_REG_14_ <= n2668;
    P3_REIP_REG_15_ <= n2673;
    P3_REIP_REG_16_ <= n2678;
    P3_REIP_REG_17_ <= n2683;
    P3_REIP_REG_18_ <= n2688;
    P3_REIP_REG_19_ <= n2693;
    P3_REIP_REG_20_ <= n2698;
    P3_REIP_REG_21_ <= n2703;
    P3_REIP_REG_22_ <= n2708;
    P3_REIP_REG_23_ <= n2713;
    P3_REIP_REG_24_ <= n2718;
    P3_REIP_REG_25_ <= n2723;
    P3_REIP_REG_26_ <= n2728;
    P3_REIP_REG_27_ <= n2733;
    P3_REIP_REG_28_ <= n2738;
    P3_REIP_REG_29_ <= n2743;
    P3_REIP_REG_30_ <= n2748;
    P3_REIP_REG_31_ <= n2753;
    P3_BYTEENABLE_REG_3_ <= n2758;
    P3_BYTEENABLE_REG_2_ <= n2763;
    P3_BYTEENABLE_REG_1_ <= n2768;
    P3_BYTEENABLE_REG_0_ <= n2773;
    P3_W_R_N_REG <= n2778;
    P3_FLUSH_REG <= n2782;
    P3_MORE_REG <= n2787;
    P3_STATEBS16_REG <= n2792;
    P3_REQUESTPENDING_REG <= n2797;
    P3_D_C_N_REG <= n2802;
    P3_M_IO_N_REG <= n2806;
    P3_CODEFETCH_REG <= n2810;
    P3_ADS_N_REG <= n2815;
    P3_READREQUEST_REG <= n2819;
    P3_MEMORYFETCH_REG <= n2824;
    P2_BE_N_REG_3_ <= n2829;
    P2_BE_N_REG_2_ <= n2834;
    P2_BE_N_REG_1_ <= n2839;
    P2_BE_N_REG_0_ <= n2844;
    P2_ADDRESS_REG_29_ <= n2849;
    P2_ADDRESS_REG_28_ <= n2854;
    P2_ADDRESS_REG_27_ <= n2859;
    P2_ADDRESS_REG_26_ <= n2864;
    P2_ADDRESS_REG_25_ <= n2869;
    P2_ADDRESS_REG_24_ <= n2874;
    P2_ADDRESS_REG_23_ <= n2879;
    P2_ADDRESS_REG_22_ <= n2884;
    P2_ADDRESS_REG_21_ <= n2889;
    P2_ADDRESS_REG_20_ <= n2894;
    P2_ADDRESS_REG_19_ <= n2899;
    P2_ADDRESS_REG_18_ <= n2904;
    P2_ADDRESS_REG_17_ <= n2909;
    P2_ADDRESS_REG_16_ <= n2914;
    P2_ADDRESS_REG_15_ <= n2919;
    P2_ADDRESS_REG_14_ <= n2924;
    P2_ADDRESS_REG_13_ <= n2929;
    P2_ADDRESS_REG_12_ <= n2934;
    P2_ADDRESS_REG_11_ <= n2939;
    P2_ADDRESS_REG_10_ <= n2944;
    P2_ADDRESS_REG_9_ <= n2949;
    P2_ADDRESS_REG_8_ <= n2954;
    P2_ADDRESS_REG_7_ <= n2959;
    P2_ADDRESS_REG_6_ <= n2964;
    P2_ADDRESS_REG_5_ <= n2969;
    P2_ADDRESS_REG_4_ <= n2974;
    P2_ADDRESS_REG_3_ <= n2979;
    P2_ADDRESS_REG_2_ <= n2984;
    P2_ADDRESS_REG_1_ <= n2989;
    P2_ADDRESS_REG_0_ <= n2994;
    P2_STATE_REG_2_ <= n2999;
    P2_STATE_REG_1_ <= n3004;
    P2_STATE_REG_0_ <= n3009;
    P2_DATAWIDTH_REG_0_ <= n3014;
    P2_DATAWIDTH_REG_1_ <= n3019;
    P2_DATAWIDTH_REG_2_ <= n3024;
    P2_DATAWIDTH_REG_3_ <= n3029;
    P2_DATAWIDTH_REG_4_ <= n3034;
    P2_DATAWIDTH_REG_5_ <= n3039;
    P2_DATAWIDTH_REG_6_ <= n3044;
    P2_DATAWIDTH_REG_7_ <= n3049;
    P2_DATAWIDTH_REG_8_ <= n3054;
    P2_DATAWIDTH_REG_9_ <= n3059;
    P2_DATAWIDTH_REG_10_ <= n3064;
    P2_DATAWIDTH_REG_11_ <= n3069;
    P2_DATAWIDTH_REG_12_ <= n3074;
    P2_DATAWIDTH_REG_13_ <= n3079;
    P2_DATAWIDTH_REG_14_ <= n3084;
    P2_DATAWIDTH_REG_15_ <= n3089;
    P2_DATAWIDTH_REG_16_ <= n3094;
    P2_DATAWIDTH_REG_17_ <= n3099;
    P2_DATAWIDTH_REG_18_ <= n3104;
    P2_DATAWIDTH_REG_19_ <= n3109;
    P2_DATAWIDTH_REG_20_ <= n3114;
    P2_DATAWIDTH_REG_21_ <= n3119;
    P2_DATAWIDTH_REG_22_ <= n3124;
    P2_DATAWIDTH_REG_23_ <= n3129;
    P2_DATAWIDTH_REG_24_ <= n3134;
    P2_DATAWIDTH_REG_25_ <= n3139;
    P2_DATAWIDTH_REG_26_ <= n3144;
    P2_DATAWIDTH_REG_27_ <= n3149;
    P2_DATAWIDTH_REG_28_ <= n3154;
    P2_DATAWIDTH_REG_29_ <= n3159;
    P2_DATAWIDTH_REG_30_ <= n3164;
    P2_DATAWIDTH_REG_31_ <= n3169;
    P2_STATE2_REG_3_ <= n3174;
    P2_STATE2_REG_2_ <= n3179;
    P2_STATE2_REG_1_ <= n3184;
    P2_STATE2_REG_0_ <= n3189;
    P2_INSTQUEUE_REG_15__7_ <= n3194;
    P2_INSTQUEUE_REG_15__6_ <= n3199;
    P2_INSTQUEUE_REG_15__5_ <= n3204;
    P2_INSTQUEUE_REG_15__4_ <= n3209;
    P2_INSTQUEUE_REG_15__3_ <= n3214;
    P2_INSTQUEUE_REG_15__2_ <= n3219;
    P2_INSTQUEUE_REG_15__1_ <= n3224;
    P2_INSTQUEUE_REG_15__0_ <= n3229;
    P2_INSTQUEUE_REG_14__7_ <= n3234;
    P2_INSTQUEUE_REG_14__6_ <= n3239;
    P2_INSTQUEUE_REG_14__5_ <= n3244;
    P2_INSTQUEUE_REG_14__4_ <= n3249;
    P2_INSTQUEUE_REG_14__3_ <= n3254;
    P2_INSTQUEUE_REG_14__2_ <= n3259;
    P2_INSTQUEUE_REG_14__1_ <= n3264;
    P2_INSTQUEUE_REG_14__0_ <= n3269;
    P2_INSTQUEUE_REG_13__7_ <= n3274;
    P2_INSTQUEUE_REG_13__6_ <= n3279;
    P2_INSTQUEUE_REG_13__5_ <= n3284;
    P2_INSTQUEUE_REG_13__4_ <= n3289;
    P2_INSTQUEUE_REG_13__3_ <= n3294;
    P2_INSTQUEUE_REG_13__2_ <= n3299;
    P2_INSTQUEUE_REG_13__1_ <= n3304;
    P2_INSTQUEUE_REG_13__0_ <= n3309;
    P2_INSTQUEUE_REG_12__7_ <= n3314;
    P2_INSTQUEUE_REG_12__6_ <= n3319;
    P2_INSTQUEUE_REG_12__5_ <= n3324;
    P2_INSTQUEUE_REG_12__4_ <= n3329;
    P2_INSTQUEUE_REG_12__3_ <= n3334;
    P2_INSTQUEUE_REG_12__2_ <= n3339;
    P2_INSTQUEUE_REG_12__1_ <= n3344;
    P2_INSTQUEUE_REG_12__0_ <= n3349;
    P2_INSTQUEUE_REG_11__7_ <= n3354;
    P2_INSTQUEUE_REG_11__6_ <= n3359;
    P2_INSTQUEUE_REG_11__5_ <= n3364;
    P2_INSTQUEUE_REG_11__4_ <= n3369;
    P2_INSTQUEUE_REG_11__3_ <= n3374;
    P2_INSTQUEUE_REG_11__2_ <= n3379;
    P2_INSTQUEUE_REG_11__1_ <= n3384;
    P2_INSTQUEUE_REG_11__0_ <= n3389;
    P2_INSTQUEUE_REG_10__7_ <= n3394;
    P2_INSTQUEUE_REG_10__6_ <= n3399;
    P2_INSTQUEUE_REG_10__5_ <= n3404;
    P2_INSTQUEUE_REG_10__4_ <= n3409;
    P2_INSTQUEUE_REG_10__3_ <= n3414;
    P2_INSTQUEUE_REG_10__2_ <= n3419;
    P2_INSTQUEUE_REG_10__1_ <= n3424;
    P2_INSTQUEUE_REG_10__0_ <= n3429;
    P2_INSTQUEUE_REG_9__7_ <= n3434;
    P2_INSTQUEUE_REG_9__6_ <= n3439;
    P2_INSTQUEUE_REG_9__5_ <= n3444;
    P2_INSTQUEUE_REG_9__4_ <= n3449;
    P2_INSTQUEUE_REG_9__3_ <= n3454;
    P2_INSTQUEUE_REG_9__2_ <= n3459;
    P2_INSTQUEUE_REG_9__1_ <= n3464;
    P2_INSTQUEUE_REG_9__0_ <= n3469;
    P2_INSTQUEUE_REG_8__7_ <= n3474;
    P2_INSTQUEUE_REG_8__6_ <= n3479;
    P2_INSTQUEUE_REG_8__5_ <= n3484;
    P2_INSTQUEUE_REG_8__4_ <= n3489;
    P2_INSTQUEUE_REG_8__3_ <= n3494;
    P2_INSTQUEUE_REG_8__2_ <= n3499;
    P2_INSTQUEUE_REG_8__1_ <= n3504;
    P2_INSTQUEUE_REG_8__0_ <= n3509;
    P2_INSTQUEUE_REG_7__7_ <= n3514;
    P2_INSTQUEUE_REG_7__6_ <= n3519;
    P2_INSTQUEUE_REG_7__5_ <= n3524;
    P2_INSTQUEUE_REG_7__4_ <= n3529;
    P2_INSTQUEUE_REG_7__3_ <= n3534;
    P2_INSTQUEUE_REG_7__2_ <= n3539;
    P2_INSTQUEUE_REG_7__1_ <= n3544;
    P2_INSTQUEUE_REG_7__0_ <= n3549;
    P2_INSTQUEUE_REG_6__7_ <= n3554;
    P2_INSTQUEUE_REG_6__6_ <= n3559;
    P2_INSTQUEUE_REG_6__5_ <= n3564;
    P2_INSTQUEUE_REG_6__4_ <= n3569;
    P2_INSTQUEUE_REG_6__3_ <= n3574;
    P2_INSTQUEUE_REG_6__2_ <= n3579;
    P2_INSTQUEUE_REG_6__1_ <= n3584;
    P2_INSTQUEUE_REG_6__0_ <= n3589;
    P2_INSTQUEUE_REG_5__7_ <= n3594;
    P2_INSTQUEUE_REG_5__6_ <= n3599;
    P2_INSTQUEUE_REG_5__5_ <= n3604;
    P2_INSTQUEUE_REG_5__4_ <= n3609;
    P2_INSTQUEUE_REG_5__3_ <= n3614;
    P2_INSTQUEUE_REG_5__2_ <= n3619;
    P2_INSTQUEUE_REG_5__1_ <= n3624;
    P2_INSTQUEUE_REG_5__0_ <= n3629;
    P2_INSTQUEUE_REG_4__7_ <= n3634;
    P2_INSTQUEUE_REG_4__6_ <= n3639;
    P2_INSTQUEUE_REG_4__5_ <= n3644;
    P2_INSTQUEUE_REG_4__4_ <= n3649;
    P2_INSTQUEUE_REG_4__3_ <= n3654;
    P2_INSTQUEUE_REG_4__2_ <= n3659;
    P2_INSTQUEUE_REG_4__1_ <= n3664;
    P2_INSTQUEUE_REG_4__0_ <= n3669;
    P2_INSTQUEUE_REG_3__7_ <= n3674;
    P2_INSTQUEUE_REG_3__6_ <= n3679;
    P2_INSTQUEUE_REG_3__5_ <= n3684;
    P2_INSTQUEUE_REG_3__4_ <= n3689;
    P2_INSTQUEUE_REG_3__3_ <= n3694;
    P2_INSTQUEUE_REG_3__2_ <= n3699;
    P2_INSTQUEUE_REG_3__1_ <= n3704;
    P2_INSTQUEUE_REG_3__0_ <= n3709;
    P2_INSTQUEUE_REG_2__7_ <= n3714;
    P2_INSTQUEUE_REG_2__6_ <= n3719;
    P2_INSTQUEUE_REG_2__5_ <= n3724;
    P2_INSTQUEUE_REG_2__4_ <= n3729;
    P2_INSTQUEUE_REG_2__3_ <= n3734;
    P2_INSTQUEUE_REG_2__2_ <= n3739;
    P2_INSTQUEUE_REG_2__1_ <= n3744;
    P2_INSTQUEUE_REG_2__0_ <= n3749;
    P2_INSTQUEUE_REG_1__7_ <= n3754;
    P2_INSTQUEUE_REG_1__6_ <= n3759;
    P2_INSTQUEUE_REG_1__5_ <= n3764;
    P2_INSTQUEUE_REG_1__4_ <= n3769;
    P2_INSTQUEUE_REG_1__3_ <= n3774;
    P2_INSTQUEUE_REG_1__2_ <= n3779;
    P2_INSTQUEUE_REG_1__1_ <= n3784;
    P2_INSTQUEUE_REG_1__0_ <= n3789;
    P2_INSTQUEUE_REG_0__7_ <= n3794;
    P2_INSTQUEUE_REG_0__6_ <= n3799;
    P2_INSTQUEUE_REG_0__5_ <= n3804;
    P2_INSTQUEUE_REG_0__4_ <= n3809;
    P2_INSTQUEUE_REG_0__3_ <= n3814;
    P2_INSTQUEUE_REG_0__2_ <= n3819;
    P2_INSTQUEUE_REG_0__1_ <= n3824;
    P2_INSTQUEUE_REG_0__0_ <= n3829;
    P2_INSTQUEUERD_ADDR_REG_4_ <= n3834;
    P2_INSTQUEUERD_ADDR_REG_3_ <= n3839;
    P2_INSTQUEUERD_ADDR_REG_2_ <= n3844;
    P2_INSTQUEUERD_ADDR_REG_1_ <= n3849;
    P2_INSTQUEUERD_ADDR_REG_0_ <= n3854;
    P2_INSTQUEUEWR_ADDR_REG_4_ <= n3859;
    P2_INSTQUEUEWR_ADDR_REG_3_ <= n3864;
    P2_INSTQUEUEWR_ADDR_REG_2_ <= n3869;
    P2_INSTQUEUEWR_ADDR_REG_1_ <= n3874;
    P2_INSTQUEUEWR_ADDR_REG_0_ <= n3879;
    P2_INSTADDRPOINTER_REG_0_ <= n3884;
    P2_INSTADDRPOINTER_REG_1_ <= n3889;
    P2_INSTADDRPOINTER_REG_2_ <= n3894;
    P2_INSTADDRPOINTER_REG_3_ <= n3899;
    P2_INSTADDRPOINTER_REG_4_ <= n3904;
    P2_INSTADDRPOINTER_REG_5_ <= n3909;
    P2_INSTADDRPOINTER_REG_6_ <= n3914;
    P2_INSTADDRPOINTER_REG_7_ <= n3919;
    P2_INSTADDRPOINTER_REG_8_ <= n3924;
    P2_INSTADDRPOINTER_REG_9_ <= n3929;
    P2_INSTADDRPOINTER_REG_10_ <= n3934;
    P2_INSTADDRPOINTER_REG_11_ <= n3939;
    P2_INSTADDRPOINTER_REG_12_ <= n3944;
    P2_INSTADDRPOINTER_REG_13_ <= n3949;
    P2_INSTADDRPOINTER_REG_14_ <= n3954;
    P2_INSTADDRPOINTER_REG_15_ <= n3959;
    P2_INSTADDRPOINTER_REG_16_ <= n3964;
    P2_INSTADDRPOINTER_REG_17_ <= n3969;
    P2_INSTADDRPOINTER_REG_18_ <= n3974;
    P2_INSTADDRPOINTER_REG_19_ <= n3979;
    P2_INSTADDRPOINTER_REG_20_ <= n3984;
    P2_INSTADDRPOINTER_REG_21_ <= n3989;
    P2_INSTADDRPOINTER_REG_22_ <= n3994;
    P2_INSTADDRPOINTER_REG_23_ <= n3999;
    P2_INSTADDRPOINTER_REG_24_ <= n4004;
    P2_INSTADDRPOINTER_REG_25_ <= n4009;
    P2_INSTADDRPOINTER_REG_26_ <= n4014;
    P2_INSTADDRPOINTER_REG_27_ <= n4019;
    P2_INSTADDRPOINTER_REG_28_ <= n4024;
    P2_INSTADDRPOINTER_REG_29_ <= n4029;
    P2_INSTADDRPOINTER_REG_30_ <= n4034;
    P2_INSTADDRPOINTER_REG_31_ <= n4039;
    P2_PHYADDRPOINTER_REG_0_ <= n4044;
    P2_PHYADDRPOINTER_REG_1_ <= n4049;
    P2_PHYADDRPOINTER_REG_2_ <= n4054;
    P2_PHYADDRPOINTER_REG_3_ <= n4059;
    P2_PHYADDRPOINTER_REG_4_ <= n4064;
    P2_PHYADDRPOINTER_REG_5_ <= n4069;
    P2_PHYADDRPOINTER_REG_6_ <= n4074;
    P2_PHYADDRPOINTER_REG_7_ <= n4079;
    P2_PHYADDRPOINTER_REG_8_ <= n4084;
    P2_PHYADDRPOINTER_REG_9_ <= n4089;
    P2_PHYADDRPOINTER_REG_10_ <= n4094;
    P2_PHYADDRPOINTER_REG_11_ <= n4099;
    P2_PHYADDRPOINTER_REG_12_ <= n4104;
    P2_PHYADDRPOINTER_REG_13_ <= n4109;
    P2_PHYADDRPOINTER_REG_14_ <= n4114;
    P2_PHYADDRPOINTER_REG_15_ <= n4119;
    P2_PHYADDRPOINTER_REG_16_ <= n4124;
    P2_PHYADDRPOINTER_REG_17_ <= n4129;
    P2_PHYADDRPOINTER_REG_18_ <= n4134;
    P2_PHYADDRPOINTER_REG_19_ <= n4139;
    P2_PHYADDRPOINTER_REG_20_ <= n4144;
    P2_PHYADDRPOINTER_REG_21_ <= n4149;
    P2_PHYADDRPOINTER_REG_22_ <= n4154;
    P2_PHYADDRPOINTER_REG_23_ <= n4159;
    P2_PHYADDRPOINTER_REG_24_ <= n4164;
    P2_PHYADDRPOINTER_REG_25_ <= n4169;
    P2_PHYADDRPOINTER_REG_26_ <= n4174;
    P2_PHYADDRPOINTER_REG_27_ <= n4179;
    P2_PHYADDRPOINTER_REG_28_ <= n4184;
    P2_PHYADDRPOINTER_REG_29_ <= n4189;
    P2_PHYADDRPOINTER_REG_30_ <= n4194;
    P2_PHYADDRPOINTER_REG_31_ <= n4199;
    P2_LWORD_REG_15_ <= n4204;
    P2_LWORD_REG_14_ <= n4209;
    P2_LWORD_REG_13_ <= n4214;
    P2_LWORD_REG_12_ <= n4219;
    P2_LWORD_REG_11_ <= n4224;
    P2_LWORD_REG_10_ <= n4229;
    P2_LWORD_REG_9_ <= n4234;
    P2_LWORD_REG_8_ <= n4239;
    P2_LWORD_REG_7_ <= n4244;
    P2_LWORD_REG_6_ <= n4249;
    P2_LWORD_REG_5_ <= n4254;
    P2_LWORD_REG_4_ <= n4259;
    P2_LWORD_REG_3_ <= n4264;
    P2_LWORD_REG_2_ <= n4269;
    P2_LWORD_REG_1_ <= n4274;
    P2_LWORD_REG_0_ <= n4279;
    P2_UWORD_REG_14_ <= n4284;
    P2_UWORD_REG_13_ <= n4289;
    P2_UWORD_REG_12_ <= n4294;
    P2_UWORD_REG_11_ <= n4299;
    P2_UWORD_REG_10_ <= n4304;
    P2_UWORD_REG_9_ <= n4309;
    P2_UWORD_REG_8_ <= n4314;
    P2_UWORD_REG_7_ <= n4319;
    P2_UWORD_REG_6_ <= n4324;
    P2_UWORD_REG_5_ <= n4329;
    P2_UWORD_REG_4_ <= n4334;
    P2_UWORD_REG_3_ <= n4339;
    P2_UWORD_REG_2_ <= n4344;
    P2_UWORD_REG_1_ <= n4349;
    P2_UWORD_REG_0_ <= n4354;
    P2_DATAO_REG_0_ <= n4359;
    P2_DATAO_REG_1_ <= n4364;
    P2_DATAO_REG_2_ <= n4369;
    P2_DATAO_REG_3_ <= n4374;
    P2_DATAO_REG_4_ <= n4379;
    P2_DATAO_REG_5_ <= n4384;
    P2_DATAO_REG_6_ <= n4389;
    P2_DATAO_REG_7_ <= n4394;
    P2_DATAO_REG_8_ <= n4399;
    P2_DATAO_REG_9_ <= n4404;
    P2_DATAO_REG_10_ <= n4409;
    P2_DATAO_REG_11_ <= n4414;
    P2_DATAO_REG_12_ <= n4419;
    P2_DATAO_REG_13_ <= n4424;
    P2_DATAO_REG_14_ <= n4429;
    P2_DATAO_REG_15_ <= n4434;
    P2_DATAO_REG_16_ <= n4439;
    P2_DATAO_REG_17_ <= n4444;
    P2_DATAO_REG_18_ <= n4449;
    P2_DATAO_REG_19_ <= n4454;
    P2_DATAO_REG_20_ <= n4459;
    P2_DATAO_REG_21_ <= n4464;
    P2_DATAO_REG_22_ <= n4469;
    P2_DATAO_REG_23_ <= n4474;
    P2_DATAO_REG_24_ <= n4479;
    P2_DATAO_REG_25_ <= n4484;
    P2_DATAO_REG_26_ <= n4489;
    P2_DATAO_REG_27_ <= n4494;
    P2_DATAO_REG_28_ <= n4499;
    P2_DATAO_REG_29_ <= n4504;
    P2_DATAO_REG_30_ <= n4509;
    P2_DATAO_REG_31_ <= n4514;
    P2_EAX_REG_0_ <= n4519;
    P2_EAX_REG_1_ <= n4524;
    P2_EAX_REG_2_ <= n4529;
    P2_EAX_REG_3_ <= n4534;
    P2_EAX_REG_4_ <= n4539;
    P2_EAX_REG_5_ <= n4544;
    P2_EAX_REG_6_ <= n4549;
    P2_EAX_REG_7_ <= n4554;
    P2_EAX_REG_8_ <= n4559;
    P2_EAX_REG_9_ <= n4564;
    P2_EAX_REG_10_ <= n4569;
    P2_EAX_REG_11_ <= n4574;
    P2_EAX_REG_12_ <= n4579;
    P2_EAX_REG_13_ <= n4584;
    P2_EAX_REG_14_ <= n4589;
    P2_EAX_REG_15_ <= n4594;
    P2_EAX_REG_16_ <= n4599;
    P2_EAX_REG_17_ <= n4604;
    P2_EAX_REG_18_ <= n4609;
    P2_EAX_REG_19_ <= n4614;
    P2_EAX_REG_20_ <= n4619;
    P2_EAX_REG_21_ <= n4624;
    P2_EAX_REG_22_ <= n4629;
    P2_EAX_REG_23_ <= n4634;
    P2_EAX_REG_24_ <= n4639;
    P2_EAX_REG_25_ <= n4644;
    P2_EAX_REG_26_ <= n4649;
    P2_EAX_REG_27_ <= n4654;
    P2_EAX_REG_28_ <= n4659;
    P2_EAX_REG_29_ <= n4664;
    P2_EAX_REG_30_ <= n4669;
    P2_EAX_REG_31_ <= n4674;
    P2_EBX_REG_0_ <= n4679;
    P2_EBX_REG_1_ <= n4684;
    P2_EBX_REG_2_ <= n4689;
    P2_EBX_REG_3_ <= n4694;
    P2_EBX_REG_4_ <= n4699;
    P2_EBX_REG_5_ <= n4704;
    P2_EBX_REG_6_ <= n4709;
    P2_EBX_REG_7_ <= n4714;
    P2_EBX_REG_8_ <= n4719;
    P2_EBX_REG_9_ <= n4724;
    P2_EBX_REG_10_ <= n4729;
    P2_EBX_REG_11_ <= n4734;
    P2_EBX_REG_12_ <= n4739;
    P2_EBX_REG_13_ <= n4744;
    P2_EBX_REG_14_ <= n4749;
    P2_EBX_REG_15_ <= n4754;
    P2_EBX_REG_16_ <= n4759;
    P2_EBX_REG_17_ <= n4764;
    P2_EBX_REG_18_ <= n4769;
    P2_EBX_REG_19_ <= n4774;
    P2_EBX_REG_20_ <= n4779;
    P2_EBX_REG_21_ <= n4784;
    P2_EBX_REG_22_ <= n4789;
    P2_EBX_REG_23_ <= n4794;
    P2_EBX_REG_24_ <= n4799;
    P2_EBX_REG_25_ <= n4804;
    P2_EBX_REG_26_ <= n4809;
    P2_EBX_REG_27_ <= n4814;
    P2_EBX_REG_28_ <= n4819;
    P2_EBX_REG_29_ <= n4824;
    P2_EBX_REG_30_ <= n4829;
    P2_EBX_REG_31_ <= n4834;
    P2_REIP_REG_0_ <= n4839;
    P2_REIP_REG_1_ <= n4844;
    P2_REIP_REG_2_ <= n4849;
    P2_REIP_REG_3_ <= n4854;
    P2_REIP_REG_4_ <= n4859;
    P2_REIP_REG_5_ <= n4864;
    P2_REIP_REG_6_ <= n4869;
    P2_REIP_REG_7_ <= n4874;
    P2_REIP_REG_8_ <= n4879;
    P2_REIP_REG_9_ <= n4884;
    P2_REIP_REG_10_ <= n4889;
    P2_REIP_REG_11_ <= n4894;
    P2_REIP_REG_12_ <= n4899;
    P2_REIP_REG_13_ <= n4904;
    P2_REIP_REG_14_ <= n4909;
    P2_REIP_REG_15_ <= n4914;
    P2_REIP_REG_16_ <= n4919;
    P2_REIP_REG_17_ <= n4924;
    P2_REIP_REG_18_ <= n4929;
    P2_REIP_REG_19_ <= n4934;
    P2_REIP_REG_20_ <= n4939;
    P2_REIP_REG_21_ <= n4944;
    P2_REIP_REG_22_ <= n4949;
    P2_REIP_REG_23_ <= n4954;
    P2_REIP_REG_24_ <= n4959;
    P2_REIP_REG_25_ <= n4964;
    P2_REIP_REG_26_ <= n4969;
    P2_REIP_REG_27_ <= n4974;
    P2_REIP_REG_28_ <= n4979;
    P2_REIP_REG_29_ <= n4984;
    P2_REIP_REG_30_ <= n4989;
    P2_REIP_REG_31_ <= n4994;
    P2_BYTEENABLE_REG_3_ <= n4999;
    P2_BYTEENABLE_REG_2_ <= n5004;
    P2_BYTEENABLE_REG_1_ <= n5009;
    P2_BYTEENABLE_REG_0_ <= n5014;
    P2_W_R_N_REG <= n5019;
    P2_FLUSH_REG <= n5024;
    P2_MORE_REG <= n5029;
    P2_STATEBS16_REG <= n5034;
    P2_REQUESTPENDING_REG <= n5039;
    P2_D_C_N_REG <= n5044;
    P2_M_IO_N_REG <= n5049;
    P2_CODEFETCH_REG <= n5054;
    P2_ADS_N_REG <= n5059;
    P2_READREQUEST_REG <= n5064;
    P2_MEMORYFETCH_REG <= n5069;
    P1_BE_N_REG_3_ <= n5074;
    P1_BE_N_REG_2_ <= n5079;
    P1_BE_N_REG_1_ <= n5084;
    P1_BE_N_REG_0_ <= n5089;
    P1_ADDRESS_REG_29_ <= n5094;
    P1_ADDRESS_REG_28_ <= n5098;
    P1_ADDRESS_REG_27_ <= n5102;
    P1_ADDRESS_REG_26_ <= n5106;
    P1_ADDRESS_REG_25_ <= n5110;
    P1_ADDRESS_REG_24_ <= n5114;
    P1_ADDRESS_REG_23_ <= n5118;
    P1_ADDRESS_REG_22_ <= n5122;
    P1_ADDRESS_REG_21_ <= n5126;
    P1_ADDRESS_REG_20_ <= n5130;
    P1_ADDRESS_REG_19_ <= n5134;
    P1_ADDRESS_REG_18_ <= n5138;
    P1_ADDRESS_REG_17_ <= n5142;
    P1_ADDRESS_REG_16_ <= n5146;
    P1_ADDRESS_REG_15_ <= n5150;
    P1_ADDRESS_REG_14_ <= n5154;
    P1_ADDRESS_REG_13_ <= n5158;
    P1_ADDRESS_REG_12_ <= n5162;
    P1_ADDRESS_REG_11_ <= n5166;
    P1_ADDRESS_REG_10_ <= n5170;
    P1_ADDRESS_REG_9_ <= n5174;
    P1_ADDRESS_REG_8_ <= n5178;
    P1_ADDRESS_REG_7_ <= n5182;
    P1_ADDRESS_REG_6_ <= n5186;
    P1_ADDRESS_REG_5_ <= n5190;
    P1_ADDRESS_REG_4_ <= n5194;
    P1_ADDRESS_REG_3_ <= n5198;
    P1_ADDRESS_REG_2_ <= n5202;
    P1_ADDRESS_REG_1_ <= n5206;
    P1_ADDRESS_REG_0_ <= n5210;
    P1_STATE_REG_2_ <= n5214;
    P1_STATE_REG_1_ <= n5219;
    P1_STATE_REG_0_ <= n5224;
    P1_DATAWIDTH_REG_0_ <= n5229;
    P1_DATAWIDTH_REG_1_ <= n5234;
    P1_DATAWIDTH_REG_2_ <= n5239;
    P1_DATAWIDTH_REG_3_ <= n5244;
    P1_DATAWIDTH_REG_4_ <= n5249;
    P1_DATAWIDTH_REG_5_ <= n5254;
    P1_DATAWIDTH_REG_6_ <= n5259;
    P1_DATAWIDTH_REG_7_ <= n5264;
    P1_DATAWIDTH_REG_8_ <= n5269;
    P1_DATAWIDTH_REG_9_ <= n5274;
    P1_DATAWIDTH_REG_10_ <= n5279;
    P1_DATAWIDTH_REG_11_ <= n5284;
    P1_DATAWIDTH_REG_12_ <= n5289;
    P1_DATAWIDTH_REG_13_ <= n5294;
    P1_DATAWIDTH_REG_14_ <= n5299;
    P1_DATAWIDTH_REG_15_ <= n5304;
    P1_DATAWIDTH_REG_16_ <= n5309;
    P1_DATAWIDTH_REG_17_ <= n5314;
    P1_DATAWIDTH_REG_18_ <= n5319;
    P1_DATAWIDTH_REG_19_ <= n5324;
    P1_DATAWIDTH_REG_20_ <= n5329;
    P1_DATAWIDTH_REG_21_ <= n5334;
    P1_DATAWIDTH_REG_22_ <= n5339;
    P1_DATAWIDTH_REG_23_ <= n5344;
    P1_DATAWIDTH_REG_24_ <= n5349;
    P1_DATAWIDTH_REG_25_ <= n5354;
    P1_DATAWIDTH_REG_26_ <= n5359;
    P1_DATAWIDTH_REG_27_ <= n5364;
    P1_DATAWIDTH_REG_28_ <= n5369;
    P1_DATAWIDTH_REG_29_ <= n5374;
    P1_DATAWIDTH_REG_30_ <= n5379;
    P1_DATAWIDTH_REG_31_ <= n5384;
    P1_STATE2_REG_3_ <= n5389;
    P1_STATE2_REG_2_ <= n5394;
    P1_STATE2_REG_1_ <= n5399;
    P1_STATE2_REG_0_ <= n5404;
    P1_INSTQUEUE_REG_15__7_ <= n5409;
    P1_INSTQUEUE_REG_15__6_ <= n5414;
    P1_INSTQUEUE_REG_15__5_ <= n5419;
    P1_INSTQUEUE_REG_15__4_ <= n5424;
    P1_INSTQUEUE_REG_15__3_ <= n5429;
    P1_INSTQUEUE_REG_15__2_ <= n5434;
    P1_INSTQUEUE_REG_15__1_ <= n5439;
    P1_INSTQUEUE_REG_15__0_ <= n5444;
    P1_INSTQUEUE_REG_14__7_ <= n5449;
    P1_INSTQUEUE_REG_14__6_ <= n5454;
    P1_INSTQUEUE_REG_14__5_ <= n5459;
    P1_INSTQUEUE_REG_14__4_ <= n5464;
    P1_INSTQUEUE_REG_14__3_ <= n5469;
    P1_INSTQUEUE_REG_14__2_ <= n5474;
    P1_INSTQUEUE_REG_14__1_ <= n5479;
    P1_INSTQUEUE_REG_14__0_ <= n5484;
    P1_INSTQUEUE_REG_13__7_ <= n5489;
    P1_INSTQUEUE_REG_13__6_ <= n5494;
    P1_INSTQUEUE_REG_13__5_ <= n5499;
    P1_INSTQUEUE_REG_13__4_ <= n5504;
    P1_INSTQUEUE_REG_13__3_ <= n5509;
    P1_INSTQUEUE_REG_13__2_ <= n5514;
    P1_INSTQUEUE_REG_13__1_ <= n5519;
    P1_INSTQUEUE_REG_13__0_ <= n5524;
    P1_INSTQUEUE_REG_12__7_ <= n5529;
    P1_INSTQUEUE_REG_12__6_ <= n5534;
    P1_INSTQUEUE_REG_12__5_ <= n5539;
    P1_INSTQUEUE_REG_12__4_ <= n5544;
    P1_INSTQUEUE_REG_12__3_ <= n5549;
    P1_INSTQUEUE_REG_12__2_ <= n5554;
    P1_INSTQUEUE_REG_12__1_ <= n5559;
    P1_INSTQUEUE_REG_12__0_ <= n5564;
    P1_INSTQUEUE_REG_11__7_ <= n5569;
    P1_INSTQUEUE_REG_11__6_ <= n5574;
    P1_INSTQUEUE_REG_11__5_ <= n5579;
    P1_INSTQUEUE_REG_11__4_ <= n5584;
    P1_INSTQUEUE_REG_11__3_ <= n5589;
    P1_INSTQUEUE_REG_11__2_ <= n5594;
    P1_INSTQUEUE_REG_11__1_ <= n5599;
    P1_INSTQUEUE_REG_11__0_ <= n5604;
    P1_INSTQUEUE_REG_10__7_ <= n5609;
    P1_INSTQUEUE_REG_10__6_ <= n5614;
    P1_INSTQUEUE_REG_10__5_ <= n5619;
    P1_INSTQUEUE_REG_10__4_ <= n5624;
    P1_INSTQUEUE_REG_10__3_ <= n5629;
    P1_INSTQUEUE_REG_10__2_ <= n5634;
    P1_INSTQUEUE_REG_10__1_ <= n5639;
    P1_INSTQUEUE_REG_10__0_ <= n5644;
    P1_INSTQUEUE_REG_9__7_ <= n5649;
    P1_INSTQUEUE_REG_9__6_ <= n5654;
    P1_INSTQUEUE_REG_9__5_ <= n5659;
    P1_INSTQUEUE_REG_9__4_ <= n5664;
    P1_INSTQUEUE_REG_9__3_ <= n5669;
    P1_INSTQUEUE_REG_9__2_ <= n5674;
    P1_INSTQUEUE_REG_9__1_ <= n5679;
    P1_INSTQUEUE_REG_9__0_ <= n5684;
    P1_INSTQUEUE_REG_8__7_ <= n5689;
    P1_INSTQUEUE_REG_8__6_ <= n5694;
    P1_INSTQUEUE_REG_8__5_ <= n5699;
    P1_INSTQUEUE_REG_8__4_ <= n5704;
    P1_INSTQUEUE_REG_8__3_ <= n5709;
    P1_INSTQUEUE_REG_8__2_ <= n5714;
    P1_INSTQUEUE_REG_8__1_ <= n5719;
    P1_INSTQUEUE_REG_8__0_ <= n5724;
    P1_INSTQUEUE_REG_7__7_ <= n5729;
    P1_INSTQUEUE_REG_7__6_ <= n5734;
    P1_INSTQUEUE_REG_7__5_ <= n5739;
    P1_INSTQUEUE_REG_7__4_ <= n5744;
    P1_INSTQUEUE_REG_7__3_ <= n5749;
    P1_INSTQUEUE_REG_7__2_ <= n5754;
    P1_INSTQUEUE_REG_7__1_ <= n5759;
    P1_INSTQUEUE_REG_7__0_ <= n5764;
    P1_INSTQUEUE_REG_6__7_ <= n5769;
    P1_INSTQUEUE_REG_6__6_ <= n5774;
    P1_INSTQUEUE_REG_6__5_ <= n5779;
    P1_INSTQUEUE_REG_6__4_ <= n5784;
    P1_INSTQUEUE_REG_6__3_ <= n5789;
    P1_INSTQUEUE_REG_6__2_ <= n5794;
    P1_INSTQUEUE_REG_6__1_ <= n5799;
    P1_INSTQUEUE_REG_6__0_ <= n5804;
    P1_INSTQUEUE_REG_5__7_ <= n5809;
    P1_INSTQUEUE_REG_5__6_ <= n5814;
    P1_INSTQUEUE_REG_5__5_ <= n5819;
    P1_INSTQUEUE_REG_5__4_ <= n5824;
    P1_INSTQUEUE_REG_5__3_ <= n5829;
    P1_INSTQUEUE_REG_5__2_ <= n5834;
    P1_INSTQUEUE_REG_5__1_ <= n5839;
    P1_INSTQUEUE_REG_5__0_ <= n5844;
    P1_INSTQUEUE_REG_4__7_ <= n5849;
    P1_INSTQUEUE_REG_4__6_ <= n5854;
    P1_INSTQUEUE_REG_4__5_ <= n5859;
    P1_INSTQUEUE_REG_4__4_ <= n5864;
    P1_INSTQUEUE_REG_4__3_ <= n5869;
    P1_INSTQUEUE_REG_4__2_ <= n5874;
    P1_INSTQUEUE_REG_4__1_ <= n5879;
    P1_INSTQUEUE_REG_4__0_ <= n5884;
    P1_INSTQUEUE_REG_3__7_ <= n5889;
    P1_INSTQUEUE_REG_3__6_ <= n5894;
    P1_INSTQUEUE_REG_3__5_ <= n5899;
    P1_INSTQUEUE_REG_3__4_ <= n5904;
    P1_INSTQUEUE_REG_3__3_ <= n5909;
    P1_INSTQUEUE_REG_3__2_ <= n5914;
    P1_INSTQUEUE_REG_3__1_ <= n5919;
    P1_INSTQUEUE_REG_3__0_ <= n5924;
    P1_INSTQUEUE_REG_2__7_ <= n5929;
    P1_INSTQUEUE_REG_2__6_ <= n5934;
    P1_INSTQUEUE_REG_2__5_ <= n5939;
    P1_INSTQUEUE_REG_2__4_ <= n5944;
    P1_INSTQUEUE_REG_2__3_ <= n5949;
    P1_INSTQUEUE_REG_2__2_ <= n5954;
    P1_INSTQUEUE_REG_2__1_ <= n5959;
    P1_INSTQUEUE_REG_2__0_ <= n5964;
    P1_INSTQUEUE_REG_1__7_ <= n5969;
    P1_INSTQUEUE_REG_1__6_ <= n5974;
    P1_INSTQUEUE_REG_1__5_ <= n5979;
    P1_INSTQUEUE_REG_1__4_ <= n5984;
    P1_INSTQUEUE_REG_1__3_ <= n5989;
    P1_INSTQUEUE_REG_1__2_ <= n5994;
    P1_INSTQUEUE_REG_1__1_ <= n5999;
    P1_INSTQUEUE_REG_1__0_ <= n6004;
    P1_INSTQUEUE_REG_0__7_ <= n6009;
    P1_INSTQUEUE_REG_0__6_ <= n6014;
    P1_INSTQUEUE_REG_0__5_ <= n6019;
    P1_INSTQUEUE_REG_0__4_ <= n6024;
    P1_INSTQUEUE_REG_0__3_ <= n6029;
    P1_INSTQUEUE_REG_0__2_ <= n6034;
    P1_INSTQUEUE_REG_0__1_ <= n6039;
    P1_INSTQUEUE_REG_0__0_ <= n6044;
    P1_INSTQUEUERD_ADDR_REG_4_ <= n6049;
    P1_INSTQUEUERD_ADDR_REG_3_ <= n6054;
    P1_INSTQUEUERD_ADDR_REG_2_ <= n6059;
    P1_INSTQUEUERD_ADDR_REG_1_ <= n6064;
    P1_INSTQUEUERD_ADDR_REG_0_ <= n6069;
    P1_INSTQUEUEWR_ADDR_REG_4_ <= n6074;
    P1_INSTQUEUEWR_ADDR_REG_3_ <= n6079;
    P1_INSTQUEUEWR_ADDR_REG_2_ <= n6084;
    P1_INSTQUEUEWR_ADDR_REG_1_ <= n6089;
    P1_INSTQUEUEWR_ADDR_REG_0_ <= n6094;
    P1_INSTADDRPOINTER_REG_0_ <= n6099;
    P1_INSTADDRPOINTER_REG_1_ <= n6104;
    P1_INSTADDRPOINTER_REG_2_ <= n6109;
    P1_INSTADDRPOINTER_REG_3_ <= n6114;
    P1_INSTADDRPOINTER_REG_4_ <= n6119;
    P1_INSTADDRPOINTER_REG_5_ <= n6124;
    P1_INSTADDRPOINTER_REG_6_ <= n6129;
    P1_INSTADDRPOINTER_REG_7_ <= n6134;
    P1_INSTADDRPOINTER_REG_8_ <= n6139;
    P1_INSTADDRPOINTER_REG_9_ <= n6144;
    P1_INSTADDRPOINTER_REG_10_ <= n6149;
    P1_INSTADDRPOINTER_REG_11_ <= n6154;
    P1_INSTADDRPOINTER_REG_12_ <= n6159;
    P1_INSTADDRPOINTER_REG_13_ <= n6164;
    P1_INSTADDRPOINTER_REG_14_ <= n6169;
    P1_INSTADDRPOINTER_REG_15_ <= n6174;
    P1_INSTADDRPOINTER_REG_16_ <= n6179;
    P1_INSTADDRPOINTER_REG_17_ <= n6184;
    P1_INSTADDRPOINTER_REG_18_ <= n6189;
    P1_INSTADDRPOINTER_REG_19_ <= n6194;
    P1_INSTADDRPOINTER_REG_20_ <= n6199;
    P1_INSTADDRPOINTER_REG_21_ <= n6204;
    P1_INSTADDRPOINTER_REG_22_ <= n6209;
    P1_INSTADDRPOINTER_REG_23_ <= n6214;
    P1_INSTADDRPOINTER_REG_24_ <= n6219;
    P1_INSTADDRPOINTER_REG_25_ <= n6224;
    P1_INSTADDRPOINTER_REG_26_ <= n6229;
    P1_INSTADDRPOINTER_REG_27_ <= n6234;
    P1_INSTADDRPOINTER_REG_28_ <= n6239;
    P1_INSTADDRPOINTER_REG_29_ <= n6244;
    P1_INSTADDRPOINTER_REG_30_ <= n6249;
    P1_INSTADDRPOINTER_REG_31_ <= n6254;
    P1_PHYADDRPOINTER_REG_0_ <= n6259;
    P1_PHYADDRPOINTER_REG_1_ <= n6264;
    P1_PHYADDRPOINTER_REG_2_ <= n6269;
    P1_PHYADDRPOINTER_REG_3_ <= n6274;
    P1_PHYADDRPOINTER_REG_4_ <= n6279;
    P1_PHYADDRPOINTER_REG_5_ <= n6284;
    P1_PHYADDRPOINTER_REG_6_ <= n6289;
    P1_PHYADDRPOINTER_REG_7_ <= n6294;
    P1_PHYADDRPOINTER_REG_8_ <= n6299;
    P1_PHYADDRPOINTER_REG_9_ <= n6304;
    P1_PHYADDRPOINTER_REG_10_ <= n6309;
    P1_PHYADDRPOINTER_REG_11_ <= n6314;
    P1_PHYADDRPOINTER_REG_12_ <= n6319;
    P1_PHYADDRPOINTER_REG_13_ <= n6324;
    P1_PHYADDRPOINTER_REG_14_ <= n6329;
    P1_PHYADDRPOINTER_REG_15_ <= n6334;
    P1_PHYADDRPOINTER_REG_16_ <= n6339;
    P1_PHYADDRPOINTER_REG_17_ <= n6344;
    P1_PHYADDRPOINTER_REG_18_ <= n6349;
    P1_PHYADDRPOINTER_REG_19_ <= n6354;
    P1_PHYADDRPOINTER_REG_20_ <= n6359;
    P1_PHYADDRPOINTER_REG_21_ <= n6364;
    P1_PHYADDRPOINTER_REG_22_ <= n6369;
    P1_PHYADDRPOINTER_REG_23_ <= n6374;
    P1_PHYADDRPOINTER_REG_24_ <= n6379;
    P1_PHYADDRPOINTER_REG_25_ <= n6384;
    P1_PHYADDRPOINTER_REG_26_ <= n6389;
    P1_PHYADDRPOINTER_REG_27_ <= n6394;
    P1_PHYADDRPOINTER_REG_28_ <= n6399;
    P1_PHYADDRPOINTER_REG_29_ <= n6404;
    P1_PHYADDRPOINTER_REG_30_ <= n6409;
    P1_PHYADDRPOINTER_REG_31_ <= n6414;
    P1_LWORD_REG_15_ <= n6419;
    P1_LWORD_REG_14_ <= n6424;
    P1_LWORD_REG_13_ <= n6429;
    P1_LWORD_REG_12_ <= n6434;
    P1_LWORD_REG_11_ <= n6439;
    P1_LWORD_REG_10_ <= n6444;
    P1_LWORD_REG_9_ <= n6449;
    P1_LWORD_REG_8_ <= n6454;
    P1_LWORD_REG_7_ <= n6459;
    P1_LWORD_REG_6_ <= n6464;
    P1_LWORD_REG_5_ <= n6469;
    P1_LWORD_REG_4_ <= n6474;
    P1_LWORD_REG_3_ <= n6479;
    P1_LWORD_REG_2_ <= n6484;
    P1_LWORD_REG_1_ <= n6489;
    P1_LWORD_REG_0_ <= n6494;
    P1_UWORD_REG_14_ <= n6499;
    P1_UWORD_REG_13_ <= n6504;
    P1_UWORD_REG_12_ <= n6509;
    P1_UWORD_REG_11_ <= n6514;
    P1_UWORD_REG_10_ <= n6519;
    P1_UWORD_REG_9_ <= n6524;
    P1_UWORD_REG_8_ <= n6529;
    P1_UWORD_REG_7_ <= n6534;
    P1_UWORD_REG_6_ <= n6539;
    P1_UWORD_REG_5_ <= n6544;
    P1_UWORD_REG_4_ <= n6549;
    P1_UWORD_REG_3_ <= n6554;
    P1_UWORD_REG_2_ <= n6559;
    P1_UWORD_REG_1_ <= n6564;
    P1_UWORD_REG_0_ <= n6569;
    P1_DATAO_REG_0_ <= n6574;
    P1_DATAO_REG_1_ <= n6579;
    P1_DATAO_REG_2_ <= n6584;
    P1_DATAO_REG_3_ <= n6589;
    P1_DATAO_REG_4_ <= n6594;
    P1_DATAO_REG_5_ <= n6599;
    P1_DATAO_REG_6_ <= n6604;
    P1_DATAO_REG_7_ <= n6609;
    P1_DATAO_REG_8_ <= n6614;
    P1_DATAO_REG_9_ <= n6619;
    P1_DATAO_REG_10_ <= n6624;
    P1_DATAO_REG_11_ <= n6629;
    P1_DATAO_REG_12_ <= n6634;
    P1_DATAO_REG_13_ <= n6639;
    P1_DATAO_REG_14_ <= n6644;
    P1_DATAO_REG_15_ <= n6649;
    P1_DATAO_REG_16_ <= n6654;
    P1_DATAO_REG_17_ <= n6659;
    P1_DATAO_REG_18_ <= n6664;
    P1_DATAO_REG_19_ <= n6669;
    P1_DATAO_REG_20_ <= n6674;
    P1_DATAO_REG_21_ <= n6679;
    P1_DATAO_REG_22_ <= n6684;
    P1_DATAO_REG_23_ <= n6689;
    P1_DATAO_REG_24_ <= n6694;
    P1_DATAO_REG_25_ <= n6699;
    P1_DATAO_REG_26_ <= n6704;
    P1_DATAO_REG_27_ <= n6709;
    P1_DATAO_REG_28_ <= n6714;
    P1_DATAO_REG_29_ <= n6719;
    P1_DATAO_REG_30_ <= n6724;
    P1_DATAO_REG_31_ <= n6729;
    P1_EAX_REG_0_ <= n6734;
    P1_EAX_REG_1_ <= n6739;
    P1_EAX_REG_2_ <= n6744;
    P1_EAX_REG_3_ <= n6749;
    P1_EAX_REG_4_ <= n6754;
    P1_EAX_REG_5_ <= n6759;
    P1_EAX_REG_6_ <= n6764;
    P1_EAX_REG_7_ <= n6769;
    P1_EAX_REG_8_ <= n6774;
    P1_EAX_REG_9_ <= n6779;
    P1_EAX_REG_10_ <= n6784;
    P1_EAX_REG_11_ <= n6789;
    P1_EAX_REG_12_ <= n6794;
    P1_EAX_REG_13_ <= n6799;
    P1_EAX_REG_14_ <= n6804;
    P1_EAX_REG_15_ <= n6809;
    P1_EAX_REG_16_ <= n6814;
    P1_EAX_REG_17_ <= n6819;
    P1_EAX_REG_18_ <= n6824;
    P1_EAX_REG_19_ <= n6829;
    P1_EAX_REG_20_ <= n6834;
    P1_EAX_REG_21_ <= n6839;
    P1_EAX_REG_22_ <= n6844;
    P1_EAX_REG_23_ <= n6849;
    P1_EAX_REG_24_ <= n6854;
    P1_EAX_REG_25_ <= n6859;
    P1_EAX_REG_26_ <= n6864;
    P1_EAX_REG_27_ <= n6869;
    P1_EAX_REG_28_ <= n6874;
    P1_EAX_REG_29_ <= n6879;
    P1_EAX_REG_30_ <= n6884;
    P1_EAX_REG_31_ <= n6889;
    P1_EBX_REG_0_ <= n6894;
    P1_EBX_REG_1_ <= n6899;
    P1_EBX_REG_2_ <= n6904;
    P1_EBX_REG_3_ <= n6909;
    P1_EBX_REG_4_ <= n6914;
    P1_EBX_REG_5_ <= n6919;
    P1_EBX_REG_6_ <= n6924;
    P1_EBX_REG_7_ <= n6929;
    P1_EBX_REG_8_ <= n6934;
    P1_EBX_REG_9_ <= n6939;
    P1_EBX_REG_10_ <= n6944;
    P1_EBX_REG_11_ <= n6949;
    P1_EBX_REG_12_ <= n6954;
    P1_EBX_REG_13_ <= n6959;
    P1_EBX_REG_14_ <= n6964;
    P1_EBX_REG_15_ <= n6969;
    P1_EBX_REG_16_ <= n6974;
    P1_EBX_REG_17_ <= n6979;
    P1_EBX_REG_18_ <= n6984;
    P1_EBX_REG_19_ <= n6989;
    P1_EBX_REG_20_ <= n6994;
    P1_EBX_REG_21_ <= n6999;
    P1_EBX_REG_22_ <= n7004;
    P1_EBX_REG_23_ <= n7009;
    P1_EBX_REG_24_ <= n7014;
    P1_EBX_REG_25_ <= n7019;
    P1_EBX_REG_26_ <= n7024;
    P1_EBX_REG_27_ <= n7029;
    P1_EBX_REG_28_ <= n7034;
    P1_EBX_REG_29_ <= n7039;
    P1_EBX_REG_30_ <= n7044;
    P1_EBX_REG_31_ <= n7049;
    P1_REIP_REG_0_ <= n7054;
    P1_REIP_REG_1_ <= n7059;
    P1_REIP_REG_2_ <= n7064;
    P1_REIP_REG_3_ <= n7069;
    P1_REIP_REG_4_ <= n7074;
    P1_REIP_REG_5_ <= n7079;
    P1_REIP_REG_6_ <= n7084;
    P1_REIP_REG_7_ <= n7089;
    P1_REIP_REG_8_ <= n7094;
    P1_REIP_REG_9_ <= n7099;
    P1_REIP_REG_10_ <= n7104;
    P1_REIP_REG_11_ <= n7109;
    P1_REIP_REG_12_ <= n7114;
    P1_REIP_REG_13_ <= n7119;
    P1_REIP_REG_14_ <= n7124;
    P1_REIP_REG_15_ <= n7129;
    P1_REIP_REG_16_ <= n7134;
    P1_REIP_REG_17_ <= n7139;
    P1_REIP_REG_18_ <= n7144;
    P1_REIP_REG_19_ <= n7149;
    P1_REIP_REG_20_ <= n7154;
    P1_REIP_REG_21_ <= n7159;
    P1_REIP_REG_22_ <= n7164;
    P1_REIP_REG_23_ <= n7169;
    P1_REIP_REG_24_ <= n7174;
    P1_REIP_REG_25_ <= n7179;
    P1_REIP_REG_26_ <= n7184;
    P1_REIP_REG_27_ <= n7189;
    P1_REIP_REG_28_ <= n7194;
    P1_REIP_REG_29_ <= n7199;
    P1_REIP_REG_30_ <= n7204;
    P1_REIP_REG_31_ <= n7209;
    P1_BYTEENABLE_REG_3_ <= n7214;
    P1_BYTEENABLE_REG_2_ <= n7219;
    P1_BYTEENABLE_REG_1_ <= n7224;
    P1_BYTEENABLE_REG_0_ <= n7229;
    P1_W_R_N_REG <= n7234;
    P1_FLUSH_REG <= n7239;
    P1_MORE_REG <= n7244;
    P1_STATEBS16_REG <= n7249;
    P1_REQUESTPENDING_REG <= n7254;
    P1_D_C_N_REG <= n7259;
    P1_M_IO_N_REG <= n7264;
    P1_CODEFETCH_REG <= n7269;
    P1_ADS_N_REG <= n7274;
    P1_READREQUEST_REG <= n7278;
    P1_MEMORYFETCH_REG <= n7283;
    Q_0 <= n67455;
    Q_1 <= n67458;
    Q_2 <= n67461;
    Q_3 <= n67464;
  end
endmodule
