library ieee;
use ieee.std_logic_1164.all;

entity sara is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y39,y40,y41,y42,y43,y44 : out std_logic );
end sara;

architecture ARC of sara is

   type states_sara is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
	s31,s32,s33,s34,s35,s36 );
   signal current_sara : states_sara;

begin
   process (clk , rst)
   procedure proc_sara is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;


   case current_sara is
   when s1 =>
      if ( x1 and x2 ) = '1' then
         y1 <= '1' ;
         current_sara <= s2;

      elsif ( x1 and not x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_sara <= s3;

      else
         current_sara <= s1;

      end if;

   when s2 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_sara <= s4;

   when s3 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y15 <= '1' ;
         y21 <= '1' ;
         current_sara <= s5;

   when s4 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_sara <= s6;

   when s5 =>
         y3 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_sara <= s7;

   when s6 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_sara <= s8;

   when s7 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y19 <= '1' ;
         current_sara <= s9;

   when s8 =>
      if ( x18 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_sara <= s10;

      else
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_sara <= s8;

      end if;

   when s9 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         y20 <= '1' ;
         current_sara <= s11;

   when s10 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_sara <= s12;

   when s11 =>
         y9 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_sara <= s1;

   when s12 =>
      if ( x17 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( x17 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( x17 and x16 and not x12 and not x13 ) = '1' then
         current_sara <= s1;

      elsif ( x17 and not x16 ) = '1' then
         current_sara <= s1;

      else
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y14 <= '1' ;
         current_sara <= s13;

      end if;

   when s13 =>
      if ( x15 ) = '1' then
         y1 <= '1' ;
         current_sara <= s2;

      elsif ( not x15 and x3 and x6 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and x3 and x6 and not x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_sara <= s15;

      elsif ( not x15 and x3 and not x6 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_sara <= s15;

      elsif ( not x15 and x3 and not x6 and not x5 and x10 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y32 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and x3 and not x6 and not x5 and not x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_sara <= s15;

      elsif ( not x15 and not x3 and x4 and x1 and x6 and x7 ) = '1' then
         y28 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and x1 and x6 and not x7 ) = '1' then
         y44 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and x8 and x13 ) = '1' then
         y9 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and x8 and not x13 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and x8 and not x13 and x16 and not x12 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and x8 and not x13 and not x16 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and not x8 and x12 and x13 ) = '1' then
         y9 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and not x8 and x12 and not x13 and x16 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and not x8 and x12 and not x13 and not x16 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and not x8 and not x12 and x16 and x13 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and not x8 and not x12 and x16 and not x13 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and x7 and not x8 and not x12 and not x16 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and not x7 and x8 ) = '1' then
         y23 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and x1 and not x6 and not x7 and not x8 ) = '1' then
         y11 <= '1' ;
         y15 <= '1' ;
         y41 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and not x1 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_sara <= s16;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and x7 and x8 ) = '1' then
         y41 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and x7 and not x8 ) = '1' then
         y40 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and not x7 and x8 ) = '1' then
         y39 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and x6 and not x7 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and x4 and not x1 and not x9 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_sara <= s17;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and not x7 and x8 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_sara <= s18;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and not x7 and not x8 and x11 ) = '1' then
         y9 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and not x7 and not x8 and not x11 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and not x7 and not x8 and not x11 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and not x7 and not x8 and not x11 and x16 and not x12 and not x13 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and x6 and not x7 and not x8 and not x11 and not x16 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and x7 and x11 ) = '1' then
         y9 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and x7 and not x11 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and x7 and not x11 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and x7 and not x11 and x16 and not x12 and not x13 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and x7 and not x11 and not x16 ) = '1' then
         current_sara <= s1;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and not x7 and x8 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_sara <= s19;

      elsif ( not x15 and not x3 and not x4 and x5 and not x6 and not x7 and not x8 ) = '1' then
         y37 <= '1' ;
         current_sara <= s14;

      elsif ( not x15 and not x3 and not x4 and not x5 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         current_sara <= s16;

      elsif ( not x15 and not x3 and not x4 and not x5 and not x9 and x6 ) = '1' then
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         current_sara <= s14;

      else
         y5 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      end if;

   when s14 =>
      if ( x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( x16 and not x12 and not x13 ) = '1' then
         current_sara <= s1;

      else
         current_sara <= s1;

      end if;

   when s15 =>
      if ( x9 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s20;

      elsif ( not x9 and x19 and x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s21;

      elsif ( not x9 and x19 and not x4 and x5 and x6 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s22;

      elsif ( not x9 and x19 and not x4 and x5 and x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_sara <= s23;

      elsif ( not x9 and x19 and not x4 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_sara <= s14;

      elsif ( not x9 and x19 and not x4 and not x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s24;

      else
         y4 <= '1' ;
         y20 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_sara <= s25;

      end if;

   when s16 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s24;

   when s17 =>
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s22;

   when s18 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_sara <= s23;

   when s19 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_sara <= s14;

   when s20 =>
      if ( x18 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         current_sara <= s26;

      else
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_sara <= s20;

      end if;

   when s21 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y19 <= '1' ;
         current_sara <= s27;

   when s22 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_sara <= s28;

   when s23 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y32 <= '1' ;
         current_sara <= s19;

   when s24 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y19 <= '1' ;
         current_sara <= s29;

   when s25 =>
      if ( x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s21;

      elsif ( not x4 and x5 and x6 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s22;

      elsif ( not x4 and x5 and x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_sara <= s23;

      elsif ( not x4 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_sara <= s14;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s24;

      end if;

   when s26 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         current_sara <= s30;

   when s27 =>
      if ( x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_sara <= s27;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         current_sara <= s31;

      end if;

   when s28 =>
      if ( x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y10 <= '1' ;
         current_sara <= s32;

      else
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_sara <= s28;

      end if;

   when s29 =>
      if ( x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_sara <= s33;

      else
         y5 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         y23 <= '1' ;
         y24 <= '1' ;
         current_sara <= s29;

      end if;

   when s30 =>
      if ( x19 and x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s21;

      elsif ( x19 and not x4 and x5 and x6 and x7 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s22;

      elsif ( x19 and not x4 and x5 and x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y27 <= '1' ;
         y30 <= '1' ;
         current_sara <= s23;

      elsif ( x19 and not x4 and x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y38 <= '1' ;
         current_sara <= s14;

      elsif ( x19 and not x4 and not x5 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         current_sara <= s24;

      else
         y4 <= '1' ;
         y20 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_sara <= s25;

      end if;

   when s31 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y23 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

   when s32 =>
         y24 <= '1' ;
         y25 <= '1' ;
         current_sara <= s34;

   when s33 =>
      if ( x5 ) = '1' then
         y5 <= '1' ;
         y23 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      else
         y5 <= '1' ;
         y23 <= '1' ;
         y32 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_sara <= s14;

      end if;

   when s34 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_sara <= s35;

   when s35 =>
         y3 <= '1' ;
         y17 <= '1' ;
         y27 <= '1' ;
         y29 <= '1' ;
         current_sara <= s36;

   when s36 =>
      if ( x14 and x16 and x12 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( x14 and x16 and not x12 and x13 ) = '1' then
         y31 <= '1' ;
         current_sara <= s1;

      elsif ( x14 and x16 and not x12 and not x13 ) = '1' then
         current_sara <= s1;

      elsif ( x14 and not x16 ) = '1' then
         current_sara <= s1;

      else
         y9 <= '1' ;
         current_sara <= s14;

      end if;

   end case;
   end proc_sara;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;

	current_sara <= s1;
      elsif (clk'event and clk ='1') then
        proc_sara;
      end if;
   end process;
end ARC;
