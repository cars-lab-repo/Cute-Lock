// Benchmark "./test_runs/structural2_16keys_5bits--s-120240927_165426/ITC99/b14_encrypted" written by ABC on Fri Sep 27 18:23:46 2024

module b14_encrypted  ( clock, 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
    ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_,
    ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_,
    ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_,
    ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG  );
  input  clock;
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, keyinput0, keyinput1, keyinput2, keyinput3,
    keyinput4;
  output ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_,
    ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_,
    ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_,
    ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG;
  reg IR_REG_0_, IR_REG_1_, IR_REG_2_, IR_REG_3_, IR_REG_4_, IR_REG_5_,
    IR_REG_6_, IR_REG_7_, IR_REG_8_, IR_REG_9_, IR_REG_10_, IR_REG_11_,
    IR_REG_12_, IR_REG_13_, IR_REG_14_, IR_REG_15_, IR_REG_16_, IR_REG_17_,
    IR_REG_18_, IR_REG_19_, IR_REG_20_, IR_REG_21_, IR_REG_22_, IR_REG_23_,
    IR_REG_24_, IR_REG_25_, IR_REG_26_, IR_REG_27_, IR_REG_28_, IR_REG_29_,
    IR_REG_30_, IR_REG_31_, D_REG_0_, D_REG_1_, D_REG_2_, D_REG_3_,
    D_REG_4_, D_REG_5_, D_REG_6_, D_REG_7_, D_REG_8_, D_REG_9_, D_REG_10_,
    D_REG_11_, D_REG_12_, D_REG_13_, D_REG_14_, D_REG_15_, D_REG_16_,
    D_REG_17_, D_REG_18_, D_REG_19_, D_REG_20_, D_REG_21_, D_REG_22_,
    D_REG_23_, D_REG_24_, D_REG_25_, D_REG_26_, D_REG_27_, D_REG_28_,
    D_REG_29_, D_REG_30_, D_REG_31_, REG0_REG_0_, REG0_REG_1_, REG0_REG_2_,
    REG0_REG_3_, REG0_REG_4_, REG0_REG_5_, REG0_REG_6_, REG0_REG_7_,
    REG0_REG_8_, REG0_REG_9_, REG0_REG_10_, REG0_REG_11_, REG0_REG_12_,
    REG0_REG_13_, REG0_REG_14_, REG0_REG_15_, REG0_REG_16_, REG0_REG_17_,
    REG0_REG_18_, REG0_REG_19_, REG0_REG_20_, REG0_REG_21_, REG0_REG_22_,
    REG0_REG_23_, REG0_REG_24_, REG0_REG_25_, REG0_REG_26_, REG0_REG_27_,
    REG0_REG_28_, REG0_REG_29_, REG0_REG_30_, REG0_REG_31_, REG1_REG_0_,
    REG1_REG_1_, REG1_REG_2_, REG1_REG_3_, REG1_REG_4_, REG1_REG_5_,
    REG1_REG_6_, REG1_REG_7_, REG1_REG_8_, REG1_REG_9_, REG1_REG_10_,
    REG1_REG_11_, REG1_REG_12_, REG1_REG_13_, REG1_REG_14_, REG1_REG_15_,
    REG1_REG_16_, REG1_REG_17_, REG1_REG_18_, REG1_REG_19_, REG1_REG_20_,
    REG1_REG_21_, REG1_REG_22_, REG1_REG_23_, REG1_REG_24_, REG1_REG_25_,
    REG1_REG_26_, REG1_REG_27_, REG1_REG_28_, REG1_REG_29_, REG1_REG_30_,
    REG1_REG_31_, REG2_REG_0_, REG2_REG_1_, REG2_REG_2_, REG2_REG_3_,
    REG2_REG_4_, REG2_REG_5_, REG2_REG_6_, REG2_REG_7_, REG2_REG_8_,
    REG2_REG_9_, REG2_REG_10_, REG2_REG_11_, REG2_REG_12_, REG2_REG_13_,
    REG2_REG_14_, REG2_REG_15_, REG2_REG_16_, REG2_REG_17_, REG2_REG_18_,
    REG2_REG_19_, REG2_REG_20_, REG2_REG_21_, REG2_REG_22_, REG2_REG_23_,
    REG2_REG_24_, REG2_REG_25_, REG2_REG_26_, REG2_REG_27_, REG2_REG_28_,
    REG2_REG_29_, REG2_REG_30_, REG2_REG_31_, ADDR_REG_19_, ADDR_REG_18_,
    ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_, ADDR_REG_14_, ADDR_REG_13_,
    ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_, ADDR_REG_9_, ADDR_REG_8_,
    ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_, ADDR_REG_4_, ADDR_REG_3_,
    ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_, DATAO_REG_0_, DATAO_REG_1_,
    DATAO_REG_2_, DATAO_REG_3_, DATAO_REG_4_, DATAO_REG_5_, DATAO_REG_6_,
    DATAO_REG_7_, DATAO_REG_8_, DATAO_REG_9_, DATAO_REG_10_, DATAO_REG_11_,
    DATAO_REG_12_, DATAO_REG_13_, DATAO_REG_14_, DATAO_REG_15_,
    DATAO_REG_16_, DATAO_REG_17_, DATAO_REG_18_, DATAO_REG_19_,
    DATAO_REG_20_, DATAO_REG_21_, DATAO_REG_22_, DATAO_REG_23_,
    DATAO_REG_24_, DATAO_REG_25_, DATAO_REG_26_, DATAO_REG_27_,
    DATAO_REG_28_, DATAO_REG_29_, DATAO_REG_30_, DATAO_REG_31_, B_REG,
    REG3_REG_15_, REG3_REG_26_, REG3_REG_6_, REG3_REG_18_, REG3_REG_2_,
    REG3_REG_11_, REG3_REG_22_, REG3_REG_13_, REG3_REG_20_, REG3_REG_0_,
    REG3_REG_9_, REG3_REG_4_, REG3_REG_24_, REG3_REG_17_, REG3_REG_5_,
    REG3_REG_16_, REG3_REG_25_, REG3_REG_12_, REG3_REG_21_, REG3_REG_1_,
    REG3_REG_8_, REG3_REG_28_, REG3_REG_19_, REG3_REG_3_, REG3_REG_10_,
    REG3_REG_23_, REG3_REG_14_, REG3_REG_27_, REG3_REG_7_, STATE_REG,
    RD_REG, WR_REG, Q_0, Q_1, Q_2, Q_3;
  wire new_R1222_U519, new_R1222_U518, new_R1222_U517, new_U3014, new_U3015,
    new_U3016, new_U3017, new_U3018, new_U3019, new_U3020, new_U3021,
    new_U3022, new_U3023, new_U3024, new_U3025, new_U3026, new_U3027,
    new_U3028, new_U3029, new_U3030, new_U3031, new_U3032, new_U3033,
    new_U3034, new_U3035, new_U3036, new_U3037, new_U3038, new_U3039,
    new_U3040, new_U3041, new_U3042, new_U3043, new_U3044, new_U3045,
    new_U3046, new_U3047, new_U3048, new_U3049, new_U3050, new_U3051,
    new_U3052, new_U3053, new_U3054, new_U3055, new_U3056, new_U3057,
    new_U3058, new_U3059, new_U3060, new_U3061, new_U3062, new_U3063,
    new_U3064, new_U3065, new_U3066, new_U3067, new_U3068, new_U3069,
    new_U3070, new_U3071, new_U3072, new_U3073, new_U3074, new_U3075,
    new_U3076, new_U3077, new_U3078, new_U3079, new_U3080, new_U3081,
    new_U3082, new_U3083, new_U3084, new_U3085, new_U3086, new_U3087,
    new_U3088, new_U3089, new_U3090, new_U3091, new_U3092, new_U3093,
    new_U3094, new_U3095, new_U3096, new_U3097, new_U3098, new_U3099,
    new_U3100, new_U3101, new_U3102, new_U3103, new_U3104, new_U3105,
    new_U3106, new_U3107, new_U3108, new_U3109, new_U3110, new_U3111,
    new_U3112, new_U3113, new_U3114, new_U3115, new_U3116, new_U3117,
    new_U3118, new_U3119, new_U3120, new_U3121, new_U3122, new_U3123,
    new_U3124, new_U3125, new_U3126, new_U3127, new_U3128, new_U3129,
    new_U3130, new_U3131, new_U3132, new_U3133, new_U3134, new_U3135,
    new_U3136, new_U3137, new_U3138, new_U3139, new_U3140, new_U3141,
    new_U3142, new_U3143, new_U3144, new_U3145, new_U3146, new_U3147,
    new_U3150, new_U3151, new_U3152, new_U3153, new_U3154, new_U3155,
    new_U3156, new_U3157, new_U3158, new_U3159, new_U3160, new_U3161,
    new_U3162, new_U3163, new_U3164, new_U3165, new_U3166, new_U3167,
    new_U3168, new_U3169, new_U3170, new_U3171, new_U3172, new_U3173,
    new_U3174, new_U3175, new_U3176, new_U3177, new_U3178, new_U3179,
    new_U3180, new_U3181, new_U3182, new_U3183, new_U3184, new_U3185,
    new_U3186, new_U3187, new_U3188, new_U3189, new_U3190, new_U3191,
    new_U3192, new_U3193, new_U3194, new_U3195, new_U3196, new_U3197,
    new_U3198, new_U3199, new_U3200, new_U3201, new_U3202, new_U3203,
    new_U3204, new_U3205, new_U3206, new_U3207, new_U3208, new_U3209,
    new_U3352, new_U3353, new_U3355, new_U3356, new_U3357, new_U3358,
    new_U3359, new_U3360, new_U3361, new_U3362, new_U3363, new_U3364,
    new_U3365, new_U3366, new_U3367, new_U3368, new_U3369, new_U3370,
    new_U3371, new_U3372, new_U3373, new_U3374, new_U3375, new_U3376,
    new_U3377, new_U3378, new_U3379, new_U3380, new_U3381, new_U3382,
    new_U3383, new_U3384, new_U3385, new_U3386, new_U3387, new_U3388,
    new_U3389, new_U3390, new_U3391, new_U3392, new_U3393, new_U3394,
    new_U3395, new_U3396, new_U3397, new_U3398, new_U3399, new_U3400,
    new_U3401, new_U3402, new_U3403, new_U3404, new_U3405, new_U3406,
    new_U3407, new_U3408, new_U3409, new_U3410, new_U3411, new_U3412,
    new_U3413, new_U3414, new_U3415, new_U3416, new_U3417, new_U3418,
    new_U3419, new_U3420, new_U3421, new_U3422, new_U3423, new_U3424,
    new_U3425, new_U3426, new_U3427, new_U3428, new_U3429, new_U3430,
    new_U3431, new_U3432, new_U3433, new_U3434, new_U3435, new_U3436,
    new_U3437, new_U3438, new_U3439, new_U3440, new_U3441, new_U3442,
    new_U3443, new_U3444, new_U3445, new_U3446, new_U3447, new_U3448,
    new_U3449, new_U3450, new_U3451, new_U3452, new_U3453, new_U3454,
    new_U3455, new_U3456, new_U3457, new_U3460, new_U3461, new_U3462,
    new_U3463, new_U3464, new_U3465, new_U3466, new_U3468, new_U3470,
    new_U3472, new_U3474, new_U3476, new_U3478, new_U3480, new_U3482,
    new_U3484, new_U3486, new_U3488, new_U3490, new_U3492, new_U3494,
    new_U3496, new_U3498, new_U3500, new_U3502, new_U3504, new_U3582,
    new_U3583, new_U3584, new_U3585, new_U3586, new_U3587, new_U3588,
    new_U3589, new_U3590, new_U3591, new_U3592, new_U3593, new_U3594,
    new_U3595, new_U3596, new_U3597, new_U3598, new_U3599, new_U3600,
    new_U3601, new_U3602, new_U3603, new_U3604, new_U3605, new_U3606,
    new_U3607, new_U3608, new_U3609, new_U3610, new_U3611, new_U3612,
    new_U3613, new_U3614, new_U3615, new_U3616, new_U3617, new_U3618,
    new_U3619, new_U3620, new_U3621, new_U3622, new_U3623, new_U3624,
    new_U3625, new_U3626, new_U3627, new_U3628, new_U3629, new_U3630,
    new_U3631, new_U3632, new_U3633, new_U3634, new_U3635, new_U3636,
    new_U3637, new_U3638, new_U3639, new_U3640, new_U3641, new_U3642,
    new_U3643, new_U3644, new_U3645, new_U3646, new_U3647, new_U3648,
    new_U3649, new_U3650, new_U3651, new_U3652, new_U3653, new_U3654,
    new_U3655, new_U3656, new_U3657, new_U3658, new_U3659, new_U3660,
    new_U3661, new_U3662, new_U3663, new_U3664, new_U3665, new_U3666,
    new_U3667, new_U3668, new_U3669, new_U3670, new_U3671, new_U3672,
    new_U3673, new_U3674, new_U3675, new_U3676, new_U3677, new_U3678,
    new_U3679, new_U3680, new_U3681, new_U3682, new_U3683, new_U3684,
    new_U3685, new_U3686, new_U3687, new_U3688, new_U3689, new_U3690,
    new_U3691, new_U3692, new_U3693, new_U3694, new_U3695, new_U3696,
    new_U3697, new_U3698, new_U3699, new_U3700, new_U3701, new_U3702,
    new_U3703, new_U3704, new_U3705, new_U3706, new_U3707, new_U3708,
    new_U3709, new_U3710, new_U3711, new_U3712, new_U3713, new_U3714,
    new_U3715, new_U3716, new_U3717, new_U3718, new_U3719, new_U3720,
    new_U3721, new_U3722, new_U3723, new_U3724, new_U3725, new_U3726,
    new_U3727, new_U3728, new_U3729, new_U3730, new_U3731, new_U3732,
    new_U3733, new_U3734, new_U3735, new_U3736, new_U3737, new_U3738,
    new_U3739, new_U3740, new_U3741, new_U3742, new_U3743, new_U3744,
    new_U3745, new_U3746, new_U3747, new_U3748, new_U3749, new_U3750,
    new_U3751, new_U3752, new_U3753, new_U3754, new_U3755, new_U3756,
    new_U3757, new_U3758, new_U3759, new_U3760, new_U3761, new_U3762,
    new_U3763, new_U3764, new_U3765, new_U3766, new_U3767, new_U3768,
    new_U3769, new_U3770, new_U3771, new_U3772, new_U3773, new_U3774,
    new_U3775, new_U3776, new_U3777, new_U3778, new_U3779, new_U3780,
    new_U3781, new_U3782, new_U3783, new_U3784, new_U3785, new_U3786,
    new_U3787, new_U3788, new_U3789, new_U3790, new_U3791, new_U3792,
    new_U3793, new_U3794, new_U3795, new_U3796, new_U3797, new_U3798,
    new_U3799, new_U3800, new_U3801, new_U3802, new_U3803, new_U3804,
    new_U3805, new_U3806, new_U3807, new_U3808, new_U3809, new_U3810,
    new_U3811, new_U3812, new_U3813, new_U3814, new_U3815, new_U3816,
    new_U3817, new_U3818, new_U3819, new_U3820, new_U3821, new_U3822,
    new_U3823, new_U3824, new_U3825, new_U3826, new_U3827, new_U3828,
    new_U3829, new_U3830, new_U3831, new_U3832, new_U3833, new_U3834,
    new_U3835, new_U3836, new_U3837, new_U3838, new_U3839, new_U3840,
    new_U3841, new_U3842, new_U3843, new_U3844, new_U3845, new_U3846,
    new_U3847, new_U3848, new_U3849, new_U3850, new_U3851, new_U3852,
    new_U3853, new_U3854, new_U3855, new_U3856, new_U3857, new_U3858,
    new_U3859, new_U3860, new_U3861, new_U3862, new_U3863, new_U3864,
    new_U3865, new_U3866, new_U3867, new_U3868, new_U3869, new_U3870,
    new_U3871, new_U3872, new_U3873, new_U3874, new_U3875, new_U3876,
    new_U3877, new_U3878, new_U3879, new_U3880, new_U3881, new_U3882,
    new_U3883, new_U3884, new_U3885, new_U3886, new_U3887, new_U3888,
    new_U3889, new_U3890, new_U3891, new_U3892, new_U3893, new_U3894,
    new_U3895, new_U3896, new_U3897, new_U3898, new_U3899, new_U3900,
    new_U3901, new_U3902, new_U3903, new_U3904, new_U3905, new_U3906,
    new_U3907, new_U3908, new_U3909, new_U3910, new_U3911, new_U3912,
    new_U3913, new_U3914, new_U3915, new_U3916, new_U3917, new_U3918,
    new_U3919, new_U3920, new_U3921, new_U3922, new_U3923, new_U3924,
    new_U3925, new_U3926, new_U3927, new_U3928, new_U3929, new_U3930,
    new_U3931, new_U3932, new_U3933, new_U3934, new_U3935, new_U3936,
    new_U3937, new_U3938, new_U3939, new_U3940, new_U3941, new_U3942,
    new_U3943, new_U3944, new_U3945, new_U3946, new_U3947, new_U3948,
    new_U3949, new_U3950, new_U3951, new_U3952, new_U3953, new_U3954,
    new_U3955, new_U3956, new_U3957, new_U3958, new_U3959, new_U3960,
    new_U3961, new_U3962, new_U3963, new_U3964, new_U3965, new_U3966,
    new_U3967, new_U3968, new_U3969, new_U3970, new_U3971, new_U3972,
    new_U3973, new_U3974, new_U3975, new_U3976, new_U3977, new_U3978,
    new_U3979, new_U3980, new_U3981, new_U3982, new_U3983, new_U3984,
    new_U3985, new_U3986, new_U3987, new_U3988, new_U3989, new_U3990,
    new_U3991, new_U3992, new_U3993, new_U3994, new_U3995, new_U3996,
    new_U3997, new_U3998, new_U3999, new_U4000, new_U4001, new_U4002,
    new_U4003, new_U4004, new_U4005, new_U4006, new_U4007, new_U4008,
    new_U4009, new_U4010, new_U4011, new_U4012, new_U4013, new_U4014,
    new_U4015, new_U4016, new_U4017, new_U4018, new_U4019, new_U4020,
    new_U4021, new_U4022, new_U4023, new_U4024, new_U4025, new_U4026,
    new_U4027, new_U4028, new_U4029, new_U4030, new_U4031, new_U4032,
    new_U4033, new_U4034, new_U4035, new_U4036, new_U4037, new_U4038,
    new_U4039, new_U4040, new_U4041, new_U4042, new_U4044, new_U4045,
    new_U4046, new_U4047, new_U4048, new_U4049, new_U4050, new_U4051,
    new_U4052, new_U4053, new_U4054, new_U4055, new_U4056, new_U4057,
    new_U4058, new_U4059, new_U4060, new_U4061, new_U4062, new_U4063,
    new_U4064, new_U4065, new_U4066, new_U4067, new_U4068, new_U4069,
    new_U4070, new_U4071, new_U4072, new_U4073, new_U4074, new_U4075,
    new_U4076, new_U4077, new_U4078, new_U4079, new_U4080, new_U4081,
    new_U4082, new_U4083, new_U4084, new_U4085, new_U4086, new_U4087,
    new_U4088, new_U4089, new_U4090, new_U4091, new_U4092, new_U4093,
    new_U4094, new_U4095, new_U4096, new_U4097, new_U4098, new_U4099,
    new_U4100, new_U4101, new_U4102, new_U4103, new_U4104, new_U4105,
    new_U4106, new_U4107, new_U4108, new_U4109, new_U4110, new_U4111,
    new_U4112, new_U4113, new_U4114, new_U4115, new_U4116, new_U4117,
    new_U4118, new_U4119, new_U4120, new_U4121, new_U4122, new_U4123,
    new_U4124, new_U4125, new_U4126, new_U4127, new_U4128, new_U4129,
    new_U4130, new_U4131, new_U4132, new_U4133, new_U4134, new_U4135,
    new_U4136, new_U4137, new_U4138, new_U4139, new_U4140, new_U4141,
    new_U4142, new_U4143, new_U4144, new_U4145, new_U4146, new_U4147,
    new_U4148, new_U4149, new_U4150, new_U4151, new_U4152, new_U4153,
    new_U4154, new_U4155, new_U4156, new_U4157, new_U4158, new_U4159,
    new_U4160, new_U4161, new_U4162, new_U4163, new_U4164, new_U4165,
    new_U4166, new_U4167, new_U4168, new_U4169, new_U4170, new_U4171,
    new_U4172, new_U4173, new_U4174, new_U4175, new_U4176, new_U4177,
    new_U4178, new_U4179, new_U4180, new_U4181, new_U4182, new_U4183,
    new_U4184, new_U4185, new_U4186, new_U4187, new_U4188, new_U4189,
    new_U4190, new_U4191, new_U4192, new_U4193, new_U4194, new_U4195,
    new_U4196, new_U4197, new_U4198, new_U4199, new_U4200, new_U4201,
    new_U4202, new_U4203, new_U4204, new_U4205, new_U4206, new_U4207,
    new_U4208, new_U4209, new_U4210, new_U4211, new_U4212, new_U4213,
    new_U4214, new_U4215, new_U4216, new_U4217, new_U4218, new_U4219,
    new_U4220, new_U4221, new_U4222, new_U4223, new_U4224, new_U4225,
    new_U4226, new_U4227, new_U4228, new_U4229, new_U4230, new_U4231,
    new_U4232, new_U4233, new_U4234, new_U4235, new_U4236, new_U4237,
    new_U4238, new_U4239, new_U4240, new_U4241, new_U4242, new_U4243,
    new_U4244, new_U4245, new_U4246, new_U4247, new_U4248, new_U4249,
    new_U4250, new_U4251, new_U4252, new_U4253, new_U4254, new_U4255,
    new_U4256, new_U4257, new_U4258, new_U4259, new_U4260, new_U4261,
    new_U4262, new_U4263, new_U4264, new_U4265, new_U4266, new_U4267,
    new_U4268, new_U4269, new_U4270, new_U4271, new_U4272, new_U4273,
    new_U4274, new_U4275, new_U4276, new_U4277, new_U4278, new_U4279,
    new_U4280, new_U4281, new_U4282, new_U4283, new_U4284, new_U4285,
    new_U4286, new_U4287, new_U4288, new_U4289, new_U4290, new_U4291,
    new_U4292, new_U4293, new_U4294, new_U4295, new_U4296, new_U4297,
    new_U4298, new_U4299, new_U4300, new_U4301, new_U4302, new_U4303,
    new_U4304, new_U4305, new_U4306, new_U4307, new_U4308, new_U4309,
    new_U4310, new_U4311, new_U4312, new_U4313, new_U4314, new_U4315,
    new_U4316, new_U4317, new_U4318, new_U4319, new_U4320, new_U4321,
    new_U4322, new_U4323, new_U4324, new_U4325, new_U4326, new_U4327,
    new_U4328, new_U4329, new_U4330, new_U4331, new_U4332, new_U4333,
    new_U4334, new_U4335, new_U4336, new_U4337, new_U4338, new_U4339,
    new_U4340, new_U4341, new_U4342, new_U4343, new_U4344, new_U4345,
    new_U4346, new_U4347, new_U4348, new_U4349, new_U4350, new_U4351,
    new_U4352, new_U4353, new_U4354, new_U4355, new_U4356, new_U4357,
    new_U4358, new_U4359, new_U4360, new_U4361, new_U4362, new_U4363,
    new_U4364, new_U4365, new_U4366, new_U4367, new_U4368, new_U4369,
    new_U4370, new_U4371, new_U4372, new_U4373, new_U4374, new_U4375,
    new_U4376, new_U4377, new_U4378, new_U4379, new_U4380, new_U4381,
    new_U4382, new_U4383, new_U4384, new_U4385, new_U4386, new_U4387,
    new_U4388, new_U4389, new_U4390, new_U4391, new_U4392, new_U4393,
    new_U4394, new_U4395, new_U4396, new_U4397, new_U4398, new_U4399,
    new_U4400, new_U4401, new_U4402, new_U4403, new_U4404, new_U4405,
    new_U4406, new_U4407, new_U4408, new_U4409, new_U4410, new_U4411,
    new_U4412, new_U4413, new_U4414, new_U4415, new_U4416, new_U4417,
    new_U4418, new_U4419, new_U4420, new_U4421, new_U4422, new_U4423,
    new_U4424, new_U4425, new_U4426, new_U4427, new_U4428, new_U4429,
    new_U4430, new_U4431, new_U4432, new_U4433, new_U4434, new_U4435,
    new_U4436, new_U4437, new_U4438, new_U4439, new_U4440, new_U4441,
    new_U4442, new_U4443, new_U4444, new_U4445, new_U4446, new_U4447,
    new_U4448, new_U4449, new_U4450, new_U4451, new_U4452, new_U4453,
    new_U4454, new_U4455, new_U4456, new_U4457, new_U4458, new_U4459,
    new_U4460, new_U4461, new_U4462, new_U4463, new_U4464, new_U4465,
    new_U4466, new_U4467, new_U4468, new_U4469, new_U4470, new_U4471,
    new_U4472, new_U4473, new_U4474, new_U4475, new_U4476, new_U4477,
    new_U4478, new_U4479, new_U4480, new_U4481, new_U4482, new_U4483,
    new_U4484, new_U4485, new_U4486, new_U4487, new_U4488, new_U4489,
    new_U4490, new_U4491, new_U4492, new_U4493, new_U4494, new_U4495,
    new_U4496, new_U4497, new_U4498, new_U4499, new_U4500, new_U4501,
    new_U4502, new_U4503, new_U4504, new_U4505, new_U4506, new_U4507,
    new_U4508, new_U4509, new_U4510, new_U4511, new_U4512, new_U4513,
    new_U4514, new_U4515, new_U4516, new_U4517, new_U4518, new_U4519,
    new_U4520, new_U4521, new_U4522, new_U4523, new_U4524, new_U4525,
    new_U4526, new_U4527, new_U4528, new_U4529, new_U4530, new_U4531,
    new_U4532, new_U4533, new_U4534, new_U4535, new_U4536, new_U4537,
    new_U4538, new_U4539, new_U4540, new_U4541, new_U4542, new_U4543,
    new_U4544, new_U4545, new_U4546, new_U4547, new_U4548, new_U4549,
    new_U4550, new_U4551, new_U4552, new_U4553, new_U4554, new_U4555,
    new_U4556, new_U4557, new_U4558, new_U4559, new_U4560, new_U4561,
    new_U4562, new_U4563, new_U4564, new_U4565, new_U4566, new_U4567,
    new_U4568, new_U4569, new_U4570, new_U4571, new_U4572, new_U4573,
    new_U4574, new_U4575, new_U4576, new_U4577, new_U4578, new_U4579,
    new_U4580, new_U4581, new_U4582, new_U4583, new_U4584, new_U4585,
    new_U4586, new_U4587, new_U4588, new_U4589, new_U4590, new_U4591,
    new_U4592, new_U4593, new_U4594, new_U4595, new_U4596, new_U4597,
    new_U4598, new_U4599, new_U4600, new_U4601, new_U4602, new_U4603,
    new_U4604, new_U4605, new_U4606, new_U4607, new_U4608, new_U4609,
    new_U4610, new_U4611, new_U4612, new_U4613, new_U4614, new_U4615,
    new_U4616, new_U4617, new_U4618, new_U4619, new_U4620, new_U4621,
    new_U4622, new_U4623, new_U4624, new_U4625, new_U4626, new_U4627,
    new_U4628, new_U4629, new_U4630, new_U4631, new_U4632, new_U4633,
    new_U4634, new_U4635, new_U4636, new_U4637, new_U4638, new_U4639,
    new_U4640, new_U4641, new_U4642, new_U4643, new_U4644, new_U4645,
    new_U4646, new_U4647, new_U4648, new_U4649, new_U4650, new_U4651,
    new_U4652, new_U4653, new_U4654, new_U4655, new_U4656, new_U4657,
    new_U4658, new_U4659, new_U4660, new_U4661, new_U4662, new_U4663,
    new_U4664, new_U4665, new_U4666, new_U4667, new_U4668, new_U4669,
    new_U4670, new_U4671, new_U4672, new_U4673, new_U4674, new_U4675,
    new_U4676, new_U4677, new_U4678, new_U4679, new_U4680, new_U4681,
    new_U4682, new_U4683, new_U4684, new_U4685, new_U4686, new_U4687,
    new_U4688, new_U4689, new_U4690, new_U4691, new_U4692, new_U4693,
    new_U4694, new_U4695, new_U4696, new_U4697, new_U4698, new_U4699,
    new_U4700, new_U4701, new_U4702, new_U4703, new_U4704, new_U4705,
    new_U4706, new_U4707, new_U4708, new_U4709, new_U4710, new_U4711,
    new_U4712, new_U4713, new_U4714, new_U4715, new_U4716, new_U4717,
    new_U4718, new_U4719, new_U4720, new_U4721, new_U4722, new_U4723,
    new_U4724, new_U4725, new_U4726, new_U4727, new_U4728, new_U4729,
    new_U4730, new_U4731, new_U4732, new_U4733, new_U4734, new_U4735,
    new_U4736, new_U4737, new_U4738, new_U4739, new_U4740, new_U4741,
    new_U4742, new_U4743, new_U4744, new_U4745, new_U4746, new_U4747,
    new_U4748, new_U4749, new_U4750, new_U4751, new_U4752, new_U4753,
    new_U4754, new_U4755, new_U4756, new_U4757, new_U4758, new_U4759,
    new_U4760, new_U4761, new_U4762, new_U4763, new_U4764, new_U4765,
    new_U4766, new_U4767, new_U4768, new_U4769, new_U4770, new_U4771,
    new_U4772, new_U4773, new_U4774, new_U4775, new_U4776, new_U4777,
    new_U4778, new_U4779, new_U4780, new_U4781, new_U4782, new_U4783,
    new_U4784, new_U4785, new_U4786, new_U4787, new_U4788, new_U4789,
    new_U4790, new_U4791, new_U4792, new_U4793, new_U4794, new_U4795,
    new_U4796, new_U4797, new_U4798, new_U4799, new_U4800, new_U4801,
    new_U4802, new_U4803, new_U4804, new_U4805, new_U4806, new_U4807,
    new_U4808, new_U4809, new_U4810, new_U4811, new_U4812, new_U4813,
    new_U4814, new_U4815, new_U4816, new_U4817, new_U4818, new_U4819,
    new_U4820, new_U4821, new_U4822, new_U4823, new_U4824, new_U4825,
    new_U4826, new_U4827, new_U4828, new_U4829, new_U4830, new_U4831,
    new_U4832, new_U4833, new_U4834, new_U4835, new_U4836, new_U4837,
    new_U4838, new_U4839, new_U4840, new_U4841, new_U4842, new_U4843,
    new_U4844, new_U4845, new_U4846, new_U4847, new_U4848, new_U4849,
    new_U4850, new_U4851, new_U4852, new_U4853, new_U4854, new_U4855,
    new_U4856, new_U4857, new_U4858, new_U4859, new_U4860, new_U4861,
    new_U4862, new_U4863, new_U4864, new_U4865, new_U4866, new_U4867,
    new_U4868, new_U4869, new_U4870, new_U4871, new_U4872, new_U4873,
    new_U4874, new_U4875, new_U4876, new_U4877, new_U4878, new_U4879,
    new_U4880, new_U4881, new_U4882, new_U4883, new_U4884, new_U4885,
    new_U4886, new_U4887, new_U4888, new_U4889, new_U4890, new_U4891,
    new_U4892, new_U4893, new_U4894, new_U4895, new_U4896, new_U4897,
    new_U4898, new_U4899, new_U4900, new_U4901, new_U4902, new_U4903,
    new_U4904, new_U4905, new_U4906, new_U4907, new_U4908, new_U4909,
    new_U4910, new_U4911, new_U4912, new_U4913, new_U4914, new_U4915,
    new_U4916, new_U4917, new_U4918, new_U4919, new_U4920, new_U4921,
    new_U4922, new_U4923, new_U4924, new_U4925, new_U4926, new_U4927,
    new_U4928, new_U4929, new_U4930, new_U4931, new_U4932, new_U4933,
    new_U4934, new_U4935, new_U4936, new_U4937, new_U4938, new_U4939,
    new_U4940, new_U4941, new_U4942, new_U4943, new_U4944, new_U4945,
    new_U4946, new_U4947, new_U4948, new_U4949, new_U4950, new_U4951,
    new_U4952, new_U4953, new_U4954, new_U4955, new_U4956, new_U4957,
    new_U4958, new_U4959, new_U4960, new_U4961, new_U4962, new_U4963,
    new_U4964, new_U4965, new_U4966, new_U4967, new_U4968, new_U4969,
    new_U4970, new_U4971, new_U4972, new_U4973, new_U4974, new_U4975,
    new_U4976, new_U4977, new_U4978, new_U4979, new_U4980, new_U4981,
    new_U4982, new_U4983, new_U4984, new_U4985, new_U4986, new_U4987,
    new_U4988, new_U4989, new_U4990, new_U4991, new_U4992, new_U4993,
    new_U4994, new_U4995, new_U4996, new_U4997, new_U4998, new_U4999,
    new_U5000, new_U5001, new_U5002, new_U5003, new_U5004, new_U5005,
    new_U5006, new_U5007, new_U5008, new_U5009, new_U5010, new_U5011,
    new_U5012, new_U5013, new_U5014, new_U5015, new_U5016, new_U5017,
    new_U5018, new_U5019, new_U5020, new_U5021, new_U5022, new_U5023,
    new_U5024, new_U5025, new_U5026, new_U5027, new_U5028, new_U5029,
    new_U5030, new_U5031, new_U5032, new_U5033, new_U5034, new_U5035,
    new_U5036, new_U5037, new_U5038, new_U5039, new_U5040, new_U5041,
    new_U5042, new_U5043, new_U5044, new_U5045, new_U5046, new_U5047,
    new_U5048, new_U5049, new_U5050, new_U5051, new_U5052, new_U5053,
    new_U5054, new_U5055, new_U5056, new_U5057, new_U5058, new_U5059,
    new_U5060, new_U5061, new_U5062, new_U5063, new_U5064, new_U5065,
    new_U5066, new_U5067, new_U5068, new_U5069, new_U5070, new_U5071,
    new_U5072, new_U5073, new_U5074, new_U5075, new_U5076, new_U5077,
    new_U5078, new_U5079, new_U5080, new_U5081, new_U5082, new_U5083,
    new_U5084, new_U5085, new_U5086, new_U5087, new_U5088, new_U5089,
    new_U5090, new_U5091, new_U5092, new_U5093, new_U5094, new_U5095,
    new_U5096, new_U5097, new_U5098, new_U5099, new_U5100, new_U5101,
    new_U5102, new_U5103, new_U5104, new_U5105, new_U5106, new_U5107,
    new_U5108, new_U5109, new_U5110, new_U5111, new_U5112, new_U5113,
    new_U5114, new_U5115, new_U5116, new_U5117, new_U5118, new_U5119,
    new_U5120, new_U5121, new_U5122, new_U5123, new_U5124, new_U5125,
    new_U5126, new_U5127, new_U5128, new_U5129, new_U5130, new_U5131,
    new_U5132, new_U5133, new_U5134, new_U5135, new_U5136, new_U5137,
    new_U5138, new_U5139, new_U5140, new_U5141, new_U5142, new_U5143,
    new_U5144, new_U5145, new_U5146, new_U5147, new_U5148, new_U5149,
    new_U5150, new_U5151, new_U5152, new_U5153, new_U5154, new_U5155,
    new_U5156, new_U5157, new_U5158, new_U5159, new_U5160, new_U5161,
    new_U5162, new_U5163, new_U5164, new_U5165, new_U5166, new_U5167,
    new_U5168, new_U5169, new_U5170, new_U5171, new_U5172, new_U5173,
    new_U5174, new_U5175, new_U5176, new_U5177, new_U5178, new_U5179,
    new_U5180, new_U5181, new_U5182, new_U5183, new_U5184, new_U5185,
    new_U5186, new_U5187, new_U5188, new_U5189, new_U5190, new_U5191,
    new_U5192, new_U5193, new_U5194, new_U5195, new_U5196, new_U5197,
    new_U5198, new_U5199, new_U5200, new_U5201, new_U5202, new_U5203,
    new_U5204, new_U5205, new_U5206, new_U5207, new_U5208, new_U5209,
    new_U5210, new_U5211, new_U5212, new_U5213, new_U5214, new_U5215,
    new_U5216, new_U5217, new_U5218, new_U5219, new_U5220, new_U5221,
    new_U5222, new_U5223, new_U5224, new_U5225, new_U5226, new_U5227,
    new_U5228, new_U5229, new_U5230, new_U5231, new_U5232, new_U5233,
    new_U5234, new_U5235, new_U5236, new_U5237, new_U5238, new_U5239,
    new_U5240, new_U5241, new_U5242, new_U5243, new_U5244, new_U5245,
    new_U5246, new_U5247, new_U5248, new_U5249, new_U5250, new_U5251,
    new_U5252, new_U5253, new_U5254, new_U5255, new_U5256, new_U5257,
    new_U5258, new_U5259, new_U5260, new_U5261, new_U5262, new_U5263,
    new_U5264, new_U5265, new_U5266, new_U5267, new_U5268, new_U5269,
    new_U5270, new_U5271, new_U5272, new_U5273, new_U5274, new_U5275,
    new_U5276, new_U5277, new_U5278, new_U5279, new_U5280, new_U5281,
    new_U5282, new_U5283, new_U5284, new_U5285, new_U5286, new_U5287,
    new_U5288, new_U5289, new_U5290, new_U5291, new_U5292, new_U5293,
    new_U5294, new_U5295, new_U5296, new_U5297, new_U5298, new_U5299,
    new_U5300, new_U5301, new_U5302, new_U5303, new_U5304, new_U5305,
    new_U5306, new_U5307, new_U5308, new_U5309, new_U5310, new_U5311,
    new_U5312, new_U5313, new_U5314, new_U5315, new_U5316, new_U5317,
    new_U5318, new_U5319, new_U5320, new_U5321, new_U5322, new_U5323,
    new_U5324, new_U5325, new_U5326, new_U5327, new_U5328, new_U5329,
    new_U5330, new_U5331, new_U5332, new_U5333, new_U5334, new_U5335,
    new_U5336, new_U5337, new_U5338, new_U5339, new_U5340, new_U5341,
    new_U5342, new_U5343, new_U5344, new_U5345, new_U5346, new_U5347,
    new_U5348, new_U5349, new_U5350, new_U5351, new_U5352, new_U5353,
    new_U5354, new_U5355, new_U5356, new_U5357, new_U5358, new_U5359,
    new_U5360, new_U5361, new_U5362, new_U5363, new_U5364, new_U5365,
    new_U5366, new_U5367, new_U5368, new_U5369, new_U5370, new_U5371,
    new_U5372, new_U5373, new_U5374, new_U5375, new_U5376, new_U5377,
    new_U5378, new_U5379, new_U5380, new_U5381, new_U5382, new_U5383,
    new_U5384, new_U5385, new_U5386, new_U5387, new_U5388, new_U5389,
    new_U5390, new_U5391, new_U5392, new_U5393, new_U5394, new_U5395,
    new_U5396, new_U5397, new_U5398, new_U5399, new_U5400, new_U5401,
    new_U5402, new_U5403, new_U5404, new_U5405, new_U5406, new_U5407,
    new_U5408, new_U5409, new_U5410, new_U5411, new_U5412, new_U5413,
    new_U5414, new_U5415, new_U5416, new_U5417, new_U5418, new_U5419,
    new_U5420, new_U5421, new_U5422, new_U5423, new_U5424, new_U5425,
    new_U5426, new_U5427, new_U5428, new_U5429, new_U5430, new_U5431,
    new_U5432, new_U5433, new_U5434, new_U5435, new_U5436, new_U5437,
    new_U5438, new_U5439, new_U5440, new_U5441, new_U5442, new_U5443,
    new_U5444, new_U5445, new_U5446, new_U5447, new_U5448, new_U5449,
    new_U5450, new_U5451, new_U5452, new_U5453, new_U5454, new_U5455,
    new_U5456, new_U5457, new_U5458, new_U5459, new_U5460, new_U5461,
    new_U5462, new_U5463, new_U5464, new_U5465, new_U5466, new_U5467,
    new_U5468, new_U5469, new_U5470, new_U5471, new_U5472, new_U5473,
    new_U5474, new_U5475, new_U5476, new_U5477, new_U5478, new_U5479,
    new_U5480, new_U5481, new_U5482, new_U5483, new_U5484, new_U5485,
    new_U5486, new_U5487, new_U5488, new_U5489, new_U5490, new_U5491,
    new_U5492, new_U5493, new_U5494, new_U5495, new_U5496, new_U5497,
    new_U5498, new_U5499, new_U5500, new_U5501, new_U5502, new_U5503,
    new_U5504, new_U5505, new_U5506, new_U5507, new_U5508, new_U5509,
    new_U5510, new_U5511, new_U5512, new_U5513, new_U5514, new_U5515,
    new_U5516, new_U5517, new_U5518, new_U5519, new_U5520, new_U5521,
    new_U5522, new_U5523, new_U5524, new_U5525, new_U5526, new_U5527,
    new_U5528, new_U5529, new_U5530, new_U5531, new_U5532, new_U5533,
    new_U5534, new_U5535, new_U5536, new_U5537, new_U5538, new_U5539,
    new_U5540, new_U5541, new_U5542, new_U5543, new_U5544, new_U5545,
    new_U5546, new_U5547, new_U5548, new_U5549, new_U5550, new_U5551,
    new_U5552, new_U5553, new_U5554, new_U5555, new_U5556, new_U5557,
    new_U5558, new_U5559, new_U5560, new_U5561, new_U5562, new_U5563,
    new_U5564, new_U5565, new_U5566, new_U5567, new_U5568, new_U5569,
    new_U5570, new_U5571, new_U5572, new_U5573, new_U5574, new_U5575,
    new_U5576, new_U5577, new_U5578, new_U5579, new_U5580, new_U5581,
    new_U5582, new_U5583, new_U5584, new_U5585, new_U5586, new_U5587,
    new_U5588, new_U5589, new_U5590, new_U5591, new_U5592, new_U5593,
    new_U5594, new_U5595, new_U5596, new_U5597, new_U5598, new_U5599,
    new_U5600, new_U5601, new_U5602, new_U5603, new_U5604, new_U5605,
    new_U5606, new_U5607, new_U5608, new_U5609, new_U5610, new_U5611,
    new_U5612, new_U5613, new_U5614, new_U5615, new_U5616, new_U5617,
    new_U5618, new_U5619, new_U5620, new_U5621, new_U5622, new_U5623,
    new_U5624, new_U5625, new_U5626, new_U5627, new_U5628, new_U5629,
    new_U5630, new_U5631, new_U5632, new_U5633, new_U5634, new_U5635,
    new_U5636, new_U5637, new_U5638, new_U5639, new_U5640, new_U5641,
    new_U5642, new_U5643, new_U5644, new_U5645, new_U5646, new_U5647,
    new_U5648, new_U5649, new_U5650, new_U5651, new_U5652, new_U5653,
    new_U5654, new_U5655, new_U5656, new_U5657, new_U5658, new_U5659,
    new_U5660, new_U5661, new_U5662, new_U5663, new_U5664, new_U5665,
    new_U5666, new_U5667, new_U5668, new_U5669, new_U5670, new_U5671,
    new_U5672, new_U5673, new_U5674, new_U5675, new_U5676, new_U5677,
    new_U5678, new_U5679, new_U5680, new_U5681, new_U5682, new_U5683,
    new_U5684, new_U5685, new_U5686, new_U5687, new_U5688, new_U5689,
    new_U5690, new_U5691, new_U5692, new_U5693, new_U5694, new_U5695,
    new_U5696, new_U5697, new_U5698, new_U5699, new_U5700, new_U5701,
    new_U5702, new_U5703, new_U5704, new_U5705, new_U5706, new_U5707,
    new_U5708, new_U5709, new_U5710, new_U5711, new_U5712, new_U5713,
    new_U5714, new_U5715, new_U5716, new_U5717, new_U5718, new_U5719,
    new_U5720, new_U5721, new_U5722, new_U5723, new_U5724, new_U5725,
    new_U5726, new_U5727, new_U5728, new_U5729, new_U5730, new_U5731,
    new_U5732, new_U5733, new_U5734, new_U5735, new_U5736, new_U5737,
    new_U5738, new_U5739, new_U5740, new_U5741, new_U5742, new_U5743,
    new_U5744, new_U5745, new_U5746, new_U5747, new_U5748, new_U5749,
    new_U5750, new_U5751, new_U5752, new_U5753, new_U5754, new_U5755,
    new_U5756, new_U5757, new_U5758, new_U5759, new_U5760, new_U5761,
    new_U5762, new_U5763, new_U5764, new_U5765, new_U5766, new_U5767,
    new_U5768, new_U5769, new_U5770, new_U5771, new_U5772, new_U5773,
    new_U5774, new_U5775, new_U5776, new_U5777, new_U5778, new_U5779,
    new_U5780, new_U5781, new_U5782, new_U5783, new_U5784, new_U5785,
    new_U5786, new_U5787, new_U5788, new_U5789, new_U5790, new_U5791,
    new_U5792, new_U5793, new_U5794, new_U5795, new_U5796, new_U5797,
    new_U5798, new_U5799, new_U5800, new_U5801, new_U5802, new_U5803,
    new_U5804, new_U5805, new_U5806, new_U5807, new_U5808, new_U5809,
    new_U5810, new_U5811, new_U5812, new_U5813, new_U5814, new_U5815,
    new_U5816, new_U5817, new_U5818, new_U5819, new_U5820, new_U5821,
    new_U5822, new_U5823, new_U5824, new_U5825, new_U5826, new_U5827,
    new_U5828, new_U5829, new_U5830, new_U5831, new_U5832, new_U5833,
    new_U5834, new_U5835, new_U5836, new_U5837, new_U5838, new_U5839,
    new_U5840, new_U5841, new_U5842, new_U5843, new_U5844, new_U5845,
    new_U5846, new_U5847, new_U5848, new_U5849, new_U5850, new_U5851,
    new_U5852, new_U5853, new_U5854, new_U5855, new_U5856, new_U5857,
    new_U5858, new_U5859, new_U5860, new_U5861, new_U5862, new_U5863,
    new_U5864, new_U5865, new_U5866, new_U5867, new_U5868, new_U5869,
    new_U5870, new_U5871, new_U5872, new_U5873, new_U5874, new_U5875,
    new_U5876, new_U5877, new_U5878, new_U5879, new_U5880, new_U5881,
    new_U5882, new_U5883, new_U5884, new_U5885, new_U5886, new_U5887,
    new_U5888, new_U5889, new_U5890, new_U5891, new_U5892, new_U5893,
    new_U5894, new_U5895, new_U5896, new_U5897, new_U5898, new_U5899,
    new_U5900, new_U5901, new_U5902, new_U5903, new_U5904, new_U5905,
    new_U5906, new_U5907, new_U5908, new_U5909, new_U5910, new_U5911,
    new_U5912, new_U5913, new_U5914, new_U5915, new_U5916, new_U5917,
    new_U5918, new_U5919, new_U5920, new_U5921, new_U5922, new_U5923,
    new_U5924, new_U5925, new_U5926, new_U5927, new_U5928, new_U5929,
    new_U5930, new_U5931, new_U5932, new_U5933, new_U5934, new_U5935,
    new_U5936, new_U5937, new_U5938, new_U5939, new_U5940, new_U5941,
    new_U5942, new_U5943, new_U5944, new_U5945, new_U5946, new_U5947,
    new_U5948, new_U5949, new_U5950, new_U5951, new_U5952, new_U5953,
    new_U5954, new_U5955, new_U5956, new_U5957, new_U5958, new_U5959,
    new_U5960, new_U5961, new_U5962, new_U5963, new_U5964, new_U5965,
    new_U5966, new_U5967, new_U5968, new_U5969, new_U5970, new_U5971,
    new_U5972, new_U5973, new_U5974, new_U5975, new_U5976, new_U5977,
    new_U5978, new_U5979, new_U5980, new_U5981, new_U5982, new_U5983,
    new_U5984, new_U5985, new_U5986, new_U5987, new_U5988, new_U5989,
    new_U5990, new_U5991, new_U5992, new_U5993, new_U5994, new_U5995,
    new_U5996, new_U5997, new_U5998, new_U5999, new_U6000, new_U6001,
    new_U6002, new_U6003, new_U6004, new_U6005, new_U6006, new_U6007,
    new_U6008, new_U6009, new_U6010, new_U6011, new_U6012, new_U6013,
    new_U6014, new_U6015, new_U6016, new_U6017, new_U6018, new_U6019,
    new_U6020, new_U6021, new_U6022, new_U6023, new_U6024, new_U6025,
    new_U6026, new_U6027, new_U6028, new_U6029, new_U6030, new_U6031,
    new_U6032, new_U6033, new_U6034, new_U6035, new_U6036, new_U6037,
    new_U6038, new_U6039, new_U6040, new_U6041, new_U6042, new_U6043,
    new_U6044, new_U6045, new_U6046, new_U6047, new_U6048, new_U6049,
    new_U6050, new_U6051, new_U6052, new_U6053, new_U6054, new_U6055,
    new_U6056, new_U6057, new_U6058, new_U6059, new_U6060, new_U6061,
    new_U6062, new_U6063, new_U6064, new_U6065, new_U6066, new_U6067,
    new_U6068, new_U6069, new_U6070, new_U6071, new_U6072, new_U6073,
    new_U6074, new_U6075, new_U6076, new_U6077, new_U6078, new_U6079,
    new_U6080, new_U6081, new_U6082, new_U6083, new_U6084, new_U6085,
    new_U6086, new_U6087, new_U6088, new_U6089, new_U6090, new_U6091,
    new_U6092, new_U6093, new_U6094, new_U6095, new_U6096, new_U6097,
    new_U6098, new_U6099, new_U6100, new_U6101, new_U6102, new_U6103,
    new_U6104, new_U6105, new_U6106, new_U6107, new_U6108, new_U6109,
    new_U6110, new_U6111, new_U6112, new_U6113, new_U6114, new_U6115,
    new_U6116, new_U6117, new_U6118, new_U6119, new_U6120, new_U6121,
    new_U6122, new_U6123, new_U6124, new_U6125, new_U6126, new_U6127,
    new_U6128, new_U6129, new_U6130, new_U6131, new_U6132, new_U6133,
    new_U6134, new_U6135, new_U6136, new_U6137, new_U6138, new_U6139,
    new_U6140, new_U6141, new_U6142, new_U6143, new_U6144, new_U6145,
    new_U6146, new_U6147, new_U6148, new_U6149, new_U6150, new_U6151,
    new_U6152, new_U6153, new_U6154, new_U6155, new_U6156, new_U6157,
    new_U6158, new_U6159, new_U6160, new_U6161, new_U6162, new_U6163,
    new_U6164, new_U6165, new_U6166, new_U6167, new_U6168, new_U6169,
    new_U6170, new_U6171, new_U6172, new_U6173, new_U6174, new_U6175,
    new_U6176, new_U6177, new_U6178, new_U6179, new_U6180, new_U6181,
    new_U6182, new_U6183, new_U6184, new_U6185, new_U6186, new_U6187,
    new_U6188, new_U6189, new_U6190, new_U6191, new_U6192, new_U6193,
    new_U6194, new_U6195, new_U6196, new_U6197, new_U6198, new_U6199,
    new_U6200, new_U6201, new_U6202, new_U6203, new_U6204, new_U6205,
    new_U6206, new_U6207, new_U6208, new_U6209, new_U6210, new_U6211,
    new_U6212, new_U6213, new_U6214, new_U6215, new_U6216, new_U6217,
    new_U6218, new_U6219, new_U6220, new_U6221, new_U6222, new_U6223,
    new_U6224, new_U6225, new_U6226, new_U6227, new_U6228, new_U6229,
    new_U6230, new_U6231, new_U6232, new_U6233, new_U6234, new_U6235,
    new_U6236, new_U6237, new_U6238, new_U6239, new_U6240, new_U6241,
    new_U6242, new_U6243, new_U6244, new_U6245, new_U6246, new_U6247,
    new_U6248, new_U6249, new_U6250, new_U6251, new_U6252, new_U6253,
    new_U6254, new_U6255, new_U6256, new_U6257, new_U6258, new_U6259,
    new_U6260, new_U6261, new_U6262, new_U6263, new_U6264, new_U6265,
    new_U6266, new_U6267, new_U6268, new_U6269, new_U6270, new_U6271,
    new_U6272, new_U6273, new_U6274, new_U6275, new_U6276, new_U6277,
    new_U6278, new_U6279, new_U6280, new_U6281, new_U6282, new_U6283,
    new_U6284, new_U6285, new_U6286, new_U6287, new_U6288, new_U6289,
    new_U6290, new_U6291, new_U6292, new_U6293, new_U6294, new_U6295,
    new_U6296, new_U6297, new_U6298, new_U6299, new_U6300, new_U6301,
    new_U6302, new_U6303, new_U6304, new_U6305, new_U6306, new_U6307,
    new_U6308, new_U6309, new_U6310, new_U6311, new_U6312, new_U6313,
    new_U6314, new_U6315, new_U6316, new_U6317, new_U6318, new_U6319,
    new_U6320, new_U6321, new_U6322, new_U6323, new_R1222_U516,
    new_R1222_U515, new_R1222_U514, new_R1222_U513, new_R1222_U512,
    new_R1222_U511, new_R1222_U510, new_R1222_U509, new_R1222_U508,
    new_R1222_U507, new_R1222_U506, new_R1222_U505, new_R1222_U504,
    new_R1222_U503, new_R1222_U502, new_R1222_U501, new_R1222_U500,
    new_R1222_U499, new_R1222_U498, new_R1222_U497, new_R1222_U496,
    new_R1222_U495, new_SUB_84_U4, new_SUB_84_U5, new_SUB_84_U6,
    new_SUB_84_U7, new_SUB_84_U8, new_SUB_84_U9, new_SUB_84_U10,
    new_SUB_84_U11, new_SUB_84_U12, new_SUB_84_U13, new_SUB_84_U14,
    new_SUB_84_U15, new_SUB_84_U16, new_SUB_84_U17, new_SUB_84_U18,
    new_SUB_84_U19, new_SUB_84_U20, new_SUB_84_U21, new_SUB_84_U22,
    new_SUB_84_U23, new_SUB_84_U24, new_SUB_84_U25, new_SUB_84_U26,
    new_SUB_84_U27, new_SUB_84_U28, new_SUB_84_U29, new_SUB_84_U30,
    new_SUB_84_U31, new_SUB_84_U32, new_SUB_84_U33, new_SUB_84_U34,
    new_SUB_84_U35, new_SUB_84_U36, new_SUB_84_U37, new_SUB_84_U38,
    new_SUB_84_U39, new_SUB_84_U40, new_SUB_84_U41, new_SUB_84_U42,
    new_SUB_84_U43, new_SUB_84_U44, new_SUB_84_U45, new_SUB_84_U46,
    new_SUB_84_U47, new_SUB_84_U48, new_SUB_84_U49, new_SUB_84_U50,
    new_SUB_84_U51, new_SUB_84_U52, new_SUB_84_U53, new_SUB_84_U54,
    new_SUB_84_U55, new_SUB_84_U56, new_SUB_84_U57, new_SUB_84_U58,
    new_SUB_84_U59, new_SUB_84_U60, new_SUB_84_U61, new_SUB_84_U62,
    new_SUB_84_U63, new_SUB_84_U64, new_SUB_84_U65, new_SUB_84_U66,
    new_SUB_84_U67, new_SUB_84_U68, new_SUB_84_U69, new_SUB_84_U70,
    new_SUB_84_U71, new_SUB_84_U72, new_SUB_84_U73, new_SUB_84_U74,
    new_SUB_84_U75, new_SUB_84_U76, new_SUB_84_U77, new_SUB_84_U78,
    new_SUB_84_U79, new_SUB_84_U80, new_SUB_84_U81, new_SUB_84_U82,
    new_SUB_84_U83, new_SUB_84_U84, new_SUB_84_U85, new_SUB_84_U86,
    new_SUB_84_U87, new_SUB_84_U88, new_SUB_84_U89, new_SUB_84_U90,
    new_SUB_84_U91, new_SUB_84_U92, new_SUB_84_U93, new_SUB_84_U94,
    new_SUB_84_U95, new_SUB_84_U96, new_SUB_84_U97, new_SUB_84_U98,
    new_SUB_84_U99, new_SUB_84_U100, new_SUB_84_U101, new_SUB_84_U102,
    new_SUB_84_U103, new_SUB_84_U104, new_SUB_84_U105, new_SUB_84_U106,
    new_SUB_84_U107, new_SUB_84_U108, new_SUB_84_U109, new_SUB_84_U110,
    new_SUB_84_U111, new_SUB_84_U112, new_SUB_84_U113, new_SUB_84_U114,
    new_SUB_84_U115, new_SUB_84_U116, new_SUB_84_U117, new_SUB_84_U118,
    new_SUB_84_U119, new_SUB_84_U120, new_SUB_84_U121, new_SUB_84_U122,
    new_SUB_84_U123, new_SUB_84_U124, new_SUB_84_U125, new_SUB_84_U126,
    new_SUB_84_U127, new_SUB_84_U128, new_SUB_84_U129, new_SUB_84_U130,
    new_SUB_84_U131, new_SUB_84_U132, new_SUB_84_U133, new_SUB_84_U134,
    new_SUB_84_U135, new_SUB_84_U136, new_SUB_84_U137, new_SUB_84_U138,
    new_SUB_84_U139, new_SUB_84_U140, new_SUB_84_U141, new_SUB_84_U142,
    new_SUB_84_U143, new_SUB_84_U144, new_SUB_84_U145, new_SUB_84_U146,
    new_SUB_84_U147, new_SUB_84_U148, new_SUB_84_U149, new_SUB_84_U150,
    new_SUB_84_U151, new_SUB_84_U152, new_SUB_84_U153, new_SUB_84_U154,
    new_SUB_84_U155, new_SUB_84_U156, new_SUB_84_U157, new_SUB_84_U158,
    new_SUB_84_U159, new_SUB_84_U160, new_SUB_84_U161, new_ADD_95_U4,
    new_ADD_95_U5, new_ADD_95_U6, new_ADD_95_U7, new_ADD_95_U8,
    new_ADD_95_U9, new_ADD_95_U10, new_ADD_95_U11, new_ADD_95_U12,
    new_ADD_95_U13, new_ADD_95_U14, new_ADD_95_U15, new_ADD_95_U16,
    new_ADD_95_U17, new_ADD_95_U18, new_ADD_95_U19, new_ADD_95_U20,
    new_ADD_95_U21, new_ADD_95_U22, new_ADD_95_U23, new_ADD_95_U24,
    new_ADD_95_U25, new_ADD_95_U26, new_ADD_95_U27, new_ADD_95_U28,
    new_ADD_95_U29, new_ADD_95_U30, new_ADD_95_U31, new_ADD_95_U32,
    new_ADD_95_U33, new_ADD_95_U34, new_ADD_95_U35, new_ADD_95_U36,
    new_ADD_95_U37, new_ADD_95_U38, new_ADD_95_U39, new_ADD_95_U40,
    new_ADD_95_U41, new_ADD_95_U42, new_ADD_95_U43, new_ADD_95_U44,
    new_ADD_95_U45, new_ADD_95_U46, new_ADD_95_U47, new_ADD_95_U48,
    new_ADD_95_U49, new_ADD_95_U50, new_ADD_95_U51, new_ADD_95_U52,
    new_ADD_95_U53, new_ADD_95_U54, new_ADD_95_U55, new_ADD_95_U56,
    new_ADD_95_U57, new_ADD_95_U58, new_ADD_95_U59, new_ADD_95_U60,
    new_ADD_95_U61, new_ADD_95_U62, new_ADD_95_U63, new_ADD_95_U64,
    new_ADD_95_U65, new_ADD_95_U66, new_ADD_95_U67, new_ADD_95_U68,
    new_ADD_95_U69, new_ADD_95_U70, new_ADD_95_U71, new_ADD_95_U72,
    new_ADD_95_U73, new_ADD_95_U74, new_ADD_95_U75, new_ADD_95_U76,
    new_ADD_95_U77, new_ADD_95_U78, new_ADD_95_U79, new_ADD_95_U80,
    new_ADD_95_U81, new_ADD_95_U82, new_ADD_95_U83, new_ADD_95_U84,
    new_ADD_95_U85, new_ADD_95_U86, new_ADD_95_U87, new_ADD_95_U88,
    new_ADD_95_U89, new_ADD_95_U90, new_ADD_95_U91, new_ADD_95_U92,
    new_ADD_95_U93, new_ADD_95_U94, new_ADD_95_U95, new_ADD_95_U96,
    new_ADD_95_U97, new_ADD_95_U98, new_ADD_95_U99, new_ADD_95_U100,
    new_ADD_95_U101, new_ADD_95_U102, new_ADD_95_U103, new_ADD_95_U104,
    new_ADD_95_U105, new_ADD_95_U106, new_ADD_95_U107, new_ADD_95_U108,
    new_ADD_95_U109, new_ADD_95_U110, new_ADD_95_U111, new_ADD_95_U112,
    new_ADD_95_U113, new_ADD_95_U114, new_ADD_95_U115, new_ADD_95_U116,
    new_ADD_95_U117, new_ADD_95_U118, new_ADD_95_U119, new_ADD_95_U120,
    new_ADD_95_U121, new_ADD_95_U122, new_ADD_95_U123, new_ADD_95_U124,
    new_ADD_95_U125, new_ADD_95_U126, new_ADD_95_U127, new_ADD_95_U128,
    new_ADD_95_U129, new_ADD_95_U130, new_ADD_95_U131, new_ADD_95_U132,
    new_ADD_95_U133, new_ADD_95_U134, new_ADD_95_U135, new_ADD_95_U136,
    new_ADD_95_U137, new_ADD_95_U138, new_ADD_95_U139, new_ADD_95_U140,
    new_ADD_95_U141, new_ADD_95_U142, new_ADD_95_U143, new_ADD_95_U144,
    new_ADD_95_U145, new_ADD_95_U146, new_ADD_95_U147, new_ADD_95_U148,
    new_ADD_95_U149, new_ADD_95_U150, new_ADD_95_U151, new_ADD_95_U152,
    new_ADD_95_U153, new_ADD_95_U154, new_ADD_95_U155, new_ADD_95_U156,
    new_ADD_95_U157, new_ADD_95_U158, new_ADD_95_U159, new_R395_U6,
    new_R395_U7, new_R395_U8, new_R395_U9, new_R395_U10, new_R395_U11,
    new_R395_U12, new_R395_U13, new_R395_U14, new_R395_U15, new_R395_U16,
    new_R395_U17, new_R395_U18, new_R395_U19, new_R395_U20, new_R395_U21,
    new_R395_U22, new_R395_U23, new_R395_U24, new_R395_U25, new_R395_U26,
    new_R395_U27, new_R395_U28, new_R395_U29, new_R395_U30, new_R395_U31,
    new_R395_U32, new_R395_U33, new_R395_U34, new_R395_U35, new_R395_U36,
    new_R395_U37, new_R395_U38, new_R395_U39, new_R395_U40, new_R395_U41,
    new_R395_U42, new_R395_U43, new_R395_U44, new_R395_U45, new_R395_U46,
    new_R395_U47, new_R395_U48, new_R395_U49, new_R395_U50, new_R395_U51,
    new_R395_U52, new_R395_U53, new_R395_U54, new_R395_U55, new_R395_U56,
    new_R395_U57, new_R395_U58, new_R395_U59, new_R395_U60, new_R395_U61,
    new_R395_U62, new_R395_U63, new_R395_U64, new_R395_U65, new_R395_U66,
    new_R395_U67, new_R395_U68, new_R395_U69, new_R395_U70, new_R395_U71,
    new_R395_U72, new_R395_U73, new_R395_U74, new_R395_U75, new_R395_U76,
    new_R395_U77, new_R395_U78, new_R395_U79, new_R395_U80, new_R395_U81,
    new_R395_U82, new_R395_U83, new_R395_U84, new_R395_U85, new_R395_U86,
    new_R395_U87, new_R395_U88, new_R395_U89, new_R395_U90, new_R395_U91,
    new_R395_U92, new_R395_U93, new_R395_U94, new_R395_U95, new_R395_U96,
    new_R395_U97, new_R395_U98, new_R395_U99, new_R395_U100, new_R395_U101,
    new_R395_U102, new_R395_U103, new_R395_U104, new_R395_U105,
    new_R395_U106, new_R395_U107, new_R395_U108, new_R395_U109,
    new_R395_U110, new_R395_U111, new_R395_U112, new_R395_U113,
    new_R395_U114, new_R395_U115, new_R395_U116, new_R395_U117,
    new_R395_U118, new_R395_U119, new_R395_U120, new_R395_U121,
    new_R395_U122, new_R395_U123, new_R395_U124, new_R395_U125,
    new_R395_U126, new_R395_U127, new_R395_U128, new_R395_U129,
    new_R395_U130, new_R395_U131, new_R395_U132, new_R395_U133,
    new_R395_U134, new_R395_U135, new_R395_U136, new_R395_U137,
    new_R395_U138, new_R395_U139, new_R395_U140, new_R395_U141,
    new_R395_U142, new_R395_U143, new_R395_U144, new_R395_U145,
    new_R395_U146, new_R395_U147, new_R395_U148, new_R395_U149,
    new_R395_U150, new_R395_U151, new_R395_U152, new_R395_U153,
    new_R395_U154, new_R395_U155, new_R395_U156, new_R395_U157,
    new_R395_U158, new_R395_U159, new_R395_U160, new_R395_U161,
    new_R395_U162, new_R395_U163, new_R395_U164, new_R395_U165,
    new_R395_U166, new_R395_U167, new_R395_U168, new_R395_U169,
    new_R395_U170, new_R395_U171, new_R395_U172, new_R395_U173,
    new_R395_U174, new_R395_U175, new_R395_U176, new_R395_U177,
    new_R395_U178, new_R395_U179, new_R395_U180, new_R395_U181,
    new_R395_U182, new_R395_U183, new_R395_U184, new_R395_U185,
    new_R395_U186, new_R395_U187, new_R395_U188, new_R1105_U4,
    new_R1105_U5, new_R1105_U6, new_R1105_U7, new_R1105_U8, new_R1105_U9,
    new_R1105_U10, new_R1105_U11, new_R1105_U12, new_R1105_U13,
    new_R1105_U14, new_R1105_U15, new_R1105_U16, new_R1105_U17,
    new_R1105_U18, new_R1105_U19, new_R1105_U20, new_R1105_U21,
    new_R1105_U22, new_R1105_U23, new_R1105_U24, new_R1105_U25,
    new_R1105_U26, new_R1105_U27, new_R1105_U28, new_R1105_U29,
    new_R1105_U30, new_R1105_U31, new_R1105_U32, new_R1105_U33,
    new_R1105_U34, new_R1105_U35, new_R1105_U36, new_R1105_U37,
    new_R1105_U38, new_R1105_U39, new_R1105_U40, new_R1105_U41,
    new_R1105_U42, new_R1105_U43, new_R1105_U44, new_R1105_U45,
    new_R1105_U46, new_R1105_U47, new_R1105_U48, new_R1105_U49,
    new_R1105_U50, new_R1105_U51, new_R1105_U52, new_R1105_U53,
    new_R1105_U54, new_R1105_U55, new_R1105_U56, new_R1105_U57,
    new_R1105_U58, new_R1105_U59, new_R1105_U60, new_R1105_U61,
    new_R1105_U62, new_R1105_U63, new_R1105_U64, new_R1105_U65,
    new_R1105_U66, new_R1105_U67, new_R1105_U68, new_R1105_U69,
    new_R1105_U70, new_R1105_U71, new_R1105_U72, new_R1105_U73,
    new_R1105_U74, new_R1105_U75, new_R1105_U76, new_R1105_U77,
    new_R1105_U78, new_R1105_U79, new_R1105_U80, new_R1105_U81,
    new_R1105_U82, new_R1105_U83, new_R1105_U84, new_R1105_U85,
    new_R1105_U86, new_R1105_U87, new_R1105_U88, new_R1105_U89,
    new_R1105_U90, new_R1105_U91, new_R1105_U92, new_R1105_U93,
    new_R1105_U94, new_R1105_U95, new_R1105_U96, new_R1105_U97,
    new_R1105_U98, new_R1105_U99, new_R1105_U100, new_R1105_U101,
    new_R1105_U102, new_R1105_U103, new_R1105_U104, new_R1105_U105,
    new_R1105_U106, new_R1105_U107, new_R1105_U108, new_R1105_U109,
    new_R1105_U110, new_R1105_U111, new_R1105_U112, new_R1105_U113,
    new_R1105_U114, new_R1105_U115, new_R1105_U116, new_R1105_U117,
    new_R1105_U118, new_R1105_U119, new_R1105_U120, new_R1105_U121,
    new_R1105_U122, new_R1105_U123, new_R1105_U124, new_R1105_U125,
    new_R1105_U126, new_R1105_U127, new_R1105_U128, new_R1105_U129,
    new_R1105_U130, new_R1105_U131, new_R1105_U132, new_R1105_U133,
    new_R1105_U134, new_R1105_U135, new_R1105_U136, new_R1105_U137,
    new_R1105_U138, new_R1105_U139, new_R1105_U140, new_R1105_U141,
    new_R1105_U142, new_R1105_U143, new_R1105_U144, new_R1105_U145,
    new_R1105_U146, new_R1105_U147, new_R1105_U148, new_R1105_U149,
    new_R1105_U150, new_R1105_U151, new_R1105_U152, new_R1105_U153,
    new_R1105_U154, new_R1105_U155, new_R1105_U156, new_R1105_U157,
    new_R1105_U158, new_R1105_U159, new_R1105_U160, new_R1105_U161,
    new_R1105_U162, new_R1105_U163, new_R1105_U164, new_R1105_U165,
    new_R1105_U166, new_R1105_U167, new_R1105_U168, new_R1105_U169,
    new_R1105_U170, new_R1105_U171, new_R1105_U172, new_R1105_U173,
    new_R1105_U174, new_R1105_U175, new_R1105_U176, new_R1105_U177,
    new_R1105_U178, new_R1105_U179, new_R1105_U180, new_R1105_U181,
    new_R1105_U182, new_R1105_U183, new_R1105_U184, new_R1105_U185,
    new_R1105_U186, new_R1105_U187, new_R1105_U188, new_R1105_U189,
    new_R1105_U190, new_R1105_U191, new_R1105_U192, new_R1105_U193,
    new_R1105_U194, new_R1105_U195, new_R1105_U196, new_R1105_U197,
    new_R1105_U198, new_R1105_U199, new_R1105_U200, new_R1105_U201,
    new_R1105_U202, new_R1105_U203, new_R1105_U204, new_R1105_U205,
    new_R1105_U206, new_R1105_U207, new_R1105_U208, new_R1105_U209,
    new_R1105_U210, new_R1105_U211, new_R1105_U212, new_R1105_U213,
    new_R1105_U214, new_R1105_U215, new_R1105_U216, new_R1105_U217,
    new_R1105_U218, new_R1105_U219, new_R1105_U220, new_R1105_U221,
    new_R1105_U222, new_R1105_U223, new_R1105_U224, new_R1105_U225,
    new_R1105_U226, new_R1105_U227, new_R1105_U228, new_R1105_U229,
    new_R1105_U230, new_R1105_U231, new_R1105_U232, new_R1105_U233,
    new_R1105_U234, new_R1105_U235, new_R1105_U236, new_R1105_U237,
    new_R1105_U238, new_R1105_U239, new_R1105_U240, new_R1105_U241,
    new_R1105_U242, new_R1105_U243, new_R1105_U244, new_R1105_U245,
    new_R1105_U246, new_R1105_U247, new_R1105_U248, new_R1105_U249,
    new_R1105_U250, new_R1105_U251, new_R1105_U252, new_R1105_U253,
    new_R1105_U254, new_R1105_U255, new_R1105_U256, new_R1105_U257,
    new_R1105_U258, new_R1105_U259, new_R1105_U260, new_R1105_U261,
    new_R1105_U262, new_R1105_U263, new_R1105_U264, new_R1105_U265,
    new_R1105_U266, new_R1105_U267, new_R1105_U268, new_R1105_U269,
    new_R1105_U270, new_R1105_U271, new_R1105_U272, new_R1105_U273,
    new_R1105_U274, new_R1105_U275, new_R1105_U276, new_R1105_U277,
    new_R1105_U278, new_R1105_U279, new_R1105_U280, new_R1105_U281,
    new_R1105_U282, new_R1105_U283, new_R1105_U284, new_R1105_U285,
    new_R1105_U286, new_R1105_U287, new_R1105_U288, new_R1105_U289,
    new_R1105_U290, new_R1105_U291, new_R1105_U292, new_R1105_U293,
    new_R1105_U294, new_R1105_U295, new_R1105_U296, new_R1105_U297,
    new_R1105_U298, new_R1105_U299, new_R1105_U300, new_R1105_U301,
    new_R1105_U302, new_R1105_U303, new_R1105_U304, new_R1105_U305,
    new_R1105_U306, new_R1105_U307, new_R1105_U308, new_R1105_U309,
    new_R1105_U310, new_R1105_U311, new_R1309_U6, new_R1309_U7,
    new_R1309_U8, new_R1309_U9, new_R1309_U10, new_R1282_U6, new_R1282_U7,
    new_R1282_U8, new_R1282_U9, new_R1282_U10, new_R1282_U11,
    new_R1282_U12, new_R1282_U13, new_R1282_U14, new_R1282_U15,
    new_R1282_U16, new_R1282_U17, new_R1282_U18, new_R1282_U19,
    new_R1282_U20, new_R1282_U21, new_R1282_U22, new_R1282_U23,
    new_R1282_U24, new_R1282_U25, new_R1282_U26, new_R1282_U27,
    new_R1282_U28, new_R1282_U29, new_R1282_U30, new_R1282_U31,
    new_R1282_U32, new_R1282_U33, new_R1282_U34, new_R1282_U35,
    new_R1282_U36, new_R1282_U37, new_R1282_U38, new_R1282_U39,
    new_R1282_U40, new_R1282_U41, new_R1282_U42, new_R1282_U43,
    new_R1282_U44, new_R1282_U45, new_R1282_U46, new_R1282_U47,
    new_R1282_U48, new_R1282_U49, new_R1282_U50, new_R1282_U51,
    new_R1282_U52, new_R1282_U53, new_R1282_U54, new_R1282_U55,
    new_R1282_U56, new_R1282_U57, new_R1282_U58, new_R1282_U59,
    new_R1282_U60, new_R1282_U61, new_R1282_U62, new_R1282_U63,
    new_R1282_U64, new_R1282_U65, new_R1282_U66, new_R1282_U67,
    new_R1282_U68, new_R1282_U69, new_R1282_U70, new_R1282_U71,
    new_R1282_U72, new_R1282_U73, new_R1282_U74, new_R1282_U75,
    new_R1282_U76, new_R1282_U77, new_R1282_U78, new_R1282_U79,
    new_R1282_U80, new_R1282_U81, new_R1282_U82, new_R1282_U83,
    new_R1282_U84, new_R1282_U85, new_R1282_U86, new_R1282_U87,
    new_R1282_U88, new_R1282_U89, new_R1282_U90, new_R1282_U91,
    new_R1282_U92, new_R1282_U93, new_R1282_U94, new_R1282_U95,
    new_R1282_U96, new_R1282_U97, new_R1282_U98, new_R1282_U99,
    new_R1282_U100, new_R1282_U101, new_R1282_U102, new_R1282_U103,
    new_R1282_U104, new_R1282_U105, new_R1282_U106, new_R1282_U107,
    new_R1282_U108, new_R1282_U109, new_R1282_U110, new_R1282_U111,
    new_R1282_U112, new_R1282_U113, new_R1282_U114, new_R1282_U115,
    new_R1282_U116, new_R1282_U117, new_R1282_U118, new_R1282_U119,
    new_R1282_U120, new_R1282_U121, new_R1282_U122, new_R1282_U123,
    new_R1282_U124, new_R1282_U125, new_R1282_U126, new_R1282_U127,
    new_R1282_U128, new_R1282_U129, new_R1282_U130, new_R1282_U131,
    new_R1282_U132, new_R1282_U133, new_R1282_U134, new_R1282_U135,
    new_R1282_U136, new_R1282_U137, new_R1282_U138, new_R1282_U139,
    new_R1282_U140, new_R1282_U141, new_R1282_U142, new_R1282_U143,
    new_R1282_U144, new_R1282_U145, new_R1282_U146, new_R1282_U147,
    new_R1282_U148, new_R1282_U149, new_R1282_U150, new_R1282_U151,
    new_R1282_U152, new_R1282_U153, new_R1282_U154, new_R1282_U155,
    new_R1282_U156, new_R1282_U157, new_R1282_U158, new_R1282_U159,
    new_R1282_U160, new_R1282_U161, new_R1282_U162, new_R1282_U163,
    new_R1282_U164, new_R1282_U165, new_R1282_U166, new_R1282_U167,
    new_R1282_U168, new_R1282_U169, new_R1282_U170, new_R1282_U171,
    new_R1282_U172, new_R1282_U173, new_R1282_U174, new_R1282_U175,
    new_R1282_U176, new_R1282_U177, new_R1282_U178, new_R1282_U179,
    new_R1282_U180, new_R1240_U4, new_R1240_U5, new_R1240_U6, new_R1240_U7,
    new_R1240_U8, new_R1240_U9, new_R1240_U10, new_R1240_U11,
    new_R1240_U12, new_R1240_U13, new_R1240_U14, new_R1240_U15,
    new_R1240_U16, new_R1240_U17, new_R1240_U18, new_R1240_U19,
    new_R1240_U20, new_R1240_U21, new_R1240_U22, new_R1240_U23,
    new_R1240_U24, new_R1240_U25, new_R1240_U26, new_R1240_U27,
    new_R1240_U28, new_R1240_U29, new_R1240_U30, new_R1240_U31,
    new_R1240_U32, new_R1240_U33, new_R1240_U34, new_R1240_U35,
    new_R1240_U36, new_R1240_U37, new_R1240_U38, new_R1240_U39,
    new_R1240_U40, new_R1240_U41, new_R1240_U42, new_R1240_U43,
    new_R1240_U44, new_R1240_U45, new_R1240_U46, new_R1240_U47,
    new_R1240_U48, new_R1240_U49, new_R1240_U50, new_R1240_U51,
    new_R1240_U52, new_R1240_U53, new_R1240_U54, new_R1240_U55,
    new_R1240_U56, new_R1240_U57, new_R1240_U58, new_R1240_U59,
    new_R1240_U60, new_R1240_U61, new_R1240_U62, new_R1240_U63,
    new_R1240_U64, new_R1240_U65, new_R1240_U66, new_R1240_U67,
    new_R1240_U68, new_R1240_U69, new_R1240_U70, new_R1240_U71,
    new_R1240_U72, new_R1240_U73, new_R1240_U74, new_R1240_U75,
    new_R1240_U76, new_R1240_U77, new_R1240_U78, new_R1240_U79,
    new_R1240_U80, new_R1240_U81, new_R1240_U82, new_R1240_U83,
    new_R1240_U84, new_R1240_U85, new_R1240_U86, new_R1240_U87,
    new_R1240_U88, new_R1240_U89, new_R1240_U90, new_R1240_U91,
    new_R1240_U92, new_R1240_U93, new_R1240_U94, new_R1240_U95,
    new_R1240_U96, new_R1240_U97, new_R1240_U98, new_R1240_U99,
    new_R1240_U100, new_R1240_U101, new_R1240_U102, new_R1240_U103,
    new_R1240_U104, new_R1240_U105, new_R1240_U106, new_R1240_U107,
    new_R1240_U108, new_R1240_U109, new_R1240_U110, new_R1240_U111,
    new_R1240_U112, new_R1240_U113, new_R1240_U114, new_R1240_U115,
    new_R1240_U116, new_R1240_U117, new_R1240_U118, new_R1240_U119,
    new_R1240_U120, new_R1240_U121, new_R1240_U122, new_R1240_U123,
    new_R1240_U124, new_R1240_U125, new_R1240_U126, new_R1240_U127,
    new_R1240_U128, new_R1240_U129, new_R1240_U130, new_R1240_U131,
    new_R1240_U132, new_R1240_U133, new_R1240_U134, new_R1240_U135,
    new_R1240_U136, new_R1240_U137, new_R1240_U138, new_R1240_U139,
    new_R1240_U140, new_R1240_U141, new_R1240_U142, new_R1240_U143,
    new_R1240_U144, new_R1240_U145, new_R1240_U146, new_R1240_U147,
    new_R1240_U148, new_R1240_U149, new_R1240_U150, new_R1240_U151,
    new_R1240_U152, new_R1240_U153, new_R1240_U154, new_R1240_U155,
    new_R1240_U156, new_R1240_U157, new_R1240_U158, new_R1240_U159,
    new_R1240_U160, new_R1240_U161, new_R1240_U162, new_R1240_U163,
    new_R1240_U164, new_R1240_U165, new_R1240_U166, new_R1240_U167,
    new_R1240_U168, new_R1240_U169, new_R1240_U170, new_R1240_U171,
    new_R1240_U172, new_R1240_U173, new_R1240_U174, new_R1240_U175,
    new_R1240_U176, new_R1240_U177, new_R1240_U178, new_R1240_U179,
    new_R1240_U180, new_R1240_U181, new_R1240_U182, new_R1240_U183,
    new_R1240_U184, new_R1240_U185, new_R1240_U186, new_R1240_U187,
    new_R1240_U188, new_R1240_U189, new_R1240_U190, new_R1240_U191,
    new_R1240_U192, new_R1240_U193, new_R1240_U194, new_R1240_U195,
    new_R1240_U196, new_R1240_U197, new_R1240_U198, new_R1240_U199,
    new_R1240_U200, new_R1240_U201, new_R1240_U202, new_R1240_U203,
    new_R1240_U204, new_R1240_U205, new_R1240_U206, new_R1240_U207,
    new_R1240_U208, new_R1240_U209, new_R1240_U210, new_R1240_U211,
    new_R1240_U212, new_R1240_U213, new_R1240_U214, new_R1240_U215,
    new_R1240_U216, new_R1240_U217, new_R1240_U218, new_R1240_U219,
    new_R1240_U220, new_R1240_U221, new_R1240_U222, new_R1240_U223,
    new_R1240_U224, new_R1240_U225, new_R1240_U226, new_R1240_U227,
    new_R1240_U228, new_R1240_U229, new_R1240_U230, new_R1240_U231,
    new_R1240_U232, new_R1240_U233, new_R1240_U234, new_R1240_U235,
    new_R1240_U236, new_R1240_U237, new_R1240_U238, new_R1240_U239,
    new_R1240_U240, new_R1240_U241, new_R1240_U242, new_R1240_U243,
    new_R1240_U244, new_R1240_U245, new_R1240_U246, new_R1240_U247,
    new_R1240_U248, new_R1240_U249, new_R1240_U250, new_R1240_U251,
    new_R1240_U252, new_R1240_U253, new_R1240_U254, new_R1240_U255,
    new_R1240_U256, new_R1240_U257, new_R1240_U258, new_R1240_U259,
    new_R1240_U260, new_R1240_U261, new_R1240_U262, new_R1240_U263,
    new_R1240_U264, new_R1240_U265, new_R1240_U266, new_R1240_U267,
    new_R1240_U268, new_R1240_U269, new_R1240_U270, new_R1240_U271,
    new_R1240_U272, new_R1240_U273, new_R1240_U274, new_R1240_U275,
    new_R1240_U276, new_R1240_U277, new_R1240_U278, new_R1240_U279,
    new_R1240_U280, new_R1240_U281, new_R1240_U282, new_R1240_U283,
    new_R1240_U284, new_R1240_U285, new_R1240_U286, new_R1240_U287,
    new_R1240_U288, new_R1240_U289, new_R1240_U290, new_R1240_U291,
    new_R1240_U292, new_R1240_U293, new_R1240_U294, new_R1240_U295,
    new_R1240_U296, new_R1240_U297, new_R1240_U298, new_R1240_U299,
    new_R1240_U300, new_R1240_U301, new_R1240_U302, new_R1240_U303,
    new_R1240_U304, new_R1240_U305, new_R1240_U306, new_R1240_U307,
    new_R1240_U308, new_R1240_U309, new_R1240_U310, new_R1240_U311,
    new_R1240_U312, new_R1240_U313, new_R1240_U314, new_R1240_U315,
    new_R1240_U316, new_R1240_U317, new_R1240_U318, new_R1240_U319,
    new_R1240_U320, new_R1240_U321, new_R1240_U322, new_R1240_U323,
    new_R1240_U324, new_R1240_U325, new_R1240_U326, new_R1240_U327,
    new_R1240_U328, new_R1240_U329, new_R1240_U330, new_R1240_U331,
    new_R1240_U332, new_R1240_U333, new_R1240_U334, new_R1240_U335,
    new_R1240_U336, new_R1240_U337, new_R1240_U338, new_R1240_U339,
    new_R1240_U340, new_R1240_U341, new_R1240_U342, new_R1240_U343,
    new_R1240_U344, new_R1240_U345, new_R1240_U346, new_R1240_U347,
    new_R1240_U348, new_R1240_U349, new_R1240_U350, new_R1240_U351,
    new_R1240_U352, new_R1240_U353, new_R1240_U354, new_R1240_U355,
    new_R1240_U356, new_R1240_U357, new_R1240_U358, new_R1240_U359,
    new_R1240_U360, new_R1240_U361, new_R1240_U362, new_R1240_U363,
    new_R1240_U364, new_R1240_U365, new_R1240_U366, new_R1240_U367,
    new_R1240_U368, new_R1240_U369, new_R1240_U370, new_R1240_U371,
    new_R1240_U372, new_R1240_U373, new_R1240_U374, new_R1240_U375,
    new_R1240_U376, new_R1240_U377, new_R1240_U378, new_R1240_U379,
    new_R1240_U380, new_R1240_U381, new_R1240_U382, new_R1240_U383,
    new_R1240_U384, new_R1240_U385, new_R1240_U386, new_R1240_U387,
    new_R1240_U388, new_R1240_U389, new_R1240_U390, new_R1240_U391,
    new_R1240_U392, new_R1240_U393, new_R1240_U394, new_R1240_U395,
    new_R1240_U396, new_R1240_U397, new_R1240_U398, new_R1240_U399,
    new_R1240_U400, new_R1240_U401, new_R1240_U402, new_R1240_U403,
    new_R1240_U404, new_R1240_U405, new_R1240_U406, new_R1240_U407,
    new_R1240_U408, new_R1240_U409, new_R1240_U410, new_R1240_U411,
    new_R1240_U412, new_R1240_U413, new_R1240_U414, new_R1240_U415,
    new_R1240_U416, new_R1240_U417, new_R1240_U418, new_R1240_U419,
    new_R1240_U420, new_R1240_U421, new_R1240_U422, new_R1240_U423,
    new_R1240_U424, new_R1240_U425, new_R1240_U426, new_R1240_U427,
    new_R1240_U428, new_R1240_U429, new_R1240_U430, new_R1240_U431,
    new_R1240_U432, new_R1240_U433, new_R1240_U434, new_R1240_U435,
    new_R1240_U436, new_R1240_U437, new_R1240_U438, new_R1240_U439,
    new_R1240_U440, new_R1240_U441, new_R1240_U442, new_R1240_U443,
    new_R1240_U444, new_R1240_U445, new_R1240_U446, new_R1240_U447,
    new_R1240_U448, new_R1240_U449, new_R1240_U450, new_R1240_U451,
    new_R1240_U452, new_R1240_U453, new_R1240_U454, new_R1240_U455,
    new_R1240_U456, new_R1240_U457, new_R1240_U458, new_R1240_U459,
    new_R1240_U460, new_R1240_U461, new_R1240_U462, new_R1240_U463,
    new_R1240_U464, new_R1240_U465, new_R1240_U466, new_R1240_U467,
    new_R1240_U468, new_R1240_U469, new_R1240_U470, new_R1240_U471,
    new_R1240_U472, new_R1240_U473, new_R1240_U474, new_R1240_U475,
    new_R1240_U476, new_R1240_U477, new_R1240_U478, new_R1240_U479,
    new_R1240_U480, new_R1240_U481, new_R1240_U482, new_R1240_U483,
    new_R1240_U484, new_R1240_U485, new_R1240_U486, new_R1240_U487,
    new_R1240_U488, new_R1240_U489, new_R1240_U490, new_R1240_U491,
    new_R1240_U492, new_R1240_U493, new_R1240_U494, new_R1240_U495,
    new_R1240_U496, new_R1240_U497, new_R1240_U498, new_R1240_U499,
    new_R1240_U500, new_R1240_U501, new_R1240_U502, new_R1240_U503,
    new_R1240_U504, new_R1240_U505, new_R1240_U506, new_R1240_U507,
    new_R1240_U508, new_R1240_U509, new_R1240_U510, new_R1240_U511,
    new_R1240_U512, new_R1240_U513, new_R1240_U514, new_R1240_U515,
    new_R1240_U516, new_R1240_U517, new_R1240_U518, new_R1240_U519,
    new_R1240_U520, new_R1240_U521, new_R1240_U522, new_R1240_U523,
    new_R1240_U524, new_R1240_U525, new_R1240_U526, new_R1240_U527,
    new_R1240_U528, new_R1240_U529, new_R1240_U530, new_R1240_U531,
    new_R1162_U4, new_R1162_U5, new_R1162_U6, new_R1162_U7, new_R1162_U8,
    new_R1162_U9, new_R1162_U10, new_R1162_U11, new_R1162_U12,
    new_R1162_U13, new_R1162_U14, new_R1162_U15, new_R1162_U16,
    new_R1162_U17, new_R1162_U18, new_R1162_U19, new_R1162_U20,
    new_R1162_U21, new_R1162_U22, new_R1162_U23, new_R1162_U24,
    new_R1162_U25, new_R1162_U26, new_R1162_U27, new_R1162_U28,
    new_R1162_U29, new_R1162_U30, new_R1162_U31, new_R1162_U32,
    new_R1162_U33, new_R1162_U34, new_R1162_U35, new_R1162_U36,
    new_R1162_U37, new_R1162_U38, new_R1162_U39, new_R1162_U40,
    new_R1162_U41, new_R1162_U42, new_R1162_U43, new_R1162_U44,
    new_R1162_U45, new_R1162_U46, new_R1162_U47, new_R1162_U48,
    new_R1162_U49, new_R1162_U50, new_R1162_U51, new_R1162_U52,
    new_R1162_U53, new_R1162_U54, new_R1162_U55, new_R1162_U56,
    new_R1162_U57, new_R1162_U58, new_R1162_U59, new_R1162_U60,
    new_R1162_U61, new_R1162_U62, new_R1162_U63, new_R1162_U64,
    new_R1162_U65, new_R1162_U66, new_R1162_U67, new_R1162_U68,
    new_R1162_U69, new_R1162_U70, new_R1162_U71, new_R1162_U72,
    new_R1162_U73, new_R1162_U74, new_R1162_U75, new_R1162_U76,
    new_R1162_U77, new_R1162_U78, new_R1162_U79, new_R1162_U80,
    new_R1162_U81, new_R1162_U82, new_R1162_U83, new_R1162_U84,
    new_R1162_U85, new_R1162_U86, new_R1162_U87, new_R1162_U88,
    new_R1162_U89, new_R1162_U90, new_R1162_U91, new_R1162_U92,
    new_R1162_U93, new_R1162_U94, new_R1162_U95, new_R1162_U96,
    new_R1162_U97, new_R1162_U98, new_R1162_U99, new_R1162_U100,
    new_R1162_U101, new_R1162_U102, new_R1162_U103, new_R1162_U104,
    new_R1162_U105, new_R1162_U106, new_R1162_U107, new_R1162_U108,
    new_R1162_U109, new_R1162_U110, new_R1162_U111, new_R1162_U112,
    new_R1162_U113, new_R1162_U114, new_R1162_U115, new_R1162_U116,
    new_R1162_U117, new_R1162_U118, new_R1162_U119, new_R1162_U120,
    new_R1162_U121, new_R1162_U122, new_R1162_U123, new_R1162_U124,
    new_R1162_U125, new_R1162_U126, new_R1162_U127, new_R1162_U128,
    new_R1162_U129, new_R1162_U130, new_R1162_U131, new_R1162_U132,
    new_R1162_U133, new_R1162_U134, new_R1162_U135, new_R1162_U136,
    new_R1162_U137, new_R1162_U138, new_R1162_U139, new_R1162_U140,
    new_R1162_U141, new_R1162_U142, new_R1162_U143, new_R1162_U144,
    new_R1162_U145, new_R1162_U146, new_R1162_U147, new_R1162_U148,
    new_R1162_U149, new_R1162_U150, new_R1162_U151, new_R1162_U152,
    new_R1162_U153, new_R1162_U154, new_R1162_U155, new_R1162_U156,
    new_R1162_U157, new_R1162_U158, new_R1162_U159, new_R1162_U160,
    new_R1162_U161, new_R1162_U162, new_R1162_U163, new_R1162_U164,
    new_R1162_U165, new_R1162_U166, new_R1162_U167, new_R1162_U168,
    new_R1162_U169, new_R1162_U170, new_R1162_U171, new_R1162_U172,
    new_R1162_U173, new_R1162_U174, new_R1162_U175, new_R1162_U176,
    new_R1162_U177, new_R1162_U178, new_R1162_U179, new_R1162_U180,
    new_R1162_U181, new_R1162_U182, new_R1162_U183, new_R1162_U184,
    new_R1162_U185, new_R1162_U186, new_R1162_U187, new_R1162_U188,
    new_R1162_U189, new_R1162_U190, new_R1162_U191, new_R1162_U192,
    new_R1162_U193, new_R1162_U194, new_R1162_U195, new_R1162_U196,
    new_R1162_U197, new_R1162_U198, new_R1162_U199, new_R1162_U200,
    new_R1162_U201, new_R1162_U202, new_R1162_U203, new_R1162_U204,
    new_R1162_U205, new_R1162_U206, new_R1162_U207, new_R1162_U208,
    new_R1162_U209, new_R1162_U210, new_R1162_U211, new_R1162_U212,
    new_R1162_U213, new_R1162_U214, new_R1162_U215, new_R1162_U216,
    new_R1162_U217, new_R1162_U218, new_R1162_U219, new_R1162_U220,
    new_R1162_U221, new_R1162_U222, new_R1162_U223, new_R1162_U224,
    new_R1162_U225, new_R1162_U226, new_R1162_U227, new_R1162_U228,
    new_R1162_U229, new_R1162_U230, new_R1162_U231, new_R1162_U232,
    new_R1162_U233, new_R1162_U234, new_R1162_U235, new_R1162_U236,
    new_R1162_U237, new_R1162_U238, new_R1162_U239, new_R1162_U240,
    new_R1162_U241, new_R1162_U242, new_R1162_U243, new_R1162_U244,
    new_R1162_U245, new_R1162_U246, new_R1162_U247, new_R1162_U248,
    new_R1162_U249, new_R1162_U250, new_R1162_U251, new_R1162_U252,
    new_R1162_U253, new_R1162_U254, new_R1162_U255, new_R1162_U256,
    new_R1162_U257, new_R1162_U258, new_R1162_U259, new_R1162_U260,
    new_R1162_U261, new_R1162_U262, new_R1162_U263, new_R1162_U264,
    new_R1162_U265, new_R1162_U266, new_R1162_U267, new_R1162_U268,
    new_R1162_U269, new_R1162_U270, new_R1162_U271, new_R1162_U272,
    new_R1162_U273, new_R1162_U274, new_R1162_U275, new_R1162_U276,
    new_R1162_U277, new_R1162_U278, new_R1162_U279, new_R1162_U280,
    new_R1162_U281, new_R1162_U282, new_R1162_U283, new_R1162_U284,
    new_R1162_U285, new_R1162_U286, new_R1162_U287, new_R1162_U288,
    new_R1162_U289, new_R1162_U290, new_R1117_U6, new_R1117_U7,
    new_R1117_U8, new_R1117_U9, new_R1117_U10, new_R1117_U11,
    new_R1117_U12, new_R1117_U13, new_R1117_U14, new_R1117_U15,
    new_R1117_U16, new_R1117_U17, new_R1117_U18, new_R1117_U19,
    new_R1117_U20, new_R1117_U21, new_R1117_U22, new_R1117_U23,
    new_R1117_U24, new_R1117_U25, new_R1117_U26, new_R1117_U27,
    new_R1117_U28, new_R1117_U29, new_R1117_U30, new_R1117_U31,
    new_R1117_U32, new_R1117_U33, new_R1117_U34, new_R1117_U35,
    new_R1117_U36, new_R1117_U37, new_R1117_U38, new_R1117_U39,
    new_R1117_U40, new_R1117_U41, new_R1117_U42, new_R1117_U43,
    new_R1117_U44, new_R1117_U45, new_R1117_U46, new_R1117_U47,
    new_R1117_U48, new_R1117_U49, new_R1117_U50, new_R1117_U51,
    new_R1117_U52, new_R1117_U53, new_R1117_U54, new_R1117_U55,
    new_R1117_U56, new_R1117_U57, new_R1117_U58, new_R1117_U59,
    new_R1117_U60, new_R1117_U61, new_R1117_U62, new_R1117_U63,
    new_R1117_U64, new_R1117_U65, new_R1117_U66, new_R1117_U67,
    new_R1117_U68, new_R1117_U69, new_R1117_U70, new_R1117_U71,
    new_R1117_U72, new_R1117_U73, new_R1117_U74, new_R1117_U75,
    new_R1117_U76, new_R1117_U77, new_R1117_U78, new_R1117_U79,
    new_R1117_U80, new_R1117_U81, new_R1117_U82, new_R1117_U83,
    new_R1117_U84, new_R1117_U85, new_R1117_U86, new_R1117_U87,
    new_R1117_U88, new_R1117_U89, new_R1117_U90, new_R1117_U91,
    new_R1117_U92, new_R1117_U93, new_R1117_U94, new_R1117_U95,
    new_R1117_U96, new_R1117_U97, new_R1117_U98, new_R1117_U99,
    new_R1117_U100, new_R1117_U101, new_R1117_U102, new_R1117_U103,
    new_R1117_U104, new_R1117_U105, new_R1117_U106, new_R1117_U107,
    new_R1117_U108, new_R1117_U109, new_R1117_U110, new_R1117_U111,
    new_R1117_U112, new_R1117_U113, new_R1117_U114, new_R1117_U115,
    new_R1117_U116, new_R1117_U117, new_R1117_U118, new_R1117_U119,
    new_R1117_U120, new_R1117_U121, new_R1117_U122, new_R1117_U123,
    new_R1117_U124, new_R1117_U125, new_R1117_U126, new_R1117_U127,
    new_R1117_U128, new_R1117_U129, new_R1117_U130, new_R1117_U131,
    new_R1117_U132, new_R1117_U133, new_R1117_U134, new_R1117_U135,
    new_R1117_U136, new_R1117_U137, new_R1117_U138, new_R1117_U139,
    new_R1117_U140, new_R1117_U141, new_R1117_U142, new_R1117_U143,
    new_R1117_U144, new_R1117_U145, new_R1117_U146, new_R1117_U147,
    new_R1117_U148, new_R1117_U149, new_R1117_U150, new_R1117_U151,
    new_R1117_U152, new_R1117_U153, new_R1117_U154, new_R1117_U155,
    new_R1117_U156, new_R1117_U157, new_R1117_U158, new_R1117_U159,
    new_R1117_U160, new_R1117_U161, new_R1117_U162, new_R1117_U163,
    new_R1117_U164, new_R1117_U165, new_R1117_U166, new_R1117_U167,
    new_R1117_U168, new_R1117_U169, new_R1117_U170, new_R1117_U171,
    new_R1117_U172, new_R1117_U173, new_R1117_U174, new_R1117_U175,
    new_R1117_U176, new_R1117_U177, new_R1117_U178, new_R1117_U179,
    new_R1117_U180, new_R1117_U181, new_R1117_U182, new_R1117_U183,
    new_R1117_U184, new_R1117_U185, new_R1117_U186, new_R1117_U187,
    new_R1117_U188, new_R1117_U189, new_R1117_U190, new_R1117_U191,
    new_R1117_U192, new_R1117_U193, new_R1117_U194, new_R1117_U195,
    new_R1117_U196, new_R1117_U197, new_R1117_U198, new_R1117_U199,
    new_R1117_U200, new_R1117_U201, new_R1117_U202, new_R1117_U203,
    new_R1117_U204, new_R1117_U205, new_R1117_U206, new_R1117_U207,
    new_R1117_U208, new_R1117_U209, new_R1117_U210, new_R1117_U211,
    new_R1117_U212, new_R1117_U213, new_R1117_U214, new_R1117_U215,
    new_R1117_U216, new_R1117_U217, new_R1117_U218, new_R1117_U219,
    new_R1117_U220, new_R1117_U221, new_R1117_U222, new_R1117_U223,
    new_R1117_U224, new_R1117_U225, new_R1117_U226, new_R1117_U227,
    new_R1117_U228, new_R1117_U229, new_R1117_U230, new_R1117_U231,
    new_R1117_U232, new_R1117_U233, new_R1117_U234, new_R1117_U235,
    new_R1117_U236, new_R1117_U237, new_R1117_U238, new_R1117_U239,
    new_R1117_U240, new_R1117_U241, new_R1117_U242, new_R1117_U243,
    new_R1117_U244, new_R1117_U245, new_R1117_U246, new_R1117_U247,
    new_R1117_U248, new_R1117_U249, new_R1117_U250, new_R1117_U251,
    new_R1117_U252, new_R1117_U253, new_R1117_U254, new_R1117_U255,
    new_R1117_U256, new_R1117_U257, new_R1117_U258, new_R1117_U259,
    new_R1117_U260, new_R1117_U261, new_R1117_U262, new_R1117_U263,
    new_R1117_U264, new_R1117_U265, new_R1117_U266, new_R1117_U267,
    new_R1117_U268, new_R1117_U269, new_R1117_U270, new_R1117_U271,
    new_R1117_U272, new_R1117_U273, new_R1117_U274, new_R1117_U275,
    new_R1117_U276, new_R1117_U277, new_R1117_U278, new_R1117_U279,
    new_R1117_U280, new_R1117_U281, new_R1117_U282, new_R1117_U283,
    new_R1117_U284, new_R1117_U285, new_R1117_U286, new_R1117_U287,
    new_R1117_U288, new_R1117_U289, new_R1117_U290, new_R1117_U291,
    new_R1117_U292, new_R1117_U293, new_R1117_U294, new_R1117_U295,
    new_R1117_U296, new_R1117_U297, new_R1117_U298, new_R1117_U299,
    new_R1117_U300, new_R1117_U301, new_R1117_U302, new_R1117_U303,
    new_R1117_U304, new_R1117_U305, new_R1117_U306, new_R1117_U307,
    new_R1117_U308, new_R1117_U309, new_R1117_U310, new_R1117_U311,
    new_R1117_U312, new_R1117_U313, new_R1117_U314, new_R1117_U315,
    new_R1117_U316, new_R1117_U317, new_R1117_U318, new_R1117_U319,
    new_R1117_U320, new_R1117_U321, new_R1117_U322, new_R1117_U323,
    new_R1117_U324, new_R1117_U325, new_R1117_U326, new_R1117_U327,
    new_R1117_U328, new_R1117_U329, new_R1117_U330, new_R1117_U331,
    new_R1117_U332, new_R1117_U333, new_R1117_U334, new_R1117_U335,
    new_R1117_U336, new_R1117_U337, new_R1117_U338, new_R1117_U339,
    new_R1117_U340, new_R1117_U341, new_R1117_U342, new_R1117_U343,
    new_R1117_U344, new_R1117_U345, new_R1117_U346, new_R1117_U347,
    new_R1117_U348, new_R1117_U349, new_R1117_U350, new_R1117_U351,
    new_R1117_U352, new_R1117_U353, new_R1117_U354, new_R1117_U355,
    new_R1117_U356, new_R1117_U357, new_R1117_U358, new_R1117_U359,
    new_R1117_U360, new_R1117_U361, new_R1117_U362, new_R1117_U363,
    new_R1117_U364, new_R1117_U365, new_R1117_U366, new_R1117_U367,
    new_R1117_U368, new_R1117_U369, new_R1117_U370, new_R1117_U371,
    new_R1117_U372, new_R1117_U373, new_R1117_U374, new_R1117_U375,
    new_R1117_U376, new_R1117_U377, new_R1117_U378, new_R1117_U379,
    new_R1117_U380, new_R1117_U381, new_R1117_U382, new_R1117_U383,
    new_R1117_U384, new_R1117_U385, new_R1117_U386, new_R1117_U387,
    new_R1117_U388, new_R1117_U389, new_R1117_U390, new_R1117_U391,
    new_R1117_U392, new_R1117_U393, new_R1117_U394, new_R1117_U395,
    new_R1117_U396, new_R1117_U397, new_R1117_U398, new_R1117_U399,
    new_R1117_U400, new_R1117_U401, new_R1117_U402, new_R1117_U403,
    new_R1117_U404, new_R1117_U405, new_R1117_U406, new_R1117_U407,
    new_R1117_U408, new_R1117_U409, new_R1117_U410, new_R1117_U411,
    new_R1117_U412, new_R1117_U413, new_R1117_U414, new_R1117_U415,
    new_R1117_U416, new_R1117_U417, new_R1117_U418, new_R1117_U419,
    new_R1117_U420, new_R1117_U421, new_R1117_U422, new_R1117_U423,
    new_R1117_U424, new_R1117_U425, new_R1117_U426, new_R1117_U427,
    new_R1117_U428, new_R1117_U429, new_R1117_U430, new_R1117_U431,
    new_R1117_U432, new_R1117_U433, new_R1117_U434, new_R1117_U435,
    new_R1117_U436, new_R1117_U437, new_R1117_U438, new_R1117_U439,
    new_R1117_U440, new_R1117_U441, new_R1117_U442, new_R1117_U443,
    new_R1117_U444, new_R1117_U445, new_R1117_U446, new_R1117_U447,
    new_R1117_U448, new_R1117_U449, new_R1117_U450, new_R1117_U451,
    new_R1117_U452, new_R1117_U453, new_R1117_U454, new_R1117_U455,
    new_R1117_U456, new_R1117_U457, new_R1117_U458, new_R1117_U459,
    new_R1117_U460, new_R1117_U461, new_R1117_U462, new_R1117_U463,
    new_R1117_U464, new_R1117_U465, new_R1117_U466, new_R1117_U467,
    new_R1117_U468, new_R1117_U469, new_R1117_U470, new_R1117_U471,
    new_R1117_U472, new_R1117_U473, new_R1117_U474, new_R1117_U475,
    new_R1117_U476, new_R1117_U477, new_R1117_U478, new_R1117_U479,
    new_R1117_U480, new_R1117_U481, new_R1117_U482, new_R1117_U483,
    new_R1117_U484, new_R1117_U485, new_R1117_U486, new_R1117_U487,
    new_R1117_U488, new_R1117_U489, new_R1117_U490, new_R1117_U491,
    new_R1117_U492, new_R1117_U493, new_R1117_U494, new_R1117_U495,
    new_R1117_U496, new_R1117_U497, new_R1117_U498, new_R1117_U499,
    new_R1117_U500, new_R1117_U501, new_R1117_U502, new_R1117_U503,
    new_R1117_U504, new_R1117_U505, new_R1117_U506, new_R1117_U507,
    new_R1117_U508, new_R1117_U509, new_R1117_U510, new_R1117_U511,
    new_R1117_U512, new_R1117_U513, new_R1117_U514, new_R1117_U515,
    new_R1375_U6, new_R1375_U7, new_R1375_U8, new_R1375_U9, new_R1375_U10,
    new_R1375_U11, new_R1375_U12, new_R1375_U13, new_R1375_U14,
    new_R1375_U15, new_R1375_U16, new_R1375_U17, new_R1375_U18,
    new_R1375_U19, new_R1375_U20, new_R1375_U21, new_R1375_U22,
    new_R1375_U23, new_R1375_U24, new_R1375_U25, new_R1375_U26,
    new_R1375_U27, new_R1375_U28, new_R1375_U29, new_R1375_U30,
    new_R1375_U31, new_R1375_U32, new_R1375_U33, new_R1375_U34,
    new_R1375_U35, new_R1375_U36, new_R1375_U37, new_R1375_U38,
    new_R1375_U39, new_R1375_U40, new_R1375_U41, new_R1375_U42,
    new_R1375_U43, new_R1375_U44, new_R1375_U45, new_R1375_U46,
    new_R1375_U47, new_R1375_U48, new_R1375_U49, new_R1375_U50,
    new_R1375_U51, new_R1375_U52, new_R1375_U53, new_R1375_U54,
    new_R1375_U55, new_R1375_U56, new_R1375_U57, new_R1375_U58,
    new_R1375_U59, new_R1375_U60, new_R1375_U61, new_R1375_U62,
    new_R1375_U63, new_R1375_U64, new_R1375_U65, new_R1375_U66,
    new_R1375_U67, new_R1375_U68, new_R1375_U69, new_R1375_U70,
    new_R1375_U71, new_R1375_U72, new_R1375_U73, new_R1375_U74,
    new_R1375_U75, new_R1375_U76, new_R1375_U77, new_R1375_U78,
    new_R1375_U79, new_R1375_U80, new_R1375_U81, new_R1375_U82,
    new_R1375_U83, new_R1375_U84, new_R1375_U85, new_R1375_U86,
    new_R1375_U87, new_R1375_U88, new_R1375_U89, new_R1375_U90,
    new_R1375_U91, new_R1375_U92, new_R1375_U93, new_R1375_U94,
    new_R1375_U95, new_R1375_U96, new_R1375_U97, new_R1375_U98,
    new_R1375_U99, new_R1375_U100, new_R1375_U101, new_R1375_U102,
    new_R1375_U103, new_R1375_U104, new_R1375_U105, new_R1375_U106,
    new_R1375_U107, new_R1375_U108, new_R1375_U109, new_R1375_U110,
    new_R1375_U111, new_R1375_U112, new_R1375_U113, new_R1375_U114,
    new_R1375_U115, new_R1375_U116, new_R1375_U117, new_R1375_U118,
    new_R1375_U119, new_R1375_U120, new_R1375_U121, new_R1375_U122,
    new_R1375_U123, new_R1375_U124, new_R1375_U125, new_R1375_U126,
    new_R1375_U127, new_R1375_U128, new_R1375_U129, new_R1375_U130,
    new_R1375_U131, new_R1375_U132, new_R1375_U133, new_R1375_U134,
    new_R1375_U135, new_R1375_U136, new_R1375_U137, new_R1375_U138,
    new_R1375_U139, new_R1375_U140, new_R1375_U141, new_R1375_U142,
    new_R1375_U143, new_R1375_U144, new_R1375_U145, new_R1375_U146,
    new_R1375_U147, new_R1375_U148, new_R1375_U149, new_R1375_U150,
    new_R1375_U151, new_R1375_U152, new_R1375_U153, new_R1375_U154,
    new_R1375_U155, new_R1375_U156, new_R1375_U157, new_R1375_U158,
    new_R1375_U159, new_R1375_U160, new_R1375_U161, new_R1375_U162,
    new_R1375_U163, new_R1375_U164, new_R1375_U165, new_R1375_U166,
    new_R1375_U167, new_R1375_U168, new_R1375_U169, new_R1375_U170,
    new_R1375_U171, new_R1375_U172, new_R1375_U173, new_R1375_U174,
    new_R1375_U175, new_R1375_U176, new_R1375_U177, new_R1375_U178,
    new_R1375_U179, new_R1375_U180, new_R1375_U181, new_R1375_U182,
    new_R1375_U183, new_R1375_U184, new_R1375_U185, new_R1375_U186,
    new_R1375_U187, new_R1375_U188, new_R1375_U189, new_R1375_U190,
    new_R1375_U191, new_R1375_U192, new_R1375_U193, new_R1375_U194,
    new_R1375_U195, new_R1375_U196, new_R1375_U197, new_R1375_U198,
    new_R1375_U199, new_R1375_U200, new_R1375_U201, new_R1375_U202,
    new_R1375_U203, new_R1375_U204, new_R1375_U205, new_R1375_U206,
    new_R1375_U207, new_R1375_U208, new_R1375_U209, new_R1375_U210,
    new_R1375_U211, new_R1375_U212, new_R1375_U213, new_R1375_U214,
    new_R1375_U215, new_R1375_U216, new_R1375_U217, new_R1375_U218,
    new_R1375_U219, new_R1375_U220, new_R1375_U221, new_R1375_U222,
    new_R1375_U223, new_R1375_U224, new_R1375_U225, new_R1352_U6,
    new_R1352_U7, new_R1207_U6, new_R1207_U7, new_R1207_U8, new_R1207_U9,
    new_R1207_U10, new_R1207_U11, new_R1207_U12, new_R1207_U13,
    new_R1207_U14, new_R1207_U15, new_R1207_U16, new_R1207_U17,
    new_R1207_U18, new_R1207_U19, new_R1207_U20, new_R1207_U21,
    new_R1207_U22, new_R1207_U23, new_R1207_U24, new_R1207_U25,
    new_R1207_U26, new_R1207_U27, new_R1207_U28, new_R1207_U29,
    new_R1207_U30, new_R1207_U31, new_R1207_U32, new_R1207_U33,
    new_R1207_U34, new_R1207_U35, new_R1207_U36, new_R1207_U37,
    new_R1207_U38, new_R1207_U39, new_R1207_U40, new_R1207_U41,
    new_R1207_U42, new_R1207_U43, new_R1207_U44, new_R1207_U45,
    new_R1207_U46, new_R1207_U47, new_R1207_U48, new_R1207_U49,
    new_R1207_U50, new_R1207_U51, new_R1207_U52, new_R1207_U53,
    new_R1207_U54, new_R1207_U55, new_R1207_U56, new_R1207_U57,
    new_R1207_U58, new_R1207_U59, new_R1207_U60, new_R1207_U61,
    new_R1207_U62, new_R1207_U63, new_R1207_U64, new_R1207_U65,
    new_R1207_U66, new_R1207_U67, new_R1207_U68, new_R1207_U69,
    new_R1207_U70, new_R1207_U71, new_R1207_U72, new_R1207_U73,
    new_R1207_U74, new_R1207_U75, new_R1207_U76, new_R1207_U77,
    new_R1207_U78, new_R1207_U79, new_R1207_U80, new_R1207_U81,
    new_R1207_U82, new_R1207_U83, new_R1207_U84, new_R1207_U85,
    new_R1207_U86, new_R1207_U87, new_R1207_U88, new_R1207_U89,
    new_R1207_U90, new_R1207_U91, new_R1207_U92, new_R1207_U93,
    new_R1207_U94, new_R1207_U95, new_R1207_U96, new_R1207_U97,
    new_R1207_U98, new_R1207_U99, new_R1207_U100, new_R1207_U101,
    new_R1207_U102, new_R1207_U103, new_R1207_U104, new_R1207_U105,
    new_R1207_U106, new_R1207_U107, new_R1207_U108, new_R1207_U109,
    new_R1207_U110, new_R1207_U111, new_R1207_U112, new_R1207_U113,
    new_R1207_U114, new_R1207_U115, new_R1207_U116, new_R1207_U117,
    new_R1207_U118, new_R1207_U119, new_R1207_U120, new_R1207_U121,
    new_R1207_U122, new_R1207_U123, new_R1207_U124, new_R1207_U125,
    new_R1207_U126, new_R1207_U127, new_R1207_U128, new_R1207_U129,
    new_R1207_U130, new_R1207_U131, new_R1207_U132, new_R1207_U133,
    new_R1207_U134, new_R1207_U135, new_R1207_U136, new_R1207_U137,
    new_R1207_U138, new_R1207_U139, new_R1207_U140, new_R1207_U141,
    new_R1207_U142, new_R1207_U143, new_R1207_U144, new_R1207_U145,
    new_R1207_U146, new_R1207_U147, new_R1207_U148, new_R1207_U149,
    new_R1207_U150, new_R1207_U151, new_R1207_U152, new_R1207_U153,
    new_R1207_U154, new_R1207_U155, new_R1207_U156, new_R1207_U157,
    new_R1207_U158, new_R1207_U159, new_R1207_U160, new_R1207_U161,
    new_R1207_U162, new_R1207_U163, new_R1207_U164, new_R1207_U165,
    new_R1207_U166, new_R1207_U167, new_R1207_U168, new_R1207_U169,
    new_R1207_U170, new_R1207_U171, new_R1207_U172, new_R1207_U173,
    new_R1207_U174, new_R1207_U175, new_R1207_U176, new_R1207_U177,
    new_R1207_U178, new_R1207_U179, new_R1207_U180, new_R1207_U181,
    new_R1207_U182, new_R1207_U183, new_R1207_U184, new_R1207_U185,
    new_R1207_U186, new_R1207_U187, new_R1207_U188, new_R1207_U189,
    new_R1207_U190, new_R1207_U191, new_R1207_U192, new_R1207_U193,
    new_R1207_U194, new_R1207_U195, new_R1207_U196, new_R1207_U197,
    new_R1207_U198, new_R1207_U199, new_R1207_U200, new_R1207_U201,
    new_R1207_U202, new_R1207_U203, new_R1207_U204, new_R1207_U205,
    new_R1207_U206, new_R1207_U207, new_R1207_U208, new_R1207_U209,
    new_R1207_U210, new_R1207_U211, new_R1207_U212, new_R1207_U213,
    new_R1207_U214, new_R1207_U215, new_R1207_U216, new_R1207_U217,
    new_R1207_U218, new_R1207_U219, new_R1207_U220, new_R1207_U221,
    new_R1207_U222, new_R1207_U223, new_R1207_U224, new_R1207_U225,
    new_R1207_U226, new_R1207_U227, new_R1207_U228, new_R1207_U229,
    new_R1207_U230, new_R1207_U231, new_R1207_U232, new_R1207_U233,
    new_R1207_U234, new_R1207_U235, new_R1207_U236, new_R1207_U237,
    new_R1207_U238, new_R1207_U239, new_R1207_U240, new_R1207_U241,
    new_R1207_U242, new_R1207_U243, new_R1207_U244, new_R1207_U245,
    new_R1207_U246, new_R1207_U247, new_R1207_U248, new_R1207_U249,
    new_R1207_U250, new_R1207_U251, new_R1207_U252, new_R1207_U253,
    new_R1207_U254, new_R1207_U255, new_R1207_U256, new_R1207_U257,
    new_R1207_U258, new_R1207_U259, new_R1207_U260, new_R1207_U261,
    new_R1207_U262, new_R1207_U263, new_R1207_U264, new_R1207_U265,
    new_R1207_U266, new_R1207_U267, new_R1207_U268, new_R1207_U269,
    new_R1207_U270, new_R1207_U271, new_R1207_U272, new_R1207_U273,
    new_R1207_U274, new_R1207_U275, new_R1207_U276, new_R1207_U277,
    new_R1207_U278, new_R1207_U279, new_R1207_U280, new_R1207_U281,
    new_R1207_U282, new_R1207_U283, new_R1207_U284, new_R1207_U285,
    new_R1207_U286, new_R1207_U287, new_R1207_U288, new_R1207_U289,
    new_R1207_U290, new_R1207_U291, new_R1207_U292, new_R1207_U293,
    new_R1207_U294, new_R1207_U295, new_R1207_U296, new_R1207_U297,
    new_R1207_U298, new_R1207_U299, new_R1207_U300, new_R1207_U301,
    new_R1207_U302, new_R1207_U303, new_R1207_U304, new_R1207_U305,
    new_R1207_U306, new_R1207_U307, new_R1207_U308, new_R1207_U309,
    new_R1207_U310, new_R1207_U311, new_R1207_U312, new_R1207_U313,
    new_R1207_U314, new_R1207_U315, new_R1207_U316, new_R1207_U317,
    new_R1207_U318, new_R1207_U319, new_R1207_U320, new_R1207_U321,
    new_R1207_U322, new_R1207_U323, new_R1207_U324, new_R1207_U325,
    new_R1207_U326, new_R1207_U327, new_R1207_U328, new_R1207_U329,
    new_R1207_U330, new_R1207_U331, new_R1207_U332, new_R1207_U333,
    new_R1207_U334, new_R1207_U335, new_R1207_U336, new_R1207_U337,
    new_R1207_U338, new_R1207_U339, new_R1207_U340, new_R1207_U341,
    new_R1207_U342, new_R1207_U343, new_R1207_U344, new_R1207_U345,
    new_R1207_U346, new_R1207_U347, new_R1207_U348, new_R1207_U349,
    new_R1207_U350, new_R1207_U351, new_R1207_U352, new_R1207_U353,
    new_R1207_U354, new_R1207_U355, new_R1207_U356, new_R1207_U357,
    new_R1207_U358, new_R1207_U359, new_R1207_U360, new_R1207_U361,
    new_R1207_U362, new_R1207_U363, new_R1207_U364, new_R1207_U365,
    new_R1207_U366, new_R1207_U367, new_R1207_U368, new_R1207_U369,
    new_R1207_U370, new_R1207_U371, new_R1207_U372, new_R1207_U373,
    new_R1207_U374, new_R1207_U375, new_R1207_U376, new_R1207_U377,
    new_R1207_U378, new_R1207_U379, new_R1207_U380, new_R1207_U381,
    new_R1207_U382, new_R1207_U383, new_R1207_U384, new_R1207_U385,
    new_R1207_U386, new_R1207_U387, new_R1207_U388, new_R1207_U389,
    new_R1207_U390, new_R1207_U391, new_R1207_U392, new_R1207_U393,
    new_R1207_U394, new_R1207_U395, new_R1207_U396, new_R1207_U397,
    new_R1207_U398, new_R1207_U399, new_R1207_U400, new_R1207_U401,
    new_R1207_U402, new_R1207_U403, new_R1207_U404, new_R1207_U405,
    new_R1207_U406, new_R1207_U407, new_R1207_U408, new_R1207_U409,
    new_R1207_U410, new_R1207_U411, new_R1207_U412, new_R1207_U413,
    new_R1207_U414, new_R1207_U415, new_R1207_U416, new_R1207_U417,
    new_R1207_U418, new_R1207_U419, new_R1207_U420, new_R1207_U421,
    new_R1207_U422, new_R1207_U423, new_R1207_U424, new_R1207_U425,
    new_R1207_U426, new_R1207_U427, new_R1207_U428, new_R1207_U429,
    new_R1207_U430, new_R1207_U431, new_R1207_U432, new_R1207_U433,
    new_R1207_U434, new_R1207_U435, new_R1207_U436, new_R1207_U437,
    new_R1207_U438, new_R1207_U439, new_R1207_U440, new_R1207_U441,
    new_R1207_U442, new_R1207_U443, new_R1207_U444, new_R1207_U445,
    new_R1207_U446, new_R1207_U447, new_R1207_U448, new_R1207_U449,
    new_R1207_U450, new_R1207_U451, new_R1207_U452, new_R1207_U453,
    new_R1207_U454, new_R1207_U455, new_R1207_U456, new_R1207_U457,
    new_R1207_U458, new_R1207_U459, new_R1207_U460, new_R1207_U461,
    new_R1207_U462, new_R1207_U463, new_R1207_U464, new_R1207_U465,
    new_R1207_U466, new_R1207_U467, new_R1207_U468, new_R1207_U469,
    new_R1207_U470, new_R1207_U471, new_R1207_U472, new_R1207_U473,
    new_R1207_U474, new_R1207_U475, new_R1207_U476, new_R1207_U477,
    new_R1207_U478, new_R1207_U479, new_R1207_U480, new_R1207_U481,
    new_R1207_U482, new_R1207_U483, new_R1207_U484, new_R1207_U485,
    new_R1207_U486, new_R1207_U487, new_R1207_U488, new_R1207_U489,
    new_R1207_U490, new_R1207_U491, new_R1207_U492, new_R1207_U493,
    new_R1207_U494, new_R1207_U495, new_R1207_U496, new_R1207_U497,
    new_R1207_U498, new_R1207_U499, new_R1207_U500, new_R1207_U501,
    new_R1207_U502, new_R1207_U503, new_R1207_U504, new_R1207_U505,
    new_R1207_U506, new_R1207_U507, new_R1207_U508, new_R1207_U509,
    new_R1207_U510, new_R1207_U511, new_R1207_U512, new_R1207_U513,
    new_R1207_U514, new_R1207_U515, new_R1207_U516, new_R1207_U517,
    new_R1207_U518, new_R1207_U519, new_R1207_U520, new_R1165_U4,
    new_R1165_U5, new_R1165_U6, new_R1165_U7, new_R1165_U8, new_R1165_U9,
    new_R1165_U10, new_R1165_U11, new_R1165_U12, new_R1165_U13,
    new_R1165_U14, new_R1165_U15, new_R1165_U16, new_R1165_U17,
    new_R1165_U18, new_R1165_U19, new_R1165_U20, new_R1165_U21,
    new_R1165_U22, new_R1165_U23, new_R1165_U24, new_R1165_U25,
    new_R1165_U26, new_R1165_U27, new_R1165_U28, new_R1165_U29,
    new_R1165_U30, new_R1165_U31, new_R1165_U32, new_R1165_U33,
    new_R1165_U34, new_R1165_U35, new_R1165_U36, new_R1165_U37,
    new_R1165_U38, new_R1165_U39, new_R1165_U40, new_R1165_U41,
    new_R1165_U42, new_R1165_U43, new_R1165_U44, new_R1165_U45,
    new_R1165_U46, new_R1165_U47, new_R1165_U48, new_R1165_U49,
    new_R1165_U50, new_R1165_U51, new_R1165_U52, new_R1165_U53,
    new_R1165_U54, new_R1165_U55, new_R1165_U56, new_R1165_U57,
    new_R1165_U58, new_R1165_U59, new_R1165_U60, new_R1165_U61,
    new_R1165_U62, new_R1165_U63, new_R1165_U64, new_R1165_U65,
    new_R1165_U66, new_R1165_U67, new_R1165_U68, new_R1165_U69,
    new_R1165_U70, new_R1165_U71, new_R1165_U72, new_R1165_U73,
    new_R1165_U74, new_R1165_U75, new_R1165_U76, new_R1165_U77,
    new_R1165_U78, new_R1165_U79, new_R1165_U80, new_R1165_U81,
    new_R1165_U82, new_R1165_U83, new_R1165_U84, new_R1165_U85,
    new_R1165_U86, new_R1165_U87, new_R1165_U88, new_R1165_U89,
    new_R1165_U90, new_R1165_U91, new_R1165_U92, new_R1165_U93,
    new_R1165_U94, new_R1165_U95, new_R1165_U96, new_R1165_U97,
    new_R1165_U98, new_R1165_U99, new_R1165_U100, new_R1165_U101,
    new_R1165_U102, new_R1165_U103, new_R1165_U104, new_R1165_U105,
    new_R1165_U106, new_R1165_U107, new_R1165_U108, new_R1165_U109,
    new_R1165_U110, new_R1165_U111, new_R1165_U112, new_R1165_U113,
    new_R1165_U114, new_R1165_U115, new_R1165_U116, new_R1165_U117,
    new_R1165_U118, new_R1165_U119, new_R1165_U120, new_R1165_U121,
    new_R1165_U122, new_R1165_U123, new_R1165_U124, new_R1165_U125,
    new_R1165_U126, new_R1165_U127, new_R1165_U128, new_R1165_U129,
    new_R1165_U130, new_R1165_U131, new_R1165_U132, new_R1165_U133,
    new_R1165_U134, new_R1165_U135, new_R1165_U136, new_R1165_U137,
    new_R1165_U138, new_R1165_U139, new_R1165_U140, new_R1165_U141,
    new_R1165_U142, new_R1165_U143, new_R1165_U144, new_R1165_U145,
    new_R1165_U146, new_R1165_U147, new_R1165_U148, new_R1165_U149,
    new_R1165_U150, new_R1165_U151, new_R1165_U152, new_R1165_U153,
    new_R1165_U154, new_R1165_U155, new_R1165_U156, new_R1165_U157,
    new_R1165_U158, new_R1165_U159, new_R1165_U160, new_R1165_U161,
    new_R1165_U162, new_R1165_U163, new_R1165_U164, new_R1165_U165,
    new_R1165_U166, new_R1165_U167, new_R1165_U168, new_R1165_U169,
    new_R1165_U170, new_R1165_U171, new_R1165_U172, new_R1165_U173,
    new_R1165_U174, new_R1165_U175, new_R1165_U176, new_R1165_U177,
    new_R1165_U178, new_R1165_U179, new_R1165_U180, new_R1165_U181,
    new_R1165_U182, new_R1165_U183, new_R1165_U184, new_R1165_U185,
    new_R1165_U186, new_R1165_U187, new_R1165_U188, new_R1165_U189,
    new_R1165_U190, new_R1165_U191, new_R1165_U192, new_R1165_U193,
    new_R1165_U194, new_R1165_U195, new_R1165_U196, new_R1165_U197,
    new_R1165_U198, new_R1165_U199, new_R1165_U200, new_R1165_U201,
    new_R1165_U202, new_R1165_U203, new_R1165_U204, new_R1165_U205,
    new_R1165_U206, new_R1165_U207, new_R1165_U208, new_R1165_U209,
    new_R1165_U210, new_R1165_U211, new_R1165_U212, new_R1165_U213,
    new_R1165_U214, new_R1165_U215, new_R1165_U216, new_R1165_U217,
    new_R1165_U218, new_R1165_U219, new_R1165_U220, new_R1165_U221,
    new_R1165_U222, new_R1165_U223, new_R1165_U224, new_R1165_U225,
    new_R1165_U226, new_R1165_U227, new_R1165_U228, new_R1165_U229,
    new_R1165_U230, new_R1165_U231, new_R1165_U232, new_R1165_U233,
    new_R1165_U234, new_R1165_U235, new_R1165_U236, new_R1165_U237,
    new_R1165_U238, new_R1165_U239, new_R1165_U240, new_R1165_U241,
    new_R1165_U242, new_R1165_U243, new_R1165_U244, new_R1165_U245,
    new_R1165_U246, new_R1165_U247, new_R1165_U248, new_R1165_U249,
    new_R1165_U250, new_R1165_U251, new_R1165_U252, new_R1165_U253,
    new_R1165_U254, new_R1165_U255, new_R1165_U256, new_R1165_U257,
    new_R1165_U258, new_R1165_U259, new_R1165_U260, new_R1165_U261,
    new_R1165_U262, new_R1165_U263, new_R1165_U264, new_R1165_U265,
    new_R1165_U266, new_R1165_U267, new_R1165_U268, new_R1165_U269,
    new_R1165_U270, new_R1165_U271, new_R1165_U272, new_R1165_U273,
    new_R1165_U274, new_R1165_U275, new_R1165_U276, new_R1165_U277,
    new_R1165_U278, new_R1165_U279, new_R1165_U280, new_R1165_U281,
    new_R1165_U282, new_R1165_U283, new_R1165_U284, new_R1165_U285,
    new_R1165_U286, new_R1165_U287, new_R1165_U288, new_R1165_U289,
    new_R1165_U290, new_R1165_U291, new_R1165_U292, new_R1165_U293,
    new_R1165_U294, new_R1165_U295, new_R1165_U296, new_R1165_U297,
    new_R1165_U298, new_R1165_U299, new_R1165_U300, new_R1165_U301,
    new_R1165_U302, new_R1165_U303, new_R1165_U304, new_R1165_U305,
    new_R1165_U306, new_R1165_U307, new_R1165_U308, new_R1165_U309,
    new_R1165_U310, new_R1165_U311, new_R1165_U312, new_R1165_U313,
    new_R1165_U314, new_R1165_U315, new_R1165_U316, new_R1165_U317,
    new_R1165_U318, new_R1165_U319, new_R1165_U320, new_R1165_U321,
    new_R1165_U322, new_R1165_U323, new_R1165_U324, new_R1165_U325,
    new_R1165_U326, new_R1165_U327, new_R1165_U328, new_R1165_U329,
    new_R1165_U330, new_R1165_U331, new_R1165_U332, new_R1165_U333,
    new_R1165_U334, new_R1165_U335, new_R1165_U336, new_R1165_U337,
    new_R1165_U338, new_R1165_U339, new_R1165_U340, new_R1165_U341,
    new_R1165_U342, new_R1165_U343, new_R1165_U344, new_R1165_U345,
    new_R1165_U346, new_R1165_U347, new_R1165_U348, new_R1165_U349,
    new_R1165_U350, new_R1165_U351, new_R1165_U352, new_R1165_U353,
    new_R1165_U354, new_R1165_U355, new_R1165_U356, new_R1165_U357,
    new_R1165_U358, new_R1165_U359, new_R1165_U360, new_R1165_U361,
    new_R1165_U362, new_R1165_U363, new_R1165_U364, new_R1165_U365,
    new_R1165_U366, new_R1165_U367, new_R1165_U368, new_R1165_U369,
    new_R1165_U370, new_R1165_U371, new_R1165_U372, new_R1165_U373,
    new_R1165_U374, new_R1165_U375, new_R1165_U376, new_R1165_U377,
    new_R1165_U378, new_R1165_U379, new_R1165_U380, new_R1165_U381,
    new_R1165_U382, new_R1165_U383, new_R1165_U384, new_R1165_U385,
    new_R1165_U386, new_R1165_U387, new_R1165_U388, new_R1165_U389,
    new_R1165_U390, new_R1165_U391, new_R1165_U392, new_R1165_U393,
    new_R1165_U394, new_R1165_U395, new_R1165_U396, new_R1165_U397,
    new_R1165_U398, new_R1165_U399, new_R1165_U400, new_R1165_U401,
    new_R1165_U402, new_R1165_U403, new_R1165_U404, new_R1165_U405,
    new_R1165_U406, new_R1165_U407, new_R1165_U408, new_R1165_U409,
    new_R1165_U410, new_R1165_U411, new_R1165_U412, new_R1165_U413,
    new_R1165_U414, new_R1165_U415, new_R1165_U416, new_R1165_U417,
    new_R1165_U418, new_R1165_U419, new_R1165_U420, new_R1165_U421,
    new_R1165_U422, new_R1165_U423, new_R1165_U424, new_R1165_U425,
    new_R1165_U426, new_R1165_U427, new_R1165_U428, new_R1165_U429,
    new_R1165_U430, new_R1165_U431, new_R1165_U432, new_R1165_U433,
    new_R1165_U434, new_R1165_U435, new_R1165_U436, new_R1165_U437,
    new_R1165_U438, new_R1165_U439, new_R1165_U440, new_R1165_U441,
    new_R1165_U442, new_R1165_U443, new_R1165_U444, new_R1165_U445,
    new_R1165_U446, new_R1165_U447, new_R1165_U448, new_R1165_U449,
    new_R1165_U450, new_R1165_U451, new_R1165_U452, new_R1165_U453,
    new_R1165_U454, new_R1165_U455, new_R1165_U456, new_R1165_U457,
    new_R1165_U458, new_R1165_U459, new_R1165_U460, new_R1165_U461,
    new_R1165_U462, new_R1165_U463, new_R1165_U464, new_R1165_U465,
    new_R1165_U466, new_R1165_U467, new_R1165_U468, new_R1165_U469,
    new_R1165_U470, new_R1165_U471, new_R1165_U472, new_R1165_U473,
    new_R1165_U474, new_R1165_U475, new_R1165_U476, new_R1165_U477,
    new_R1165_U478, new_R1165_U479, new_R1165_U480, new_R1165_U481,
    new_R1165_U482, new_R1165_U483, new_R1165_U484, new_R1165_U485,
    new_R1165_U486, new_R1165_U487, new_R1165_U488, new_R1165_U489,
    new_R1165_U490, new_R1165_U491, new_R1165_U492, new_R1165_U493,
    new_R1165_U494, new_R1165_U495, new_R1165_U496, new_R1165_U497,
    new_R1165_U498, new_R1165_U499, new_R1165_U500, new_R1165_U501,
    new_R1165_U502, new_R1165_U503, new_R1165_U504, new_R1165_U505,
    new_R1165_U506, new_R1165_U507, new_R1165_U508, new_R1165_U509,
    new_R1165_U510, new_R1165_U511, new_R1165_U512, new_R1165_U513,
    new_R1165_U514, new_R1165_U515, new_R1165_U516, new_R1165_U517,
    new_R1165_U518, new_R1165_U519, new_R1165_U520, new_R1165_U521,
    new_R1165_U522, new_R1165_U523, new_R1165_U524, new_R1165_U525,
    new_R1165_U526, new_R1165_U527, new_R1165_U528, new_R1165_U529,
    new_R1165_U530, new_R1165_U531, new_R1165_U532, new_R1165_U533,
    new_R1165_U534, new_R1165_U535, new_R1165_U536, new_R1165_U537,
    new_R1165_U538, new_R1165_U539, new_R1165_U540, new_R1165_U541,
    new_R1165_U542, new_R1165_U543, new_R1165_U544, new_R1165_U545,
    new_R1165_U546, new_R1165_U547, new_R1165_U548, new_R1165_U549,
    new_R1165_U550, new_R1165_U551, new_R1165_U552, new_R1165_U553,
    new_R1165_U554, new_R1165_U555, new_R1165_U556, new_R1165_U557,
    new_R1165_U558, new_R1165_U559, new_R1165_U560, new_R1165_U561,
    new_R1165_U562, new_R1165_U563, new_R1165_U564, new_R1165_U565,
    new_R1165_U566, new_R1165_U567, new_R1165_U568, new_R1165_U569,
    new_R1165_U570, new_R1165_U571, new_R1165_U572, new_R1165_U573,
    new_R1165_U574, new_R1165_U575, new_R1165_U576, new_R1165_U577,
    new_R1165_U578, new_R1165_U579, new_R1165_U580, new_R1165_U581,
    new_R1165_U582, new_R1165_U583, new_R1165_U584, new_R1165_U585,
    new_R1165_U586, new_R1165_U587, new_R1165_U588, new_R1165_U589,
    new_R1165_U590, new_R1165_U591, new_R1165_U592, new_R1165_U593,
    new_R1165_U594, new_R1165_U595, new_R1165_U596, new_R1165_U597,
    new_R1165_U598, new_R1165_U599, new_R1165_U600, new_R1165_U601,
    new_R1165_U602, new_R1165_U603, new_R1165_U604, new_R1165_U605,
    new_R1165_U606, new_R1165_U607, new_R1165_U608, new_R1165_U609,
    new_R1165_U610, new_R1165_U611, new_R1165_U612, new_R1165_U613,
    new_R1150_U6, new_R1150_U7, new_R1150_U8, new_R1150_U9, new_R1150_U10,
    new_R1150_U11, new_R1150_U12, new_R1150_U13, new_R1150_U14,
    new_R1150_U15, new_R1150_U16, new_R1150_U17, new_R1150_U18,
    new_R1150_U19, new_R1150_U20, new_R1150_U21, new_R1150_U22,
    new_R1150_U23, new_R1150_U24, new_R1150_U25, new_R1150_U26,
    new_R1150_U27, new_R1150_U28, new_R1150_U29, new_R1150_U30,
    new_R1150_U31, new_R1150_U32, new_R1150_U33, new_R1150_U34,
    new_R1150_U35, new_R1150_U36, new_R1150_U37, new_R1150_U38,
    new_R1150_U39, new_R1150_U40, new_R1150_U41, new_R1150_U42,
    new_R1150_U43, new_R1150_U44, new_R1150_U45, new_R1150_U46,
    new_R1150_U47, new_R1150_U48, new_R1150_U49, new_R1150_U50,
    new_R1150_U51, new_R1150_U52, new_R1150_U53, new_R1150_U54,
    new_R1150_U55, new_R1150_U56, new_R1150_U57, new_R1150_U58,
    new_R1150_U59, new_R1150_U60, new_R1150_U61, new_R1150_U62,
    new_R1150_U63, new_R1150_U64, new_R1150_U65, new_R1150_U66,
    new_R1150_U67, new_R1150_U68, new_R1150_U69, new_R1150_U70,
    new_R1150_U71, new_R1150_U72, new_R1150_U73, new_R1150_U74,
    new_R1150_U75, new_R1150_U76, new_R1150_U77, new_R1150_U78,
    new_R1150_U79, new_R1150_U80, new_R1150_U81, new_R1150_U82,
    new_R1150_U83, new_R1150_U84, new_R1150_U85, new_R1150_U86,
    new_R1150_U87, new_R1150_U88, new_R1150_U89, new_R1150_U90,
    new_R1150_U91, new_R1150_U92, new_R1150_U93, new_R1150_U94,
    new_R1150_U95, new_R1150_U96, new_R1150_U97, new_R1150_U98,
    new_R1150_U99, new_R1150_U100, new_R1150_U101, new_R1150_U102,
    new_R1150_U103, new_R1150_U104, new_R1150_U105, new_R1150_U106,
    new_R1150_U107, new_R1150_U108, new_R1150_U109, new_R1150_U110,
    new_R1150_U111, new_R1150_U112, new_R1150_U113, new_R1150_U114,
    new_R1150_U115, new_R1150_U116, new_R1150_U117, new_R1150_U118,
    new_R1150_U119, new_R1150_U120, new_R1150_U121, new_R1150_U122,
    new_R1150_U123, new_R1150_U124, new_R1150_U125, new_R1150_U126,
    new_R1150_U127, new_R1150_U128, new_R1150_U129, new_R1150_U130,
    new_R1150_U131, new_R1150_U132, new_R1150_U133, new_R1150_U134,
    new_R1150_U135, new_R1150_U136, new_R1150_U137, new_R1150_U138,
    new_R1150_U139, new_R1150_U140, new_R1150_U141, new_R1150_U142,
    new_R1150_U143, new_R1150_U144, new_R1150_U145, new_R1150_U146,
    new_R1150_U147, new_R1150_U148, new_R1150_U149, new_R1150_U150,
    new_R1150_U151, new_R1150_U152, new_R1150_U153, new_R1150_U154,
    new_R1150_U155, new_R1150_U156, new_R1150_U157, new_R1150_U158,
    new_R1150_U159, new_R1150_U160, new_R1150_U161, new_R1150_U162,
    new_R1150_U163, new_R1150_U164, new_R1150_U165, new_R1150_U166,
    new_R1150_U167, new_R1150_U168, new_R1150_U169, new_R1150_U170,
    new_R1150_U171, new_R1150_U172, new_R1150_U173, new_R1150_U174,
    new_R1150_U175, new_R1150_U176, new_R1150_U177, new_R1150_U178,
    new_R1150_U179, new_R1150_U180, new_R1150_U181, new_R1150_U182,
    new_R1150_U183, new_R1150_U184, new_R1150_U185, new_R1150_U186,
    new_R1150_U187, new_R1150_U188, new_R1150_U189, new_R1150_U190,
    new_R1150_U191, new_R1150_U192, new_R1150_U193, new_R1150_U194,
    new_R1150_U195, new_R1150_U196, new_R1150_U197, new_R1150_U198,
    new_R1150_U199, new_R1150_U200, new_R1150_U201, new_R1150_U202,
    new_R1150_U203, new_R1150_U204, new_R1150_U205, new_R1150_U206,
    new_R1150_U207, new_R1150_U208, new_R1150_U209, new_R1150_U210,
    new_R1150_U211, new_R1150_U212, new_R1150_U213, new_R1150_U214,
    new_R1150_U215, new_R1150_U216, new_R1150_U217, new_R1150_U218,
    new_R1150_U219, new_R1150_U220, new_R1150_U221, new_R1150_U222,
    new_R1150_U223, new_R1150_U224, new_R1150_U225, new_R1150_U226,
    new_R1150_U227, new_R1150_U228, new_R1150_U229, new_R1150_U230,
    new_R1150_U231, new_R1150_U232, new_R1150_U233, new_R1150_U234,
    new_R1150_U235, new_R1150_U236, new_R1150_U237, new_R1150_U238,
    new_R1150_U239, new_R1150_U240, new_R1150_U241, new_R1150_U242,
    new_R1150_U243, new_R1150_U244, new_R1150_U245, new_R1150_U246,
    new_R1150_U247, new_R1150_U248, new_R1150_U249, new_R1150_U250,
    new_R1150_U251, new_R1150_U252, new_R1150_U253, new_R1150_U254,
    new_R1150_U255, new_R1150_U256, new_R1150_U257, new_R1150_U258,
    new_R1150_U259, new_R1150_U260, new_R1150_U261, new_R1150_U262,
    new_R1150_U263, new_R1150_U264, new_R1150_U265, new_R1150_U266,
    new_R1150_U267, new_R1150_U268, new_R1150_U269, new_R1150_U270,
    new_R1150_U271, new_R1150_U272, new_R1150_U273, new_R1150_U274,
    new_R1150_U275, new_R1150_U276, new_R1150_U277, new_R1150_U278,
    new_R1150_U279, new_R1150_U280, new_R1150_U281, new_R1150_U282,
    new_R1150_U283, new_R1150_U284, new_R1150_U285, new_R1150_U286,
    new_R1150_U287, new_R1150_U288, new_R1150_U289, new_R1150_U290,
    new_R1150_U291, new_R1150_U292, new_R1150_U293, new_R1150_U294,
    new_R1150_U295, new_R1150_U296, new_R1150_U297, new_R1150_U298,
    new_R1150_U299, new_R1150_U300, new_R1150_U301, new_R1150_U302,
    new_R1150_U303, new_R1150_U304, new_R1150_U305, new_R1150_U306,
    new_R1150_U307, new_R1150_U308, new_R1150_U309, new_R1150_U310,
    new_R1150_U311, new_R1150_U312, new_R1150_U313, new_R1150_U314,
    new_R1150_U315, new_R1150_U316, new_R1150_U317, new_R1150_U318,
    new_R1150_U319, new_R1150_U320, new_R1150_U321, new_R1150_U322,
    new_R1150_U323, new_R1150_U324, new_R1150_U325, new_R1150_U326,
    new_R1150_U327, new_R1150_U328, new_R1150_U329, new_R1150_U330,
    new_R1150_U331, new_R1150_U332, new_R1150_U333, new_R1150_U334,
    new_R1150_U335, new_R1150_U336, new_R1150_U337, new_R1150_U338,
    new_R1150_U339, new_R1150_U340, new_R1150_U341, new_R1150_U342,
    new_R1150_U343, new_R1150_U344, new_R1150_U345, new_R1150_U346,
    new_R1150_U347, new_R1150_U348, new_R1150_U349, new_R1150_U350,
    new_R1150_U351, new_R1150_U352, new_R1150_U353, new_R1150_U354,
    new_R1150_U355, new_R1150_U356, new_R1150_U357, new_R1150_U358,
    new_R1150_U359, new_R1150_U360, new_R1150_U361, new_R1150_U362,
    new_R1150_U363, new_R1150_U364, new_R1150_U365, new_R1150_U366,
    new_R1150_U367, new_R1150_U368, new_R1150_U369, new_R1150_U370,
    new_R1150_U371, new_R1150_U372, new_R1150_U373, new_R1150_U374,
    new_R1150_U375, new_R1150_U376, new_R1150_U377, new_R1150_U378,
    new_R1150_U379, new_R1150_U380, new_R1150_U381, new_R1150_U382,
    new_R1150_U383, new_R1150_U384, new_R1150_U385, new_R1150_U386,
    new_R1150_U387, new_R1150_U388, new_R1150_U389, new_R1150_U390,
    new_R1150_U391, new_R1150_U392, new_R1150_U393, new_R1150_U394,
    new_R1150_U395, new_R1150_U396, new_R1150_U397, new_R1150_U398,
    new_R1150_U399, new_R1150_U400, new_R1150_U401, new_R1150_U402,
    new_R1150_U403, new_R1150_U404, new_R1150_U405, new_R1150_U406,
    new_R1150_U407, new_R1150_U408, new_R1150_U409, new_R1150_U410,
    new_R1150_U411, new_R1150_U412, new_R1150_U413, new_R1150_U414,
    new_R1150_U415, new_R1150_U416, new_R1150_U417, new_R1150_U418,
    new_R1150_U419, new_R1150_U420, new_R1150_U421, new_R1150_U422,
    new_R1150_U423, new_R1150_U424, new_R1150_U425, new_R1150_U426,
    new_R1150_U427, new_R1150_U428, new_R1150_U429, new_R1150_U430,
    new_R1150_U431, new_R1150_U432, new_R1150_U433, new_R1150_U434,
    new_R1150_U435, new_R1150_U436, new_R1150_U437, new_R1150_U438,
    new_R1150_U439, new_R1150_U440, new_R1150_U441, new_R1150_U442,
    new_R1150_U443, new_R1150_U444, new_R1150_U445, new_R1150_U446,
    new_R1150_U447, new_R1150_U448, new_R1150_U449, new_R1150_U450,
    new_R1150_U451, new_R1150_U452, new_R1150_U453, new_R1150_U454,
    new_R1150_U455, new_R1150_U456, new_R1150_U457, new_R1150_U458,
    new_R1150_U459, new_R1150_U460, new_R1150_U461, new_R1150_U462,
    new_R1150_U463, new_R1150_U464, new_R1150_U465, new_R1150_U466,
    new_R1150_U467, new_R1150_U468, new_R1150_U469, new_R1150_U470,
    new_R1150_U471, new_R1150_U472, new_R1150_U473, new_R1150_U474,
    new_R1150_U475, new_R1150_U476, new_R1150_U477, new_R1150_U478,
    new_R1150_U479, new_R1150_U480, new_R1150_U481, new_R1150_U482,
    new_R1150_U483, new_R1150_U484, new_R1150_U485, new_R1150_U486,
    new_R1150_U487, new_R1150_U488, new_R1150_U489, new_R1150_U490,
    new_R1150_U491, new_R1150_U492, new_R1150_U493, new_R1150_U494,
    new_R1150_U495, new_R1150_U496, new_R1150_U497, new_R1150_U498,
    new_R1150_U499, new_R1150_U500, new_R1150_U501, new_R1150_U502,
    new_R1150_U503, new_R1150_U504, new_R1150_U505, new_R1150_U506,
    new_R1150_U507, new_R1150_U508, new_R1150_U509, new_R1150_U510,
    new_R1150_U511, new_R1192_U6, new_R1192_U7, new_R1192_U8, new_R1192_U9,
    new_R1192_U10, new_R1192_U11, new_R1192_U12, new_R1192_U13,
    new_R1192_U14, new_R1192_U15, new_R1192_U16, new_R1192_U17,
    new_R1192_U18, new_R1192_U19, new_R1192_U20, new_R1192_U21,
    new_R1192_U22, new_R1192_U23, new_R1192_U24, new_R1192_U25,
    new_R1192_U26, new_R1192_U27, new_R1192_U28, new_R1192_U29,
    new_R1192_U30, new_R1192_U31, new_R1192_U32, new_R1192_U33,
    new_R1192_U34, new_R1192_U35, new_R1192_U36, new_R1192_U37,
    new_R1192_U38, new_R1192_U39, new_R1192_U40, new_R1192_U41,
    new_R1192_U42, new_R1192_U43, new_R1192_U44, new_R1192_U45,
    new_R1192_U46, new_R1192_U47, new_R1192_U48, new_R1192_U49,
    new_R1192_U50, new_R1192_U51, new_R1192_U52, new_R1192_U53,
    new_R1192_U54, new_R1192_U55, new_R1192_U56, new_R1192_U57,
    new_R1192_U58, new_R1192_U59, new_R1192_U60, new_R1192_U61,
    new_R1192_U62, new_R1192_U63, new_R1192_U64, new_R1192_U65,
    new_R1192_U66, new_R1192_U67, new_R1192_U68, new_R1192_U69,
    new_R1192_U70, new_R1192_U71, new_R1192_U72, new_R1192_U73,
    new_R1192_U74, new_R1192_U75, new_R1192_U76, new_R1192_U77,
    new_R1192_U78, new_R1192_U79, new_R1192_U80, new_R1192_U81,
    new_R1192_U82, new_R1192_U83, new_R1192_U84, new_R1192_U85,
    new_R1192_U86, new_R1192_U87, new_R1192_U88, new_R1192_U89,
    new_R1192_U90, new_R1192_U91, new_R1192_U92, new_R1192_U93,
    new_R1192_U94, new_R1192_U95, new_R1192_U96, new_R1192_U97,
    new_R1192_U98, new_R1192_U99, new_R1192_U100, new_R1192_U101,
    new_R1192_U102, new_R1192_U103, new_R1192_U104, new_R1192_U105,
    new_R1192_U106, new_R1192_U107, new_R1192_U108, new_R1192_U109,
    new_R1192_U110, new_R1192_U111, new_R1192_U112, new_R1192_U113,
    new_R1192_U114, new_R1192_U115, new_R1192_U116, new_R1192_U117,
    new_R1192_U118, new_R1192_U119, new_R1192_U120, new_R1192_U121,
    new_R1192_U122, new_R1192_U123, new_R1192_U124, new_R1192_U125,
    new_R1192_U126, new_R1192_U127, new_R1192_U128, new_R1192_U129,
    new_R1192_U130, new_R1192_U131, new_R1192_U132, new_R1192_U133,
    new_R1192_U134, new_R1192_U135, new_R1192_U136, new_R1192_U137,
    new_R1192_U138, new_R1192_U139, new_R1192_U140, new_R1192_U141,
    new_R1192_U142, new_R1192_U143, new_R1192_U144, new_R1192_U145,
    new_R1192_U146, new_R1192_U147, new_R1192_U148, new_R1192_U149,
    new_R1192_U150, new_R1192_U151, new_R1192_U152, new_R1192_U153,
    new_R1192_U154, new_R1192_U155, new_R1192_U156, new_R1192_U157,
    new_R1192_U158, new_R1192_U159, new_R1192_U160, new_R1192_U161,
    new_R1192_U162, new_R1192_U163, new_R1192_U164, new_R1192_U165,
    new_R1192_U166, new_R1192_U167, new_R1192_U168, new_R1192_U169,
    new_R1192_U170, new_R1192_U171, new_R1192_U172, new_R1192_U173,
    new_R1192_U174, new_R1192_U175, new_R1192_U176, new_R1192_U177,
    new_R1192_U178, new_R1192_U179, new_R1192_U180, new_R1192_U181,
    new_R1192_U182, new_R1192_U183, new_R1192_U184, new_R1192_U185,
    new_R1192_U186, new_R1192_U187, new_R1192_U188, new_R1192_U189,
    new_R1192_U190, new_R1192_U191, new_R1192_U192, new_R1192_U193,
    new_R1192_U194, new_R1192_U195, new_R1192_U196, new_R1192_U197,
    new_R1192_U198, new_R1192_U199, new_R1192_U200, new_R1192_U201,
    new_R1192_U202, new_R1192_U203, new_R1192_U204, new_R1192_U205,
    new_R1192_U206, new_R1192_U207, new_R1192_U208, new_R1192_U209,
    new_R1192_U210, new_R1192_U211, new_R1192_U212, new_R1192_U213,
    new_R1192_U214, new_R1192_U215, new_R1192_U216, new_R1192_U217,
    new_R1192_U218, new_R1192_U219, new_R1192_U220, new_R1192_U221,
    new_R1192_U222, new_R1192_U223, new_R1192_U224, new_R1192_U225,
    new_R1192_U226, new_R1192_U227, new_R1192_U228, new_R1192_U229,
    new_R1192_U230, new_R1192_U231, new_R1192_U232, new_R1192_U233,
    new_R1192_U234, new_R1192_U235, new_R1192_U236, new_R1192_U237,
    new_R1192_U238, new_R1192_U239, new_R1192_U240, new_R1192_U241,
    new_R1192_U242, new_R1192_U243, new_R1192_U244, new_R1192_U245,
    new_R1192_U246, new_R1192_U247, new_R1192_U248, new_R1192_U249,
    new_R1192_U250, new_R1192_U251, new_R1192_U252, new_R1192_U253,
    new_R1192_U254, new_R1192_U255, new_R1192_U256, new_R1192_U257,
    new_R1192_U258, new_R1192_U259, new_R1192_U260, new_R1192_U261,
    new_R1192_U262, new_R1192_U263, new_R1192_U264, new_R1192_U265,
    new_R1192_U266, new_R1192_U267, new_R1192_U268, new_R1192_U269,
    new_R1192_U270, new_R1192_U271, new_R1192_U272, new_R1192_U273,
    new_R1192_U274, new_R1192_U275, new_R1192_U276, new_R1192_U277,
    new_R1192_U278, new_R1192_U279, new_R1192_U280, new_R1192_U281,
    new_R1192_U282, new_R1192_U283, new_R1192_U284, new_R1192_U285,
    new_R1192_U286, new_R1192_U287, new_R1192_U288, new_R1192_U289,
    new_R1192_U290, new_R1192_U291, new_R1192_U292, new_R1192_U293,
    new_R1192_U294, new_R1192_U295, new_R1192_U296, new_R1192_U297,
    new_R1192_U298, new_R1192_U299, new_R1192_U300, new_R1192_U301,
    new_R1192_U302, new_R1192_U303, new_R1192_U304, new_R1192_U305,
    new_R1192_U306, new_R1192_U307, new_R1192_U308, new_R1192_U309,
    new_R1192_U310, new_R1192_U311, new_R1192_U312, new_R1192_U313,
    new_R1192_U314, new_R1192_U315, new_R1192_U316, new_R1192_U317,
    new_R1192_U318, new_R1192_U319, new_R1192_U320, new_R1192_U321,
    new_R1192_U322, new_R1192_U323, new_R1192_U324, new_R1192_U325,
    new_R1192_U326, new_R1192_U327, new_R1192_U328, new_R1192_U329,
    new_R1192_U330, new_R1192_U331, new_R1192_U332, new_R1192_U333,
    new_R1192_U334, new_R1192_U335, new_R1192_U336, new_R1192_U337,
    new_R1192_U338, new_R1192_U339, new_R1192_U340, new_R1192_U341,
    new_R1192_U342, new_R1192_U343, new_R1192_U344, new_R1192_U345,
    new_R1192_U346, new_R1192_U347, new_R1192_U348, new_R1192_U349,
    new_R1192_U350, new_R1192_U351, new_R1192_U352, new_R1192_U353,
    new_R1192_U354, new_R1192_U355, new_R1192_U356, new_R1192_U357,
    new_R1192_U358, new_R1192_U359, new_R1192_U360, new_R1192_U361,
    new_R1192_U362, new_R1192_U363, new_R1192_U364, new_R1192_U365,
    new_R1192_U366, new_R1192_U367, new_R1192_U368, new_R1192_U369,
    new_R1192_U370, new_R1192_U371, new_R1192_U372, new_R1192_U373,
    new_R1192_U374, new_R1192_U375, new_R1192_U376, new_R1192_U377,
    new_R1192_U378, new_R1192_U379, new_R1192_U380, new_R1192_U381,
    new_R1192_U382, new_R1192_U383, new_R1192_U384, new_R1192_U385,
    new_R1192_U386, new_R1192_U387, new_R1192_U388, new_R1192_U389,
    new_R1192_U390, new_R1192_U391, new_R1192_U392, new_R1192_U393,
    new_R1192_U394, new_R1192_U395, new_R1192_U396, new_R1192_U397,
    new_R1192_U398, new_R1192_U399, new_R1192_U400, new_R1192_U401,
    new_R1192_U402, new_R1192_U403, new_R1192_U404, new_R1192_U405,
    new_R1192_U406, new_R1192_U407, new_R1192_U408, new_R1192_U409,
    new_R1192_U410, new_R1192_U411, new_R1192_U412, new_R1192_U413,
    new_R1192_U414, new_R1192_U415, new_R1192_U416, new_R1192_U417,
    new_R1192_U418, new_R1192_U419, new_R1192_U420, new_R1192_U421,
    new_R1192_U422, new_R1192_U423, new_R1192_U424, new_R1192_U425,
    new_R1192_U426, new_R1192_U427, new_R1192_U428, new_R1192_U429,
    new_R1192_U430, new_R1192_U431, new_R1192_U432, new_R1192_U433,
    new_R1192_U434, new_R1192_U435, new_R1192_U436, new_R1192_U437,
    new_R1192_U438, new_R1192_U439, new_R1192_U440, new_R1192_U441,
    new_R1192_U442, new_R1192_U443, new_R1192_U444, new_R1192_U445,
    new_R1192_U446, new_R1192_U447, new_R1192_U448, new_R1192_U449,
    new_R1192_U450, new_R1192_U451, new_R1192_U452, new_R1192_U453,
    new_R1192_U454, new_R1192_U455, new_R1192_U456, new_R1192_U457,
    new_R1192_U458, new_R1192_U459, new_R1192_U460, new_R1192_U461,
    new_R1192_U462, new_R1192_U463, new_R1192_U464, new_R1192_U465,
    new_R1192_U466, new_R1192_U467, new_R1192_U468, new_R1192_U469,
    new_R1192_U470, new_R1192_U471, new_R1192_U472, new_R1192_U473,
    new_R1192_U474, new_R1192_U475, new_R1192_U476, new_R1192_U477,
    new_R1192_U478, new_R1192_U479, new_R1192_U480, new_R1192_U481,
    new_R1192_U482, new_R1192_U483, new_R1192_U484, new_R1192_U485,
    new_R1192_U486, new_R1192_U487, new_R1192_U488, new_R1192_U489,
    new_R1192_U490, new_R1192_U491, new_R1192_U492, new_R1192_U493,
    new_R1192_U494, new_R1192_U495, new_R1192_U496, new_R1192_U497,
    new_R1192_U498, new_R1192_U499, new_R1192_U500, new_R1192_U501,
    new_R1192_U502, new_R1192_U503, new_R1192_U504, new_R1192_U505,
    new_R1192_U506, new_R1192_U507, new_R1192_U508, new_R1192_U509,
    new_R1192_U510, new_R1192_U511, new_R1192_U512, new_R1192_U513,
    new_R1192_U514, new_R1192_U515, new_R1192_U516, new_R1192_U517,
    new_R1192_U518, new_R1192_U519, new_R1192_U520, new_R1347_U6,
    new_R1347_U7, new_R1347_U8, new_R1347_U9, new_R1347_U10, new_R1347_U11,
    new_R1347_U12, new_R1347_U13, new_R1347_U14, new_R1347_U15,
    new_R1347_U16, new_R1347_U17, new_R1347_U18, new_R1347_U19,
    new_R1347_U20, new_R1347_U21, new_R1347_U22, new_R1347_U23,
    new_R1347_U24, new_R1347_U25, new_R1347_U26, new_R1347_U27,
    new_R1347_U28, new_R1347_U29, new_R1347_U30, new_R1347_U31,
    new_R1347_U32, new_R1347_U33, new_R1347_U34, new_R1347_U35,
    new_R1347_U36, new_R1347_U37, new_R1347_U38, new_R1347_U39,
    new_R1347_U40, new_R1347_U41, new_R1347_U42, new_R1347_U43,
    new_R1347_U44, new_R1347_U45, new_R1347_U46, new_R1347_U47,
    new_R1347_U48, new_R1347_U49, new_R1347_U50, new_R1347_U51,
    new_R1347_U52, new_R1347_U53, new_R1347_U54, new_R1347_U55,
    new_R1347_U56, new_R1347_U57, new_R1347_U58, new_R1347_U59,
    new_R1347_U60, new_R1347_U61, new_R1347_U62, new_R1347_U63,
    new_R1347_U64, new_R1347_U65, new_R1347_U66, new_R1347_U67,
    new_R1347_U68, new_R1347_U69, new_R1347_U70, new_R1347_U71,
    new_R1347_U72, new_R1347_U73, new_R1347_U74, new_R1347_U75,
    new_R1347_U76, new_R1347_U77, new_R1347_U78, new_R1347_U79,
    new_R1347_U80, new_R1347_U81, new_R1347_U82, new_R1347_U83,
    new_R1347_U84, new_R1347_U85, new_R1347_U86, new_R1347_U87,
    new_R1347_U88, new_R1347_U89, new_R1347_U90, new_R1347_U91,
    new_R1347_U92, new_R1347_U93, new_R1347_U94, new_R1347_U95,
    new_R1347_U96, new_R1347_U97, new_R1347_U98, new_R1347_U99,
    new_R1347_U100, new_R1347_U101, new_R1347_U102, new_R1347_U103,
    new_R1347_U104, new_R1347_U105, new_R1347_U106, new_R1347_U107,
    new_R1347_U108, new_R1347_U109, new_R1347_U110, new_R1347_U111,
    new_R1347_U112, new_R1347_U113, new_R1347_U114, new_R1347_U115,
    new_R1347_U116, new_R1347_U117, new_R1347_U118, new_R1347_U119,
    new_R1347_U120, new_R1347_U121, new_R1347_U122, new_R1347_U123,
    new_R1347_U124, new_R1347_U125, new_R1347_U126, new_R1347_U127,
    new_R1347_U128, new_R1347_U129, new_R1347_U130, new_R1347_U131,
    new_R1347_U132, new_R1347_U133, new_R1347_U134, new_R1347_U135,
    new_R1347_U136, new_R1347_U137, new_R1347_U138, new_R1347_U139,
    new_R1347_U140, new_R1347_U141, new_R1347_U142, new_R1347_U143,
    new_R1347_U144, new_R1347_U145, new_R1347_U146, new_R1347_U147,
    new_R1347_U148, new_R1347_U149, new_R1347_U150, new_R1347_U151,
    new_R1347_U152, new_R1347_U153, new_R1347_U154, new_R1347_U155,
    new_R1347_U156, new_R1347_U157, new_R1347_U158, new_R1347_U159,
    new_R1347_U160, new_R1347_U161, new_R1347_U162, new_R1347_U163,
    new_R1347_U164, new_R1347_U165, new_R1347_U166, new_R1347_U167,
    new_R1347_U168, new_R1347_U169, new_R1347_U170, new_R1347_U171,
    new_R1347_U172, new_R1347_U173, new_R1347_U174, new_R1347_U175,
    new_R1347_U176, new_R1347_U177, new_R1347_U178, new_R1347_U179,
    new_R1347_U180, new_R1347_U181, new_R1347_U182, new_R1347_U183,
    new_R1347_U184, new_R1347_U185, new_R1347_U186, new_R1347_U187,
    new_R1347_U188, new_R1347_U189, new_R1347_U190, new_R1347_U191,
    new_R1347_U192, new_R1347_U193, new_R1347_U194, new_R1347_U195,
    new_R1347_U196, new_R1347_U197, new_R1347_U198, new_R1347_U199,
    new_R1347_U200, new_R1347_U201, new_R1347_U202, new_R1347_U203,
    new_R1347_U204, new_R1347_U205, new_R1347_U206, new_R1347_U207,
    new_R1347_U208, new_R1347_U209, new_R1347_U210, new_R1347_U211,
    new_R1347_U212, new_R1171_U4, new_R1171_U5, new_R1171_U6, new_R1171_U7,
    new_R1171_U8, new_R1171_U9, new_R1171_U10, new_R1171_U11,
    new_R1171_U12, new_R1171_U13, new_R1171_U14, new_R1171_U15,
    new_R1171_U16, new_R1171_U17, new_R1171_U18, new_R1171_U19,
    new_R1171_U20, new_R1171_U21, new_R1171_U22, new_R1171_U23,
    new_R1171_U24, new_R1171_U25, new_R1171_U26, new_R1171_U27,
    new_R1171_U28, new_R1171_U29, new_R1171_U30, new_R1171_U31,
    new_R1171_U32, new_R1171_U33, new_R1171_U34, new_R1171_U35,
    new_R1171_U36, new_R1171_U37, new_R1171_U38, new_R1171_U39,
    new_R1171_U40, new_R1171_U41, new_R1171_U42, new_R1171_U43,
    new_R1171_U44, new_R1171_U45, new_R1171_U46, new_R1171_U47,
    new_R1171_U48, new_R1171_U49, new_R1171_U50, new_R1171_U51,
    new_R1171_U52, new_R1171_U53, new_R1171_U54, new_R1171_U55,
    new_R1171_U56, new_R1171_U57, new_R1171_U58, new_R1171_U59,
    new_R1171_U60, new_R1171_U61, new_R1171_U62, new_R1171_U63,
    new_R1171_U64, new_R1171_U65, new_R1171_U66, new_R1171_U67,
    new_R1171_U68, new_R1171_U69, new_R1171_U70, new_R1171_U71,
    new_R1171_U72, new_R1171_U73, new_R1171_U74, new_R1171_U75,
    new_R1171_U76, new_R1171_U77, new_R1171_U78, new_R1171_U79,
    new_R1171_U80, new_R1171_U81, new_R1171_U82, new_R1171_U83,
    new_R1171_U84, new_R1171_U85, new_R1171_U86, new_R1171_U87,
    new_R1171_U88, new_R1171_U89, new_R1171_U90, new_R1171_U91,
    new_R1171_U92, new_R1171_U93, new_R1171_U94, new_R1171_U95,
    new_R1171_U96, new_R1171_U97, new_R1171_U98, new_R1171_U99,
    new_R1171_U100, new_R1171_U101, new_R1171_U102, new_R1171_U103,
    new_R1171_U104, new_R1171_U105, new_R1171_U106, new_R1171_U107,
    new_R1171_U108, new_R1171_U109, new_R1171_U110, new_R1171_U111,
    new_R1171_U112, new_R1171_U113, new_R1171_U114, new_R1171_U115,
    new_R1171_U116, new_R1171_U117, new_R1171_U118, new_R1171_U119,
    new_R1171_U120, new_R1171_U121, new_R1171_U122, new_R1171_U123,
    new_R1171_U124, new_R1171_U125, new_R1171_U126, new_R1171_U127,
    new_R1171_U128, new_R1171_U129, new_R1171_U130, new_R1171_U131,
    new_R1171_U132, new_R1171_U133, new_R1171_U134, new_R1171_U135,
    new_R1171_U136, new_R1171_U137, new_R1171_U138, new_R1171_U139,
    new_R1171_U140, new_R1171_U141, new_R1171_U142, new_R1171_U143,
    new_R1171_U144, new_R1171_U145, new_R1171_U146, new_R1171_U147,
    new_R1171_U148, new_R1171_U149, new_R1171_U150, new_R1171_U151,
    new_R1171_U152, new_R1171_U153, new_R1171_U154, new_R1171_U155,
    new_R1171_U156, new_R1171_U157, new_R1171_U158, new_R1171_U159,
    new_R1171_U160, new_R1171_U161, new_R1171_U162, new_R1171_U163,
    new_R1171_U164, new_R1171_U165, new_R1171_U166, new_R1171_U167,
    new_R1171_U168, new_R1171_U169, new_R1171_U170, new_R1171_U171,
    new_R1171_U172, new_R1171_U173, new_R1171_U174, new_R1171_U175,
    new_R1171_U176, new_R1171_U177, new_R1171_U178, new_R1171_U179,
    new_R1171_U180, new_R1171_U181, new_R1171_U182, new_R1171_U183,
    new_R1171_U184, new_R1171_U185, new_R1171_U186, new_R1171_U187,
    new_R1171_U188, new_R1171_U189, new_R1171_U190, new_R1171_U191,
    new_R1171_U192, new_R1171_U193, new_R1171_U194, new_R1171_U195,
    new_R1171_U196, new_R1171_U197, new_R1171_U198, new_R1171_U199,
    new_R1171_U200, new_R1171_U201, new_R1171_U202, new_R1171_U203,
    new_R1171_U204, new_R1171_U205, new_R1171_U206, new_R1171_U207,
    new_R1171_U208, new_R1171_U209, new_R1171_U210, new_R1171_U211,
    new_R1171_U212, new_R1171_U213, new_R1171_U214, new_R1171_U215,
    new_R1171_U216, new_R1171_U217, new_R1171_U218, new_R1171_U219,
    new_R1171_U220, new_R1171_U221, new_R1171_U222, new_R1171_U223,
    new_R1171_U224, new_R1171_U225, new_R1171_U226, new_R1171_U227,
    new_R1171_U228, new_R1171_U229, new_R1171_U230, new_R1171_U231,
    new_R1171_U232, new_R1171_U233, new_R1171_U234, new_R1171_U235,
    new_R1171_U236, new_R1171_U237, new_R1171_U238, new_R1171_U239,
    new_R1171_U240, new_R1171_U241, new_R1171_U242, new_R1171_U243,
    new_R1171_U244, new_R1171_U245, new_R1171_U246, new_R1171_U247,
    new_R1171_U248, new_R1171_U249, new_R1171_U250, new_R1171_U251,
    new_R1171_U252, new_R1171_U253, new_R1171_U254, new_R1171_U255,
    new_R1171_U256, new_R1171_U257, new_R1171_U258, new_R1171_U259,
    new_R1171_U260, new_R1171_U261, new_R1171_U262, new_R1171_U263,
    new_R1171_U264, new_R1171_U265, new_R1171_U266, new_R1171_U267,
    new_R1171_U268, new_R1171_U269, new_R1171_U270, new_R1171_U271,
    new_R1171_U272, new_R1171_U273, new_R1171_U274, new_R1171_U275,
    new_R1171_U276, new_R1171_U277, new_R1171_U278, new_R1171_U279,
    new_R1171_U280, new_R1171_U281, new_R1171_U282, new_R1171_U283,
    new_R1171_U284, new_R1171_U285, new_R1171_U286, new_R1171_U287,
    new_R1171_U288, new_R1171_U289, new_R1171_U290, new_R1171_U291,
    new_R1171_U292, new_R1171_U293, new_R1171_U294, new_R1171_U295,
    new_R1171_U296, new_R1171_U297, new_R1171_U298, new_R1171_U299,
    new_R1171_U300, new_R1171_U301, new_R1171_U302, new_R1171_U303,
    new_R1171_U304, new_R1171_U305, new_R1171_U306, new_R1171_U307,
    new_R1171_U308, new_R1171_U309, new_R1171_U310, new_R1171_U311,
    new_R1171_U312, new_R1171_U313, new_R1171_U314, new_R1171_U315,
    new_R1171_U316, new_R1171_U317, new_R1171_U318, new_R1171_U319,
    new_R1171_U320, new_R1171_U321, new_R1171_U322, new_R1171_U323,
    new_R1171_U324, new_R1171_U325, new_R1171_U326, new_R1171_U327,
    new_R1171_U328, new_R1171_U329, new_R1171_U330, new_R1171_U331,
    new_R1171_U332, new_R1171_U333, new_R1171_U334, new_R1171_U335,
    new_R1171_U336, new_R1171_U337, new_R1171_U338, new_R1171_U339,
    new_R1171_U340, new_R1171_U341, new_R1171_U342, new_R1171_U343,
    new_R1171_U344, new_R1171_U345, new_R1171_U346, new_R1171_U347,
    new_R1171_U348, new_R1171_U349, new_R1171_U350, new_R1171_U351,
    new_R1171_U352, new_R1171_U353, new_R1171_U354, new_R1171_U355,
    new_R1171_U356, new_R1171_U357, new_R1171_U358, new_R1171_U359,
    new_R1171_U360, new_R1171_U361, new_R1171_U362, new_R1171_U363,
    new_R1171_U364, new_R1171_U365, new_R1171_U366, new_R1171_U367,
    new_R1171_U368, new_R1171_U369, new_R1171_U370, new_R1171_U371,
    new_R1171_U372, new_R1171_U373, new_R1171_U374, new_R1171_U375,
    new_R1171_U376, new_R1171_U377, new_R1171_U378, new_R1171_U379,
    new_R1171_U380, new_R1171_U381, new_R1171_U382, new_R1171_U383,
    new_R1171_U384, new_R1171_U385, new_R1171_U386, new_R1171_U387,
    new_R1171_U388, new_R1171_U389, new_R1171_U390, new_R1171_U391,
    new_R1171_U392, new_R1171_U393, new_R1171_U394, new_R1171_U395,
    new_R1171_U396, new_R1171_U397, new_R1171_U398, new_R1171_U399,
    new_R1171_U400, new_R1171_U401, new_R1171_U402, new_R1171_U403,
    new_R1171_U404, new_R1171_U405, new_R1171_U406, new_R1171_U407,
    new_R1171_U408, new_R1171_U409, new_R1171_U410, new_R1171_U411,
    new_R1171_U412, new_R1171_U413, new_R1171_U414, new_R1171_U415,
    new_R1171_U416, new_R1171_U417, new_R1171_U418, new_R1171_U419,
    new_R1171_U420, new_R1171_U421, new_R1171_U422, new_R1171_U423,
    new_R1171_U424, new_R1171_U425, new_R1171_U426, new_R1171_U427,
    new_R1171_U428, new_R1171_U429, new_R1171_U430, new_R1171_U431,
    new_R1171_U432, new_R1171_U433, new_R1171_U434, new_R1171_U435,
    new_R1171_U436, new_R1171_U437, new_R1171_U438, new_R1171_U439,
    new_R1171_U440, new_R1171_U441, new_R1171_U442, new_R1171_U443,
    new_R1171_U444, new_R1171_U445, new_R1171_U446, new_R1171_U447,
    new_R1171_U448, new_R1171_U449, new_R1171_U450, new_R1171_U451,
    new_R1171_U452, new_R1171_U453, new_R1171_U454, new_R1171_U455,
    new_R1171_U456, new_R1171_U457, new_R1171_U458, new_R1171_U459,
    new_R1171_U460, new_R1171_U461, new_R1171_U462, new_R1171_U463,
    new_R1171_U464, new_R1171_U465, new_R1171_U466, new_R1171_U467,
    new_R1171_U468, new_R1171_U469, new_R1171_U470, new_R1171_U471,
    new_R1171_U472, new_R1171_U473, new_R1171_U474, new_R1171_U475,
    new_R1171_U476, new_R1171_U477, new_R1171_U478, new_R1171_U479,
    new_R1171_U480, new_R1171_U481, new_R1171_U482, new_R1171_U483,
    new_R1171_U484, new_R1171_U485, new_R1171_U486, new_R1171_U487,
    new_R1171_U488, new_R1171_U489, new_R1171_U490, new_R1171_U491,
    new_R1171_U492, new_R1171_U493, new_R1171_U494, new_R1171_U495,
    new_R1171_U496, new_R1171_U497, new_R1171_U498, new_R1171_U499,
    new_R1171_U500, new_R1171_U501, new_R1171_U502, new_R1171_U503,
    new_R1171_U504, new_R1171_U505, new_R1171_U506, new_R1171_U507,
    new_R1171_U508, new_R1171_U509, new_R1171_U510, new_R1171_U511,
    new_R1171_U512, new_R1171_U513, new_R1171_U514, new_R1171_U515,
    new_R1171_U516, new_R1171_U517, new_R1171_U518, new_R1171_U519,
    new_R1171_U520, new_R1171_U521, new_R1171_U522, new_R1171_U523,
    new_R1171_U524, new_R1171_U525, new_R1171_U526, new_R1171_U527,
    new_R1171_U528, new_R1171_U529, new_R1171_U530, new_R1171_U531,
    new_R1138_U4, new_R1138_U5, new_R1138_U6, new_R1138_U7, new_R1138_U8,
    new_R1138_U9, new_R1138_U10, new_R1138_U11, new_R1138_U12,
    new_R1138_U13, new_R1138_U14, new_R1138_U15, new_R1138_U16,
    new_R1138_U17, new_R1138_U18, new_R1138_U19, new_R1138_U20,
    new_R1138_U21, new_R1138_U22, new_R1138_U23, new_R1138_U24,
    new_R1138_U25, new_R1138_U26, new_R1138_U27, new_R1138_U28,
    new_R1138_U29, new_R1138_U30, new_R1138_U31, new_R1138_U32,
    new_R1138_U33, new_R1138_U34, new_R1138_U35, new_R1138_U36,
    new_R1138_U37, new_R1138_U38, new_R1138_U39, new_R1138_U40,
    new_R1138_U41, new_R1138_U42, new_R1138_U43, new_R1138_U44,
    new_R1138_U45, new_R1138_U46, new_R1138_U47, new_R1138_U48,
    new_R1138_U49, new_R1138_U50, new_R1138_U51, new_R1138_U52,
    new_R1138_U53, new_R1138_U54, new_R1138_U55, new_R1138_U56,
    new_R1138_U57, new_R1138_U58, new_R1138_U59, new_R1138_U60,
    new_R1138_U61, new_R1138_U62, new_R1138_U63, new_R1138_U64,
    new_R1138_U65, new_R1138_U66, new_R1138_U67, new_R1138_U68,
    new_R1138_U69, new_R1138_U70, new_R1138_U71, new_R1138_U72,
    new_R1138_U73, new_R1138_U74, new_R1138_U75, new_R1138_U76,
    new_R1138_U77, new_R1138_U78, new_R1138_U79, new_R1138_U80,
    new_R1138_U81, new_R1138_U82, new_R1138_U83, new_R1138_U84,
    new_R1138_U85, new_R1138_U86, new_R1138_U87, new_R1138_U88,
    new_R1138_U89, new_R1138_U90, new_R1138_U91, new_R1138_U92,
    new_R1138_U93, new_R1138_U94, new_R1138_U95, new_R1138_U96,
    new_R1138_U97, new_R1138_U98, new_R1138_U99, new_R1138_U100,
    new_R1138_U101, new_R1138_U102, new_R1138_U103, new_R1138_U104,
    new_R1138_U105, new_R1138_U106, new_R1138_U107, new_R1138_U108,
    new_R1138_U109, new_R1138_U110, new_R1138_U111, new_R1138_U112,
    new_R1138_U113, new_R1138_U114, new_R1138_U115, new_R1138_U116,
    new_R1138_U117, new_R1138_U118, new_R1138_U119, new_R1138_U120,
    new_R1138_U121, new_R1138_U122, new_R1138_U123, new_R1138_U124,
    new_R1138_U125, new_R1138_U126, new_R1138_U127, new_R1138_U128,
    new_R1138_U129, new_R1138_U130, new_R1138_U131, new_R1138_U132,
    new_R1138_U133, new_R1138_U134, new_R1138_U135, new_R1138_U136,
    new_R1138_U137, new_R1138_U138, new_R1138_U139, new_R1138_U140,
    new_R1138_U141, new_R1138_U142, new_R1138_U143, new_R1138_U144,
    new_R1138_U145, new_R1138_U146, new_R1138_U147, new_R1138_U148,
    new_R1138_U149, new_R1138_U150, new_R1138_U151, new_R1138_U152,
    new_R1138_U153, new_R1138_U154, new_R1138_U155, new_R1138_U156,
    new_R1138_U157, new_R1138_U158, new_R1138_U159, new_R1138_U160,
    new_R1138_U161, new_R1138_U162, new_R1138_U163, new_R1138_U164,
    new_R1138_U165, new_R1138_U166, new_R1138_U167, new_R1138_U168,
    new_R1138_U169, new_R1138_U170, new_R1138_U171, new_R1138_U172,
    new_R1138_U173, new_R1138_U174, new_R1138_U175, new_R1138_U176,
    new_R1138_U177, new_R1138_U178, new_R1138_U179, new_R1138_U180,
    new_R1138_U181, new_R1138_U182, new_R1138_U183, new_R1138_U184,
    new_R1138_U185, new_R1138_U186, new_R1138_U187, new_R1138_U188,
    new_R1138_U189, new_R1138_U190, new_R1138_U191, new_R1138_U192,
    new_R1138_U193, new_R1138_U194, new_R1138_U195, new_R1138_U196,
    new_R1138_U197, new_R1138_U198, new_R1138_U199, new_R1138_U200,
    new_R1138_U201, new_R1138_U202, new_R1138_U203, new_R1138_U204,
    new_R1138_U205, new_R1138_U206, new_R1138_U207, new_R1138_U208,
    new_R1138_U209, new_R1138_U210, new_R1138_U211, new_R1138_U212,
    new_R1138_U213, new_R1138_U214, new_R1138_U215, new_R1138_U216,
    new_R1138_U217, new_R1138_U218, new_R1138_U219, new_R1138_U220,
    new_R1138_U221, new_R1138_U222, new_R1138_U223, new_R1138_U224,
    new_R1138_U225, new_R1138_U226, new_R1138_U227, new_R1138_U228,
    new_R1138_U229, new_R1138_U230, new_R1138_U231, new_R1138_U232,
    new_R1138_U233, new_R1138_U234, new_R1138_U235, new_R1138_U236,
    new_R1138_U237, new_R1138_U238, new_R1138_U239, new_R1138_U240,
    new_R1138_U241, new_R1138_U242, new_R1138_U243, new_R1138_U244,
    new_R1138_U245, new_R1138_U246, new_R1138_U247, new_R1138_U248,
    new_R1138_U249, new_R1138_U250, new_R1138_U251, new_R1138_U252,
    new_R1138_U253, new_R1138_U254, new_R1138_U255, new_R1138_U256,
    new_R1138_U257, new_R1138_U258, new_R1138_U259, new_R1138_U260,
    new_R1138_U261, new_R1138_U262, new_R1138_U263, new_R1138_U264,
    new_R1138_U265, new_R1138_U266, new_R1138_U267, new_R1138_U268,
    new_R1138_U269, new_R1138_U270, new_R1138_U271, new_R1138_U272,
    new_R1138_U273, new_R1138_U274, new_R1138_U275, new_R1138_U276,
    new_R1138_U277, new_R1138_U278, new_R1138_U279, new_R1138_U280,
    new_R1138_U281, new_R1138_U282, new_R1138_U283, new_R1138_U284,
    new_R1138_U285, new_R1138_U286, new_R1138_U287, new_R1138_U288,
    new_R1138_U289, new_R1138_U290, new_R1138_U291, new_R1138_U292,
    new_R1138_U293, new_R1138_U294, new_R1138_U295, new_R1138_U296,
    new_R1138_U297, new_R1138_U298, new_R1138_U299, new_R1138_U300,
    new_R1138_U301, new_R1138_U302, new_R1138_U303, new_R1138_U304,
    new_R1138_U305, new_R1138_U306, new_R1138_U307, new_R1138_U308,
    new_R1138_U309, new_R1138_U310, new_R1138_U311, new_R1138_U312,
    new_R1138_U313, new_R1138_U314, new_R1138_U315, new_R1138_U316,
    new_R1138_U317, new_R1138_U318, new_R1138_U319, new_R1138_U320,
    new_R1138_U321, new_R1138_U322, new_R1138_U323, new_R1138_U324,
    new_R1138_U325, new_R1138_U326, new_R1138_U327, new_R1138_U328,
    new_R1138_U329, new_R1138_U330, new_R1138_U331, new_R1138_U332,
    new_R1138_U333, new_R1138_U334, new_R1138_U335, new_R1138_U336,
    new_R1138_U337, new_R1138_U338, new_R1138_U339, new_R1138_U340,
    new_R1138_U341, new_R1138_U342, new_R1138_U343, new_R1138_U344,
    new_R1138_U345, new_R1138_U346, new_R1138_U347, new_R1138_U348,
    new_R1138_U349, new_R1138_U350, new_R1138_U351, new_R1138_U352,
    new_R1138_U353, new_R1138_U354, new_R1138_U355, new_R1138_U356,
    new_R1138_U357, new_R1138_U358, new_R1138_U359, new_R1138_U360,
    new_R1138_U361, new_R1138_U362, new_R1138_U363, new_R1138_U364,
    new_R1138_U365, new_R1138_U366, new_R1138_U367, new_R1138_U368,
    new_R1138_U369, new_R1138_U370, new_R1138_U371, new_R1138_U372,
    new_R1138_U373, new_R1138_U374, new_R1138_U375, new_R1138_U376,
    new_R1138_U377, new_R1138_U378, new_R1138_U379, new_R1138_U380,
    new_R1138_U381, new_R1138_U382, new_R1138_U383, new_R1138_U384,
    new_R1138_U385, new_R1138_U386, new_R1138_U387, new_R1138_U388,
    new_R1138_U389, new_R1138_U390, new_R1138_U391, new_R1138_U392,
    new_R1138_U393, new_R1138_U394, new_R1138_U395, new_R1138_U396,
    new_R1138_U397, new_R1138_U398, new_R1138_U399, new_R1138_U400,
    new_R1138_U401, new_R1138_U402, new_R1138_U403, new_R1138_U404,
    new_R1138_U405, new_R1138_U406, new_R1138_U407, new_R1138_U408,
    new_R1138_U409, new_R1138_U410, new_R1138_U411, new_R1138_U412,
    new_R1138_U413, new_R1138_U414, new_R1138_U415, new_R1138_U416,
    new_R1138_U417, new_R1138_U418, new_R1138_U419, new_R1138_U420,
    new_R1138_U421, new_R1138_U422, new_R1138_U423, new_R1138_U424,
    new_R1138_U425, new_R1138_U426, new_R1138_U427, new_R1138_U428,
    new_R1138_U429, new_R1138_U430, new_R1138_U431, new_R1138_U432,
    new_R1138_U433, new_R1138_U434, new_R1138_U435, new_R1138_U436,
    new_R1138_U437, new_R1138_U438, new_R1138_U439, new_R1138_U440,
    new_R1138_U441, new_R1138_U442, new_R1138_U443, new_R1138_U444,
    new_R1138_U445, new_R1138_U446, new_R1138_U447, new_R1138_U448,
    new_R1138_U449, new_R1138_U450, new_R1138_U451, new_R1138_U452,
    new_R1138_U453, new_R1138_U454, new_R1138_U455, new_R1138_U456,
    new_R1138_U457, new_R1138_U458, new_R1138_U459, new_R1138_U460,
    new_R1138_U461, new_R1138_U462, new_R1138_U463, new_R1138_U464,
    new_R1138_U465, new_R1138_U466, new_R1138_U467, new_R1138_U468,
    new_R1138_U469, new_R1138_U470, new_R1138_U471, new_R1138_U472,
    new_R1138_U473, new_R1138_U474, new_R1138_U475, new_R1138_U476,
    new_R1138_U477, new_R1138_U478, new_R1138_U479, new_R1138_U480,
    new_R1138_U481, new_R1138_U482, new_R1138_U483, new_R1138_U484,
    new_R1138_U485, new_R1138_U486, new_R1138_U487, new_R1138_U488,
    new_R1138_U489, new_R1138_U490, new_R1138_U491, new_R1138_U492,
    new_R1138_U493, new_R1138_U494, new_R1138_U495, new_R1138_U496,
    new_R1138_U497, new_R1138_U498, new_R1138_U499, new_R1138_U500,
    new_R1138_U501, new_R1138_U502, new_R1138_U503, new_R1138_U504,
    new_R1138_U505, new_R1138_U506, new_R1138_U507, new_R1138_U508,
    new_R1138_U509, new_R1138_U510, new_R1138_U511, new_R1138_U512,
    new_R1138_U513, new_R1138_U514, new_R1138_U515, new_R1138_U516,
    new_R1138_U517, new_R1138_U518, new_R1138_U519, new_R1138_U520,
    new_R1138_U521, new_R1138_U522, new_R1138_U523, new_R1138_U524,
    new_R1138_U525, new_R1138_U526, new_R1138_U527, new_R1138_U528,
    new_R1138_U529, new_R1138_U530, new_R1138_U531, new_R1222_U4,
    new_R1222_U5, new_R1222_U6, new_R1222_U7, new_R1222_U8, new_R1222_U9,
    new_R1222_U10, new_R1222_U11, new_R1222_U12, new_R1222_U13,
    new_R1222_U14, new_R1222_U15, new_R1222_U16, new_R1222_U17,
    new_R1222_U18, new_R1222_U19, new_R1222_U20, new_R1222_U21,
    new_R1222_U22, new_R1222_U23, new_R1222_U24, new_R1222_U25,
    new_R1222_U26, new_R1222_U27, new_R1222_U28, new_R1222_U29,
    new_R1222_U30, new_R1222_U31, new_R1222_U32, new_R1222_U33,
    new_R1222_U34, new_R1222_U35, new_R1222_U36, new_R1222_U37,
    new_R1222_U38, new_R1222_U39, new_R1222_U40, new_R1222_U41,
    new_R1222_U42, new_R1222_U43, new_R1222_U44, new_R1222_U45,
    new_R1222_U46, new_R1222_U47, new_R1222_U48, new_R1222_U49,
    new_R1222_U50, new_R1222_U51, new_R1222_U52, new_R1222_U53,
    new_R1222_U54, new_R1222_U55, new_R1222_U56, new_R1222_U57,
    new_R1222_U58, new_R1222_U59, new_R1222_U60, new_R1222_U61,
    new_R1222_U62, new_R1222_U63, new_R1222_U64, new_R1222_U65,
    new_R1222_U66, new_R1222_U67, new_R1222_U68, new_R1222_U69,
    new_R1222_U70, new_R1222_U71, new_R1222_U72, new_R1222_U73,
    new_R1222_U74, new_R1222_U75, new_R1222_U76, new_R1222_U77,
    new_R1222_U78, new_R1222_U79, new_R1222_U80, new_R1222_U81,
    new_R1222_U82, new_R1222_U83, new_R1222_U84, new_R1222_U85,
    new_R1222_U86, new_R1222_U87, new_R1222_U88, new_R1222_U89,
    new_R1222_U90, new_R1222_U91, new_R1222_U92, new_R1222_U93,
    new_R1222_U94, new_R1222_U95, new_R1222_U96, new_R1222_U97,
    new_R1222_U98, new_R1222_U99, new_R1222_U100, new_R1222_U101,
    new_R1222_U102, new_R1222_U103, new_R1222_U104, new_R1222_U105,
    new_R1222_U106, new_R1222_U107, new_R1222_U108, new_R1222_U109,
    new_R1222_U110, new_R1222_U111, new_R1222_U112, new_R1222_U113,
    new_R1222_U114, new_R1222_U115, new_R1222_U116, new_R1222_U117,
    new_R1222_U118, new_R1222_U119, new_R1222_U120, new_R1222_U121,
    new_R1222_U122, new_R1222_U123, new_R1222_U124, new_R1222_U125,
    new_R1222_U126, new_R1222_U127, new_R1222_U128, new_R1222_U129,
    new_R1222_U130, new_R1222_U131, new_R1222_U132, new_R1222_U133,
    new_R1222_U134, new_R1222_U135, new_R1222_U136, new_R1222_U137,
    new_R1222_U138, new_R1222_U139, new_R1222_U140, new_R1222_U141,
    new_R1222_U142, new_R1222_U143, new_R1222_U144, new_R1222_U145,
    new_R1222_U146, new_R1222_U147, new_R1222_U148, new_R1222_U149,
    new_R1222_U150, new_R1222_U151, new_R1222_U152, new_R1222_U153,
    new_R1222_U154, new_R1222_U155, new_R1222_U156, new_R1222_U157,
    new_R1222_U158, new_R1222_U159, new_R1222_U160, new_R1222_U161,
    new_R1222_U162, new_R1222_U163, new_R1222_U164, new_R1222_U165,
    new_R1222_U166, new_R1222_U167, new_R1222_U168, new_R1222_U169,
    new_R1222_U170, new_R1222_U171, new_R1222_U172, new_R1222_U173,
    new_R1222_U174, new_R1222_U175, new_R1222_U176, new_R1222_U177,
    new_R1222_U178, new_R1222_U179, new_R1222_U180, new_R1222_U181,
    new_R1222_U182, new_R1222_U183, new_R1222_U184, new_R1222_U185,
    new_R1222_U186, new_R1222_U187, new_R1222_U188, new_R1222_U189,
    new_R1222_U190, new_R1222_U191, new_R1222_U192, new_R1222_U193,
    new_R1222_U194, new_R1222_U195, new_R1222_U196, new_R1222_U197,
    new_R1222_U198, new_R1222_U199, new_R1222_U200, new_R1222_U201,
    new_R1222_U202, new_R1222_U203, new_R1222_U204, new_R1222_U205,
    new_R1222_U206, new_R1222_U207, new_R1222_U208, new_R1222_U209,
    new_R1222_U210, new_R1222_U211, new_R1222_U212, new_R1222_U213,
    new_R1222_U214, new_R1222_U215, new_R1222_U216, new_R1222_U217,
    new_R1222_U218, new_R1222_U219, new_R1222_U220, new_R1222_U221,
    new_R1222_U222, new_R1222_U223, new_R1222_U224, new_R1222_U225,
    new_R1222_U226, new_R1222_U227, new_R1222_U228, new_R1222_U229,
    new_R1222_U230, new_R1222_U231, new_R1222_U232, new_R1222_U233,
    new_R1222_U234, new_R1222_U235, new_R1222_U236, new_R1222_U237,
    new_R1222_U238, new_R1222_U239, new_R1222_U240, new_R1222_U241,
    new_R1222_U242, new_R1222_U243, new_R1222_U244, new_R1222_U245,
    new_R1222_U246, new_R1222_U247, new_R1222_U248, new_R1222_U249,
    new_R1222_U250, new_R1222_U251, new_R1222_U252, new_R1222_U253,
    new_R1222_U254, new_R1222_U255, new_R1222_U256, new_R1222_U257,
    new_R1222_U258, new_R1222_U259, new_R1222_U260, new_R1222_U261,
    new_R1222_U262, new_R1222_U263, new_R1222_U264, new_R1222_U265,
    new_R1222_U266, new_R1222_U267, new_R1222_U268, new_R1222_U269,
    new_R1222_U270, new_R1222_U271, new_R1222_U272, new_R1222_U273,
    new_R1222_U274, new_R1222_U275, new_R1222_U276, new_R1222_U277,
    new_R1222_U278, new_R1222_U279, new_R1222_U280, new_R1222_U281,
    new_R1222_U282, new_R1222_U283, new_R1222_U284, new_R1222_U285,
    new_R1222_U286, new_R1222_U287, new_R1222_U288, new_R1222_U289,
    new_R1222_U290, new_R1222_U291, new_R1222_U292, new_R1222_U293,
    new_R1222_U294, new_R1222_U295, new_R1222_U296, new_R1222_U297,
    new_R1222_U298, new_R1222_U299, new_R1222_U300, new_R1222_U301,
    new_R1222_U302, new_R1222_U303, new_R1222_U304, new_R1222_U305,
    new_R1222_U306, new_R1222_U307, new_R1222_U308, new_R1222_U309,
    new_R1222_U310, new_R1222_U311, new_R1222_U312, new_R1222_U313,
    new_R1222_U314, new_R1222_U315, new_R1222_U316, new_R1222_U317,
    new_R1222_U318, new_R1222_U319, new_R1222_U320, new_R1222_U321,
    new_R1222_U322, new_R1222_U323, new_R1222_U324, new_R1222_U325,
    new_R1222_U326, new_R1222_U327, new_R1222_U328, new_R1222_U329,
    new_R1222_U330, new_R1222_U331, new_R1222_U332, new_R1222_U333,
    new_R1222_U334, new_R1222_U335, new_R1222_U336, new_R1222_U337,
    new_R1222_U338, new_R1222_U339, new_R1222_U340, new_R1222_U341,
    new_R1222_U342, new_R1222_U343, new_R1222_U344, new_R1222_U345,
    new_R1222_U346, new_R1222_U347, new_R1222_U348, new_R1222_U349,
    new_R1222_U350, new_R1222_U351, new_R1222_U352, new_R1222_U353,
    new_R1222_U354, new_R1222_U355, new_R1222_U356, new_R1222_U357,
    new_R1222_U358, new_R1222_U359, new_R1222_U360, new_R1222_U361,
    new_R1222_U362, new_R1222_U363, new_R1222_U364, new_R1222_U365,
    new_R1222_U366, new_R1222_U367, new_R1222_U368, new_R1222_U369,
    new_R1222_U370, new_R1222_U371, new_R1222_U372, new_R1222_U373,
    new_R1222_U374, new_R1222_U375, new_R1222_U376, new_R1222_U377,
    new_R1222_U378, new_R1222_U379, new_R1222_U380, new_R1222_U381,
    new_R1222_U382, new_R1222_U383, new_R1222_U384, new_R1222_U385,
    new_R1222_U386, new_R1222_U387, new_R1222_U388, new_R1222_U389,
    new_R1222_U390, new_R1222_U391, new_R1222_U392, new_R1222_U393,
    new_R1222_U394, new_R1222_U395, new_R1222_U396, new_R1222_U397,
    new_R1222_U398, new_R1222_U399, new_R1222_U400, new_R1222_U401,
    new_R1222_U402, new_R1222_U403, new_R1222_U404, new_R1222_U405,
    new_R1222_U406, new_R1222_U407, new_R1222_U408, new_R1222_U409,
    new_R1222_U410, new_R1222_U411, new_R1222_U412, new_R1222_U413,
    new_R1222_U414, new_R1222_U415, new_R1222_U416, new_R1222_U417,
    new_R1222_U418, new_R1222_U419, new_R1222_U420, new_R1222_U421,
    new_R1222_U422, new_R1222_U423, new_R1222_U424, new_R1222_U425,
    new_R1222_U426, new_R1222_U427, new_R1222_U428, new_R1222_U429,
    new_R1222_U430, new_R1222_U431, new_R1222_U432, new_R1222_U433,
    new_R1222_U434, new_R1222_U435, new_R1222_U436, new_R1222_U437,
    new_R1222_U438, new_R1222_U439, new_R1222_U440, new_R1222_U441,
    new_R1222_U442, new_R1222_U443, new_R1222_U444, new_R1222_U445,
    new_R1222_U446, new_R1222_U447, new_R1222_U448, new_R1222_U449,
    new_R1222_U450, new_R1222_U451, new_R1222_U452, new_R1222_U453,
    new_R1222_U454, new_R1222_U455, new_R1222_U456, new_R1222_U457,
    new_R1222_U458, new_R1222_U459, new_R1222_U460, new_R1222_U461,
    new_R1222_U462, new_R1222_U463, new_R1222_U464, new_R1222_U465,
    new_R1222_U466, new_R1222_U467, new_R1222_U468, new_R1222_U469,
    new_R1222_U470, new_R1222_U471, new_R1222_U472, new_R1222_U473,
    new_R1222_U474, new_R1222_U475, new_R1222_U476, new_R1222_U477,
    new_R1222_U478, new_R1222_U479, new_R1222_U480, new_R1222_U481,
    new_R1222_U482, new_R1222_U483, new_R1222_U484, new_R1222_U485,
    new_R1222_U486, new_R1222_U487, new_R1222_U488, new_R1222_U489,
    new_R1222_U490, new_R1222_U491, new_R1222_U492, new_R1222_U493,
    new_R1222_U494, new_not_keyinput0, new_not_keyinput1,
    new_not_keyinput2, new_not_keyinput3, new_not_keyinput4, new_not_0,
    new_and_1, new_not_2, new_and_3, new_not_4, new_and_5, new_not_6,
    new_and_7, new_not_9, new_and_10, new_not_11, new_and_12, new_not_13,
    new_and_14, new_not_16, new_and_17, new_not_18, new_and_19,
    new_not_Q_0, new_not_Q_1, new_not_Q_2, new_not_Q_3, new_count_state_1,
    new_count_state_2, new_count_state_3, new_count_state_4,
    new_count_state_5, new_count_state_6, new_count_state_7,
    new_count_state_8, new_count_state_9, new_count_state_10,
    new_count_state_11, new_count_state_12, new_count_state_13,
    new_count_state_14, new_count_state_15, new_y_mux_key0_and_0,
    new_y_mux_key0_and_1, new_y_mux_key0, new_y_mux_key1_and_0,
    new_y_mux_key1_and_1, new_y_mux_key1, new_y_mux_key2_and_0,
    new_y_mux_key2_and_1, new_y_mux_key2, new_y_mux_key3_and_0,
    new_y_mux_key3_and_1, new_y_mux_key3, new_y_mux_key4_and_0,
    new_y_mux_key4_and_1, new_y_mux_key4, new_y_mux_key5_and_0,
    new_y_mux_key5_and_1, new_y_mux_key5, new_y_mux_key6_and_0,
    new_y_mux_key6_and_1, new_y_mux_key6, new_y_mux_key7_and_0,
    new_y_mux_key7_and_1, new_y_mux_key7, new_y_mux_key8_and_0,
    new_y_mux_key8_and_1, new_y_mux_key8, new_y_mux_key9_and_0,
    new_y_mux_key9_and_1, new_y_mux_key9, new_y_mux_key10_and_0,
    new_y_mux_key10_and_1, new_y_mux_key10, new_y_mux_key11_and_0,
    new_y_mux_key11_and_1, new_y_mux_key11, new_y_mux_key12_and_0,
    new_y_mux_key12_and_1, new_y_mux_key12, new_y_mux_key13_and_0,
    new_y_mux_key13_and_1, new_y_mux_key13, new_y_mux_key14_and_0,
    new_y_mux_key14_and_1, new_y_mux_key14, new_y_mux_key15_and_0,
    new_y_mux_key15_and_1, new_y_mux_key15, new__state_1, new__state_2,
    new__state_3, new__state_4, new__state_5, new__state_6, new__state_7,
    new__state_8, new__state_9, new__state_10, new__state_11,
    new__state_12, new__state_13, new__state_14, new__state_15,
    new__state_17, new__state_18, new__state_19, new__state_20,
    new__state_21, new__state_22, new__state_23, new__state_25,
    new__state_26, new__state_27, new__state_29, new_s__state_1,
    new_not_s__state_1, new_I0__state_1, new_I1__state_1,
    new_and_mux__state_1, new_and_mux__state_1_2, new_y_mux_16,
    new_s__state_3, new_not_s__state_3, new_I0__state_3, new_I1__state_3,
    new_and_mux__state_3, new_and_mux__state_3_2, new_y_mux_17,
    new_s__state_5, new_not_s__state_5, new_I0__state_5, new_I1__state_5,
    new_and_mux__state_5, new_and_mux__state_5_2, new_y_mux_18,
    new_s__state_7, new_not_s__state_7, new_I0__state_7, new_I1__state_7,
    new_and_mux__state_7, new_and_mux__state_7_2, new_y_mux_19,
    new_s__state_9, new_not_s__state_9, new_I0__state_9, new_I1__state_9,
    new_and_mux__state_9, new_and_mux__state_9_2, new_y_mux_20,
    new_s__state_11, new_not_s__state_11, new_I0__state_11,
    new_I1__state_11, new_and_mux__state_11, new_and_mux__state_11_2,
    new_y_mux_21, new_s__state_13, new_not_s__state_13, new_I0__state_13,
    new_I1__state_13, new_and_mux__state_13, new_and_mux__state_13_2,
    new_y_mux_22, new_s__state_15, new_not_s__state_15, new_I0__state_15,
    new_I1__state_15, new_and_mux__state_15, new_and_mux__state_15_2,
    new_y_mux_23, new_s__state_17, new_not_s__state_17, new_I0__state_17,
    new_I1__state_17, new_and_mux__state_17, new_and_mux__state_17_2,
    new_y_mux_24, new_s__state_19, new_not_s__state_19, new_I0__state_19,
    new_I1__state_19, new_and_mux__state_19, new_and_mux__state_19_2,
    new_y_mux_25, new_s__state_21, new_not_s__state_21, new_I0__state_21,
    new_I1__state_21, new_and_mux__state_21, new_and_mux__state_21_2,
    new_y_mux_26, new_s__state_23, new_not_s__state_23, new_I0__state_23,
    new_I1__state_23, new_and_mux__state_23, new_and_mux__state_23_2,
    new_y_mux_27, new_s__state_25, new_not_s__state_25, new_I0__state_25,
    new_I1__state_25, new_and_mux__state_25, new_and_mux__state_25_2,
    new_y_mux_28, new_s__state_27, new_not_s__state_27, new_I0__state_27,
    new_I1__state_27, new_and_mux__state_27, new_and_mux__state_27_2,
    new_y_mux_29, new_s__state_29, new_not_s__state_29, new_I0__state_29,
    new_I1__state_29, new_and_mux__state_29, new_and_mux__state_29_2, n184,
    n189, n194, n199, n204, n209, n214, n219, n224, n229, n234, n239, n244,
    n249, n254, n259, n264, n269, n274, n279, n284, n289, n294, n299, n304,
    n309, n314, n319, n324, n329, n334, n339, n344, n349, n354, n359, n364,
    n369, n374, n379, n384, n389, n394, n399, n404, n409, n414, n419, n424,
    n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484,
    n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544,
    n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599, n604,
    n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n664,
    n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719, n724,
    n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784,
    n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839, n844,
    n849, n854, n859, n864, n869, n874, n879, n884, n889, n894, n899, n904,
    n909, n914, n919, n924, n929, n934, n939, n944, n949, n954, n959, n964,
    n969, n974, n979, n984, n988, n992, n996, n1000, n1004, n1008, n1012,
    n1016, n1020, n1024, n1028, n1032, n1036, n1040, n1044, n1048, n1052,
    n1056, n1060, n1064, n1068, n1072, n1076, n1080, n1084, n1088, n1092,
    n1096, n1100, n1104, n1108, n1112, n1116, n1120, n1124, n1128, n1132,
    n1136, n1140, n1144, n1148, n1152, n1156, n1160, n1164, n1168, n1172,
    n1176, n1180, n1184, n1188, n1192, n1197, n1202, n1207, n1212, n1217,
    n1222, n1227, n1232, n1237, n1242, n1247, n1252, n1257, n1262, n1267,
    n1272, n1277, n1282, n1287, n1292, n1297, n1302, n1307, n1312, n1317,
    n1322, n1327, n1332, n1337, n1342, n1347, n1351, n20702, n20705,
    n20708, n20711;
  assign new_R1222_U519 = ~new_U3464 | ~new_R1222_U42;
  assign new_R1222_U518 = ~new_U3074 | ~new_R1222_U41;
  assign new_R1222_U517 = ~new_U3486 | ~new_R1222_U71;
  assign new_U3014 = new_U4201 & new_U3431;
  assign new_U3015 = new_U4011 & new_U3456;
  assign new_U3016 = new_U3454 & new_U3455;
  assign new_U3017 = new_U3659 & new_U3654;
  assign new_U3018 = new_U3462 & new_U3463;
  assign new_U3019 = new_U5826 & new_U3462;
  assign new_U3020 = new_U5823 & new_U3463;
  assign new_U3021 = new_U5823 & new_U5826;
  assign new_U3022 = new_U5613 & new_U3355;
  assign new_U3023 = new_U3047 & STATE_REG;
  assign new_U3024 = new_U5808 & new_U5820 & new_U5805;
  assign new_U3025 = new_U3845 & new_U3421;
  assign new_U3026 = new_U4042 & new_U5799;
  assign new_U3027 = new_U4010 & new_U5820;
  assign new_U3028 = new_U3908 & new_U4028;
  assign new_U3029 = new_U3357 & STATE_REG;
  assign new_U3030 = new_U4019 & new_U4044;
  assign new_U3031 = new_U4044 & new_U4021;
  assign new_U3032 = new_U4012 & new_U4044;
  assign new_U3033 = new_U4020 & new_U4044;
  assign new_U3034 = new_U4042 & new_U3454;
  assign new_U3035 = new_U4028 & new_U5799;
  assign new_U3036 = new_U4044 & new_U3026;
  assign new_U3037 = new_U4028 & new_U3454;
  assign new_U3038 = new_U5802 & new_U4938;
  assign new_U3039 = new_U3025 & new_U5802;
  assign new_U3040 = new_U5799 & new_U4938;
  assign new_U3041 = new_U3025 & new_U5799;
  assign new_U3042 = new_U3016 & new_U4938;
  assign new_U3043 = new_U3025 & new_U3016;
  assign new_U3044 = new_U3023 & new_U3421;
  assign new_U3045 = new_U5170 & STATE_REG;
  assign new_U3046 = new_U3023 & new_U5172;
  assign new_U3047 = new_U5748 & new_U3355;
  assign new_U3048 = new_U3660 & new_U3017;
  assign new_U3049 = new_U4765 & new_U4766 & new_U4762 & new_U4759 & new_U4758;
  assign new_U3050 = ~new_U4698 | ~new_U4695 | ~new_U4696 | ~new_U4697;
  assign new_U3051 = ~new_U4717 | ~new_U4714 | ~new_U4715 | ~new_U4716;
  assign new_U3052 = ~new_U4733 | ~new_U4734 | ~new_U4736 | ~new_U4735;
  assign new_U3053 = ~new_U4772 | ~new_U4773 | ~new_U4774;
  assign new_U3054 = ~new_U4679 | ~new_U4676 | ~new_U4677 | ~new_U4678;
  assign new_U3055 = ~new_U4660 | ~new_U4657 | ~new_U4658 | ~new_U4659;
  assign new_U3056 = ~new_U4752 | ~new_U4753 | ~new_U4754;
  assign new_U3057 = ~new_U4258 | ~new_U4259 | ~new_U4261 | ~new_U4260;
  assign new_U3058 = ~new_U4603 | ~new_U4600 | ~new_U4601 | ~new_U4602;
  assign new_U3059 = ~new_U4372 | ~new_U4373 | ~new_U4375 | ~new_U4374;
  assign new_U3060 = ~new_U4391 | ~new_U4392 | ~new_U4394 | ~new_U4393;
  assign new_U3061 = ~new_U4239 | ~new_U4240 | ~new_U4242 | ~new_U4241;
  assign new_U3062 = ~new_U4641 | ~new_U4638 | ~new_U4639 | ~new_U4640;
  assign new_U3063 = ~new_U4622 | ~new_U4619 | ~new_U4620 | ~new_U4621;
  assign new_U3064 = ~new_U4277 | ~new_U4278 | ~new_U4280 | ~new_U4279;
  assign new_U3065 = ~new_U4215 | ~new_U4216 | ~new_U4218 | ~new_U4217;
  assign new_U3066 = ~new_U4505 | ~new_U4506 | ~new_U4508 | ~new_U4507;
  assign new_U3067 = ~new_U4315 | ~new_U4316 | ~new_U4318 | ~new_U4317;
  assign new_U3068 = ~new_U4296 | ~new_U4297 | ~new_U4299 | ~new_U4298;
  assign new_U3069 = ~new_U4410 | ~new_U4411 | ~new_U4413 | ~new_U4412;
  assign new_U3070 = ~new_U4486 | ~new_U4487 | ~new_U4489 | ~new_U4488;
  assign new_U3071 = ~new_U4467 | ~new_U4468 | ~new_U4470 | ~new_U4469;
  assign new_U3072 = ~new_U4584 | ~new_U4581 | ~new_U4582 | ~new_U4583;
  assign new_U3073 = ~new_U4562 | ~new_U4563 | ~new_U4565 | ~new_U4564;
  assign new_U3074 = ~new_U4220 | ~new_U4221 | ~new_U4223 | ~new_U4222;
  assign new_U3075 = ~new_U4196 | ~new_U4197 | ~new_U4199 | ~new_U4198;
  assign new_U3076 = ~new_U4448 | ~new_U4449 | ~new_U4451 | ~new_U4450;
  assign new_U3077 = ~new_U4429 | ~new_U4430 | ~new_U4432 | ~new_U4431;
  assign new_U3078 = ~new_U4543 | ~new_U4544 | ~new_U4546 | ~new_U4545;
  assign new_U3079 = ~new_U4524 | ~new_U4525 | ~new_U4527 | ~new_U4526;
  assign new_U3080 = ~new_U4353 | ~new_U4354 | ~new_U4356 | ~new_U4355;
  assign new_U3081 = ~new_U4334 | ~new_U4335 | ~new_U4337 | ~new_U4336;
  assign new_U3082 = ~new_U5538 | ~new_U5537;
  assign new_U3083 = ~new_U5540 | ~new_U5539;
  assign new_U3084 = ~new_U5546 | ~new_U5545 | ~new_U5544;
  assign new_U3085 = ~new_U5549 | ~new_U5548 | ~new_U5547;
  assign new_U3086 = ~new_U5551 | ~new_U5552 | ~new_U5550;
  assign new_U3087 = ~new_U5555 | ~new_U5554 | ~new_U5553;
  assign new_U3088 = ~new_U5557 | ~new_U5558 | ~new_U5556;
  assign new_U3089 = ~new_U5561 | ~new_U5560 | ~new_U5559;
  assign new_U3090 = ~new_U5563 | ~new_U5564 | ~new_U5562;
  assign new_U3091 = ~new_U5567 | ~new_U5566 | ~new_U5565;
  assign new_U3092 = ~new_U5569 | ~new_U5570 | ~new_U5568;
  assign new_U3093 = ~new_U5573 | ~new_U5572 | ~new_U5571;
  assign new_U3094 = ~new_U5578 | ~new_U5579 | ~new_U5577;
  assign new_U3095 = ~new_U5582 | ~new_U5581 | ~new_U5580;
  assign new_U3096 = ~new_U5585 | ~new_U5584 | ~new_U5583;
  assign new_U3097 = ~new_U5588 | ~new_U5587 | ~new_U5586;
  assign new_U3098 = ~new_U5591 | ~new_U5590 | ~new_U5589;
  assign new_U3099 = ~new_U5594 | ~new_U5593 | ~new_U5592;
  assign new_U3100 = ~new_U5597 | ~new_U5596 | ~new_U5595;
  assign new_U3101 = ~new_U5600 | ~new_U5599 | ~new_U5598;
  assign new_U3102 = ~new_U5603 | ~new_U5602 | ~new_U5601;
  assign new_U3103 = ~new_U5606 | ~new_U5605 | ~new_U5604;
  assign new_U3104 = ~new_U5521 | ~new_U5520 | ~new_U5519;
  assign new_U3105 = ~new_U5524 | ~new_U5523 | ~new_U5522;
  assign new_U3106 = ~new_U5527 | ~new_U5526 | ~new_U5525;
  assign new_U3107 = ~new_U5530 | ~new_U5529 | ~new_U5528;
  assign new_U3108 = ~new_U5533 | ~new_U5532 | ~new_U5531;
  assign new_U3109 = ~new_U5536 | ~new_U5535 | ~new_U5534;
  assign new_U3110 = ~new_U5543 | ~new_U5542 | ~new_U5541;
  assign new_U3111 = ~new_U5576 | ~new_U5575 | ~new_U5574;
  assign new_U3112 = ~new_U5609 | ~new_U5608 | ~new_U5607;
  assign new_U3113 = ~new_U5611 | ~new_U5610;
  assign new_U3114 = ~new_U3926 | ~new_U5441;
  assign new_U3115 = ~new_U3927 | ~new_U5444;
  assign new_U3116 = ~new_U5450 | ~new_U3929;
  assign new_U3117 = ~new_U5453 | ~new_U3931;
  assign new_U3118 = ~new_U5456 | ~new_U3933;
  assign new_U3119 = ~new_U5459 | ~new_U3935;
  assign new_U3120 = ~new_U5462 | ~new_U3937;
  assign new_U3121 = ~new_U5465 | ~new_U3939;
  assign new_U3122 = ~new_U5468 | ~new_U3941;
  assign new_U3123 = ~new_U5471 | ~new_U3943;
  assign new_U3124 = ~new_U5474 | ~new_U3945;
  assign new_U3125 = ~new_U5477 | ~new_U3947;
  assign new_U3126 = ~new_U5484 | ~new_U3950;
  assign new_U3127 = ~new_U5487 | ~new_U3951;
  assign new_U3128 = ~new_U5490 | ~new_U3952;
  assign new_U3129 = ~new_U5493 | ~new_U3953;
  assign new_U3130 = ~new_U5496 | ~new_U3954;
  assign new_U3131 = ~new_U5499 | ~new_U3955;
  assign new_U3132 = ~new_U5502 | ~new_U3956;
  assign new_U3133 = ~new_U5505 | ~new_U3957;
  assign new_U3134 = ~new_U5508 | ~new_U3958;
  assign new_U3135 = ~new_U5511 | ~new_U3959;
  assign new_U3136 = ~new_U5424 | ~new_U3920;
  assign new_U3137 = ~new_U5427 | ~new_U3921;
  assign new_U3138 = ~new_U5430 | ~new_U3922;
  assign new_U3139 = ~new_U5433 | ~new_U3923;
  assign new_U3140 = ~new_U5436 | ~new_U3924;
  assign new_U3141 = ~new_U5439 | ~new_U3925;
  assign new_U3142 = ~new_U5448 | ~new_U3928;
  assign new_U3143 = ~new_U5481 | ~new_U3949;
  assign new_U3144 = ~new_U5514 | ~new_U3960;
  assign new_U3145 = ~new_U5517 | ~new_U3961;
  assign new_U3146 = ~new_U4201 | ~new_U5748;
  assign new_U3147 = ~new_U5808 | ~new_U3372;
  assign n1347 = ~new_U4062 | ~STATE_REG;
  assign n1342 = ~STATE_REG;
  assign new_U3150 = ~new_U5693 | ~new_U5692;
  assign new_U3151 = ~new_U5695 | ~new_U5694;
  assign new_U3152 = ~new_U5697 | ~new_U5696;
  assign new_U3153 = ~new_U5699 | ~new_U5698;
  assign new_U3154 = ~new_U5701 | ~new_U5700;
  assign new_U3155 = ~new_U5703 | ~new_U5702;
  assign new_U3156 = ~new_U5705 | ~new_U5704;
  assign new_U3157 = ~new_U5707 | ~new_U5706;
  assign new_U3158 = ~new_U5709 | ~new_U5708;
  assign new_U3159 = ~new_U5713 | ~new_U5712;
  assign new_U3160 = ~new_U5715 | ~new_U5714;
  assign new_U3161 = ~new_U5717 | ~new_U5716;
  assign new_U3162 = ~new_U5719 | ~new_U5718;
  assign new_U3163 = ~new_U5721 | ~new_U5720;
  assign new_U3164 = ~new_U5723 | ~new_U5722;
  assign new_U3165 = ~new_U5725 | ~new_U5724;
  assign new_U3166 = ~new_U5727 | ~new_U5726;
  assign new_U3167 = ~new_U5729 | ~new_U5728;
  assign new_U3168 = ~new_U5731 | ~new_U5730;
  assign new_U3169 = ~new_U5679 | ~new_U5678;
  assign new_U3170 = ~new_U5681 | ~new_U5680;
  assign new_U3171 = ~new_U5683 | ~new_U5682;
  assign new_U3172 = ~new_U5685 | ~new_U5684;
  assign new_U3173 = ~new_U5687 | ~new_U5686;
  assign new_U3174 = ~new_U5689 | ~new_U5688;
  assign new_U3175 = ~new_U5691 | ~new_U5690;
  assign new_U3176 = ~new_U5711 | ~new_U5710;
  assign new_U3177 = ~new_U5733 | ~new_U5732;
  assign new_U3178 = ~new_U3966 | ~new_U5735;
  assign new_U3179 = ~new_U5634 | ~new_U5633;
  assign new_U3180 = ~new_U5636 | ~new_U5635;
  assign new_U3181 = ~new_U5638 | ~new_U5637;
  assign new_U3182 = ~new_U5640 | ~new_U5639;
  assign new_U3183 = ~new_U5642 | ~new_U5641;
  assign new_U3184 = ~new_U5644 | ~new_U5643;
  assign new_U3185 = ~new_U5646 | ~new_U5645;
  assign new_U3186 = ~new_U5648 | ~new_U5647;
  assign new_U3187 = ~new_U5650 | ~new_U5649;
  assign new_U3188 = ~new_U5654 | ~new_U5653;
  assign new_U3189 = ~new_U5656 | ~new_U5655;
  assign new_U3190 = ~new_U5658 | ~new_U5657;
  assign new_U3191 = ~new_U5660 | ~new_U5659;
  assign new_U3192 = ~new_U5662 | ~new_U5661;
  assign new_U3193 = ~new_U5664 | ~new_U5663;
  assign new_U3194 = ~new_U5666 | ~new_U5665;
  assign new_U3195 = ~new_U5668 | ~new_U5667;
  assign new_U3196 = ~new_U5670 | ~new_U5669;
  assign new_U3197 = ~new_U5672 | ~new_U5671;
  assign new_U3198 = ~new_U5620 | ~new_U5619;
  assign new_U3199 = ~new_U5622 | ~new_U5621;
  assign new_U3200 = ~new_U5624 | ~new_U5623;
  assign new_U3201 = ~new_U5626 | ~new_U5625;
  assign new_U3202 = ~new_U5628 | ~new_U5627;
  assign new_U3203 = ~new_U5630 | ~new_U5629;
  assign new_U3204 = ~new_U5632 | ~new_U5631;
  assign new_U3205 = ~new_U5652 | ~new_U5651;
  assign new_U3206 = ~new_U5674 | ~new_U5673;
  assign new_U3207 = ~new_U3965 | ~new_U5675;
  assign new_U3208 = new_U5612 & new_U3355;
  assign new_U3209 = ~new_U5422 | ~new_U6259 | ~new_U6258;
  assign n1337 = ~new_U5418 | ~new_U5417 | ~new_U5419 | ~new_U5416 | ~new_U5415;
  assign n1332 = ~new_U5409 | ~new_U5408 | ~new_U5410 | ~new_U5407 | ~new_U5406;
  assign n1327 = ~new_U5400 | ~new_U5399 | ~new_U5401 | ~new_U5398 | ~new_U5397;
  assign n1322 = ~new_U5391 | ~new_U5390 | ~new_U5392 | ~new_U5389 | ~new_U5388;
  assign n1317 = ~new_U5382 | ~new_U5381 | ~new_U5383 | ~new_U5380 | ~new_U5379;
  assign n1312 = ~new_U5372 | ~new_U3918 | ~new_U5371;
  assign n1307 = ~new_U5364 | ~new_U5363 | ~new_U5365 | ~new_U5362 | ~new_U5361;
  assign n1302 = ~new_U5355 | ~new_U5354 | ~new_U5356 | ~new_U5353 | ~new_U5352;
  assign n1297 = ~new_U5346 | ~new_U5345 | ~new_U5347 | ~new_U5344 | ~new_U5343;
  assign n1292 = ~new_U5336 | ~new_U3916 | ~new_U5335;
  assign n1287 = ~new_U5328 | ~new_U5327 | ~new_U5329 | ~new_U5326 | ~new_U5325;
  assign n1282 = ~new_U5319 | ~new_U5318 | ~new_U5320 | ~new_U5317 | ~new_U5316;
  assign n1277 = ~new_U5310 | ~new_U5309 | ~new_U5311 | ~new_U5308 | ~new_U5307;
  assign n1272 = ~new_U5301 | ~new_U5300 | ~new_U5302 | ~new_U5299 | ~new_U5298;
  assign n1267 = ~new_U3915 | ~new_U5291 | ~new_U5290 | ~new_U5289;
  assign n1262 = ~new_U5283 | ~new_U5282 | ~new_U5284 | ~new_U5281 | ~new_U5280;
  assign n1257 = ~new_U5274 | ~new_U5273 | ~new_U5275 | ~new_U5272 | ~new_U5271;
  assign n1252 = ~new_U5264 | ~new_U3914 | ~new_U5263 | ~new_U5262;
  assign n1247 = ~new_U5256 | ~new_U5255 | ~new_U5257 | ~new_U5254 | ~new_U5253;
  assign n1242 = ~new_U3912 | ~new_U3913 | ~new_U5246;
  assign n1237 = ~new_U5239 | ~new_U5238 | ~new_U5240 | ~new_U5237 | ~new_U5236;
  assign n1232 = ~new_U5230 | ~new_U5229 | ~new_U5231 | ~new_U5228 | ~new_U5227;
  assign n1227 = ~new_U5221 | ~new_U5220 | ~new_U5222 | ~new_U5219 | ~new_U5218;
  assign n1222 = ~new_U5212 | ~new_U5211 | ~new_U5213 | ~new_U5210 | ~new_U5209;
  assign n1217 = ~new_U5202 | ~new_U3909 | ~new_U5201;
  assign n1212 = ~new_U5194 | ~new_U5193 | ~new_U5195 | ~new_U5192 | ~new_U5191;
  assign n1207 = ~new_U5185 | ~new_U5184 | ~new_U5186 | ~new_U5183 | ~new_U5182;
  assign n1202 = ~new_U5176 | ~new_U5175 | ~new_U5177 | ~new_U5174 | ~new_U5173;
  assign n1197 = ~new_U5163 | ~new_U5162 | ~new_U5164 | ~new_U5161 | ~new_U5160;
  assign n1192 = ~new_U3904 | ~new_U5147;
  assign n1060 = ~new_U3890 | ~new_U3889;
  assign n1056 = ~new_U3888 | ~new_U3887;
  assign n1052 = ~new_U3886 | ~new_U3885;
  assign n1048 = ~new_U3883 | ~new_U3882;
  assign n1044 = ~new_U3881 | ~new_U3880;
  assign n1040 = ~new_U3878 | ~new_U3877;
  assign n1036 = ~new_U3876 | ~new_U3875;
  assign n1032 = ~new_U3874 | ~new_U3873;
  assign n1028 = ~new_U5050 | ~new_U5054 | ~new_U3872 | ~new_U3871;
  assign n1024 = ~new_U5040 | ~new_U5044 | ~new_U3870 | ~new_U3869;
  assign n1020 = ~new_U5030 | ~new_U5034 | ~new_U3868 | ~new_U3867;
  assign n1016 = ~new_U5020 | ~new_U5024 | ~new_U3866 | ~new_U3865;
  assign n1012 = ~new_U5010 | ~new_U5014 | ~new_U3864 | ~new_U3863;
  assign n1008 = ~new_U5000 | ~new_U5004 | ~new_U3862 | ~new_U3861;
  assign n1004 = ~new_U4990 | ~new_U4994 | ~new_U3860 | ~new_U3859;
  assign n1000 = ~new_U4980 | ~new_U4984 | ~new_U3858 | ~new_U3857;
  assign n996 = ~new_U4970 | ~new_U4974 | ~new_U3856 | ~new_U3855;
  assign n992 = ~new_U4960 | ~new_U4964 | ~new_U3854 | ~new_U3853;
  assign n988 = ~new_U3852 | ~new_U3850;
  assign n984 = ~new_U3848 | ~new_U3846;
  assign n979 = ~new_U4004 | ~new_U4937 | ~new_U4936;
  assign n974 = ~new_U4003 | ~new_U4935 | ~new_U4934;
  assign n964 = ~new_U4000 | ~new_U4927 | ~new_U3836 | ~new_U3837;
  assign n959 = ~new_U3999 | ~new_U4922 | ~new_U3834 | ~new_U3835;
  assign n954 = ~new_U3998 | ~new_U4917 | ~new_U3832 | ~new_U3833;
  assign n949 = ~new_U3997 | ~new_U4912 | ~new_U3830 | ~new_U3831;
  assign n944 = ~new_U3996 | ~new_U4907 | ~new_U3828 | ~new_U3829;
  assign n939 = ~new_U3995 | ~new_U4902 | ~new_U3826 | ~new_U3827;
  assign n934 = ~new_U3994 | ~new_U4897 | ~new_U3824 | ~new_U3825;
  assign n929 = ~new_U3993 | ~new_U4892 | ~new_U3822 | ~new_U3823;
  assign n924 = ~new_U3992 | ~new_U4887 | ~new_U3820 | ~new_U3821;
  assign n919 = ~new_U3991 | ~new_U4882 | ~new_U3818 | ~new_U3819;
  assign n914 = ~new_U3990 | ~new_U4877 | ~new_U3816 | ~new_U3817;
  assign n909 = ~new_U3989 | ~new_U4872 | ~new_U3814 | ~new_U3815;
  assign n904 = ~new_U3988 | ~new_U4867 | ~new_U3812 | ~new_U3813;
  assign n899 = ~new_U3987 | ~new_U4862 | ~new_U3810 | ~new_U3811;
  assign n894 = ~new_U3986 | ~new_U3809 | ~new_U3808;
  assign n889 = ~new_U3985 | ~new_U4852 | ~new_U3806 | ~new_U3807;
  assign n884 = ~new_U3984 | ~new_U3805 | ~new_U3804;
  assign n879 = ~new_U3983 | ~new_U3803 | ~new_U3802;
  assign n874 = ~new_U3982 | ~new_U3801 | ~new_U3800;
  assign n869 = ~new_U3981 | ~new_U3799 | ~new_U3798;
  assign n864 = ~new_U3980 | ~new_U3797 | ~new_U3796;
  assign n859 = ~new_U3979 | ~new_U3795 | ~new_U3794;
  assign n854 = ~new_U3978 | ~new_U3793 | ~new_U3792;
  assign n849 = ~new_U3977 | ~new_U3791 | ~new_U3790;
  assign n844 = ~new_U3789 | ~new_U3788;
  assign n839 = ~new_U3787 | ~new_U3786;
  assign n834 = ~new_U3785 | ~new_U3784;
  assign n829 = ~new_U3783 | ~new_U3782;
  assign n824 = ~new_U3781 | ~new_U3780;
  assign n499 = D_REG_31_ & new_U3968;
  assign n494 = D_REG_30_ & new_U3968;
  assign n489 = D_REG_29_ & new_U3968;
  assign n484 = D_REG_28_ & new_U3968;
  assign n479 = D_REG_27_ & new_U3968;
  assign n474 = D_REG_26_ & new_U3968;
  assign n469 = D_REG_25_ & new_U3968;
  assign n464 = D_REG_24_ & new_U3968;
  assign n459 = D_REG_23_ & new_U3968;
  assign n454 = D_REG_22_ & new_U3968;
  assign n449 = D_REG_21_ & new_U3968;
  assign n444 = D_REG_20_ & new_U3968;
  assign n439 = D_REG_19_ & new_U3968;
  assign n434 = D_REG_18_ & new_U3968;
  assign n429 = D_REG_17_ & new_U3968;
  assign n424 = D_REG_16_ & new_U3968;
  assign n419 = D_REG_15_ & new_U3968;
  assign n414 = D_REG_14_ & new_U3968;
  assign n409 = D_REG_13_ & new_U3968;
  assign n404 = D_REG_12_ & new_U3968;
  assign n399 = D_REG_11_ & new_U3968;
  assign n394 = D_REG_10_ & new_U3968;
  assign n389 = D_REG_9_ & new_U3968;
  assign n384 = D_REG_8_ & new_U3968;
  assign n379 = D_REG_7_ & new_U3968;
  assign n374 = D_REG_6_ & new_U3968;
  assign n369 = D_REG_5_ & new_U3968;
  assign n364 = D_REG_4_ & new_U3968;
  assign n359 = D_REG_3_ & new_U3968;
  assign n354 = D_REG_2_ & new_U3968;
  assign n339 = ~new_U3645 | ~new_U4159;
  assign n334 = ~new_U3644 | ~new_U4156;
  assign n329 = ~new_U3643 | ~new_U4153;
  assign n324 = ~new_U3642 | ~new_U4150;
  assign n319 = ~new_U3641 | ~new_U4147;
  assign n314 = ~new_U3640 | ~new_U4144;
  assign n309 = ~new_U3639 | ~new_U4141;
  assign n304 = ~new_U3638 | ~new_U4138;
  assign n299 = ~new_U3637 | ~new_U4135;
  assign n294 = ~new_U3636 | ~new_U4132;
  assign n289 = ~new_U3635 | ~new_U4129;
  assign n284 = ~new_U3634 | ~new_U4126;
  assign n279 = ~new_U3633 | ~new_U4123;
  assign n274 = ~new_U3632 | ~new_U4120;
  assign n269 = ~new_U3631 | ~new_U4117;
  assign n264 = ~new_U3630 | ~new_U4114;
  assign n259 = ~new_U3629 | ~new_U4111;
  assign n254 = ~new_U3628 | ~new_U4108;
  assign n249 = ~new_U3627 | ~new_U4105;
  assign n244 = ~new_U3626 | ~new_U4102;
  assign n239 = ~new_U3625 | ~new_U4099;
  assign n234 = ~new_U3624 | ~new_U4096;
  assign n229 = ~new_U3623 | ~new_U4093;
  assign n224 = ~new_U3622 | ~new_U4090;
  assign n219 = ~new_U3621 | ~new_U4087;
  assign n214 = ~new_U3620 | ~new_U4084;
  assign n209 = ~new_U3619 | ~new_U4081;
  assign n204 = ~new_U3618 | ~new_U4078;
  assign n199 = ~new_U3617 | ~new_U4075;
  assign n194 = ~new_U3616 | ~new_U4072;
  assign n189 = ~new_U3615 | ~new_U4069;
  assign new_U3352 = ~new_U3614 | ~new_U4066;
  assign new_U3353 = ~new_U4055 | ~new_U5805;
  assign n969 = ~new_U4001 | ~new_U4931 | ~new_U4933 | ~new_U4932 | ~new_U4930;
  assign new_U3355 = ~new_U3434 | ~new_U3433 | ~new_U3432;
  assign new_U3356 = ~new_U4059 | ~new_U5748;
  assign new_U3357 = ~STATE_REG | ~new_U3967;
  assign new_U3358 = ~new_U3432 | ~new_U5757;
  assign new_U3359 = ~B_REG;
  assign new_U3360 = ~new_U3432 | ~new_U5810 | ~new_U5809;
  assign new_U3361 = ~new_U5820 | ~new_U3456;
  assign new_U3362 = ~new_U4201 | ~new_U3461;
  assign new_U3363 = ~new_U3460 | ~new_U3461 | ~new_U3456;
  assign new_U3364 = ~new_U3460 | ~new_U5817 | ~new_U3456;
  assign new_U3365 = ~new_U3460 | ~new_U3457;
  assign new_U3366 = ~new_U4056 | ~new_U3461;
  assign new_U3367 = ~new_U4056 | ~new_U5817;
  assign new_U3368 = ~new_U4201 | ~new_U5817;
  assign new_U3369 = ~new_U4015 | ~new_U5808;
  assign new_U3370 = ~new_U3457 | ~new_U5817 | ~new_U5820;
  assign new_U3371 = ~new_U4011 | ~new_U5805;
  assign new_U3372 = ~new_U5805 | ~new_U3461;
  assign new_U3373 = ~new_U3457 | ~new_U3456;
  assign new_U3374 = ~new_U5808 | ~new_U3460;
  assign new_U3375 = ~new_U3646 | ~new_U3647 | ~new_U4208 | ~new_U4207 | ~new_U4206;
  assign new_U3376 = ~REG2_REG_0_;
  assign new_U3377 = ~new_U3664 | ~new_U3662 | ~new_U4226 | ~new_U4225;
  assign new_U3378 = ~new_U3668 | ~new_U3666 | ~new_U4245 | ~new_U4244;
  assign new_U3379 = ~new_U3672 | ~new_U3670 | ~new_U4264 | ~new_U4263;
  assign new_U3380 = ~new_U3676 | ~new_U3674 | ~new_U4283 | ~new_U4282;
  assign new_U3381 = ~new_U3680 | ~new_U3678 | ~new_U4302 | ~new_U4301;
  assign new_U3382 = ~new_U3684 | ~new_U3682 | ~new_U4321 | ~new_U4320;
  assign new_U3383 = ~new_U3688 | ~new_U3686 | ~new_U4340 | ~new_U4339;
  assign new_U3384 = ~new_U3692 | ~new_U3690 | ~new_U4359 | ~new_U4358;
  assign new_U3385 = ~new_U3696 | ~new_U3694 | ~new_U4378 | ~new_U4377;
  assign new_U3386 = ~new_U3700 | ~new_U3698 | ~new_U4397 | ~new_U4396;
  assign new_U3387 = ~new_U3704 | ~new_U3702 | ~new_U4416 | ~new_U4415;
  assign new_U3388 = ~new_U3708 | ~new_U3706 | ~new_U4435 | ~new_U4434;
  assign new_U3389 = ~new_U3712 | ~new_U3710 | ~new_U4454 | ~new_U4453;
  assign new_U3390 = ~new_U3716 | ~new_U3714 | ~new_U4473 | ~new_U4472;
  assign new_U3391 = ~new_U3720 | ~new_U3718 | ~new_U4492 | ~new_U4491;
  assign new_U3392 = ~new_U3724 | ~new_U3722 | ~new_U4511 | ~new_U4510;
  assign new_U3393 = ~new_U3728 | ~new_U3726 | ~new_U4530 | ~new_U4529;
  assign new_U3394 = ~new_U3732 | ~new_U3730 | ~new_U4549 | ~new_U4548;
  assign new_U3395 = ~new_U3736 | ~new_U3734 | ~new_U4568 | ~new_U4567;
  assign new_U3396 = ~DATAI_20_ | ~new_U3969;
  assign new_U3397 = ~new_U3740 | ~new_U3738 | ~new_U4587 | ~new_U4586;
  assign new_U3398 = ~DATAI_21_ | ~new_U3969;
  assign new_U3399 = ~new_U3744 | ~new_U3742 | ~new_U4606 | ~new_U4605;
  assign new_U3400 = ~DATAI_22_ | ~new_U3969;
  assign new_U3401 = ~new_U3748 | ~new_U3746 | ~new_U4625 | ~new_U4624;
  assign new_U3402 = ~DATAI_23_ | ~new_U3969;
  assign new_U3403 = ~new_U3752 | ~new_U3750 | ~new_U4644 | ~new_U4643;
  assign new_U3404 = ~DATAI_24_ | ~new_U3969;
  assign new_U3405 = ~new_U3756 | ~new_U3754 | ~new_U4663 | ~new_U4662;
  assign new_U3406 = ~DATAI_25_ | ~new_U3969;
  assign new_U3407 = ~new_U3760 | ~new_U3758 | ~new_U4682 | ~new_U4681;
  assign new_U3408 = ~DATAI_26_ | ~new_U3969;
  assign new_U3409 = ~new_U3764 | ~new_U3762 | ~new_U4701 | ~new_U4700;
  assign new_U3410 = ~DATAI_27_ | ~new_U3969;
  assign new_U3411 = ~new_U3768 | ~new_U3766 | ~new_U4720 | ~new_U4719;
  assign new_U3412 = ~DATAI_28_ | ~new_U3969;
  assign new_U3413 = ~new_U3772 | ~new_U3770 | ~new_U4739 | ~new_U4738;
  assign new_U3414 = ~DATAI_29_ | ~new_U3969;
  assign new_U3415 = ~DATAI_30_ | ~new_U3969;
  assign new_U3416 = ~DATAI_31_ | ~new_U3969;
  assign new_U3417 = ~new_U3023 | ~new_U4784;
  assign new_U3418 = ~new_U5808 | ~new_U5820 | ~new_U4010;
  assign new_U3419 = ~new_U3457 | ~new_U3461 | ~new_U5820;
  assign new_U3420 = ~new_U3024 | ~new_U5817;
  assign new_U3421 = ~new_U3356 | ~new_U4063;
  assign new_U3422 = ~new_U4054 | ~STATE_REG;
  assign new_U3423 = ~new_U3015 | ~new_U3016;
  assign new_U3424 = ~new_R395_U6;
  assign new_U3425 = ~new_U3901 | ~new_U3900;
  assign new_U3426 = ~new_U3023 | ~new_U4021;
  assign new_U3427 = ~new_U3905 | ~new_U3017;
  assign new_U3428 = ~new_U3015 | ~new_U3023;
  assign new_U3429 = ~new_U3907 | ~new_U5158;
  assign new_U3430 = ~new_U5808 | ~new_U3461;
  assign new_U3431 = ~new_U5747 | ~new_U5746;
  assign new_U3432 = ~new_U5753 | ~new_U5752;
  assign new_U3433 = ~new_U5756 | ~new_U5755;
  assign new_U3434 = ~new_U5750 | ~new_U5749;
  assign new_U3435 = ~new_U5759 | ~new_U5758;
  assign new_U3436 = ~new_U5761 | ~new_U5760;
  assign new_U3437 = ~new_U5763 | ~new_U5762;
  assign new_U3438 = ~new_U5765 | ~new_U5764;
  assign new_U3439 = ~new_U5767 | ~new_U5766;
  assign new_U3440 = ~new_U5769 | ~new_U5768;
  assign new_U3441 = ~new_U5771 | ~new_U5770;
  assign new_U3442 = ~new_U5773 | ~new_U5772;
  assign new_U3443 = ~new_U5775 | ~new_U5774;
  assign new_U3444 = ~new_U5777 | ~new_U5776;
  assign new_U3445 = ~new_U5779 | ~new_U5778;
  assign new_U3446 = ~new_U5781 | ~new_U5780;
  assign new_U3447 = ~new_U5783 | ~new_U5782;
  assign new_U3448 = ~new_U5785 | ~new_U5784;
  assign new_U3449 = ~new_U5787 | ~new_U5786;
  assign new_U3450 = ~new_U5789 | ~new_U5788;
  assign new_U3451 = ~new_U5791 | ~new_U5790;
  assign new_U3452 = ~new_U5793 | ~new_U5792;
  assign new_U3453 = ~new_U5795 | ~new_U5794;
  assign new_U3454 = ~new_U5798 | ~new_U5797;
  assign new_U3455 = ~new_U5801 | ~new_U5800;
  assign new_U3456 = ~new_U5804 | ~new_U5803;
  assign new_U3457 = ~new_U5807 | ~new_U5806;
  assign n344 = ~new_U5812 | ~new_U5811;
  assign n349 = ~new_U5814 | ~new_U5813;
  assign new_U3460 = ~new_U5819 | ~new_U5818;
  assign new_U3461 = ~new_U5816 | ~new_U5815;
  assign new_U3462 = ~new_U5822 | ~new_U5821;
  assign new_U3463 = ~new_U5825 | ~new_U5824;
  assign new_U3464 = ~new_U5828 | ~new_U5827;
  assign new_U3465 = ~new_U5836 | ~new_U5835;
  assign new_U3466 = ~new_U5833 | ~new_U5832;
  assign n504 = ~new_U5839 | ~new_U5838;
  assign new_U3468 = ~new_U5841 | ~new_U5840;
  assign n509 = ~new_U5844 | ~new_U5843;
  assign new_U3470 = ~new_U5846 | ~new_U5845;
  assign n514 = ~new_U5849 | ~new_U5848;
  assign new_U3472 = ~new_U5851 | ~new_U5850;
  assign n519 = ~new_U5854 | ~new_U5853;
  assign new_U3474 = ~new_U5856 | ~new_U5855;
  assign n524 = ~new_U5859 | ~new_U5858;
  assign new_U3476 = ~new_U5861 | ~new_U5860;
  assign n529 = ~new_U5864 | ~new_U5863;
  assign new_U3478 = ~new_U5866 | ~new_U5865;
  assign n534 = ~new_U5869 | ~new_U5868;
  assign new_U3480 = ~new_U5871 | ~new_U5870;
  assign n539 = ~new_U5874 | ~new_U5873;
  assign new_U3482 = ~new_U5876 | ~new_U5875;
  assign n544 = ~new_U5879 | ~new_U5878;
  assign new_U3484 = ~new_U5881 | ~new_U5880;
  assign n549 = ~new_U5884 | ~new_U5883;
  assign new_U3486 = ~new_U5886 | ~new_U5885;
  assign n554 = ~new_U5889 | ~new_U5888;
  assign new_U3488 = ~new_U5891 | ~new_U5890;
  assign n559 = ~new_U5894 | ~new_U5893;
  assign new_U3490 = ~new_U5896 | ~new_U5895;
  assign n564 = ~new_U5899 | ~new_U5898;
  assign new_U3492 = ~new_U5901 | ~new_U5900;
  assign n569 = ~new_U5904 | ~new_U5903;
  assign new_U3494 = ~new_U5906 | ~new_U5905;
  assign n574 = ~new_U5909 | ~new_U5908;
  assign new_U3496 = ~new_U5911 | ~new_U5910;
  assign n579 = ~new_U5914 | ~new_U5913;
  assign new_U3498 = ~new_U5916 | ~new_U5915;
  assign n584 = ~new_U5919 | ~new_U5918;
  assign new_U3500 = ~new_U5921 | ~new_U5920;
  assign n589 = ~new_U5924 | ~new_U5923;
  assign new_U3502 = ~new_U5926 | ~new_U5925;
  assign n594 = ~new_U5929 | ~new_U5928;
  assign new_U3504 = ~new_U5931 | ~new_U5930;
  assign n599 = ~new_U5934 | ~new_U5933;
  assign n604 = ~new_U5936 | ~new_U5935;
  assign n609 = ~new_U5938 | ~new_U5937;
  assign n614 = ~new_U5940 | ~new_U5939;
  assign n619 = ~new_U5942 | ~new_U5941;
  assign n624 = ~new_U5944 | ~new_U5943;
  assign n629 = ~new_U5946 | ~new_U5945;
  assign n634 = ~new_U5948 | ~new_U5947;
  assign n639 = ~new_U5950 | ~new_U5949;
  assign n644 = ~new_U5952 | ~new_U5951;
  assign n649 = ~new_U5954 | ~new_U5953;
  assign n654 = ~new_U5956 | ~new_U5955;
  assign n659 = ~new_U5958 | ~new_U5957;
  assign n664 = ~new_U5960 | ~new_U5959;
  assign n669 = ~new_U5962 | ~new_U5961;
  assign n674 = ~new_U5964 | ~new_U5963;
  assign n679 = ~new_U5966 | ~new_U5965;
  assign n684 = ~new_U5968 | ~new_U5967;
  assign n689 = ~new_U5970 | ~new_U5969;
  assign n694 = ~new_U5972 | ~new_U5971;
  assign n699 = ~new_U5974 | ~new_U5973;
  assign n704 = ~new_U5976 | ~new_U5975;
  assign n709 = ~new_U5978 | ~new_U5977;
  assign n714 = ~new_U5980 | ~new_U5979;
  assign n719 = ~new_U5982 | ~new_U5981;
  assign n724 = ~new_U5984 | ~new_U5983;
  assign n729 = ~new_U5986 | ~new_U5985;
  assign n734 = ~new_U5988 | ~new_U5987;
  assign n739 = ~new_U5990 | ~new_U5989;
  assign n744 = ~new_U5992 | ~new_U5991;
  assign n749 = ~new_U5994 | ~new_U5993;
  assign n754 = ~new_U5996 | ~new_U5995;
  assign n759 = ~new_U5998 | ~new_U5997;
  assign n764 = ~new_U6000 | ~new_U5999;
  assign n769 = ~new_U6002 | ~new_U6001;
  assign n774 = ~new_U6004 | ~new_U6003;
  assign n779 = ~new_U6006 | ~new_U6005;
  assign n784 = ~new_U6008 | ~new_U6007;
  assign n789 = ~new_U6010 | ~new_U6009;
  assign n794 = ~new_U6012 | ~new_U6011;
  assign n799 = ~new_U6014 | ~new_U6013;
  assign n804 = ~new_U6016 | ~new_U6015;
  assign n809 = ~new_U6018 | ~new_U6017;
  assign n814 = ~new_U6020 | ~new_U6019;
  assign n819 = ~new_U6022 | ~new_U6021;
  assign n1064 = ~new_U6088 | ~new_U6087;
  assign n1068 = ~new_U6090 | ~new_U6089;
  assign n1072 = ~new_U6092 | ~new_U6091;
  assign n1076 = ~new_U6094 | ~new_U6093;
  assign n1080 = ~new_U6096 | ~new_U6095;
  assign n1084 = ~new_U6098 | ~new_U6097;
  assign n1088 = ~new_U6100 | ~new_U6099;
  assign n1092 = ~new_U6102 | ~new_U6101;
  assign n1096 = ~new_U6104 | ~new_U6103;
  assign n1100 = ~new_U6106 | ~new_U6105;
  assign n1104 = ~new_U6108 | ~new_U6107;
  assign n1108 = ~new_U6110 | ~new_U6109;
  assign n1112 = ~new_U6112 | ~new_U6111;
  assign n1116 = ~new_U6114 | ~new_U6113;
  assign n1120 = ~new_U6116 | ~new_U6115;
  assign n1124 = ~new_U6118 | ~new_U6117;
  assign n1128 = ~new_U6120 | ~new_U6119;
  assign n1132 = ~new_U6122 | ~new_U6121;
  assign n1136 = ~new_U6124 | ~new_U6123;
  assign n1140 = ~new_U6126 | ~new_U6125;
  assign n1144 = ~new_U6128 | ~new_U6127;
  assign n1148 = ~new_U6130 | ~new_U6129;
  assign n1152 = ~new_U6132 | ~new_U6131;
  assign n1156 = ~new_U6134 | ~new_U6133;
  assign n1160 = ~new_U6136 | ~new_U6135;
  assign n1164 = ~new_U6138 | ~new_U6137;
  assign n1168 = ~new_U6140 | ~new_U6139;
  assign n1172 = ~new_U6142 | ~new_U6141;
  assign n1176 = ~new_U6144 | ~new_U6143;
  assign n1180 = ~new_U6146 | ~new_U6145;
  assign n1184 = ~new_U6148 | ~new_U6147;
  assign n1188 = ~new_U6150 | ~new_U6149;
  assign new_U3582 = ~new_U6261 | ~new_U6260;
  assign new_U3583 = ~new_U6263 | ~new_U6262;
  assign new_U3584 = ~new_U6265 | ~new_U6264;
  assign new_U3585 = ~new_U6267 | ~new_U6266;
  assign new_U3586 = ~new_U6269 | ~new_U6268;
  assign new_U3587 = ~new_U6271 | ~new_U6270;
  assign new_U3588 = ~new_U6273 | ~new_U6272;
  assign new_U3589 = ~new_U6275 | ~new_U6274;
  assign new_U3590 = ~new_U6277 | ~new_U6276;
  assign new_U3591 = ~new_U6279 | ~new_U6278;
  assign new_U3592 = ~new_U6281 | ~new_U6280;
  assign new_U3593 = ~new_U6283 | ~new_U6282;
  assign new_U3594 = ~new_U6285 | ~new_U6284;
  assign new_U3595 = ~new_U6287 | ~new_U6286;
  assign new_U3596 = ~new_U6289 | ~new_U6288;
  assign new_U3597 = ~new_U6291 | ~new_U6290;
  assign new_U3598 = ~new_U6293 | ~new_U6292;
  assign new_U3599 = ~new_U6295 | ~new_U6294;
  assign new_U3600 = ~new_U6297 | ~new_U6296;
  assign new_U3601 = ~new_U6299 | ~new_U6298;
  assign new_U3602 = ~new_U6301 | ~new_U6300;
  assign new_U3603 = ~new_U6303 | ~new_U6302;
  assign new_U3604 = ~new_U6305 | ~new_U6304;
  assign new_U3605 = ~new_U6307 | ~new_U6306;
  assign new_U3606 = ~new_U6309 | ~new_U6308;
  assign new_U3607 = ~new_U6311 | ~new_U6310;
  assign new_U3608 = ~new_U6313 | ~new_U6312;
  assign new_U3609 = ~new_U6315 | ~new_U6314;
  assign new_U3610 = ~new_U6317 | ~new_U6316;
  assign new_U3611 = ~new_U6319 | ~new_U6318;
  assign new_U3612 = ~new_U6321 | ~new_U6320;
  assign new_U3613 = ~new_U6323 | ~new_U6322;
  assign new_U3614 = new_U4067 & new_U4065;
  assign new_U3615 = new_U4070 & new_U4068;
  assign new_U3616 = new_U4073 & new_U4071;
  assign new_U3617 = new_U4076 & new_U4074;
  assign new_U3618 = new_U4079 & new_U4077;
  assign new_U3619 = new_U4082 & new_U4080;
  assign new_U3620 = new_U4085 & new_U4083;
  assign new_U3621 = new_U4088 & new_U4086;
  assign new_U3622 = new_U4091 & new_U4089;
  assign new_U3623 = new_U4094 & new_U4092;
  assign new_U3624 = new_U4097 & new_U4095;
  assign new_U3625 = new_U4100 & new_U4098;
  assign new_U3626 = new_U4103 & new_U4101;
  assign new_U3627 = new_U4106 & new_U4104;
  assign new_U3628 = new_U4109 & new_U4107;
  assign new_U3629 = new_U4112 & new_U4110;
  assign new_U3630 = new_U4115 & new_U4113;
  assign new_U3631 = new_U4118 & new_U4116;
  assign new_U3632 = new_U4121 & new_U4119;
  assign new_U3633 = new_U4124 & new_U4122;
  assign new_U3634 = new_U4127 & new_U4125;
  assign new_U3635 = new_U4130 & new_U4128;
  assign new_U3636 = new_U4133 & new_U4131;
  assign new_U3637 = new_U4136 & new_U4134;
  assign new_U3638 = new_U4139 & new_U4137;
  assign new_U3639 = new_U4142 & new_U4140;
  assign new_U3640 = new_U4145 & new_U4143;
  assign new_U3641 = new_U4148 & new_U4146;
  assign new_U3642 = new_U4151 & new_U4149;
  assign new_U3643 = new_U4154 & new_U4152;
  assign new_U3644 = new_U4157 & new_U4155;
  assign new_U3645 = new_U4160 & new_U4158;
  assign new_U3646 = new_U4203 & new_U4202;
  assign new_U3647 = new_U4205 & new_U4204;
  assign new_U3648 = new_U4212 & new_U4210;
  assign new_U3649 = new_U3648 & new_U4213 & new_U4211;
  assign new_U3650 = new_U4164 & new_U4165 & new_U4167 & new_U4166;
  assign new_U3651 = new_U4168 & new_U4169 & new_U4171 & new_U4170;
  assign new_U3652 = new_U4172 & new_U4173 & new_U4175 & new_U4174;
  assign new_U3653 = new_U4178 & new_U4177 & new_U4176;
  assign new_U3654 = new_U3650 & new_U3651 & new_U3653 & new_U3652;
  assign new_U3655 = new_U4179 & new_U4180 & new_U4182 & new_U4181;
  assign new_U3656 = new_U4183 & new_U4184 & new_U4186 & new_U4185;
  assign new_U3657 = new_U4187 & new_U4188 & new_U4190 & new_U4189;
  assign new_U3658 = new_U4193 & new_U4192 & new_U4191;
  assign new_U3659 = new_U3655 & new_U3656 & new_U3658 & new_U3657;
  assign new_U3660 = new_U5834 & new_U4195;
  assign new_U3661 = new_U5837 & new_U3023;
  assign new_U3662 = new_U4228 & new_U4227;
  assign new_U3663 = new_U4230 & new_U4229;
  assign new_U3664 = new_U3663 & new_U4232 & new_U4231;
  assign new_U3665 = new_U4234 & new_U4237 & new_U4235 & new_U4236;
  assign new_U3666 = new_U4247 & new_U4246;
  assign new_U3667 = new_U4249 & new_U4248;
  assign new_U3668 = new_U3667 & new_U4251 & new_U4250;
  assign new_U3669 = new_U4253 & new_U4256 & new_U4254 & new_U4255;
  assign new_U3670 = new_U4266 & new_U4265;
  assign new_U3671 = new_U4268 & new_U4267;
  assign new_U3672 = new_U3671 & new_U4270 & new_U4269;
  assign new_U3673 = new_U4272 & new_U4275 & new_U4273 & new_U4274;
  assign new_U3674 = new_U4285 & new_U4284;
  assign new_U3675 = new_U4287 & new_U4286;
  assign new_U3676 = new_U3675 & new_U4289 & new_U4288;
  assign new_U3677 = new_U4291 & new_U4294 & new_U4292 & new_U4293;
  assign new_U3678 = new_U4304 & new_U4303;
  assign new_U3679 = new_U4306 & new_U4305;
  assign new_U3680 = new_U3679 & new_U4308 & new_U4307;
  assign new_U3681 = new_U4310 & new_U4313 & new_U4311 & new_U4312;
  assign new_U3682 = new_U4323 & new_U4322;
  assign new_U3683 = new_U4325 & new_U4324;
  assign new_U3684 = new_U3683 & new_U4327 & new_U4326;
  assign new_U3685 = new_U4329 & new_U4332 & new_U4330 & new_U4331;
  assign new_U3686 = new_U4342 & new_U4341;
  assign new_U3687 = new_U4344 & new_U4343;
  assign new_U3688 = new_U3687 & new_U4346 & new_U4345;
  assign new_U3689 = new_U4348 & new_U4351 & new_U4349 & new_U4350;
  assign new_U3690 = new_U4361 & new_U4360;
  assign new_U3691 = new_U4363 & new_U4362;
  assign new_U3692 = new_U3691 & new_U4365 & new_U4364;
  assign new_U3693 = new_U4367 & new_U4370 & new_U4368 & new_U4369;
  assign new_U3694 = new_U4380 & new_U4379;
  assign new_U3695 = new_U4382 & new_U4381;
  assign new_U3696 = new_U3695 & new_U4384 & new_U4383;
  assign new_U3697 = new_U4386 & new_U4389 & new_U4387 & new_U4388;
  assign new_U3698 = new_U4399 & new_U4398;
  assign new_U3699 = new_U4401 & new_U4400;
  assign new_U3700 = new_U3699 & new_U4403 & new_U4402;
  assign new_U3701 = new_U4405 & new_U4408 & new_U4406 & new_U4407;
  assign new_U3702 = new_U4418 & new_U4417;
  assign new_U3703 = new_U4420 & new_U4419;
  assign new_U3704 = new_U3703 & new_U4422 & new_U4421;
  assign new_U3705 = new_U4424 & new_U4427 & new_U4425 & new_U4426;
  assign new_U3706 = new_U4437 & new_U4436;
  assign new_U3707 = new_U4439 & new_U4438;
  assign new_U3708 = new_U3707 & new_U4441 & new_U4440;
  assign new_U3709 = new_U4443 & new_U4446 & new_U4444 & new_U4445;
  assign new_U3710 = new_U4456 & new_U4455;
  assign new_U3711 = new_U4458 & new_U4457;
  assign new_U3712 = new_U3711 & new_U4460 & new_U4459;
  assign new_U3713 = new_U4462 & new_U4465 & new_U4463 & new_U4464;
  assign new_U3714 = new_U4475 & new_U4474;
  assign new_U3715 = new_U4477 & new_U4476;
  assign new_U3716 = new_U3715 & new_U4479 & new_U4478;
  assign new_U3717 = new_U4481 & new_U4484 & new_U4482 & new_U4483;
  assign new_U3718 = new_U4494 & new_U4493;
  assign new_U3719 = new_U4496 & new_U4495;
  assign new_U3720 = new_U3719 & new_U4498 & new_U4497;
  assign new_U3721 = new_U4500 & new_U4503 & new_U4501 & new_U4502;
  assign new_U3722 = new_U4513 & new_U4512;
  assign new_U3723 = new_U4515 & new_U4514;
  assign new_U3724 = new_U3723 & new_U4517 & new_U4516;
  assign new_U3725 = new_U4519 & new_U4522 & new_U4520 & new_U4521;
  assign new_U3726 = new_U4532 & new_U4531;
  assign new_U3727 = new_U4534 & new_U4533;
  assign new_U3728 = new_U3727 & new_U4536 & new_U4535;
  assign new_U3729 = new_U4538 & new_U4541 & new_U4539 & new_U4540;
  assign new_U3730 = new_U4551 & new_U4550;
  assign new_U3731 = new_U4553 & new_U4552;
  assign new_U3732 = new_U3731 & new_U4555 & new_U4554;
  assign new_U3733 = new_U4557 & new_U4560 & new_U4558 & new_U4559;
  assign new_U3734 = new_U4570 & new_U4569;
  assign new_U3735 = new_U4572 & new_U4571;
  assign new_U3736 = new_U3735 & new_U4574 & new_U4573;
  assign new_U3737 = new_U4576 & new_U4579 & new_U4577 & new_U4578;
  assign new_U3738 = new_U4589 & new_U4588;
  assign new_U3739 = new_U4591 & new_U4590;
  assign new_U3740 = new_U3739 & new_U4593 & new_U4592;
  assign new_U3741 = new_U4595 & new_U4598 & new_U4596 & new_U4597;
  assign new_U3742 = new_U4608 & new_U4607;
  assign new_U3743 = new_U4610 & new_U4609;
  assign new_U3744 = new_U3743 & new_U4612 & new_U4611;
  assign new_U3745 = new_U4614 & new_U4617 & new_U4615 & new_U4616;
  assign new_U3746 = new_U4627 & new_U4626;
  assign new_U3747 = new_U4629 & new_U4628;
  assign new_U3748 = new_U3747 & new_U4631 & new_U4630;
  assign new_U3749 = new_U4633 & new_U4636 & new_U4634 & new_U4635;
  assign new_U3750 = new_U4646 & new_U4645;
  assign new_U3751 = new_U4648 & new_U4647;
  assign new_U3752 = new_U3751 & new_U4650 & new_U4649;
  assign new_U3753 = new_U4652 & new_U4655 & new_U4653 & new_U4654;
  assign new_U3754 = new_U4665 & new_U4664;
  assign new_U3755 = new_U4667 & new_U4666;
  assign new_U3756 = new_U3755 & new_U4669 & new_U4668;
  assign new_U3757 = new_U4671 & new_U4674 & new_U4672 & new_U4673;
  assign new_U3758 = new_U4684 & new_U4683;
  assign new_U3759 = new_U4686 & new_U4685;
  assign new_U3760 = new_U3759 & new_U4688 & new_U4687;
  assign new_U3761 = new_U4690 & new_U4693 & new_U4691 & new_U4692;
  assign new_U3762 = new_U4703 & new_U4702;
  assign new_U3763 = new_U4705 & new_U4704;
  assign new_U3764 = new_U3763 & new_U4707 & new_U4706;
  assign new_U3765 = new_U4709 & new_U4712 & new_U4710 & new_U4711;
  assign new_U3766 = new_U4722 & new_U4721;
  assign new_U3767 = new_U4724 & new_U4723;
  assign new_U3768 = new_U3767 & new_U4726 & new_U4725;
  assign new_U3769 = new_U4728 & new_U4731 & new_U4729 & new_U4730;
  assign new_U3770 = new_U4741 & new_U4740;
  assign new_U3771 = new_U4743 & new_U4742;
  assign new_U3772 = new_U3771 & new_U4745 & new_U4744;
  assign new_U3773 = new_U4747 & new_U4750 & new_U4748 & new_U4749;
  assign new_U3774 = new_U4757 & new_U4042;
  assign new_U3775 = new_U4760 & new_U4761 & new_U4764 & new_U4763;
  assign new_U3776 = new_U4768 & new_U4769 & new_U4770;
  assign new_U3777 = new_U4042 & new_U4757;
  assign new_U3778 = new_U3023 & new_U3465;
  assign new_U3779 = new_U3466 & new_U5837 & new_U4025;
  assign new_U3780 = new_U4787 & new_U4786 & new_U4785;
  assign new_U3781 = new_U3972 & new_U4789 & new_U4788;
  assign new_U3782 = new_U4792 & new_U4791 & new_U4790;
  assign new_U3783 = new_U3973 & new_U4794 & new_U4793;
  assign new_U3784 = new_U4797 & new_U4796 & new_U4795;
  assign new_U3785 = new_U3974 & new_U4799 & new_U4798;
  assign new_U3786 = new_U4802 & new_U4801 & new_U4800;
  assign new_U3787 = new_U3975 & new_U4804 & new_U4803;
  assign new_U3788 = new_U4807 & new_U4806 & new_U4805;
  assign new_U3789 = new_U3976 & new_U4809 & new_U4808;
  assign new_U3790 = new_U4812 & new_U4811 & new_U4810;
  assign new_U3791 = new_U4814 & new_U4813;
  assign new_U3792 = new_U4817 & new_U4816 & new_U4815;
  assign new_U3793 = new_U4819 & new_U4818;
  assign new_U3794 = new_U4822 & new_U4821 & new_U4820;
  assign new_U3795 = new_U4824 & new_U4823;
  assign new_U3796 = new_U4827 & new_U4826 & new_U4825;
  assign new_U3797 = new_U4829 & new_U4828;
  assign new_U3798 = new_U4832 & new_U4831 & new_U4830;
  assign new_U3799 = new_U4834 & new_U4833;
  assign new_U3800 = new_U4837 & new_U4836 & new_U4835;
  assign new_U3801 = new_U4839 & new_U4838;
  assign new_U3802 = new_U4842 & new_U4841 & new_U4840;
  assign new_U3803 = new_U4844 & new_U4843;
  assign new_U3804 = new_U4847 & new_U4846 & new_U4845;
  assign new_U3805 = new_U4849 & new_U4848;
  assign new_U3806 = new_U4851 & new_U4850;
  assign new_U3807 = new_U4854 & new_U4853;
  assign new_U3808 = new_U4857 & new_U4856 & new_U4855;
  assign new_U3809 = new_U4859 & new_U4858;
  assign new_U3810 = new_U4861 & new_U4860;
  assign new_U3811 = new_U4864 & new_U4863;
  assign new_U3812 = new_U4866 & new_U4865;
  assign new_U3813 = new_U4869 & new_U4868;
  assign new_U3814 = new_U4871 & new_U4870;
  assign new_U3815 = new_U4874 & new_U4873;
  assign new_U3816 = new_U4876 & new_U4875;
  assign new_U3817 = new_U4879 & new_U4878;
  assign new_U3818 = new_U4881 & new_U4880;
  assign new_U3819 = new_U4884 & new_U4883;
  assign new_U3820 = new_U4886 & new_U4885;
  assign new_U3821 = new_U4889 & new_U4888;
  assign new_U3822 = new_U4891 & new_U4890;
  assign new_U3823 = new_U4894 & new_U4893;
  assign new_U3824 = new_U4896 & new_U4895;
  assign new_U3825 = new_U4899 & new_U4898;
  assign new_U3826 = new_U4901 & new_U4900;
  assign new_U3827 = new_U4904 & new_U4903;
  assign new_U3828 = new_U4906 & new_U4905;
  assign new_U3829 = new_U4909 & new_U4908;
  assign new_U3830 = new_U4911 & new_U4910;
  assign new_U3831 = new_U4914 & new_U4913;
  assign new_U3832 = new_U4916 & new_U4915;
  assign new_U3833 = new_U4919 & new_U4918;
  assign new_U3834 = new_U4921 & new_U4920;
  assign new_U3835 = new_U4924 & new_U4923;
  assign new_U3836 = new_U4926 & new_U4925;
  assign new_U3837 = new_U4929 & new_U4928;
  assign new_U3838 = new_U5739 & new_U5738 & new_U5737;
  assign new_U3839 = new_U3367 & new_U3419 & new_U3370;
  assign new_U3840 = new_U3366 & new_U3368 & new_U3362;
  assign new_U3841 = new_U3363 & new_U3364;
  assign new_U3842 = new_U3841 & new_U3420;
  assign new_U3843 = new_U3353 & new_U3418;
  assign new_U3844 = new_U3040 & new_U3461;
  assign new_U3845 = new_U3431 & STATE_REG;
  assign new_U3846 = new_U4941 & new_U4943 & new_U4940 & new_U4939;
  assign new_U3847 = new_U4947 & new_U4944;
  assign new_U3848 = new_U4946 & new_U4945 & new_U3847;
  assign new_U3849 = new_U3040 & new_U3444;
  assign new_U3850 = new_U4950 & new_U4951 & new_U4949 & new_U4948;
  assign new_U3851 = new_U4955 & new_U4952;
  assign new_U3852 = new_U4954 & new_U4953 & new_U3851;
  assign new_U3853 = new_U4961 & new_U4962;
  assign new_U3854 = new_U4965 & new_U4963;
  assign new_U3855 = new_U4971 & new_U4972;
  assign new_U3856 = new_U4975 & new_U4973;
  assign new_U3857 = new_U4981 & new_U4982;
  assign new_U3858 = new_U4985 & new_U4983;
  assign new_U3859 = new_U4991 & new_U4992;
  assign new_U3860 = new_U4995 & new_U4993;
  assign new_U3861 = new_U5001 & new_U5002;
  assign new_U3862 = new_U5005 & new_U5003;
  assign new_U3863 = new_U5011 & new_U5012;
  assign new_U3864 = new_U5015 & new_U5013;
  assign new_U3865 = new_U5021 & new_U5022;
  assign new_U3866 = new_U5025 & new_U5023;
  assign new_U3867 = new_U5031 & new_U5032;
  assign new_U3868 = new_U5035 & new_U5033;
  assign new_U3869 = new_U5041 & new_U5042;
  assign new_U3870 = new_U5045 & new_U5043;
  assign new_U3871 = new_U5051 & new_U5052;
  assign new_U3872 = new_U5055 & new_U5053;
  assign new_U3873 = new_U5060 & new_U5061 & new_U5062;
  assign new_U3874 = new_U5065 & new_U5064 & new_U5063;
  assign new_U3875 = new_U5070 & new_U5071 & new_U5072;
  assign new_U3876 = new_U5075 & new_U5074 & new_U5073;
  assign new_U3877 = new_U5080 & new_U5081 & new_U5082;
  assign new_U3878 = new_U5085 & new_U5084 & new_U5083;
  assign new_U3879 = new_U5090 & new_U4053;
  assign new_U3880 = new_U3879 & new_U5092 & new_U5091;
  assign new_U3881 = new_U5095 & new_U5094 & new_U5093;
  assign new_U3882 = new_U5100 & new_U5101 & new_U5102;
  assign new_U3883 = new_U5105 & new_U5104 & new_U5103;
  assign new_U3884 = new_U5110 & new_U4053;
  assign new_U3885 = new_U3884 & new_U5112 & new_U5111;
  assign new_U3886 = new_U5115 & new_U5114 & new_U5113;
  assign new_U3887 = new_U5120 & new_U5121 & new_U5122;
  assign new_U3888 = new_U5125 & new_U5124 & new_U5123;
  assign new_U3889 = new_U5130 & new_U5131 & new_U5132;
  assign new_U3890 = new_U5135 & new_U5134 & new_U5133;
  assign new_U3891 = new_U6201 & new_U6204 & new_U6210 & new_U6207;
  assign new_U3892 = new_U6213 & new_U6216 & new_U6222 & new_U6219;
  assign new_U3893 = new_U6225 & new_U6228 & new_U6234 & new_U6231;
  assign new_U3894 = new_U6237 & new_U6240 & new_U6246 & new_U6243;
  assign new_U3895 = new_U6165 & new_U6168 & new_U6174 & new_U6171;
  assign new_U3896 = new_U6162 & new_U6159 & new_U6156;
  assign new_U3897 = new_U6183 & new_U6186 & new_U6192 & new_U6189;
  assign new_U3898 = new_U6180 & new_U6177;
  assign new_U3899 = new_U6198 & new_U6195;
  assign new_U3900 = new_U3898 & new_U3897 & new_U6153 & new_U3895 & new_U3896;
  assign new_U3901 = new_U3899 & new_U3891 & new_U3892 & new_U3894 & new_U3893;
  assign new_U3902 = new_U5140 & new_U5141 & new_U6255 & new_U6254;
  assign new_U3903 = new_U3356 & STATE_REG;
  assign new_U3904 = new_U5148 & new_U5146;
  assign new_U3905 = new_U3465 & new_U3466;
  assign new_U3906 = new_U4008 & new_U3371 & new_U3420;
  assign new_U3907 = new_U5748 & new_U3356 & new_U4025;
  assign new_U3908 = new_U3023 & new_U5157;
  assign new_U3909 = new_U3910 & new_U5200;
  assign new_U3910 = new_U5204 & new_U5203;
  assign new_U3911 = new_U4049 & new_U3075;
  assign new_U3912 = new_U5245 & new_U5244;
  assign new_U3913 = new_U5248 & new_U5247;
  assign new_U3914 = new_U5266 & new_U5265;
  assign new_U3915 = new_U5293 & new_U5292;
  assign new_U3916 = new_U3917 & new_U5334;
  assign new_U3917 = new_U5338 & new_U5337;
  assign new_U3918 = new_U3919 & new_U5370;
  assign new_U3919 = new_U5374 & new_U5373;
  assign new_U3920 = new_U5425 & new_U3431 & new_U5423;
  assign new_U3921 = new_U5428 & new_U3431 & new_U5426;
  assign new_U3922 = new_U5431 & new_U3431 & new_U5429;
  assign new_U3923 = new_U5434 & new_U3431 & new_U5432;
  assign new_U3924 = new_U5437 & new_U3431 & new_U5435;
  assign new_U3925 = new_U5440 & new_U3431 & new_U5438;
  assign new_U3926 = new_U5442 & new_U5443;
  assign new_U3927 = new_U5445 & new_U5446;
  assign new_U3928 = new_U5449 & new_U3431 & new_U5447;
  assign new_U3929 = new_U5452 & new_U3930;
  assign new_U3930 = new_U3431 & new_U5451;
  assign new_U3931 = new_U5455 & new_U3932;
  assign new_U3932 = new_U3431 & new_U5454;
  assign new_U3933 = new_U5458 & new_U3934;
  assign new_U3934 = new_U3431 & new_U5457;
  assign new_U3935 = new_U5461 & new_U3936;
  assign new_U3936 = new_U3431 & new_U5460;
  assign new_U3937 = new_U5464 & new_U3938;
  assign new_U3938 = new_U3431 & new_U5463;
  assign new_U3939 = new_U5467 & new_U3940;
  assign new_U3940 = new_U3431 & new_U5466;
  assign new_U3941 = new_U5470 & new_U3942;
  assign new_U3942 = new_U3431 & new_U5469;
  assign new_U3943 = new_U5473 & new_U3944;
  assign new_U3944 = new_U3431 & new_U5472;
  assign new_U3945 = new_U5476 & new_U3946;
  assign new_U3946 = new_U3431 & new_U5475;
  assign new_U3947 = new_U5479 & new_U3948;
  assign new_U3948 = new_U3431 & new_U5478;
  assign new_U3949 = new_U5482 & new_U3431 & new_U5480;
  assign new_U3950 = new_U5485 & new_U3431 & new_U5483;
  assign new_U3951 = new_U5488 & new_U3431 & new_U5486;
  assign new_U3952 = new_U5491 & new_U3431 & new_U5489;
  assign new_U3953 = new_U5494 & new_U3431 & new_U5492;
  assign new_U3954 = new_U5497 & new_U3431 & new_U5495;
  assign new_U3955 = new_U5500 & new_U3431 & new_U5498;
  assign new_U3956 = new_U5503 & new_U3431 & new_U5501;
  assign new_U3957 = new_U5506 & new_U3431 & new_U5504;
  assign new_U3958 = new_U5509 & new_U3431 & new_U5507;
  assign new_U3959 = new_U5512 & new_U3431 & new_U5510;
  assign new_U3960 = new_U5515 & new_U3431 & new_U5513;
  assign new_U3961 = new_U5518 & new_U3431 & new_U5516;
  assign new_U3962 = new_U5808 & new_U5805;
  assign new_U3963 = new_U3365 & new_U3430;
  assign new_U3964 = new_U5616 & new_U4026;
  assign new_U3965 = new_U5676 & new_U5677;
  assign new_U3966 = new_U5736 & new_U5734;
  assign new_U3967 = ~IR_REG_31_;
  assign new_U3968 = ~new_U3023 | ~new_U3360;
  assign new_U3969 = ~new_U5802 | ~new_U5799;
  assign new_U3970 = ~new_U3661 | ~new_U3048;
  assign new_U3971 = ~new_U3778 | ~new_U3048;
  assign new_U3972 = new_U6024 & new_U6023;
  assign new_U3973 = new_U6026 & new_U6025;
  assign new_U3974 = new_U6028 & new_U6027;
  assign new_U3975 = new_U6030 & new_U6029;
  assign new_U3976 = new_U6032 & new_U6031;
  assign new_U3977 = new_U6034 & new_U6033;
  assign new_U3978 = new_U6036 & new_U6035;
  assign new_U3979 = new_U6038 & new_U6037;
  assign new_U3980 = new_U6040 & new_U6039;
  assign new_U3981 = new_U6042 & new_U6041;
  assign new_U3982 = new_U6044 & new_U6043;
  assign new_U3983 = new_U6046 & new_U6045;
  assign new_U3984 = new_U6048 & new_U6047;
  assign new_U3985 = new_U6050 & new_U6049;
  assign new_U3986 = new_U6052 & new_U6051;
  assign new_U3987 = new_U6054 & new_U6053;
  assign new_U3988 = new_U6056 & new_U6055;
  assign new_U3989 = new_U6058 & new_U6057;
  assign new_U3990 = new_U6060 & new_U6059;
  assign new_U3991 = new_U6062 & new_U6061;
  assign new_U3992 = new_U6064 & new_U6063;
  assign new_U3993 = new_U6066 & new_U6065;
  assign new_U3994 = new_U6068 & new_U6067;
  assign new_U3995 = new_U6070 & new_U6069;
  assign new_U3996 = new_U6072 & new_U6071;
  assign new_U3997 = new_U6074 & new_U6073;
  assign new_U3998 = new_U6076 & new_U6075;
  assign new_U3999 = new_U6078 & new_U6077;
  assign new_U4000 = new_U6080 & new_U6079;
  assign new_U4001 = new_U6082 & new_U6081;
  assign new_U4002 = ~new_U3777 | ~new_U3053;
  assign new_U4003 = new_U6084 & new_U6083;
  assign new_U4004 = new_U6086 & new_U6085;
  assign new_U4005 = ~new_R1375_U26;
  assign new_U4006 = new_U6251 & new_U6250;
  assign new_U4007 = ~new_R1347_U13;
  assign new_U4008 = ~new_U4013 | ~new_U5805;
  assign new_U4009 = ~new_R1352_U6;
  assign new_U4010 = ~new_U3372;
  assign new_U4011 = ~new_U3370;
  assign new_U4012 = ~new_U3419;
  assign new_U4013 = ~new_U3367;
  assign new_U4014 = ~new_U3366;
  assign new_U4015 = ~new_U3368;
  assign new_U4016 = ~new_U3362;
  assign new_U4017 = ~new_U3364;
  assign new_U4018 = ~new_U3363;
  assign new_U4019 = ~new_U3420;
  assign new_U4020 = ~new_U3418;
  assign new_U4021 = ~new_U3353;
  assign new_U4022 = ~new_U3371;
  assign new_U4023 = ~new_U4008;
  assign new_U4024 = ~new_U3369;
  assign new_U4025 = ~new_U4042 | ~new_U4782;
  assign new_U4026 = ~new_U3962 | ~new_U3355;
  assign new_U4027 = ~new_U3969;
  assign new_U4028 = ~new_U3427;
  assign new_U4029 = ~new_U3412;
  assign new_U4030 = ~new_U3410;
  assign new_U4031 = ~new_U3408;
  assign new_U4032 = ~new_U3406;
  assign new_U4033 = ~new_U3404;
  assign new_U4034 = ~new_U3402;
  assign new_U4035 = ~new_U3400;
  assign new_U4036 = ~new_U3398;
  assign new_U4037 = ~new_U3396;
  assign new_U4038 = ~new_U3416;
  assign new_U4039 = ~new_U3415;
  assign new_U4040 = ~new_U3414;
  assign new_U4041 = ~new_U3423;
  assign new_U4042 = ~new_U3373;
  assign n1351 = ~new_U3422;
  assign new_U4044 = ~new_U3417;
  assign new_U4045 = ~new_U3971;
  assign new_U4046 = ~new_U3970;
  assign new_U4047 = ~new_U3968;
  assign new_U4048 = ~new_U4002;
  assign new_U4049 = ~new_U3428;
  assign new_U4050 = ~new_U3429 | ~STATE_REG;
  assign new_U4051 = ~new_U4020 | ~new_U3023;
  assign new_U4052 = ~new_U3426;
  assign new_U4053 = ~n1351 | ~new_U3209;
  assign new_U4054 = ~new_U3356;
  assign new_U4055 = ~new_U3374;
  assign new_U4056 = ~new_U3365;
  assign new_U4057 = ~new_U3430;
  assign new_U4058 = ~new_U3358;
  assign new_U4059 = ~new_U3355;
  assign new_U4060 = ~new_U3047 | ~new_U3373;
  assign new_U4061 = ~new_U5748 | ~new_U4060;
  assign new_U4062 = ~new_U4061 | ~new_U3969;
  assign new_U4063 = ~n1347;
  assign new_U4064 = ~new_U3357;
  assign new_U4065 = ~DATAI_0_ | ~n1342;
  assign new_U4066 = ~new_U3029 | ~IR_REG_0_;
  assign new_U4067 = ~new_U4064 | ~IR_REG_0_;
  assign new_U4068 = ~DATAI_1_ | ~n1342;
  assign new_U4069 = ~new_U3029 | ~new_SUB_84_U48;
  assign new_U4070 = ~new_U4064 | ~IR_REG_1_;
  assign new_U4071 = ~DATAI_2_ | ~n1342;
  assign new_U4072 = ~new_U3029 | ~new_SUB_84_U20;
  assign new_U4073 = ~new_U4064 | ~IR_REG_2_;
  assign new_U4074 = ~DATAI_3_ | ~n1342;
  assign new_U4075 = ~new_U3029 | ~new_SUB_84_U21;
  assign new_U4076 = ~new_U4064 | ~IR_REG_3_;
  assign new_U4077 = ~DATAI_4_ | ~n1342;
  assign new_U4078 = ~new_U3029 | ~new_SUB_84_U70;
  assign new_U4079 = ~new_U4064 | ~IR_REG_4_;
  assign new_U4080 = ~DATAI_5_ | ~n1342;
  assign new_U4081 = ~new_U3029 | ~new_SUB_84_U22;
  assign new_U4082 = ~new_U4064 | ~IR_REG_5_;
  assign new_U4083 = ~DATAI_6_ | ~n1342;
  assign new_U4084 = ~new_U3029 | ~new_SUB_84_U23;
  assign new_U4085 = ~new_U4064 | ~IR_REG_6_;
  assign new_U4086 = ~DATAI_7_ | ~n1342;
  assign new_U4087 = ~new_U3029 | ~new_SUB_84_U24;
  assign new_U4088 = ~new_U4064 | ~IR_REG_7_;
  assign new_U4089 = ~DATAI_8_ | ~n1342;
  assign new_U4090 = ~new_U3029 | ~new_SUB_84_U68;
  assign new_U4091 = ~new_U4064 | ~IR_REG_8_;
  assign new_U4092 = ~DATAI_9_ | ~n1342;
  assign new_U4093 = ~new_U3029 | ~new_SUB_84_U25;
  assign new_U4094 = ~new_U4064 | ~IR_REG_9_;
  assign new_U4095 = ~DATAI_10_ | ~n1342;
  assign new_U4096 = ~new_U3029 | ~new_SUB_84_U6;
  assign new_U4097 = ~new_U4064 | ~IR_REG_10_;
  assign new_U4098 = ~DATAI_11_ | ~n1342;
  assign new_U4099 = ~new_U3029 | ~new_SUB_84_U7;
  assign new_U4100 = ~new_U4064 | ~IR_REG_11_;
  assign new_U4101 = ~DATAI_12_ | ~n1342;
  assign new_U4102 = ~new_U3029 | ~new_SUB_84_U89;
  assign new_U4103 = ~new_U4064 | ~IR_REG_12_;
  assign new_U4104 = ~DATAI_13_ | ~n1342;
  assign new_U4105 = ~new_U3029 | ~new_SUB_84_U8;
  assign new_U4106 = ~new_U4064 | ~IR_REG_13_;
  assign new_U4107 = ~DATAI_14_ | ~n1342;
  assign new_U4108 = ~new_U3029 | ~new_SUB_84_U9;
  assign new_U4109 = ~new_U4064 | ~IR_REG_14_;
  assign new_U4110 = ~DATAI_15_ | ~n1342;
  assign new_U4111 = ~new_U3029 | ~new_SUB_84_U10;
  assign new_U4112 = ~new_U4064 | ~IR_REG_15_;
  assign new_U4113 = ~DATAI_16_ | ~n1342;
  assign new_U4114 = ~new_U3029 | ~new_SUB_84_U87;
  assign new_U4115 = ~new_U4064 | ~IR_REG_16_;
  assign new_U4116 = ~DATAI_17_ | ~n1342;
  assign new_U4117 = ~new_U3029 | ~new_SUB_84_U11;
  assign new_U4118 = ~new_U4064 | ~IR_REG_17_;
  assign new_U4119 = ~DATAI_18_ | ~n1342;
  assign new_U4120 = ~new_U3029 | ~new_SUB_84_U12;
  assign new_U4121 = ~new_U4064 | ~IR_REG_18_;
  assign new_U4122 = ~DATAI_19_ | ~n1342;
  assign new_U4123 = ~new_SUB_84_U13 | ~new_U3029;
  assign new_U4124 = ~IR_REG_19_ | ~new_U4064;
  assign new_U4125 = ~DATAI_20_ | ~n1342;
  assign new_U4126 = ~new_SUB_84_U83 | ~new_U3029;
  assign new_U4127 = ~IR_REG_20_ | ~new_U4064;
  assign new_U4128 = ~DATAI_21_ | ~n1342;
  assign new_U4129 = ~new_U3029 | ~new_SUB_84_U14;
  assign new_U4130 = ~new_U4064 | ~IR_REG_21_;
  assign new_U4131 = ~DATAI_22_ | ~n1342;
  assign new_U4132 = ~new_U3029 | ~new_SUB_84_U15;
  assign new_U4133 = ~new_U4064 | ~IR_REG_22_;
  assign new_U4134 = ~DATAI_23_ | ~n1342;
  assign new_U4135 = ~new_U3029 | ~new_SUB_84_U81;
  assign new_U4136 = ~new_U4064 | ~IR_REG_23_;
  assign new_U4137 = ~DATAI_24_ | ~n1342;
  assign new_U4138 = ~new_U3029 | ~new_SUB_84_U78;
  assign new_U4139 = ~new_U4064 | ~IR_REG_24_;
  assign new_U4140 = ~DATAI_25_ | ~n1342;
  assign new_U4141 = ~new_U3029 | ~new_SUB_84_U16;
  assign new_U4142 = ~new_U4064 | ~IR_REG_25_;
  assign new_U4143 = ~DATAI_26_ | ~n1342;
  assign new_U4144 = ~new_U3029 | ~new_SUB_84_U17;
  assign new_U4145 = ~new_U4064 | ~IR_REG_26_;
  assign new_U4146 = ~DATAI_27_ | ~n1342;
  assign new_U4147 = ~new_U3029 | ~new_SUB_84_U76;
  assign new_U4148 = ~new_U4064 | ~IR_REG_27_;
  assign new_U4149 = ~DATAI_28_ | ~n1342;
  assign new_U4150 = ~new_U3029 | ~new_SUB_84_U18;
  assign new_U4151 = ~new_U4064 | ~IR_REG_28_;
  assign new_U4152 = ~DATAI_29_ | ~n1342;
  assign new_U4153 = ~new_SUB_84_U19 | ~new_U3029;
  assign new_U4154 = ~IR_REG_29_ | ~new_U4064;
  assign new_U4155 = ~DATAI_30_ | ~n1342;
  assign new_U4156 = ~new_SUB_84_U73 | ~new_U3029;
  assign new_U4157 = ~IR_REG_30_ | ~new_U4064;
  assign new_U4158 = ~DATAI_31_ | ~n1342;
  assign new_U4159 = ~new_SUB_84_U49 | ~new_U3029;
  assign new_U4160 = ~IR_REG_31_ | ~new_U4064;
  assign new_U4161 = ~new_U3360;
  assign new_U4162 = ~new_U3358 | ~new_U5751;
  assign new_U4163 = ~new_U3358 | ~new_U5757;
  assign new_U4164 = ~new_U4161 | ~D_REG_10_;
  assign new_U4165 = ~new_U4161 | ~D_REG_11_;
  assign new_U4166 = ~new_U4161 | ~D_REG_12_;
  assign new_U4167 = ~new_U4161 | ~D_REG_13_;
  assign new_U4168 = ~new_U4161 | ~D_REG_14_;
  assign new_U4169 = ~new_U4161 | ~D_REG_15_;
  assign new_U4170 = ~new_U4161 | ~D_REG_16_;
  assign new_U4171 = ~new_U4161 | ~D_REG_17_;
  assign new_U4172 = ~new_U4161 | ~D_REG_18_;
  assign new_U4173 = ~new_U4161 | ~D_REG_19_;
  assign new_U4174 = ~new_U4161 | ~D_REG_20_;
  assign new_U4175 = ~new_U4161 | ~D_REG_21_;
  assign new_U4176 = ~new_U4161 | ~D_REG_22_;
  assign new_U4177 = ~new_U4161 | ~D_REG_23_;
  assign new_U4178 = ~new_U4161 | ~D_REG_24_;
  assign new_U4179 = ~new_U4161 | ~D_REG_25_;
  assign new_U4180 = ~new_U4161 | ~D_REG_26_;
  assign new_U4181 = ~new_U4161 | ~D_REG_27_;
  assign new_U4182 = ~new_U4161 | ~D_REG_28_;
  assign new_U4183 = ~new_U4161 | ~D_REG_29_;
  assign new_U4184 = ~new_U4161 | ~D_REG_2_;
  assign new_U4185 = ~new_U4161 | ~D_REG_30_;
  assign new_U4186 = ~new_U4161 | ~D_REG_31_;
  assign new_U4187 = ~new_U4161 | ~D_REG_3_;
  assign new_U4188 = ~new_U4161 | ~D_REG_4_;
  assign new_U4189 = ~new_U4161 | ~D_REG_5_;
  assign new_U4190 = ~new_U4161 | ~D_REG_6_;
  assign new_U4191 = ~new_U4161 | ~D_REG_7_;
  assign new_U4192 = ~new_U4161 | ~D_REG_8_;
  assign new_U4193 = ~new_U4161 | ~D_REG_9_;
  assign new_U4194 = ~new_U5820 | ~new_U5817;
  assign new_U4195 = ~new_U5830 | ~new_U5831 | ~new_U4194 | ~new_U3374;
  assign new_U4196 = ~new_U3019 | ~REG2_REG_1_;
  assign new_U4197 = ~new_U3020 | ~REG1_REG_1_;
  assign new_U4198 = ~new_U3021 | ~REG0_REG_1_;
  assign new_U4199 = ~REG3_REG_1_ | ~new_U3018;
  assign new_U4200 = ~new_U3075;
  assign new_U4201 = ~new_U3361;
  assign new_U4202 = ~new_U4016 | ~new_R1150_U31;
  assign new_U4203 = ~new_U4018 | ~new_R1117_U30;
  assign new_U4204 = ~new_U4017 | ~new_R1138_U108;
  assign new_U4205 = ~new_U4014 | ~new_R1192_U32;
  assign new_U4206 = ~new_U4013 | ~new_R1207_U32;
  assign new_U4207 = ~new_U4024 | ~new_R1171_U108;
  assign new_U4208 = ~new_U4022 | ~new_R1240_U108;
  assign new_U4209 = ~new_U3375;
  assign new_U4210 = ~new_R1222_U104 | ~new_U3027;
  assign new_U4211 = ~new_U3026 | ~new_U3075;
  assign new_U4212 = ~new_U3464 | ~new_U3024;
  assign new_U4213 = ~new_U3464 | ~new_U4021;
  assign new_U4214 = ~new_U3649 | ~new_U4209;
  assign new_U4215 = ~REG2_REG_2_ | ~new_U3019;
  assign new_U4216 = ~REG1_REG_2_ | ~new_U3020;
  assign new_U4217 = ~REG0_REG_2_ | ~new_U3021;
  assign new_U4218 = ~REG3_REG_2_ | ~new_U3018;
  assign new_U4219 = ~new_U3065;
  assign new_U4220 = ~REG0_REG_0_ | ~new_U3021;
  assign new_U4221 = ~REG1_REG_0_ | ~new_U3020;
  assign new_U4222 = ~REG2_REG_0_ | ~new_U3019;
  assign new_U4223 = ~REG3_REG_0_ | ~new_U3018;
  assign new_U4224 = ~new_U3074;
  assign new_U4225 = ~new_U3034 | ~new_U3074;
  assign new_U4226 = ~new_R1150_U114 | ~new_U4016;
  assign new_U4227 = ~new_R1117_U113 | ~new_U4018;
  assign new_U4228 = ~new_R1138_U107 | ~new_U4017;
  assign new_U4229 = ~new_R1192_U114 | ~new_U4014;
  assign new_U4230 = ~new_R1207_U114 | ~new_U4013;
  assign new_U4231 = ~new_R1171_U107 | ~new_U4024;
  assign new_U4232 = ~new_R1240_U107 | ~new_U4022;
  assign new_U4233 = ~new_U3377;
  assign new_U4234 = ~new_R1222_U103 | ~new_U3027;
  assign new_U4235 = ~new_U3026 | ~new_U3065;
  assign new_U4236 = ~new_R1282_U31 | ~new_U3024;
  assign new_U4237 = ~new_U3468 | ~new_U4021;
  assign new_U4238 = ~new_U3665 | ~new_U4233;
  assign new_U4239 = ~REG2_REG_3_ | ~new_U3019;
  assign new_U4240 = ~REG1_REG_3_ | ~new_U3020;
  assign new_U4241 = ~REG0_REG_3_ | ~new_U3021;
  assign new_U4242 = ~new_ADD_95_U4 | ~new_U3018;
  assign new_U4243 = ~new_U3061;
  assign new_U4244 = ~new_U3034 | ~new_U3075;
  assign new_U4245 = ~new_R1150_U124 | ~new_U4016;
  assign new_U4246 = ~new_R1117_U123 | ~new_U4018;
  assign new_U4247 = ~new_R1138_U24 | ~new_U4017;
  assign new_U4248 = ~new_R1192_U124 | ~new_U4014;
  assign new_U4249 = ~new_R1207_U124 | ~new_U4013;
  assign new_U4250 = ~new_R1171_U24 | ~new_U4024;
  assign new_U4251 = ~new_R1240_U24 | ~new_U4022;
  assign new_U4252 = ~new_U3378;
  assign new_U4253 = ~new_R1222_U23 | ~new_U3027;
  assign new_U4254 = ~new_U3026 | ~new_U3061;
  assign new_U4255 = ~new_R1282_U6 | ~new_U3024;
  assign new_U4256 = ~new_U3470 | ~new_U4021;
  assign new_U4257 = ~new_U3669 | ~new_U4252;
  assign new_U4258 = ~REG2_REG_4_ | ~new_U3019;
  assign new_U4259 = ~REG1_REG_4_ | ~new_U3020;
  assign new_U4260 = ~REG0_REG_4_ | ~new_U3021;
  assign new_U4261 = ~new_ADD_95_U51 | ~new_U3018;
  assign new_U4262 = ~new_U3057;
  assign new_U4263 = ~new_U3034 | ~new_U3065;
  assign new_U4264 = ~new_R1150_U28 | ~new_U4016;
  assign new_U4265 = ~new_R1117_U27 | ~new_U4018;
  assign new_U4266 = ~new_R1138_U113 | ~new_U4017;
  assign new_U4267 = ~new_R1192_U29 | ~new_U4014;
  assign new_U4268 = ~new_R1207_U29 | ~new_U4013;
  assign new_U4269 = ~new_R1171_U113 | ~new_U4024;
  assign new_U4270 = ~new_R1240_U113 | ~new_U4022;
  assign new_U4271 = ~new_U3379;
  assign new_U4272 = ~new_R1222_U109 | ~new_U3027;
  assign new_U4273 = ~new_U3026 | ~new_U3057;
  assign new_U4274 = ~new_R1282_U7 | ~new_U3024;
  assign new_U4275 = ~new_U3472 | ~new_U4021;
  assign new_U4276 = ~new_U3673 | ~new_U4271;
  assign new_U4277 = ~REG2_REG_5_ | ~new_U3019;
  assign new_U4278 = ~REG1_REG_5_ | ~new_U3020;
  assign new_U4279 = ~REG0_REG_5_ | ~new_U3021;
  assign new_U4280 = ~new_ADD_95_U50 | ~new_U3018;
  assign new_U4281 = ~new_U3064;
  assign new_U4282 = ~new_U3034 | ~new_U3061;
  assign new_U4283 = ~new_R1150_U123 | ~new_U4016;
  assign new_U4284 = ~new_R1117_U122 | ~new_U4018;
  assign new_U4285 = ~new_R1138_U112 | ~new_U4017;
  assign new_U4286 = ~new_R1192_U123 | ~new_U4014;
  assign new_U4287 = ~new_R1207_U123 | ~new_U4013;
  assign new_U4288 = ~new_R1171_U112 | ~new_U4024;
  assign new_U4289 = ~new_R1240_U112 | ~new_U4022;
  assign new_U4290 = ~new_U3380;
  assign new_U4291 = ~new_R1222_U108 | ~new_U3027;
  assign new_U4292 = ~new_U3026 | ~new_U3064;
  assign new_U4293 = ~new_R1282_U8 | ~new_U3024;
  assign new_U4294 = ~new_U3474 | ~new_U4021;
  assign new_U4295 = ~new_U3677 | ~new_U4290;
  assign new_U4296 = ~REG2_REG_6_ | ~new_U3019;
  assign new_U4297 = ~REG1_REG_6_ | ~new_U3020;
  assign new_U4298 = ~REG0_REG_6_ | ~new_U3021;
  assign new_U4299 = ~new_ADD_95_U49 | ~new_U3018;
  assign new_U4300 = ~new_U3068;
  assign new_U4301 = ~new_U3034 | ~new_U3057;
  assign new_U4302 = ~new_R1150_U122 | ~new_U4016;
  assign new_U4303 = ~new_R1117_U121 | ~new_U4018;
  assign new_U4304 = ~new_R1138_U25 | ~new_U4017;
  assign new_U4305 = ~new_R1192_U122 | ~new_U4014;
  assign new_U4306 = ~new_R1207_U122 | ~new_U4013;
  assign new_U4307 = ~new_R1171_U25 | ~new_U4024;
  assign new_U4308 = ~new_R1240_U25 | ~new_U4022;
  assign new_U4309 = ~new_U3381;
  assign new_U4310 = ~new_R1222_U24 | ~new_U3027;
  assign new_U4311 = ~new_U3026 | ~new_U3068;
  assign new_U4312 = ~new_R1282_U9 | ~new_U3024;
  assign new_U4313 = ~new_U3476 | ~new_U4021;
  assign new_U4314 = ~new_U3681 | ~new_U4309;
  assign new_U4315 = ~REG2_REG_7_ | ~new_U3019;
  assign new_U4316 = ~REG1_REG_7_ | ~new_U3020;
  assign new_U4317 = ~REG0_REG_7_ | ~new_U3021;
  assign new_U4318 = ~new_ADD_95_U48 | ~new_U3018;
  assign new_U4319 = ~new_U3067;
  assign new_U4320 = ~new_U3034 | ~new_U3064;
  assign new_U4321 = ~new_R1150_U29 | ~new_U4016;
  assign new_U4322 = ~new_R1117_U28 | ~new_U4018;
  assign new_U4323 = ~new_R1138_U111 | ~new_U4017;
  assign new_U4324 = ~new_R1192_U30 | ~new_U4014;
  assign new_U4325 = ~new_R1207_U30 | ~new_U4013;
  assign new_U4326 = ~new_R1171_U111 | ~new_U4024;
  assign new_U4327 = ~new_R1240_U111 | ~new_U4022;
  assign new_U4328 = ~new_U3382;
  assign new_U4329 = ~new_R1222_U107 | ~new_U3027;
  assign new_U4330 = ~new_U3026 | ~new_U3067;
  assign new_U4331 = ~new_R1282_U10 | ~new_U3024;
  assign new_U4332 = ~new_U3478 | ~new_U4021;
  assign new_U4333 = ~new_U3685 | ~new_U4328;
  assign new_U4334 = ~REG2_REG_8_ | ~new_U3019;
  assign new_U4335 = ~REG1_REG_8_ | ~new_U3020;
  assign new_U4336 = ~REG0_REG_8_ | ~new_U3021;
  assign new_U4337 = ~new_ADD_95_U47 | ~new_U3018;
  assign new_U4338 = ~new_U3081;
  assign new_U4339 = ~new_U3034 | ~new_U3068;
  assign new_U4340 = ~new_R1150_U121 | ~new_U4016;
  assign new_U4341 = ~new_R1117_U120 | ~new_U4018;
  assign new_U4342 = ~new_R1138_U26 | ~new_U4017;
  assign new_U4343 = ~new_R1192_U121 | ~new_U4014;
  assign new_U4344 = ~new_R1207_U121 | ~new_U4013;
  assign new_U4345 = ~new_R1171_U26 | ~new_U4024;
  assign new_U4346 = ~new_R1240_U26 | ~new_U4022;
  assign new_U4347 = ~new_U3383;
  assign new_U4348 = ~new_R1222_U25 | ~new_U3027;
  assign new_U4349 = ~new_U3026 | ~new_U3081;
  assign new_U4350 = ~new_R1282_U11 | ~new_U3024;
  assign new_U4351 = ~new_U3480 | ~new_U4021;
  assign new_U4352 = ~new_U3689 | ~new_U4347;
  assign new_U4353 = ~REG2_REG_9_ | ~new_U3019;
  assign new_U4354 = ~REG1_REG_9_ | ~new_U3020;
  assign new_U4355 = ~REG0_REG_9_ | ~new_U3021;
  assign new_U4356 = ~new_ADD_95_U46 | ~new_U3018;
  assign new_U4357 = ~new_U3080;
  assign new_U4358 = ~new_U3034 | ~new_U3067;
  assign new_U4359 = ~new_R1150_U30 | ~new_U4016;
  assign new_U4360 = ~new_R1117_U29 | ~new_U4018;
  assign new_U4361 = ~new_R1138_U110 | ~new_U4017;
  assign new_U4362 = ~new_R1192_U31 | ~new_U4014;
  assign new_U4363 = ~new_R1207_U31 | ~new_U4013;
  assign new_U4364 = ~new_R1171_U110 | ~new_U4024;
  assign new_U4365 = ~new_R1240_U110 | ~new_U4022;
  assign new_U4366 = ~new_U3384;
  assign new_U4367 = ~new_R1222_U106 | ~new_U3027;
  assign new_U4368 = ~new_U3026 | ~new_U3080;
  assign new_U4369 = ~new_R1282_U36 | ~new_U3024;
  assign new_U4370 = ~new_U3482 | ~new_U4021;
  assign new_U4371 = ~new_U3693 | ~new_U4366;
  assign new_U4372 = ~REG2_REG_10_ | ~new_U3019;
  assign new_U4373 = ~REG1_REG_10_ | ~new_U3020;
  assign new_U4374 = ~REG0_REG_10_ | ~new_U3021;
  assign new_U4375 = ~new_ADD_95_U70 | ~new_U3018;
  assign new_U4376 = ~new_U3059;
  assign new_U4377 = ~new_U3034 | ~new_U3081;
  assign new_U4378 = ~new_R1150_U120 | ~new_U4016;
  assign new_U4379 = ~new_R1117_U119 | ~new_U4018;
  assign new_U4380 = ~new_R1138_U109 | ~new_U4017;
  assign new_U4381 = ~new_R1192_U120 | ~new_U4014;
  assign new_U4382 = ~new_R1207_U120 | ~new_U4013;
  assign new_U4383 = ~new_R1171_U109 | ~new_U4024;
  assign new_U4384 = ~new_R1240_U109 | ~new_U4022;
  assign new_U4385 = ~new_U3385;
  assign new_U4386 = ~new_R1222_U105 | ~new_U3027;
  assign new_U4387 = ~new_U3026 | ~new_U3059;
  assign new_U4388 = ~new_R1282_U33 | ~new_U3024;
  assign new_U4389 = ~new_U3484 | ~new_U4021;
  assign new_U4390 = ~new_U3697 | ~new_U4385;
  assign new_U4391 = ~REG2_REG_11_ | ~new_U3019;
  assign new_U4392 = ~REG1_REG_11_ | ~new_U3020;
  assign new_U4393 = ~REG0_REG_11_ | ~new_U3021;
  assign new_U4394 = ~new_ADD_95_U69 | ~new_U3018;
  assign new_U4395 = ~new_U3060;
  assign new_U4396 = ~new_U3034 | ~new_U3080;
  assign new_U4397 = ~new_R1150_U130 | ~new_U4016;
  assign new_U4398 = ~new_R1117_U129 | ~new_U4018;
  assign new_U4399 = ~new_R1138_U18 | ~new_U4017;
  assign new_U4400 = ~new_R1192_U130 | ~new_U4014;
  assign new_U4401 = ~new_R1207_U130 | ~new_U4013;
  assign new_U4402 = ~new_R1171_U18 | ~new_U4024;
  assign new_U4403 = ~new_R1240_U18 | ~new_U4022;
  assign new_U4404 = ~new_U3386;
  assign new_U4405 = ~new_R1222_U17 | ~new_U3027;
  assign new_U4406 = ~new_U3026 | ~new_U3060;
  assign new_U4407 = ~new_R1282_U94 | ~new_U3024;
  assign new_U4408 = ~new_U3486 | ~new_U4021;
  assign new_U4409 = ~new_U3701 | ~new_U4404;
  assign new_U4410 = ~REG2_REG_12_ | ~new_U3019;
  assign new_U4411 = ~REG1_REG_12_ | ~new_U3020;
  assign new_U4412 = ~REG0_REG_12_ | ~new_U3021;
  assign new_U4413 = ~new_ADD_95_U68 | ~new_U3018;
  assign new_U4414 = ~new_U3069;
  assign new_U4415 = ~new_U3034 | ~new_U3059;
  assign new_U4416 = ~new_R1150_U23 | ~new_U4016;
  assign new_U4417 = ~new_R1117_U23 | ~new_U4018;
  assign new_U4418 = ~new_R1138_U127 | ~new_U4017;
  assign new_U4419 = ~new_R1192_U24 | ~new_U4014;
  assign new_U4420 = ~new_R1207_U24 | ~new_U4013;
  assign new_U4421 = ~new_R1171_U127 | ~new_U4024;
  assign new_U4422 = ~new_R1240_U127 | ~new_U4022;
  assign new_U4423 = ~new_U3387;
  assign new_U4424 = ~new_R1222_U123 | ~new_U3027;
  assign new_U4425 = ~new_U3026 | ~new_U3069;
  assign new_U4426 = ~new_R1282_U91 | ~new_U3024;
  assign new_U4427 = ~new_U3488 | ~new_U4021;
  assign new_U4428 = ~new_U3705 | ~new_U4423;
  assign new_U4429 = ~REG2_REG_13_ | ~new_U3019;
  assign new_U4430 = ~REG1_REG_13_ | ~new_U3020;
  assign new_U4431 = ~REG0_REG_13_ | ~new_U3021;
  assign new_U4432 = ~new_ADD_95_U67 | ~new_U3018;
  assign new_U4433 = ~new_U3077;
  assign new_U4434 = ~new_U3034 | ~new_U3060;
  assign new_U4435 = ~new_R1150_U119 | ~new_U4016;
  assign new_U4436 = ~new_R1117_U118 | ~new_U4018;
  assign new_U4437 = ~new_R1138_U126 | ~new_U4017;
  assign new_U4438 = ~new_R1192_U119 | ~new_U4014;
  assign new_U4439 = ~new_R1207_U119 | ~new_U4013;
  assign new_U4440 = ~new_R1171_U126 | ~new_U4024;
  assign new_U4441 = ~new_R1240_U126 | ~new_U4022;
  assign new_U4442 = ~new_U3388;
  assign new_U4443 = ~new_R1222_U122 | ~new_U3027;
  assign new_U4444 = ~new_U3026 | ~new_U3077;
  assign new_U4445 = ~new_R1282_U89 | ~new_U3024;
  assign new_U4446 = ~new_U3490 | ~new_U4021;
  assign new_U4447 = ~new_U3709 | ~new_U4442;
  assign new_U4448 = ~REG2_REG_14_ | ~new_U3019;
  assign new_U4449 = ~REG1_REG_14_ | ~new_U3020;
  assign new_U4450 = ~REG0_REG_14_ | ~new_U3021;
  assign new_U4451 = ~new_ADD_95_U66 | ~new_U3018;
  assign new_U4452 = ~new_U3076;
  assign new_U4453 = ~new_U3034 | ~new_U3069;
  assign new_U4454 = ~new_R1150_U118 | ~new_U4016;
  assign new_U4455 = ~new_R1117_U117 | ~new_U4018;
  assign new_U4456 = ~new_R1138_U19 | ~new_U4017;
  assign new_U4457 = ~new_R1192_U118 | ~new_U4014;
  assign new_U4458 = ~new_R1207_U118 | ~new_U4013;
  assign new_U4459 = ~new_R1171_U19 | ~new_U4024;
  assign new_U4460 = ~new_R1240_U19 | ~new_U4022;
  assign new_U4461 = ~new_U3389;
  assign new_U4462 = ~new_R1222_U18 | ~new_U3027;
  assign new_U4463 = ~new_U3026 | ~new_U3076;
  assign new_U4464 = ~new_R1282_U86 | ~new_U3024;
  assign new_U4465 = ~new_U3492 | ~new_U4021;
  assign new_U4466 = ~new_U3713 | ~new_U4461;
  assign new_U4467 = ~REG2_REG_15_ | ~new_U3019;
  assign new_U4468 = ~REG1_REG_15_ | ~new_U3020;
  assign new_U4469 = ~REG0_REG_15_ | ~new_U3021;
  assign new_U4470 = ~new_ADD_95_U65 | ~new_U3018;
  assign new_U4471 = ~new_U3071;
  assign new_U4472 = ~new_U3034 | ~new_U3077;
  assign new_U4473 = ~new_R1150_U129 | ~new_U4016;
  assign new_U4474 = ~new_R1117_U128 | ~new_U4018;
  assign new_U4475 = ~new_R1138_U125 | ~new_U4017;
  assign new_U4476 = ~new_R1192_U129 | ~new_U4014;
  assign new_U4477 = ~new_R1207_U129 | ~new_U4013;
  assign new_U4478 = ~new_R1171_U125 | ~new_U4024;
  assign new_U4479 = ~new_R1240_U125 | ~new_U4022;
  assign new_U4480 = ~new_U3390;
  assign new_U4481 = ~new_R1222_U121 | ~new_U3027;
  assign new_U4482 = ~new_U3026 | ~new_U3071;
  assign new_U4483 = ~new_R1282_U84 | ~new_U3024;
  assign new_U4484 = ~new_U3494 | ~new_U4021;
  assign new_U4485 = ~new_U3717 | ~new_U4480;
  assign new_U4486 = ~REG2_REG_16_ | ~new_U3019;
  assign new_U4487 = ~REG1_REG_16_ | ~new_U3020;
  assign new_U4488 = ~REG0_REG_16_ | ~new_U3021;
  assign new_U4489 = ~new_ADD_95_U64 | ~new_U3018;
  assign new_U4490 = ~new_U3070;
  assign new_U4491 = ~new_U3034 | ~new_U3076;
  assign new_U4492 = ~new_R1150_U128 | ~new_U4016;
  assign new_U4493 = ~new_R1117_U127 | ~new_U4018;
  assign new_U4494 = ~new_R1138_U124 | ~new_U4017;
  assign new_U4495 = ~new_R1192_U128 | ~new_U4014;
  assign new_U4496 = ~new_R1207_U128 | ~new_U4013;
  assign new_U4497 = ~new_R1171_U124 | ~new_U4024;
  assign new_U4498 = ~new_R1240_U124 | ~new_U4022;
  assign new_U4499 = ~new_U3391;
  assign new_U4500 = ~new_R1222_U120 | ~new_U3027;
  assign new_U4501 = ~new_U3026 | ~new_U3070;
  assign new_U4502 = ~new_R1282_U81 | ~new_U3024;
  assign new_U4503 = ~new_U3496 | ~new_U4021;
  assign new_U4504 = ~new_U3721 | ~new_U4499;
  assign new_U4505 = ~REG2_REG_17_ | ~new_U3019;
  assign new_U4506 = ~REG1_REG_17_ | ~new_U3020;
  assign new_U4507 = ~REG0_REG_17_ | ~new_U3021;
  assign new_U4508 = ~new_ADD_95_U63 | ~new_U3018;
  assign new_U4509 = ~new_U3066;
  assign new_U4510 = ~new_U3034 | ~new_U3071;
  assign new_U4511 = ~new_R1150_U24 | ~new_U4016;
  assign new_U4512 = ~new_R1117_U24 | ~new_U4018;
  assign new_U4513 = ~new_R1138_U123 | ~new_U4017;
  assign new_U4514 = ~new_R1192_U25 | ~new_U4014;
  assign new_U4515 = ~new_R1207_U25 | ~new_U4013;
  assign new_U4516 = ~new_R1171_U123 | ~new_U4024;
  assign new_U4517 = ~new_R1240_U123 | ~new_U4022;
  assign new_U4518 = ~new_U3392;
  assign new_U4519 = ~new_R1222_U119 | ~new_U3027;
  assign new_U4520 = ~new_U3026 | ~new_U3066;
  assign new_U4521 = ~new_R1282_U79 | ~new_U3024;
  assign new_U4522 = ~new_U3498 | ~new_U4021;
  assign new_U4523 = ~new_U3725 | ~new_U4518;
  assign new_U4524 = ~REG2_REG_18_ | ~new_U3019;
  assign new_U4525 = ~REG1_REG_18_ | ~new_U3020;
  assign new_U4526 = ~REG0_REG_18_ | ~new_U3021;
  assign new_U4527 = ~new_ADD_95_U62 | ~new_U3018;
  assign new_U4528 = ~new_U3079;
  assign new_U4529 = ~new_U3034 | ~new_U3070;
  assign new_U4530 = ~new_R1150_U117 | ~new_U4016;
  assign new_U4531 = ~new_R1117_U116 | ~new_U4018;
  assign new_U4532 = ~new_R1138_U20 | ~new_U4017;
  assign new_U4533 = ~new_R1192_U117 | ~new_U4014;
  assign new_U4534 = ~new_R1207_U117 | ~new_U4013;
  assign new_U4535 = ~new_R1171_U20 | ~new_U4024;
  assign new_U4536 = ~new_R1240_U20 | ~new_U4022;
  assign new_U4537 = ~new_U3393;
  assign new_U4538 = ~new_R1222_U19 | ~new_U3027;
  assign new_U4539 = ~new_U3026 | ~new_U3079;
  assign new_U4540 = ~new_R1282_U76 | ~new_U3024;
  assign new_U4541 = ~new_U3500 | ~new_U4021;
  assign new_U4542 = ~new_U3729 | ~new_U4537;
  assign new_U4543 = ~REG2_REG_19_ | ~new_U3019;
  assign new_U4544 = ~REG1_REG_19_ | ~new_U3020;
  assign new_U4545 = ~REG0_REG_19_ | ~new_U3021;
  assign new_U4546 = ~new_ADD_95_U61 | ~new_U3018;
  assign new_U4547 = ~new_U3078;
  assign new_U4548 = ~new_U3034 | ~new_U3066;
  assign new_U4549 = ~new_R1150_U116 | ~new_U4016;
  assign new_U4550 = ~new_R1117_U115 | ~new_U4018;
  assign new_U4551 = ~new_R1138_U122 | ~new_U4017;
  assign new_U4552 = ~new_R1192_U116 | ~new_U4014;
  assign new_U4553 = ~new_R1207_U116 | ~new_U4013;
  assign new_U4554 = ~new_R1171_U122 | ~new_U4024;
  assign new_U4555 = ~new_R1240_U122 | ~new_U4022;
  assign new_U4556 = ~new_U3394;
  assign new_U4557 = ~new_R1222_U118 | ~new_U3027;
  assign new_U4558 = ~new_U3026 | ~new_U3078;
  assign new_U4559 = ~new_R1282_U74 | ~new_U3024;
  assign new_U4560 = ~new_U3502 | ~new_U4021;
  assign new_U4561 = ~new_U3733 | ~new_U4556;
  assign new_U4562 = ~REG2_REG_20_ | ~new_U3019;
  assign new_U4563 = ~REG1_REG_20_ | ~new_U3020;
  assign new_U4564 = ~REG0_REG_20_ | ~new_U3021;
  assign new_U4565 = ~new_ADD_95_U60 | ~new_U3018;
  assign new_U4566 = ~new_U3073;
  assign new_U4567 = ~new_U3034 | ~new_U3079;
  assign new_U4568 = ~new_R1150_U115 | ~new_U4016;
  assign new_U4569 = ~new_R1117_U114 | ~new_U4018;
  assign new_U4570 = ~new_R1138_U121 | ~new_U4017;
  assign new_U4571 = ~new_R1192_U115 | ~new_U4014;
  assign new_U4572 = ~new_R1207_U115 | ~new_U4013;
  assign new_U4573 = ~new_R1171_U121 | ~new_U4024;
  assign new_U4574 = ~new_R1240_U121 | ~new_U4022;
  assign new_U4575 = ~new_U3395;
  assign new_U4576 = ~new_R1222_U117 | ~new_U3027;
  assign new_U4577 = ~new_U3026 | ~new_U3073;
  assign new_U4578 = ~new_R1282_U71 | ~new_U3024;
  assign new_U4579 = ~new_U3504 | ~new_U4021;
  assign new_U4580 = ~new_U3737 | ~new_U4575;
  assign new_U4581 = ~REG2_REG_21_ | ~new_U3019;
  assign new_U4582 = ~REG1_REG_21_ | ~new_U3020;
  assign new_U4583 = ~REG0_REG_21_ | ~new_U3021;
  assign new_U4584 = ~new_ADD_95_U59 | ~new_U3018;
  assign new_U4585 = ~new_U3072;
  assign new_U4586 = ~new_U3034 | ~new_U3078;
  assign new_U4587 = ~new_R1150_U113 | ~new_U4016;
  assign new_U4588 = ~new_R1117_U112 | ~new_U4018;
  assign new_U4589 = ~new_R1138_U21 | ~new_U4017;
  assign new_U4590 = ~new_R1192_U113 | ~new_U4014;
  assign new_U4591 = ~new_R1207_U113 | ~new_U4013;
  assign new_U4592 = ~new_R1171_U21 | ~new_U4024;
  assign new_U4593 = ~new_R1240_U21 | ~new_U4022;
  assign new_U4594 = ~new_U3397;
  assign new_U4595 = ~new_R1222_U20 | ~new_U3027;
  assign new_U4596 = ~new_U3026 | ~new_U3072;
  assign new_U4597 = ~new_R1282_U67 | ~new_U3024;
  assign new_U4598 = ~new_U4037 | ~new_U4021;
  assign new_U4599 = ~new_U3741 | ~new_U4594;
  assign new_U4600 = ~REG2_REG_22_ | ~new_U3019;
  assign new_U4601 = ~REG1_REG_22_ | ~new_U3020;
  assign new_U4602 = ~REG0_REG_22_ | ~new_U3021;
  assign new_U4603 = ~new_ADD_95_U58 | ~new_U3018;
  assign new_U4604 = ~new_U3058;
  assign new_U4605 = ~new_U3034 | ~new_U3073;
  assign new_U4606 = ~new_R1150_U127 | ~new_U4016;
  assign new_U4607 = ~new_R1117_U126 | ~new_U4018;
  assign new_U4608 = ~new_R1138_U22 | ~new_U4017;
  assign new_U4609 = ~new_R1192_U127 | ~new_U4014;
  assign new_U4610 = ~new_R1207_U127 | ~new_U4013;
  assign new_U4611 = ~new_R1171_U22 | ~new_U4024;
  assign new_U4612 = ~new_R1240_U22 | ~new_U4022;
  assign new_U4613 = ~new_U3399;
  assign new_U4614 = ~new_R1222_U21 | ~new_U3027;
  assign new_U4615 = ~new_U3026 | ~new_U3058;
  assign new_U4616 = ~new_R1282_U64 | ~new_U3024;
  assign new_U4617 = ~new_U4036 | ~new_U4021;
  assign new_U4618 = ~new_U3745 | ~new_U4613;
  assign new_U4619 = ~REG2_REG_23_ | ~new_U3019;
  assign new_U4620 = ~REG1_REG_23_ | ~new_U3020;
  assign new_U4621 = ~REG0_REG_23_ | ~new_U3021;
  assign new_U4622 = ~new_ADD_95_U57 | ~new_U3018;
  assign new_U4623 = ~new_U3063;
  assign new_U4624 = ~new_U3034 | ~new_U3072;
  assign new_U4625 = ~new_R1150_U126 | ~new_U4016;
  assign new_U4626 = ~new_R1117_U125 | ~new_U4018;
  assign new_U4627 = ~new_R1138_U120 | ~new_U4017;
  assign new_U4628 = ~new_R1192_U126 | ~new_U4014;
  assign new_U4629 = ~new_R1207_U126 | ~new_U4013;
  assign new_U4630 = ~new_R1171_U120 | ~new_U4024;
  assign new_U4631 = ~new_R1240_U120 | ~new_U4022;
  assign new_U4632 = ~new_U3401;
  assign new_U4633 = ~new_R1222_U116 | ~new_U3027;
  assign new_U4634 = ~new_U3026 | ~new_U3063;
  assign new_U4635 = ~new_R1282_U62 | ~new_U3024;
  assign new_U4636 = ~new_U4035 | ~new_U4021;
  assign new_U4637 = ~new_U3749 | ~new_U4632;
  assign new_U4638 = ~REG2_REG_24_ | ~new_U3019;
  assign new_U4639 = ~REG1_REG_24_ | ~new_U3020;
  assign new_U4640 = ~REG0_REG_24_ | ~new_U3021;
  assign new_U4641 = ~new_ADD_95_U56 | ~new_U3018;
  assign new_U4642 = ~new_U3062;
  assign new_U4643 = ~new_U3034 | ~new_U3058;
  assign new_U4644 = ~new_R1150_U25 | ~new_U4016;
  assign new_U4645 = ~new_R1117_U25 | ~new_U4018;
  assign new_U4646 = ~new_R1138_U119 | ~new_U4017;
  assign new_U4647 = ~new_R1192_U26 | ~new_U4014;
  assign new_U4648 = ~new_R1207_U26 | ~new_U4013;
  assign new_U4649 = ~new_R1171_U119 | ~new_U4024;
  assign new_U4650 = ~new_R1240_U119 | ~new_U4022;
  assign new_U4651 = ~new_U3403;
  assign new_U4652 = ~new_R1222_U115 | ~new_U3027;
  assign new_U4653 = ~new_U3026 | ~new_U3062;
  assign new_U4654 = ~new_R1282_U59 | ~new_U3024;
  assign new_U4655 = ~new_U4034 | ~new_U4021;
  assign new_U4656 = ~new_U3753 | ~new_U4651;
  assign new_U4657 = ~REG2_REG_25_ | ~new_U3019;
  assign new_U4658 = ~REG1_REG_25_ | ~new_U3020;
  assign new_U4659 = ~REG0_REG_25_ | ~new_U3021;
  assign new_U4660 = ~new_ADD_95_U55 | ~new_U3018;
  assign new_U4661 = ~new_U3055;
  assign new_U4662 = ~new_U3034 | ~new_U3063;
  assign new_U4663 = ~new_R1150_U112 | ~new_U4016;
  assign new_U4664 = ~new_R1117_U111 | ~new_U4018;
  assign new_U4665 = ~new_R1138_U118 | ~new_U4017;
  assign new_U4666 = ~new_R1192_U112 | ~new_U4014;
  assign new_U4667 = ~new_R1207_U112 | ~new_U4013;
  assign new_U4668 = ~new_R1171_U118 | ~new_U4024;
  assign new_U4669 = ~new_R1240_U118 | ~new_U4022;
  assign new_U4670 = ~new_U3405;
  assign new_U4671 = ~new_R1222_U114 | ~new_U3027;
  assign new_U4672 = ~new_U3026 | ~new_U3055;
  assign new_U4673 = ~new_R1282_U57 | ~new_U3024;
  assign new_U4674 = ~new_U4033 | ~new_U4021;
  assign new_U4675 = ~new_U3757 | ~new_U4670;
  assign new_U4676 = ~REG2_REG_26_ | ~new_U3019;
  assign new_U4677 = ~REG1_REG_26_ | ~new_U3020;
  assign new_U4678 = ~REG0_REG_26_ | ~new_U3021;
  assign new_U4679 = ~new_ADD_95_U54 | ~new_U3018;
  assign new_U4680 = ~new_U3054;
  assign new_U4681 = ~new_U3034 | ~new_U3062;
  assign new_U4682 = ~new_R1150_U111 | ~new_U4016;
  assign new_U4683 = ~new_R1117_U110 | ~new_U4018;
  assign new_U4684 = ~new_R1138_U117 | ~new_U4017;
  assign new_U4685 = ~new_R1192_U111 | ~new_U4014;
  assign new_U4686 = ~new_R1207_U111 | ~new_U4013;
  assign new_U4687 = ~new_R1171_U117 | ~new_U4024;
  assign new_U4688 = ~new_R1240_U117 | ~new_U4022;
  assign new_U4689 = ~new_U3407;
  assign new_U4690 = ~new_R1222_U113 | ~new_U3027;
  assign new_U4691 = ~new_U3026 | ~new_U3054;
  assign new_U4692 = ~new_R1282_U54 | ~new_U3024;
  assign new_U4693 = ~new_U4032 | ~new_U4021;
  assign new_U4694 = ~new_U3761 | ~new_U4689;
  assign new_U4695 = ~REG2_REG_27_ | ~new_U3019;
  assign new_U4696 = ~REG1_REG_27_ | ~new_U3020;
  assign new_U4697 = ~REG0_REG_27_ | ~new_U3021;
  assign new_U4698 = ~new_ADD_95_U53 | ~new_U3018;
  assign new_U4699 = ~new_U3050;
  assign new_U4700 = ~new_U3034 | ~new_U3055;
  assign new_U4701 = ~new_R1150_U125 | ~new_U4016;
  assign new_U4702 = ~new_R1117_U124 | ~new_U4018;
  assign new_U4703 = ~new_R1138_U23 | ~new_U4017;
  assign new_U4704 = ~new_R1192_U125 | ~new_U4014;
  assign new_U4705 = ~new_R1207_U125 | ~new_U4013;
  assign new_U4706 = ~new_R1171_U23 | ~new_U4024;
  assign new_U4707 = ~new_R1240_U23 | ~new_U4022;
  assign new_U4708 = ~new_U3409;
  assign new_U4709 = ~new_R1222_U22 | ~new_U3027;
  assign new_U4710 = ~new_U3026 | ~new_U3050;
  assign new_U4711 = ~new_R1282_U52 | ~new_U3024;
  assign new_U4712 = ~new_U4031 | ~new_U4021;
  assign new_U4713 = ~new_U3765 | ~new_U4708;
  assign new_U4714 = ~REG2_REG_28_ | ~new_U3019;
  assign new_U4715 = ~REG1_REG_28_ | ~new_U3020;
  assign new_U4716 = ~REG0_REG_28_ | ~new_U3021;
  assign new_U4717 = ~new_ADD_95_U52 | ~new_U3018;
  assign new_U4718 = ~new_U3051;
  assign new_U4719 = ~new_U3034 | ~new_U3054;
  assign new_U4720 = ~new_R1150_U26 | ~new_U4016;
  assign new_U4721 = ~new_R1117_U31 | ~new_U4018;
  assign new_U4722 = ~new_R1138_U116 | ~new_U4017;
  assign new_U4723 = ~new_R1192_U27 | ~new_U4014;
  assign new_U4724 = ~new_R1207_U27 | ~new_U4013;
  assign new_U4725 = ~new_R1171_U116 | ~new_U4024;
  assign new_U4726 = ~new_R1240_U116 | ~new_U4022;
  assign new_U4727 = ~new_U3411;
  assign new_U4728 = ~new_R1222_U112 | ~new_U3027;
  assign new_U4729 = ~new_U3026 | ~new_U3051;
  assign new_U4730 = ~new_R1282_U49 | ~new_U3024;
  assign new_U4731 = ~new_U4030 | ~new_U4021;
  assign new_U4732 = ~new_U3769 | ~new_U4727;
  assign new_U4733 = ~new_ADD_95_U5 | ~new_U3018;
  assign new_U4734 = ~REG2_REG_29_ | ~new_U3019;
  assign new_U4735 = ~REG1_REG_29_ | ~new_U3020;
  assign new_U4736 = ~REG0_REG_29_ | ~new_U3021;
  assign new_U4737 = ~new_U3052;
  assign new_U4738 = ~new_U3034 | ~new_U3050;
  assign new_U4739 = ~new_R1150_U110 | ~new_U4016;
  assign new_U4740 = ~new_R1117_U109 | ~new_U4018;
  assign new_U4741 = ~new_R1138_U115 | ~new_U4017;
  assign new_U4742 = ~new_R1192_U110 | ~new_U4014;
  assign new_U4743 = ~new_R1207_U110 | ~new_U4013;
  assign new_U4744 = ~new_R1171_U115 | ~new_U4024;
  assign new_U4745 = ~new_R1240_U115 | ~new_U4022;
  assign new_U4746 = ~new_U3413;
  assign new_U4747 = ~new_R1222_U111 | ~new_U3027;
  assign new_U4748 = ~new_U3026 | ~new_U3052;
  assign new_U4749 = ~new_R1282_U47 | ~new_U3024;
  assign new_U4750 = ~new_U4029 | ~new_U4021;
  assign new_U4751 = ~new_U3773 | ~new_U4746;
  assign new_U4752 = ~REG2_REG_30_ | ~new_U3019;
  assign new_U4753 = ~REG1_REG_30_ | ~new_U3020;
  assign new_U4754 = ~REG0_REG_30_ | ~new_U3021;
  assign new_U4755 = ~new_U3056;
  assign new_U4756 = ~new_U5799 | ~new_U3359;
  assign new_U4757 = ~new_U3969 | ~new_U4756;
  assign new_U4758 = ~new_U3774 | ~new_U3056;
  assign new_U4759 = ~new_U3034 | ~new_U3051;
  assign new_U4760 = ~new_R1150_U27 | ~new_U4016;
  assign new_U4761 = ~new_R1117_U26 | ~new_U4018;
  assign new_U4762 = ~new_R1138_U114 | ~new_U4017;
  assign new_U4763 = ~new_R1192_U28 | ~new_U4014;
  assign new_U4764 = ~new_R1207_U28 | ~new_U4013;
  assign new_U4765 = ~new_R1171_U114 | ~new_U4024;
  assign new_U4766 = ~new_R1240_U114 | ~new_U4022;
  assign new_U4767 = ~new_U3838 | ~new_U3049 | ~new_U5740;
  assign new_U4768 = ~new_R1222_U110 | ~new_U3027;
  assign new_U4769 = ~new_R1282_U44 | ~new_U3024;
  assign new_U4770 = ~new_U4040 | ~new_U4021;
  assign new_U4771 = ~new_U3775 | ~new_U3776 | ~new_U3049;
  assign new_U4772 = ~REG2_REG_31_ | ~new_U3019;
  assign new_U4773 = ~REG1_REG_31_ | ~new_U3020;
  assign new_U4774 = ~REG0_REG_31_ | ~new_U3021;
  assign new_U4775 = ~new_U3053;
  assign new_U4776 = ~new_R1282_U42 | ~new_U3024;
  assign new_U4777 = ~new_U4039 | ~new_U4021;
  assign new_U4778 = ~new_U4776 | ~new_U4777 | ~new_U4002;
  assign new_U4779 = ~new_R1282_U39 | ~new_U3024;
  assign new_U4780 = ~new_U4038 | ~new_U4021;
  assign new_U4781 = ~new_U4779 | ~new_U4780 | ~new_U4002;
  assign new_U4782 = ~new_U5820 | ~new_U5817;
  assign new_U4783 = ~new_U3779 | ~new_U3017;
  assign new_U4784 = ~new_U3418 | ~new_U4783;
  assign new_U4785 = ~new_U3036 | ~new_U3075;
  assign new_U4786 = ~new_U3033 | ~REG3_REG_0_;
  assign new_U4787 = ~new_U3032 | ~new_R1222_U104;
  assign new_U4788 = ~new_U3031 | ~new_U3464;
  assign new_U4789 = ~new_U3030 | ~new_U3464;
  assign new_U4790 = ~new_U3036 | ~new_U3065;
  assign new_U4791 = ~new_U3033 | ~REG3_REG_1_;
  assign new_U4792 = ~new_U3032 | ~new_R1222_U103;
  assign new_U4793 = ~new_U3031 | ~new_U3468;
  assign new_U4794 = ~new_U3030 | ~new_R1282_U31;
  assign new_U4795 = ~new_U3036 | ~new_U3061;
  assign new_U4796 = ~new_U3033 | ~REG3_REG_2_;
  assign new_U4797 = ~new_U3032 | ~new_R1222_U23;
  assign new_U4798 = ~new_U3031 | ~new_U3470;
  assign new_U4799 = ~new_U3030 | ~new_R1282_U6;
  assign new_U4800 = ~new_U3036 | ~new_U3057;
  assign new_U4801 = ~new_U3033 | ~new_ADD_95_U4;
  assign new_U4802 = ~new_U3032 | ~new_R1222_U109;
  assign new_U4803 = ~new_U3031 | ~new_U3472;
  assign new_U4804 = ~new_U3030 | ~new_R1282_U7;
  assign new_U4805 = ~new_U3036 | ~new_U3064;
  assign new_U4806 = ~new_U3033 | ~new_ADD_95_U51;
  assign new_U4807 = ~new_U3032 | ~new_R1222_U108;
  assign new_U4808 = ~new_U3031 | ~new_U3474;
  assign new_U4809 = ~new_U3030 | ~new_R1282_U8;
  assign new_U4810 = ~new_U3036 | ~new_U3068;
  assign new_U4811 = ~new_U3033 | ~new_ADD_95_U50;
  assign new_U4812 = ~new_U3032 | ~new_R1222_U24;
  assign new_U4813 = ~new_U3031 | ~new_U3476;
  assign new_U4814 = ~new_U3030 | ~new_R1282_U9;
  assign new_U4815 = ~new_U3036 | ~new_U3067;
  assign new_U4816 = ~new_U3033 | ~new_ADD_95_U49;
  assign new_U4817 = ~new_U3032 | ~new_R1222_U107;
  assign new_U4818 = ~new_U3031 | ~new_U3478;
  assign new_U4819 = ~new_U3030 | ~new_R1282_U10;
  assign new_U4820 = ~new_U3036 | ~new_U3081;
  assign new_U4821 = ~new_U3033 | ~new_ADD_95_U48;
  assign new_U4822 = ~new_U3032 | ~new_R1222_U25;
  assign new_U4823 = ~new_U3031 | ~new_U3480;
  assign new_U4824 = ~new_U3030 | ~new_R1282_U11;
  assign new_U4825 = ~new_U3036 | ~new_U3080;
  assign new_U4826 = ~new_U3033 | ~new_ADD_95_U47;
  assign new_U4827 = ~new_U3032 | ~new_R1222_U106;
  assign new_U4828 = ~new_U3031 | ~new_U3482;
  assign new_U4829 = ~new_U3030 | ~new_R1282_U36;
  assign new_U4830 = ~new_U3036 | ~new_U3059;
  assign new_U4831 = ~new_U3033 | ~new_ADD_95_U46;
  assign new_U4832 = ~new_U3032 | ~new_R1222_U105;
  assign new_U4833 = ~new_U3031 | ~new_U3484;
  assign new_U4834 = ~new_U3030 | ~new_R1282_U33;
  assign new_U4835 = ~new_U3036 | ~new_U3060;
  assign new_U4836 = ~new_U3033 | ~new_ADD_95_U70;
  assign new_U4837 = ~new_U3032 | ~new_R1222_U17;
  assign new_U4838 = ~new_U3031 | ~new_U3486;
  assign new_U4839 = ~new_U3030 | ~new_R1282_U94;
  assign new_U4840 = ~new_U3036 | ~new_U3069;
  assign new_U4841 = ~new_U3033 | ~new_ADD_95_U69;
  assign new_U4842 = ~new_U3032 | ~new_R1222_U123;
  assign new_U4843 = ~new_U3031 | ~new_U3488;
  assign new_U4844 = ~new_U3030 | ~new_R1282_U91;
  assign new_U4845 = ~new_U3036 | ~new_U3077;
  assign new_U4846 = ~new_U3033 | ~new_ADD_95_U68;
  assign new_U4847 = ~new_U3032 | ~new_R1222_U122;
  assign new_U4848 = ~new_U3031 | ~new_U3490;
  assign new_U4849 = ~new_U3030 | ~new_R1282_U89;
  assign new_U4850 = ~new_U3036 | ~new_U3076;
  assign new_U4851 = ~new_U3033 | ~new_ADD_95_U67;
  assign new_U4852 = ~new_U3032 | ~new_R1222_U18;
  assign new_U4853 = ~new_U3031 | ~new_U3492;
  assign new_U4854 = ~new_U3030 | ~new_R1282_U86;
  assign new_U4855 = ~new_U3036 | ~new_U3071;
  assign new_U4856 = ~new_U3033 | ~new_ADD_95_U66;
  assign new_U4857 = ~new_U3032 | ~new_R1222_U121;
  assign new_U4858 = ~new_U3031 | ~new_U3494;
  assign new_U4859 = ~new_U3030 | ~new_R1282_U84;
  assign new_U4860 = ~new_U3036 | ~new_U3070;
  assign new_U4861 = ~new_U3033 | ~new_ADD_95_U65;
  assign new_U4862 = ~new_U3032 | ~new_R1222_U120;
  assign new_U4863 = ~new_U3031 | ~new_U3496;
  assign new_U4864 = ~new_U3030 | ~new_R1282_U81;
  assign new_U4865 = ~new_U3036 | ~new_U3066;
  assign new_U4866 = ~new_U3033 | ~new_ADD_95_U64;
  assign new_U4867 = ~new_U3032 | ~new_R1222_U119;
  assign new_U4868 = ~new_U3031 | ~new_U3498;
  assign new_U4869 = ~new_U3030 | ~new_R1282_U79;
  assign new_U4870 = ~new_U3036 | ~new_U3079;
  assign new_U4871 = ~new_U3033 | ~new_ADD_95_U63;
  assign new_U4872 = ~new_U3032 | ~new_R1222_U19;
  assign new_U4873 = ~new_U3031 | ~new_U3500;
  assign new_U4874 = ~new_U3030 | ~new_R1282_U76;
  assign new_U4875 = ~new_U3036 | ~new_U3078;
  assign new_U4876 = ~new_U3033 | ~new_ADD_95_U62;
  assign new_U4877 = ~new_U3032 | ~new_R1222_U118;
  assign new_U4878 = ~new_U3031 | ~new_U3502;
  assign new_U4879 = ~new_U3030 | ~new_R1282_U74;
  assign new_U4880 = ~new_U3036 | ~new_U3073;
  assign new_U4881 = ~new_U3033 | ~new_ADD_95_U61;
  assign new_U4882 = ~new_U3032 | ~new_R1222_U117;
  assign new_U4883 = ~new_U3031 | ~new_U3504;
  assign new_U4884 = ~new_U3030 | ~new_R1282_U71;
  assign new_U4885 = ~new_U3036 | ~new_U3072;
  assign new_U4886 = ~new_U3033 | ~new_ADD_95_U60;
  assign new_U4887 = ~new_U3032 | ~new_R1222_U20;
  assign new_U4888 = ~new_U3031 | ~new_U4037;
  assign new_U4889 = ~new_U3030 | ~new_R1282_U67;
  assign new_U4890 = ~new_U3036 | ~new_U3058;
  assign new_U4891 = ~new_U3033 | ~new_ADD_95_U59;
  assign new_U4892 = ~new_U3032 | ~new_R1222_U21;
  assign new_U4893 = ~new_U3031 | ~new_U4036;
  assign new_U4894 = ~new_U3030 | ~new_R1282_U64;
  assign new_U4895 = ~new_U3036 | ~new_U3063;
  assign new_U4896 = ~new_U3033 | ~new_ADD_95_U58;
  assign new_U4897 = ~new_U3032 | ~new_R1222_U116;
  assign new_U4898 = ~new_U3031 | ~new_U4035;
  assign new_U4899 = ~new_U3030 | ~new_R1282_U62;
  assign new_U4900 = ~new_U3036 | ~new_U3062;
  assign new_U4901 = ~new_U3033 | ~new_ADD_95_U57;
  assign new_U4902 = ~new_U3032 | ~new_R1222_U115;
  assign new_U4903 = ~new_U3031 | ~new_U4034;
  assign new_U4904 = ~new_U3030 | ~new_R1282_U59;
  assign new_U4905 = ~new_U3036 | ~new_U3055;
  assign new_U4906 = ~new_U3033 | ~new_ADD_95_U56;
  assign new_U4907 = ~new_U3032 | ~new_R1222_U114;
  assign new_U4908 = ~new_U3031 | ~new_U4033;
  assign new_U4909 = ~new_U3030 | ~new_R1282_U57;
  assign new_U4910 = ~new_U3036 | ~new_U3054;
  assign new_U4911 = ~new_U3033 | ~new_ADD_95_U55;
  assign new_U4912 = ~new_U3032 | ~new_R1222_U113;
  assign new_U4913 = ~new_U3031 | ~new_U4032;
  assign new_U4914 = ~new_U3030 | ~new_R1282_U54;
  assign new_U4915 = ~new_U3036 | ~new_U3050;
  assign new_U4916 = ~new_U3033 | ~new_ADD_95_U54;
  assign new_U4917 = ~new_U3032 | ~new_R1222_U22;
  assign new_U4918 = ~new_U3031 | ~new_U4031;
  assign new_U4919 = ~new_U3030 | ~new_R1282_U52;
  assign new_U4920 = ~new_U3036 | ~new_U3051;
  assign new_U4921 = ~new_U3033 | ~new_ADD_95_U53;
  assign new_U4922 = ~new_U3032 | ~new_R1222_U112;
  assign new_U4923 = ~new_U3031 | ~new_U4030;
  assign new_U4924 = ~new_U3030 | ~new_R1282_U49;
  assign new_U4925 = ~new_U3036 | ~new_U3052;
  assign new_U4926 = ~new_U3033 | ~new_ADD_95_U52;
  assign new_U4927 = ~new_U3032 | ~new_R1222_U111;
  assign new_U4928 = ~new_U3031 | ~new_U4029;
  assign new_U4929 = ~new_U3030 | ~new_R1282_U47;
  assign new_U4930 = ~new_U3033 | ~new_ADD_95_U5;
  assign new_U4931 = ~new_U3032 | ~new_R1222_U110;
  assign new_U4932 = ~new_U3031 | ~new_U4040;
  assign new_U4933 = ~new_U3030 | ~new_R1282_U44;
  assign new_U4934 = ~new_U3031 | ~new_U4039;
  assign new_U4935 = ~new_U3030 | ~new_R1282_U42;
  assign new_U4936 = ~new_U3031 | ~new_U4038;
  assign new_U4937 = ~new_U3030 | ~new_R1282_U39;
  assign new_U4938 = ~new_U3839 | ~new_U3840 | ~new_U3843 | ~new_U3842;
  assign new_U4939 = ~new_R1105_U4 | ~new_U3042 | ~new_U3044;
  assign new_U4940 = ~new_U3844 | ~new_U3044;
  assign new_U4941 = ~new_R1162_U4 | ~new_U3038 | ~new_U3044;
  assign new_U4942 = ~new_U3421;
  assign new_U4943 = ~new_U3043 | ~new_R1105_U4;
  assign new_U4944 = ~REG3_REG_19_ | ~n1342;
  assign new_U4945 = ~new_U3041 | ~new_U3461;
  assign new_U4946 = ~new_U3039 | ~new_R1162_U4;
  assign new_U4947 = ~ADDR_REG_19_ | ~new_U4942;
  assign new_U4948 = ~new_R1105_U55 | ~new_U3042 | ~new_U3044;
  assign new_U4949 = ~new_U3849 | ~new_U3044;
  assign new_U4950 = ~new_R1162_U62 | ~new_U3038 | ~new_U3044;
  assign new_U4951 = ~new_R1105_U55 | ~new_U3043;
  assign new_U4952 = ~REG3_REG_18_ | ~n1342;
  assign new_U4953 = ~new_U3041 | ~new_U3444;
  assign new_U4954 = ~new_R1162_U62 | ~new_U3039;
  assign new_U4955 = ~ADDR_REG_18_ | ~new_U4942;
  assign new_U4956 = ~new_R1105_U56 | ~new_U3042;
  assign new_U4957 = ~new_U3040 | ~new_U3445;
  assign new_U4958 = ~new_R1162_U63 | ~new_U3038;
  assign new_U4959 = ~new_U4958 | ~new_U4957 | ~new_U4956;
  assign new_U4960 = ~new_U3044 | ~new_U4959;
  assign new_U4961 = ~new_R1105_U56 | ~new_U3043;
  assign new_U4962 = ~REG3_REG_17_ | ~n1342;
  assign new_U4963 = ~new_U3041 | ~new_U3445;
  assign new_U4964 = ~new_R1162_U63 | ~new_U3039;
  assign new_U4965 = ~ADDR_REG_17_ | ~new_U4942;
  assign new_U4966 = ~new_R1105_U57 | ~new_U3042;
  assign new_U4967 = ~new_U3040 | ~new_U3446;
  assign new_U4968 = ~new_R1162_U64 | ~new_U3038;
  assign new_U4969 = ~new_U4968 | ~new_U4967 | ~new_U4966;
  assign new_U4970 = ~new_U3044 | ~new_U4969;
  assign new_U4971 = ~new_R1105_U57 | ~new_U3043;
  assign new_U4972 = ~REG3_REG_16_ | ~n1342;
  assign new_U4973 = ~new_U3041 | ~new_U3446;
  assign new_U4974 = ~new_R1162_U64 | ~new_U3039;
  assign new_U4975 = ~ADDR_REG_16_ | ~new_U4942;
  assign new_U4976 = ~new_R1105_U58 | ~new_U3042;
  assign new_U4977 = ~new_U3040 | ~new_U3447;
  assign new_U4978 = ~new_R1162_U65 | ~new_U3038;
  assign new_U4979 = ~new_U4978 | ~new_U4977 | ~new_U4976;
  assign new_U4980 = ~new_U3044 | ~new_U4979;
  assign new_U4981 = ~new_R1105_U58 | ~new_U3043;
  assign new_U4982 = ~REG3_REG_15_ | ~n1342;
  assign new_U4983 = ~new_U3041 | ~new_U3447;
  assign new_U4984 = ~new_R1162_U65 | ~new_U3039;
  assign new_U4985 = ~ADDR_REG_15_ | ~new_U4942;
  assign new_U4986 = ~new_R1105_U59 | ~new_U3042;
  assign new_U4987 = ~new_U3040 | ~new_U3448;
  assign new_U4988 = ~new_R1162_U66 | ~new_U3038;
  assign new_U4989 = ~new_U4988 | ~new_U4987 | ~new_U4986;
  assign new_U4990 = ~new_U3044 | ~new_U4989;
  assign new_U4991 = ~new_R1105_U59 | ~new_U3043;
  assign new_U4992 = ~REG3_REG_14_ | ~n1342;
  assign new_U4993 = ~new_U3041 | ~new_U3448;
  assign new_U4994 = ~new_R1162_U66 | ~new_U3039;
  assign new_U4995 = ~ADDR_REG_14_ | ~new_U4942;
  assign new_U4996 = ~new_R1105_U60 | ~new_U3042;
  assign new_U4997 = ~new_U3040 | ~new_U3449;
  assign new_U4998 = ~new_R1162_U67 | ~new_U3038;
  assign new_U4999 = ~new_U4998 | ~new_U4997 | ~new_U4996;
  assign new_U5000 = ~new_U3044 | ~new_U4999;
  assign new_U5001 = ~new_R1105_U60 | ~new_U3043;
  assign new_U5002 = ~REG3_REG_13_ | ~n1342;
  assign new_U5003 = ~new_U3041 | ~new_U3449;
  assign new_U5004 = ~new_R1162_U67 | ~new_U3039;
  assign new_U5005 = ~ADDR_REG_13_ | ~new_U4942;
  assign new_U5006 = ~new_R1105_U61 | ~new_U3042;
  assign new_U5007 = ~new_U3040 | ~new_U3450;
  assign new_U5008 = ~new_R1162_U68 | ~new_U3038;
  assign new_U5009 = ~new_U5008 | ~new_U5007 | ~new_U5006;
  assign new_U5010 = ~new_U3044 | ~new_U5009;
  assign new_U5011 = ~new_R1105_U61 | ~new_U3043;
  assign new_U5012 = ~REG3_REG_12_ | ~n1342;
  assign new_U5013 = ~new_U3041 | ~new_U3450;
  assign new_U5014 = ~new_R1162_U68 | ~new_U3039;
  assign new_U5015 = ~ADDR_REG_12_ | ~new_U4942;
  assign new_U5016 = ~new_R1105_U62 | ~new_U3042;
  assign new_U5017 = ~new_U3040 | ~new_U3451;
  assign new_U5018 = ~new_R1162_U69 | ~new_U3038;
  assign new_U5019 = ~new_U5018 | ~new_U5017 | ~new_U5016;
  assign new_U5020 = ~new_U3044 | ~new_U5019;
  assign new_U5021 = ~new_R1105_U62 | ~new_U3043;
  assign new_U5022 = ~REG3_REG_11_ | ~n1342;
  assign new_U5023 = ~new_U3041 | ~new_U3451;
  assign new_U5024 = ~new_R1162_U69 | ~new_U3039;
  assign new_U5025 = ~ADDR_REG_11_ | ~new_U4942;
  assign new_U5026 = ~new_R1105_U63 | ~new_U3042;
  assign new_U5027 = ~new_U3040 | ~new_U3452;
  assign new_U5028 = ~new_R1162_U70 | ~new_U3038;
  assign new_U5029 = ~new_U5028 | ~new_U5027 | ~new_U5026;
  assign new_U5030 = ~new_U3044 | ~new_U5029;
  assign new_U5031 = ~new_R1105_U63 | ~new_U3043;
  assign new_U5032 = ~REG3_REG_10_ | ~n1342;
  assign new_U5033 = ~new_U3041 | ~new_U3452;
  assign new_U5034 = ~new_R1162_U70 | ~new_U3039;
  assign new_U5035 = ~ADDR_REG_10_ | ~new_U4942;
  assign new_U5036 = ~new_R1105_U47 | ~new_U3042;
  assign new_U5037 = ~new_U3040 | ~new_U3435;
  assign new_U5038 = ~new_R1162_U54 | ~new_U3038;
  assign new_U5039 = ~new_U5038 | ~new_U5037 | ~new_U5036;
  assign new_U5040 = ~new_U3044 | ~new_U5039;
  assign new_U5041 = ~new_R1105_U47 | ~new_U3043;
  assign new_U5042 = ~REG3_REG_9_ | ~n1342;
  assign new_U5043 = ~new_U3041 | ~new_U3435;
  assign new_U5044 = ~new_R1162_U54 | ~new_U3039;
  assign new_U5045 = ~ADDR_REG_9_ | ~new_U4942;
  assign new_U5046 = ~new_R1105_U48 | ~new_U3042;
  assign new_U5047 = ~new_U3040 | ~new_U3436;
  assign new_U5048 = ~new_R1162_U55 | ~new_U3038;
  assign new_U5049 = ~new_U5048 | ~new_U5047 | ~new_U5046;
  assign new_U5050 = ~new_U3044 | ~new_U5049;
  assign new_U5051 = ~new_R1105_U48 | ~new_U3043;
  assign new_U5052 = ~REG3_REG_8_ | ~n1342;
  assign new_U5053 = ~new_U3041 | ~new_U3436;
  assign new_U5054 = ~new_R1162_U55 | ~new_U3039;
  assign new_U5055 = ~ADDR_REG_8_ | ~new_U4942;
  assign new_U5056 = ~new_R1105_U49 | ~new_U3042;
  assign new_U5057 = ~new_U3040 | ~new_U3437;
  assign new_U5058 = ~new_R1162_U56 | ~new_U3038;
  assign new_U5059 = ~new_U5058 | ~new_U5057 | ~new_U5056;
  assign new_U5060 = ~new_U3044 | ~new_U5059;
  assign new_U5061 = ~new_R1105_U49 | ~new_U3043;
  assign new_U5062 = ~REG3_REG_7_ | ~n1342;
  assign new_U5063 = ~new_U3041 | ~new_U3437;
  assign new_U5064 = ~new_R1162_U56 | ~new_U3039;
  assign new_U5065 = ~ADDR_REG_7_ | ~new_U4942;
  assign new_U5066 = ~new_R1105_U50 | ~new_U3042;
  assign new_U5067 = ~new_U3040 | ~new_U3438;
  assign new_U5068 = ~new_R1162_U57 | ~new_U3038;
  assign new_U5069 = ~new_U5068 | ~new_U5067 | ~new_U5066;
  assign new_U5070 = ~new_U3044 | ~new_U5069;
  assign new_U5071 = ~new_R1105_U50 | ~new_U3043;
  assign new_U5072 = ~REG3_REG_6_ | ~n1342;
  assign new_U5073 = ~new_U3041 | ~new_U3438;
  assign new_U5074 = ~new_R1162_U57 | ~new_U3039;
  assign new_U5075 = ~ADDR_REG_6_ | ~new_U4942;
  assign new_U5076 = ~new_R1105_U51 | ~new_U3042;
  assign new_U5077 = ~new_U3040 | ~new_U3439;
  assign new_U5078 = ~new_R1162_U58 | ~new_U3038;
  assign new_U5079 = ~new_U5078 | ~new_U5077 | ~new_U5076;
  assign new_U5080 = ~new_U3044 | ~new_U5079;
  assign new_U5081 = ~new_R1105_U51 | ~new_U3043;
  assign new_U5082 = ~REG3_REG_5_ | ~n1342;
  assign new_U5083 = ~new_U3041 | ~new_U3439;
  assign new_U5084 = ~new_R1162_U58 | ~new_U3039;
  assign new_U5085 = ~ADDR_REG_5_ | ~new_U4942;
  assign new_U5086 = ~new_R1105_U52 | ~new_U3042;
  assign new_U5087 = ~new_U3040 | ~new_U3440;
  assign new_U5088 = ~new_R1162_U59 | ~new_U3038;
  assign new_U5089 = ~new_U5088 | ~new_U5087 | ~new_U5086;
  assign new_U5090 = ~new_U3044 | ~new_U5089;
  assign new_U5091 = ~new_R1105_U52 | ~new_U3043;
  assign new_U5092 = ~REG3_REG_4_ | ~n1342;
  assign new_U5093 = ~new_U3041 | ~new_U3440;
  assign new_U5094 = ~new_R1162_U59 | ~new_U3039;
  assign new_U5095 = ~ADDR_REG_4_ | ~new_U4942;
  assign new_U5096 = ~new_R1105_U53 | ~new_U3042;
  assign new_U5097 = ~new_U3040 | ~new_U3441;
  assign new_U5098 = ~new_R1162_U60 | ~new_U3038;
  assign new_U5099 = ~new_U5098 | ~new_U5097 | ~new_U5096;
  assign new_U5100 = ~new_U3044 | ~new_U5099;
  assign new_U5101 = ~new_R1105_U53 | ~new_U3043;
  assign new_U5102 = ~REG3_REG_3_ | ~n1342;
  assign new_U5103 = ~new_U3041 | ~new_U3441;
  assign new_U5104 = ~new_R1162_U60 | ~new_U3039;
  assign new_U5105 = ~ADDR_REG_3_ | ~new_U4942;
  assign new_U5106 = ~new_R1105_U54 | ~new_U3042;
  assign new_U5107 = ~new_U3040 | ~new_U3442;
  assign new_U5108 = ~new_R1162_U61 | ~new_U3038;
  assign new_U5109 = ~new_U5108 | ~new_U5107 | ~new_U5106;
  assign new_U5110 = ~new_U3044 | ~new_U5109;
  assign new_U5111 = ~new_R1105_U54 | ~new_U3043;
  assign new_U5112 = ~REG3_REG_2_ | ~n1342;
  assign new_U5113 = ~new_U3041 | ~new_U3442;
  assign new_U5114 = ~new_R1162_U61 | ~new_U3039;
  assign new_U5115 = ~ADDR_REG_2_ | ~new_U4942;
  assign new_U5116 = ~new_R1105_U5 | ~new_U3042;
  assign new_U5117 = ~new_U3040 | ~new_U3443;
  assign new_U5118 = ~new_R1162_U5 | ~new_U3038;
  assign new_U5119 = ~new_U5118 | ~new_U5117 | ~new_U5116;
  assign new_U5120 = ~new_U3044 | ~new_U5119;
  assign new_U5121 = ~new_R1105_U5 | ~new_U3043;
  assign new_U5122 = ~REG3_REG_1_ | ~n1342;
  assign new_U5123 = ~new_U3041 | ~new_U3443;
  assign new_U5124 = ~new_R1162_U5 | ~new_U3039;
  assign new_U5125 = ~ADDR_REG_1_ | ~new_U4942;
  assign new_U5126 = ~new_R1105_U46 | ~new_U3042;
  assign new_U5127 = ~new_U3040 | ~new_U3453;
  assign new_U5128 = ~new_R1162_U53 | ~new_U3038;
  assign new_U5129 = ~new_U5128 | ~new_U5127 | ~new_U5126;
  assign new_U5130 = ~new_U3044 | ~new_U5129;
  assign new_U5131 = ~new_R1105_U46 | ~new_U3043;
  assign new_U5132 = ~REG3_REG_0_ | ~n1342;
  assign new_U5133 = ~new_U3041 | ~new_U3453;
  assign new_U5134 = ~new_R1162_U53 | ~new_U3039;
  assign new_U5135 = ~ADDR_REG_0_ | ~new_U4942;
  assign new_U5136 = ~new_U3903 | ~new_U6257 | ~new_U6256;
  assign new_U5137 = ~new_U3425;
  assign new_U5138 = ~new_U5137 | ~new_U4055;
  assign new_U5139 = ~new_U4006 | ~new_U5138;
  assign new_U5140 = ~new_U4020 | ~new_U3424;
  assign new_U5141 = ~new_U4012 | ~new_U4005;
  assign new_U5142 = ~new_U3902 | ~new_U6253 | ~new_U6252;
  assign new_U5143 = ~new_U4005 | ~new_U3461 | ~new_U3014;
  assign new_U5144 = ~new_U3431 | ~new_U5142;
  assign new_U5145 = ~new_U5144 | ~new_U5143;
  assign new_U5146 = ~new_R395_U6 | ~new_U4041 | ~new_U3023;
  assign new_U5147 = ~new_U5145 | ~STATE_REG;
  assign new_U5148 = ~B_REG | ~new_U5136;
  assign new_U5149 = ~new_U3037 | ~new_U3076;
  assign new_U5150 = ~new_U3035 | ~new_U3070;
  assign new_U5151 = ~new_ADD_95_U65 | ~new_U3427;
  assign new_U5152 = ~new_U5151 | ~new_U5150 | ~new_U5149;
  assign new_U5153 = ~new_U3362 | ~new_U3364 | ~new_U3363;
  assign new_U5154 = ~new_U3419 | ~new_U3366;
  assign new_U5155 = ~new_U5805 | ~new_U5154;
  assign new_U5156 = ~new_U5808 | ~new_U5153;
  assign new_U5157 = ~new_U3906 | ~new_U5155 | ~new_U5156 | ~new_U3369;
  assign new_U5158 = ~new_U5157 | ~new_U3427;
  assign new_U5159 = ~new_U3429;
  assign new_U5160 = ~new_U3496 | ~new_U5744;
  assign new_U5161 = ~new_ADD_95_U65 | ~new_U5743;
  assign new_U5162 = ~new_U4049 | ~new_U5152;
  assign new_U5163 = ~new_R1165_U109 | ~new_U3028;
  assign new_U5164 = ~REG3_REG_15_ | ~n1342;
  assign new_U5165 = ~new_U3037 | ~new_U3055;
  assign new_U5166 = ~new_U3035 | ~new_U3050;
  assign new_U5167 = ~new_ADD_95_U54 | ~new_U3427;
  assign new_U5168 = ~new_U5167 | ~new_U5166 | ~new_U5165;
  assign new_U5169 = ~new_U4021 | ~new_U3427;
  assign new_U5170 = ~new_U5159 | ~new_U5169;
  assign new_U5171 = ~new_U4028 | ~new_U4021;
  assign new_U5172 = ~new_U3418 | ~new_U5171;
  assign new_U5173 = ~new_U3046 | ~new_U4031;
  assign new_U5174 = ~new_U3045 | ~new_ADD_95_U54;
  assign new_U5175 = ~new_U4049 | ~new_U5168;
  assign new_U5176 = ~new_R1165_U15 | ~new_U3028;
  assign new_U5177 = ~REG3_REG_26_ | ~n1342;
  assign new_U5178 = ~new_U3037 | ~new_U3064;
  assign new_U5179 = ~new_U3035 | ~new_U3067;
  assign new_U5180 = ~new_ADD_95_U49 | ~new_U3427;
  assign new_U5181 = ~new_U5180 | ~new_U5179 | ~new_U5178;
  assign new_U5182 = ~new_U3478 | ~new_U5744;
  assign new_U5183 = ~new_ADD_95_U49 | ~new_U5743;
  assign new_U5184 = ~new_U4049 | ~new_U5181;
  assign new_U5185 = ~new_R1165_U94 | ~new_U3028;
  assign new_U5186 = ~REG3_REG_6_ | ~n1342;
  assign new_U5187 = ~new_U3037 | ~new_U3066;
  assign new_U5188 = ~new_U3035 | ~new_U3078;
  assign new_U5189 = ~new_ADD_95_U62 | ~new_U3427;
  assign new_U5190 = ~new_U5189 | ~new_U5188 | ~new_U5187;
  assign new_U5191 = ~new_U3502 | ~new_U5744;
  assign new_U5192 = ~new_ADD_95_U62 | ~new_U5743;
  assign new_U5193 = ~new_U4049 | ~new_U5190;
  assign new_U5194 = ~new_R1165_U107 | ~new_U3028;
  assign new_U5195 = ~REG3_REG_18_ | ~n1342;
  assign new_U5196 = ~new_U3037 | ~new_U3075;
  assign new_U5197 = ~new_U3035 | ~new_U3061;
  assign new_U5198 = ~REG3_REG_2_ | ~new_U3427;
  assign new_U5199 = ~new_U5198 | ~new_U5197 | ~new_U5196;
  assign new_U5200 = ~new_U3470 | ~new_U5744;
  assign new_U5201 = ~REG3_REG_2_ | ~new_U5743;
  assign new_U5202 = ~new_U4049 | ~new_U5199;
  assign new_U5203 = ~new_R1165_U97 | ~new_U3028;
  assign new_U5204 = ~REG3_REG_2_ | ~n1342;
  assign new_U5205 = ~new_U3037 | ~new_U3059;
  assign new_U5206 = ~new_U3035 | ~new_U3069;
  assign new_U5207 = ~new_ADD_95_U69 | ~new_U3427;
  assign new_U5208 = ~new_U5207 | ~new_U5206 | ~new_U5205;
  assign new_U5209 = ~new_U3488 | ~new_U5744;
  assign new_U5210 = ~new_ADD_95_U69 | ~new_U5743;
  assign new_U5211 = ~new_U4049 | ~new_U5208;
  assign new_U5212 = ~new_R1165_U112 | ~new_U3028;
  assign new_U5213 = ~REG3_REG_11_ | ~n1342;
  assign new_U5214 = ~new_U3037 | ~new_U3072;
  assign new_U5215 = ~new_U3035 | ~new_U3063;
  assign new_U5216 = ~new_ADD_95_U58 | ~new_U3427;
  assign new_U5217 = ~new_U5216 | ~new_U5215 | ~new_U5214;
  assign new_U5218 = ~new_U3046 | ~new_U4035;
  assign new_U5219 = ~new_U3045 | ~new_ADD_95_U58;
  assign new_U5220 = ~new_U4049 | ~new_U5217;
  assign new_U5221 = ~new_R1165_U103 | ~new_U3028;
  assign new_U5222 = ~REG3_REG_22_ | ~n1342;
  assign new_U5223 = ~new_U3037 | ~new_U3069;
  assign new_U5224 = ~new_U3035 | ~new_U3076;
  assign new_U5225 = ~new_ADD_95_U67 | ~new_U3427;
  assign new_U5226 = ~new_U5225 | ~new_U5224 | ~new_U5223;
  assign new_U5227 = ~new_U3492 | ~new_U5744;
  assign new_U5228 = ~new_ADD_95_U67 | ~new_U5743;
  assign new_U5229 = ~new_U4049 | ~new_U5226;
  assign new_U5230 = ~new_R1165_U12 | ~new_U3028;
  assign new_U5231 = ~REG3_REG_13_ | ~n1342;
  assign new_U5232 = ~new_U3037 | ~new_U3078;
  assign new_U5233 = ~new_U3035 | ~new_U3072;
  assign new_U5234 = ~new_ADD_95_U60 | ~new_U3427;
  assign new_U5235 = ~new_U5234 | ~new_U5233 | ~new_U5232;
  assign new_U5236 = ~new_U3046 | ~new_U4037;
  assign new_U5237 = ~new_U3045 | ~new_ADD_95_U60;
  assign new_U5238 = ~new_U4049 | ~new_U5235;
  assign new_U5239 = ~new_R1165_U104 | ~new_U3028;
  assign new_U5240 = ~REG3_REG_20_ | ~n1342;
  assign new_U5241 = ~new_U3428 | ~new_U3426;
  assign new_U5242 = ~new_U5241 | ~new_U3427;
  assign new_U5243 = ~new_U4050 | ~new_U5242;
  assign new_U5244 = ~new_U3911 | ~new_U3035;
  assign new_U5245 = ~new_U3464 | ~new_U5744;
  assign new_U5246 = ~REG3_REG_0_ | ~new_U5243;
  assign new_U5247 = ~new_R1165_U91 | ~new_U3028;
  assign new_U5248 = ~REG3_REG_0_ | ~n1342;
  assign new_U5249 = ~new_U3037 | ~new_U3081;
  assign new_U5250 = ~new_U3035 | ~new_U3059;
  assign new_U5251 = ~new_ADD_95_U46 | ~new_U3427;
  assign new_U5252 = ~new_U5251 | ~new_U5250 | ~new_U5249;
  assign new_U5253 = ~new_U3484 | ~new_U5744;
  assign new_U5254 = ~new_ADD_95_U46 | ~new_U5743;
  assign new_U5255 = ~new_U4049 | ~new_U5252;
  assign new_U5256 = ~new_R1165_U92 | ~new_U3028;
  assign new_U5257 = ~REG3_REG_9_ | ~n1342;
  assign new_U5258 = ~new_U3037 | ~new_U3061;
  assign new_U5259 = ~new_U3035 | ~new_U3064;
  assign new_U5260 = ~new_ADD_95_U51 | ~new_U3427;
  assign new_U5261 = ~new_U5260 | ~new_U5259 | ~new_U5258;
  assign new_U5262 = ~new_U3474 | ~new_U5744;
  assign new_U5263 = ~new_ADD_95_U51 | ~new_U5743;
  assign new_U5264 = ~new_U4049 | ~new_U5261;
  assign new_U5265 = ~new_R1165_U96 | ~new_U3028;
  assign new_U5266 = ~REG3_REG_4_ | ~n1342;
  assign new_U5267 = ~new_U3037 | ~new_U3063;
  assign new_U5268 = ~new_U3035 | ~new_U3055;
  assign new_U5269 = ~new_ADD_95_U56 | ~new_U3427;
  assign new_U5270 = ~new_U5269 | ~new_U5268 | ~new_U5267;
  assign new_U5271 = ~new_U3046 | ~new_U4033;
  assign new_U5272 = ~new_U3045 | ~new_ADD_95_U56;
  assign new_U5273 = ~new_U4049 | ~new_U5270;
  assign new_U5274 = ~new_R1165_U101 | ~new_U3028;
  assign new_U5275 = ~REG3_REG_24_ | ~n1342;
  assign new_U5276 = ~new_U3037 | ~new_U3070;
  assign new_U5277 = ~new_U3035 | ~new_U3079;
  assign new_U5278 = ~new_ADD_95_U63 | ~new_U3427;
  assign new_U5279 = ~new_U5278 | ~new_U5277 | ~new_U5276;
  assign new_U5280 = ~new_U3500 | ~new_U5744;
  assign new_U5281 = ~new_ADD_95_U63 | ~new_U5743;
  assign new_U5282 = ~new_U4049 | ~new_U5279;
  assign new_U5283 = ~new_R1165_U13 | ~new_U3028;
  assign new_U5284 = ~REG3_REG_17_ | ~n1342;
  assign new_U5285 = ~new_U3037 | ~new_U3057;
  assign new_U5286 = ~new_U3035 | ~new_U3068;
  assign new_U5287 = ~new_ADD_95_U50 | ~new_U3427;
  assign new_U5288 = ~new_U5287 | ~new_U5286 | ~new_U5285;
  assign new_U5289 = ~new_U3476 | ~new_U5744;
  assign new_U5290 = ~new_ADD_95_U50 | ~new_U5743;
  assign new_U5291 = ~new_U4049 | ~new_U5288;
  assign new_U5292 = ~new_R1165_U95 | ~new_U3028;
  assign new_U5293 = ~REG3_REG_5_ | ~n1342;
  assign new_U5294 = ~new_U3037 | ~new_U3071;
  assign new_U5295 = ~new_U3035 | ~new_U3066;
  assign new_U5296 = ~new_ADD_95_U64 | ~new_U3427;
  assign new_U5297 = ~new_U5296 | ~new_U5295 | ~new_U5294;
  assign new_U5298 = ~new_U3498 | ~new_U5744;
  assign new_U5299 = ~new_ADD_95_U64 | ~new_U5743;
  assign new_U5300 = ~new_U4049 | ~new_U5297;
  assign new_U5301 = ~new_R1165_U108 | ~new_U3028;
  assign new_U5302 = ~REG3_REG_16_ | ~n1342;
  assign new_U5303 = ~new_U3037 | ~new_U3062;
  assign new_U5304 = ~new_U3035 | ~new_U3054;
  assign new_U5305 = ~new_ADD_95_U55 | ~new_U3427;
  assign new_U5306 = ~new_U5305 | ~new_U5304 | ~new_U5303;
  assign new_U5307 = ~new_U3046 | ~new_U4032;
  assign new_U5308 = ~new_U3045 | ~new_ADD_95_U55;
  assign new_U5309 = ~new_U4049 | ~new_U5306;
  assign new_U5310 = ~new_R1165_U100 | ~new_U3028;
  assign new_U5311 = ~REG3_REG_25_ | ~n1342;
  assign new_U5312 = ~new_U3037 | ~new_U3060;
  assign new_U5313 = ~new_U3035 | ~new_U3077;
  assign new_U5314 = ~new_ADD_95_U68 | ~new_U3427;
  assign new_U5315 = ~new_U5314 | ~new_U5313 | ~new_U5312;
  assign new_U5316 = ~new_U3490 | ~new_U5744;
  assign new_U5317 = ~new_ADD_95_U68 | ~new_U5743;
  assign new_U5318 = ~new_U4049 | ~new_U5315;
  assign new_U5319 = ~new_R1165_U111 | ~new_U3028;
  assign new_U5320 = ~REG3_REG_12_ | ~n1342;
  assign new_U5321 = ~new_U3037 | ~new_U3073;
  assign new_U5322 = ~new_U3035 | ~new_U3058;
  assign new_U5323 = ~new_ADD_95_U59 | ~new_U3427;
  assign new_U5324 = ~new_U5323 | ~new_U5322 | ~new_U5321;
  assign new_U5325 = ~new_U3046 | ~new_U4036;
  assign new_U5326 = ~new_U3045 | ~new_ADD_95_U59;
  assign new_U5327 = ~new_U4049 | ~new_U5324;
  assign new_U5328 = ~new_R1165_U14 | ~new_U3028;
  assign new_U5329 = ~REG3_REG_21_ | ~n1342;
  assign new_U5330 = ~new_U3037 | ~new_U3074;
  assign new_U5331 = ~new_U3035 | ~new_U3065;
  assign new_U5332 = ~REG3_REG_1_ | ~new_U3427;
  assign new_U5333 = ~new_U5332 | ~new_U5331 | ~new_U5330;
  assign new_U5334 = ~new_U3468 | ~new_U5744;
  assign new_U5335 = ~REG3_REG_1_ | ~new_U5743;
  assign new_U5336 = ~new_U4049 | ~new_U5333;
  assign new_U5337 = ~new_R1165_U105 | ~new_U3028;
  assign new_U5338 = ~REG3_REG_1_ | ~n1342;
  assign new_U5339 = ~new_U3037 | ~new_U3067;
  assign new_U5340 = ~new_U3035 | ~new_U3080;
  assign new_U5341 = ~new_ADD_95_U47 | ~new_U3427;
  assign new_U5342 = ~new_U5341 | ~new_U5340 | ~new_U5339;
  assign new_U5343 = ~new_U3482 | ~new_U5744;
  assign new_U5344 = ~new_ADD_95_U47 | ~new_U5743;
  assign new_U5345 = ~new_U4049 | ~new_U5342;
  assign new_U5346 = ~new_R1165_U93 | ~new_U3028;
  assign new_U5347 = ~REG3_REG_8_ | ~n1342;
  assign new_U5348 = ~new_U3037 | ~new_U3050;
  assign new_U5349 = ~new_U3035 | ~new_U3052;
  assign new_U5350 = ~new_ADD_95_U52 | ~new_U3427;
  assign new_U5351 = ~new_U5350 | ~new_U5349 | ~new_U5348;
  assign new_U5352 = ~new_U3046 | ~new_U4029;
  assign new_U5353 = ~new_U3045 | ~new_ADD_95_U52;
  assign new_U5354 = ~new_U4049 | ~new_U5351;
  assign new_U5355 = ~new_R1165_U98 | ~new_U3028;
  assign new_U5356 = ~REG3_REG_28_ | ~n1342;
  assign new_U5357 = ~new_U3037 | ~new_U3079;
  assign new_U5358 = ~new_U3035 | ~new_U3073;
  assign new_U5359 = ~new_ADD_95_U61 | ~new_U3427;
  assign new_U5360 = ~new_U5359 | ~new_U5358 | ~new_U5357;
  assign new_U5361 = ~new_U3504 | ~new_U5744;
  assign new_U5362 = ~new_ADD_95_U61 | ~new_U5743;
  assign new_U5363 = ~new_U4049 | ~new_U5360;
  assign new_U5364 = ~new_R1165_U106 | ~new_U3028;
  assign new_U5365 = ~REG3_REG_19_ | ~n1342;
  assign new_U5366 = ~new_U3037 | ~new_U3065;
  assign new_U5367 = ~new_U3035 | ~new_U3057;
  assign new_U5368 = ~new_ADD_95_U4 | ~new_U3427;
  assign new_U5369 = ~new_U5368 | ~new_U5367 | ~new_U5366;
  assign new_U5370 = ~new_U3472 | ~new_U5744;
  assign new_U5371 = ~new_ADD_95_U4 | ~new_U5743;
  assign new_U5372 = ~new_U4049 | ~new_U5369;
  assign new_U5373 = ~new_R1165_U16 | ~new_U3028;
  assign new_U5374 = ~REG3_REG_3_ | ~n1342;
  assign new_U5375 = ~new_U3037 | ~new_U3080;
  assign new_U5376 = ~new_U3035 | ~new_U3060;
  assign new_U5377 = ~new_ADD_95_U70 | ~new_U3427;
  assign new_U5378 = ~new_U5377 | ~new_U5376 | ~new_U5375;
  assign new_U5379 = ~new_U3486 | ~new_U5744;
  assign new_U5380 = ~new_ADD_95_U70 | ~new_U5743;
  assign new_U5381 = ~new_U4049 | ~new_U5378;
  assign new_U5382 = ~new_R1165_U113 | ~new_U3028;
  assign new_U5383 = ~REG3_REG_10_ | ~n1342;
  assign new_U5384 = ~new_U3037 | ~new_U3058;
  assign new_U5385 = ~new_U3035 | ~new_U3062;
  assign new_U5386 = ~new_ADD_95_U57 | ~new_U3427;
  assign new_U5387 = ~new_U5386 | ~new_U5385 | ~new_U5384;
  assign new_U5388 = ~new_U3046 | ~new_U4034;
  assign new_U5389 = ~new_U3045 | ~new_ADD_95_U57;
  assign new_U5390 = ~new_U4049 | ~new_U5387;
  assign new_U5391 = ~new_R1165_U102 | ~new_U3028;
  assign new_U5392 = ~REG3_REG_23_ | ~n1342;
  assign new_U5393 = ~new_U3037 | ~new_U3077;
  assign new_U5394 = ~new_U3035 | ~new_U3071;
  assign new_U5395 = ~new_ADD_95_U66 | ~new_U3427;
  assign new_U5396 = ~new_U5395 | ~new_U5394 | ~new_U5393;
  assign new_U5397 = ~new_U3494 | ~new_U5744;
  assign new_U5398 = ~new_ADD_95_U66 | ~new_U5743;
  assign new_U5399 = ~new_U4049 | ~new_U5396;
  assign new_U5400 = ~new_R1165_U110 | ~new_U3028;
  assign new_U5401 = ~REG3_REG_14_ | ~n1342;
  assign new_U5402 = ~new_U3037 | ~new_U3054;
  assign new_U5403 = ~new_U3035 | ~new_U3051;
  assign new_U5404 = ~new_ADD_95_U53 | ~new_U3427;
  assign new_U5405 = ~new_U5404 | ~new_U5403 | ~new_U5402;
  assign new_U5406 = ~new_U3046 | ~new_U4030;
  assign new_U5407 = ~new_U3045 | ~new_ADD_95_U53;
  assign new_U5408 = ~new_U4049 | ~new_U5405;
  assign new_U5409 = ~new_R1165_U99 | ~new_U3028;
  assign new_U5410 = ~REG3_REG_27_ | ~n1342;
  assign new_U5411 = ~new_U3037 | ~new_U3068;
  assign new_U5412 = ~new_U3035 | ~new_U3081;
  assign new_U5413 = ~new_ADD_95_U48 | ~new_U3427;
  assign new_U5414 = ~new_U5413 | ~new_U5412 | ~new_U5411;
  assign new_U5415 = ~new_U3480 | ~new_U5744;
  assign new_U5416 = ~new_ADD_95_U48 | ~new_U5743;
  assign new_U5417 = ~new_U4049 | ~new_U5414;
  assign new_U5418 = ~new_R1165_U17 | ~new_U3028;
  assign new_U5419 = ~REG3_REG_7_ | ~n1342;
  assign new_U5420 = ~new_U3455 | ~new_U3376;
  assign new_U5421 = ~new_U3454 | ~new_U5420;
  assign new_U5422 = ~new_R1165_U91 | ~new_U5802 | ~new_U3454;
  assign new_U5423 = ~new_U3014 | ~new_U3484;
  assign new_U5424 = ~new_U3582 | ~new_U3460;
  assign new_U5425 = ~new_U5805 | ~new_U3080;
  assign new_U5426 = ~new_U3014 | ~new_U3482;
  assign new_U5427 = ~new_U3583 | ~new_U3460;
  assign new_U5428 = ~new_U5805 | ~new_U3081;
  assign new_U5429 = ~new_U3014 | ~new_U3480;
  assign new_U5430 = ~new_U3584 | ~new_U3460;
  assign new_U5431 = ~new_U5805 | ~new_U3067;
  assign new_U5432 = ~new_U3014 | ~new_U3478;
  assign new_U5433 = ~new_U3585 | ~new_U3460;
  assign new_U5434 = ~new_U5805 | ~new_U3068;
  assign new_U5435 = ~new_U3014 | ~new_U3476;
  assign new_U5436 = ~new_U3586 | ~new_U3460;
  assign new_U5437 = ~new_U5805 | ~new_U3064;
  assign new_U5438 = ~new_U3014 | ~new_U3474;
  assign new_U5439 = ~new_U3587 | ~new_U3460;
  assign new_U5440 = ~new_U5805 | ~new_U3057;
  assign new_U5441 = ~new_U3588 | ~new_U3460;
  assign new_U5442 = ~new_U3014 | ~new_U4038;
  assign new_U5443 = ~new_U5805 | ~new_U3053;
  assign new_U5444 = ~new_U3589 | ~new_U3460;
  assign new_U5445 = ~new_U3014 | ~new_U4039;
  assign new_U5446 = ~new_U5805 | ~new_U3056;
  assign new_U5447 = ~new_U3014 | ~new_U3472;
  assign new_U5448 = ~new_U3590 | ~new_U3460;
  assign new_U5449 = ~new_U5805 | ~new_U3061;
  assign new_U5450 = ~new_U3591 | ~new_U3460;
  assign new_U5451 = ~new_U3014 | ~new_U4040;
  assign new_U5452 = ~new_U5805 | ~new_U3052;
  assign new_U5453 = ~new_U3592 | ~new_U3460;
  assign new_U5454 = ~new_U3014 | ~new_U4029;
  assign new_U5455 = ~new_U5805 | ~new_U3051;
  assign new_U5456 = ~new_U3593 | ~new_U3460;
  assign new_U5457 = ~new_U3014 | ~new_U4030;
  assign new_U5458 = ~new_U5805 | ~new_U3050;
  assign new_U5459 = ~new_U3594 | ~new_U3460;
  assign new_U5460 = ~new_U3014 | ~new_U4031;
  assign new_U5461 = ~new_U5805 | ~new_U3054;
  assign new_U5462 = ~new_U3595 | ~new_U3460;
  assign new_U5463 = ~new_U3014 | ~new_U4032;
  assign new_U5464 = ~new_U5805 | ~new_U3055;
  assign new_U5465 = ~new_U3596 | ~new_U3460;
  assign new_U5466 = ~new_U3014 | ~new_U4033;
  assign new_U5467 = ~new_U5805 | ~new_U3062;
  assign new_U5468 = ~new_U3597 | ~new_U3460;
  assign new_U5469 = ~new_U3014 | ~new_U4034;
  assign new_U5470 = ~new_U5805 | ~new_U3063;
  assign new_U5471 = ~new_U3598 | ~new_U3460;
  assign new_U5472 = ~new_U3014 | ~new_U4035;
  assign new_U5473 = ~new_U5805 | ~new_U3058;
  assign new_U5474 = ~new_U3599 | ~new_U3460;
  assign new_U5475 = ~new_U3014 | ~new_U4036;
  assign new_U5476 = ~new_U5805 | ~new_U3072;
  assign new_U5477 = ~new_U3600 | ~new_U3460;
  assign new_U5478 = ~new_U3014 | ~new_U4037;
  assign new_U5479 = ~new_U5805 | ~new_U3073;
  assign new_U5480 = ~new_U3014 | ~new_U3470;
  assign new_U5481 = ~new_U3601 | ~new_U3460;
  assign new_U5482 = ~new_U5805 | ~new_U3065;
  assign new_U5483 = ~new_U3014 | ~new_U3504;
  assign new_U5484 = ~new_U3602 | ~new_U3460;
  assign new_U5485 = ~new_U5805 | ~new_U3078;
  assign new_U5486 = ~new_U3014 | ~new_U3502;
  assign new_U5487 = ~new_U3603 | ~new_U3460;
  assign new_U5488 = ~new_U5805 | ~new_U3079;
  assign new_U5489 = ~new_U3014 | ~new_U3500;
  assign new_U5490 = ~new_U3604 | ~new_U3460;
  assign new_U5491 = ~new_U5805 | ~new_U3066;
  assign new_U5492 = ~new_U3014 | ~new_U3498;
  assign new_U5493 = ~new_U3605 | ~new_U3460;
  assign new_U5494 = ~new_U5805 | ~new_U3070;
  assign new_U5495 = ~new_U3014 | ~new_U3496;
  assign new_U5496 = ~new_U3606 | ~new_U3460;
  assign new_U5497 = ~new_U5805 | ~new_U3071;
  assign new_U5498 = ~new_U3014 | ~new_U3494;
  assign new_U5499 = ~new_U3607 | ~new_U3460;
  assign new_U5500 = ~new_U5805 | ~new_U3076;
  assign new_U5501 = ~new_U3014 | ~new_U3492;
  assign new_U5502 = ~new_U3608 | ~new_U3460;
  assign new_U5503 = ~new_U5805 | ~new_U3077;
  assign new_U5504 = ~new_U3014 | ~new_U3490;
  assign new_U5505 = ~new_U3609 | ~new_U3460;
  assign new_U5506 = ~new_U5805 | ~new_U3069;
  assign new_U5507 = ~new_U3014 | ~new_U3488;
  assign new_U5508 = ~new_U3610 | ~new_U3460;
  assign new_U5509 = ~new_U5805 | ~new_U3060;
  assign new_U5510 = ~new_U3014 | ~new_U3486;
  assign new_U5511 = ~new_U3611 | ~new_U3460;
  assign new_U5512 = ~new_U5805 | ~new_U3059;
  assign new_U5513 = ~new_U3014 | ~new_U3468;
  assign new_U5514 = ~new_U3612 | ~new_U3460;
  assign new_U5515 = ~new_U5805 | ~new_U3075;
  assign new_U5516 = ~new_U3014 | ~new_U3464;
  assign new_U5517 = ~new_U3613 | ~new_U3460;
  assign new_U5518 = ~new_U5805 | ~new_U3074;
  assign new_U5519 = ~new_U3484 | ~new_U3361;
  assign new_U5520 = ~new_U3014 | ~new_U3080;
  assign new_U5521 = ~new_U5748 | ~new_U3081;
  assign new_U5522 = ~new_U3482 | ~new_U3361;
  assign new_U5523 = ~new_U3014 | ~new_U3081;
  assign new_U5524 = ~new_U5748 | ~new_U3067;
  assign new_U5525 = ~new_U3480 | ~new_U3361;
  assign new_U5526 = ~new_U3014 | ~new_U3067;
  assign new_U5527 = ~new_U5748 | ~new_U3068;
  assign new_U5528 = ~new_U3478 | ~new_U3361;
  assign new_U5529 = ~new_U3014 | ~new_U3068;
  assign new_U5530 = ~new_U5748 | ~new_U3064;
  assign new_U5531 = ~new_U3476 | ~new_U3361;
  assign new_U5532 = ~new_U3014 | ~new_U3064;
  assign new_U5533 = ~new_U5748 | ~new_U3057;
  assign new_U5534 = ~new_U3474 | ~new_U3361;
  assign new_U5535 = ~new_U3014 | ~new_U3057;
  assign new_U5536 = ~new_U5748 | ~new_U3061;
  assign new_U5537 = ~new_U4038 | ~new_U3361;
  assign new_U5538 = ~new_U3014 | ~new_U3053;
  assign new_U5539 = ~new_U4039 | ~new_U3361;
  assign new_U5540 = ~new_U3014 | ~new_U3056;
  assign new_U5541 = ~new_U3472 | ~new_U3361;
  assign new_U5542 = ~new_U3014 | ~new_U3061;
  assign new_U5543 = ~new_U5748 | ~new_U3065;
  assign new_U5544 = ~new_U4040 | ~new_U3361;
  assign new_U5545 = ~new_U3014 | ~new_U3052;
  assign new_U5546 = ~new_U5748 | ~new_U3051;
  assign new_U5547 = ~new_U4029 | ~new_U3361;
  assign new_U5548 = ~new_U3014 | ~new_U3051;
  assign new_U5549 = ~new_U5748 | ~new_U3050;
  assign new_U5550 = ~new_U4030 | ~new_U3361;
  assign new_U5551 = ~new_U3014 | ~new_U3050;
  assign new_U5552 = ~new_U5748 | ~new_U3054;
  assign new_U5553 = ~new_U4031 | ~new_U3361;
  assign new_U5554 = ~new_U3014 | ~new_U3054;
  assign new_U5555 = ~new_U5748 | ~new_U3055;
  assign new_U5556 = ~new_U4032 | ~new_U3361;
  assign new_U5557 = ~new_U3014 | ~new_U3055;
  assign new_U5558 = ~new_U5748 | ~new_U3062;
  assign new_U5559 = ~new_U4033 | ~new_U3361;
  assign new_U5560 = ~new_U3014 | ~new_U3062;
  assign new_U5561 = ~new_U5748 | ~new_U3063;
  assign new_U5562 = ~new_U4034 | ~new_U3361;
  assign new_U5563 = ~new_U3014 | ~new_U3063;
  assign new_U5564 = ~new_U5748 | ~new_U3058;
  assign new_U5565 = ~new_U4035 | ~new_U3361;
  assign new_U5566 = ~new_U3014 | ~new_U3058;
  assign new_U5567 = ~new_U5748 | ~new_U3072;
  assign new_U5568 = ~new_U4036 | ~new_U3361;
  assign new_U5569 = ~new_U3014 | ~new_U3072;
  assign new_U5570 = ~new_U5748 | ~new_U3073;
  assign new_U5571 = ~new_U4037 | ~new_U3361;
  assign new_U5572 = ~new_U3014 | ~new_U3073;
  assign new_U5573 = ~new_U5748 | ~new_U3078;
  assign new_U5574 = ~new_U3470 | ~new_U3361;
  assign new_U5575 = ~new_U3014 | ~new_U3065;
  assign new_U5576 = ~new_U5748 | ~new_U3075;
  assign new_U5577 = ~new_U3504 | ~new_U3361;
  assign new_U5578 = ~new_U3014 | ~new_U3078;
  assign new_U5579 = ~new_U5748 | ~new_U3079;
  assign new_U5580 = ~new_U3502 | ~new_U3361;
  assign new_U5581 = ~new_U3014 | ~new_U3079;
  assign new_U5582 = ~new_U5748 | ~new_U3066;
  assign new_U5583 = ~new_U3500 | ~new_U3361;
  assign new_U5584 = ~new_U3014 | ~new_U3066;
  assign new_U5585 = ~new_U5748 | ~new_U3070;
  assign new_U5586 = ~new_U3498 | ~new_U3361;
  assign new_U5587 = ~new_U3014 | ~new_U3070;
  assign new_U5588 = ~new_U5748 | ~new_U3071;
  assign new_U5589 = ~new_U3496 | ~new_U3361;
  assign new_U5590 = ~new_U3014 | ~new_U3071;
  assign new_U5591 = ~new_U5748 | ~new_U3076;
  assign new_U5592 = ~new_U3494 | ~new_U3361;
  assign new_U5593 = ~new_U3014 | ~new_U3076;
  assign new_U5594 = ~new_U5748 | ~new_U3077;
  assign new_U5595 = ~new_U3492 | ~new_U3361;
  assign new_U5596 = ~new_U3014 | ~new_U3077;
  assign new_U5597 = ~new_U5748 | ~new_U3069;
  assign new_U5598 = ~new_U3490 | ~new_U3361;
  assign new_U5599 = ~new_U3014 | ~new_U3069;
  assign new_U5600 = ~new_U5748 | ~new_U3060;
  assign new_U5601 = ~new_U3488 | ~new_U3361;
  assign new_U5602 = ~new_U3014 | ~new_U3060;
  assign new_U5603 = ~new_U5748 | ~new_U3059;
  assign new_U5604 = ~new_U3486 | ~new_U3361;
  assign new_U5605 = ~new_U3014 | ~new_U3059;
  assign new_U5606 = ~new_U5748 | ~new_U3080;
  assign new_U5607 = ~new_U3468 | ~new_U3361;
  assign new_U5608 = ~new_U3014 | ~new_U3075;
  assign new_U5609 = ~new_U5748 | ~new_U3074;
  assign new_U5610 = ~new_U3464 | ~new_U3361;
  assign new_U5611 = ~new_U3014 | ~new_U3074;
  assign new_U5612 = ~new_U3963 | ~new_U4026;
  assign new_U5613 = ~new_U3370 | ~new_U3419;
  assign new_U5614 = ~new_U3367 | ~new_U3366 | ~new_U3374 | ~new_U3368;
  assign new_U5615 = ~new_U5614 | ~new_U3355;
  assign new_U5616 = ~new_U4057 | ~new_U3355;
  assign new_U5617 = ~new_U5616 | ~new_U5615;
  assign new_U5618 = ~new_U3964 | ~new_U5615;
  assign new_U5619 = ~new_U3484 | ~new_U5618;
  assign new_U5620 = ~new_U3022 | ~new_U3080;
  assign new_U5621 = ~new_U3482 | ~new_U5618;
  assign new_U5622 = ~new_U3022 | ~new_U3081;
  assign new_U5623 = ~new_U3480 | ~new_U5618;
  assign new_U5624 = ~new_U3022 | ~new_U3067;
  assign new_U5625 = ~new_U3478 | ~new_U5618;
  assign new_U5626 = ~new_U3022 | ~new_U3068;
  assign new_U5627 = ~new_U3476 | ~new_U5618;
  assign new_U5628 = ~new_U3022 | ~new_U3064;
  assign new_U5629 = ~new_U3474 | ~new_U5618;
  assign new_U5630 = ~new_U3022 | ~new_U3057;
  assign new_U5631 = ~new_U3472 | ~new_U5618;
  assign new_U5632 = ~new_U3022 | ~new_U3061;
  assign new_U5633 = ~new_U4029 | ~new_U5618;
  assign new_U5634 = ~new_U3022 | ~new_U3051;
  assign new_U5635 = ~new_U4030 | ~new_U5618;
  assign new_U5636 = ~new_U3022 | ~new_U3050;
  assign new_U5637 = ~new_U4031 | ~new_U5618;
  assign new_U5638 = ~new_U3022 | ~new_U3054;
  assign new_U5639 = ~new_U4032 | ~new_U5618;
  assign new_U5640 = ~new_U3022 | ~new_U3055;
  assign new_U5641 = ~new_U4033 | ~new_U5618;
  assign new_U5642 = ~new_U3022 | ~new_U3062;
  assign new_U5643 = ~new_U4034 | ~new_U5618;
  assign new_U5644 = ~new_U3022 | ~new_U3063;
  assign new_U5645 = ~new_U4035 | ~new_U5618;
  assign new_U5646 = ~new_U3022 | ~new_U3058;
  assign new_U5647 = ~new_U4036 | ~new_U5618;
  assign new_U5648 = ~new_U3022 | ~new_U3072;
  assign new_U5649 = ~new_U4037 | ~new_U5618;
  assign new_U5650 = ~new_U3022 | ~new_U3073;
  assign new_U5651 = ~new_U3470 | ~new_U5618;
  assign new_U5652 = ~new_U3022 | ~new_U3065;
  assign new_U5653 = ~new_U3504 | ~new_U5618;
  assign new_U5654 = ~new_U3022 | ~new_U3078;
  assign new_U5655 = ~new_U3502 | ~new_U5618;
  assign new_U5656 = ~new_U3022 | ~new_U3079;
  assign new_U5657 = ~new_U3500 | ~new_U5618;
  assign new_U5658 = ~new_U3022 | ~new_U3066;
  assign new_U5659 = ~new_U3498 | ~new_U5618;
  assign new_U5660 = ~new_U3022 | ~new_U3070;
  assign new_U5661 = ~new_U3496 | ~new_U5618;
  assign new_U5662 = ~new_U3022 | ~new_U3071;
  assign new_U5663 = ~new_U3494 | ~new_U5618;
  assign new_U5664 = ~new_U3022 | ~new_U3076;
  assign new_U5665 = ~new_U3492 | ~new_U5618;
  assign new_U5666 = ~new_U3022 | ~new_U3077;
  assign new_U5667 = ~new_U3490 | ~new_U5618;
  assign new_U5668 = ~new_U3022 | ~new_U3069;
  assign new_U5669 = ~new_U3488 | ~new_U5618;
  assign new_U5670 = ~new_U3022 | ~new_U3060;
  assign new_U5671 = ~new_U3486 | ~new_U5618;
  assign new_U5672 = ~new_U3022 | ~new_U3059;
  assign new_U5673 = ~new_U3468 | ~new_U5618;
  assign new_U5674 = ~new_U3022 | ~new_U3075;
  assign new_U5675 = ~new_U3464 | ~new_U5618;
  assign new_U5676 = ~new_U3022 | ~new_U3074;
  assign new_U5677 = ~REG1_REG_0_ | ~new_U4059;
  assign new_U5678 = ~new_U3022 | ~new_U3484;
  assign new_U5679 = ~new_U5617 | ~new_U3080;
  assign new_U5680 = ~new_U3022 | ~new_U3482;
  assign new_U5681 = ~new_U5617 | ~new_U3081;
  assign new_U5682 = ~new_U3022 | ~new_U3480;
  assign new_U5683 = ~new_U5617 | ~new_U3067;
  assign new_U5684 = ~new_U3022 | ~new_U3478;
  assign new_U5685 = ~new_U5617 | ~new_U3068;
  assign new_U5686 = ~new_U3022 | ~new_U3476;
  assign new_U5687 = ~new_U5617 | ~new_U3064;
  assign new_U5688 = ~new_U3022 | ~new_U3474;
  assign new_U5689 = ~new_U5617 | ~new_U3057;
  assign new_U5690 = ~new_U3022 | ~new_U3472;
  assign new_U5691 = ~new_U5617 | ~new_U3061;
  assign new_U5692 = ~new_U3022 | ~new_U4029;
  assign new_U5693 = ~new_U5617 | ~new_U3051;
  assign new_U5694 = ~new_U3022 | ~new_U4030;
  assign new_U5695 = ~new_U5617 | ~new_U3050;
  assign new_U5696 = ~new_U3022 | ~new_U4031;
  assign new_U5697 = ~new_U5617 | ~new_U3054;
  assign new_U5698 = ~new_U3022 | ~new_U4032;
  assign new_U5699 = ~new_U5617 | ~new_U3055;
  assign new_U5700 = ~new_U3022 | ~new_U4033;
  assign new_U5701 = ~new_U5617 | ~new_U3062;
  assign new_U5702 = ~new_U3022 | ~new_U4034;
  assign new_U5703 = ~new_U5617 | ~new_U3063;
  assign new_U5704 = ~new_U3022 | ~new_U4035;
  assign new_U5705 = ~new_U5617 | ~new_U3058;
  assign new_U5706 = ~new_U3022 | ~new_U4036;
  assign new_U5707 = ~new_U5617 | ~new_U3072;
  assign new_U5708 = ~new_U3022 | ~new_U4037;
  assign new_U5709 = ~new_U5617 | ~new_U3073;
  assign new_U5710 = ~new_U3022 | ~new_U3470;
  assign new_U5711 = ~new_U5617 | ~new_U3065;
  assign new_U5712 = ~new_U3022 | ~new_U3504;
  assign new_U5713 = ~new_U5617 | ~new_U3078;
  assign new_U5714 = ~new_U3022 | ~new_U3502;
  assign new_U5715 = ~new_U5617 | ~new_U3079;
  assign new_U5716 = ~new_U3022 | ~new_U3500;
  assign new_U5717 = ~new_U5617 | ~new_U3066;
  assign new_U5718 = ~new_U3022 | ~new_U3498;
  assign new_U5719 = ~new_U5617 | ~new_U3070;
  assign new_U5720 = ~new_U3022 | ~new_U3496;
  assign new_U5721 = ~new_U5617 | ~new_U3071;
  assign new_U5722 = ~new_U3022 | ~new_U3494;
  assign new_U5723 = ~new_U5617 | ~new_U3076;
  assign new_U5724 = ~new_U3022 | ~new_U3492;
  assign new_U5725 = ~new_U5617 | ~new_U3077;
  assign new_U5726 = ~new_U3022 | ~new_U3490;
  assign new_U5727 = ~new_U5617 | ~new_U3069;
  assign new_U5728 = ~new_U3022 | ~new_U3488;
  assign new_U5729 = ~new_U5617 | ~new_U3060;
  assign new_U5730 = ~new_U3022 | ~new_U3486;
  assign new_U5731 = ~new_U5617 | ~new_U3059;
  assign new_U5732 = ~new_U3022 | ~new_U3468;
  assign new_U5733 = ~new_U5617 | ~new_U3075;
  assign new_U5734 = ~new_U3022 | ~new_U3464;
  assign new_U5735 = ~new_U5617 | ~new_U3074;
  assign new_U5736 = ~new_U4059 | ~new_U3453;
  assign new_U5737 = ~new_R1207_U28 | ~new_U4013;
  assign new_U5738 = ~new_R1192_U28 | ~new_U4014;
  assign new_U5739 = ~new_R1150_U27 | ~new_U4016;
  assign new_U5740 = ~new_R1117_U26 | ~new_U4018;
  assign new_U5741 = ~new_U4052 | ~new_U3427;
  assign new_U5742 = ~new_U4028 | ~new_U4052;
  assign new_U5743 = ~new_U5741 | ~new_U4050;
  assign new_U5744 = ~new_U5742 | ~new_U4051;
  assign new_U5745 = ~new_U5754 | ~new_U5751;
  assign new_U5746 = ~IR_REG_23_ | ~new_U3967;
  assign new_U5747 = ~IR_REG_31_ | ~new_SUB_84_U81;
  assign new_U5748 = ~new_U3431;
  assign new_U5749 = ~IR_REG_24_ | ~new_U3967;
  assign new_U5750 = ~IR_REG_31_ | ~new_SUB_84_U78;
  assign new_U5751 = ~new_U3434;
  assign new_U5752 = ~IR_REG_26_ | ~new_U3967;
  assign new_U5753 = ~IR_REG_31_ | ~new_SUB_84_U17;
  assign new_U5754 = ~new_U3432;
  assign new_U5755 = ~IR_REG_25_ | ~new_U3967;
  assign new_U5756 = ~IR_REG_31_ | ~new_SUB_84_U16;
  assign new_U5757 = ~new_U3433;
  assign new_U5758 = ~IR_REG_9_ | ~new_U3967;
  assign new_U5759 = ~IR_REG_31_ | ~new_SUB_84_U25;
  assign new_U5760 = ~IR_REG_8_ | ~new_U3967;
  assign new_U5761 = ~IR_REG_31_ | ~new_SUB_84_U68;
  assign new_U5762 = ~IR_REG_7_ | ~new_U3967;
  assign new_U5763 = ~IR_REG_31_ | ~new_SUB_84_U24;
  assign new_U5764 = ~IR_REG_6_ | ~new_U3967;
  assign new_U5765 = ~IR_REG_31_ | ~new_SUB_84_U23;
  assign new_U5766 = ~IR_REG_5_ | ~new_U3967;
  assign new_U5767 = ~IR_REG_31_ | ~new_SUB_84_U22;
  assign new_U5768 = ~IR_REG_4_ | ~new_U3967;
  assign new_U5769 = ~IR_REG_31_ | ~new_SUB_84_U70;
  assign new_U5770 = ~IR_REG_3_ | ~new_U3967;
  assign new_U5771 = ~IR_REG_31_ | ~new_SUB_84_U21;
  assign new_U5772 = ~IR_REG_2_ | ~new_U3967;
  assign new_U5773 = ~IR_REG_31_ | ~new_SUB_84_U20;
  assign new_U5774 = ~IR_REG_1_ | ~new_U3967;
  assign new_U5775 = ~IR_REG_31_ | ~new_SUB_84_U48;
  assign new_U5776 = ~IR_REG_18_ | ~new_U3967;
  assign new_U5777 = ~IR_REG_31_ | ~new_SUB_84_U12;
  assign new_U5778 = ~IR_REG_17_ | ~new_U3967;
  assign new_U5779 = ~IR_REG_31_ | ~new_SUB_84_U11;
  assign new_U5780 = ~IR_REG_16_ | ~new_U3967;
  assign new_U5781 = ~IR_REG_31_ | ~new_SUB_84_U87;
  assign new_U5782 = ~IR_REG_15_ | ~new_U3967;
  assign new_U5783 = ~IR_REG_31_ | ~new_SUB_84_U10;
  assign new_U5784 = ~IR_REG_14_ | ~new_U3967;
  assign new_U5785 = ~IR_REG_31_ | ~new_SUB_84_U9;
  assign new_U5786 = ~IR_REG_13_ | ~new_U3967;
  assign new_U5787 = ~IR_REG_31_ | ~new_SUB_84_U8;
  assign new_U5788 = ~IR_REG_12_ | ~new_U3967;
  assign new_U5789 = ~IR_REG_31_ | ~new_SUB_84_U89;
  assign new_U5790 = ~IR_REG_11_ | ~new_U3967;
  assign new_U5791 = ~IR_REG_31_ | ~new_SUB_84_U7;
  assign new_U5792 = ~IR_REG_10_ | ~new_U3967;
  assign new_U5793 = ~IR_REG_31_ | ~new_SUB_84_U6;
  assign new_U5794 = ~IR_REG_0_ | ~new_U3967;
  assign new_U5795 = ~IR_REG_31_ | ~IR_REG_0_;
  assign new_U5796 = ~new_U3453;
  assign new_U5797 = ~IR_REG_28_ | ~new_U3967;
  assign new_U5798 = ~IR_REG_31_ | ~new_SUB_84_U18;
  assign new_U5799 = ~new_U3454;
  assign new_U5800 = ~IR_REG_27_ | ~new_U3967;
  assign new_U5801 = ~IR_REG_31_ | ~new_SUB_84_U76;
  assign new_U5802 = ~new_U3455;
  assign new_U5803 = ~IR_REG_22_ | ~new_U3967;
  assign new_U5804 = ~IR_REG_31_ | ~new_SUB_84_U15;
  assign new_U5805 = ~new_U3456;
  assign new_U5806 = ~IR_REG_21_ | ~new_U3967;
  assign new_U5807 = ~IR_REG_31_ | ~new_SUB_84_U14;
  assign new_U5808 = ~new_U3457;
  assign new_U5809 = ~new_U3434 | ~new_U3359;
  assign new_U5810 = ~B_REG | ~new_U4058 | ~new_U5751;
  assign new_U5811 = ~D_REG_0_ | ~new_U3968;
  assign new_U5812 = ~new_U4047 | ~new_U4162;
  assign new_U5813 = ~D_REG_1_ | ~new_U3968;
  assign new_U5814 = ~new_U4047 | ~new_U4163;
  assign new_U5815 = ~IR_REG_19_ | ~new_U3967;
  assign new_U5816 = ~IR_REG_31_ | ~new_SUB_84_U13;
  assign new_U5817 = ~new_U3461;
  assign new_U5818 = ~IR_REG_20_ | ~new_U3967;
  assign new_U5819 = ~IR_REG_31_ | ~new_SUB_84_U83;
  assign new_U5820 = ~new_U3460;
  assign new_U5821 = ~IR_REG_30_ | ~new_U3967;
  assign new_U5822 = ~IR_REG_31_ | ~new_SUB_84_U73;
  assign new_U5823 = ~new_U3462;
  assign new_U5824 = ~IR_REG_29_ | ~new_U3967;
  assign new_U5825 = ~IR_REG_31_ | ~new_SUB_84_U19;
  assign new_U5826 = ~new_U3463;
  assign new_U5827 = ~DATAI_0_ | ~new_U3969;
  assign new_U5828 = ~new_U4027 | ~new_U3453;
  assign new_U5829 = ~new_U3464;
  assign new_U5830 = ~new_U3456 | ~new_U5808;
  assign new_U5831 = ~new_U3457 | ~new_U5805;
  assign new_U5832 = ~D_REG_1_ | ~new_U4161;
  assign new_U5833 = ~new_U4163 | ~new_U3360;
  assign new_U5834 = ~new_U3466;
  assign new_U5835 = ~new_U5745 | ~new_U3360;
  assign new_U5836 = ~D_REG_0_ | ~new_U4161;
  assign new_U5837 = ~new_U3465;
  assign new_U5838 = ~REG0_REG_0_ | ~new_U3970;
  assign new_U5839 = ~new_U4046 | ~new_U4214;
  assign new_U5840 = ~DATAI_1_ | ~new_U3969;
  assign new_U5841 = ~new_U4027 | ~new_U3443;
  assign new_U5842 = ~new_U3468;
  assign new_U5843 = ~REG0_REG_1_ | ~new_U3970;
  assign new_U5844 = ~new_U4046 | ~new_U4238;
  assign new_U5845 = ~DATAI_2_ | ~new_U3969;
  assign new_U5846 = ~new_U4027 | ~new_U3442;
  assign new_U5847 = ~new_U3470;
  assign new_U5848 = ~REG0_REG_2_ | ~new_U3970;
  assign new_U5849 = ~new_U4046 | ~new_U4257;
  assign new_U5850 = ~DATAI_3_ | ~new_U3969;
  assign new_U5851 = ~new_U4027 | ~new_U3441;
  assign new_U5852 = ~new_U3472;
  assign new_U5853 = ~REG0_REG_3_ | ~new_U3970;
  assign new_U5854 = ~new_U4046 | ~new_U4276;
  assign new_U5855 = ~DATAI_4_ | ~new_U3969;
  assign new_U5856 = ~new_U4027 | ~new_U3440;
  assign new_U5857 = ~new_U3474;
  assign new_U5858 = ~REG0_REG_4_ | ~new_U3970;
  assign new_U5859 = ~new_U4046 | ~new_U4295;
  assign new_U5860 = ~DATAI_5_ | ~new_U3969;
  assign new_U5861 = ~new_U4027 | ~new_U3439;
  assign new_U5862 = ~new_U3476;
  assign new_U5863 = ~REG0_REG_5_ | ~new_U3970;
  assign new_U5864 = ~new_U4046 | ~new_U4314;
  assign new_U5865 = ~DATAI_6_ | ~new_U3969;
  assign new_U5866 = ~new_U4027 | ~new_U3438;
  assign new_U5867 = ~new_U3478;
  assign new_U5868 = ~REG0_REG_6_ | ~new_U3970;
  assign new_U5869 = ~new_U4046 | ~new_U4333;
  assign new_U5870 = ~DATAI_7_ | ~new_U3969;
  assign new_U5871 = ~new_U4027 | ~new_U3437;
  assign new_U5872 = ~new_U3480;
  assign new_U5873 = ~REG0_REG_7_ | ~new_U3970;
  assign new_U5874 = ~new_U4046 | ~new_U4352;
  assign new_U5875 = ~DATAI_8_ | ~new_U3969;
  assign new_U5876 = ~new_U4027 | ~new_U3436;
  assign new_U5877 = ~new_U3482;
  assign new_U5878 = ~REG0_REG_8_ | ~new_U3970;
  assign new_U5879 = ~new_U4046 | ~new_U4371;
  assign new_U5880 = ~DATAI_9_ | ~new_U3969;
  assign new_U5881 = ~new_U4027 | ~new_U3435;
  assign new_U5882 = ~new_U3484;
  assign new_U5883 = ~REG0_REG_9_ | ~new_U3970;
  assign new_U5884 = ~new_U4046 | ~new_U4390;
  assign new_U5885 = ~DATAI_10_ | ~new_U3969;
  assign new_U5886 = ~new_U4027 | ~new_U3452;
  assign new_U5887 = ~new_U3486;
  assign new_U5888 = ~REG0_REG_10_ | ~new_U3970;
  assign new_U5889 = ~new_U4046 | ~new_U4409;
  assign new_U5890 = ~DATAI_11_ | ~new_U3969;
  assign new_U5891 = ~new_U4027 | ~new_U3451;
  assign new_U5892 = ~new_U3488;
  assign new_U5893 = ~REG0_REG_11_ | ~new_U3970;
  assign new_U5894 = ~new_U4046 | ~new_U4428;
  assign new_U5895 = ~DATAI_12_ | ~new_U3969;
  assign new_U5896 = ~new_U4027 | ~new_U3450;
  assign new_U5897 = ~new_U3490;
  assign new_U5898 = ~REG0_REG_12_ | ~new_U3970;
  assign new_U5899 = ~new_U4046 | ~new_U4447;
  assign new_U5900 = ~DATAI_13_ | ~new_U3969;
  assign new_U5901 = ~new_U4027 | ~new_U3449;
  assign new_U5902 = ~new_U3492;
  assign new_U5903 = ~REG0_REG_13_ | ~new_U3970;
  assign new_U5904 = ~new_U4046 | ~new_U4466;
  assign new_U5905 = ~DATAI_14_ | ~new_U3969;
  assign new_U5906 = ~new_U4027 | ~new_U3448;
  assign new_U5907 = ~new_U3494;
  assign new_U5908 = ~REG0_REG_14_ | ~new_U3970;
  assign new_U5909 = ~new_U4046 | ~new_U4485;
  assign new_U5910 = ~DATAI_15_ | ~new_U3969;
  assign new_U5911 = ~new_U4027 | ~new_U3447;
  assign new_U5912 = ~new_U3496;
  assign new_U5913 = ~REG0_REG_15_ | ~new_U3970;
  assign new_U5914 = ~new_U4046 | ~new_U4504;
  assign new_U5915 = ~DATAI_16_ | ~new_U3969;
  assign new_U5916 = ~new_U4027 | ~new_U3446;
  assign new_U5917 = ~new_U3498;
  assign new_U5918 = ~REG0_REG_16_ | ~new_U3970;
  assign new_U5919 = ~new_U4046 | ~new_U4523;
  assign new_U5920 = ~DATAI_17_ | ~new_U3969;
  assign new_U5921 = ~new_U4027 | ~new_U3445;
  assign new_U5922 = ~new_U3500;
  assign new_U5923 = ~REG0_REG_17_ | ~new_U3970;
  assign new_U5924 = ~new_U4046 | ~new_U4542;
  assign new_U5925 = ~DATAI_18_ | ~new_U3969;
  assign new_U5926 = ~new_U4027 | ~new_U3444;
  assign new_U5927 = ~new_U3502;
  assign new_U5928 = ~REG0_REG_18_ | ~new_U3970;
  assign new_U5929 = ~new_U4046 | ~new_U4561;
  assign new_U5930 = ~DATAI_19_ | ~new_U3969;
  assign new_U5931 = ~new_U4027 | ~new_U3461;
  assign new_U5932 = ~new_U3504;
  assign new_U5933 = ~REG0_REG_19_ | ~new_U3970;
  assign new_U5934 = ~new_U4046 | ~new_U4580;
  assign new_U5935 = ~REG0_REG_20_ | ~new_U3970;
  assign new_U5936 = ~new_U4046 | ~new_U4599;
  assign new_U5937 = ~REG0_REG_21_ | ~new_U3970;
  assign new_U5938 = ~new_U4046 | ~new_U4618;
  assign new_U5939 = ~REG0_REG_22_ | ~new_U3970;
  assign new_U5940 = ~new_U4046 | ~new_U4637;
  assign new_U5941 = ~REG0_REG_23_ | ~new_U3970;
  assign new_U5942 = ~new_U4046 | ~new_U4656;
  assign new_U5943 = ~REG0_REG_24_ | ~new_U3970;
  assign new_U5944 = ~new_U4046 | ~new_U4675;
  assign new_U5945 = ~REG0_REG_25_ | ~new_U3970;
  assign new_U5946 = ~new_U4046 | ~new_U4694;
  assign new_U5947 = ~REG0_REG_26_ | ~new_U3970;
  assign new_U5948 = ~new_U4046 | ~new_U4713;
  assign new_U5949 = ~REG0_REG_27_ | ~new_U3970;
  assign new_U5950 = ~new_U4046 | ~new_U4732;
  assign new_U5951 = ~REG0_REG_28_ | ~new_U3970;
  assign new_U5952 = ~new_U4046 | ~new_U4751;
  assign new_U5953 = ~REG0_REG_29_ | ~new_U3970;
  assign new_U5954 = ~new_U4046 | ~new_U4771;
  assign new_U5955 = ~REG0_REG_30_ | ~new_U3970;
  assign new_U5956 = ~new_U4046 | ~new_U4778;
  assign new_U5957 = ~REG0_REG_31_ | ~new_U3970;
  assign new_U5958 = ~new_U4046 | ~new_U4781;
  assign new_U5959 = ~REG1_REG_0_ | ~new_U3971;
  assign new_U5960 = ~new_U4045 | ~new_U4214;
  assign new_U5961 = ~REG1_REG_1_ | ~new_U3971;
  assign new_U5962 = ~new_U4045 | ~new_U4238;
  assign new_U5963 = ~REG1_REG_2_ | ~new_U3971;
  assign new_U5964 = ~new_U4045 | ~new_U4257;
  assign new_U5965 = ~REG1_REG_3_ | ~new_U3971;
  assign new_U5966 = ~new_U4045 | ~new_U4276;
  assign new_U5967 = ~REG1_REG_4_ | ~new_U3971;
  assign new_U5968 = ~new_U4045 | ~new_U4295;
  assign new_U5969 = ~REG1_REG_5_ | ~new_U3971;
  assign new_U5970 = ~new_U4045 | ~new_U4314;
  assign new_U5971 = ~REG1_REG_6_ | ~new_U3971;
  assign new_U5972 = ~new_U4045 | ~new_U4333;
  assign new_U5973 = ~REG1_REG_7_ | ~new_U3971;
  assign new_U5974 = ~new_U4045 | ~new_U4352;
  assign new_U5975 = ~REG1_REG_8_ | ~new_U3971;
  assign new_U5976 = ~new_U4045 | ~new_U4371;
  assign new_U5977 = ~REG1_REG_9_ | ~new_U3971;
  assign new_U5978 = ~new_U4045 | ~new_U4390;
  assign new_U5979 = ~REG1_REG_10_ | ~new_U3971;
  assign new_U5980 = ~new_U4045 | ~new_U4409;
  assign new_U5981 = ~REG1_REG_11_ | ~new_U3971;
  assign new_U5982 = ~new_U4045 | ~new_U4428;
  assign new_U5983 = ~REG1_REG_12_ | ~new_U3971;
  assign new_U5984 = ~new_U4045 | ~new_U4447;
  assign new_U5985 = ~REG1_REG_13_ | ~new_U3971;
  assign new_U5986 = ~new_U4045 | ~new_U4466;
  assign new_U5987 = ~REG1_REG_14_ | ~new_U3971;
  assign new_U5988 = ~new_U4045 | ~new_U4485;
  assign new_U5989 = ~REG1_REG_15_ | ~new_U3971;
  assign new_U5990 = ~new_U4045 | ~new_U4504;
  assign new_U5991 = ~REG1_REG_16_ | ~new_U3971;
  assign new_U5992 = ~new_U4045 | ~new_U4523;
  assign new_U5993 = ~REG1_REG_17_ | ~new_U3971;
  assign new_U5994 = ~new_U4045 | ~new_U4542;
  assign new_U5995 = ~REG1_REG_18_ | ~new_U3971;
  assign new_U5996 = ~new_U4045 | ~new_U4561;
  assign new_U5997 = ~REG1_REG_19_ | ~new_U3971;
  assign new_U5998 = ~new_U4045 | ~new_U4580;
  assign new_U5999 = ~REG1_REG_20_ | ~new_U3971;
  assign new_U6000 = ~new_U4045 | ~new_U4599;
  assign new_U6001 = ~REG1_REG_21_ | ~new_U3971;
  assign new_U6002 = ~new_U4045 | ~new_U4618;
  assign new_U6003 = ~REG1_REG_22_ | ~new_U3971;
  assign new_U6004 = ~new_U4045 | ~new_U4637;
  assign new_U6005 = ~REG1_REG_23_ | ~new_U3971;
  assign new_U6006 = ~new_U4045 | ~new_U4656;
  assign new_U6007 = ~REG1_REG_24_ | ~new_U3971;
  assign new_U6008 = ~new_U4045 | ~new_U4675;
  assign new_U6009 = ~REG1_REG_25_ | ~new_U3971;
  assign new_U6010 = ~new_U4045 | ~new_U4694;
  assign new_U6011 = ~REG1_REG_26_ | ~new_U3971;
  assign new_U6012 = ~new_U4045 | ~new_U4713;
  assign new_U6013 = ~REG1_REG_27_ | ~new_U3971;
  assign new_U6014 = ~new_U4045 | ~new_U4732;
  assign new_U6015 = ~REG1_REG_28_ | ~new_U3971;
  assign new_U6016 = ~new_U4045 | ~new_U4751;
  assign new_U6017 = ~REG1_REG_29_ | ~new_U3971;
  assign new_U6018 = ~new_U4045 | ~new_U4771;
  assign new_U6019 = ~REG1_REG_30_ | ~new_U3971;
  assign new_U6020 = ~new_U4045 | ~new_U4778;
  assign new_U6021 = ~REG1_REG_31_ | ~new_U3971;
  assign new_U6022 = ~new_U4045 | ~new_U4781;
  assign new_U6023 = ~REG2_REG_0_ | ~new_U3417;
  assign new_U6024 = ~new_U4044 | ~new_U3375;
  assign new_U6025 = ~REG2_REG_1_ | ~new_U3417;
  assign new_U6026 = ~new_U4044 | ~new_U3377;
  assign new_U6027 = ~REG2_REG_2_ | ~new_U3417;
  assign new_U6028 = ~new_U4044 | ~new_U3378;
  assign new_U6029 = ~REG2_REG_3_ | ~new_U3417;
  assign new_U6030 = ~new_U4044 | ~new_U3379;
  assign new_U6031 = ~REG2_REG_4_ | ~new_U3417;
  assign new_U6032 = ~new_U4044 | ~new_U3380;
  assign new_U6033 = ~REG2_REG_5_ | ~new_U3417;
  assign new_U6034 = ~new_U4044 | ~new_U3381;
  assign new_U6035 = ~REG2_REG_6_ | ~new_U3417;
  assign new_U6036 = ~new_U4044 | ~new_U3382;
  assign new_U6037 = ~REG2_REG_7_ | ~new_U3417;
  assign new_U6038 = ~new_U4044 | ~new_U3383;
  assign new_U6039 = ~REG2_REG_8_ | ~new_U3417;
  assign new_U6040 = ~new_U4044 | ~new_U3384;
  assign new_U6041 = ~REG2_REG_9_ | ~new_U3417;
  assign new_U6042 = ~new_U4044 | ~new_U3385;
  assign new_U6043 = ~REG2_REG_10_ | ~new_U3417;
  assign new_U6044 = ~new_U4044 | ~new_U3386;
  assign new_U6045 = ~REG2_REG_11_ | ~new_U3417;
  assign new_U6046 = ~new_U4044 | ~new_U3387;
  assign new_U6047 = ~REG2_REG_12_ | ~new_U3417;
  assign new_U6048 = ~new_U4044 | ~new_U3388;
  assign new_U6049 = ~REG2_REG_13_ | ~new_U3417;
  assign new_U6050 = ~new_U4044 | ~new_U3389;
  assign new_U6051 = ~REG2_REG_14_ | ~new_U3417;
  assign new_U6052 = ~new_U4044 | ~new_U3390;
  assign new_U6053 = ~REG2_REG_15_ | ~new_U3417;
  assign new_U6054 = ~new_U4044 | ~new_U3391;
  assign new_U6055 = ~REG2_REG_16_ | ~new_U3417;
  assign new_U6056 = ~new_U4044 | ~new_U3392;
  assign new_U6057 = ~REG2_REG_17_ | ~new_U3417;
  assign new_U6058 = ~new_U4044 | ~new_U3393;
  assign new_U6059 = ~REG2_REG_18_ | ~new_U3417;
  assign new_U6060 = ~new_U4044 | ~new_U3394;
  assign new_U6061 = ~REG2_REG_19_ | ~new_U3417;
  assign new_U6062 = ~new_U4044 | ~new_U3395;
  assign new_U6063 = ~REG2_REG_20_ | ~new_U3417;
  assign new_U6064 = ~new_U4044 | ~new_U3397;
  assign new_U6065 = ~REG2_REG_21_ | ~new_U3417;
  assign new_U6066 = ~new_U4044 | ~new_U3399;
  assign new_U6067 = ~REG2_REG_22_ | ~new_U3417;
  assign new_U6068 = ~new_U4044 | ~new_U3401;
  assign new_U6069 = ~REG2_REG_23_ | ~new_U3417;
  assign new_U6070 = ~new_U4044 | ~new_U3403;
  assign new_U6071 = ~REG2_REG_24_ | ~new_U3417;
  assign new_U6072 = ~new_U4044 | ~new_U3405;
  assign new_U6073 = ~REG2_REG_25_ | ~new_U3417;
  assign new_U6074 = ~new_U4044 | ~new_U3407;
  assign new_U6075 = ~REG2_REG_26_ | ~new_U3417;
  assign new_U6076 = ~new_U4044 | ~new_U3409;
  assign new_U6077 = ~REG2_REG_27_ | ~new_U3417;
  assign new_U6078 = ~new_U4044 | ~new_U3411;
  assign new_U6079 = ~REG2_REG_28_ | ~new_U3417;
  assign new_U6080 = ~new_U4044 | ~new_U3413;
  assign new_U6081 = ~REG2_REG_29_ | ~new_U3417;
  assign new_U6082 = ~new_U4044 | ~new_U4767;
  assign new_U6083 = ~REG2_REG_30_ | ~new_U3417;
  assign new_U6084 = ~new_U4048 | ~new_U4044;
  assign new_U6085 = ~REG2_REG_31_ | ~new_U3417;
  assign new_U6086 = ~new_U4048 | ~new_U4044;
  assign new_U6087 = ~DATAO_REG_0_ | ~new_U3422;
  assign new_U6088 = ~n1351 | ~new_U3074;
  assign new_U6089 = ~DATAO_REG_1_ | ~new_U3422;
  assign new_U6090 = ~n1351 | ~new_U3075;
  assign new_U6091 = ~DATAO_REG_2_ | ~new_U3422;
  assign new_U6092 = ~n1351 | ~new_U3065;
  assign new_U6093 = ~DATAO_REG_3_ | ~new_U3422;
  assign new_U6094 = ~n1351 | ~new_U3061;
  assign new_U6095 = ~DATAO_REG_4_ | ~new_U3422;
  assign new_U6096 = ~n1351 | ~new_U3057;
  assign new_U6097 = ~DATAO_REG_5_ | ~new_U3422;
  assign new_U6098 = ~n1351 | ~new_U3064;
  assign new_U6099 = ~DATAO_REG_6_ | ~new_U3422;
  assign new_U6100 = ~n1351 | ~new_U3068;
  assign new_U6101 = ~DATAO_REG_7_ | ~new_U3422;
  assign new_U6102 = ~n1351 | ~new_U3067;
  assign new_U6103 = ~DATAO_REG_8_ | ~new_U3422;
  assign new_U6104 = ~n1351 | ~new_U3081;
  assign new_U6105 = ~DATAO_REG_9_ | ~new_U3422;
  assign new_U6106 = ~n1351 | ~new_U3080;
  assign new_U6107 = ~DATAO_REG_10_ | ~new_U3422;
  assign new_U6108 = ~n1351 | ~new_U3059;
  assign new_U6109 = ~DATAO_REG_11_ | ~new_U3422;
  assign new_U6110 = ~n1351 | ~new_U3060;
  assign new_U6111 = ~DATAO_REG_12_ | ~new_U3422;
  assign new_U6112 = ~n1351 | ~new_U3069;
  assign new_U6113 = ~DATAO_REG_13_ | ~new_U3422;
  assign new_U6114 = ~n1351 | ~new_U3077;
  assign new_U6115 = ~DATAO_REG_14_ | ~new_U3422;
  assign new_U6116 = ~n1351 | ~new_U3076;
  assign new_U6117 = ~DATAO_REG_15_ | ~new_U3422;
  assign new_U6118 = ~n1351 | ~new_U3071;
  assign new_U6119 = ~DATAO_REG_16_ | ~new_U3422;
  assign new_U6120 = ~n1351 | ~new_U3070;
  assign new_U6121 = ~DATAO_REG_17_ | ~new_U3422;
  assign new_U6122 = ~n1351 | ~new_U3066;
  assign new_U6123 = ~DATAO_REG_18_ | ~new_U3422;
  assign new_U6124 = ~n1351 | ~new_U3079;
  assign new_U6125 = ~DATAO_REG_19_ | ~new_U3422;
  assign new_U6126 = ~n1351 | ~new_U3078;
  assign new_U6127 = ~DATAO_REG_20_ | ~new_U3422;
  assign new_U6128 = ~n1351 | ~new_U3073;
  assign new_U6129 = ~DATAO_REG_21_ | ~new_U3422;
  assign new_U6130 = ~n1351 | ~new_U3072;
  assign new_U6131 = ~DATAO_REG_22_ | ~new_U3422;
  assign new_U6132 = ~n1351 | ~new_U3058;
  assign new_U6133 = ~DATAO_REG_23_ | ~new_U3422;
  assign new_U6134 = ~n1351 | ~new_U3063;
  assign new_U6135 = ~DATAO_REG_24_ | ~new_U3422;
  assign new_U6136 = ~n1351 | ~new_U3062;
  assign new_U6137 = ~DATAO_REG_25_ | ~new_U3422;
  assign new_U6138 = ~n1351 | ~new_U3055;
  assign new_U6139 = ~DATAO_REG_26_ | ~new_U3422;
  assign new_U6140 = ~n1351 | ~new_U3054;
  assign new_U6141 = ~DATAO_REG_27_ | ~new_U3422;
  assign new_U6142 = ~n1351 | ~new_U3050;
  assign new_U6143 = ~DATAO_REG_28_ | ~new_U3422;
  assign new_U6144 = ~n1351 | ~new_U3051;
  assign new_U6145 = ~DATAO_REG_29_ | ~new_U3422;
  assign new_U6146 = ~n1351 | ~new_U3052;
  assign new_U6147 = ~DATAO_REG_30_ | ~new_U3422;
  assign new_U6148 = ~n1351 | ~new_U3056;
  assign new_U6149 = ~DATAO_REG_31_ | ~new_U3422;
  assign new_U6150 = ~n1351 | ~new_U3053;
  assign new_U6151 = ~new_U4040 | ~new_U3052;
  assign new_U6152 = ~new_U3414 | ~new_U4737;
  assign new_U6153 = ~new_U6152 | ~new_U6151;
  assign new_U6154 = ~new_U4038 | ~new_U3053;
  assign new_U6155 = ~new_U3416 | ~new_U4775;
  assign new_U6156 = ~new_U6155 | ~new_U6154;
  assign new_U6157 = ~new_U4039 | ~new_U3056;
  assign new_U6158 = ~new_U3415 | ~new_U4755;
  assign new_U6159 = ~new_U6158 | ~new_U6157;
  assign new_U6160 = ~new_U4037 | ~new_U3073;
  assign new_U6161 = ~new_U3396 | ~new_U4566;
  assign new_U6162 = ~new_U6161 | ~new_U6160;
  assign new_U6163 = ~new_U5892 | ~new_U4395;
  assign new_U6164 = ~new_U3488 | ~new_U3060;
  assign new_U6165 = ~new_U6164 | ~new_U6163;
  assign new_U6166 = ~new_U5887 | ~new_U4376;
  assign new_U6167 = ~new_U3486 | ~new_U3059;
  assign new_U6168 = ~new_U6167 | ~new_U6166;
  assign new_U6169 = ~new_U5857 | ~new_U4262;
  assign new_U6170 = ~new_U3474 | ~new_U3057;
  assign new_U6171 = ~new_U6170 | ~new_U6169;
  assign new_U6172 = ~new_U5932 | ~new_U4547;
  assign new_U6173 = ~new_U3504 | ~new_U3078;
  assign new_U6174 = ~new_U6173 | ~new_U6172;
  assign new_U6175 = ~new_U4032 | ~new_U3055;
  assign new_U6176 = ~new_U3406 | ~new_U4661;
  assign new_U6177 = ~new_U6176 | ~new_U6175;
  assign new_U6178 = ~new_U4031 | ~new_U3054;
  assign new_U6179 = ~new_U3408 | ~new_U4680;
  assign new_U6180 = ~new_U6179 | ~new_U6178;
  assign new_U6181 = ~new_U4036 | ~new_U3072;
  assign new_U6182 = ~new_U3398 | ~new_U4585;
  assign new_U6183 = ~new_U6182 | ~new_U6181;
  assign new_U6184 = ~new_U4035 | ~new_U3058;
  assign new_U6185 = ~new_U3400 | ~new_U4604;
  assign new_U6186 = ~new_U6185 | ~new_U6184;
  assign new_U6187 = ~new_U4034 | ~new_U3063;
  assign new_U6188 = ~new_U3402 | ~new_U4623;
  assign new_U6189 = ~new_U6188 | ~new_U6187;
  assign new_U6190 = ~new_U4033 | ~new_U3062;
  assign new_U6191 = ~new_U3404 | ~new_U4642;
  assign new_U6192 = ~new_U6191 | ~new_U6190;
  assign new_U6193 = ~new_U4030 | ~new_U3050;
  assign new_U6194 = ~new_U3410 | ~new_U4699;
  assign new_U6195 = ~new_U6194 | ~new_U6193;
  assign new_U6196 = ~new_U4029 | ~new_U3051;
  assign new_U6197 = ~new_U3412 | ~new_U4718;
  assign new_U6198 = ~new_U6197 | ~new_U6196;
  assign new_U6199 = ~new_U5877 | ~new_U4338;
  assign new_U6200 = ~new_U3482 | ~new_U3081;
  assign new_U6201 = ~new_U6200 | ~new_U6199;
  assign new_U6202 = ~new_U5882 | ~new_U4357;
  assign new_U6203 = ~new_U3484 | ~new_U3080;
  assign new_U6204 = ~new_U6203 | ~new_U6202;
  assign new_U6205 = ~new_U5927 | ~new_U4528;
  assign new_U6206 = ~new_U3502 | ~new_U3079;
  assign new_U6207 = ~new_U6206 | ~new_U6205;
  assign new_U6208 = ~new_U5902 | ~new_U4433;
  assign new_U6209 = ~new_U3492 | ~new_U3077;
  assign new_U6210 = ~new_U6209 | ~new_U6208;
  assign new_U6211 = ~new_U5907 | ~new_U4452;
  assign new_U6212 = ~new_U3494 | ~new_U3076;
  assign new_U6213 = ~new_U6212 | ~new_U6211;
  assign new_U6214 = ~new_U5842 | ~new_U4200;
  assign new_U6215 = ~new_U3468 | ~new_U3075;
  assign new_U6216 = ~new_U6215 | ~new_U6214;
  assign new_U6217 = ~new_U5829 | ~new_U4224;
  assign new_U6218 = ~new_U3464 | ~new_U3074;
  assign new_U6219 = ~new_U6218 | ~new_U6217;
  assign new_U6220 = ~new_U5912 | ~new_U4471;
  assign new_U6221 = ~new_U3496 | ~new_U3071;
  assign new_U6222 = ~new_U6221 | ~new_U6220;
  assign new_U6223 = ~new_U5917 | ~new_U4490;
  assign new_U6224 = ~new_U3498 | ~new_U3070;
  assign new_U6225 = ~new_U6224 | ~new_U6223;
  assign new_U6226 = ~new_U5897 | ~new_U4414;
  assign new_U6227 = ~new_U3490 | ~new_U3069;
  assign new_U6228 = ~new_U6227 | ~new_U6226;
  assign new_U6229 = ~new_U5867 | ~new_U4300;
  assign new_U6230 = ~new_U3478 | ~new_U3068;
  assign new_U6231 = ~new_U6230 | ~new_U6229;
  assign new_U6232 = ~new_U5872 | ~new_U4319;
  assign new_U6233 = ~new_U3480 | ~new_U3067;
  assign new_U6234 = ~new_U6233 | ~new_U6232;
  assign new_U6235 = ~new_U5922 | ~new_U4509;
  assign new_U6236 = ~new_U3500 | ~new_U3066;
  assign new_U6237 = ~new_U6236 | ~new_U6235;
  assign new_U6238 = ~new_U5847 | ~new_U4219;
  assign new_U6239 = ~new_U3470 | ~new_U3065;
  assign new_U6240 = ~new_U6239 | ~new_U6238;
  assign new_U6241 = ~new_U5862 | ~new_U4281;
  assign new_U6242 = ~new_U3476 | ~new_U3064;
  assign new_U6243 = ~new_U6242 | ~new_U6241;
  assign new_U6244 = ~new_U5852 | ~new_U4243;
  assign new_U6245 = ~new_U3472 | ~new_U3061;
  assign new_U6246 = ~new_U6245 | ~new_U6244;
  assign new_U6247 = ~new_U4042 | ~new_U3424;
  assign new_U6248 = ~new_R1375_U26 | ~new_U3373;
  assign new_U6249 = ~new_U6248 | ~new_U6247;
  assign new_U6250 = ~new_U6249 | ~new_U5820;
  assign new_U6251 = ~new_U3460 | ~new_R395_U6 | ~new_U4042;
  assign new_U6252 = ~new_U5817 | ~new_U5139;
  assign new_U6253 = ~new_U3461 | ~new_U4055 | ~new_U3425;
  assign new_U6254 = ~new_U4014 | ~new_U4007;
  assign new_U6255 = ~new_U4023 | ~new_R1347_U13;
  assign new_U6256 = ~new_U5748 | ~new_U3423;
  assign new_U6257 = ~new_U3456 | ~new_U3431;
  assign new_U6258 = ~new_U3453 | ~new_U5421;
  assign new_U6259 = ~new_U5796 | ~new_U3016 | ~REG2_REG_0_;
  assign new_U6260 = ~new_U3080 | ~new_R1352_U6;
  assign new_U6261 = ~new_U3080 | ~new_U4009;
  assign new_U6262 = ~new_U3081 | ~new_R1352_U6;
  assign new_U6263 = ~new_U3081 | ~new_U4009;
  assign new_U6264 = ~new_U3067 | ~new_R1352_U6;
  assign new_U6265 = ~new_U3067 | ~new_U4009;
  assign new_U6266 = ~new_U3068 | ~new_R1352_U6;
  assign new_U6267 = ~new_U3068 | ~new_U4009;
  assign new_U6268 = ~new_U3064 | ~new_R1352_U6;
  assign new_U6269 = ~new_U3064 | ~new_U4009;
  assign new_U6270 = ~new_U3057 | ~new_R1352_U6;
  assign new_U6271 = ~new_U3057 | ~new_U4009;
  assign new_U6272 = ~new_R1309_U8 | ~new_R1352_U6;
  assign new_U6273 = ~new_U3053 | ~new_U4009;
  assign new_U6274 = ~new_R1309_U6 | ~new_R1352_U6;
  assign new_U6275 = ~new_U3056 | ~new_U4009;
  assign new_U6276 = ~new_U3061 | ~new_R1352_U6;
  assign new_U6277 = ~new_U3061 | ~new_U4009;
  assign new_U6278 = ~new_U3052 | ~new_R1352_U6;
  assign new_U6279 = ~new_U3052 | ~new_U4009;
  assign new_U6280 = ~new_U3051 | ~new_R1352_U6;
  assign new_U6281 = ~new_U3051 | ~new_U4009;
  assign new_U6282 = ~new_U3050 | ~new_R1352_U6;
  assign new_U6283 = ~new_U3050 | ~new_U4009;
  assign new_U6284 = ~new_U3054 | ~new_R1352_U6;
  assign new_U6285 = ~new_U3054 | ~new_U4009;
  assign new_U6286 = ~new_U3055 | ~new_R1352_U6;
  assign new_U6287 = ~new_U3055 | ~new_U4009;
  assign new_U6288 = ~new_U3062 | ~new_R1352_U6;
  assign new_U6289 = ~new_U3062 | ~new_U4009;
  assign new_U6290 = ~new_U3063 | ~new_R1352_U6;
  assign new_U6291 = ~new_U3063 | ~new_U4009;
  assign new_U6292 = ~new_U3058 | ~new_R1352_U6;
  assign new_U6293 = ~new_U3058 | ~new_U4009;
  assign new_U6294 = ~new_U3072 | ~new_R1352_U6;
  assign new_U6295 = ~new_U3072 | ~new_U4009;
  assign new_U6296 = ~new_U3073 | ~new_R1352_U6;
  assign new_U6297 = ~new_U3073 | ~new_U4009;
  assign new_U6298 = ~new_U3065 | ~new_R1352_U6;
  assign new_U6299 = ~new_U3065 | ~new_U4009;
  assign new_U6300 = ~new_U3078 | ~new_R1352_U6;
  assign new_U6301 = ~new_U3078 | ~new_U4009;
  assign new_U6302 = ~new_U3079 | ~new_R1352_U6;
  assign new_U6303 = ~new_U3079 | ~new_U4009;
  assign new_U6304 = ~new_U3066 | ~new_R1352_U6;
  assign new_U6305 = ~new_U3066 | ~new_U4009;
  assign new_U6306 = ~new_U3070 | ~new_R1352_U6;
  assign new_U6307 = ~new_U3070 | ~new_U4009;
  assign new_U6308 = ~new_U3071 | ~new_R1352_U6;
  assign new_U6309 = ~new_U3071 | ~new_U4009;
  assign new_U6310 = ~new_U3076 | ~new_R1352_U6;
  assign new_U6311 = ~new_U3076 | ~new_U4009;
  assign new_U6312 = ~new_U3077 | ~new_R1352_U6;
  assign new_U6313 = ~new_U3077 | ~new_U4009;
  assign new_U6314 = ~new_U3069 | ~new_R1352_U6;
  assign new_U6315 = ~new_U3069 | ~new_U4009;
  assign new_U6316 = ~new_U3060 | ~new_R1352_U6;
  assign new_U6317 = ~new_U3060 | ~new_U4009;
  assign new_U6318 = ~new_U3059 | ~new_R1352_U6;
  assign new_U6319 = ~new_U3059 | ~new_U4009;
  assign new_U6320 = ~new_U3075 | ~new_R1352_U6;
  assign new_U6321 = ~new_U3075 | ~new_U4009;
  assign new_U6322 = ~new_U3074 | ~new_R1352_U6;
  assign new_U6323 = ~new_U3074 | ~new_U4009;
  assign new_R1222_U516 = ~new_U3059 | ~new_R1222_U70;
  assign new_R1222_U515 = ~new_R1222_U378 | ~new_R1222_U513;
  assign new_R1222_U514 = ~new_R1222_U179 | ~new_R1222_U359;
  assign new_R1222_U513 = ~new_R1222_U512 | ~new_R1222_U511;
  assign new_R1222_U512 = ~new_U3488 | ~new_R1222_U75;
  assign new_R1222_U511 = ~new_U3060 | ~new_R1222_U74;
  assign new_R1222_U510 = ~new_R1222_U508 | ~new_R1222_U334;
  assign new_R1222_U509 = ~new_R1222_U358 | ~new_R1222_U102;
  assign new_R1222_U508 = ~new_R1222_U507 | ~new_R1222_U506;
  assign new_R1222_U507 = ~new_U3490 | ~new_R1222_U73;
  assign new_R1222_U506 = ~new_U3069 | ~new_R1222_U72;
  assign new_R1222_U505 = ~new_U3492 | ~new_R1222_U78;
  assign new_R1222_U504 = ~new_U3077 | ~new_R1222_U77;
  assign new_R1222_U503 = ~new_R1222_U254 | ~new_R1222_U501;
  assign new_R1222_U502 = ~new_R1222_U177 | ~new_R1222_U178;
  assign new_R1222_U501 = ~new_R1222_U500 | ~new_R1222_U499;
  assign new_R1222_U500 = ~new_U3494 | ~new_R1222_U80;
  assign new_R1222_U499 = ~new_U3076 | ~new_R1222_U79;
  assign new_R1222_U498 = ~new_U3494 | ~new_R1222_U80;
  assign new_R1222_U497 = ~new_U3076 | ~new_R1222_U79;
  assign new_R1222_U496 = ~new_R1222_U257 | ~new_R1222_U494;
  assign new_R1222_U495 = ~new_R1222_U175 | ~new_R1222_U176;
  assign new_SUB_84_U4 = ~IR_REG_25_ & ~IR_REG_24_ & ~IR_REG_26_ & ~IR_REG_27_;
  assign new_SUB_84_U5 = new_SUB_84_U55 & new_SUB_84_U54;
  assign new_SUB_84_U6 = new_SUB_84_U138 & new_SUB_84_U103;
  assign new_SUB_84_U7 = new_SUB_84_U137 & new_SUB_84_U46;
  assign new_SUB_84_U8 = new_SUB_84_U136 & new_SUB_84_U32;
  assign new_SUB_84_U9 = new_SUB_84_U134 & new_SUB_84_U106;
  assign new_SUB_84_U10 = new_SUB_84_U133 & new_SUB_84_U43;
  assign new_SUB_84_U11 = new_SUB_84_U132 & new_SUB_84_U38;
  assign new_SUB_84_U12 = new_SUB_84_U130 & new_SUB_84_U122;
  assign new_SUB_84_U13 = new_SUB_84_U129 & new_SUB_84_U39;
  assign new_SUB_84_U14 = new_SUB_84_U128 & new_SUB_84_U40;
  assign new_SUB_84_U15 = new_SUB_84_U126 & new_SUB_84_U80;
  assign new_SUB_84_U16 = new_SUB_84_U120 & new_SUB_84_U36;
  assign new_SUB_84_U17 = new_SUB_84_U118 & new_SUB_84_U75;
  assign new_SUB_84_U18 = new_SUB_84_U115 & new_SUB_84_U109;
  assign new_SUB_84_U19 = new_SUB_84_U113 & new_SUB_84_U33;
  assign new_SUB_84_U20 = new_SUB_84_U112 & new_SUB_84_U29;
  assign new_SUB_84_U21 = new_SUB_84_U102 & new_SUB_84_U30;
  assign new_SUB_84_U22 = new_SUB_84_U101 & new_SUB_84_U26;
  assign new_SUB_84_U23 = new_SUB_84_U99 & new_SUB_84_U93;
  assign new_SUB_84_U24 = new_SUB_84_U98 & new_SUB_84_U27;
  assign new_SUB_84_U25 = new_SUB_84_U97 & new_SUB_84_U45;
  assign new_SUB_84_U26 = ~new_SUB_84_U51 | ~new_SUB_84_U50;
  assign new_SUB_84_U27 = ~new_SUB_84_U53 | ~new_SUB_84_U92;
  assign new_SUB_84_U28 = ~IR_REG_6_;
  assign new_SUB_84_U29 = IR_REG_2_ | IR_REG_1_ | IR_REG_0_;
  assign new_SUB_84_U30 = ~new_SUB_84_U90 | ~new_SUB_84_U31;
  assign new_SUB_84_U31 = ~IR_REG_3_;
  assign new_SUB_84_U32 = ~new_SUB_84_U56 | ~new_SUB_84_U57 | ~new_SUB_84_U59 | ~new_SUB_84_U58;
  assign new_SUB_84_U33 = ~new_SUB_84_U5 | ~new_SUB_84_U60 | ~new_SUB_84_U105 | ~new_SUB_84_U4;
  assign new_SUB_84_U34 = ~new_SUB_84_U105 | ~new_SUB_84_U5;
  assign new_SUB_84_U35 = ~IR_REG_28_;
  assign new_SUB_84_U36 = ~new_SUB_84_U61 | ~new_SUB_84_U108;
  assign new_SUB_84_U37 = ~IR_REG_26_;
  assign new_SUB_84_U38 = ~new_SUB_84_U62 | ~new_SUB_84_U105;
  assign new_SUB_84_U39 = ~new_SUB_84_U63 | ~new_SUB_84_U121;
  assign new_SUB_84_U40 = ~new_SUB_84_U64 | ~new_SUB_84_U123;
  assign new_SUB_84_U41 = ~IR_REG_22_;
  assign new_SUB_84_U42 = ~IR_REG_18_;
  assign new_SUB_84_U43 = ~new_SUB_84_U65 | ~new_SUB_84_U105;
  assign new_SUB_84_U44 = ~IR_REG_14_;
  assign new_SUB_84_U45 = ~new_SUB_84_U52 | ~new_SUB_84_U92;
  assign new_SUB_84_U46 = ~new_SUB_84_U66 | ~new_SUB_84_U95;
  assign new_SUB_84_U47 = ~IR_REG_10_;
  assign new_SUB_84_U48 = ~new_SUB_84_U157 | ~new_SUB_84_U156;
  assign new_SUB_84_U49 = ~new_SUB_84_U145 | ~new_SUB_84_U144;
  assign new_SUB_84_U50 = ~IR_REG_0_ & ~IR_REG_2_ & ~IR_REG_1_;
  assign new_SUB_84_U51 = ~IR_REG_4_ & ~IR_REG_5_ & ~IR_REG_3_;
  assign new_SUB_84_U52 = ~IR_REG_9_ & ~IR_REG_8_ & ~IR_REG_6_ & ~IR_REG_7_;
  assign new_SUB_84_U53 = ~IR_REG_6_ & ~IR_REG_7_;
  assign new_SUB_84_U54 = ~IR_REG_15_ & ~IR_REG_14_ & ~IR_REG_16_ & ~IR_REG_17_ & ~IR_REG_18_;
  assign new_SUB_84_U55 = ~IR_REG_20_ & ~IR_REG_19_ & ~IR_REG_21_ & ~IR_REG_22_ & ~IR_REG_23_;
  assign new_SUB_84_U56 = ~IR_REG_13_ & ~IR_REG_12_ & ~IR_REG_10_ & ~IR_REG_11_;
  assign new_SUB_84_U57 = ~IR_REG_0_ & ~IR_REG_2_ & ~IR_REG_1_;
  assign new_SUB_84_U58 = ~IR_REG_6_ & ~IR_REG_5_ & ~IR_REG_3_ & ~IR_REG_4_;
  assign new_SUB_84_U59 = ~IR_REG_8_ & ~IR_REG_9_ & ~IR_REG_7_;
  assign new_SUB_84_U60 = ~IR_REG_28_ & ~IR_REG_29_;
  assign new_SUB_84_U61 = ~IR_REG_24_ & ~IR_REG_25_;
  assign new_SUB_84_U62 = ~IR_REG_17_ & ~IR_REG_16_ & ~IR_REG_14_ & ~IR_REG_15_;
  assign new_SUB_84_U63 = ~IR_REG_18_ & ~IR_REG_19_;
  assign new_SUB_84_U64 = ~IR_REG_20_ & ~IR_REG_21_;
  assign new_SUB_84_U65 = ~IR_REG_14_ & ~IR_REG_15_;
  assign new_SUB_84_U66 = ~IR_REG_10_ & ~IR_REG_11_;
  assign new_SUB_84_U67 = ~IR_REG_8_;
  assign new_SUB_84_U68 = new_SUB_84_U141 & new_SUB_84_U140;
  assign new_SUB_84_U69 = ~IR_REG_4_;
  assign new_SUB_84_U70 = new_SUB_84_U143 & new_SUB_84_U142;
  assign new_SUB_84_U71 = ~IR_REG_31_;
  assign new_SUB_84_U72 = ~IR_REG_30_;
  assign new_SUB_84_U73 = new_SUB_84_U147 & new_SUB_84_U146;
  assign new_SUB_84_U74 = ~IR_REG_27_;
  assign new_SUB_84_U75 = ~new_SUB_84_U116 | ~new_SUB_84_U37;
  assign new_SUB_84_U76 = new_SUB_84_U149 & new_SUB_84_U148;
  assign new_SUB_84_U77 = ~IR_REG_24_;
  assign new_SUB_84_U78 = new_SUB_84_U151 & new_SUB_84_U150;
  assign new_SUB_84_U79 = ~IR_REG_23_;
  assign new_SUB_84_U80 = ~new_SUB_84_U124 | ~new_SUB_84_U41;
  assign new_SUB_84_U81 = new_SUB_84_U153 & new_SUB_84_U152;
  assign new_SUB_84_U82 = ~IR_REG_20_;
  assign new_SUB_84_U83 = new_SUB_84_U155 & new_SUB_84_U154;
  assign new_SUB_84_U84 = ~IR_REG_1_;
  assign new_SUB_84_U85 = ~IR_REG_0_;
  assign new_SUB_84_U86 = ~IR_REG_16_;
  assign new_SUB_84_U87 = new_SUB_84_U159 & new_SUB_84_U158;
  assign new_SUB_84_U88 = ~IR_REG_12_;
  assign new_SUB_84_U89 = new_SUB_84_U161 & new_SUB_84_U160;
  assign new_SUB_84_U90 = ~new_SUB_84_U29;
  assign new_SUB_84_U91 = ~new_SUB_84_U30;
  assign new_SUB_84_U92 = ~new_SUB_84_U26;
  assign new_SUB_84_U93 = ~new_SUB_84_U92 | ~new_SUB_84_U28;
  assign new_SUB_84_U94 = ~new_SUB_84_U27;
  assign new_SUB_84_U95 = ~new_SUB_84_U45;
  assign new_SUB_84_U96 = ~new_SUB_84_U94 | ~new_SUB_84_U67;
  assign new_SUB_84_U97 = ~IR_REG_9_ | ~new_SUB_84_U96;
  assign new_SUB_84_U98 = ~IR_REG_7_ | ~new_SUB_84_U93;
  assign new_SUB_84_U99 = ~IR_REG_6_ | ~new_SUB_84_U26;
  assign new_SUB_84_U100 = ~new_SUB_84_U91 | ~new_SUB_84_U69;
  assign new_SUB_84_U101 = ~IR_REG_5_ | ~new_SUB_84_U100;
  assign new_SUB_84_U102 = ~IR_REG_3_ | ~new_SUB_84_U29;
  assign new_SUB_84_U103 = ~new_SUB_84_U95 | ~new_SUB_84_U47;
  assign new_SUB_84_U104 = ~new_SUB_84_U46;
  assign new_SUB_84_U105 = ~new_SUB_84_U32;
  assign new_SUB_84_U106 = ~new_SUB_84_U105 | ~new_SUB_84_U44;
  assign new_SUB_84_U107 = ~new_SUB_84_U43;
  assign new_SUB_84_U108 = ~new_SUB_84_U34;
  assign new_SUB_84_U109 = ~new_SUB_84_U35 | ~new_SUB_84_U5 | ~new_SUB_84_U105 | ~new_SUB_84_U4;
  assign new_SUB_84_U110 = ~new_SUB_84_U33;
  assign new_SUB_84_U111 = IR_REG_1_ | IR_REG_0_;
  assign new_SUB_84_U112 = ~IR_REG_2_ | ~new_SUB_84_U111;
  assign new_SUB_84_U113 = ~IR_REG_29_ | ~new_SUB_84_U109;
  assign new_SUB_84_U114 = ~new_SUB_84_U108 | ~new_SUB_84_U4;
  assign new_SUB_84_U115 = ~IR_REG_28_ | ~new_SUB_84_U114;
  assign new_SUB_84_U116 = ~new_SUB_84_U36;
  assign new_SUB_84_U117 = ~new_SUB_84_U75;
  assign new_SUB_84_U118 = ~IR_REG_26_ | ~new_SUB_84_U36;
  assign new_SUB_84_U119 = ~new_SUB_84_U108 | ~new_SUB_84_U77;
  assign new_SUB_84_U120 = ~IR_REG_25_ | ~new_SUB_84_U119;
  assign new_SUB_84_U121 = ~new_SUB_84_U38;
  assign new_SUB_84_U122 = ~new_SUB_84_U121 | ~new_SUB_84_U42;
  assign new_SUB_84_U123 = ~new_SUB_84_U39;
  assign new_SUB_84_U124 = ~new_SUB_84_U40;
  assign new_SUB_84_U125 = ~new_SUB_84_U80;
  assign new_SUB_84_U126 = ~IR_REG_22_ | ~new_SUB_84_U40;
  assign new_SUB_84_U127 = ~new_SUB_84_U123 | ~new_SUB_84_U82;
  assign new_SUB_84_U128 = ~IR_REG_21_ | ~new_SUB_84_U127;
  assign new_SUB_84_U129 = ~IR_REG_19_ | ~new_SUB_84_U122;
  assign new_SUB_84_U130 = ~IR_REG_18_ | ~new_SUB_84_U38;
  assign new_SUB_84_U131 = ~new_SUB_84_U107 | ~new_SUB_84_U86;
  assign new_SUB_84_U132 = ~IR_REG_17_ | ~new_SUB_84_U131;
  assign new_SUB_84_U133 = ~IR_REG_15_ | ~new_SUB_84_U106;
  assign new_SUB_84_U134 = ~IR_REG_14_ | ~new_SUB_84_U32;
  assign new_SUB_84_U135 = ~new_SUB_84_U104 | ~new_SUB_84_U88;
  assign new_SUB_84_U136 = ~IR_REG_13_ | ~new_SUB_84_U135;
  assign new_SUB_84_U137 = ~IR_REG_11_ | ~new_SUB_84_U103;
  assign new_SUB_84_U138 = ~IR_REG_10_ | ~new_SUB_84_U45;
  assign new_SUB_84_U139 = ~new_SUB_84_U110 | ~new_SUB_84_U72;
  assign new_SUB_84_U140 = ~IR_REG_8_ | ~new_SUB_84_U27;
  assign new_SUB_84_U141 = ~new_SUB_84_U94 | ~new_SUB_84_U67;
  assign new_SUB_84_U142 = ~IR_REG_4_ | ~new_SUB_84_U30;
  assign new_SUB_84_U143 = ~new_SUB_84_U91 | ~new_SUB_84_U69;
  assign new_SUB_84_U144 = ~new_SUB_84_U139 | ~new_SUB_84_U71;
  assign new_SUB_84_U145 = ~IR_REG_31_ | ~new_SUB_84_U110 | ~new_SUB_84_U72;
  assign new_SUB_84_U146 = ~IR_REG_30_ | ~new_SUB_84_U33;
  assign new_SUB_84_U147 = ~new_SUB_84_U110 | ~new_SUB_84_U72;
  assign new_SUB_84_U148 = ~IR_REG_27_ | ~new_SUB_84_U75;
  assign new_SUB_84_U149 = ~new_SUB_84_U117 | ~new_SUB_84_U74;
  assign new_SUB_84_U150 = ~IR_REG_24_ | ~new_SUB_84_U34;
  assign new_SUB_84_U151 = ~new_SUB_84_U108 | ~new_SUB_84_U77;
  assign new_SUB_84_U152 = ~IR_REG_23_ | ~new_SUB_84_U80;
  assign new_SUB_84_U153 = ~new_SUB_84_U125 | ~new_SUB_84_U79;
  assign new_SUB_84_U154 = ~IR_REG_20_ | ~new_SUB_84_U39;
  assign new_SUB_84_U155 = ~new_SUB_84_U123 | ~new_SUB_84_U82;
  assign new_SUB_84_U156 = ~IR_REG_1_ | ~new_SUB_84_U85;
  assign new_SUB_84_U157 = ~IR_REG_0_ | ~new_SUB_84_U84;
  assign new_SUB_84_U158 = ~IR_REG_16_ | ~new_SUB_84_U43;
  assign new_SUB_84_U159 = ~new_SUB_84_U107 | ~new_SUB_84_U86;
  assign new_SUB_84_U160 = ~IR_REG_12_ | ~new_SUB_84_U46;
  assign new_SUB_84_U161 = ~new_SUB_84_U104 | ~new_SUB_84_U88;
  assign new_ADD_95_U4 = ~REG3_REG_3_;
  assign new_ADD_95_U5 = new_ADD_95_U76 & new_ADD_95_U107;
  assign new_ADD_95_U6 = ~REG3_REG_7_;
  assign new_ADD_95_U7 = ~REG3_REG_6_;
  assign new_ADD_95_U8 = ~REG3_REG_5_;
  assign new_ADD_95_U9 = ~REG3_REG_4_;
  assign new_ADD_95_U10 = ~REG3_REG_5_ | ~REG3_REG_4_ | ~REG3_REG_6_ | ~REG3_REG_7_ | ~REG3_REG_3_;
  assign new_ADD_95_U11 = ~REG3_REG_8_;
  assign new_ADD_95_U12 = ~REG3_REG_9_;
  assign new_ADD_95_U13 = ~new_ADD_95_U71 | ~new_ADD_95_U88;
  assign new_ADD_95_U14 = ~REG3_REG_11_;
  assign new_ADD_95_U15 = ~REG3_REG_10_;
  assign new_ADD_95_U16 = ~new_ADD_95_U72 | ~new_ADD_95_U90;
  assign new_ADD_95_U17 = ~REG3_REG_13_;
  assign new_ADD_95_U18 = ~REG3_REG_12_;
  assign new_ADD_95_U19 = ~new_ADD_95_U73 | ~new_ADD_95_U92;
  assign new_ADD_95_U20 = ~REG3_REG_15_;
  assign new_ADD_95_U21 = ~REG3_REG_14_;
  assign new_ADD_95_U22 = ~new_ADD_95_U74 | ~new_ADD_95_U94;
  assign new_ADD_95_U23 = ~REG3_REG_17_;
  assign new_ADD_95_U24 = ~REG3_REG_16_;
  assign new_ADD_95_U25 = ~new_ADD_95_U75 | ~new_ADD_95_U96;
  assign new_ADD_95_U26 = ~REG3_REG_18_;
  assign new_ADD_95_U27 = ~REG3_REG_18_ | ~new_ADD_95_U98;
  assign new_ADD_95_U28 = ~REG3_REG_19_;
  assign new_ADD_95_U29 = ~REG3_REG_19_ | ~new_ADD_95_U99;
  assign new_ADD_95_U30 = ~REG3_REG_20_;
  assign new_ADD_95_U31 = ~REG3_REG_20_ | ~new_ADD_95_U100;
  assign new_ADD_95_U32 = ~REG3_REG_21_;
  assign new_ADD_95_U33 = ~REG3_REG_21_ | ~new_ADD_95_U101;
  assign new_ADD_95_U34 = ~REG3_REG_22_;
  assign new_ADD_95_U35 = ~REG3_REG_22_ | ~new_ADD_95_U102;
  assign new_ADD_95_U36 = ~REG3_REG_23_;
  assign new_ADD_95_U37 = ~REG3_REG_23_ | ~new_ADD_95_U103;
  assign new_ADD_95_U38 = ~REG3_REG_24_;
  assign new_ADD_95_U39 = ~REG3_REG_24_ | ~new_ADD_95_U104;
  assign new_ADD_95_U40 = ~REG3_REG_25_;
  assign new_ADD_95_U41 = ~REG3_REG_25_ | ~new_ADD_95_U105;
  assign new_ADD_95_U42 = ~REG3_REG_26_;
  assign new_ADD_95_U43 = ~REG3_REG_26_ | ~new_ADD_95_U106;
  assign new_ADD_95_U44 = ~REG3_REG_28_;
  assign new_ADD_95_U45 = ~REG3_REG_27_;
  assign new_ADD_95_U46 = ~new_ADD_95_U111 | ~new_ADD_95_U110;
  assign new_ADD_95_U47 = ~new_ADD_95_U113 | ~new_ADD_95_U112;
  assign new_ADD_95_U48 = ~new_ADD_95_U115 | ~new_ADD_95_U114;
  assign new_ADD_95_U49 = ~new_ADD_95_U117 | ~new_ADD_95_U116;
  assign new_ADD_95_U50 = ~new_ADD_95_U119 | ~new_ADD_95_U118;
  assign new_ADD_95_U51 = ~new_ADD_95_U121 | ~new_ADD_95_U120;
  assign new_ADD_95_U52 = ~new_ADD_95_U123 | ~new_ADD_95_U122;
  assign new_ADD_95_U53 = ~new_ADD_95_U125 | ~new_ADD_95_U124;
  assign new_ADD_95_U54 = ~new_ADD_95_U127 | ~new_ADD_95_U126;
  assign new_ADD_95_U55 = ~new_ADD_95_U129 | ~new_ADD_95_U128;
  assign new_ADD_95_U56 = ~new_ADD_95_U131 | ~new_ADD_95_U130;
  assign new_ADD_95_U57 = ~new_ADD_95_U133 | ~new_ADD_95_U132;
  assign new_ADD_95_U58 = ~new_ADD_95_U135 | ~new_ADD_95_U134;
  assign new_ADD_95_U59 = ~new_ADD_95_U137 | ~new_ADD_95_U136;
  assign new_ADD_95_U60 = ~new_ADD_95_U139 | ~new_ADD_95_U138;
  assign new_ADD_95_U61 = ~new_ADD_95_U141 | ~new_ADD_95_U140;
  assign new_ADD_95_U62 = ~new_ADD_95_U143 | ~new_ADD_95_U142;
  assign new_ADD_95_U63 = ~new_ADD_95_U145 | ~new_ADD_95_U144;
  assign new_ADD_95_U64 = ~new_ADD_95_U147 | ~new_ADD_95_U146;
  assign new_ADD_95_U65 = ~new_ADD_95_U149 | ~new_ADD_95_U148;
  assign new_ADD_95_U66 = ~new_ADD_95_U151 | ~new_ADD_95_U150;
  assign new_ADD_95_U67 = ~new_ADD_95_U153 | ~new_ADD_95_U152;
  assign new_ADD_95_U68 = ~new_ADD_95_U155 | ~new_ADD_95_U154;
  assign new_ADD_95_U69 = ~new_ADD_95_U157 | ~new_ADD_95_U156;
  assign new_ADD_95_U70 = ~new_ADD_95_U159 | ~new_ADD_95_U158;
  assign new_ADD_95_U71 = REG3_REG_8_ & REG3_REG_9_;
  assign new_ADD_95_U72 = REG3_REG_11_ & REG3_REG_10_;
  assign new_ADD_95_U73 = REG3_REG_13_ & REG3_REG_12_;
  assign new_ADD_95_U74 = REG3_REG_15_ & REG3_REG_14_;
  assign new_ADD_95_U75 = REG3_REG_17_ & REG3_REG_16_;
  assign new_ADD_95_U76 = REG3_REG_28_ & REG3_REG_27_;
  assign new_ADD_95_U77 = ~REG3_REG_8_ | ~new_ADD_95_U88;
  assign new_ADD_95_U78 = ~REG3_REG_3_ | ~REG3_REG_6_ | ~REG3_REG_4_ | ~REG3_REG_5_;
  assign new_ADD_95_U79 = ~REG3_REG_4_ | ~REG3_REG_5_ | ~REG3_REG_3_;
  assign new_ADD_95_U80 = ~REG3_REG_4_ | ~REG3_REG_3_;
  assign new_ADD_95_U81 = ~REG3_REG_27_ | ~new_ADD_95_U107;
  assign new_ADD_95_U82 = ~REG3_REG_16_ | ~new_ADD_95_U96;
  assign new_ADD_95_U83 = ~REG3_REG_14_ | ~new_ADD_95_U94;
  assign new_ADD_95_U84 = ~REG3_REG_12_ | ~new_ADD_95_U92;
  assign new_ADD_95_U85 = ~REG3_REG_10_ | ~new_ADD_95_U90;
  assign new_ADD_95_U86 = ~new_ADD_95_U80;
  assign new_ADD_95_U87 = ~new_ADD_95_U78;
  assign new_ADD_95_U88 = ~new_ADD_95_U10;
  assign new_ADD_95_U89 = ~new_ADD_95_U77;
  assign new_ADD_95_U90 = ~new_ADD_95_U13;
  assign new_ADD_95_U91 = ~new_ADD_95_U85;
  assign new_ADD_95_U92 = ~new_ADD_95_U16;
  assign new_ADD_95_U93 = ~new_ADD_95_U84;
  assign new_ADD_95_U94 = ~new_ADD_95_U19;
  assign new_ADD_95_U95 = ~new_ADD_95_U83;
  assign new_ADD_95_U96 = ~new_ADD_95_U22;
  assign new_ADD_95_U97 = ~new_ADD_95_U82;
  assign new_ADD_95_U98 = ~new_ADD_95_U25;
  assign new_ADD_95_U99 = ~new_ADD_95_U27;
  assign new_ADD_95_U100 = ~new_ADD_95_U29;
  assign new_ADD_95_U101 = ~new_ADD_95_U31;
  assign new_ADD_95_U102 = ~new_ADD_95_U33;
  assign new_ADD_95_U103 = ~new_ADD_95_U35;
  assign new_ADD_95_U104 = ~new_ADD_95_U37;
  assign new_ADD_95_U105 = ~new_ADD_95_U39;
  assign new_ADD_95_U106 = ~new_ADD_95_U41;
  assign new_ADD_95_U107 = ~new_ADD_95_U43;
  assign new_ADD_95_U108 = ~new_ADD_95_U81;
  assign new_ADD_95_U109 = ~new_ADD_95_U79;
  assign new_ADD_95_U110 = ~REG3_REG_9_ | ~new_ADD_95_U77;
  assign new_ADD_95_U111 = ~new_ADD_95_U89 | ~new_ADD_95_U12;
  assign new_ADD_95_U112 = ~REG3_REG_8_ | ~new_ADD_95_U10;
  assign new_ADD_95_U113 = ~new_ADD_95_U88 | ~new_ADD_95_U11;
  assign new_ADD_95_U114 = ~REG3_REG_7_ | ~new_ADD_95_U78;
  assign new_ADD_95_U115 = ~new_ADD_95_U87 | ~new_ADD_95_U6;
  assign new_ADD_95_U116 = ~REG3_REG_6_ | ~new_ADD_95_U79;
  assign new_ADD_95_U117 = ~new_ADD_95_U109 | ~new_ADD_95_U7;
  assign new_ADD_95_U118 = ~REG3_REG_5_ | ~new_ADD_95_U80;
  assign new_ADD_95_U119 = ~new_ADD_95_U86 | ~new_ADD_95_U8;
  assign new_ADD_95_U120 = ~REG3_REG_4_ | ~new_ADD_95_U4;
  assign new_ADD_95_U121 = ~REG3_REG_3_ | ~new_ADD_95_U9;
  assign new_ADD_95_U122 = ~REG3_REG_28_ | ~new_ADD_95_U81;
  assign new_ADD_95_U123 = ~new_ADD_95_U108 | ~new_ADD_95_U44;
  assign new_ADD_95_U124 = ~REG3_REG_27_ | ~new_ADD_95_U43;
  assign new_ADD_95_U125 = ~new_ADD_95_U107 | ~new_ADD_95_U45;
  assign new_ADD_95_U126 = ~REG3_REG_26_ | ~new_ADD_95_U41;
  assign new_ADD_95_U127 = ~new_ADD_95_U106 | ~new_ADD_95_U42;
  assign new_ADD_95_U128 = ~REG3_REG_25_ | ~new_ADD_95_U39;
  assign new_ADD_95_U129 = ~new_ADD_95_U105 | ~new_ADD_95_U40;
  assign new_ADD_95_U130 = ~REG3_REG_24_ | ~new_ADD_95_U37;
  assign new_ADD_95_U131 = ~new_ADD_95_U104 | ~new_ADD_95_U38;
  assign new_ADD_95_U132 = ~REG3_REG_23_ | ~new_ADD_95_U35;
  assign new_ADD_95_U133 = ~new_ADD_95_U103 | ~new_ADD_95_U36;
  assign new_ADD_95_U134 = ~REG3_REG_22_ | ~new_ADD_95_U33;
  assign new_ADD_95_U135 = ~new_ADD_95_U102 | ~new_ADD_95_U34;
  assign new_ADD_95_U136 = ~REG3_REG_21_ | ~new_ADD_95_U31;
  assign new_ADD_95_U137 = ~new_ADD_95_U101 | ~new_ADD_95_U32;
  assign new_ADD_95_U138 = ~REG3_REG_20_ | ~new_ADD_95_U29;
  assign new_ADD_95_U139 = ~new_ADD_95_U100 | ~new_ADD_95_U30;
  assign new_ADD_95_U140 = ~REG3_REG_19_ | ~new_ADD_95_U27;
  assign new_ADD_95_U141 = ~new_ADD_95_U99 | ~new_ADD_95_U28;
  assign new_ADD_95_U142 = ~REG3_REG_18_ | ~new_ADD_95_U25;
  assign new_ADD_95_U143 = ~new_ADD_95_U98 | ~new_ADD_95_U26;
  assign new_ADD_95_U144 = ~REG3_REG_17_ | ~new_ADD_95_U82;
  assign new_ADD_95_U145 = ~new_ADD_95_U97 | ~new_ADD_95_U23;
  assign new_ADD_95_U146 = ~REG3_REG_16_ | ~new_ADD_95_U22;
  assign new_ADD_95_U147 = ~new_ADD_95_U96 | ~new_ADD_95_U24;
  assign new_ADD_95_U148 = ~REG3_REG_15_ | ~new_ADD_95_U83;
  assign new_ADD_95_U149 = ~new_ADD_95_U95 | ~new_ADD_95_U20;
  assign new_ADD_95_U150 = ~REG3_REG_14_ | ~new_ADD_95_U19;
  assign new_ADD_95_U151 = ~new_ADD_95_U94 | ~new_ADD_95_U21;
  assign new_ADD_95_U152 = ~REG3_REG_13_ | ~new_ADD_95_U84;
  assign new_ADD_95_U153 = ~new_ADD_95_U93 | ~new_ADD_95_U17;
  assign new_ADD_95_U154 = ~REG3_REG_12_ | ~new_ADD_95_U16;
  assign new_ADD_95_U155 = ~new_ADD_95_U92 | ~new_ADD_95_U18;
  assign new_ADD_95_U156 = ~REG3_REG_11_ | ~new_ADD_95_U85;
  assign new_ADD_95_U157 = ~new_ADD_95_U91 | ~new_ADD_95_U14;
  assign new_ADD_95_U158 = ~REG3_REG_10_ | ~new_ADD_95_U13;
  assign new_ADD_95_U159 = ~new_ADD_95_U90 | ~new_ADD_95_U15;
  assign new_R395_U6 = ~new_R395_U99 | ~new_R395_U183;
  assign new_R395_U7 = ~new_U3111;
  assign new_R395_U8 = ~new_U3110;
  assign new_R395_U9 = ~new_U3109;
  assign new_R395_U10 = ~new_U3143;
  assign new_R395_U11 = ~new_U3142;
  assign new_R395_U12 = ~new_U3141;
  assign new_R395_U13 = ~new_U3140;
  assign new_R395_U14 = ~new_U3139;
  assign new_R395_U15 = ~new_U3138;
  assign new_R395_U16 = ~new_U3108;
  assign new_R395_U17 = ~new_U3107;
  assign new_R395_U18 = ~new_U3106;
  assign new_R395_U19 = ~new_U3105;
  assign new_R395_U20 = ~new_U3104;
  assign new_R395_U21 = ~new_U3103;
  assign new_R395_U22 = ~new_U3137;
  assign new_R395_U23 = ~new_U3136;
  assign new_R395_U24 = ~new_U3135;
  assign new_R395_U25 = ~new_U3134;
  assign new_R395_U26 = ~new_U3133;
  assign new_R395_U27 = ~new_U3132;
  assign new_R395_U28 = ~new_U3102;
  assign new_R395_U29 = ~new_U3101;
  assign new_R395_U30 = ~new_U3100;
  assign new_R395_U31 = ~new_U3099;
  assign new_R395_U32 = ~new_U3131;
  assign new_R395_U33 = ~new_U3130;
  assign new_R395_U34 = ~new_U3098;
  assign new_R395_U35 = ~new_U3097;
  assign new_R395_U36 = ~new_U3129;
  assign new_R395_U37 = ~new_U3128;
  assign new_R395_U38 = ~new_U3096;
  assign new_R395_U39 = ~new_U3095;
  assign new_R395_U40 = ~new_U3127;
  assign new_R395_U41 = ~new_U3126;
  assign new_R395_U42 = ~new_U3094;
  assign new_R395_U43 = ~new_U3093;
  assign new_R395_U44 = ~new_U3125;
  assign new_R395_U45 = ~new_U3124;
  assign new_R395_U46 = ~new_U3092;
  assign new_R395_U47 = ~new_U3091;
  assign new_R395_U48 = ~new_U3123;
  assign new_R395_U49 = ~new_U3122;
  assign new_R395_U50 = ~new_U3090;
  assign new_R395_U51 = ~new_U3089;
  assign new_R395_U52 = ~new_U3121;
  assign new_R395_U53 = ~new_U3120;
  assign new_R395_U54 = ~new_U3088;
  assign new_R395_U55 = ~new_U3087;
  assign new_R395_U56 = ~new_U3119;
  assign new_R395_U57 = ~new_U3118;
  assign new_R395_U58 = ~new_U3086;
  assign new_R395_U59 = ~new_U3085;
  assign new_R395_U60 = ~new_U3117;
  assign new_R395_U61 = ~new_U3116;
  assign new_R395_U62 = ~new_U3084;
  assign new_R395_U63 = ~new_U3083;
  assign new_R395_U64 = ~new_U3115;
  assign new_R395_U65 = ~new_U3114;
  assign new_R395_U66 = ~new_U3146;
  assign new_R395_U67 = new_R395_U102 & new_R395_U103 & new_R395_U104;
  assign new_R395_U68 = new_R395_U184 & new_R395_U109 & new_R395_U108;
  assign new_R395_U69 = new_U3142 & new_R395_U8;
  assign new_R395_U70 = new_R395_U106 & new_R395_U110 & new_R395_U107;
  assign new_R395_U71 = new_R395_U116 & new_R395_U115 & new_R395_U111;
  assign new_R395_U72 = new_U3107 & new_R395_U14;
  assign new_R395_U73 = new_R395_U74 & new_R395_U113 & new_R395_U117 & new_R395_U114;
  assign new_R395_U74 = new_R395_U123 & new_R395_U122 & new_R395_U118;
  assign new_R395_U75 = new_U3136 & new_R395_U20;
  assign new_R395_U76 = new_R395_U77 & new_R395_U120 & new_R395_U124 & new_R395_U121;
  assign new_R395_U77 = new_R395_U130 & new_R395_U129 & new_R395_U125;
  assign new_R395_U78 = new_U3101 & new_R395_U26;
  assign new_R395_U79 = new_R395_U127 & new_R395_U80 & new_R395_U128;
  assign new_R395_U80 = new_R395_U132 & new_R395_U131;
  assign new_R395_U81 = new_R395_U134 & new_R395_U135;
  assign new_R395_U82 = new_R395_U137 & new_R395_U138;
  assign new_R395_U83 = new_R395_U140 & new_R395_U141;
  assign new_R395_U84 = new_R395_U143 & new_R395_U144;
  assign new_R395_U85 = new_R395_U146 & new_R395_U147;
  assign new_R395_U86 = new_R395_U149 & new_R395_U150;
  assign new_R395_U87 = new_R395_U152 & new_R395_U153;
  assign new_R395_U88 = new_R395_U155 & new_R395_U156;
  assign new_R395_U89 = new_R395_U158 & new_R395_U159;
  assign new_R395_U90 = new_R395_U161 & new_R395_U162;
  assign new_R395_U91 = new_R395_U164 & new_R395_U165;
  assign new_R395_U92 = new_R395_U167 & new_R395_U168;
  assign new_R395_U93 = new_R395_U170 & new_R395_U171;
  assign new_R395_U94 = new_R395_U173 & new_R395_U174;
  assign new_R395_U95 = new_R395_U176 & new_R395_U177;
  assign new_R395_U96 = new_R395_U179 & new_R395_U180;
  assign new_R395_U97 = new_R395_U182 & new_R395_U186 & new_R395_U185;
  assign new_R395_U98 = ~new_U3082;
  assign new_R395_U99 = new_R395_U188 & new_R395_U187;
  assign new_R395_U100 = ~new_U3144;
  assign new_R395_U101 = ~new_U3145;
  assign new_R395_U102 = ~new_U3113 | ~new_R395_U101 | ~new_R395_U100;
  assign new_R395_U103 = ~new_U3112 | ~new_R395_U100;
  assign new_R395_U104 = ~new_U3111 | ~new_R395_U10;
  assign new_R395_U105 = ~new_R395_U68 | ~new_R395_U67;
  assign new_R395_U106 = ~new_R395_U7 | ~new_R395_U108 | ~new_U3143 | ~new_R395_U109;
  assign new_R395_U107 = ~new_R395_U69 | ~new_R395_U109;
  assign new_R395_U108 = ~new_U3110 | ~new_R395_U11;
  assign new_R395_U109 = ~new_U3109 | ~new_R395_U12;
  assign new_R395_U110 = ~new_U3141 | ~new_R395_U9;
  assign new_R395_U111 = ~new_U3140 | ~new_R395_U16;
  assign new_R395_U112 = ~new_R395_U70 | ~new_R395_U105 | ~new_R395_U71;
  assign new_R395_U113 = ~new_R395_U13 | ~new_R395_U115 | ~new_U3108 | ~new_R395_U116;
  assign new_R395_U114 = ~new_R395_U72 | ~new_R395_U116;
  assign new_R395_U115 = ~new_U3139 | ~new_R395_U17;
  assign new_R395_U116 = ~new_U3138 | ~new_R395_U18;
  assign new_R395_U117 = ~new_U3106 | ~new_R395_U15;
  assign new_R395_U118 = ~new_U3105 | ~new_R395_U22;
  assign new_R395_U119 = ~new_R395_U112 | ~new_R395_U73;
  assign new_R395_U120 = ~new_R395_U19 | ~new_R395_U122 | ~new_U3137 | ~new_R395_U123;
  assign new_R395_U121 = ~new_R395_U75 | ~new_R395_U123;
  assign new_R395_U122 = ~new_U3104 | ~new_R395_U23;
  assign new_R395_U123 = ~new_U3103 | ~new_R395_U24;
  assign new_R395_U124 = ~new_U3135 | ~new_R395_U21;
  assign new_R395_U125 = ~new_U3134 | ~new_R395_U28;
  assign new_R395_U126 = ~new_R395_U119 | ~new_R395_U76;
  assign new_R395_U127 = ~new_R395_U25 | ~new_R395_U129 | ~new_U3102 | ~new_R395_U130;
  assign new_R395_U128 = ~new_R395_U78 | ~new_R395_U130;
  assign new_R395_U129 = ~new_U3133 | ~new_R395_U29;
  assign new_R395_U130 = ~new_U3132 | ~new_R395_U30;
  assign new_R395_U131 = ~new_U3100 | ~new_R395_U27;
  assign new_R395_U132 = ~new_U3099 | ~new_R395_U32;
  assign new_R395_U133 = ~new_R395_U126 | ~new_R395_U79;
  assign new_R395_U134 = ~new_U3131 | ~new_R395_U31;
  assign new_R395_U135 = ~new_U3130 | ~new_R395_U34;
  assign new_R395_U136 = ~new_R395_U81 | ~new_R395_U133;
  assign new_R395_U137 = ~new_U3098 | ~new_R395_U33;
  assign new_R395_U138 = ~new_U3097 | ~new_R395_U36;
  assign new_R395_U139 = ~new_R395_U82 | ~new_R395_U136;
  assign new_R395_U140 = ~new_U3129 | ~new_R395_U35;
  assign new_R395_U141 = ~new_U3128 | ~new_R395_U38;
  assign new_R395_U142 = ~new_R395_U83 | ~new_R395_U139;
  assign new_R395_U143 = ~new_U3096 | ~new_R395_U37;
  assign new_R395_U144 = ~new_U3095 | ~new_R395_U40;
  assign new_R395_U145 = ~new_R395_U84 | ~new_R395_U142;
  assign new_R395_U146 = ~new_U3127 | ~new_R395_U39;
  assign new_R395_U147 = ~new_U3126 | ~new_R395_U42;
  assign new_R395_U148 = ~new_R395_U85 | ~new_R395_U145;
  assign new_R395_U149 = ~new_U3094 | ~new_R395_U41;
  assign new_R395_U150 = ~new_U3093 | ~new_R395_U44;
  assign new_R395_U151 = ~new_R395_U86 | ~new_R395_U148;
  assign new_R395_U152 = ~new_U3125 | ~new_R395_U43;
  assign new_R395_U153 = ~new_U3124 | ~new_R395_U46;
  assign new_R395_U154 = ~new_R395_U87 | ~new_R395_U151;
  assign new_R395_U155 = ~new_U3092 | ~new_R395_U45;
  assign new_R395_U156 = ~new_U3091 | ~new_R395_U48;
  assign new_R395_U157 = ~new_R395_U88 | ~new_R395_U154;
  assign new_R395_U158 = ~new_U3123 | ~new_R395_U47;
  assign new_R395_U159 = ~new_U3122 | ~new_R395_U50;
  assign new_R395_U160 = ~new_R395_U89 | ~new_R395_U157;
  assign new_R395_U161 = ~new_U3090 | ~new_R395_U49;
  assign new_R395_U162 = ~new_U3089 | ~new_R395_U52;
  assign new_R395_U163 = ~new_R395_U90 | ~new_R395_U160;
  assign new_R395_U164 = ~new_U3121 | ~new_R395_U51;
  assign new_R395_U165 = ~new_U3120 | ~new_R395_U54;
  assign new_R395_U166 = ~new_R395_U91 | ~new_R395_U163;
  assign new_R395_U167 = ~new_U3088 | ~new_R395_U53;
  assign new_R395_U168 = ~new_U3087 | ~new_R395_U56;
  assign new_R395_U169 = ~new_R395_U92 | ~new_R395_U166;
  assign new_R395_U170 = ~new_U3119 | ~new_R395_U55;
  assign new_R395_U171 = ~new_U3118 | ~new_R395_U58;
  assign new_R395_U172 = ~new_R395_U93 | ~new_R395_U169;
  assign new_R395_U173 = ~new_U3086 | ~new_R395_U57;
  assign new_R395_U174 = ~new_U3085 | ~new_R395_U60;
  assign new_R395_U175 = ~new_R395_U94 | ~new_R395_U172;
  assign new_R395_U176 = ~new_U3117 | ~new_R395_U59;
  assign new_R395_U177 = ~new_U3116 | ~new_R395_U62;
  assign new_R395_U178 = ~new_R395_U95 | ~new_R395_U175;
  assign new_R395_U179 = ~new_U3084 | ~new_R395_U61;
  assign new_R395_U180 = ~new_U3083 | ~new_R395_U64;
  assign new_R395_U181 = ~new_R395_U96 | ~new_R395_U178;
  assign new_R395_U182 = ~new_U3115 | ~new_R395_U63;
  assign new_R395_U183 = ~new_R395_U97 | ~new_R395_U181;
  assign new_R395_U184 = ~new_R395_U101 | ~new_U3113 | ~new_U3112;
  assign new_R395_U185 = ~new_U3114 | ~new_R395_U98;
  assign new_R395_U186 = ~new_U3082 | ~new_R395_U65;
  assign new_R395_U187 = ~new_R395_U98 | ~new_U3146 | ~new_U3114;
  assign new_R395_U188 = ~new_U3082 | ~new_R395_U66 | ~new_R395_U65;
  assign new_R1105_U4 = new_R1105_U179 & new_R1105_U175;
  assign new_R1105_U5 = ~new_R1105_U83 | ~new_R1105_U180;
  assign new_R1105_U6 = ~REG2_REG_0_;
  assign new_R1105_U7 = ~new_U3453;
  assign new_R1105_U8 = ~REG2_REG_1_;
  assign new_R1105_U9 = ~new_U3453 | ~REG2_REG_0_;
  assign new_R1105_U10 = ~new_U3443;
  assign new_R1105_U11 = ~REG2_REG_2_;
  assign new_R1105_U12 = ~new_U3442;
  assign new_R1105_U13 = ~REG2_REG_3_;
  assign new_R1105_U14 = ~new_U3441;
  assign new_R1105_U15 = ~REG2_REG_4_;
  assign new_R1105_U16 = ~new_U3440;
  assign new_R1105_U17 = ~REG2_REG_5_;
  assign new_R1105_U18 = ~new_U3439;
  assign new_R1105_U19 = ~REG2_REG_6_;
  assign new_R1105_U20 = ~new_U3438;
  assign new_R1105_U21 = ~REG2_REG_7_;
  assign new_R1105_U22 = ~new_U3437;
  assign new_R1105_U23 = ~REG2_REG_8_;
  assign new_R1105_U24 = ~new_U3436;
  assign new_R1105_U25 = ~new_U3435;
  assign new_R1105_U26 = ~REG2_REG_9_;
  assign new_R1105_U27 = ~REG2_REG_10_;
  assign new_R1105_U28 = ~new_U3452;
  assign new_R1105_U29 = ~REG2_REG_11_;
  assign new_R1105_U30 = ~new_U3451;
  assign new_R1105_U31 = ~REG2_REG_12_;
  assign new_R1105_U32 = ~new_U3450;
  assign new_R1105_U33 = ~REG2_REG_13_;
  assign new_R1105_U34 = ~new_U3449;
  assign new_R1105_U35 = ~REG2_REG_14_;
  assign new_R1105_U36 = ~new_U3448;
  assign new_R1105_U37 = ~REG2_REG_15_;
  assign new_R1105_U38 = ~new_U3447;
  assign new_R1105_U39 = ~REG2_REG_16_;
  assign new_R1105_U40 = ~new_U3446;
  assign new_R1105_U41 = ~REG2_REG_17_;
  assign new_R1105_U42 = ~new_U3445;
  assign new_R1105_U43 = ~REG2_REG_18_;
  assign new_R1105_U44 = ~new_U3444;
  assign new_R1105_U45 = ~new_R1105_U170 | ~new_R1105_U169;
  assign new_R1105_U46 = ~new_R1105_U311 | ~new_R1105_U310;
  assign new_R1105_U47 = ~new_R1105_U187 | ~new_R1105_U186;
  assign new_R1105_U48 = ~new_R1105_U194 | ~new_R1105_U193;
  assign new_R1105_U49 = ~new_R1105_U201 | ~new_R1105_U200;
  assign new_R1105_U50 = ~new_R1105_U208 | ~new_R1105_U207;
  assign new_R1105_U51 = ~new_R1105_U215 | ~new_R1105_U214;
  assign new_R1105_U52 = ~new_R1105_U222 | ~new_R1105_U221;
  assign new_R1105_U53 = ~new_R1105_U229 | ~new_R1105_U228;
  assign new_R1105_U54 = ~new_R1105_U236 | ~new_R1105_U235;
  assign new_R1105_U55 = ~new_R1105_U253 | ~new_R1105_U252;
  assign new_R1105_U56 = ~new_R1105_U260 | ~new_R1105_U259;
  assign new_R1105_U57 = ~new_R1105_U267 | ~new_R1105_U266;
  assign new_R1105_U58 = ~new_R1105_U274 | ~new_R1105_U273;
  assign new_R1105_U59 = ~new_R1105_U281 | ~new_R1105_U280;
  assign new_R1105_U60 = ~new_R1105_U288 | ~new_R1105_U287;
  assign new_R1105_U61 = ~new_R1105_U295 | ~new_R1105_U294;
  assign new_R1105_U62 = ~new_R1105_U302 | ~new_R1105_U301;
  assign new_R1105_U63 = ~new_R1105_U309 | ~new_R1105_U308;
  assign new_R1105_U64 = new_R1105_U174 & new_R1105_U243 & new_R1105_U242;
  assign new_R1105_U65 = new_R1105_U178 & new_R1105_U246;
  assign new_R1105_U66 = new_R1105_U182 & new_R1105_U181;
  assign new_R1105_U67 = ~new_R1105_U134 | ~new_R1105_U133;
  assign new_R1105_U68 = new_R1105_U189 & new_R1105_U188;
  assign new_R1105_U69 = ~new_R1105_U130 | ~new_R1105_U129;
  assign new_R1105_U70 = new_R1105_U196 & new_R1105_U195;
  assign new_R1105_U71 = ~new_R1105_U126 | ~new_R1105_U125;
  assign new_R1105_U72 = new_R1105_U203 & new_R1105_U202;
  assign new_R1105_U73 = ~new_R1105_U122 | ~new_R1105_U121;
  assign new_R1105_U74 = new_R1105_U210 & new_R1105_U209;
  assign new_R1105_U75 = ~new_R1105_U118 | ~new_R1105_U117;
  assign new_R1105_U76 = new_R1105_U217 & new_R1105_U216;
  assign new_R1105_U77 = ~new_R1105_U114 | ~new_R1105_U113;
  assign new_R1105_U78 = new_R1105_U224 & new_R1105_U223;
  assign new_R1105_U79 = ~new_R1105_U110 | ~new_R1105_U109;
  assign new_R1105_U80 = new_R1105_U231 & new_R1105_U230;
  assign new_R1105_U81 = ~new_R1105_U82 | ~new_R1105_U106;
  assign new_R1105_U82 = ~new_U3443 | ~new_R1105_U104;
  assign new_R1105_U83 = new_R1105_U241 & new_R1105_U240;
  assign new_R1105_U84 = ~new_U3461;
  assign new_R1105_U85 = ~REG2_REG_19_;
  assign new_R1105_U86 = new_R1105_U248 & new_R1105_U247;
  assign new_R1105_U87 = new_R1105_U255 & new_R1105_U254;
  assign new_R1105_U88 = ~new_R1105_U166 | ~new_R1105_U165;
  assign new_R1105_U89 = new_R1105_U262 & new_R1105_U261;
  assign new_R1105_U90 = ~new_R1105_U162 | ~new_R1105_U161;
  assign new_R1105_U91 = new_R1105_U269 & new_R1105_U268;
  assign new_R1105_U92 = ~new_R1105_U158 | ~new_R1105_U157;
  assign new_R1105_U93 = new_R1105_U276 & new_R1105_U275;
  assign new_R1105_U94 = ~new_R1105_U154 | ~new_R1105_U153;
  assign new_R1105_U95 = new_R1105_U283 & new_R1105_U282;
  assign new_R1105_U96 = ~new_R1105_U150 | ~new_R1105_U149;
  assign new_R1105_U97 = new_R1105_U290 & new_R1105_U289;
  assign new_R1105_U98 = ~new_R1105_U146 | ~new_R1105_U145;
  assign new_R1105_U99 = new_R1105_U297 & new_R1105_U296;
  assign new_R1105_U100 = ~new_R1105_U142 | ~new_R1105_U141;
  assign new_R1105_U101 = new_R1105_U304 & new_R1105_U303;
  assign new_R1105_U102 = ~new_R1105_U138 | ~new_R1105_U137;
  assign new_R1105_U103 = ~new_R1105_U82;
  assign new_R1105_U104 = ~new_R1105_U9;
  assign new_R1105_U105 = ~new_R1105_U10 | ~new_R1105_U9;
  assign new_R1105_U106 = ~REG2_REG_1_ | ~new_R1105_U105;
  assign new_R1105_U107 = ~new_R1105_U81;
  assign new_R1105_U108 = REG2_REG_2_ | new_U3442;
  assign new_R1105_U109 = ~new_R1105_U108 | ~new_R1105_U81;
  assign new_R1105_U110 = ~new_U3442 | ~REG2_REG_2_;
  assign new_R1105_U111 = ~new_R1105_U79;
  assign new_R1105_U112 = REG2_REG_3_ | new_U3441;
  assign new_R1105_U113 = ~new_R1105_U112 | ~new_R1105_U79;
  assign new_R1105_U114 = ~new_U3441 | ~REG2_REG_3_;
  assign new_R1105_U115 = ~new_R1105_U77;
  assign new_R1105_U116 = REG2_REG_4_ | new_U3440;
  assign new_R1105_U117 = ~new_R1105_U116 | ~new_R1105_U77;
  assign new_R1105_U118 = ~new_U3440 | ~REG2_REG_4_;
  assign new_R1105_U119 = ~new_R1105_U75;
  assign new_R1105_U120 = REG2_REG_5_ | new_U3439;
  assign new_R1105_U121 = ~new_R1105_U120 | ~new_R1105_U75;
  assign new_R1105_U122 = ~new_U3439 | ~REG2_REG_5_;
  assign new_R1105_U123 = ~new_R1105_U73;
  assign new_R1105_U124 = REG2_REG_6_ | new_U3438;
  assign new_R1105_U125 = ~new_R1105_U124 | ~new_R1105_U73;
  assign new_R1105_U126 = ~new_U3438 | ~REG2_REG_6_;
  assign new_R1105_U127 = ~new_R1105_U71;
  assign new_R1105_U128 = REG2_REG_7_ | new_U3437;
  assign new_R1105_U129 = ~new_R1105_U128 | ~new_R1105_U71;
  assign new_R1105_U130 = ~new_U3437 | ~REG2_REG_7_;
  assign new_R1105_U131 = ~new_R1105_U69;
  assign new_R1105_U132 = REG2_REG_8_ | new_U3436;
  assign new_R1105_U133 = ~new_R1105_U132 | ~new_R1105_U69;
  assign new_R1105_U134 = ~new_U3436 | ~REG2_REG_8_;
  assign new_R1105_U135 = ~new_R1105_U67;
  assign new_R1105_U136 = REG2_REG_9_ | new_U3435;
  assign new_R1105_U137 = ~new_R1105_U136 | ~new_R1105_U67;
  assign new_R1105_U138 = ~REG2_REG_9_ | ~new_U3435;
  assign new_R1105_U139 = ~new_R1105_U102;
  assign new_R1105_U140 = REG2_REG_10_ | new_U3452;
  assign new_R1105_U141 = ~new_R1105_U140 | ~new_R1105_U102;
  assign new_R1105_U142 = ~new_U3452 | ~REG2_REG_10_;
  assign new_R1105_U143 = ~new_R1105_U100;
  assign new_R1105_U144 = REG2_REG_11_ | new_U3451;
  assign new_R1105_U145 = ~new_R1105_U144 | ~new_R1105_U100;
  assign new_R1105_U146 = ~new_U3451 | ~REG2_REG_11_;
  assign new_R1105_U147 = ~new_R1105_U98;
  assign new_R1105_U148 = REG2_REG_12_ | new_U3450;
  assign new_R1105_U149 = ~new_R1105_U148 | ~new_R1105_U98;
  assign new_R1105_U150 = ~new_U3450 | ~REG2_REG_12_;
  assign new_R1105_U151 = ~new_R1105_U96;
  assign new_R1105_U152 = REG2_REG_13_ | new_U3449;
  assign new_R1105_U153 = ~new_R1105_U152 | ~new_R1105_U96;
  assign new_R1105_U154 = ~new_U3449 | ~REG2_REG_13_;
  assign new_R1105_U155 = ~new_R1105_U94;
  assign new_R1105_U156 = REG2_REG_14_ | new_U3448;
  assign new_R1105_U157 = ~new_R1105_U156 | ~new_R1105_U94;
  assign new_R1105_U158 = ~new_U3448 | ~REG2_REG_14_;
  assign new_R1105_U159 = ~new_R1105_U92;
  assign new_R1105_U160 = REG2_REG_15_ | new_U3447;
  assign new_R1105_U161 = ~new_R1105_U160 | ~new_R1105_U92;
  assign new_R1105_U162 = ~new_U3447 | ~REG2_REG_15_;
  assign new_R1105_U163 = ~new_R1105_U90;
  assign new_R1105_U164 = REG2_REG_16_ | new_U3446;
  assign new_R1105_U165 = ~new_R1105_U164 | ~new_R1105_U90;
  assign new_R1105_U166 = ~new_U3446 | ~REG2_REG_16_;
  assign new_R1105_U167 = ~new_R1105_U88;
  assign new_R1105_U168 = REG2_REG_17_ | new_U3445;
  assign new_R1105_U169 = ~new_R1105_U168 | ~new_R1105_U88;
  assign new_R1105_U170 = ~new_U3445 | ~REG2_REG_17_;
  assign new_R1105_U171 = ~new_R1105_U45;
  assign new_R1105_U172 = REG2_REG_18_ | new_U3444;
  assign new_R1105_U173 = ~new_R1105_U172 | ~new_R1105_U45;
  assign new_R1105_U174 = ~new_U3444 | ~REG2_REG_18_;
  assign new_R1105_U175 = ~new_R1105_U64 | ~new_R1105_U173;
  assign new_R1105_U176 = ~new_U3444 | ~REG2_REG_18_;
  assign new_R1105_U177 = ~new_R1105_U171 | ~new_R1105_U176;
  assign new_R1105_U178 = new_U3444 | REG2_REG_18_;
  assign new_R1105_U179 = ~new_R1105_U65 | ~new_R1105_U177;
  assign new_R1105_U180 = ~new_R1105_U239 | ~new_R1105_U10;
  assign new_R1105_U181 = ~new_U3435 | ~new_R1105_U26;
  assign new_R1105_U182 = ~REG2_REG_9_ | ~new_R1105_U25;
  assign new_R1105_U183 = ~new_U3435 | ~new_R1105_U26;
  assign new_R1105_U184 = ~REG2_REG_9_ | ~new_R1105_U25;
  assign new_R1105_U185 = ~new_R1105_U184 | ~new_R1105_U183;
  assign new_R1105_U186 = ~new_R1105_U66 | ~new_R1105_U67;
  assign new_R1105_U187 = ~new_R1105_U135 | ~new_R1105_U185;
  assign new_R1105_U188 = ~new_U3436 | ~new_R1105_U23;
  assign new_R1105_U189 = ~REG2_REG_8_ | ~new_R1105_U24;
  assign new_R1105_U190 = ~new_U3436 | ~new_R1105_U23;
  assign new_R1105_U191 = ~REG2_REG_8_ | ~new_R1105_U24;
  assign new_R1105_U192 = ~new_R1105_U191 | ~new_R1105_U190;
  assign new_R1105_U193 = ~new_R1105_U68 | ~new_R1105_U69;
  assign new_R1105_U194 = ~new_R1105_U131 | ~new_R1105_U192;
  assign new_R1105_U195 = ~new_U3437 | ~new_R1105_U21;
  assign new_R1105_U196 = ~REG2_REG_7_ | ~new_R1105_U22;
  assign new_R1105_U197 = ~new_U3437 | ~new_R1105_U21;
  assign new_R1105_U198 = ~REG2_REG_7_ | ~new_R1105_U22;
  assign new_R1105_U199 = ~new_R1105_U198 | ~new_R1105_U197;
  assign new_R1105_U200 = ~new_R1105_U70 | ~new_R1105_U71;
  assign new_R1105_U201 = ~new_R1105_U127 | ~new_R1105_U199;
  assign new_R1105_U202 = ~new_U3438 | ~new_R1105_U19;
  assign new_R1105_U203 = ~REG2_REG_6_ | ~new_R1105_U20;
  assign new_R1105_U204 = ~new_U3438 | ~new_R1105_U19;
  assign new_R1105_U205 = ~REG2_REG_6_ | ~new_R1105_U20;
  assign new_R1105_U206 = ~new_R1105_U205 | ~new_R1105_U204;
  assign new_R1105_U207 = ~new_R1105_U72 | ~new_R1105_U73;
  assign new_R1105_U208 = ~new_R1105_U123 | ~new_R1105_U206;
  assign new_R1105_U209 = ~new_U3439 | ~new_R1105_U17;
  assign new_R1105_U210 = ~REG2_REG_5_ | ~new_R1105_U18;
  assign new_R1105_U211 = ~new_U3439 | ~new_R1105_U17;
  assign new_R1105_U212 = ~REG2_REG_5_ | ~new_R1105_U18;
  assign new_R1105_U213 = ~new_R1105_U212 | ~new_R1105_U211;
  assign new_R1105_U214 = ~new_R1105_U74 | ~new_R1105_U75;
  assign new_R1105_U215 = ~new_R1105_U119 | ~new_R1105_U213;
  assign new_R1105_U216 = ~new_U3440 | ~new_R1105_U15;
  assign new_R1105_U217 = ~REG2_REG_4_ | ~new_R1105_U16;
  assign new_R1105_U218 = ~new_U3440 | ~new_R1105_U15;
  assign new_R1105_U219 = ~REG2_REG_4_ | ~new_R1105_U16;
  assign new_R1105_U220 = ~new_R1105_U219 | ~new_R1105_U218;
  assign new_R1105_U221 = ~new_R1105_U76 | ~new_R1105_U77;
  assign new_R1105_U222 = ~new_R1105_U115 | ~new_R1105_U220;
  assign new_R1105_U223 = ~new_U3441 | ~new_R1105_U13;
  assign new_R1105_U224 = ~REG2_REG_3_ | ~new_R1105_U14;
  assign new_R1105_U225 = ~new_U3441 | ~new_R1105_U13;
  assign new_R1105_U226 = ~REG2_REG_3_ | ~new_R1105_U14;
  assign new_R1105_U227 = ~new_R1105_U226 | ~new_R1105_U225;
  assign new_R1105_U228 = ~new_R1105_U78 | ~new_R1105_U79;
  assign new_R1105_U229 = ~new_R1105_U111 | ~new_R1105_U227;
  assign new_R1105_U230 = ~new_U3442 | ~new_R1105_U11;
  assign new_R1105_U231 = ~REG2_REG_2_ | ~new_R1105_U12;
  assign new_R1105_U232 = ~new_U3442 | ~new_R1105_U11;
  assign new_R1105_U233 = ~REG2_REG_2_ | ~new_R1105_U12;
  assign new_R1105_U234 = ~new_R1105_U233 | ~new_R1105_U232;
  assign new_R1105_U235 = ~new_R1105_U80 | ~new_R1105_U81;
  assign new_R1105_U236 = ~new_R1105_U107 | ~new_R1105_U234;
  assign new_R1105_U237 = ~REG2_REG_1_ | ~new_R1105_U9;
  assign new_R1105_U238 = ~new_R1105_U104 | ~new_R1105_U8;
  assign new_R1105_U239 = ~new_R1105_U238 | ~new_R1105_U237;
  assign new_R1105_U240 = ~new_R1105_U8 | ~new_U3443 | ~new_R1105_U9;
  assign new_R1105_U241 = ~new_R1105_U103 | ~REG2_REG_1_;
  assign new_R1105_U242 = ~new_U3461 | ~new_R1105_U85;
  assign new_R1105_U243 = ~REG2_REG_19_ | ~new_R1105_U84;
  assign new_R1105_U244 = ~new_U3461 | ~new_R1105_U85;
  assign new_R1105_U245 = ~REG2_REG_19_ | ~new_R1105_U84;
  assign new_R1105_U246 = ~new_R1105_U245 | ~new_R1105_U244;
  assign new_R1105_U247 = ~new_U3444 | ~new_R1105_U43;
  assign new_R1105_U248 = ~REG2_REG_18_ | ~new_R1105_U44;
  assign new_R1105_U249 = ~new_U3444 | ~new_R1105_U43;
  assign new_R1105_U250 = ~REG2_REG_18_ | ~new_R1105_U44;
  assign new_R1105_U251 = ~new_R1105_U250 | ~new_R1105_U249;
  assign new_R1105_U252 = ~new_R1105_U86 | ~new_R1105_U45;
  assign new_R1105_U253 = ~new_R1105_U251 | ~new_R1105_U171;
  assign new_R1105_U254 = ~new_U3445 | ~new_R1105_U41;
  assign new_R1105_U255 = ~REG2_REG_17_ | ~new_R1105_U42;
  assign new_R1105_U256 = ~new_U3445 | ~new_R1105_U41;
  assign new_R1105_U257 = ~REG2_REG_17_ | ~new_R1105_U42;
  assign new_R1105_U258 = ~new_R1105_U257 | ~new_R1105_U256;
  assign new_R1105_U259 = ~new_R1105_U87 | ~new_R1105_U88;
  assign new_R1105_U260 = ~new_R1105_U167 | ~new_R1105_U258;
  assign new_R1105_U261 = ~new_U3446 | ~new_R1105_U39;
  assign new_R1105_U262 = ~REG2_REG_16_ | ~new_R1105_U40;
  assign new_R1105_U263 = ~new_U3446 | ~new_R1105_U39;
  assign new_R1105_U264 = ~REG2_REG_16_ | ~new_R1105_U40;
  assign new_R1105_U265 = ~new_R1105_U264 | ~new_R1105_U263;
  assign new_R1105_U266 = ~new_R1105_U89 | ~new_R1105_U90;
  assign new_R1105_U267 = ~new_R1105_U163 | ~new_R1105_U265;
  assign new_R1105_U268 = ~new_U3447 | ~new_R1105_U37;
  assign new_R1105_U269 = ~REG2_REG_15_ | ~new_R1105_U38;
  assign new_R1105_U270 = ~new_U3447 | ~new_R1105_U37;
  assign new_R1105_U271 = ~REG2_REG_15_ | ~new_R1105_U38;
  assign new_R1105_U272 = ~new_R1105_U271 | ~new_R1105_U270;
  assign new_R1105_U273 = ~new_R1105_U91 | ~new_R1105_U92;
  assign new_R1105_U274 = ~new_R1105_U159 | ~new_R1105_U272;
  assign new_R1105_U275 = ~new_U3448 | ~new_R1105_U35;
  assign new_R1105_U276 = ~REG2_REG_14_ | ~new_R1105_U36;
  assign new_R1105_U277 = ~new_U3448 | ~new_R1105_U35;
  assign new_R1105_U278 = ~REG2_REG_14_ | ~new_R1105_U36;
  assign new_R1105_U279 = ~new_R1105_U278 | ~new_R1105_U277;
  assign new_R1105_U280 = ~new_R1105_U93 | ~new_R1105_U94;
  assign new_R1105_U281 = ~new_R1105_U155 | ~new_R1105_U279;
  assign new_R1105_U282 = ~new_U3449 | ~new_R1105_U33;
  assign new_R1105_U283 = ~REG2_REG_13_ | ~new_R1105_U34;
  assign new_R1105_U284 = ~new_U3449 | ~new_R1105_U33;
  assign new_R1105_U285 = ~REG2_REG_13_ | ~new_R1105_U34;
  assign new_R1105_U286 = ~new_R1105_U285 | ~new_R1105_U284;
  assign new_R1105_U287 = ~new_R1105_U95 | ~new_R1105_U96;
  assign new_R1105_U288 = ~new_R1105_U151 | ~new_R1105_U286;
  assign new_R1105_U289 = ~new_U3450 | ~new_R1105_U31;
  assign new_R1105_U290 = ~REG2_REG_12_ | ~new_R1105_U32;
  assign new_R1105_U291 = ~new_U3450 | ~new_R1105_U31;
  assign new_R1105_U292 = ~REG2_REG_12_ | ~new_R1105_U32;
  assign new_R1105_U293 = ~new_R1105_U292 | ~new_R1105_U291;
  assign new_R1105_U294 = ~new_R1105_U97 | ~new_R1105_U98;
  assign new_R1105_U295 = ~new_R1105_U147 | ~new_R1105_U293;
  assign new_R1105_U296 = ~new_U3451 | ~new_R1105_U29;
  assign new_R1105_U297 = ~REG2_REG_11_ | ~new_R1105_U30;
  assign new_R1105_U298 = ~new_U3451 | ~new_R1105_U29;
  assign new_R1105_U299 = ~REG2_REG_11_ | ~new_R1105_U30;
  assign new_R1105_U300 = ~new_R1105_U299 | ~new_R1105_U298;
  assign new_R1105_U301 = ~new_R1105_U99 | ~new_R1105_U100;
  assign new_R1105_U302 = ~new_R1105_U143 | ~new_R1105_U300;
  assign new_R1105_U303 = ~new_U3452 | ~new_R1105_U27;
  assign new_R1105_U304 = ~REG2_REG_10_ | ~new_R1105_U28;
  assign new_R1105_U305 = ~new_U3452 | ~new_R1105_U27;
  assign new_R1105_U306 = ~REG2_REG_10_ | ~new_R1105_U28;
  assign new_R1105_U307 = ~new_R1105_U306 | ~new_R1105_U305;
  assign new_R1105_U308 = ~new_R1105_U101 | ~new_R1105_U102;
  assign new_R1105_U309 = ~new_R1105_U139 | ~new_R1105_U307;
  assign new_R1105_U310 = ~new_U3453 | ~new_R1105_U6;
  assign new_R1105_U311 = ~REG2_REG_0_ | ~new_R1105_U7;
  assign new_R1309_U6 = ~new_U3056;
  assign new_R1309_U7 = ~new_U3053;
  assign new_R1309_U8 = new_R1309_U10 & new_R1309_U9;
  assign new_R1309_U9 = ~new_U3053 | ~new_R1309_U6;
  assign new_R1309_U10 = ~new_U3056 | ~new_R1309_U7;
  assign new_R1282_U6 = new_R1282_U130 & new_R1282_U12;
  assign new_R1282_U7 = new_R1282_U106 & new_R1282_U96;
  assign new_R1282_U8 = new_R1282_U105 & new_R1282_U13;
  assign new_R1282_U9 = new_R1282_U104 & new_R1282_U98;
  assign new_R1282_U10 = new_R1282_U103 & new_R1282_U14;
  assign new_R1282_U11 = new_R1282_U102 & new_R1282_U35;
  assign new_R1282_U12 = new_U3470 | new_U3468 | new_U3464;
  assign new_R1282_U13 = ~new_R1282_U95 | ~new_R1282_U19 | ~new_R1282_U20;
  assign new_R1282_U14 = ~new_R1282_U97 | ~new_R1282_U17 | ~new_R1282_U18;
  assign new_R1282_U15 = ~new_R1282_U99 | ~new_R1282_U34 | ~new_R1282_U16;
  assign new_R1282_U16 = ~new_U3480;
  assign new_R1282_U17 = ~new_U3478;
  assign new_R1282_U18 = ~new_U3476;
  assign new_R1282_U19 = ~new_U3474;
  assign new_R1282_U20 = ~new_U3472;
  assign new_R1282_U21 = ~new_R1282_U101 | ~new_R1282_U32 | ~new_R1282_U92;
  assign new_R1282_U22 = ~new_R1282_U108 | ~new_R1282_U87 | ~new_R1282_U90;
  assign new_R1282_U23 = ~new_R1282_U110 | ~new_R1282_U82 | ~new_R1282_U85;
  assign new_R1282_U24 = ~new_R1282_U112 | ~new_R1282_U77 | ~new_R1282_U80;
  assign new_R1282_U25 = ~new_R1282_U114 | ~new_R1282_U72 | ~new_R1282_U75;
  assign new_R1282_U26 = ~new_R1282_U116 | ~new_R1282_U65 | ~new_R1282_U70;
  assign new_R1282_U27 = ~new_R1282_U118 | ~new_R1282_U60 | ~new_R1282_U63;
  assign new_R1282_U28 = ~new_R1282_U120 | ~new_R1282_U55 | ~new_R1282_U58;
  assign new_R1282_U29 = ~new_R1282_U122 | ~new_R1282_U50 | ~new_R1282_U53;
  assign new_R1282_U30 = ~new_R1282_U124 | ~new_R1282_U45 | ~new_R1282_U48;
  assign new_R1282_U31 = ~new_R1282_U160 | ~new_R1282_U159;
  assign new_R1282_U32 = ~new_U3484;
  assign new_R1282_U33 = new_R1282_U132 & new_R1282_U131;
  assign new_R1282_U34 = ~new_U3482;
  assign new_R1282_U35 = ~new_R1282_U99 | ~new_R1282_U16;
  assign new_R1282_U36 = new_R1282_U134 & new_R1282_U133;
  assign new_R1282_U37 = ~new_U4038;
  assign new_R1282_U38 = ~new_R1282_U126 | ~new_R1282_U40 | ~new_R1282_U43;
  assign new_R1282_U39 = new_R1282_U136 & new_R1282_U135;
  assign new_R1282_U40 = ~new_U4039;
  assign new_R1282_U41 = ~new_R1282_U126 | ~new_R1282_U43;
  assign new_R1282_U42 = new_R1282_U138 & new_R1282_U137;
  assign new_R1282_U43 = ~new_U4040;
  assign new_R1282_U44 = new_R1282_U140 & new_R1282_U139;
  assign new_R1282_U45 = ~new_U4029;
  assign new_R1282_U46 = ~new_R1282_U124 | ~new_R1282_U48;
  assign new_R1282_U47 = new_R1282_U142 & new_R1282_U141;
  assign new_R1282_U48 = ~new_U4030;
  assign new_R1282_U49 = new_R1282_U144 & new_R1282_U143;
  assign new_R1282_U50 = ~new_U4031;
  assign new_R1282_U51 = ~new_R1282_U122 | ~new_R1282_U53;
  assign new_R1282_U52 = new_R1282_U146 & new_R1282_U145;
  assign new_R1282_U53 = ~new_U4032;
  assign new_R1282_U54 = new_R1282_U148 & new_R1282_U147;
  assign new_R1282_U55 = ~new_U4033;
  assign new_R1282_U56 = ~new_R1282_U120 | ~new_R1282_U58;
  assign new_R1282_U57 = new_R1282_U150 & new_R1282_U149;
  assign new_R1282_U58 = ~new_U4034;
  assign new_R1282_U59 = new_R1282_U152 & new_R1282_U151;
  assign new_R1282_U60 = ~new_U4035;
  assign new_R1282_U61 = ~new_R1282_U118 | ~new_R1282_U63;
  assign new_R1282_U62 = new_R1282_U154 & new_R1282_U153;
  assign new_R1282_U63 = ~new_U4036;
  assign new_R1282_U64 = new_R1282_U156 & new_R1282_U155;
  assign new_R1282_U65 = ~new_U4037;
  assign new_R1282_U66 = ~new_R1282_U116 | ~new_R1282_U70;
  assign new_R1282_U67 = new_R1282_U158 & new_R1282_U157;
  assign new_R1282_U68 = ~new_U3468;
  assign new_R1282_U69 = ~new_U3464;
  assign new_R1282_U70 = ~new_U3504;
  assign new_R1282_U71 = new_R1282_U162 & new_R1282_U161;
  assign new_R1282_U72 = ~new_U3502;
  assign new_R1282_U73 = ~new_R1282_U114 | ~new_R1282_U75;
  assign new_R1282_U74 = new_R1282_U164 & new_R1282_U163;
  assign new_R1282_U75 = ~new_U3500;
  assign new_R1282_U76 = new_R1282_U166 & new_R1282_U165;
  assign new_R1282_U77 = ~new_U3498;
  assign new_R1282_U78 = ~new_R1282_U112 | ~new_R1282_U80;
  assign new_R1282_U79 = new_R1282_U168 & new_R1282_U167;
  assign new_R1282_U80 = ~new_U3496;
  assign new_R1282_U81 = new_R1282_U170 & new_R1282_U169;
  assign new_R1282_U82 = ~new_U3494;
  assign new_R1282_U83 = ~new_R1282_U110 | ~new_R1282_U85;
  assign new_R1282_U84 = new_R1282_U172 & new_R1282_U171;
  assign new_R1282_U85 = ~new_U3492;
  assign new_R1282_U86 = new_R1282_U174 & new_R1282_U173;
  assign new_R1282_U87 = ~new_U3490;
  assign new_R1282_U88 = ~new_R1282_U108 | ~new_R1282_U90;
  assign new_R1282_U89 = new_R1282_U176 & new_R1282_U175;
  assign new_R1282_U90 = ~new_U3488;
  assign new_R1282_U91 = new_R1282_U178 & new_R1282_U177;
  assign new_R1282_U92 = ~new_U3486;
  assign new_R1282_U93 = ~new_R1282_U101 | ~new_R1282_U32;
  assign new_R1282_U94 = new_R1282_U180 & new_R1282_U179;
  assign new_R1282_U95 = ~new_R1282_U12;
  assign new_R1282_U96 = ~new_R1282_U95 | ~new_R1282_U20;
  assign new_R1282_U97 = ~new_R1282_U13;
  assign new_R1282_U98 = ~new_R1282_U97 | ~new_R1282_U18;
  assign new_R1282_U99 = ~new_R1282_U14;
  assign new_R1282_U100 = ~new_R1282_U35;
  assign new_R1282_U101 = ~new_R1282_U15;
  assign new_R1282_U102 = ~new_U3480 | ~new_R1282_U14;
  assign new_R1282_U103 = ~new_U3478 | ~new_R1282_U98;
  assign new_R1282_U104 = ~new_U3476 | ~new_R1282_U13;
  assign new_R1282_U105 = ~new_U3474 | ~new_R1282_U96;
  assign new_R1282_U106 = ~new_U3472 | ~new_R1282_U12;
  assign new_R1282_U107 = ~new_R1282_U93;
  assign new_R1282_U108 = ~new_R1282_U21;
  assign new_R1282_U109 = ~new_R1282_U88;
  assign new_R1282_U110 = ~new_R1282_U22;
  assign new_R1282_U111 = ~new_R1282_U83;
  assign new_R1282_U112 = ~new_R1282_U23;
  assign new_R1282_U113 = ~new_R1282_U78;
  assign new_R1282_U114 = ~new_R1282_U24;
  assign new_R1282_U115 = ~new_R1282_U73;
  assign new_R1282_U116 = ~new_R1282_U25;
  assign new_R1282_U117 = ~new_R1282_U66;
  assign new_R1282_U118 = ~new_R1282_U26;
  assign new_R1282_U119 = ~new_R1282_U61;
  assign new_R1282_U120 = ~new_R1282_U27;
  assign new_R1282_U121 = ~new_R1282_U56;
  assign new_R1282_U122 = ~new_R1282_U28;
  assign new_R1282_U123 = ~new_R1282_U51;
  assign new_R1282_U124 = ~new_R1282_U29;
  assign new_R1282_U125 = ~new_R1282_U46;
  assign new_R1282_U126 = ~new_R1282_U30;
  assign new_R1282_U127 = ~new_R1282_U41;
  assign new_R1282_U128 = ~new_R1282_U38;
  assign new_R1282_U129 = new_U3468 | new_U3464;
  assign new_R1282_U130 = ~new_U3470 | ~new_R1282_U129;
  assign new_R1282_U131 = ~new_U3484 | ~new_R1282_U15;
  assign new_R1282_U132 = ~new_R1282_U101 | ~new_R1282_U32;
  assign new_R1282_U133 = ~new_U3482 | ~new_R1282_U35;
  assign new_R1282_U134 = ~new_R1282_U100 | ~new_R1282_U34;
  assign new_R1282_U135 = ~new_U4038 | ~new_R1282_U38;
  assign new_R1282_U136 = ~new_R1282_U128 | ~new_R1282_U37;
  assign new_R1282_U137 = ~new_U4039 | ~new_R1282_U41;
  assign new_R1282_U138 = ~new_R1282_U127 | ~new_R1282_U40;
  assign new_R1282_U139 = ~new_U4040 | ~new_R1282_U30;
  assign new_R1282_U140 = ~new_R1282_U126 | ~new_R1282_U43;
  assign new_R1282_U141 = ~new_U4029 | ~new_R1282_U46;
  assign new_R1282_U142 = ~new_R1282_U125 | ~new_R1282_U45;
  assign new_R1282_U143 = ~new_U4030 | ~new_R1282_U29;
  assign new_R1282_U144 = ~new_R1282_U124 | ~new_R1282_U48;
  assign new_R1282_U145 = ~new_U4031 | ~new_R1282_U51;
  assign new_R1282_U146 = ~new_R1282_U123 | ~new_R1282_U50;
  assign new_R1282_U147 = ~new_U4032 | ~new_R1282_U28;
  assign new_R1282_U148 = ~new_R1282_U122 | ~new_R1282_U53;
  assign new_R1282_U149 = ~new_U4033 | ~new_R1282_U56;
  assign new_R1282_U150 = ~new_R1282_U121 | ~new_R1282_U55;
  assign new_R1282_U151 = ~new_U4034 | ~new_R1282_U27;
  assign new_R1282_U152 = ~new_R1282_U120 | ~new_R1282_U58;
  assign new_R1282_U153 = ~new_U4035 | ~new_R1282_U61;
  assign new_R1282_U154 = ~new_R1282_U119 | ~new_R1282_U60;
  assign new_R1282_U155 = ~new_U4036 | ~new_R1282_U26;
  assign new_R1282_U156 = ~new_R1282_U118 | ~new_R1282_U63;
  assign new_R1282_U157 = ~new_U4037 | ~new_R1282_U66;
  assign new_R1282_U158 = ~new_R1282_U117 | ~new_R1282_U65;
  assign new_R1282_U159 = ~new_U3468 | ~new_R1282_U69;
  assign new_R1282_U160 = ~new_U3464 | ~new_R1282_U68;
  assign new_R1282_U161 = ~new_U3504 | ~new_R1282_U25;
  assign new_R1282_U162 = ~new_R1282_U116 | ~new_R1282_U70;
  assign new_R1282_U163 = ~new_U3502 | ~new_R1282_U73;
  assign new_R1282_U164 = ~new_R1282_U115 | ~new_R1282_U72;
  assign new_R1282_U165 = ~new_U3500 | ~new_R1282_U24;
  assign new_R1282_U166 = ~new_R1282_U114 | ~new_R1282_U75;
  assign new_R1282_U167 = ~new_U3498 | ~new_R1282_U78;
  assign new_R1282_U168 = ~new_R1282_U113 | ~new_R1282_U77;
  assign new_R1282_U169 = ~new_U3496 | ~new_R1282_U23;
  assign new_R1282_U170 = ~new_R1282_U112 | ~new_R1282_U80;
  assign new_R1282_U171 = ~new_U3494 | ~new_R1282_U83;
  assign new_R1282_U172 = ~new_R1282_U111 | ~new_R1282_U82;
  assign new_R1282_U173 = ~new_U3492 | ~new_R1282_U22;
  assign new_R1282_U174 = ~new_R1282_U110 | ~new_R1282_U85;
  assign new_R1282_U175 = ~new_U3490 | ~new_R1282_U88;
  assign new_R1282_U176 = ~new_R1282_U109 | ~new_R1282_U87;
  assign new_R1282_U177 = ~new_U3488 | ~new_R1282_U21;
  assign new_R1282_U178 = ~new_R1282_U108 | ~new_R1282_U90;
  assign new_R1282_U179 = ~new_U3486 | ~new_R1282_U93;
  assign new_R1282_U180 = ~new_R1282_U107 | ~new_R1282_U92;
  assign new_R1240_U4 = new_R1240_U196 & new_R1240_U195;
  assign new_R1240_U5 = new_R1240_U197 & new_R1240_U198;
  assign new_R1240_U6 = new_R1240_U210 & new_R1240_U209;
  assign new_R1240_U7 = new_R1240_U250 & new_R1240_U249;
  assign new_R1240_U8 = new_R1240_U258 & new_R1240_U257;
  assign new_R1240_U9 = new_R1240_U274 & new_R1240_U273;
  assign new_R1240_U10 = new_R1240_U282 & new_R1240_U281;
  assign new_R1240_U11 = new_R1240_U10 & new_R1240_U283;
  assign new_R1240_U12 = new_R1240_U7 & new_R1240_U217;
  assign new_R1240_U13 = new_R1240_U8 & new_R1240_U262;
  assign new_R1240_U14 = new_R1240_U11 & new_R1240_U292;
  assign new_R1240_U15 = new_R1240_U13 & new_R1240_U267;
  assign new_R1240_U16 = new_R1240_U9 & new_R1240_U14;
  assign new_R1240_U17 = new_R1240_U299 & new_R1240_U305;
  assign new_R1240_U18 = new_R1240_U359 & new_R1240_U356;
  assign new_R1240_U19 = new_R1240_U352 & new_R1240_U349;
  assign new_R1240_U20 = new_R1240_U343 & new_R1240_U340;
  assign new_R1240_U21 = new_R1240_U334 & new_R1240_U331;
  assign new_R1240_U22 = new_R1240_U328 & new_R1240_U326;
  assign new_R1240_U23 = new_R1240_U321 & new_R1240_U318;
  assign new_R1240_U24 = new_R1240_U248 & new_R1240_U245;
  assign new_R1240_U25 = new_R1240_U240 & new_R1240_U237;
  assign new_R1240_U26 = new_R1240_U226 & new_R1240_U223;
  assign new_R1240_U27 = ~new_U3470;
  assign new_R1240_U28 = ~new_U3065;
  assign new_R1240_U29 = ~new_U3472;
  assign new_R1240_U30 = ~new_U3061;
  assign new_R1240_U31 = ~new_U3474;
  assign new_R1240_U32 = ~new_U3057;
  assign new_R1240_U33 = ~new_U3064;
  assign new_R1240_U34 = ~new_U3057 | ~new_U3474;
  assign new_R1240_U35 = ~new_U3476;
  assign new_R1240_U36 = ~new_U3468 | ~new_U3075;
  assign new_R1240_U37 = ~new_U3464;
  assign new_R1240_U38 = ~new_U3074;
  assign new_R1240_U39 = ~new_R1240_U131 | ~new_R1240_U200;
  assign new_R1240_U40 = ~new_U3478;
  assign new_R1240_U41 = ~new_U3068;
  assign new_R1240_U42 = ~new_U3067;
  assign new_R1240_U43 = ~new_U3068 | ~new_U3478;
  assign new_R1240_U44 = ~new_U3480;
  assign new_R1240_U45 = ~new_R1240_U214 | ~new_R1240_U213;
  assign new_R1240_U46 = ~new_U3482;
  assign new_R1240_U47 = ~new_U3081;
  assign new_R1240_U48 = ~new_U3080;
  assign new_R1240_U49 = ~new_U3484;
  assign new_R1240_U50 = ~new_R1240_U65 | ~new_R1240_U218;
  assign new_R1240_U51 = ~new_R1240_U133 | ~new_R1240_U132;
  assign new_R1240_U52 = ~new_R1240_U136 | ~new_R1240_U232;
  assign new_R1240_U53 = ~new_R1240_U229 | ~new_R1240_U228;
  assign new_R1240_U54 = ~new_U4030;
  assign new_R1240_U55 = ~new_U3050;
  assign new_R1240_U56 = ~new_U3054;
  assign new_R1240_U57 = ~new_U4031;
  assign new_R1240_U58 = ~new_U4033;
  assign new_R1240_U59 = ~new_U3062;
  assign new_R1240_U60 = ~new_U3062 | ~new_U4033;
  assign new_R1240_U61 = ~new_U4035;
  assign new_R1240_U62 = ~new_U3058;
  assign new_R1240_U63 = ~new_U3496;
  assign new_R1240_U64 = ~new_U3071;
  assign new_R1240_U65 = ~new_U3081 | ~new_U3482;
  assign new_R1240_U66 = ~new_U3486;
  assign new_R1240_U67 = ~new_U3059;
  assign new_R1240_U68 = ~new_U3490;
  assign new_R1240_U69 = ~new_U3069;
  assign new_R1240_U70 = ~new_U3488;
  assign new_R1240_U71 = ~new_U3060;
  assign new_R1240_U72 = ~new_U3060 | ~new_U3488;
  assign new_R1240_U73 = ~new_U3492;
  assign new_R1240_U74 = ~new_U3077;
  assign new_R1240_U75 = ~new_U3494;
  assign new_R1240_U76 = ~new_U3076;
  assign new_R1240_U77 = ~new_R1240_U380 | ~new_R1240_U267;
  assign new_R1240_U78 = ~new_U3504;
  assign new_R1240_U79 = ~new_U3078;
  assign new_R1240_U80 = ~new_U3078 | ~new_U3504;
  assign new_R1240_U81 = ~new_U4037;
  assign new_R1240_U82 = ~new_U3502;
  assign new_R1240_U83 = ~new_U3079;
  assign new_R1240_U84 = ~new_U3079 | ~new_U3502;
  assign new_R1240_U85 = ~new_U4036;
  assign new_R1240_U86 = ~new_U3072;
  assign new_R1240_U87 = ~new_U3498;
  assign new_R1240_U88 = ~new_U3070;
  assign new_R1240_U89 = ~new_U3066;
  assign new_R1240_U90 = ~new_U3070 | ~new_U3498;
  assign new_R1240_U91 = ~new_U3500;
  assign new_R1240_U92 = ~new_U4034;
  assign new_R1240_U93 = ~new_U3063;
  assign new_R1240_U94 = ~new_R1240_U146 | ~new_R1240_U388;
  assign new_R1240_U95 = ~new_U4032;
  assign new_R1240_U96 = ~new_U3055;
  assign new_R1240_U97 = ~new_R1240_U397 | ~new_R1240_U396 | ~new_R1240_U306;
  assign new_R1240_U98 = ~new_U3051;
  assign new_R1240_U99 = ~new_U4029;
  assign new_R1240_U100 = ~new_R1240_U60 | ~new_R1240_U314;
  assign new_R1240_U101 = ~new_R1240_U385 | ~new_R1240_U294;
  assign new_R1240_U102 = ~new_R1240_U278 | ~new_R1240_U277;
  assign new_R1240_U103 = ~new_U3073;
  assign new_R1240_U104 = ~new_R1240_U84 | ~new_R1240_U323;
  assign new_R1240_U105 = ~new_R1240_U382 | ~new_R1240_U383 | ~new_R1240_U271;
  assign new_R1240_U106 = ~new_R1240_U72 | ~new_R1240_U345;
  assign new_R1240_U107 = ~new_R1240_U484 | ~new_R1240_U483;
  assign new_R1240_U108 = ~new_R1240_U531 | ~new_R1240_U530;
  assign new_R1240_U109 = ~new_R1240_U402 | ~new_R1240_U401;
  assign new_R1240_U110 = ~new_R1240_U407 | ~new_R1240_U406;
  assign new_R1240_U111 = ~new_R1240_U414 | ~new_R1240_U413;
  assign new_R1240_U112 = ~new_R1240_U421 | ~new_R1240_U420;
  assign new_R1240_U113 = ~new_R1240_U426 | ~new_R1240_U425;
  assign new_R1240_U114 = ~new_R1240_U435 | ~new_R1240_U434;
  assign new_R1240_U115 = ~new_R1240_U442 | ~new_R1240_U441;
  assign new_R1240_U116 = ~new_R1240_U449 | ~new_R1240_U448;
  assign new_R1240_U117 = ~new_R1240_U456 | ~new_R1240_U455;
  assign new_R1240_U118 = ~new_R1240_U461 | ~new_R1240_U460;
  assign new_R1240_U119 = ~new_R1240_U468 | ~new_R1240_U467;
  assign new_R1240_U120 = ~new_R1240_U475 | ~new_R1240_U474;
  assign new_R1240_U121 = ~new_R1240_U489 | ~new_R1240_U488;
  assign new_R1240_U122 = ~new_R1240_U494 | ~new_R1240_U493;
  assign new_R1240_U123 = ~new_R1240_U501 | ~new_R1240_U500;
  assign new_R1240_U124 = ~new_R1240_U508 | ~new_R1240_U507;
  assign new_R1240_U125 = ~new_R1240_U515 | ~new_R1240_U514;
  assign new_R1240_U126 = ~new_R1240_U522 | ~new_R1240_U521;
  assign new_R1240_U127 = ~new_R1240_U527 | ~new_R1240_U526;
  assign new_R1240_U128 = new_R1240_U129 & new_R1240_U197;
  assign new_R1240_U129 = new_U3065 & new_U3470;
  assign new_R1240_U130 = new_U3472 & new_U3061;
  assign new_R1240_U131 = new_U3464 & new_U3074;
  assign new_R1240_U132 = new_R1240_U203 & new_R1240_U204 & new_R1240_U206;
  assign new_R1240_U133 = new_R1240_U374 & new_R1240_U373 & new_R1240_U207;
  assign new_R1240_U134 = new_R1240_U43 & new_R1240_U409 & new_R1240_U408;
  assign new_R1240_U135 = new_R1240_U225 & new_R1240_U6;
  assign new_R1240_U136 = new_R1240_U233 & new_R1240_U231;
  assign new_R1240_U137 = new_R1240_U34 & new_R1240_U416 & new_R1240_U415;
  assign new_R1240_U138 = new_R1240_U239 & new_R1240_U4;
  assign new_R1240_U139 = new_R1240_U247 & new_R1240_U198;
  assign new_R1240_U140 = new_R1240_U252 & new_R1240_U188;
  assign new_R1240_U141 = new_R1240_U6 & new_R1240_U12;
  assign new_R1240_U142 = new_R1240_U378 & new_R1240_U255;
  assign new_R1240_U143 = new_R1240_U270 & new_R1240_U15;
  assign new_R1240_U144 = new_R1240_U260 & new_R1240_U189;
  assign new_R1240_U145 = new_R1240_U296 & new_R1240_U16;
  assign new_R1240_U146 = new_R1240_U389 & new_R1240_U297;
  assign new_R1240_U147 = new_R1240_U309 & new_R1240_U185;
  assign new_R1240_U148 = new_R1240_U395 & new_R1240_U393 & new_R1240_U310;
  assign new_R1240_U149 = new_R1240_U17 & new_R1240_U185;
  assign new_R1240_U150 = new_R1240_U97 & new_R1240_U304;
  assign new_R1240_U151 = new_R1240_U190 & new_R1240_U451 & new_R1240_U450;
  assign new_R1240_U152 = new_R1240_U320 & new_R1240_U185;
  assign new_R1240_U153 = new_R1240_U176 & new_R1240_U288;
  assign new_R1240_U154 = new_R1240_U80 & new_R1240_U482 & new_R1240_U481;
  assign new_R1240_U155 = new_R1240_U333 & new_R1240_U10;
  assign new_R1240_U156 = new_R1240_U90 & new_R1240_U496 & new_R1240_U495;
  assign new_R1240_U157 = new_R1240_U342 & new_R1240_U9;
  assign new_R1240_U158 = new_R1240_U189 & new_R1240_U517 & new_R1240_U516;
  assign new_R1240_U159 = new_R1240_U351 & new_R1240_U8;
  assign new_R1240_U160 = new_R1240_U188 & new_R1240_U529 & new_R1240_U528;
  assign new_R1240_U161 = new_R1240_U358 & new_R1240_U7;
  assign new_R1240_U162 = ~new_R1240_U375 | ~new_R1240_U215;
  assign new_R1240_U163 = ~new_R1240_U230 | ~new_R1240_U242;
  assign new_R1240_U164 = ~new_U3052;
  assign new_R1240_U165 = ~new_U4040;
  assign new_R1240_U166 = new_R1240_U430 & new_R1240_U429;
  assign new_R1240_U167 = ~new_R1240_U372 | ~new_R1240_U312 | ~new_R1240_U186;
  assign new_R1240_U168 = new_R1240_U437 & new_R1240_U436;
  assign new_R1240_U169 = ~new_R1240_U148 | ~new_R1240_U394;
  assign new_R1240_U170 = new_R1240_U444 & new_R1240_U443;
  assign new_R1240_U171 = ~new_R1240_U150 | ~new_R1240_U307;
  assign new_R1240_U172 = ~new_R1240_U301 | ~new_R1240_U300;
  assign new_R1240_U173 = new_R1240_U463 & new_R1240_U462;
  assign new_R1240_U174 = new_R1240_U470 & new_R1240_U469;
  assign new_R1240_U175 = ~new_R1240_U386 | ~new_R1240_U384;
  assign new_R1240_U176 = new_R1240_U477 & new_R1240_U476;
  assign new_R1240_U177 = ~new_U3074 | ~new_U3464;
  assign new_R1240_U178 = ~new_R1240_U36 | ~new_R1240_U335;
  assign new_R1240_U179 = ~new_R1240_U376 | ~new_R1240_U279;
  assign new_R1240_U180 = new_R1240_U503 & new_R1240_U502;
  assign new_R1240_U181 = ~new_R1240_U77 | ~new_R1240_U379;
  assign new_R1240_U182 = new_R1240_U510 & new_R1240_U509;
  assign new_R1240_U183 = ~new_R1240_U265 | ~new_R1240_U264;
  assign new_R1240_U184 = ~new_R1240_U142 | ~new_R1240_U377;
  assign new_R1240_U185 = ~new_R1240_U391 | ~new_R1240_U390;
  assign new_R1240_U186 = ~new_U3051 | ~new_R1240_U169;
  assign new_R1240_U187 = ~new_R1240_U34;
  assign new_R1240_U188 = ~new_U3484 | ~new_U3080;
  assign new_R1240_U189 = ~new_U3069 | ~new_U3490;
  assign new_R1240_U190 = ~new_U3055 | ~new_U4032;
  assign new_R1240_U191 = ~new_R1240_U72;
  assign new_R1240_U192 = ~new_R1240_U84;
  assign new_R1240_U193 = ~new_R1240_U60;
  assign new_R1240_U194 = ~new_R1240_U65;
  assign new_R1240_U195 = new_U3064 | new_U3476;
  assign new_R1240_U196 = new_U3057 | new_U3474;
  assign new_R1240_U197 = new_U3472 | new_U3061;
  assign new_R1240_U198 = new_U3470 | new_U3065;
  assign new_R1240_U199 = ~new_R1240_U177;
  assign new_R1240_U200 = new_U3468 | new_U3075;
  assign new_R1240_U201 = ~new_R1240_U39;
  assign new_R1240_U202 = ~new_R1240_U36;
  assign new_R1240_U203 = ~new_R1240_U4 | ~new_R1240_U128;
  assign new_R1240_U204 = ~new_R1240_U130 | ~new_R1240_U4;
  assign new_R1240_U205 = ~new_R1240_U35 | ~new_R1240_U34;
  assign new_R1240_U206 = ~new_U3064 | ~new_R1240_U205;
  assign new_R1240_U207 = ~new_U3476 | ~new_R1240_U187;
  assign new_R1240_U208 = ~new_R1240_U51;
  assign new_R1240_U209 = new_U3067 | new_U3480;
  assign new_R1240_U210 = new_U3068 | new_U3478;
  assign new_R1240_U211 = ~new_R1240_U43;
  assign new_R1240_U212 = ~new_R1240_U44 | ~new_R1240_U43;
  assign new_R1240_U213 = ~new_U3067 | ~new_R1240_U212;
  assign new_R1240_U214 = ~new_U3480 | ~new_R1240_U211;
  assign new_R1240_U215 = ~new_R1240_U6 | ~new_R1240_U51;
  assign new_R1240_U216 = ~new_R1240_U162;
  assign new_R1240_U217 = new_U3482 | new_U3081;
  assign new_R1240_U218 = ~new_R1240_U217 | ~new_R1240_U162;
  assign new_R1240_U219 = ~new_R1240_U50;
  assign new_R1240_U220 = new_U3080 | new_U3484;
  assign new_R1240_U221 = new_U3478 | new_U3068;
  assign new_R1240_U222 = ~new_R1240_U221 | ~new_R1240_U51;
  assign new_R1240_U223 = ~new_R1240_U134 | ~new_R1240_U222;
  assign new_R1240_U224 = ~new_R1240_U208 | ~new_R1240_U43;
  assign new_R1240_U225 = ~new_U3480 | ~new_U3067;
  assign new_R1240_U226 = ~new_R1240_U135 | ~new_R1240_U224;
  assign new_R1240_U227 = new_U3068 | new_U3478;
  assign new_R1240_U228 = ~new_R1240_U202 | ~new_R1240_U198;
  assign new_R1240_U229 = ~new_U3065 | ~new_U3470;
  assign new_R1240_U230 = ~new_R1240_U53;
  assign new_R1240_U231 = ~new_R1240_U201 | ~new_R1240_U5;
  assign new_R1240_U232 = ~new_R1240_U53 | ~new_R1240_U197;
  assign new_R1240_U233 = ~new_U3061 | ~new_U3472;
  assign new_R1240_U234 = ~new_R1240_U52;
  assign new_R1240_U235 = new_U3474 | new_U3057;
  assign new_R1240_U236 = ~new_R1240_U235 | ~new_R1240_U52;
  assign new_R1240_U237 = ~new_R1240_U137 | ~new_R1240_U236;
  assign new_R1240_U238 = ~new_R1240_U234 | ~new_R1240_U34;
  assign new_R1240_U239 = ~new_U3476 | ~new_U3064;
  assign new_R1240_U240 = ~new_R1240_U138 | ~new_R1240_U238;
  assign new_R1240_U241 = new_U3057 | new_U3474;
  assign new_R1240_U242 = ~new_R1240_U201 | ~new_R1240_U198;
  assign new_R1240_U243 = ~new_R1240_U163;
  assign new_R1240_U244 = ~new_U3061 | ~new_U3472;
  assign new_R1240_U245 = ~new_R1240_U39 | ~new_R1240_U36 | ~new_R1240_U428 | ~new_R1240_U427;
  assign new_R1240_U246 = ~new_R1240_U36 | ~new_R1240_U39;
  assign new_R1240_U247 = ~new_U3065 | ~new_U3470;
  assign new_R1240_U248 = ~new_R1240_U139 | ~new_R1240_U246;
  assign new_R1240_U249 = new_U3080 | new_U3484;
  assign new_R1240_U250 = new_U3059 | new_U3486;
  assign new_R1240_U251 = ~new_R1240_U194 | ~new_R1240_U7;
  assign new_R1240_U252 = ~new_U3059 | ~new_U3486;
  assign new_R1240_U253 = ~new_R1240_U140 | ~new_R1240_U251;
  assign new_R1240_U254 = new_U3486 | new_U3059;
  assign new_R1240_U255 = ~new_R1240_U254 | ~new_R1240_U253;
  assign new_R1240_U256 = ~new_R1240_U184;
  assign new_R1240_U257 = new_U3077 | new_U3492;
  assign new_R1240_U258 = new_U3069 | new_U3490;
  assign new_R1240_U259 = ~new_R1240_U191 | ~new_R1240_U8;
  assign new_R1240_U260 = ~new_U3077 | ~new_U3492;
  assign new_R1240_U261 = ~new_R1240_U144 | ~new_R1240_U259;
  assign new_R1240_U262 = new_U3488 | new_U3060;
  assign new_R1240_U263 = new_U3492 | new_U3077;
  assign new_R1240_U264 = ~new_R1240_U13 | ~new_R1240_U184;
  assign new_R1240_U265 = ~new_R1240_U263 | ~new_R1240_U261;
  assign new_R1240_U266 = ~new_R1240_U183;
  assign new_R1240_U267 = new_U3494 | new_U3076;
  assign new_R1240_U268 = ~new_U3076 | ~new_U3494;
  assign new_R1240_U269 = ~new_R1240_U181;
  assign new_R1240_U270 = new_U3496 | new_U3071;
  assign new_R1240_U271 = ~new_U3071 | ~new_U3496;
  assign new_R1240_U272 = ~new_R1240_U105;
  assign new_R1240_U273 = new_U3066 | new_U3500;
  assign new_R1240_U274 = new_U3070 | new_U3498;
  assign new_R1240_U275 = ~new_R1240_U90;
  assign new_R1240_U276 = ~new_R1240_U91 | ~new_R1240_U90;
  assign new_R1240_U277 = ~new_U3066 | ~new_R1240_U276;
  assign new_R1240_U278 = ~new_U3500 | ~new_R1240_U275;
  assign new_R1240_U279 = ~new_R1240_U9 | ~new_R1240_U105;
  assign new_R1240_U280 = ~new_R1240_U179;
  assign new_R1240_U281 = new_U3073 | new_U4037;
  assign new_R1240_U282 = new_U3078 | new_U3504;
  assign new_R1240_U283 = new_U3072 | new_U4036;
  assign new_R1240_U284 = ~new_R1240_U80;
  assign new_R1240_U285 = ~new_U4037 | ~new_R1240_U284;
  assign new_R1240_U286 = ~new_R1240_U285 | ~new_R1240_U103;
  assign new_R1240_U287 = ~new_R1240_U80 | ~new_R1240_U81;
  assign new_R1240_U288 = ~new_R1240_U287 | ~new_R1240_U286;
  assign new_R1240_U289 = ~new_R1240_U192 | ~new_R1240_U11;
  assign new_R1240_U290 = ~new_U3072 | ~new_U4036;
  assign new_R1240_U291 = ~new_R1240_U290 | ~new_R1240_U289 | ~new_R1240_U288;
  assign new_R1240_U292 = new_U3502 | new_U3079;
  assign new_R1240_U293 = new_U4036 | new_U3072;
  assign new_R1240_U294 = ~new_R1240_U293 | ~new_R1240_U291;
  assign new_R1240_U295 = ~new_R1240_U175;
  assign new_R1240_U296 = new_U4035 | new_U3058;
  assign new_R1240_U297 = ~new_U3058 | ~new_U4035;
  assign new_R1240_U298 = ~new_R1240_U94;
  assign new_R1240_U299 = new_U4034 | new_U3063;
  assign new_R1240_U300 = ~new_R1240_U299 | ~new_R1240_U94;
  assign new_R1240_U301 = ~new_U3063 | ~new_U4034;
  assign new_R1240_U302 = ~new_R1240_U172;
  assign new_R1240_U303 = new_U3055 | new_U4032;
  assign new_R1240_U304 = ~new_R1240_U193 | ~new_R1240_U185;
  assign new_R1240_U305 = new_U4033 | new_U3062;
  assign new_R1240_U306 = new_U4031 | new_U3054;
  assign new_R1240_U307 = ~new_R1240_U149 | ~new_R1240_U392;
  assign new_R1240_U308 = ~new_R1240_U171;
  assign new_R1240_U309 = new_U4030 | new_U3050;
  assign new_R1240_U310 = ~new_U3050 | ~new_U4030;
  assign new_R1240_U311 = ~new_R1240_U169;
  assign new_R1240_U312 = ~new_U4029 | ~new_R1240_U169;
  assign new_R1240_U313 = ~new_R1240_U167;
  assign new_R1240_U314 = ~new_R1240_U305 | ~new_R1240_U172;
  assign new_R1240_U315 = ~new_R1240_U100;
  assign new_R1240_U316 = new_U4032 | new_U3055;
  assign new_R1240_U317 = ~new_R1240_U316 | ~new_R1240_U100;
  assign new_R1240_U318 = ~new_R1240_U151 | ~new_R1240_U317;
  assign new_R1240_U319 = ~new_R1240_U315 | ~new_R1240_U190;
  assign new_R1240_U320 = ~new_U4031 | ~new_U3054;
  assign new_R1240_U321 = ~new_R1240_U152 | ~new_R1240_U319;
  assign new_R1240_U322 = new_U3055 | new_U4032;
  assign new_R1240_U323 = ~new_R1240_U292 | ~new_R1240_U179;
  assign new_R1240_U324 = ~new_R1240_U104;
  assign new_R1240_U325 = ~new_R1240_U10 | ~new_R1240_U104;
  assign new_R1240_U326 = ~new_R1240_U153 | ~new_R1240_U325;
  assign new_R1240_U327 = ~new_R1240_U325 | ~new_R1240_U288;
  assign new_R1240_U328 = ~new_R1240_U480 | ~new_R1240_U327;
  assign new_R1240_U329 = new_U3504 | new_U3078;
  assign new_R1240_U330 = ~new_R1240_U329 | ~new_R1240_U104;
  assign new_R1240_U331 = ~new_R1240_U154 | ~new_R1240_U330;
  assign new_R1240_U332 = ~new_R1240_U324 | ~new_R1240_U80;
  assign new_R1240_U333 = ~new_U3073 | ~new_U4037;
  assign new_R1240_U334 = ~new_R1240_U155 | ~new_R1240_U332;
  assign new_R1240_U335 = new_U3468 | new_U3075;
  assign new_R1240_U336 = ~new_R1240_U178;
  assign new_R1240_U337 = new_U3078 | new_U3504;
  assign new_R1240_U338 = new_U3498 | new_U3070;
  assign new_R1240_U339 = ~new_R1240_U338 | ~new_R1240_U105;
  assign new_R1240_U340 = ~new_R1240_U156 | ~new_R1240_U339;
  assign new_R1240_U341 = ~new_R1240_U272 | ~new_R1240_U90;
  assign new_R1240_U342 = ~new_U3500 | ~new_U3066;
  assign new_R1240_U343 = ~new_R1240_U157 | ~new_R1240_U341;
  assign new_R1240_U344 = new_U3070 | new_U3498;
  assign new_R1240_U345 = ~new_R1240_U262 | ~new_R1240_U184;
  assign new_R1240_U346 = ~new_R1240_U106;
  assign new_R1240_U347 = new_U3490 | new_U3069;
  assign new_R1240_U348 = ~new_R1240_U347 | ~new_R1240_U106;
  assign new_R1240_U349 = ~new_R1240_U158 | ~new_R1240_U348;
  assign new_R1240_U350 = ~new_R1240_U346 | ~new_R1240_U189;
  assign new_R1240_U351 = ~new_U3077 | ~new_U3492;
  assign new_R1240_U352 = ~new_R1240_U159 | ~new_R1240_U350;
  assign new_R1240_U353 = new_U3069 | new_U3490;
  assign new_R1240_U354 = new_U3484 | new_U3080;
  assign new_R1240_U355 = ~new_R1240_U354 | ~new_R1240_U50;
  assign new_R1240_U356 = ~new_R1240_U160 | ~new_R1240_U355;
  assign new_R1240_U357 = ~new_R1240_U219 | ~new_R1240_U188;
  assign new_R1240_U358 = ~new_U3059 | ~new_U3486;
  assign new_R1240_U359 = ~new_R1240_U161 | ~new_R1240_U357;
  assign new_R1240_U360 = ~new_R1240_U220 | ~new_R1240_U188;
  assign new_R1240_U361 = ~new_R1240_U217 | ~new_R1240_U65;
  assign new_R1240_U362 = ~new_R1240_U227 | ~new_R1240_U43;
  assign new_R1240_U363 = ~new_R1240_U241 | ~new_R1240_U34;
  assign new_R1240_U364 = ~new_R1240_U244 | ~new_R1240_U197;
  assign new_R1240_U365 = ~new_R1240_U322 | ~new_R1240_U190;
  assign new_R1240_U366 = ~new_R1240_U305 | ~new_R1240_U60;
  assign new_R1240_U367 = ~new_R1240_U337 | ~new_R1240_U80;
  assign new_R1240_U368 = ~new_R1240_U292 | ~new_R1240_U84;
  assign new_R1240_U369 = ~new_R1240_U344 | ~new_R1240_U90;
  assign new_R1240_U370 = ~new_R1240_U353 | ~new_R1240_U189;
  assign new_R1240_U371 = ~new_R1240_U262 | ~new_R1240_U72;
  assign new_R1240_U372 = ~new_U4029 | ~new_U3051;
  assign new_R1240_U373 = ~new_R1240_U5 | ~new_R1240_U202 | ~new_R1240_U4;
  assign new_R1240_U374 = ~new_R1240_U201 | ~new_R1240_U5 | ~new_R1240_U4;
  assign new_R1240_U375 = ~new_R1240_U45;
  assign new_R1240_U376 = ~new_R1240_U102;
  assign new_R1240_U377 = ~new_R1240_U141 | ~new_R1240_U51;
  assign new_R1240_U378 = ~new_R1240_U12 | ~new_R1240_U45;
  assign new_R1240_U379 = ~new_R1240_U15 | ~new_R1240_U184;
  assign new_R1240_U380 = ~new_R1240_U268 | ~new_R1240_U265;
  assign new_R1240_U381 = ~new_R1240_U77;
  assign new_R1240_U382 = ~new_R1240_U143 | ~new_R1240_U184;
  assign new_R1240_U383 = ~new_R1240_U381 | ~new_R1240_U270;
  assign new_R1240_U384 = ~new_R1240_U16 | ~new_R1240_U105;
  assign new_R1240_U385 = ~new_R1240_U14 | ~new_R1240_U102;
  assign new_R1240_U386 = ~new_R1240_U101;
  assign new_R1240_U387 = ~new_R1240_U97;
  assign new_R1240_U388 = ~new_R1240_U145 | ~new_R1240_U105;
  assign new_R1240_U389 = ~new_R1240_U101 | ~new_R1240_U296;
  assign new_R1240_U390 = ~new_U3054 | ~new_R1240_U303;
  assign new_R1240_U391 = ~new_U4031 | ~new_R1240_U303;
  assign new_R1240_U392 = ~new_R1240_U298 | ~new_R1240_U301;
  assign new_R1240_U393 = ~new_R1240_U309 | ~new_R1240_U193 | ~new_R1240_U185;
  assign new_R1240_U394 = ~new_R1240_U147 | ~new_R1240_U17 | ~new_R1240_U392;
  assign new_R1240_U395 = ~new_R1240_U387 | ~new_R1240_U309;
  assign new_R1240_U396 = ~new_R1240_U57 | ~new_R1240_U190;
  assign new_R1240_U397 = ~new_R1240_U56 | ~new_R1240_U190;
  assign new_R1240_U398 = ~new_U3080 | ~new_R1240_U49;
  assign new_R1240_U399 = ~new_U3484 | ~new_R1240_U48;
  assign new_R1240_U400 = ~new_R1240_U399 | ~new_R1240_U398;
  assign new_R1240_U401 = ~new_R1240_U360 | ~new_R1240_U50;
  assign new_R1240_U402 = ~new_R1240_U400 | ~new_R1240_U219;
  assign new_R1240_U403 = ~new_U3081 | ~new_R1240_U46;
  assign new_R1240_U404 = ~new_U3482 | ~new_R1240_U47;
  assign new_R1240_U405 = ~new_R1240_U404 | ~new_R1240_U403;
  assign new_R1240_U406 = ~new_R1240_U361 | ~new_R1240_U162;
  assign new_R1240_U407 = ~new_R1240_U216 | ~new_R1240_U405;
  assign new_R1240_U408 = ~new_U3067 | ~new_R1240_U44;
  assign new_R1240_U409 = ~new_U3480 | ~new_R1240_U42;
  assign new_R1240_U410 = ~new_U3068 | ~new_R1240_U40;
  assign new_R1240_U411 = ~new_U3478 | ~new_R1240_U41;
  assign new_R1240_U412 = ~new_R1240_U411 | ~new_R1240_U410;
  assign new_R1240_U413 = ~new_R1240_U362 | ~new_R1240_U51;
  assign new_R1240_U414 = ~new_R1240_U412 | ~new_R1240_U208;
  assign new_R1240_U415 = ~new_U3064 | ~new_R1240_U35;
  assign new_R1240_U416 = ~new_U3476 | ~new_R1240_U33;
  assign new_R1240_U417 = ~new_U3057 | ~new_R1240_U31;
  assign new_R1240_U418 = ~new_U3474 | ~new_R1240_U32;
  assign new_R1240_U419 = ~new_R1240_U418 | ~new_R1240_U417;
  assign new_R1240_U420 = ~new_R1240_U363 | ~new_R1240_U52;
  assign new_R1240_U421 = ~new_R1240_U419 | ~new_R1240_U234;
  assign new_R1240_U422 = ~new_U3061 | ~new_R1240_U29;
  assign new_R1240_U423 = ~new_U3472 | ~new_R1240_U30;
  assign new_R1240_U424 = ~new_R1240_U423 | ~new_R1240_U422;
  assign new_R1240_U425 = ~new_R1240_U364 | ~new_R1240_U163;
  assign new_R1240_U426 = ~new_R1240_U243 | ~new_R1240_U424;
  assign new_R1240_U427 = ~new_U3065 | ~new_R1240_U27;
  assign new_R1240_U428 = ~new_U3470 | ~new_R1240_U28;
  assign new_R1240_U429 = ~new_U3052 | ~new_R1240_U165;
  assign new_R1240_U430 = ~new_U4040 | ~new_R1240_U164;
  assign new_R1240_U431 = ~new_U3052 | ~new_R1240_U165;
  assign new_R1240_U432 = ~new_U4040 | ~new_R1240_U164;
  assign new_R1240_U433 = ~new_R1240_U432 | ~new_R1240_U431;
  assign new_R1240_U434 = ~new_R1240_U166 | ~new_R1240_U167;
  assign new_R1240_U435 = ~new_R1240_U313 | ~new_R1240_U433;
  assign new_R1240_U436 = ~new_U3051 | ~new_R1240_U99;
  assign new_R1240_U437 = ~new_U4029 | ~new_R1240_U98;
  assign new_R1240_U438 = ~new_U3051 | ~new_R1240_U99;
  assign new_R1240_U439 = ~new_U4029 | ~new_R1240_U98;
  assign new_R1240_U440 = ~new_R1240_U439 | ~new_R1240_U438;
  assign new_R1240_U441 = ~new_R1240_U168 | ~new_R1240_U169;
  assign new_R1240_U442 = ~new_R1240_U311 | ~new_R1240_U440;
  assign new_R1240_U443 = ~new_U3050 | ~new_R1240_U54;
  assign new_R1240_U444 = ~new_U4030 | ~new_R1240_U55;
  assign new_R1240_U445 = ~new_U3050 | ~new_R1240_U54;
  assign new_R1240_U446 = ~new_U4030 | ~new_R1240_U55;
  assign new_R1240_U447 = ~new_R1240_U446 | ~new_R1240_U445;
  assign new_R1240_U448 = ~new_R1240_U170 | ~new_R1240_U171;
  assign new_R1240_U449 = ~new_R1240_U308 | ~new_R1240_U447;
  assign new_R1240_U450 = ~new_U3054 | ~new_R1240_U57;
  assign new_R1240_U451 = ~new_U4031 | ~new_R1240_U56;
  assign new_R1240_U452 = ~new_U3055 | ~new_R1240_U95;
  assign new_R1240_U453 = ~new_U4032 | ~new_R1240_U96;
  assign new_R1240_U454 = ~new_R1240_U453 | ~new_R1240_U452;
  assign new_R1240_U455 = ~new_R1240_U365 | ~new_R1240_U100;
  assign new_R1240_U456 = ~new_R1240_U454 | ~new_R1240_U315;
  assign new_R1240_U457 = ~new_U3062 | ~new_R1240_U58;
  assign new_R1240_U458 = ~new_U4033 | ~new_R1240_U59;
  assign new_R1240_U459 = ~new_R1240_U458 | ~new_R1240_U457;
  assign new_R1240_U460 = ~new_R1240_U366 | ~new_R1240_U172;
  assign new_R1240_U461 = ~new_R1240_U302 | ~new_R1240_U459;
  assign new_R1240_U462 = ~new_U3063 | ~new_R1240_U92;
  assign new_R1240_U463 = ~new_U4034 | ~new_R1240_U93;
  assign new_R1240_U464 = ~new_U3063 | ~new_R1240_U92;
  assign new_R1240_U465 = ~new_U4034 | ~new_R1240_U93;
  assign new_R1240_U466 = ~new_R1240_U465 | ~new_R1240_U464;
  assign new_R1240_U467 = ~new_R1240_U173 | ~new_R1240_U94;
  assign new_R1240_U468 = ~new_R1240_U466 | ~new_R1240_U298;
  assign new_R1240_U469 = ~new_U3058 | ~new_R1240_U61;
  assign new_R1240_U470 = ~new_U4035 | ~new_R1240_U62;
  assign new_R1240_U471 = ~new_U3058 | ~new_R1240_U61;
  assign new_R1240_U472 = ~new_U4035 | ~new_R1240_U62;
  assign new_R1240_U473 = ~new_R1240_U472 | ~new_R1240_U471;
  assign new_R1240_U474 = ~new_R1240_U174 | ~new_R1240_U175;
  assign new_R1240_U475 = ~new_R1240_U295 | ~new_R1240_U473;
  assign new_R1240_U476 = ~new_U3072 | ~new_R1240_U85;
  assign new_R1240_U477 = ~new_U4036 | ~new_R1240_U86;
  assign new_R1240_U478 = ~new_U3072 | ~new_R1240_U85;
  assign new_R1240_U479 = ~new_U4036 | ~new_R1240_U86;
  assign new_R1240_U480 = ~new_R1240_U479 | ~new_R1240_U478;
  assign new_R1240_U481 = ~new_U3073 | ~new_R1240_U81;
  assign new_R1240_U482 = ~new_U4037 | ~new_R1240_U103;
  assign new_R1240_U483 = ~new_R1240_U199 | ~new_R1240_U178;
  assign new_R1240_U484 = ~new_R1240_U336 | ~new_R1240_U177;
  assign new_R1240_U485 = ~new_U3078 | ~new_R1240_U78;
  assign new_R1240_U486 = ~new_U3504 | ~new_R1240_U79;
  assign new_R1240_U487 = ~new_R1240_U486 | ~new_R1240_U485;
  assign new_R1240_U488 = ~new_R1240_U367 | ~new_R1240_U104;
  assign new_R1240_U489 = ~new_R1240_U487 | ~new_R1240_U324;
  assign new_R1240_U490 = ~new_U3079 | ~new_R1240_U82;
  assign new_R1240_U491 = ~new_U3502 | ~new_R1240_U83;
  assign new_R1240_U492 = ~new_R1240_U491 | ~new_R1240_U490;
  assign new_R1240_U493 = ~new_R1240_U368 | ~new_R1240_U179;
  assign new_R1240_U494 = ~new_R1240_U280 | ~new_R1240_U492;
  assign new_R1240_U495 = ~new_U3066 | ~new_R1240_U91;
  assign new_R1240_U496 = ~new_U3500 | ~new_R1240_U89;
  assign new_R1240_U497 = ~new_U3070 | ~new_R1240_U87;
  assign new_R1240_U498 = ~new_U3498 | ~new_R1240_U88;
  assign new_R1240_U499 = ~new_R1240_U498 | ~new_R1240_U497;
  assign new_R1240_U500 = ~new_R1240_U369 | ~new_R1240_U105;
  assign new_R1240_U501 = ~new_R1240_U499 | ~new_R1240_U272;
  assign new_R1240_U502 = ~new_U3071 | ~new_R1240_U63;
  assign new_R1240_U503 = ~new_U3496 | ~new_R1240_U64;
  assign new_R1240_U504 = ~new_U3071 | ~new_R1240_U63;
  assign new_R1240_U505 = ~new_U3496 | ~new_R1240_U64;
  assign new_R1240_U506 = ~new_R1240_U505 | ~new_R1240_U504;
  assign new_R1240_U507 = ~new_R1240_U180 | ~new_R1240_U181;
  assign new_R1240_U508 = ~new_R1240_U269 | ~new_R1240_U506;
  assign new_R1240_U509 = ~new_U3076 | ~new_R1240_U75;
  assign new_R1240_U510 = ~new_U3494 | ~new_R1240_U76;
  assign new_R1240_U511 = ~new_U3076 | ~new_R1240_U75;
  assign new_R1240_U512 = ~new_U3494 | ~new_R1240_U76;
  assign new_R1240_U513 = ~new_R1240_U512 | ~new_R1240_U511;
  assign new_R1240_U514 = ~new_R1240_U182 | ~new_R1240_U183;
  assign new_R1240_U515 = ~new_R1240_U266 | ~new_R1240_U513;
  assign new_R1240_U516 = ~new_U3077 | ~new_R1240_U73;
  assign new_R1240_U517 = ~new_U3492 | ~new_R1240_U74;
  assign new_R1240_U518 = ~new_U3069 | ~new_R1240_U68;
  assign new_R1240_U519 = ~new_U3490 | ~new_R1240_U69;
  assign new_R1240_U520 = ~new_R1240_U519 | ~new_R1240_U518;
  assign new_R1240_U521 = ~new_R1240_U370 | ~new_R1240_U106;
  assign new_R1240_U522 = ~new_R1240_U520 | ~new_R1240_U346;
  assign new_R1240_U523 = ~new_U3060 | ~new_R1240_U70;
  assign new_R1240_U524 = ~new_U3488 | ~new_R1240_U71;
  assign new_R1240_U525 = ~new_R1240_U524 | ~new_R1240_U523;
  assign new_R1240_U526 = ~new_R1240_U371 | ~new_R1240_U184;
  assign new_R1240_U527 = ~new_R1240_U256 | ~new_R1240_U525;
  assign new_R1240_U528 = ~new_U3059 | ~new_R1240_U66;
  assign new_R1240_U529 = ~new_U3486 | ~new_R1240_U67;
  assign new_R1240_U530 = ~new_U3074 | ~new_R1240_U37;
  assign new_R1240_U531 = ~new_U3464 | ~new_R1240_U38;
  assign new_R1162_U4 = new_R1162_U165 & new_R1162_U161;
  assign new_R1162_U5 = ~new_R1162_U84 | ~new_R1162_U166;
  assign new_R1162_U6 = ~REG1_REG_0_;
  assign new_R1162_U7 = ~new_U3453;
  assign new_R1162_U8 = ~new_U3443;
  assign new_R1162_U9 = ~new_U3453 | ~REG1_REG_0_;
  assign new_R1162_U10 = ~REG1_REG_1_;
  assign new_R1162_U11 = ~REG1_REG_2_;
  assign new_R1162_U12 = ~new_U3442;
  assign new_R1162_U13 = ~new_R1162_U103 | ~new_R1162_U102;
  assign new_R1162_U14 = ~new_U3441;
  assign new_R1162_U15 = ~REG1_REG_3_;
  assign new_R1162_U16 = ~REG1_REG_4_;
  assign new_R1162_U17 = ~new_U3440;
  assign new_R1162_U18 = ~new_R1162_U110 | ~new_R1162_U109;
  assign new_R1162_U19 = ~new_U3439;
  assign new_R1162_U20 = ~REG1_REG_5_;
  assign new_R1162_U21 = ~REG1_REG_6_;
  assign new_R1162_U22 = ~new_U3438;
  assign new_R1162_U23 = ~REG1_REG_7_;
  assign new_R1162_U24 = ~new_U3437;
  assign new_R1162_U25 = ~new_R1162_U121 | ~new_R1162_U120;
  assign new_R1162_U26 = ~new_U3436;
  assign new_R1162_U27 = ~REG1_REG_8_;
  assign new_R1162_U28 = ~new_U3435;
  assign new_R1162_U29 = ~REG1_REG_9_;
  assign new_R1162_U30 = ~new_R1162_U128 | ~new_R1162_U127;
  assign new_R1162_U31 = ~new_U3452;
  assign new_R1162_U32 = ~REG1_REG_10_;
  assign new_R1162_U33 = ~REG1_REG_11_;
  assign new_R1162_U34 = ~new_U3451;
  assign new_R1162_U35 = ~REG1_REG_12_;
  assign new_R1162_U36 = ~new_U3450;
  assign new_R1162_U37 = ~new_R1162_U139 | ~new_R1162_U138;
  assign new_R1162_U38 = ~new_U3449;
  assign new_R1162_U39 = ~REG1_REG_13_;
  assign new_R1162_U40 = ~new_R1162_U142 | ~new_R1162_U141;
  assign new_R1162_U41 = ~new_U3448;
  assign new_R1162_U42 = ~REG1_REG_14_;
  assign new_R1162_U43 = ~new_R1162_U145 | ~new_R1162_U144;
  assign new_R1162_U44 = ~new_U3447;
  assign new_R1162_U45 = ~REG1_REG_15_;
  assign new_R1162_U46 = ~REG1_REG_16_;
  assign new_R1162_U47 = ~new_U3446;
  assign new_R1162_U48 = ~REG1_REG_17_;
  assign new_R1162_U49 = ~new_U3445;
  assign new_R1162_U50 = ~REG1_REG_18_;
  assign new_R1162_U51 = ~new_U3444;
  assign new_R1162_U52 = ~new_R1162_U156 | ~new_R1162_U155;
  assign new_R1162_U53 = ~new_R1162_U290 | ~new_R1162_U289;
  assign new_R1162_U54 = ~new_R1162_U173 | ~new_R1162_U172;
  assign new_R1162_U55 = ~new_R1162_U179 | ~new_R1162_U178;
  assign new_R1162_U56 = ~new_R1162_U186 | ~new_R1162_U185;
  assign new_R1162_U57 = ~new_R1162_U193 | ~new_R1162_U192;
  assign new_R1162_U58 = ~new_R1162_U199 | ~new_R1162_U198;
  assign new_R1162_U59 = ~new_R1162_U206 | ~new_R1162_U205;
  assign new_R1162_U60 = ~new_R1162_U212 | ~new_R1162_U211;
  assign new_R1162_U61 = ~new_R1162_U219 | ~new_R1162_U218;
  assign new_R1162_U62 = ~new_R1162_U236 | ~new_R1162_U235;
  assign new_R1162_U63 = ~new_R1162_U243 | ~new_R1162_U242;
  assign new_R1162_U64 = ~new_R1162_U250 | ~new_R1162_U249;
  assign new_R1162_U65 = ~new_R1162_U256 | ~new_R1162_U255;
  assign new_R1162_U66 = ~new_R1162_U262 | ~new_R1162_U261;
  assign new_R1162_U67 = ~new_R1162_U268 | ~new_R1162_U267;
  assign new_R1162_U68 = ~new_R1162_U275 | ~new_R1162_U274;
  assign new_R1162_U69 = ~new_R1162_U282 | ~new_R1162_U281;
  assign new_R1162_U70 = ~new_R1162_U288 | ~new_R1162_U287;
  assign new_R1162_U71 = new_R1162_U160 & new_R1162_U226 & new_R1162_U225;
  assign new_R1162_U72 = new_R1162_U164 & new_R1162_U229;
  assign new_R1162_U73 = new_R1162_U168 & new_R1162_U167;
  assign new_R1162_U74 = ~new_R1162_U124 | ~new_R1162_U123;
  assign new_R1162_U75 = new_R1162_U181 & new_R1162_U180;
  assign new_R1162_U76 = ~new_R1162_U117 | ~new_R1162_U116;
  assign new_R1162_U77 = new_R1162_U188 & new_R1162_U187;
  assign new_R1162_U78 = ~new_R1162_U113 | ~new_R1162_U112;
  assign new_R1162_U79 = new_R1162_U201 & new_R1162_U200;
  assign new_R1162_U80 = ~new_R1162_U106 | ~new_R1162_U105;
  assign new_R1162_U81 = new_R1162_U214 & new_R1162_U213;
  assign new_R1162_U82 = ~new_R1162_U83 | ~new_R1162_U99;
  assign new_R1162_U83 = ~REG1_REG_1_ | ~new_R1162_U97;
  assign new_R1162_U84 = new_R1162_U224 & new_R1162_U223;
  assign new_R1162_U85 = ~new_U3461;
  assign new_R1162_U86 = ~REG1_REG_19_;
  assign new_R1162_U87 = new_R1162_U231 & new_R1162_U230;
  assign new_R1162_U88 = new_R1162_U238 & new_R1162_U237;
  assign new_R1162_U89 = ~new_R1162_U152 | ~new_R1162_U151;
  assign new_R1162_U90 = new_R1162_U245 & new_R1162_U244;
  assign new_R1162_U91 = ~new_R1162_U148 | ~new_R1162_U147;
  assign new_R1162_U92 = new_R1162_U270 & new_R1162_U269;
  assign new_R1162_U93 = ~new_R1162_U135 | ~new_R1162_U134;
  assign new_R1162_U94 = new_R1162_U277 & new_R1162_U276;
  assign new_R1162_U95 = ~new_R1162_U131 | ~new_R1162_U130;
  assign new_R1162_U96 = ~new_R1162_U83;
  assign new_R1162_U97 = ~new_R1162_U9;
  assign new_R1162_U98 = ~new_R1162_U10 | ~new_R1162_U9;
  assign new_R1162_U99 = ~new_U3443 | ~new_R1162_U98;
  assign new_R1162_U100 = ~new_R1162_U82;
  assign new_R1162_U101 = REG1_REG_2_ | new_U3442;
  assign new_R1162_U102 = ~new_R1162_U101 | ~new_R1162_U82;
  assign new_R1162_U103 = ~new_U3442 | ~REG1_REG_2_;
  assign new_R1162_U104 = ~new_R1162_U13;
  assign new_R1162_U105 = ~new_U3441 | ~new_R1162_U208;
  assign new_R1162_U106 = ~REG1_REG_3_ | ~new_R1162_U13;
  assign new_R1162_U107 = ~new_R1162_U80;
  assign new_R1162_U108 = REG1_REG_4_ | new_U3440;
  assign new_R1162_U109 = ~new_R1162_U108 | ~new_R1162_U80;
  assign new_R1162_U110 = ~new_U3440 | ~REG1_REG_4_;
  assign new_R1162_U111 = ~new_R1162_U18;
  assign new_R1162_U112 = ~new_U3439 | ~new_R1162_U195;
  assign new_R1162_U113 = ~REG1_REG_5_ | ~new_R1162_U18;
  assign new_R1162_U114 = ~new_R1162_U78;
  assign new_R1162_U115 = REG1_REG_6_ | new_U3438;
  assign new_R1162_U116 = ~new_R1162_U115 | ~new_R1162_U78;
  assign new_R1162_U117 = ~new_U3438 | ~REG1_REG_6_;
  assign new_R1162_U118 = ~new_R1162_U76;
  assign new_R1162_U119 = REG1_REG_7_ | new_U3437;
  assign new_R1162_U120 = ~new_R1162_U119 | ~new_R1162_U76;
  assign new_R1162_U121 = ~new_U3437 | ~REG1_REG_7_;
  assign new_R1162_U122 = ~new_R1162_U25;
  assign new_R1162_U123 = ~new_U3436 | ~new_R1162_U175;
  assign new_R1162_U124 = ~REG1_REG_8_ | ~new_R1162_U25;
  assign new_R1162_U125 = ~new_R1162_U74;
  assign new_R1162_U126 = REG1_REG_9_ | new_U3435;
  assign new_R1162_U127 = ~new_R1162_U126 | ~new_R1162_U74;
  assign new_R1162_U128 = ~REG1_REG_9_ | ~new_U3435;
  assign new_R1162_U129 = ~new_R1162_U30;
  assign new_R1162_U130 = ~new_U3452 | ~new_R1162_U284;
  assign new_R1162_U131 = ~REG1_REG_10_ | ~new_R1162_U30;
  assign new_R1162_U132 = ~new_R1162_U95;
  assign new_R1162_U133 = REG1_REG_11_ | new_U3451;
  assign new_R1162_U134 = ~new_R1162_U133 | ~new_R1162_U95;
  assign new_R1162_U135 = ~new_U3451 | ~REG1_REG_11_;
  assign new_R1162_U136 = ~new_R1162_U93;
  assign new_R1162_U137 = REG1_REG_12_ | new_U3450;
  assign new_R1162_U138 = ~new_R1162_U137 | ~new_R1162_U93;
  assign new_R1162_U139 = ~new_U3450 | ~REG1_REG_12_;
  assign new_R1162_U140 = ~new_R1162_U37;
  assign new_R1162_U141 = ~new_U3449 | ~new_R1162_U264;
  assign new_R1162_U142 = ~REG1_REG_13_ | ~new_R1162_U37;
  assign new_R1162_U143 = ~new_R1162_U40;
  assign new_R1162_U144 = ~new_U3448 | ~new_R1162_U258;
  assign new_R1162_U145 = ~REG1_REG_14_ | ~new_R1162_U40;
  assign new_R1162_U146 = ~new_R1162_U43;
  assign new_R1162_U147 = ~new_U3447 | ~new_R1162_U252;
  assign new_R1162_U148 = ~REG1_REG_15_ | ~new_R1162_U43;
  assign new_R1162_U149 = ~new_R1162_U91;
  assign new_R1162_U150 = REG1_REG_16_ | new_U3446;
  assign new_R1162_U151 = ~new_R1162_U150 | ~new_R1162_U91;
  assign new_R1162_U152 = ~new_U3446 | ~REG1_REG_16_;
  assign new_R1162_U153 = ~new_R1162_U89;
  assign new_R1162_U154 = REG1_REG_17_ | new_U3445;
  assign new_R1162_U155 = ~new_R1162_U154 | ~new_R1162_U89;
  assign new_R1162_U156 = ~new_U3445 | ~REG1_REG_17_;
  assign new_R1162_U157 = ~new_R1162_U52;
  assign new_R1162_U158 = REG1_REG_18_ | new_U3444;
  assign new_R1162_U159 = ~new_R1162_U158 | ~new_R1162_U52;
  assign new_R1162_U160 = ~new_U3444 | ~REG1_REG_18_;
  assign new_R1162_U161 = ~new_R1162_U71 | ~new_R1162_U159;
  assign new_R1162_U162 = ~new_U3444 | ~REG1_REG_18_;
  assign new_R1162_U163 = ~new_R1162_U157 | ~new_R1162_U162;
  assign new_R1162_U164 = new_U3444 | REG1_REG_18_;
  assign new_R1162_U165 = ~new_R1162_U72 | ~new_R1162_U163;
  assign new_R1162_U166 = ~new_R1162_U222 | ~new_R1162_U10;
  assign new_R1162_U167 = ~new_U3435 | ~new_R1162_U29;
  assign new_R1162_U168 = ~REG1_REG_9_ | ~new_R1162_U28;
  assign new_R1162_U169 = ~new_U3435 | ~new_R1162_U29;
  assign new_R1162_U170 = ~REG1_REG_9_ | ~new_R1162_U28;
  assign new_R1162_U171 = ~new_R1162_U170 | ~new_R1162_U169;
  assign new_R1162_U172 = ~new_R1162_U73 | ~new_R1162_U74;
  assign new_R1162_U173 = ~new_R1162_U125 | ~new_R1162_U171;
  assign new_R1162_U174 = ~REG1_REG_8_ | ~new_R1162_U25;
  assign new_R1162_U175 = ~new_R1162_U122 | ~new_R1162_U27;
  assign new_R1162_U176 = ~REG1_REG_8_ | ~new_R1162_U25;
  assign new_R1162_U177 = ~new_R1162_U175 | ~new_R1162_U176;
  assign new_R1162_U178 = ~new_R1162_U26 | ~new_R1162_U175 | ~new_R1162_U174;
  assign new_R1162_U179 = ~new_R1162_U177 | ~new_U3436;
  assign new_R1162_U180 = ~new_U3437 | ~new_R1162_U23;
  assign new_R1162_U181 = ~REG1_REG_7_ | ~new_R1162_U24;
  assign new_R1162_U182 = ~new_U3437 | ~new_R1162_U23;
  assign new_R1162_U183 = ~REG1_REG_7_ | ~new_R1162_U24;
  assign new_R1162_U184 = ~new_R1162_U183 | ~new_R1162_U182;
  assign new_R1162_U185 = ~new_R1162_U75 | ~new_R1162_U76;
  assign new_R1162_U186 = ~new_R1162_U118 | ~new_R1162_U184;
  assign new_R1162_U187 = ~new_U3438 | ~new_R1162_U21;
  assign new_R1162_U188 = ~REG1_REG_6_ | ~new_R1162_U22;
  assign new_R1162_U189 = ~new_U3438 | ~new_R1162_U21;
  assign new_R1162_U190 = ~REG1_REG_6_ | ~new_R1162_U22;
  assign new_R1162_U191 = ~new_R1162_U190 | ~new_R1162_U189;
  assign new_R1162_U192 = ~new_R1162_U77 | ~new_R1162_U78;
  assign new_R1162_U193 = ~new_R1162_U114 | ~new_R1162_U191;
  assign new_R1162_U194 = ~REG1_REG_5_ | ~new_R1162_U18;
  assign new_R1162_U195 = ~new_R1162_U111 | ~new_R1162_U20;
  assign new_R1162_U196 = ~REG1_REG_5_ | ~new_R1162_U18;
  assign new_R1162_U197 = ~new_R1162_U195 | ~new_R1162_U196;
  assign new_R1162_U198 = ~new_R1162_U19 | ~new_R1162_U195 | ~new_R1162_U194;
  assign new_R1162_U199 = ~new_R1162_U197 | ~new_U3439;
  assign new_R1162_U200 = ~new_U3440 | ~new_R1162_U16;
  assign new_R1162_U201 = ~REG1_REG_4_ | ~new_R1162_U17;
  assign new_R1162_U202 = ~new_U3440 | ~new_R1162_U16;
  assign new_R1162_U203 = ~REG1_REG_4_ | ~new_R1162_U17;
  assign new_R1162_U204 = ~new_R1162_U203 | ~new_R1162_U202;
  assign new_R1162_U205 = ~new_R1162_U79 | ~new_R1162_U80;
  assign new_R1162_U206 = ~new_R1162_U107 | ~new_R1162_U204;
  assign new_R1162_U207 = ~REG1_REG_3_ | ~new_R1162_U13;
  assign new_R1162_U208 = ~new_R1162_U104 | ~new_R1162_U15;
  assign new_R1162_U209 = ~REG1_REG_3_ | ~new_R1162_U13;
  assign new_R1162_U210 = ~new_R1162_U208 | ~new_R1162_U209;
  assign new_R1162_U211 = ~new_R1162_U14 | ~new_R1162_U208 | ~new_R1162_U207;
  assign new_R1162_U212 = ~new_R1162_U210 | ~new_U3441;
  assign new_R1162_U213 = ~new_U3442 | ~new_R1162_U11;
  assign new_R1162_U214 = ~REG1_REG_2_ | ~new_R1162_U12;
  assign new_R1162_U215 = ~new_U3442 | ~new_R1162_U11;
  assign new_R1162_U216 = ~REG1_REG_2_ | ~new_R1162_U12;
  assign new_R1162_U217 = ~new_R1162_U216 | ~new_R1162_U215;
  assign new_R1162_U218 = ~new_R1162_U81 | ~new_R1162_U82;
  assign new_R1162_U219 = ~new_R1162_U100 | ~new_R1162_U217;
  assign new_R1162_U220 = ~new_U3443 | ~new_R1162_U9;
  assign new_R1162_U221 = ~new_R1162_U97 | ~new_R1162_U8;
  assign new_R1162_U222 = ~new_R1162_U221 | ~new_R1162_U220;
  assign new_R1162_U223 = ~new_R1162_U8 | ~REG1_REG_1_ | ~new_R1162_U9;
  assign new_R1162_U224 = ~new_R1162_U96 | ~new_U3443;
  assign new_R1162_U225 = ~new_U3461 | ~new_R1162_U86;
  assign new_R1162_U226 = ~REG1_REG_19_ | ~new_R1162_U85;
  assign new_R1162_U227 = ~new_U3461 | ~new_R1162_U86;
  assign new_R1162_U228 = ~REG1_REG_19_ | ~new_R1162_U85;
  assign new_R1162_U229 = ~new_R1162_U228 | ~new_R1162_U227;
  assign new_R1162_U230 = ~new_U3444 | ~new_R1162_U50;
  assign new_R1162_U231 = ~REG1_REG_18_ | ~new_R1162_U51;
  assign new_R1162_U232 = ~new_U3444 | ~new_R1162_U50;
  assign new_R1162_U233 = ~REG1_REG_18_ | ~new_R1162_U51;
  assign new_R1162_U234 = ~new_R1162_U233 | ~new_R1162_U232;
  assign new_R1162_U235 = ~new_R1162_U87 | ~new_R1162_U52;
  assign new_R1162_U236 = ~new_R1162_U234 | ~new_R1162_U157;
  assign new_R1162_U237 = ~new_U3445 | ~new_R1162_U48;
  assign new_R1162_U238 = ~REG1_REG_17_ | ~new_R1162_U49;
  assign new_R1162_U239 = ~new_U3445 | ~new_R1162_U48;
  assign new_R1162_U240 = ~REG1_REG_17_ | ~new_R1162_U49;
  assign new_R1162_U241 = ~new_R1162_U240 | ~new_R1162_U239;
  assign new_R1162_U242 = ~new_R1162_U88 | ~new_R1162_U89;
  assign new_R1162_U243 = ~new_R1162_U153 | ~new_R1162_U241;
  assign new_R1162_U244 = ~new_U3446 | ~new_R1162_U46;
  assign new_R1162_U245 = ~REG1_REG_16_ | ~new_R1162_U47;
  assign new_R1162_U246 = ~new_U3446 | ~new_R1162_U46;
  assign new_R1162_U247 = ~REG1_REG_16_ | ~new_R1162_U47;
  assign new_R1162_U248 = ~new_R1162_U247 | ~new_R1162_U246;
  assign new_R1162_U249 = ~new_R1162_U90 | ~new_R1162_U91;
  assign new_R1162_U250 = ~new_R1162_U149 | ~new_R1162_U248;
  assign new_R1162_U251 = ~REG1_REG_15_ | ~new_R1162_U43;
  assign new_R1162_U252 = ~new_R1162_U146 | ~new_R1162_U45;
  assign new_R1162_U253 = ~REG1_REG_15_ | ~new_R1162_U43;
  assign new_R1162_U254 = ~new_R1162_U252 | ~new_R1162_U253;
  assign new_R1162_U255 = ~new_R1162_U44 | ~new_R1162_U252 | ~new_R1162_U251;
  assign new_R1162_U256 = ~new_R1162_U254 | ~new_U3447;
  assign new_R1162_U257 = ~REG1_REG_14_ | ~new_R1162_U40;
  assign new_R1162_U258 = ~new_R1162_U143 | ~new_R1162_U42;
  assign new_R1162_U259 = ~REG1_REG_14_ | ~new_R1162_U40;
  assign new_R1162_U260 = ~new_R1162_U258 | ~new_R1162_U259;
  assign new_R1162_U261 = ~new_R1162_U41 | ~new_R1162_U258 | ~new_R1162_U257;
  assign new_R1162_U262 = ~new_R1162_U260 | ~new_U3448;
  assign new_R1162_U263 = ~REG1_REG_13_ | ~new_R1162_U37;
  assign new_R1162_U264 = ~new_R1162_U140 | ~new_R1162_U39;
  assign new_R1162_U265 = ~REG1_REG_13_ | ~new_R1162_U37;
  assign new_R1162_U266 = ~new_R1162_U264 | ~new_R1162_U265;
  assign new_R1162_U267 = ~new_R1162_U38 | ~new_R1162_U264 | ~new_R1162_U263;
  assign new_R1162_U268 = ~new_R1162_U266 | ~new_U3449;
  assign new_R1162_U269 = ~new_U3450 | ~new_R1162_U35;
  assign new_R1162_U270 = ~REG1_REG_12_ | ~new_R1162_U36;
  assign new_R1162_U271 = ~new_U3450 | ~new_R1162_U35;
  assign new_R1162_U272 = ~REG1_REG_12_ | ~new_R1162_U36;
  assign new_R1162_U273 = ~new_R1162_U272 | ~new_R1162_U271;
  assign new_R1162_U274 = ~new_R1162_U92 | ~new_R1162_U93;
  assign new_R1162_U275 = ~new_R1162_U136 | ~new_R1162_U273;
  assign new_R1162_U276 = ~new_U3451 | ~new_R1162_U33;
  assign new_R1162_U277 = ~REG1_REG_11_ | ~new_R1162_U34;
  assign new_R1162_U278 = ~new_U3451 | ~new_R1162_U33;
  assign new_R1162_U279 = ~REG1_REG_11_ | ~new_R1162_U34;
  assign new_R1162_U280 = ~new_R1162_U279 | ~new_R1162_U278;
  assign new_R1162_U281 = ~new_R1162_U94 | ~new_R1162_U95;
  assign new_R1162_U282 = ~new_R1162_U132 | ~new_R1162_U280;
  assign new_R1162_U283 = ~REG1_REG_10_ | ~new_R1162_U30;
  assign new_R1162_U284 = ~new_R1162_U129 | ~new_R1162_U32;
  assign new_R1162_U285 = ~REG1_REG_10_ | ~new_R1162_U30;
  assign new_R1162_U286 = ~new_R1162_U284 | ~new_R1162_U285;
  assign new_R1162_U287 = ~new_R1162_U31 | ~new_R1162_U284 | ~new_R1162_U283;
  assign new_R1162_U288 = ~new_R1162_U286 | ~new_U3452;
  assign new_R1162_U289 = ~new_U3453 | ~new_R1162_U6;
  assign new_R1162_U290 = ~REG1_REG_0_ | ~new_R1162_U7;
  assign new_R1117_U6 = new_R1117_U228 & new_R1117_U227;
  assign new_R1117_U7 = new_R1117_U208 & new_R1117_U261;
  assign new_R1117_U8 = new_R1117_U263 & new_R1117_U262;
  assign new_R1117_U9 = new_R1117_U209 & new_R1117_U272;
  assign new_R1117_U10 = new_R1117_U274 & new_R1117_U273;
  assign new_R1117_U11 = new_R1117_U186 & new_R1117_U290;
  assign new_R1117_U12 = new_R1117_U292 & new_R1117_U291;
  assign new_R1117_U13 = new_R1117_U304 & new_R1117_U211;
  assign new_R1117_U14 = new_R1117_U231 & new_R1117_U226 & new_R1117_U213;
  assign new_R1117_U15 = new_R1117_U236 & new_R1117_U214;
  assign new_R1117_U16 = new_R1117_U7 & new_R1117_U241;
  assign new_R1117_U17 = new_R1117_U9 & new_R1117_U277;
  assign new_R1117_U18 = new_R1117_U11 & new_R1117_U295;
  assign new_R1117_U19 = new_R1117_U16 & new_R1117_U268;
  assign new_R1117_U20 = new_R1117_U288 & new_R1117_U286;
  assign new_R1117_U21 = new_R1117_U20 & new_R1117_U18;
  assign new_R1117_U22 = new_R1117_U421 & new_R1117_U420;
  assign new_R1117_U23 = ~new_R1117_U328 | ~new_R1117_U331;
  assign new_R1117_U24 = ~new_R1117_U319 | ~new_R1117_U322;
  assign new_R1117_U25 = ~new_R1117_U453 | ~new_R1117_U454 | ~new_R1117_U383 | ~new_R1117_U382;
  assign new_R1117_U26 = ~new_R1117_U150 | ~new_R1117_U203;
  assign new_R1117_U27 = ~new_R1117_U259 | ~new_R1117_U371;
  assign new_R1117_U28 = ~new_R1117_U252 | ~new_R1117_U255;
  assign new_R1117_U29 = ~new_R1117_U244 | ~new_R1117_U246;
  assign new_R1117_U30 = ~new_R1117_U192 | ~new_R1117_U334;
  assign new_R1117_U31 = new_R1117_U373 & new_R1117_U379;
  assign new_R1117_U32 = ~new_U3067;
  assign new_R1117_U33 = ~new_U3067 | ~new_R1117_U38;
  assign new_R1117_U34 = ~new_U3081;
  assign new_R1117_U35 = ~new_U3476;
  assign new_R1117_U36 = ~new_U3478;
  assign new_R1117_U37 = ~new_U3474;
  assign new_R1117_U38 = ~new_U3480;
  assign new_R1117_U39 = ~new_U3482;
  assign new_R1117_U40 = ~new_U3065;
  assign new_R1117_U41 = ~new_U3065 | ~new_R1117_U43;
  assign new_R1117_U42 = ~new_U3061;
  assign new_R1117_U43 = ~new_U3470;
  assign new_R1117_U44 = ~new_U3464;
  assign new_R1117_U45 = ~new_U3075;
  assign new_R1117_U46 = ~new_U3472;
  assign new_R1117_U47 = ~new_U3068;
  assign new_R1117_U48 = ~new_U3064;
  assign new_R1117_U49 = ~new_U3057;
  assign new_R1117_U50 = ~new_U3057 | ~new_R1117_U37;
  assign new_R1117_U51 = ~new_R1117_U232 | ~new_R1117_U230;
  assign new_R1117_U52 = ~new_U3484;
  assign new_R1117_U53 = ~new_U3080;
  assign new_R1117_U54 = ~new_R1117_U51 | ~new_R1117_U233;
  assign new_R1117_U55 = ~new_R1117_U50 | ~new_R1117_U248;
  assign new_R1117_U56 = ~new_R1117_U335 | ~new_R1117_U220 | ~new_R1117_U204;
  assign new_R1117_U57 = ~new_U4029;
  assign new_R1117_U58 = ~new_U3054;
  assign new_R1117_U59 = ~new_U3054 | ~new_R1117_U99;
  assign new_R1117_U60 = ~new_U3050;
  assign new_R1117_U61 = ~new_U3062;
  assign new_R1117_U62 = ~new_U4033;
  assign new_R1117_U63 = ~new_U3063;
  assign new_R1117_U64 = ~new_U3058;
  assign new_R1117_U65 = ~new_U3072;
  assign new_R1117_U66 = ~new_U4034;
  assign new_R1117_U67 = ~new_U4035;
  assign new_R1117_U68 = ~new_U3072 | ~new_R1117_U69;
  assign new_R1117_U69 = ~new_U4036;
  assign new_R1117_U70 = ~new_U3073;
  assign new_R1117_U71 = ~new_U3078;
  assign new_R1117_U72 = ~new_U4037;
  assign new_R1117_U73 = ~new_U3078 | ~new_R1117_U74;
  assign new_R1117_U74 = ~new_U3504;
  assign new_R1117_U75 = ~new_U3079;
  assign new_R1117_U76 = ~new_U3066;
  assign new_R1117_U77 = ~new_U3500;
  assign new_R1117_U78 = ~new_U3498;
  assign new_R1117_U79 = ~new_U3496;
  assign new_R1117_U80 = ~new_U3494;
  assign new_R1117_U81 = ~new_U3077;
  assign new_R1117_U82 = ~new_U3492;
  assign new_R1117_U83 = ~new_U3490;
  assign new_R1117_U84 = ~new_U3060;
  assign new_R1117_U85 = ~new_U3059;
  assign new_R1117_U86 = ~new_U3488;
  assign new_R1117_U87 = ~new_U3486;
  assign new_R1117_U88 = ~new_U3080 | ~new_R1117_U52;
  assign new_R1117_U89 = ~new_U3069;
  assign new_R1117_U90 = ~new_R1117_U339 | ~new_R1117_U268;
  assign new_R1117_U91 = ~new_U3070;
  assign new_R1117_U92 = ~new_U3071;
  assign new_R1117_U93 = ~new_U3076;
  assign new_R1117_U94 = ~new_U3076 | ~new_R1117_U80;
  assign new_R1117_U95 = ~new_R1117_U278 | ~new_R1117_U276;
  assign new_R1117_U96 = ~new_U3502;
  assign new_R1117_U97 = ~new_U4032;
  assign new_R1117_U98 = ~new_U3055;
  assign new_R1117_U99 = ~new_U4031;
  assign new_R1117_U100 = ~new_U4030;
  assign new_R1117_U101 = ~new_U3051;
  assign new_R1117_U102 = ~new_R1117_U431 | ~new_R1117_U211;
  assign new_R1117_U103 = ~new_R1117_U346 | ~new_R1117_U297;
  assign new_R1117_U104 = ~new_R1117_U157 | ~new_R1117_U356;
  assign new_R1117_U105 = ~new_R1117_U344 | ~new_R1117_U289;
  assign new_R1117_U106 = ~new_R1117_U94 | ~new_R1117_U315;
  assign new_R1117_U107 = ~new_R1117_U360 | ~new_R1117_U88;
  assign new_R1117_U108 = ~new_U3074;
  assign new_R1117_U109 = ~new_R1117_U428 | ~new_R1117_U427;
  assign new_R1117_U110 = ~new_R1117_U444 | ~new_R1117_U443;
  assign new_R1117_U111 = ~new_R1117_U449 | ~new_R1117_U448;
  assign new_R1117_U112 = ~new_R1117_U467 | ~new_R1117_U466;
  assign new_R1117_U113 = ~new_R1117_U472 | ~new_R1117_U471;
  assign new_R1117_U114 = ~new_R1117_U477 | ~new_R1117_U476;
  assign new_R1117_U115 = ~new_R1117_U482 | ~new_R1117_U481;
  assign new_R1117_U116 = ~new_R1117_U487 | ~new_R1117_U486;
  assign new_R1117_U117 = ~new_R1117_U503 | ~new_R1117_U502;
  assign new_R1117_U118 = ~new_R1117_U508 | ~new_R1117_U507;
  assign new_R1117_U119 = ~new_R1117_U387 | ~new_R1117_U386;
  assign new_R1117_U120 = ~new_R1117_U396 | ~new_R1117_U395;
  assign new_R1117_U121 = ~new_R1117_U403 | ~new_R1117_U402;
  assign new_R1117_U122 = ~new_R1117_U407 | ~new_R1117_U406;
  assign new_R1117_U123 = ~new_R1117_U416 | ~new_R1117_U415;
  assign new_R1117_U124 = ~new_R1117_U439 | ~new_R1117_U438;
  assign new_R1117_U125 = ~new_R1117_U458 | ~new_R1117_U457;
  assign new_R1117_U126 = ~new_R1117_U462 | ~new_R1117_U461;
  assign new_R1117_U127 = ~new_R1117_U494 | ~new_R1117_U493;
  assign new_R1117_U128 = ~new_R1117_U498 | ~new_R1117_U497;
  assign new_R1117_U129 = ~new_R1117_U515 | ~new_R1117_U514;
  assign new_R1117_U130 = new_R1117_U222 & new_R1117_U212;
  assign new_R1117_U131 = new_R1117_U225 & new_R1117_U224;
  assign new_R1117_U132 = new_R1117_U15 & new_R1117_U14;
  assign new_R1117_U133 = new_R1117_U239 & new_R1117_U238;
  assign new_R1117_U134 = new_R1117_U338 & new_R1117_U133;
  assign new_R1117_U135 = new_R1117_U33 & new_R1117_U389 & new_R1117_U388;
  assign new_R1117_U136 = new_R1117_U392 & new_R1117_U214;
  assign new_R1117_U137 = new_R1117_U254 & new_R1117_U6;
  assign new_R1117_U138 = new_R1117_U399 & new_R1117_U213;
  assign new_R1117_U139 = new_R1117_U41 & new_R1117_U409 & new_R1117_U408;
  assign new_R1117_U140 = new_R1117_U412 & new_R1117_U212;
  assign new_R1117_U141 = new_R1117_U270 & new_R1117_U19;
  assign new_R1117_U142 = new_R1117_U17 & new_R1117_U282;
  assign new_R1117_U143 = new_R1117_U343 & new_R1117_U283;
  assign new_R1117_U144 = new_R1117_U21 & new_R1117_U298;
  assign new_R1117_U145 = new_R1117_U348 & new_R1117_U299;
  assign new_R1117_U146 = new_R1117_U307 & new_R1117_U306;
  assign new_R1117_U147 = new_R1117_U419 & new_R1117_U308;
  assign new_R1117_U148 = new_R1117_U307 & new_R1117_U22;
  assign new_R1117_U149 = new_R1117_U309 & new_R1117_U148 & new_R1117_U306;
  assign new_R1117_U150 = new_R1117_U375 & new_R1117_U179;
  assign new_R1117_U151 = ~new_R1117_U425 | ~new_R1117_U424;
  assign new_R1117_U152 = new_R1117_U211 & new_R1117_U102;
  assign new_R1117_U153 = ~new_R1117_U441 | ~new_R1117_U440;
  assign new_R1117_U154 = ~new_R1117_U446 | ~new_R1117_U445;
  assign new_R1117_U155 = new_U3058 & new_R1117_U67;
  assign new_R1117_U156 = new_R1117_U20 & new_R1117_U295;
  assign new_R1117_U157 = new_R1117_U349 & new_R1117_U68;
  assign new_R1117_U158 = new_R1117_U12 & new_R1117_U311;
  assign new_R1117_U159 = ~new_R1117_U464 | ~new_R1117_U463;
  assign new_R1117_U160 = ~new_R1117_U469 | ~new_R1117_U468;
  assign new_R1117_U161 = ~new_R1117_U474 | ~new_R1117_U473;
  assign new_R1117_U162 = ~new_R1117_U479 | ~new_R1117_U478;
  assign new_R1117_U163 = ~new_R1117_U484 | ~new_R1117_U483;
  assign new_R1117_U164 = new_R1117_U321 & new_R1117_U10;
  assign new_R1117_U165 = new_R1117_U490 & new_R1117_U209;
  assign new_R1117_U166 = ~new_R1117_U500 | ~new_R1117_U499;
  assign new_R1117_U167 = ~new_R1117_U505 | ~new_R1117_U504;
  assign new_R1117_U168 = new_R1117_U330 & new_R1117_U8;
  assign new_R1117_U169 = new_R1117_U511 & new_R1117_U208;
  assign new_R1117_U170 = new_R1117_U385 & new_R1117_U384;
  assign new_R1117_U171 = ~new_R1117_U134 | ~new_R1117_U337;
  assign new_R1117_U172 = new_R1117_U394 & new_R1117_U393;
  assign new_R1117_U173 = new_R1117_U401 & new_R1117_U400;
  assign new_R1117_U174 = new_R1117_U405 & new_R1117_U404;
  assign new_R1117_U175 = ~new_R1117_U131 | ~new_R1117_U368;
  assign new_R1117_U176 = new_R1117_U414 & new_R1117_U413;
  assign new_R1117_U177 = ~new_U4040;
  assign new_R1117_U178 = ~new_U3052;
  assign new_R1117_U179 = new_R1117_U423 & new_R1117_U422;
  assign new_R1117_U180 = ~new_R1117_U146 | ~new_R1117_U376;
  assign new_R1117_U181 = new_R1117_U435 & new_R1117_U434;
  assign new_R1117_U182 = new_R1117_U437 & new_R1117_U436;
  assign new_R1117_U183 = ~new_R1117_U302 | ~new_R1117_U301;
  assign new_R1117_U184 = ~new_R1117_U145 | ~new_R1117_U358;
  assign new_R1117_U185 = ~new_R1117_U347 | ~new_R1117_U354;
  assign new_R1117_U186 = ~new_U4035 | ~new_R1117_U64;
  assign new_R1117_U187 = new_R1117_U456 & new_R1117_U455;
  assign new_R1117_U188 = new_R1117_U460 & new_R1117_U459;
  assign new_R1117_U189 = ~new_R1117_U345 | ~new_R1117_U352;
  assign new_R1117_U190 = ~new_R1117_U350 | ~new_R1117_U73;
  assign new_R1117_U191 = ~new_U3468;
  assign new_R1117_U192 = ~new_U3464 | ~new_R1117_U108;
  assign new_R1117_U193 = ~new_R1117_U380 | ~new_R1117_U336;
  assign new_R1117_U194 = ~new_R1117_U143 | ~new_R1117_U342;
  assign new_R1117_U195 = ~new_R1117_U95 | ~new_R1117_U279;
  assign new_R1117_U196 = new_R1117_U492 & new_R1117_U491;
  assign new_R1117_U197 = new_R1117_U496 & new_R1117_U495;
  assign new_R1117_U198 = ~new_R1117_U366 | ~new_R1117_U341 | ~new_R1117_U271;
  assign new_R1117_U199 = ~new_R1117_U364 | ~new_R1117_U90;
  assign new_R1117_U200 = ~new_R1117_U362 | ~new_R1117_U267;
  assign new_R1117_U201 = new_R1117_U513 & new_R1117_U512;
  assign new_R1117_U202 = ~new_R1117_U102;
  assign new_R1117_U203 = ~new_R1117_U147 | ~new_R1117_U180;
  assign new_R1117_U204 = ~new_R1117_U192 | ~new_R1117_U191;
  assign new_R1117_U205 = ~new_R1117_U59;
  assign new_R1117_U206 = ~new_R1117_U41;
  assign new_R1117_U207 = ~new_R1117_U33;
  assign new_R1117_U208 = ~new_U3486 | ~new_R1117_U85;
  assign new_R1117_U209 = ~new_U3496 | ~new_R1117_U92;
  assign new_R1117_U210 = ~new_R1117_U186;
  assign new_R1117_U211 = ~new_U4031 | ~new_R1117_U58;
  assign new_R1117_U212 = ~new_U3470 | ~new_R1117_U40;
  assign new_R1117_U213 = ~new_U3476 | ~new_R1117_U48;
  assign new_R1117_U214 = ~new_U3480 | ~new_R1117_U32;
  assign new_R1117_U215 = ~new_R1117_U94;
  assign new_R1117_U216 = ~new_R1117_U68;
  assign new_R1117_U217 = ~new_R1117_U50;
  assign new_R1117_U218 = ~new_R1117_U88;
  assign new_R1117_U219 = ~new_R1117_U192;
  assign new_R1117_U220 = ~new_U3075 | ~new_R1117_U192;
  assign new_R1117_U221 = ~new_R1117_U56;
  assign new_R1117_U222 = ~new_U3472 | ~new_R1117_U42;
  assign new_R1117_U223 = ~new_R1117_U42 | ~new_R1117_U41;
  assign new_R1117_U224 = ~new_R1117_U223 | ~new_R1117_U46;
  assign new_R1117_U225 = ~new_U3061 | ~new_R1117_U206;
  assign new_R1117_U226 = ~new_U3478 | ~new_R1117_U47;
  assign new_R1117_U227 = ~new_U3068 | ~new_R1117_U36;
  assign new_R1117_U228 = ~new_U3064 | ~new_R1117_U35;
  assign new_R1117_U229 = ~new_R1117_U217 | ~new_R1117_U213;
  assign new_R1117_U230 = ~new_R1117_U6 | ~new_R1117_U229;
  assign new_R1117_U231 = ~new_U3474 | ~new_R1117_U49;
  assign new_R1117_U232 = ~new_U3478 | ~new_R1117_U47;
  assign new_R1117_U233 = ~new_R1117_U14 | ~new_R1117_U175;
  assign new_R1117_U234 = ~new_R1117_U51;
  assign new_R1117_U235 = ~new_R1117_U54;
  assign new_R1117_U236 = ~new_U3482 | ~new_R1117_U34;
  assign new_R1117_U237 = ~new_R1117_U34 | ~new_R1117_U33;
  assign new_R1117_U238 = ~new_R1117_U237 | ~new_R1117_U39;
  assign new_R1117_U239 = ~new_U3081 | ~new_R1117_U207;
  assign new_R1117_U240 = ~new_R1117_U171;
  assign new_R1117_U241 = ~new_U3484 | ~new_R1117_U53;
  assign new_R1117_U242 = ~new_R1117_U241 | ~new_R1117_U88;
  assign new_R1117_U243 = ~new_R1117_U235 | ~new_R1117_U33;
  assign new_R1117_U244 = ~new_R1117_U136 | ~new_R1117_U243;
  assign new_R1117_U245 = ~new_R1117_U54 | ~new_R1117_U214;
  assign new_R1117_U246 = ~new_R1117_U135 | ~new_R1117_U245;
  assign new_R1117_U247 = ~new_R1117_U33 | ~new_R1117_U214;
  assign new_R1117_U248 = ~new_R1117_U231 | ~new_R1117_U175;
  assign new_R1117_U249 = ~new_R1117_U55;
  assign new_R1117_U250 = ~new_U3064 | ~new_R1117_U35;
  assign new_R1117_U251 = ~new_R1117_U249 | ~new_R1117_U250;
  assign new_R1117_U252 = ~new_R1117_U138 | ~new_R1117_U251;
  assign new_R1117_U253 = ~new_R1117_U55 | ~new_R1117_U213;
  assign new_R1117_U254 = ~new_U3478 | ~new_R1117_U47;
  assign new_R1117_U255 = ~new_R1117_U137 | ~new_R1117_U253;
  assign new_R1117_U256 = ~new_U3064 | ~new_R1117_U35;
  assign new_R1117_U257 = ~new_R1117_U213 | ~new_R1117_U256;
  assign new_R1117_U258 = ~new_R1117_U231 | ~new_R1117_U50;
  assign new_R1117_U259 = ~new_R1117_U140 | ~new_R1117_U372;
  assign new_R1117_U260 = ~new_R1117_U41 | ~new_R1117_U212;
  assign new_R1117_U261 = ~new_U3488 | ~new_R1117_U84;
  assign new_R1117_U262 = ~new_U3060 | ~new_R1117_U86;
  assign new_R1117_U263 = ~new_U3059 | ~new_R1117_U87;
  assign new_R1117_U264 = ~new_R1117_U218 | ~new_R1117_U7;
  assign new_R1117_U265 = ~new_R1117_U8 | ~new_R1117_U264;
  assign new_R1117_U266 = ~new_U3488 | ~new_R1117_U84;
  assign new_R1117_U267 = ~new_R1117_U266 | ~new_R1117_U265;
  assign new_R1117_U268 = ~new_U3490 | ~new_R1117_U89;
  assign new_R1117_U269 = ~new_U3069 | ~new_R1117_U83;
  assign new_R1117_U270 = ~new_U3492 | ~new_R1117_U81;
  assign new_R1117_U271 = ~new_U3077 | ~new_R1117_U82;
  assign new_R1117_U272 = ~new_U3498 | ~new_R1117_U91;
  assign new_R1117_U273 = ~new_U3070 | ~new_R1117_U78;
  assign new_R1117_U274 = ~new_U3071 | ~new_R1117_U79;
  assign new_R1117_U275 = ~new_R1117_U215 | ~new_R1117_U9;
  assign new_R1117_U276 = ~new_R1117_U10 | ~new_R1117_U275;
  assign new_R1117_U277 = ~new_U3494 | ~new_R1117_U93;
  assign new_R1117_U278 = ~new_U3498 | ~new_R1117_U91;
  assign new_R1117_U279 = ~new_R1117_U17 | ~new_R1117_U198;
  assign new_R1117_U280 = ~new_R1117_U95;
  assign new_R1117_U281 = ~new_R1117_U195;
  assign new_R1117_U282 = ~new_U3500 | ~new_R1117_U76;
  assign new_R1117_U283 = ~new_U3066 | ~new_R1117_U77;
  assign new_R1117_U284 = ~new_R1117_U194;
  assign new_R1117_U285 = ~new_U3502 | ~new_R1117_U75;
  assign new_R1117_U286 = ~new_U3504 | ~new_R1117_U71;
  assign new_R1117_U287 = ~new_R1117_U73;
  assign new_R1117_U288 = ~new_U4037 | ~new_R1117_U70;
  assign new_R1117_U289 = ~new_U3073 | ~new_R1117_U72;
  assign new_R1117_U290 = ~new_U4034 | ~new_R1117_U63;
  assign new_R1117_U291 = ~new_U3063 | ~new_R1117_U66;
  assign new_R1117_U292 = ~new_U3058 | ~new_R1117_U67;
  assign new_R1117_U293 = ~new_R1117_U216 | ~new_R1117_U11;
  assign new_R1117_U294 = ~new_R1117_U12 | ~new_R1117_U293;
  assign new_R1117_U295 = ~new_U4036 | ~new_R1117_U65;
  assign new_R1117_U296 = ~new_U4034 | ~new_R1117_U63;
  assign new_R1117_U297 = ~new_R1117_U296 | ~new_R1117_U294;
  assign new_R1117_U298 = ~new_U4033 | ~new_R1117_U61;
  assign new_R1117_U299 = ~new_U3062 | ~new_R1117_U62;
  assign new_R1117_U300 = ~new_U4032 | ~new_R1117_U98;
  assign new_R1117_U301 = ~new_R1117_U300 | ~new_R1117_U184;
  assign new_R1117_U302 = ~new_U3055 | ~new_R1117_U97;
  assign new_R1117_U303 = ~new_R1117_U183;
  assign new_R1117_U304 = ~new_U4030 | ~new_R1117_U60;
  assign new_R1117_U305 = ~new_R1117_U60 | ~new_R1117_U59;
  assign new_R1117_U306 = ~new_R1117_U305 | ~new_R1117_U100;
  assign new_R1117_U307 = ~new_U3050 | ~new_R1117_U205;
  assign new_R1117_U308 = ~new_U4029 | ~new_R1117_U101;
  assign new_R1117_U309 = ~new_U3051 | ~new_R1117_U57;
  assign new_R1117_U310 = ~new_R1117_U59 | ~new_R1117_U211;
  assign new_R1117_U311 = ~new_U4034 | ~new_R1117_U63;
  assign new_R1117_U312 = ~new_U3058 | ~new_R1117_U67;
  assign new_R1117_U313 = ~new_R1117_U186 | ~new_R1117_U312;
  assign new_R1117_U314 = ~new_R1117_U295 | ~new_R1117_U68;
  assign new_R1117_U315 = ~new_R1117_U277 | ~new_R1117_U198;
  assign new_R1117_U316 = ~new_R1117_U106;
  assign new_R1117_U317 = ~new_U3071 | ~new_R1117_U79;
  assign new_R1117_U318 = ~new_R1117_U316 | ~new_R1117_U317;
  assign new_R1117_U319 = ~new_R1117_U165 | ~new_R1117_U318;
  assign new_R1117_U320 = ~new_R1117_U106 | ~new_R1117_U209;
  assign new_R1117_U321 = ~new_U3498 | ~new_R1117_U91;
  assign new_R1117_U322 = ~new_R1117_U164 | ~new_R1117_U320;
  assign new_R1117_U323 = ~new_U3071 | ~new_R1117_U79;
  assign new_R1117_U324 = ~new_R1117_U209 | ~new_R1117_U323;
  assign new_R1117_U325 = ~new_R1117_U277 | ~new_R1117_U94;
  assign new_R1117_U326 = ~new_U3059 | ~new_R1117_U87;
  assign new_R1117_U327 = ~new_R1117_U361 | ~new_R1117_U326;
  assign new_R1117_U328 = ~new_R1117_U169 | ~new_R1117_U327;
  assign new_R1117_U329 = ~new_R1117_U107 | ~new_R1117_U208;
  assign new_R1117_U330 = ~new_U3488 | ~new_R1117_U84;
  assign new_R1117_U331 = ~new_R1117_U168 | ~new_R1117_U329;
  assign new_R1117_U332 = ~new_U3059 | ~new_R1117_U87;
  assign new_R1117_U333 = ~new_R1117_U208 | ~new_R1117_U332;
  assign new_R1117_U334 = ~new_U3074 | ~new_R1117_U44;
  assign new_R1117_U335 = ~new_U3075 | ~new_R1117_U191;
  assign new_R1117_U336 = ~new_U3079 | ~new_R1117_U96;
  assign new_R1117_U337 = ~new_R1117_U132 | ~new_R1117_U175;
  assign new_R1117_U338 = ~new_R1117_U234 | ~new_R1117_U15;
  assign new_R1117_U339 = ~new_R1117_U269 | ~new_R1117_U267;
  assign new_R1117_U340 = ~new_R1117_U90;
  assign new_R1117_U341 = ~new_R1117_U340 | ~new_R1117_U270;
  assign new_R1117_U342 = ~new_R1117_U142 | ~new_R1117_U198;
  assign new_R1117_U343 = ~new_R1117_U280 | ~new_R1117_U282;
  assign new_R1117_U344 = ~new_R1117_U287 | ~new_R1117_U288;
  assign new_R1117_U345 = ~new_R1117_U105;
  assign new_R1117_U346 = ~new_R1117_U18 | ~new_R1117_U105;
  assign new_R1117_U347 = ~new_R1117_U103;
  assign new_R1117_U348 = ~new_R1117_U103 | ~new_R1117_U298;
  assign new_R1117_U349 = ~new_R1117_U105 | ~new_R1117_U295;
  assign new_R1117_U350 = ~new_R1117_U286 | ~new_R1117_U193;
  assign new_R1117_U351 = ~new_R1117_U190;
  assign new_R1117_U352 = ~new_R1117_U20 | ~new_R1117_U193;
  assign new_R1117_U353 = ~new_R1117_U189;
  assign new_R1117_U354 = ~new_R1117_U21 | ~new_R1117_U193;
  assign new_R1117_U355 = ~new_R1117_U185;
  assign new_R1117_U356 = ~new_R1117_U156 | ~new_R1117_U193;
  assign new_R1117_U357 = ~new_R1117_U104;
  assign new_R1117_U358 = ~new_R1117_U144 | ~new_R1117_U193;
  assign new_R1117_U359 = ~new_R1117_U184;
  assign new_R1117_U360 = ~new_R1117_U241 | ~new_R1117_U171;
  assign new_R1117_U361 = ~new_R1117_U107;
  assign new_R1117_U362 = ~new_R1117_U16 | ~new_R1117_U171;
  assign new_R1117_U363 = ~new_R1117_U200;
  assign new_R1117_U364 = ~new_R1117_U19 | ~new_R1117_U171;
  assign new_R1117_U365 = ~new_R1117_U199;
  assign new_R1117_U366 = ~new_R1117_U141 | ~new_R1117_U171;
  assign new_R1117_U367 = ~new_R1117_U198;
  assign new_R1117_U368 = ~new_R1117_U130 | ~new_R1117_U56;
  assign new_R1117_U369 = ~new_R1117_U175;
  assign new_R1117_U370 = ~new_R1117_U212 | ~new_R1117_U56;
  assign new_R1117_U371 = ~new_R1117_U139 | ~new_R1117_U370;
  assign new_R1117_U372 = ~new_R1117_U221 | ~new_R1117_U41;
  assign new_R1117_U373 = ~new_R1117_U152 | ~new_R1117_U183;
  assign new_R1117_U374 = ~new_R1117_U13 | ~new_R1117_U183;
  assign new_R1117_U375 = ~new_R1117_U149 | ~new_R1117_U374;
  assign new_R1117_U376 = ~new_R1117_U13 | ~new_R1117_U183;
  assign new_R1117_U377 = ~new_R1117_U180;
  assign new_R1117_U378 = ~new_R1117_U202 | ~new_R1117_U183;
  assign new_R1117_U379 = ~new_R1117_U181 | ~new_R1117_U378;
  assign new_R1117_U380 = ~new_R1117_U285 | ~new_R1117_U194;
  assign new_R1117_U381 = ~new_R1117_U193;
  assign new_R1117_U382 = ~new_R1117_U155 | ~new_R1117_U452;
  assign new_R1117_U383 = ~new_R1117_U158 | ~new_R1117_U357;
  assign new_R1117_U384 = ~new_U3484 | ~new_R1117_U53;
  assign new_R1117_U385 = ~new_U3080 | ~new_R1117_U52;
  assign new_R1117_U386 = ~new_R1117_U242 | ~new_R1117_U171;
  assign new_R1117_U387 = ~new_R1117_U240 | ~new_R1117_U170;
  assign new_R1117_U388 = ~new_U3482 | ~new_R1117_U34;
  assign new_R1117_U389 = ~new_U3081 | ~new_R1117_U39;
  assign new_R1117_U390 = ~new_U3482 | ~new_R1117_U34;
  assign new_R1117_U391 = ~new_U3081 | ~new_R1117_U39;
  assign new_R1117_U392 = ~new_R1117_U391 | ~new_R1117_U390;
  assign new_R1117_U393 = ~new_U3480 | ~new_R1117_U32;
  assign new_R1117_U394 = ~new_U3067 | ~new_R1117_U38;
  assign new_R1117_U395 = ~new_R1117_U247 | ~new_R1117_U54;
  assign new_R1117_U396 = ~new_R1117_U172 | ~new_R1117_U235;
  assign new_R1117_U397 = ~new_U3478 | ~new_R1117_U47;
  assign new_R1117_U398 = ~new_U3068 | ~new_R1117_U36;
  assign new_R1117_U399 = ~new_R1117_U398 | ~new_R1117_U397;
  assign new_R1117_U400 = ~new_U3476 | ~new_R1117_U48;
  assign new_R1117_U401 = ~new_U3064 | ~new_R1117_U35;
  assign new_R1117_U402 = ~new_R1117_U257 | ~new_R1117_U55;
  assign new_R1117_U403 = ~new_R1117_U173 | ~new_R1117_U249;
  assign new_R1117_U404 = ~new_U3474 | ~new_R1117_U49;
  assign new_R1117_U405 = ~new_U3057 | ~new_R1117_U37;
  assign new_R1117_U406 = ~new_R1117_U175 | ~new_R1117_U258;
  assign new_R1117_U407 = ~new_R1117_U369 | ~new_R1117_U174;
  assign new_R1117_U408 = ~new_U3472 | ~new_R1117_U42;
  assign new_R1117_U409 = ~new_U3061 | ~new_R1117_U46;
  assign new_R1117_U410 = ~new_U3472 | ~new_R1117_U42;
  assign new_R1117_U411 = ~new_U3061 | ~new_R1117_U46;
  assign new_R1117_U412 = ~new_R1117_U411 | ~new_R1117_U410;
  assign new_R1117_U413 = ~new_U3470 | ~new_R1117_U40;
  assign new_R1117_U414 = ~new_U3065 | ~new_R1117_U43;
  assign new_R1117_U415 = ~new_R1117_U260 | ~new_R1117_U56;
  assign new_R1117_U416 = ~new_R1117_U176 | ~new_R1117_U221;
  assign new_R1117_U417 = ~new_U4040 | ~new_R1117_U178;
  assign new_R1117_U418 = ~new_U3052 | ~new_R1117_U177;
  assign new_R1117_U419 = ~new_R1117_U418 | ~new_R1117_U417;
  assign new_R1117_U420 = ~new_U4040 | ~new_R1117_U178;
  assign new_R1117_U421 = ~new_U3052 | ~new_R1117_U177;
  assign new_R1117_U422 = ~new_R1117_U57 | ~new_U3051 | ~new_R1117_U419;
  assign new_R1117_U423 = ~new_U4029 | ~new_R1117_U22 | ~new_R1117_U101;
  assign new_R1117_U424 = ~new_U4029 | ~new_R1117_U101;
  assign new_R1117_U425 = ~new_U3051 | ~new_R1117_U57;
  assign new_R1117_U426 = ~new_R1117_U151;
  assign new_R1117_U427 = ~new_R1117_U377 | ~new_R1117_U426;
  assign new_R1117_U428 = ~new_R1117_U151 | ~new_R1117_U180;
  assign new_R1117_U429 = ~new_U4030 | ~new_R1117_U60;
  assign new_R1117_U430 = ~new_U3050 | ~new_R1117_U100;
  assign new_R1117_U431 = ~new_R1117_U430 | ~new_R1117_U429;
  assign new_R1117_U432 = ~new_U4030 | ~new_R1117_U60;
  assign new_R1117_U433 = ~new_U3050 | ~new_R1117_U100;
  assign new_R1117_U434 = ~new_R1117_U59 | ~new_R1117_U433 | ~new_R1117_U432;
  assign new_R1117_U435 = ~new_R1117_U431 | ~new_R1117_U205;
  assign new_R1117_U436 = ~new_U4031 | ~new_R1117_U58;
  assign new_R1117_U437 = ~new_U3054 | ~new_R1117_U99;
  assign new_R1117_U438 = ~new_R1117_U310 | ~new_R1117_U183;
  assign new_R1117_U439 = ~new_R1117_U303 | ~new_R1117_U182;
  assign new_R1117_U440 = ~new_U4032 | ~new_R1117_U98;
  assign new_R1117_U441 = ~new_U3055 | ~new_R1117_U97;
  assign new_R1117_U442 = ~new_R1117_U153;
  assign new_R1117_U443 = ~new_R1117_U359 | ~new_R1117_U442;
  assign new_R1117_U444 = ~new_R1117_U153 | ~new_R1117_U184;
  assign new_R1117_U445 = ~new_U4033 | ~new_R1117_U61;
  assign new_R1117_U446 = ~new_U3062 | ~new_R1117_U62;
  assign new_R1117_U447 = ~new_R1117_U154;
  assign new_R1117_U448 = ~new_R1117_U355 | ~new_R1117_U447;
  assign new_R1117_U449 = ~new_R1117_U154 | ~new_R1117_U185;
  assign new_R1117_U450 = ~new_U4034 | ~new_R1117_U63;
  assign new_R1117_U451 = ~new_U3063 | ~new_R1117_U66;
  assign new_R1117_U452 = ~new_R1117_U451 | ~new_R1117_U450;
  assign new_R1117_U453 = ~new_R1117_U186 | ~new_R1117_U452 | ~new_R1117_U104;
  assign new_R1117_U454 = ~new_R1117_U210 | ~new_R1117_U12 | ~new_R1117_U311;
  assign new_R1117_U455 = ~new_U4035 | ~new_R1117_U64;
  assign new_R1117_U456 = ~new_U3058 | ~new_R1117_U67;
  assign new_R1117_U457 = ~new_R1117_U104 | ~new_R1117_U313;
  assign new_R1117_U458 = ~new_R1117_U187 | ~new_R1117_U357;
  assign new_R1117_U459 = ~new_U4036 | ~new_R1117_U65;
  assign new_R1117_U460 = ~new_U3072 | ~new_R1117_U69;
  assign new_R1117_U461 = ~new_R1117_U189 | ~new_R1117_U314;
  assign new_R1117_U462 = ~new_R1117_U353 | ~new_R1117_U188;
  assign new_R1117_U463 = ~new_U4037 | ~new_R1117_U70;
  assign new_R1117_U464 = ~new_U3073 | ~new_R1117_U72;
  assign new_R1117_U465 = ~new_R1117_U159;
  assign new_R1117_U466 = ~new_R1117_U351 | ~new_R1117_U465;
  assign new_R1117_U467 = ~new_R1117_U159 | ~new_R1117_U190;
  assign new_R1117_U468 = ~new_U3468 | ~new_R1117_U45;
  assign new_R1117_U469 = ~new_U3075 | ~new_R1117_U191;
  assign new_R1117_U470 = ~new_R1117_U160;
  assign new_R1117_U471 = ~new_R1117_U219 | ~new_R1117_U470;
  assign new_R1117_U472 = ~new_R1117_U160 | ~new_R1117_U192;
  assign new_R1117_U473 = ~new_U3504 | ~new_R1117_U71;
  assign new_R1117_U474 = ~new_U3078 | ~new_R1117_U74;
  assign new_R1117_U475 = ~new_R1117_U161;
  assign new_R1117_U476 = ~new_R1117_U381 | ~new_R1117_U475;
  assign new_R1117_U477 = ~new_R1117_U161 | ~new_R1117_U193;
  assign new_R1117_U478 = ~new_U3502 | ~new_R1117_U75;
  assign new_R1117_U479 = ~new_U3079 | ~new_R1117_U96;
  assign new_R1117_U480 = ~new_R1117_U162;
  assign new_R1117_U481 = ~new_R1117_U284 | ~new_R1117_U480;
  assign new_R1117_U482 = ~new_R1117_U162 | ~new_R1117_U194;
  assign new_R1117_U483 = ~new_U3500 | ~new_R1117_U76;
  assign new_R1117_U484 = ~new_U3066 | ~new_R1117_U77;
  assign new_R1117_U485 = ~new_R1117_U163;
  assign new_R1117_U486 = ~new_R1117_U281 | ~new_R1117_U485;
  assign new_R1117_U487 = ~new_R1117_U163 | ~new_R1117_U195;
  assign new_R1117_U488 = ~new_U3498 | ~new_R1117_U91;
  assign new_R1117_U489 = ~new_U3070 | ~new_R1117_U78;
  assign new_R1117_U490 = ~new_R1117_U489 | ~new_R1117_U488;
  assign new_R1117_U491 = ~new_U3496 | ~new_R1117_U92;
  assign new_R1117_U492 = ~new_U3071 | ~new_R1117_U79;
  assign new_R1117_U493 = ~new_R1117_U324 | ~new_R1117_U106;
  assign new_R1117_U494 = ~new_R1117_U196 | ~new_R1117_U316;
  assign new_R1117_U495 = ~new_U3494 | ~new_R1117_U93;
  assign new_R1117_U496 = ~new_U3076 | ~new_R1117_U80;
  assign new_R1117_U497 = ~new_R1117_U198 | ~new_R1117_U325;
  assign new_R1117_U498 = ~new_R1117_U367 | ~new_R1117_U197;
  assign new_R1117_U499 = ~new_U3492 | ~new_R1117_U81;
  assign new_R1117_U500 = ~new_U3077 | ~new_R1117_U82;
  assign new_R1117_U501 = ~new_R1117_U166;
  assign new_R1117_U502 = ~new_R1117_U365 | ~new_R1117_U501;
  assign new_R1117_U503 = ~new_R1117_U166 | ~new_R1117_U199;
  assign new_R1117_U504 = ~new_U3490 | ~new_R1117_U89;
  assign new_R1117_U505 = ~new_U3069 | ~new_R1117_U83;
  assign new_R1117_U506 = ~new_R1117_U167;
  assign new_R1117_U507 = ~new_R1117_U363 | ~new_R1117_U506;
  assign new_R1117_U508 = ~new_R1117_U167 | ~new_R1117_U200;
  assign new_R1117_U509 = ~new_U3488 | ~new_R1117_U84;
  assign new_R1117_U510 = ~new_U3060 | ~new_R1117_U86;
  assign new_R1117_U511 = ~new_R1117_U510 | ~new_R1117_U509;
  assign new_R1117_U512 = ~new_U3486 | ~new_R1117_U85;
  assign new_R1117_U513 = ~new_U3059 | ~new_R1117_U87;
  assign new_R1117_U514 = ~new_R1117_U107 | ~new_R1117_U333;
  assign new_R1117_U515 = ~new_R1117_U201 | ~new_R1117_U361;
  assign new_R1375_U6 = new_R1375_U164 & new_R1375_U163;
  assign new_R1375_U7 = new_R1375_U172 & new_R1375_U173;
  assign new_R1375_U8 = new_R1375_U171 & new_R1375_U96 & new_R1375_U7 & new_R1375_U174;
  assign new_R1375_U9 = new_R1375_U97 & new_R1375_U8;
  assign new_R1375_U10 = new_R1375_U98 & new_R1375_U9;
  assign new_R1375_U11 = new_R1375_U181 & new_R1375_U182;
  assign new_R1375_U12 = new_R1375_U23 & new_R1375_U183;
  assign new_R1375_U13 = new_R1375_U186 & new_R1375_U185 & new_R1375_U184;
  assign new_R1375_U14 = new_R1375_U152 & new_R1375_U103 & new_R1375_U13 & new_R1375_U191;
  assign new_R1375_U15 = new_R1375_U157 & new_R1375_U155 & new_R1375_U154 & new_R1375_U153;
  assign new_R1375_U16 = new_R1375_U169 & new_R1375_U24 & new_R1375_U158 & new_R1375_U165 & new_R1375_U168;
  assign new_R1375_U17 = new_R1375_U109 & new_R1375_U24 & new_R1375_U10 & new_R1375_U179;
  assign new_R1375_U18 = new_R1375_U100 & new_R1375_U22;
  assign new_R1375_U19 = new_R1375_U10 & new_R1375_U165;
  assign new_R1375_U20 = new_R1375_U34 & new_R1375_U154 & new_U4030 & new_R1375_U155;
  assign new_R1375_U21 = new_R1375_U27 & new_R1375_U155 & new_U4029 & new_R1375_U154;
  assign new_R1375_U22 = new_R1375_U99 & new_R1375_U10 & new_R1375_U12;
  assign new_R1375_U23 = new_R1375_U178 & new_R1375_U179 & new_R1375_U11 & new_R1375_U180;
  assign new_R1375_U24 = new_R1375_U161 & new_R1375_U162 & new_R1375_U160;
  assign new_R1375_U25 = new_R1375_U100 & new_R1375_U165;
  assign new_R1375_U26 = ~new_R1375_U141 | ~new_R1375_U144 | ~new_R1375_U149 | ~new_R1375_U147 | ~new_R1375_U146;
  assign new_R1375_U27 = ~new_U3051;
  assign new_R1375_U28 = ~new_U3054;
  assign new_R1375_U29 = ~new_U4032;
  assign new_R1375_U30 = ~new_U4031;
  assign new_R1375_U31 = ~new_U4038;
  assign new_R1375_U32 = ~new_U3056;
  assign new_R1375_U33 = ~new_U3052;
  assign new_R1375_U34 = ~new_U3050;
  assign new_R1375_U35 = ~new_U3057;
  assign new_R1375_U36 = ~new_U3061;
  assign new_R1375_U37 = ~new_U3065;
  assign new_R1375_U38 = ~new_U3478;
  assign new_R1375_U39 = ~new_U3064;
  assign new_R1375_U40 = ~new_U4034;
  assign new_R1375_U41 = ~new_U4033;
  assign new_R1375_U42 = ~new_U3058;
  assign new_R1375_U43 = ~new_U3077;
  assign new_R1375_U44 = ~new_U3071;
  assign new_R1375_U45 = ~new_U3073;
  assign new_R1375_U46 = ~new_U3072;
  assign new_R1375_U47 = ~new_U3502;
  assign new_R1375_U48 = ~new_U3066;
  assign new_R1375_U49 = ~new_U3079;
  assign new_R1375_U50 = ~new_U3078;
  assign new_R1375_U51 = ~new_U3070;
  assign new_R1375_U52 = ~new_U3076;
  assign new_R1375_U53 = ~new_U3069;
  assign new_R1375_U54 = ~new_U3068;
  assign new_R1375_U55 = ~new_U3490;
  assign new_R1375_U56 = ~new_U3060;
  assign new_R1375_U57 = ~new_U3059;
  assign new_R1375_U58 = ~new_U3067;
  assign new_R1375_U59 = ~new_U3081;
  assign new_R1375_U60 = ~new_U3080;
  assign new_R1375_U61 = ~new_U3063;
  assign new_R1375_U62 = ~new_U3055;
  assign new_R1375_U63 = ~new_U3062;
  assign new_R1375_U64 = ~new_U3468;
  assign new_R1375_U65 = ~new_U3075;
  assign new_R1375_U66 = ~new_U3053;
  assign new_R1375_U67 = ~new_U3488;
  assign new_R1375_U68 = ~new_U3484;
  assign new_R1375_U69 = ~new_U3496;
  assign new_R1375_U70 = ~new_U3476;
  assign new_R1375_U71 = ~new_U3472;
  assign new_R1375_U72 = ~new_U3504;
  assign new_R1375_U73 = ~new_U3492;
  assign new_R1375_U74 = ~new_U3480;
  assign new_R1375_U75 = ~new_U4037;
  assign new_R1375_U76 = ~new_U3498;
  assign new_R1375_U77 = ~new_U3494;
  assign new_R1375_U78 = ~new_U3486;
  assign new_R1375_U79 = ~new_U3482;
  assign new_R1375_U80 = ~new_U3474;
  assign new_R1375_U81 = ~new_U3470;
  assign new_R1375_U82 = ~new_U4036;
  assign new_R1375_U83 = ~new_U4035;
  assign new_R1375_U84 = ~new_U3500;
  assign new_R1375_U85 = ~new_U4030;
  assign new_R1375_U86 = ~new_U4029;
  assign new_R1375_U87 = ~new_U4040;
  assign new_R1375_U88 = ~new_U4039;
  assign new_R1375_U89 = ~new_R1375_U198 | ~new_R1375_U197;
  assign new_R1375_U90 = new_U4032 & new_R1375_U62;
  assign new_R1375_U91 = new_U3063 & new_R1375_U40;
  assign new_R1375_U92 = new_U3064 & new_R1375_U70;
  assign new_R1375_U93 = new_U3058 & new_R1375_U83;
  assign new_R1375_U94 = new_U3060 & new_R1375_U67;
  assign new_R1375_U95 = new_U3066 & new_R1375_U84;
  assign new_R1375_U96 = new_R1375_U169 & new_R1375_U168;
  assign new_R1375_U97 = new_R1375_U175 & new_R1375_U167;
  assign new_R1375_U98 = new_R1375_U176 & new_R1375_U166;
  assign new_R1375_U99 = new_R1375_U165 & new_R1375_U152;
  assign new_R1375_U100 = new_R1375_U24 & new_R1375_U158;
  assign new_R1375_U101 = new_R1375_U15 & new_R1375_U65;
  assign new_R1375_U102 = new_R1375_U13 & new_U3468;
  assign new_R1375_U103 = new_R1375_U189 & new_R1375_U190;
  assign new_R1375_U104 = new_R1375_U192 & new_R1375_U156;
  assign new_R1375_U105 = new_R1375_U15 & new_R1375_U12 & new_R1375_U100 & new_R1375_U14 & new_R1375_U10;
  assign new_R1375_U106 = new_R1375_U156 & new_R1375_U53;
  assign new_R1375_U107 = new_R1375_U15 & new_R1375_U166;
  assign new_R1375_U108 = new_R1375_U15 & new_R1375_U56;
  assign new_R1375_U109 = new_R1375_U158 & new_R1375_U165 & new_R1375_U178;
  assign new_R1375_U110 = new_R1375_U15 & new_R1375_U60;
  assign new_R1375_U111 = new_R1375_U15 & new_R1375_U44;
  assign new_R1375_U112 = new_U3496 & new_R1375_U8;
  assign new_R1375_U113 = new_R1375_U156 & new_R1375_U54;
  assign new_R1375_U114 = new_U3478 & new_R1375_U15;
  assign new_R1375_U115 = new_R1375_U156 & new_R1375_U39;
  assign new_R1375_U116 = new_R1375_U15 & new_R1375_U12 & new_R1375_U100 & new_R1375_U19 & new_U3476;
  assign new_R1375_U117 = new_R1375_U156 & new_R1375_U184 & new_R1375_U36;
  assign new_R1375_U118 = new_R1375_U15 & new_R1375_U50;
  assign new_R1375_U119 = new_R1375_U15 & new_R1375_U43;
  assign new_R1375_U120 = new_R1375_U15 & new_R1375_U58;
  assign new_R1375_U121 = new_U3480 & new_R1375_U11;
  assign new_R1375_U122 = new_R1375_U156 & new_R1375_U169 & new_R1375_U45;
  assign new_R1375_U123 = new_R1375_U156 & new_R1375_U51;
  assign new_R1375_U124 = new_R1375_U15 & new_R1375_U171;
  assign new_R1375_U125 = new_U3498 & new_R1375_U7;
  assign new_R1375_U126 = new_R1375_U156 & new_R1375_U52;
  assign new_R1375_U127 = new_R1375_U15 & new_R1375_U167;
  assign new_R1375_U128 = new_U3494 & new_R1375_U8;
  assign new_R1375_U129 = new_R1375_U156 & new_R1375_U57;
  assign new_R1375_U130 = new_R1375_U15 & new_R1375_U178 & new_R1375_U100 & new_R1375_U19 & new_U3486;
  assign new_R1375_U131 = new_R1375_U156 & new_R1375_U181 & new_R1375_U59;
  assign new_R1375_U132 = new_R1375_U15 & new_R1375_U35;
  assign new_R1375_U133 = new_R1375_U156 & new_R1375_U37 & new_R1375_U185 & new_R1375_U184;
  assign new_R1375_U134 = new_R1375_U218 & new_R1375_U217;
  assign new_R1375_U135 = new_R1375_U219 & new_R1375_U156;
  assign new_R1375_U136 = new_R1375_U156 & new_R1375_U172 & new_R1375_U49;
  assign new_R1375_U137 = new_R1375_U15 & new_R1375_U48;
  assign new_R1375_U138 = new_U3500 & new_R1375_U7;
  assign new_R1375_U139 = new_R1375_U199 & new_R1375_U193;
  assign new_R1375_U140 = new_R1375_U200 & new_R1375_U201 & new_R1375_U202;
  assign new_R1375_U141 = new_R1375_U140 & new_R1375_U139 & new_R1375_U187 & new_R1375_U150;
  assign new_R1375_U142 = new_R1375_U204 & new_R1375_U203;
  assign new_R1375_U143 = new_R1375_U208 & new_R1375_U207;
  assign new_R1375_U144 = new_R1375_U209 & new_R1375_U143 & new_R1375_U142 & new_R1375_U206 & new_R1375_U205;
  assign new_R1375_U145 = new_R1375_U211 & new_R1375_U210;
  assign new_R1375_U146 = new_R1375_U145 & new_R1375_U213 & new_R1375_U212;
  assign new_R1375_U147 = new_R1375_U216 & new_R1375_U215 & new_R1375_U214;
  assign new_R1375_U148 = new_R1375_U223 & new_R1375_U224 & new_R1375_U225;
  assign new_R1375_U149 = new_R1375_U148 & new_R1375_U222 & new_R1375_U221 & new_R1375_U220;
  assign new_R1375_U150 = ~new_R1375_U156 | ~new_R1375_U196 | ~new_R1375_U15;
  assign new_R1375_U151 = ~new_U3478 | ~new_R1375_U54;
  assign new_R1375_U152 = ~new_R1375_U92 | ~new_R1375_U151;
  assign new_R1375_U153 = ~new_U4038 | ~new_R1375_U66;
  assign new_R1375_U154 = ~new_U3056 | ~new_R1375_U88;
  assign new_R1375_U155 = ~new_U3052 | ~new_R1375_U87;
  assign new_R1375_U156 = ~new_U3051 | ~new_R1375_U86;
  assign new_R1375_U157 = ~new_U3050 | ~new_R1375_U85;
  assign new_R1375_U158 = ~new_U3054 | ~new_R1375_U30;
  assign new_R1375_U159 = ~new_U4033 | ~new_R1375_U63;
  assign new_R1375_U160 = ~new_R1375_U91 | ~new_R1375_U159;
  assign new_R1375_U161 = ~new_U3055 | ~new_R1375_U29;
  assign new_R1375_U162 = ~new_U3062 | ~new_R1375_U41;
  assign new_R1375_U163 = ~new_U4034 | ~new_R1375_U61;
  assign new_R1375_U164 = ~new_U4033 | ~new_R1375_U63;
  assign new_R1375_U165 = ~new_R1375_U93 | ~new_R1375_U6;
  assign new_R1375_U166 = ~new_U3077 | ~new_R1375_U73;
  assign new_R1375_U167 = ~new_U3071 | ~new_R1375_U69;
  assign new_R1375_U168 = ~new_U3073 | ~new_R1375_U75;
  assign new_R1375_U169 = ~new_U3072 | ~new_R1375_U82;
  assign new_R1375_U170 = ~new_U3502 | ~new_R1375_U49;
  assign new_R1375_U171 = ~new_R1375_U95 | ~new_R1375_U170;
  assign new_R1375_U172 = ~new_U3078 | ~new_R1375_U72;
  assign new_R1375_U173 = ~new_U3079 | ~new_R1375_U47;
  assign new_R1375_U174 = ~new_U3070 | ~new_R1375_U76;
  assign new_R1375_U175 = ~new_U3076 | ~new_R1375_U77;
  assign new_R1375_U176 = ~new_U3069 | ~new_R1375_U55;
  assign new_R1375_U177 = ~new_U3490 | ~new_R1375_U53;
  assign new_R1375_U178 = ~new_R1375_U94 | ~new_R1375_U177;
  assign new_R1375_U179 = ~new_U3059 | ~new_R1375_U78;
  assign new_R1375_U180 = ~new_U3067 | ~new_R1375_U74;
  assign new_R1375_U181 = ~new_U3080 | ~new_R1375_U68;
  assign new_R1375_U182 = ~new_U3081 | ~new_R1375_U79;
  assign new_R1375_U183 = ~new_U3068 | ~new_R1375_U38;
  assign new_R1375_U184 = ~new_U3057 | ~new_R1375_U80;
  assign new_R1375_U185 = ~new_U3061 | ~new_R1375_U71;
  assign new_R1375_U186 = ~new_U3065 | ~new_R1375_U81;
  assign new_R1375_U187 = ~new_R1375_U101 | ~new_R1375_U156 | ~new_R1375_U102 | ~new_R1375_U18;
  assign new_R1375_U188 = ~new_U3464 | ~new_U3147;
  assign new_R1375_U189 = ~new_U3074 | ~new_R1375_U188;
  assign new_R1375_U190 = ~new_U3075 | ~new_R1375_U64;
  assign new_R1375_U191 = new_U3464 | new_U3147;
  assign new_R1375_U192 = ~new_U3058 | ~new_R1375_U83;
  assign new_R1375_U193 = ~new_R1375_U104 | ~new_R1375_U105;
  assign new_R1375_U194 = ~new_R1375_U90 | ~new_R1375_U158;
  assign new_R1375_U195 = ~new_U4031 | ~new_R1375_U28;
  assign new_R1375_U196 = ~new_R1375_U195 | ~new_R1375_U194;
  assign new_R1375_U197 = ~new_R1375_U33 | ~new_R1375_U154 | ~new_U4040;
  assign new_R1375_U198 = ~new_U4039 | ~new_R1375_U32;
  assign new_R1375_U199 = ~new_U3053 | ~new_R1375_U31;
  assign new_R1375_U200 = ~new_R1375_U106 | ~new_R1375_U107 | ~new_R1375_U25 | ~new_U3490 | ~new_R1375_U9;
  assign new_R1375_U201 = ~new_R1375_U108 | ~new_R1375_U156 | ~new_R1375_U100 | ~new_R1375_U19 | ~new_U3488;
  assign new_R1375_U202 = ~new_R1375_U110 | ~new_R1375_U156 | ~new_U3484 | ~new_R1375_U17;
  assign new_R1375_U203 = ~new_R1375_U111 | ~new_R1375_U156 | ~new_R1375_U112 | ~new_R1375_U25;
  assign new_R1375_U204 = ~new_R1375_U113 | ~new_R1375_U114 | ~new_R1375_U25 | ~new_R1375_U10 | ~new_R1375_U23;
  assign new_R1375_U205 = ~new_R1375_U115 | ~new_R1375_U116;
  assign new_R1375_U206 = ~new_R1375_U117 | ~new_R1375_U15 | ~new_R1375_U18 | ~new_U3472;
  assign new_R1375_U207 = ~new_R1375_U118 | ~new_R1375_U156 | ~new_U3504 | ~new_R1375_U16;
  assign new_R1375_U208 = ~new_R1375_U119 | ~new_R1375_U156 | ~new_R1375_U25 | ~new_U3492 | ~new_R1375_U9;
  assign new_R1375_U209 = ~new_R1375_U120 | ~new_R1375_U156 | ~new_R1375_U121 | ~new_R1375_U17;
  assign new_R1375_U210 = ~new_R1375_U122 | ~new_R1375_U15 | ~new_R1375_U25 | ~new_U4037;
  assign new_R1375_U211 = ~new_R1375_U123 | ~new_R1375_U124 | ~new_R1375_U125 | ~new_R1375_U16;
  assign new_R1375_U212 = ~new_R1375_U126 | ~new_R1375_U127 | ~new_R1375_U128 | ~new_R1375_U25;
  assign new_R1375_U213 = ~new_R1375_U129 | ~new_R1375_U130;
  assign new_R1375_U214 = ~new_R1375_U131 | ~new_R1375_U15 | ~new_R1375_U17 | ~new_U3482;
  assign new_R1375_U215 = ~new_R1375_U132 | ~new_R1375_U156 | ~new_U3474 | ~new_R1375_U18;
  assign new_R1375_U216 = ~new_R1375_U133 | ~new_R1375_U15 | ~new_R1375_U100 | ~new_U3470 | ~new_R1375_U22;
  assign new_R1375_U217 = ~new_U4036 | ~new_R1375_U46;
  assign new_R1375_U218 = ~new_U4035 | ~new_R1375_U42;
  assign new_R1375_U219 = ~new_R1375_U134 | ~new_R1375_U6;
  assign new_R1375_U220 = ~new_R1375_U135 | ~new_R1375_U25 | ~new_R1375_U15;
  assign new_R1375_U221 = ~new_R1375_U136 | ~new_R1375_U15 | ~new_U3502 | ~new_R1375_U16;
  assign new_R1375_U222 = ~new_R1375_U137 | ~new_R1375_U156 | ~new_R1375_U138 | ~new_R1375_U16;
  assign new_R1375_U223 = ~new_R1375_U156 | ~new_R1375_U20 | ~new_R1375_U153;
  assign new_R1375_U224 = ~new_R1375_U21 | ~new_R1375_U153;
  assign new_R1375_U225 = ~new_R1375_U89 | ~new_R1375_U153;
  assign new_R1352_U6 = new_U3056 & new_R1352_U7;
  assign new_R1352_U7 = ~new_U3053;
  assign new_R1207_U6 = new_R1207_U231 & new_R1207_U230;
  assign new_R1207_U7 = new_R1207_U211 & new_R1207_U264;
  assign new_R1207_U8 = new_R1207_U266 & new_R1207_U265;
  assign new_R1207_U9 = new_R1207_U212 & new_R1207_U275;
  assign new_R1207_U10 = new_R1207_U277 & new_R1207_U276;
  assign new_R1207_U11 = new_R1207_U106 & new_R1207_U293;
  assign new_R1207_U12 = new_R1207_U295 & new_R1207_U294;
  assign new_R1207_U13 = new_R1207_U234 & new_R1207_U229 & new_R1207_U216;
  assign new_R1207_U14 = new_R1207_U239 & new_R1207_U217;
  assign new_R1207_U15 = new_R1207_U7 & new_R1207_U244;
  assign new_R1207_U16 = new_R1207_U9 & new_R1207_U280;
  assign new_R1207_U17 = new_R1207_U11 & new_R1207_U298;
  assign new_R1207_U18 = new_R1207_U15 & new_R1207_U271;
  assign new_R1207_U19 = new_R1207_U291 & new_R1207_U289;
  assign new_R1207_U20 = new_R1207_U19 & new_R1207_U17;
  assign new_R1207_U21 = new_R1207_U20 & new_R1207_U301;
  assign new_R1207_U22 = new_R1207_U457 & new_R1207_U106;
  assign new_R1207_U23 = new_R1207_U423 & new_R1207_U422;
  assign new_R1207_U24 = ~new_R1207_U334 | ~new_R1207_U337;
  assign new_R1207_U25 = ~new_R1207_U325 | ~new_R1207_U328;
  assign new_R1207_U26 = ~new_R1207_U359 | ~new_R1207_U387 | ~new_R1207_U388 | ~new_R1207_U459 | ~new_R1207_U458;
  assign new_R1207_U27 = new_R1207_U344 & new_R1207_U313;
  assign new_R1207_U28 = ~new_R1207_U343 | ~new_R1207_U182 | ~new_R1207_U206;
  assign new_R1207_U29 = ~new_R1207_U262 | ~new_R1207_U383;
  assign new_R1207_U30 = ~new_R1207_U255 | ~new_R1207_U258;
  assign new_R1207_U31 = ~new_R1207_U247 | ~new_R1207_U249;
  assign new_R1207_U32 = ~new_R1207_U195 | ~new_R1207_U340;
  assign new_R1207_U33 = ~new_U3067;
  assign new_R1207_U34 = ~new_U3067 | ~new_R1207_U39;
  assign new_R1207_U35 = ~new_U3081;
  assign new_R1207_U36 = ~new_U3476;
  assign new_R1207_U37 = ~new_U3478;
  assign new_R1207_U38 = ~new_U3474;
  assign new_R1207_U39 = ~new_U3480;
  assign new_R1207_U40 = ~new_U3482;
  assign new_R1207_U41 = ~new_U3065;
  assign new_R1207_U42 = ~new_U3065 | ~new_R1207_U44;
  assign new_R1207_U43 = ~new_U3061;
  assign new_R1207_U44 = ~new_U3470;
  assign new_R1207_U45 = ~new_U3464;
  assign new_R1207_U46 = ~new_U3075;
  assign new_R1207_U47 = ~new_U3472;
  assign new_R1207_U48 = ~new_U3068;
  assign new_R1207_U49 = ~new_U3064;
  assign new_R1207_U50 = ~new_U3057;
  assign new_R1207_U51 = ~new_U3057 | ~new_R1207_U38;
  assign new_R1207_U52 = ~new_R1207_U235 | ~new_R1207_U233;
  assign new_R1207_U53 = ~new_U3484;
  assign new_R1207_U54 = ~new_U3080;
  assign new_R1207_U55 = ~new_R1207_U52 | ~new_R1207_U236;
  assign new_R1207_U56 = ~new_R1207_U51 | ~new_R1207_U251;
  assign new_R1207_U57 = ~new_R1207_U341 | ~new_R1207_U223 | ~new_R1207_U207;
  assign new_R1207_U58 = ~new_U4031;
  assign new_R1207_U59 = ~new_U4030;
  assign new_R1207_U60 = ~new_U3055;
  assign new_R1207_U61 = ~new_U4032;
  assign new_R1207_U62 = ~new_U3062;
  assign new_R1207_U63 = ~new_U4033;
  assign new_R1207_U64 = ~new_U3063;
  assign new_R1207_U65 = ~new_U3058;
  assign new_R1207_U66 = ~new_U3072;
  assign new_R1207_U67 = ~new_U4034;
  assign new_R1207_U68 = ~new_U4035;
  assign new_R1207_U69 = ~new_U3072 | ~new_R1207_U70;
  assign new_R1207_U70 = ~new_U4036;
  assign new_R1207_U71 = ~new_U3073;
  assign new_R1207_U72 = ~new_U3078;
  assign new_R1207_U73 = ~new_U4037;
  assign new_R1207_U74 = ~new_U3078 | ~new_R1207_U75;
  assign new_R1207_U75 = ~new_U3504;
  assign new_R1207_U76 = ~new_U3079;
  assign new_R1207_U77 = ~new_U3066;
  assign new_R1207_U78 = ~new_U3500;
  assign new_R1207_U79 = ~new_U3498;
  assign new_R1207_U80 = ~new_U3496;
  assign new_R1207_U81 = ~new_U3494;
  assign new_R1207_U82 = ~new_U3077;
  assign new_R1207_U83 = ~new_U3492;
  assign new_R1207_U84 = ~new_U3490;
  assign new_R1207_U85 = ~new_U3060;
  assign new_R1207_U86 = ~new_U3059;
  assign new_R1207_U87 = ~new_U3488;
  assign new_R1207_U88 = ~new_U3486;
  assign new_R1207_U89 = ~new_U3080 | ~new_R1207_U53;
  assign new_R1207_U90 = ~new_U3069;
  assign new_R1207_U91 = ~new_R1207_U347 | ~new_R1207_U271;
  assign new_R1207_U92 = ~new_U3070;
  assign new_R1207_U93 = ~new_U3071;
  assign new_R1207_U94 = ~new_U3076;
  assign new_R1207_U95 = ~new_U3076 | ~new_R1207_U81;
  assign new_R1207_U96 = ~new_R1207_U281 | ~new_R1207_U279;
  assign new_R1207_U97 = ~new_U3502;
  assign new_R1207_U98 = ~new_U3054;
  assign new_R1207_U99 = ~new_U3054 | ~new_R1207_U58;
  assign new_R1207_U100 = ~new_U3050;
  assign new_R1207_U101 = ~new_U4029;
  assign new_R1207_U102 = ~new_U3051;
  assign new_R1207_U103 = ~new_R1207_U356 | ~new_R1207_U302;
  assign new_R1207_U104 = ~new_R1207_U354 | ~new_R1207_U300;
  assign new_R1207_U105 = ~new_R1207_U352 | ~new_R1207_U292;
  assign new_R1207_U106 = ~new_U4035 | ~new_R1207_U65;
  assign new_R1207_U107 = ~new_R1207_U95 | ~new_R1207_U321;
  assign new_R1207_U108 = ~new_R1207_U372 | ~new_R1207_U89;
  assign new_R1207_U109 = ~new_U3074;
  assign new_R1207_U110 = ~new_R1207_U433 | ~new_R1207_U432;
  assign new_R1207_U111 = ~new_R1207_U449 | ~new_R1207_U448;
  assign new_R1207_U112 = ~new_R1207_U454 | ~new_R1207_U453;
  assign new_R1207_U113 = ~new_R1207_U472 | ~new_R1207_U471;
  assign new_R1207_U114 = ~new_R1207_U477 | ~new_R1207_U476;
  assign new_R1207_U115 = ~new_R1207_U482 | ~new_R1207_U481;
  assign new_R1207_U116 = ~new_R1207_U487 | ~new_R1207_U486;
  assign new_R1207_U117 = ~new_R1207_U492 | ~new_R1207_U491;
  assign new_R1207_U118 = ~new_R1207_U508 | ~new_R1207_U507;
  assign new_R1207_U119 = ~new_R1207_U513 | ~new_R1207_U512;
  assign new_R1207_U120 = ~new_R1207_U392 | ~new_R1207_U391;
  assign new_R1207_U121 = ~new_R1207_U401 | ~new_R1207_U400;
  assign new_R1207_U122 = ~new_R1207_U408 | ~new_R1207_U407;
  assign new_R1207_U123 = ~new_R1207_U412 | ~new_R1207_U411;
  assign new_R1207_U124 = ~new_R1207_U421 | ~new_R1207_U420;
  assign new_R1207_U125 = ~new_R1207_U444 | ~new_R1207_U443;
  assign new_R1207_U126 = ~new_R1207_U463 | ~new_R1207_U462;
  assign new_R1207_U127 = ~new_R1207_U467 | ~new_R1207_U466;
  assign new_R1207_U128 = ~new_R1207_U499 | ~new_R1207_U498;
  assign new_R1207_U129 = ~new_R1207_U503 | ~new_R1207_U502;
  assign new_R1207_U130 = ~new_R1207_U520 | ~new_R1207_U519;
  assign new_R1207_U131 = new_R1207_U225 & new_R1207_U215;
  assign new_R1207_U132 = new_R1207_U228 & new_R1207_U227;
  assign new_R1207_U133 = new_R1207_U14 & new_R1207_U13;
  assign new_R1207_U134 = new_R1207_U242 & new_R1207_U241;
  assign new_R1207_U135 = new_R1207_U346 & new_R1207_U134;
  assign new_R1207_U136 = new_R1207_U34 & new_R1207_U394 & new_R1207_U393;
  assign new_R1207_U137 = new_R1207_U397 & new_R1207_U217;
  assign new_R1207_U138 = new_R1207_U257 & new_R1207_U6;
  assign new_R1207_U139 = new_R1207_U404 & new_R1207_U216;
  assign new_R1207_U140 = new_R1207_U42 & new_R1207_U414 & new_R1207_U413;
  assign new_R1207_U141 = new_R1207_U417 & new_R1207_U215;
  assign new_R1207_U142 = new_R1207_U273 & new_R1207_U18;
  assign new_R1207_U143 = new_R1207_U16 & new_R1207_U285;
  assign new_R1207_U144 = new_R1207_U351 & new_R1207_U286;
  assign new_R1207_U145 = new_R1207_U21 & new_R1207_U303;
  assign new_R1207_U146 = new_R1207_U358 & new_R1207_U304;
  assign new_R1207_U147 = new_R1207_U305 & new_R1207_U214;
  assign new_R1207_U148 = new_R1207_U308 & new_R1207_U309;
  assign new_R1207_U149 = new_R1207_U311 & new_R1207_U426;
  assign new_R1207_U150 = new_R1207_U308 & new_R1207_U309;
  assign new_R1207_U151 = new_R1207_U23 & new_R1207_U312;
  assign new_R1207_U152 = ~new_R1207_U430 | ~new_R1207_U429;
  assign new_R1207_U153 = new_R1207_U436 & new_R1207_U214;
  assign new_R1207_U154 = new_R1207_U214 & new_R1207_U186;
  assign new_R1207_U155 = ~new_R1207_U446 | ~new_R1207_U445;
  assign new_R1207_U156 = ~new_R1207_U451 | ~new_R1207_U450;
  assign new_R1207_U157 = new_R1207_U22 & new_R1207_U298;
  assign new_R1207_U158 = new_R1207_U213 & new_R1207_U317;
  assign new_R1207_U159 = new_U3058 & new_R1207_U68;
  assign new_R1207_U160 = new_R1207_U19 & new_R1207_U298;
  assign new_R1207_U161 = new_R1207_U12 & new_R1207_U360 & new_R1207_U317;
  assign new_R1207_U162 = ~new_R1207_U469 | ~new_R1207_U468;
  assign new_R1207_U163 = ~new_R1207_U474 | ~new_R1207_U473;
  assign new_R1207_U164 = ~new_R1207_U479 | ~new_R1207_U478;
  assign new_R1207_U165 = ~new_R1207_U484 | ~new_R1207_U483;
  assign new_R1207_U166 = ~new_R1207_U489 | ~new_R1207_U488;
  assign new_R1207_U167 = new_R1207_U327 & new_R1207_U10;
  assign new_R1207_U168 = new_R1207_U495 & new_R1207_U212;
  assign new_R1207_U169 = ~new_R1207_U505 | ~new_R1207_U504;
  assign new_R1207_U170 = ~new_R1207_U510 | ~new_R1207_U509;
  assign new_R1207_U171 = new_R1207_U336 & new_R1207_U8;
  assign new_R1207_U172 = new_R1207_U516 & new_R1207_U211;
  assign new_R1207_U173 = new_R1207_U390 & new_R1207_U389;
  assign new_R1207_U174 = ~new_R1207_U135 | ~new_R1207_U345;
  assign new_R1207_U175 = new_R1207_U399 & new_R1207_U398;
  assign new_R1207_U176 = new_R1207_U406 & new_R1207_U405;
  assign new_R1207_U177 = new_R1207_U410 & new_R1207_U409;
  assign new_R1207_U178 = ~new_R1207_U132 | ~new_R1207_U380;
  assign new_R1207_U179 = new_R1207_U419 & new_R1207_U418;
  assign new_R1207_U180 = ~new_U4040;
  assign new_R1207_U181 = ~new_U3052;
  assign new_R1207_U182 = new_R1207_U428 & new_R1207_U427;
  assign new_R1207_U183 = ~new_R1207_U148 | ~new_R1207_U306;
  assign new_R1207_U184 = new_R1207_U440 & new_R1207_U439;
  assign new_R1207_U185 = new_R1207_U442 & new_R1207_U441;
  assign new_R1207_U186 = ~new_R1207_U146 | ~new_R1207_U370;
  assign new_R1207_U187 = ~new_R1207_U357 | ~new_R1207_U367;
  assign new_R1207_U188 = ~new_R1207_U355 | ~new_R1207_U365;
  assign new_R1207_U189 = new_R1207_U461 & new_R1207_U460;
  assign new_R1207_U190 = ~new_R1207_U69 | ~new_R1207_U315;
  assign new_R1207_U191 = new_R1207_U465 & new_R1207_U464;
  assign new_R1207_U192 = ~new_R1207_U353 | ~new_R1207_U363;
  assign new_R1207_U193 = ~new_R1207_U361 | ~new_R1207_U74;
  assign new_R1207_U194 = ~new_U3468;
  assign new_R1207_U195 = ~new_U3464 | ~new_R1207_U109;
  assign new_R1207_U196 = ~new_R1207_U385 | ~new_R1207_U342;
  assign new_R1207_U197 = ~new_R1207_U144 | ~new_R1207_U350;
  assign new_R1207_U198 = ~new_R1207_U96 | ~new_R1207_U282;
  assign new_R1207_U199 = new_R1207_U497 & new_R1207_U496;
  assign new_R1207_U200 = new_R1207_U501 & new_R1207_U500;
  assign new_R1207_U201 = ~new_R1207_U378 | ~new_R1207_U349 | ~new_R1207_U274;
  assign new_R1207_U202 = ~new_R1207_U376 | ~new_R1207_U91;
  assign new_R1207_U203 = ~new_R1207_U374 | ~new_R1207_U270;
  assign new_R1207_U204 = new_R1207_U518 & new_R1207_U517;
  assign new_R1207_U205 = ~new_R1207_U153 | ~new_R1207_U186;
  assign new_R1207_U206 = ~new_R1207_U149 | ~new_R1207_U183;
  assign new_R1207_U207 = ~new_R1207_U195 | ~new_R1207_U194;
  assign new_R1207_U208 = ~new_R1207_U99;
  assign new_R1207_U209 = ~new_R1207_U42;
  assign new_R1207_U210 = ~new_R1207_U34;
  assign new_R1207_U211 = ~new_U3486 | ~new_R1207_U86;
  assign new_R1207_U212 = ~new_U3496 | ~new_R1207_U93;
  assign new_R1207_U213 = ~new_R1207_U106;
  assign new_R1207_U214 = ~new_U4031 | ~new_R1207_U98;
  assign new_R1207_U215 = ~new_U3470 | ~new_R1207_U41;
  assign new_R1207_U216 = ~new_U3476 | ~new_R1207_U49;
  assign new_R1207_U217 = ~new_U3480 | ~new_R1207_U33;
  assign new_R1207_U218 = ~new_R1207_U95;
  assign new_R1207_U219 = ~new_R1207_U69;
  assign new_R1207_U220 = ~new_R1207_U51;
  assign new_R1207_U221 = ~new_R1207_U89;
  assign new_R1207_U222 = ~new_R1207_U195;
  assign new_R1207_U223 = ~new_U3075 | ~new_R1207_U195;
  assign new_R1207_U224 = ~new_R1207_U57;
  assign new_R1207_U225 = ~new_U3472 | ~new_R1207_U43;
  assign new_R1207_U226 = ~new_R1207_U43 | ~new_R1207_U42;
  assign new_R1207_U227 = ~new_R1207_U226 | ~new_R1207_U47;
  assign new_R1207_U228 = ~new_U3061 | ~new_R1207_U209;
  assign new_R1207_U229 = ~new_U3478 | ~new_R1207_U48;
  assign new_R1207_U230 = ~new_U3068 | ~new_R1207_U37;
  assign new_R1207_U231 = ~new_U3064 | ~new_R1207_U36;
  assign new_R1207_U232 = ~new_R1207_U220 | ~new_R1207_U216;
  assign new_R1207_U233 = ~new_R1207_U6 | ~new_R1207_U232;
  assign new_R1207_U234 = ~new_U3474 | ~new_R1207_U50;
  assign new_R1207_U235 = ~new_U3478 | ~new_R1207_U48;
  assign new_R1207_U236 = ~new_R1207_U13 | ~new_R1207_U178;
  assign new_R1207_U237 = ~new_R1207_U52;
  assign new_R1207_U238 = ~new_R1207_U55;
  assign new_R1207_U239 = ~new_U3482 | ~new_R1207_U35;
  assign new_R1207_U240 = ~new_R1207_U35 | ~new_R1207_U34;
  assign new_R1207_U241 = ~new_R1207_U240 | ~new_R1207_U40;
  assign new_R1207_U242 = ~new_U3081 | ~new_R1207_U210;
  assign new_R1207_U243 = ~new_R1207_U174;
  assign new_R1207_U244 = ~new_U3484 | ~new_R1207_U54;
  assign new_R1207_U245 = ~new_R1207_U244 | ~new_R1207_U89;
  assign new_R1207_U246 = ~new_R1207_U238 | ~new_R1207_U34;
  assign new_R1207_U247 = ~new_R1207_U137 | ~new_R1207_U246;
  assign new_R1207_U248 = ~new_R1207_U55 | ~new_R1207_U217;
  assign new_R1207_U249 = ~new_R1207_U136 | ~new_R1207_U248;
  assign new_R1207_U250 = ~new_R1207_U34 | ~new_R1207_U217;
  assign new_R1207_U251 = ~new_R1207_U234 | ~new_R1207_U178;
  assign new_R1207_U252 = ~new_R1207_U56;
  assign new_R1207_U253 = ~new_U3064 | ~new_R1207_U36;
  assign new_R1207_U254 = ~new_R1207_U252 | ~new_R1207_U253;
  assign new_R1207_U255 = ~new_R1207_U139 | ~new_R1207_U254;
  assign new_R1207_U256 = ~new_R1207_U56 | ~new_R1207_U216;
  assign new_R1207_U257 = ~new_U3478 | ~new_R1207_U48;
  assign new_R1207_U258 = ~new_R1207_U138 | ~new_R1207_U256;
  assign new_R1207_U259 = ~new_U3064 | ~new_R1207_U36;
  assign new_R1207_U260 = ~new_R1207_U216 | ~new_R1207_U259;
  assign new_R1207_U261 = ~new_R1207_U234 | ~new_R1207_U51;
  assign new_R1207_U262 = ~new_R1207_U141 | ~new_R1207_U384;
  assign new_R1207_U263 = ~new_R1207_U42 | ~new_R1207_U215;
  assign new_R1207_U264 = ~new_U3488 | ~new_R1207_U85;
  assign new_R1207_U265 = ~new_U3060 | ~new_R1207_U87;
  assign new_R1207_U266 = ~new_U3059 | ~new_R1207_U88;
  assign new_R1207_U267 = ~new_R1207_U221 | ~new_R1207_U7;
  assign new_R1207_U268 = ~new_R1207_U8 | ~new_R1207_U267;
  assign new_R1207_U269 = ~new_U3488 | ~new_R1207_U85;
  assign new_R1207_U270 = ~new_R1207_U269 | ~new_R1207_U268;
  assign new_R1207_U271 = ~new_U3490 | ~new_R1207_U90;
  assign new_R1207_U272 = ~new_U3069 | ~new_R1207_U84;
  assign new_R1207_U273 = ~new_U3492 | ~new_R1207_U82;
  assign new_R1207_U274 = ~new_U3077 | ~new_R1207_U83;
  assign new_R1207_U275 = ~new_U3498 | ~new_R1207_U92;
  assign new_R1207_U276 = ~new_U3070 | ~new_R1207_U79;
  assign new_R1207_U277 = ~new_U3071 | ~new_R1207_U80;
  assign new_R1207_U278 = ~new_R1207_U218 | ~new_R1207_U9;
  assign new_R1207_U279 = ~new_R1207_U10 | ~new_R1207_U278;
  assign new_R1207_U280 = ~new_U3494 | ~new_R1207_U94;
  assign new_R1207_U281 = ~new_U3498 | ~new_R1207_U92;
  assign new_R1207_U282 = ~new_R1207_U16 | ~new_R1207_U201;
  assign new_R1207_U283 = ~new_R1207_U96;
  assign new_R1207_U284 = ~new_R1207_U198;
  assign new_R1207_U285 = ~new_U3500 | ~new_R1207_U77;
  assign new_R1207_U286 = ~new_U3066 | ~new_R1207_U78;
  assign new_R1207_U287 = ~new_R1207_U197;
  assign new_R1207_U288 = ~new_U3502 | ~new_R1207_U76;
  assign new_R1207_U289 = ~new_U3504 | ~new_R1207_U72;
  assign new_R1207_U290 = ~new_R1207_U74;
  assign new_R1207_U291 = ~new_U4037 | ~new_R1207_U71;
  assign new_R1207_U292 = ~new_U3073 | ~new_R1207_U73;
  assign new_R1207_U293 = ~new_U4034 | ~new_R1207_U64;
  assign new_R1207_U294 = ~new_U3063 | ~new_R1207_U67;
  assign new_R1207_U295 = ~new_U3058 | ~new_R1207_U68;
  assign new_R1207_U296 = ~new_R1207_U219 | ~new_R1207_U11;
  assign new_R1207_U297 = ~new_R1207_U12 | ~new_R1207_U296;
  assign new_R1207_U298 = ~new_U4036 | ~new_R1207_U66;
  assign new_R1207_U299 = ~new_U4034 | ~new_R1207_U64;
  assign new_R1207_U300 = ~new_R1207_U299 | ~new_R1207_U297;
  assign new_R1207_U301 = ~new_U4033 | ~new_R1207_U62;
  assign new_R1207_U302 = ~new_U3062 | ~new_R1207_U63;
  assign new_R1207_U303 = ~new_U4032 | ~new_R1207_U60;
  assign new_R1207_U304 = ~new_U3055 | ~new_R1207_U61;
  assign new_R1207_U305 = ~new_U4030 | ~new_R1207_U100;
  assign new_R1207_U306 = ~new_R1207_U147 | ~new_R1207_U186;
  assign new_R1207_U307 = ~new_R1207_U100 | ~new_R1207_U99;
  assign new_R1207_U308 = ~new_R1207_U307 | ~new_R1207_U59;
  assign new_R1207_U309 = ~new_U3050 | ~new_R1207_U208;
  assign new_R1207_U310 = ~new_R1207_U183;
  assign new_R1207_U311 = ~new_U4029 | ~new_R1207_U102;
  assign new_R1207_U312 = ~new_U3051 | ~new_R1207_U101;
  assign new_R1207_U313 = ~new_R1207_U154 | ~new_R1207_U205;
  assign new_R1207_U314 = ~new_R1207_U99 | ~new_R1207_U214;
  assign new_R1207_U315 = ~new_R1207_U298 | ~new_R1207_U192;
  assign new_R1207_U316 = ~new_R1207_U190;
  assign new_R1207_U317 = ~new_U4034 | ~new_R1207_U64;
  assign new_R1207_U318 = ~new_U3058 | ~new_R1207_U68;
  assign new_R1207_U319 = ~new_R1207_U106 | ~new_R1207_U318;
  assign new_R1207_U320 = ~new_R1207_U298 | ~new_R1207_U69;
  assign new_R1207_U321 = ~new_R1207_U280 | ~new_R1207_U201;
  assign new_R1207_U322 = ~new_R1207_U107;
  assign new_R1207_U323 = ~new_U3071 | ~new_R1207_U80;
  assign new_R1207_U324 = ~new_R1207_U322 | ~new_R1207_U323;
  assign new_R1207_U325 = ~new_R1207_U168 | ~new_R1207_U324;
  assign new_R1207_U326 = ~new_R1207_U107 | ~new_R1207_U212;
  assign new_R1207_U327 = ~new_U3498 | ~new_R1207_U92;
  assign new_R1207_U328 = ~new_R1207_U167 | ~new_R1207_U326;
  assign new_R1207_U329 = ~new_U3071 | ~new_R1207_U80;
  assign new_R1207_U330 = ~new_R1207_U212 | ~new_R1207_U329;
  assign new_R1207_U331 = ~new_R1207_U280 | ~new_R1207_U95;
  assign new_R1207_U332 = ~new_U3059 | ~new_R1207_U88;
  assign new_R1207_U333 = ~new_R1207_U373 | ~new_R1207_U332;
  assign new_R1207_U334 = ~new_R1207_U172 | ~new_R1207_U333;
  assign new_R1207_U335 = ~new_R1207_U108 | ~new_R1207_U211;
  assign new_R1207_U336 = ~new_U3488 | ~new_R1207_U85;
  assign new_R1207_U337 = ~new_R1207_U171 | ~new_R1207_U335;
  assign new_R1207_U338 = ~new_U3059 | ~new_R1207_U88;
  assign new_R1207_U339 = ~new_R1207_U211 | ~new_R1207_U338;
  assign new_R1207_U340 = ~new_U3074 | ~new_R1207_U45;
  assign new_R1207_U341 = ~new_U3075 | ~new_R1207_U194;
  assign new_R1207_U342 = ~new_U3079 | ~new_R1207_U97;
  assign new_R1207_U343 = ~new_R1207_U151 | ~new_R1207_U150 | ~new_R1207_U306;
  assign new_R1207_U344 = ~new_R1207_U184 | ~new_R1207_U205;
  assign new_R1207_U345 = ~new_R1207_U133 | ~new_R1207_U178;
  assign new_R1207_U346 = ~new_R1207_U237 | ~new_R1207_U14;
  assign new_R1207_U347 = ~new_R1207_U272 | ~new_R1207_U270;
  assign new_R1207_U348 = ~new_R1207_U91;
  assign new_R1207_U349 = ~new_R1207_U348 | ~new_R1207_U273;
  assign new_R1207_U350 = ~new_R1207_U143 | ~new_R1207_U201;
  assign new_R1207_U351 = ~new_R1207_U283 | ~new_R1207_U285;
  assign new_R1207_U352 = ~new_R1207_U290 | ~new_R1207_U291;
  assign new_R1207_U353 = ~new_R1207_U105;
  assign new_R1207_U354 = ~new_R1207_U17 | ~new_R1207_U105;
  assign new_R1207_U355 = ~new_R1207_U104;
  assign new_R1207_U356 = ~new_R1207_U104 | ~new_R1207_U301;
  assign new_R1207_U357 = ~new_R1207_U103;
  assign new_R1207_U358 = ~new_R1207_U103 | ~new_R1207_U303;
  assign new_R1207_U359 = ~new_R1207_U157 | ~new_R1207_U192;
  assign new_R1207_U360 = ~new_R1207_U105 | ~new_R1207_U298;
  assign new_R1207_U361 = ~new_R1207_U289 | ~new_R1207_U196;
  assign new_R1207_U362 = ~new_R1207_U193;
  assign new_R1207_U363 = ~new_R1207_U19 | ~new_R1207_U196;
  assign new_R1207_U364 = ~new_R1207_U192;
  assign new_R1207_U365 = ~new_R1207_U20 | ~new_R1207_U196;
  assign new_R1207_U366 = ~new_R1207_U188;
  assign new_R1207_U367 = ~new_R1207_U21 | ~new_R1207_U196;
  assign new_R1207_U368 = ~new_R1207_U187;
  assign new_R1207_U369 = ~new_R1207_U160 | ~new_R1207_U196;
  assign new_R1207_U370 = ~new_R1207_U145 | ~new_R1207_U196;
  assign new_R1207_U371 = ~new_R1207_U186;
  assign new_R1207_U372 = ~new_R1207_U244 | ~new_R1207_U174;
  assign new_R1207_U373 = ~new_R1207_U108;
  assign new_R1207_U374 = ~new_R1207_U15 | ~new_R1207_U174;
  assign new_R1207_U375 = ~new_R1207_U203;
  assign new_R1207_U376 = ~new_R1207_U18 | ~new_R1207_U174;
  assign new_R1207_U377 = ~new_R1207_U202;
  assign new_R1207_U378 = ~new_R1207_U142 | ~new_R1207_U174;
  assign new_R1207_U379 = ~new_R1207_U201;
  assign new_R1207_U380 = ~new_R1207_U131 | ~new_R1207_U57;
  assign new_R1207_U381 = ~new_R1207_U178;
  assign new_R1207_U382 = ~new_R1207_U215 | ~new_R1207_U57;
  assign new_R1207_U383 = ~new_R1207_U140 | ~new_R1207_U382;
  assign new_R1207_U384 = ~new_R1207_U224 | ~new_R1207_U42;
  assign new_R1207_U385 = ~new_R1207_U288 | ~new_R1207_U197;
  assign new_R1207_U386 = ~new_R1207_U196;
  assign new_R1207_U387 = ~new_R1207_U158 | ~new_R1207_U12;
  assign new_R1207_U388 = ~new_R1207_U159 | ~new_R1207_U457;
  assign new_R1207_U389 = ~new_U3484 | ~new_R1207_U54;
  assign new_R1207_U390 = ~new_U3080 | ~new_R1207_U53;
  assign new_R1207_U391 = ~new_R1207_U245 | ~new_R1207_U174;
  assign new_R1207_U392 = ~new_R1207_U243 | ~new_R1207_U173;
  assign new_R1207_U393 = ~new_U3482 | ~new_R1207_U35;
  assign new_R1207_U394 = ~new_U3081 | ~new_R1207_U40;
  assign new_R1207_U395 = ~new_U3482 | ~new_R1207_U35;
  assign new_R1207_U396 = ~new_U3081 | ~new_R1207_U40;
  assign new_R1207_U397 = ~new_R1207_U396 | ~new_R1207_U395;
  assign new_R1207_U398 = ~new_U3480 | ~new_R1207_U33;
  assign new_R1207_U399 = ~new_U3067 | ~new_R1207_U39;
  assign new_R1207_U400 = ~new_R1207_U250 | ~new_R1207_U55;
  assign new_R1207_U401 = ~new_R1207_U175 | ~new_R1207_U238;
  assign new_R1207_U402 = ~new_U3478 | ~new_R1207_U48;
  assign new_R1207_U403 = ~new_U3068 | ~new_R1207_U37;
  assign new_R1207_U404 = ~new_R1207_U403 | ~new_R1207_U402;
  assign new_R1207_U405 = ~new_U3476 | ~new_R1207_U49;
  assign new_R1207_U406 = ~new_U3064 | ~new_R1207_U36;
  assign new_R1207_U407 = ~new_R1207_U260 | ~new_R1207_U56;
  assign new_R1207_U408 = ~new_R1207_U176 | ~new_R1207_U252;
  assign new_R1207_U409 = ~new_U3474 | ~new_R1207_U50;
  assign new_R1207_U410 = ~new_U3057 | ~new_R1207_U38;
  assign new_R1207_U411 = ~new_R1207_U178 | ~new_R1207_U261;
  assign new_R1207_U412 = ~new_R1207_U381 | ~new_R1207_U177;
  assign new_R1207_U413 = ~new_U3472 | ~new_R1207_U43;
  assign new_R1207_U414 = ~new_U3061 | ~new_R1207_U47;
  assign new_R1207_U415 = ~new_U3472 | ~new_R1207_U43;
  assign new_R1207_U416 = ~new_U3061 | ~new_R1207_U47;
  assign new_R1207_U417 = ~new_R1207_U416 | ~new_R1207_U415;
  assign new_R1207_U418 = ~new_U3470 | ~new_R1207_U41;
  assign new_R1207_U419 = ~new_U3065 | ~new_R1207_U44;
  assign new_R1207_U420 = ~new_R1207_U263 | ~new_R1207_U57;
  assign new_R1207_U421 = ~new_R1207_U179 | ~new_R1207_U224;
  assign new_R1207_U422 = ~new_U4040 | ~new_R1207_U181;
  assign new_R1207_U423 = ~new_U3052 | ~new_R1207_U180;
  assign new_R1207_U424 = ~new_U4040 | ~new_R1207_U181;
  assign new_R1207_U425 = ~new_U3052 | ~new_R1207_U180;
  assign new_R1207_U426 = ~new_R1207_U425 | ~new_R1207_U424;
  assign new_R1207_U427 = ~new_R1207_U102 | ~new_U4029 | ~new_R1207_U23;
  assign new_R1207_U428 = ~new_U3051 | ~new_R1207_U426 | ~new_R1207_U101;
  assign new_R1207_U429 = ~new_U4029 | ~new_R1207_U102;
  assign new_R1207_U430 = ~new_U3051 | ~new_R1207_U101;
  assign new_R1207_U431 = ~new_R1207_U152;
  assign new_R1207_U432 = ~new_R1207_U310 | ~new_R1207_U431;
  assign new_R1207_U433 = ~new_R1207_U152 | ~new_R1207_U183;
  assign new_R1207_U434 = ~new_U4030 | ~new_R1207_U100;
  assign new_R1207_U435 = ~new_U3050 | ~new_R1207_U59;
  assign new_R1207_U436 = ~new_R1207_U435 | ~new_R1207_U434;
  assign new_R1207_U437 = ~new_U4030 | ~new_R1207_U100;
  assign new_R1207_U438 = ~new_U3050 | ~new_R1207_U59;
  assign new_R1207_U439 = ~new_R1207_U99 | ~new_R1207_U438 | ~new_R1207_U437;
  assign new_R1207_U440 = ~new_R1207_U436 | ~new_R1207_U208;
  assign new_R1207_U441 = ~new_U4031 | ~new_R1207_U98;
  assign new_R1207_U442 = ~new_U3054 | ~new_R1207_U58;
  assign new_R1207_U443 = ~new_R1207_U186 | ~new_R1207_U314;
  assign new_R1207_U444 = ~new_R1207_U371 | ~new_R1207_U185;
  assign new_R1207_U445 = ~new_U4032 | ~new_R1207_U60;
  assign new_R1207_U446 = ~new_U3055 | ~new_R1207_U61;
  assign new_R1207_U447 = ~new_R1207_U155;
  assign new_R1207_U448 = ~new_R1207_U368 | ~new_R1207_U447;
  assign new_R1207_U449 = ~new_R1207_U155 | ~new_R1207_U187;
  assign new_R1207_U450 = ~new_U4033 | ~new_R1207_U62;
  assign new_R1207_U451 = ~new_U3062 | ~new_R1207_U63;
  assign new_R1207_U452 = ~new_R1207_U156;
  assign new_R1207_U453 = ~new_R1207_U366 | ~new_R1207_U452;
  assign new_R1207_U454 = ~new_R1207_U156 | ~new_R1207_U188;
  assign new_R1207_U455 = ~new_U4034 | ~new_R1207_U64;
  assign new_R1207_U456 = ~new_U3063 | ~new_R1207_U67;
  assign new_R1207_U457 = ~new_R1207_U456 | ~new_R1207_U455;
  assign new_R1207_U458 = ~new_R1207_U69 | ~new_R1207_U161 | ~new_R1207_U369;
  assign new_R1207_U459 = ~new_R1207_U22 | ~new_R1207_U219;
  assign new_R1207_U460 = ~new_U4035 | ~new_R1207_U65;
  assign new_R1207_U461 = ~new_U3058 | ~new_R1207_U68;
  assign new_R1207_U462 = ~new_R1207_U319 | ~new_R1207_U190;
  assign new_R1207_U463 = ~new_R1207_U316 | ~new_R1207_U189;
  assign new_R1207_U464 = ~new_U4036 | ~new_R1207_U66;
  assign new_R1207_U465 = ~new_U3072 | ~new_R1207_U70;
  assign new_R1207_U466 = ~new_R1207_U192 | ~new_R1207_U320;
  assign new_R1207_U467 = ~new_R1207_U364 | ~new_R1207_U191;
  assign new_R1207_U468 = ~new_U4037 | ~new_R1207_U71;
  assign new_R1207_U469 = ~new_U3073 | ~new_R1207_U73;
  assign new_R1207_U470 = ~new_R1207_U162;
  assign new_R1207_U471 = ~new_R1207_U362 | ~new_R1207_U470;
  assign new_R1207_U472 = ~new_R1207_U162 | ~new_R1207_U193;
  assign new_R1207_U473 = ~new_U3468 | ~new_R1207_U46;
  assign new_R1207_U474 = ~new_U3075 | ~new_R1207_U194;
  assign new_R1207_U475 = ~new_R1207_U163;
  assign new_R1207_U476 = ~new_R1207_U222 | ~new_R1207_U475;
  assign new_R1207_U477 = ~new_R1207_U163 | ~new_R1207_U195;
  assign new_R1207_U478 = ~new_U3504 | ~new_R1207_U72;
  assign new_R1207_U479 = ~new_U3078 | ~new_R1207_U75;
  assign new_R1207_U480 = ~new_R1207_U164;
  assign new_R1207_U481 = ~new_R1207_U386 | ~new_R1207_U480;
  assign new_R1207_U482 = ~new_R1207_U164 | ~new_R1207_U196;
  assign new_R1207_U483 = ~new_U3502 | ~new_R1207_U76;
  assign new_R1207_U484 = ~new_U3079 | ~new_R1207_U97;
  assign new_R1207_U485 = ~new_R1207_U165;
  assign new_R1207_U486 = ~new_R1207_U287 | ~new_R1207_U485;
  assign new_R1207_U487 = ~new_R1207_U165 | ~new_R1207_U197;
  assign new_R1207_U488 = ~new_U3500 | ~new_R1207_U77;
  assign new_R1207_U489 = ~new_U3066 | ~new_R1207_U78;
  assign new_R1207_U490 = ~new_R1207_U166;
  assign new_R1207_U491 = ~new_R1207_U284 | ~new_R1207_U490;
  assign new_R1207_U492 = ~new_R1207_U166 | ~new_R1207_U198;
  assign new_R1207_U493 = ~new_U3498 | ~new_R1207_U92;
  assign new_R1207_U494 = ~new_U3070 | ~new_R1207_U79;
  assign new_R1207_U495 = ~new_R1207_U494 | ~new_R1207_U493;
  assign new_R1207_U496 = ~new_U3496 | ~new_R1207_U93;
  assign new_R1207_U497 = ~new_U3071 | ~new_R1207_U80;
  assign new_R1207_U498 = ~new_R1207_U330 | ~new_R1207_U107;
  assign new_R1207_U499 = ~new_R1207_U199 | ~new_R1207_U322;
  assign new_R1207_U500 = ~new_U3494 | ~new_R1207_U94;
  assign new_R1207_U501 = ~new_U3076 | ~new_R1207_U81;
  assign new_R1207_U502 = ~new_R1207_U201 | ~new_R1207_U331;
  assign new_R1207_U503 = ~new_R1207_U379 | ~new_R1207_U200;
  assign new_R1207_U504 = ~new_U3492 | ~new_R1207_U82;
  assign new_R1207_U505 = ~new_U3077 | ~new_R1207_U83;
  assign new_R1207_U506 = ~new_R1207_U169;
  assign new_R1207_U507 = ~new_R1207_U377 | ~new_R1207_U506;
  assign new_R1207_U508 = ~new_R1207_U169 | ~new_R1207_U202;
  assign new_R1207_U509 = ~new_U3490 | ~new_R1207_U90;
  assign new_R1207_U510 = ~new_U3069 | ~new_R1207_U84;
  assign new_R1207_U511 = ~new_R1207_U170;
  assign new_R1207_U512 = ~new_R1207_U375 | ~new_R1207_U511;
  assign new_R1207_U513 = ~new_R1207_U170 | ~new_R1207_U203;
  assign new_R1207_U514 = ~new_U3488 | ~new_R1207_U85;
  assign new_R1207_U515 = ~new_U3060 | ~new_R1207_U87;
  assign new_R1207_U516 = ~new_R1207_U515 | ~new_R1207_U514;
  assign new_R1207_U517 = ~new_U3486 | ~new_R1207_U86;
  assign new_R1207_U518 = ~new_U3059 | ~new_R1207_U88;
  assign new_R1207_U519 = ~new_R1207_U108 | ~new_R1207_U339;
  assign new_R1207_U520 = ~new_R1207_U204 | ~new_R1207_U373;
  assign new_R1165_U4 = new_R1165_U216 & new_R1165_U215;
  assign new_R1165_U5 = new_R1165_U226 & new_R1165_U225;
  assign new_R1165_U6 = new_R1165_U252 & new_R1165_U251;
  assign new_R1165_U7 = new_R1165_U268 & new_R1165_U267;
  assign new_R1165_U8 = new_R1165_U280 & new_R1165_U279;
  assign new_R1165_U9 = new_R1165_U298 & new_R1165_U297;
  assign new_R1165_U10 = new_R1165_U6 & new_R1165_U256;
  assign new_R1165_U11 = new_R1165_U5 & new_R1165_U223;
  assign new_R1165_U12 = new_R1165_U343 & new_R1165_U340;
  assign new_R1165_U13 = new_R1165_U334 & new_R1165_U331;
  assign new_R1165_U14 = new_R1165_U327 & new_R1165_U324;
  assign new_R1165_U15 = new_R1165_U318 & new_R1165_U315;
  assign new_R1165_U16 = new_R1165_U245 & new_R1165_U242;
  assign new_R1165_U17 = new_R1165_U238 & new_R1165_U235;
  assign new_R1165_U18 = ~new_U3208;
  assign new_R1165_U19 = ~new_U3170;
  assign new_R1165_U20 = ~new_U3172;
  assign new_R1165_U21 = ~new_U3172 | ~new_R1165_U64;
  assign new_R1165_U22 = ~new_U3171;
  assign new_R1165_U23 = ~new_U3173;
  assign new_R1165_U24 = ~new_U3173 | ~new_R1165_U66;
  assign new_R1165_U25 = ~new_U3174;
  assign new_R1165_U26 = ~new_U3176;
  assign new_R1165_U27 = ~new_U3176 | ~new_R1165_U68;
  assign new_R1165_U28 = ~new_U3175;
  assign new_R1165_U29 = ~new_U3177;
  assign new_R1165_U30 = ~new_U3178;
  assign new_R1165_U31 = ~new_U3178 | ~new_U3208;
  assign new_R1165_U32 = ~new_U3169;
  assign new_R1165_U33 = ~new_R1165_U360 | ~new_R1165_U230 | ~new_R1165_U229;
  assign new_R1165_U34 = ~new_R1165_U364 | ~new_R1165_U24;
  assign new_R1165_U35 = ~new_R1165_U357 | ~new_R1165_U358 | ~new_R1165_U213;
  assign new_R1165_U36 = ~new_U3162;
  assign new_R1165_U37 = ~new_U3162 | ~new_R1165_U72;
  assign new_R1165_U38 = ~new_U3161;
  assign new_R1165_U39 = ~new_U3166;
  assign new_R1165_U40 = ~new_U3167;
  assign new_R1165_U41 = ~new_U3167 | ~new_R1165_U76;
  assign new_R1165_U42 = ~new_U3165;
  assign new_R1165_U43 = ~new_U3168;
  assign new_R1165_U44 = ~new_U3168 | ~new_R1165_U77;
  assign new_R1165_U45 = ~new_U3164;
  assign new_R1165_U46 = ~new_U3163;
  assign new_R1165_U47 = ~new_U3160;
  assign new_R1165_U48 = ~new_U3158;
  assign new_R1165_U49 = ~new_U3159;
  assign new_R1165_U50 = ~new_U3159 | ~new_R1165_U81;
  assign new_R1165_U51 = ~new_U3157;
  assign new_R1165_U52 = ~new_U3156;
  assign new_R1165_U53 = ~new_U3155;
  assign new_R1165_U54 = ~new_U3153;
  assign new_R1165_U55 = ~new_U3154;
  assign new_R1165_U56 = ~new_U3154 | ~new_R1165_U86;
  assign new_R1165_U57 = ~new_U3152;
  assign new_R1165_U58 = ~new_U3151;
  assign new_R1165_U59 = ~new_R1165_U50 | ~new_R1165_U320;
  assign new_R1165_U60 = ~new_R1165_U265 | ~new_R1165_U264;
  assign new_R1165_U61 = ~new_R1165_U41 | ~new_R1165_U336;
  assign new_R1165_U62 = ~new_R1165_U377 | ~new_R1165_U376;
  assign new_R1165_U63 = ~new_R1165_U400 | ~new_R1165_U399;
  assign new_R1165_U64 = ~new_R1165_U409 | ~new_R1165_U408;
  assign new_R1165_U65 = ~new_R1165_U406 | ~new_R1165_U405;
  assign new_R1165_U66 = ~new_R1165_U403 | ~new_R1165_U402;
  assign new_R1165_U67 = ~new_R1165_U385 | ~new_R1165_U384;
  assign new_R1165_U68 = ~new_R1165_U397 | ~new_R1165_U396;
  assign new_R1165_U69 = ~new_R1165_U394 | ~new_R1165_U393;
  assign new_R1165_U70 = ~new_R1165_U388 | ~new_R1165_U387;
  assign new_R1165_U71 = ~new_R1165_U391 | ~new_R1165_U390;
  assign new_R1165_U72 = ~new_R1165_U473 | ~new_R1165_U472;
  assign new_R1165_U73 = ~new_R1165_U470 | ~new_R1165_U469;
  assign new_R1165_U74 = ~new_R1165_U458 | ~new_R1165_U457;
  assign new_R1165_U75 = ~new_R1165_U455 | ~new_R1165_U454;
  assign new_R1165_U76 = ~new_R1165_U452 | ~new_R1165_U451;
  assign new_R1165_U77 = ~new_R1165_U461 | ~new_R1165_U460;
  assign new_R1165_U78 = ~new_R1165_U464 | ~new_R1165_U463;
  assign new_R1165_U79 = ~new_R1165_U467 | ~new_R1165_U466;
  assign new_R1165_U80 = ~new_R1165_U476 | ~new_R1165_U475;
  assign new_R1165_U81 = ~new_R1165_U485 | ~new_R1165_U484;
  assign new_R1165_U82 = ~new_R1165_U479 | ~new_R1165_U478;
  assign new_R1165_U83 = ~new_R1165_U482 | ~new_R1165_U481;
  assign new_R1165_U84 = ~new_R1165_U488 | ~new_R1165_U487;
  assign new_R1165_U85 = ~new_R1165_U491 | ~new_R1165_U490;
  assign new_R1165_U86 = ~new_R1165_U500 | ~new_R1165_U499;
  assign new_R1165_U87 = ~new_R1165_U494 | ~new_R1165_U493;
  assign new_R1165_U88 = ~new_R1165_U497 | ~new_R1165_U496;
  assign new_R1165_U89 = ~new_R1165_U449 | ~new_R1165_U448;
  assign new_R1165_U90 = ~new_R1165_U506 | ~new_R1165_U505;
  assign new_R1165_U91 = ~new_R1165_U613 | ~new_R1165_U612;
  assign new_R1165_U92 = ~new_R1165_U412 | ~new_R1165_U411;
  assign new_R1165_U93 = ~new_R1165_U419 | ~new_R1165_U418;
  assign new_R1165_U94 = ~new_R1165_U426 | ~new_R1165_U425;
  assign new_R1165_U95 = ~new_R1165_U433 | ~new_R1165_U432;
  assign new_R1165_U96 = ~new_R1165_U440 | ~new_R1165_U439;
  assign new_R1165_U97 = ~new_R1165_U447 | ~new_R1165_U446;
  assign new_R1165_U98 = ~new_R1165_U509 | ~new_R1165_U508;
  assign new_R1165_U99 = ~new_R1165_U516 | ~new_R1165_U515;
  assign new_R1165_U100 = ~new_R1165_U523 | ~new_R1165_U522;
  assign new_R1165_U101 = ~new_R1165_U528 | ~new_R1165_U527;
  assign new_R1165_U102 = ~new_R1165_U535 | ~new_R1165_U534;
  assign new_R1165_U103 = ~new_R1165_U542 | ~new_R1165_U541;
  assign new_R1165_U104 = ~new_R1165_U549 | ~new_R1165_U548;
  assign new_R1165_U105 = ~new_R1165_U556 | ~new_R1165_U555;
  assign new_R1165_U106 = ~new_R1165_U561 | ~new_R1165_U560;
  assign new_R1165_U107 = ~new_R1165_U568 | ~new_R1165_U567;
  assign new_R1165_U108 = ~new_R1165_U575 | ~new_R1165_U574;
  assign new_R1165_U109 = ~new_R1165_U582 | ~new_R1165_U581;
  assign new_R1165_U110 = ~new_R1165_U589 | ~new_R1165_U588;
  assign new_R1165_U111 = ~new_R1165_U596 | ~new_R1165_U595;
  assign new_R1165_U112 = ~new_R1165_U601 | ~new_R1165_U600;
  assign new_R1165_U113 = ~new_R1165_U608 | ~new_R1165_U607;
  assign new_R1165_U114 = new_R1165_U71 & new_R1165_U209;
  assign new_R1165_U115 = new_R1165_U219 & new_R1165_U218;
  assign new_R1165_U116 = new_R1165_U11 & new_R1165_U231;
  assign new_R1165_U117 = new_R1165_U362 & new_R1165_U232;
  assign new_R1165_U118 = new_R1165_U21 & new_R1165_U421 & new_R1165_U420;
  assign new_R1165_U119 = new_R1165_U237 & new_R1165_U5;
  assign new_R1165_U120 = new_R1165_U27 & new_R1165_U442 & new_R1165_U441;
  assign new_R1165_U121 = new_R1165_U244 & new_R1165_U4;
  assign new_R1165_U122 = new_R1165_U254 & new_R1165_U203;
  assign new_R1165_U123 = new_R1165_U249 & new_R1165_U10;
  assign new_R1165_U124 = new_R1165_U363 & new_R1165_U258;
  assign new_R1165_U125 = new_R1165_U272 & new_R1165_U271;
  assign new_R1165_U126 = new_R1165_U284 & new_R1165_U8;
  assign new_R1165_U127 = new_R1165_U282 & new_R1165_U204;
  assign new_R1165_U128 = new_R1165_U302 & new_R1165_U9;
  assign new_R1165_U129 = new_R1165_U300 & new_R1165_U205;
  assign new_R1165_U130 = new_R1165_U305 & new_R1165_U308;
  assign new_R1165_U131 = ~new_R1165_U503 | ~new_R1165_U502;
  assign new_R1165_U132 = new_R1165_U205 & new_R1165_U518 & new_R1165_U517;
  assign new_R1165_U133 = new_R1165_U56 & new_R1165_U205;
  assign new_R1165_U134 = new_R1165_U317 & new_R1165_U9;
  assign new_R1165_U135 = new_R1165_U204 & new_R1165_U544 & new_R1165_U543;
  assign new_R1165_U136 = new_R1165_U326 & new_R1165_U8;
  assign new_R1165_U137 = new_R1165_U37 & new_R1165_U570 & new_R1165_U569;
  assign new_R1165_U138 = new_R1165_U333 & new_R1165_U7;
  assign new_R1165_U139 = new_R1165_U203 & new_R1165_U591 & new_R1165_U590;
  assign new_R1165_U140 = new_R1165_U342 & new_R1165_U6;
  assign new_R1165_U141 = ~new_R1165_U610 | ~new_R1165_U609;
  assign new_R1165_U142 = ~new_U3198;
  assign new_R1165_U143 = new_R1165_U380 & new_R1165_U379;
  assign new_R1165_U144 = ~new_U3203;
  assign new_R1165_U145 = ~new_U3206;
  assign new_R1165_U146 = ~new_U3207;
  assign new_R1165_U147 = ~new_U3204;
  assign new_R1165_U148 = ~new_U3205;
  assign new_R1165_U149 = ~new_U3199;
  assign new_R1165_U150 = ~new_U3202;
  assign new_R1165_U151 = ~new_U3200;
  assign new_R1165_U152 = ~new_U3201;
  assign new_R1165_U153 = ~new_R1165_U117 | ~new_R1165_U368;
  assign new_R1165_U154 = new_R1165_U414 & new_R1165_U413;
  assign new_R1165_U155 = ~new_R1165_U361 | ~new_R1165_U366;
  assign new_R1165_U156 = new_R1165_U428 & new_R1165_U427;
  assign new_R1165_U157 = ~new_R1165_U370 | ~new_R1165_U354;
  assign new_R1165_U158 = new_R1165_U435 & new_R1165_U434;
  assign new_R1165_U159 = ~new_R1165_U115 | ~new_R1165_U220;
  assign new_R1165_U160 = ~new_U3180;
  assign new_R1165_U161 = ~new_U3196;
  assign new_R1165_U162 = ~new_U3194;
  assign new_R1165_U163 = ~new_U3195;
  assign new_R1165_U164 = ~new_U3197;
  assign new_R1165_U165 = ~new_U3193;
  assign new_R1165_U166 = ~new_U3192;
  assign new_R1165_U167 = ~new_U3190;
  assign new_R1165_U168 = ~new_U3191;
  assign new_R1165_U169 = ~new_U3189;
  assign new_R1165_U170 = ~new_U3186;
  assign new_R1165_U171 = ~new_U3187;
  assign new_R1165_U172 = ~new_U3188;
  assign new_R1165_U173 = ~new_U3185;
  assign new_R1165_U174 = ~new_U3184;
  assign new_R1165_U175 = ~new_U3181;
  assign new_R1165_U176 = ~new_U3182;
  assign new_R1165_U177 = ~new_U3183;
  assign new_R1165_U178 = ~new_U3150;
  assign new_R1165_U179 = ~new_U3179;
  assign new_R1165_U180 = new_R1165_U511 & new_R1165_U510;
  assign new_R1165_U181 = ~new_R1165_U305 | ~new_R1165_U304;
  assign new_R1165_U182 = ~new_R1165_U56 | ~new_R1165_U311;
  assign new_R1165_U183 = ~new_R1165_U295 | ~new_R1165_U294;
  assign new_R1165_U184 = new_R1165_U530 & new_R1165_U529;
  assign new_R1165_U185 = ~new_R1165_U291 | ~new_R1165_U290;
  assign new_R1165_U186 = new_R1165_U537 & new_R1165_U536;
  assign new_R1165_U187 = ~new_R1165_U287 | ~new_R1165_U286;
  assign new_R1165_U188 = new_R1165_U551 & new_R1165_U550;
  assign new_R1165_U189 = ~new_R1165_U31 | ~new_R1165_U210;
  assign new_R1165_U190 = ~new_R1165_U277 | ~new_R1165_U276;
  assign new_R1165_U191 = new_R1165_U563 & new_R1165_U562;
  assign new_R1165_U192 = ~new_R1165_U125 | ~new_R1165_U273;
  assign new_R1165_U193 = new_R1165_U577 & new_R1165_U576;
  assign new_R1165_U194 = ~new_R1165_U261 | ~new_R1165_U260;
  assign new_R1165_U195 = new_R1165_U584 & new_R1165_U583;
  assign new_R1165_U196 = ~new_R1165_U124 | ~new_R1165_U374;
  assign new_R1165_U197 = ~new_R1165_U372 | ~new_R1165_U44;
  assign new_R1165_U198 = new_R1165_U603 & new_R1165_U602;
  assign new_R1165_U199 = ~new_R1165_U355 | ~new_R1165_U247 | ~new_R1165_U201;
  assign new_R1165_U200 = ~new_R1165_U310 | ~new_R1165_U181;
  assign new_R1165_U201 = ~new_R1165_U62 | ~new_R1165_U153;
  assign new_R1165_U202 = ~new_R1165_U27;
  assign new_R1165_U203 = ~new_U3166 | ~new_R1165_U74;
  assign new_R1165_U204 = ~new_U3158 | ~new_R1165_U83;
  assign new_R1165_U205 = ~new_U3153 | ~new_R1165_U88;
  assign new_R1165_U206 = ~new_R1165_U41;
  assign new_R1165_U207 = ~new_R1165_U50;
  assign new_R1165_U208 = ~new_R1165_U56;
  assign new_R1165_U209 = new_U3208 | new_U3178;
  assign new_R1165_U210 = ~new_R1165_U71 | ~new_R1165_U209;
  assign new_R1165_U211 = ~new_R1165_U31;
  assign new_R1165_U212 = ~new_R1165_U189;
  assign new_R1165_U213 = ~new_U3177 | ~new_R1165_U70;
  assign new_R1165_U214 = ~new_R1165_U35;
  assign new_R1165_U215 = ~new_R1165_U395 | ~new_R1165_U28;
  assign new_R1165_U216 = ~new_R1165_U398 | ~new_R1165_U26;
  assign new_R1165_U217 = ~new_R1165_U28 | ~new_R1165_U27;
  assign new_R1165_U218 = ~new_R1165_U69 | ~new_R1165_U217;
  assign new_R1165_U219 = ~new_U3175 | ~new_R1165_U202;
  assign new_R1165_U220 = ~new_R1165_U4 | ~new_R1165_U35;
  assign new_R1165_U221 = ~new_R1165_U159;
  assign new_R1165_U222 = ~new_R1165_U386 | ~new_R1165_U25;
  assign new_R1165_U223 = ~new_R1165_U404 | ~new_R1165_U23;
  assign new_R1165_U224 = ~new_R1165_U24;
  assign new_R1165_U225 = ~new_R1165_U407 | ~new_R1165_U22;
  assign new_R1165_U226 = ~new_R1165_U410 | ~new_R1165_U20;
  assign new_R1165_U227 = ~new_R1165_U21;
  assign new_R1165_U228 = ~new_R1165_U22 | ~new_R1165_U21;
  assign new_R1165_U229 = ~new_R1165_U65 | ~new_R1165_U228;
  assign new_R1165_U230 = ~new_U3171 | ~new_R1165_U227;
  assign new_R1165_U231 = ~new_R1165_U401 | ~new_R1165_U19;
  assign new_R1165_U232 = ~new_U3170 | ~new_R1165_U63;
  assign new_R1165_U233 = ~new_R1165_U410 | ~new_R1165_U20;
  assign new_R1165_U234 = ~new_R1165_U233 | ~new_R1165_U34;
  assign new_R1165_U235 = ~new_R1165_U118 | ~new_R1165_U234;
  assign new_R1165_U236 = ~new_R1165_U365 | ~new_R1165_U21;
  assign new_R1165_U237 = ~new_U3171 | ~new_R1165_U65;
  assign new_R1165_U238 = ~new_R1165_U119 | ~new_R1165_U236;
  assign new_R1165_U239 = ~new_R1165_U410 | ~new_R1165_U20;
  assign new_R1165_U240 = ~new_R1165_U398 | ~new_R1165_U26;
  assign new_R1165_U241 = ~new_R1165_U240 | ~new_R1165_U35;
  assign new_R1165_U242 = ~new_R1165_U120 | ~new_R1165_U241;
  assign new_R1165_U243 = ~new_R1165_U214 | ~new_R1165_U27;
  assign new_R1165_U244 = ~new_U3175 | ~new_R1165_U69;
  assign new_R1165_U245 = ~new_R1165_U121 | ~new_R1165_U243;
  assign new_R1165_U246 = ~new_R1165_U398 | ~new_R1165_U26;
  assign new_R1165_U247 = ~new_U3169 | ~new_R1165_U153;
  assign new_R1165_U248 = ~new_R1165_U199;
  assign new_R1165_U249 = ~new_R1165_U462 | ~new_R1165_U43;
  assign new_R1165_U250 = ~new_R1165_U44;
  assign new_R1165_U251 = ~new_R1165_U456 | ~new_R1165_U42;
  assign new_R1165_U252 = ~new_R1165_U459 | ~new_R1165_U39;
  assign new_R1165_U253 = ~new_R1165_U206 | ~new_R1165_U6;
  assign new_R1165_U254 = ~new_U3165 | ~new_R1165_U75;
  assign new_R1165_U255 = ~new_R1165_U122 | ~new_R1165_U253;
  assign new_R1165_U256 = ~new_R1165_U453 | ~new_R1165_U40;
  assign new_R1165_U257 = ~new_R1165_U456 | ~new_R1165_U42;
  assign new_R1165_U258 = ~new_R1165_U257 | ~new_R1165_U255;
  assign new_R1165_U259 = ~new_R1165_U465 | ~new_R1165_U45;
  assign new_R1165_U260 = ~new_R1165_U259 | ~new_R1165_U196;
  assign new_R1165_U261 = ~new_U3164 | ~new_R1165_U78;
  assign new_R1165_U262 = ~new_R1165_U194;
  assign new_R1165_U263 = ~new_R1165_U468 | ~new_R1165_U46;
  assign new_R1165_U264 = ~new_R1165_U263 | ~new_R1165_U194;
  assign new_R1165_U265 = ~new_U3163 | ~new_R1165_U79;
  assign new_R1165_U266 = ~new_R1165_U60;
  assign new_R1165_U267 = ~new_R1165_U471 | ~new_R1165_U38;
  assign new_R1165_U268 = ~new_R1165_U474 | ~new_R1165_U36;
  assign new_R1165_U269 = ~new_R1165_U37;
  assign new_R1165_U270 = ~new_R1165_U38 | ~new_R1165_U37;
  assign new_R1165_U271 = ~new_R1165_U73 | ~new_R1165_U270;
  assign new_R1165_U272 = ~new_U3161 | ~new_R1165_U269;
  assign new_R1165_U273 = ~new_R1165_U7 | ~new_R1165_U60;
  assign new_R1165_U274 = ~new_R1165_U192;
  assign new_R1165_U275 = ~new_R1165_U477 | ~new_R1165_U47;
  assign new_R1165_U276 = ~new_R1165_U275 | ~new_R1165_U192;
  assign new_R1165_U277 = ~new_U3160 | ~new_R1165_U80;
  assign new_R1165_U278 = ~new_R1165_U190;
  assign new_R1165_U279 = ~new_R1165_U480 | ~new_R1165_U51;
  assign new_R1165_U280 = ~new_R1165_U483 | ~new_R1165_U48;
  assign new_R1165_U281 = ~new_R1165_U207 | ~new_R1165_U8;
  assign new_R1165_U282 = ~new_U3157 | ~new_R1165_U82;
  assign new_R1165_U283 = ~new_R1165_U127 | ~new_R1165_U281;
  assign new_R1165_U284 = ~new_R1165_U486 | ~new_R1165_U49;
  assign new_R1165_U285 = ~new_R1165_U480 | ~new_R1165_U51;
  assign new_R1165_U286 = ~new_R1165_U126 | ~new_R1165_U190;
  assign new_R1165_U287 = ~new_R1165_U285 | ~new_R1165_U283;
  assign new_R1165_U288 = ~new_R1165_U187;
  assign new_R1165_U289 = ~new_R1165_U489 | ~new_R1165_U52;
  assign new_R1165_U290 = ~new_R1165_U289 | ~new_R1165_U187;
  assign new_R1165_U291 = ~new_U3156 | ~new_R1165_U84;
  assign new_R1165_U292 = ~new_R1165_U185;
  assign new_R1165_U293 = ~new_R1165_U492 | ~new_R1165_U53;
  assign new_R1165_U294 = ~new_R1165_U293 | ~new_R1165_U185;
  assign new_R1165_U295 = ~new_U3155 | ~new_R1165_U85;
  assign new_R1165_U296 = ~new_R1165_U183;
  assign new_R1165_U297 = ~new_R1165_U495 | ~new_R1165_U57;
  assign new_R1165_U298 = ~new_R1165_U498 | ~new_R1165_U54;
  assign new_R1165_U299 = ~new_R1165_U208 | ~new_R1165_U9;
  assign new_R1165_U300 = ~new_U3152 | ~new_R1165_U87;
  assign new_R1165_U301 = ~new_R1165_U129 | ~new_R1165_U299;
  assign new_R1165_U302 = ~new_R1165_U501 | ~new_R1165_U55;
  assign new_R1165_U303 = ~new_R1165_U495 | ~new_R1165_U57;
  assign new_R1165_U304 = ~new_R1165_U128 | ~new_R1165_U183;
  assign new_R1165_U305 = ~new_R1165_U303 | ~new_R1165_U301;
  assign new_R1165_U306 = ~new_R1165_U181;
  assign new_R1165_U307 = ~new_R1165_U450 | ~new_R1165_U58;
  assign new_R1165_U308 = ~new_U3151 | ~new_R1165_U89;
  assign new_R1165_U309 = ~new_U3151 | ~new_R1165_U89;
  assign new_R1165_U310 = ~new_R1165_U450 | ~new_R1165_U58;
  assign new_R1165_U311 = ~new_R1165_U302 | ~new_R1165_U183;
  assign new_R1165_U312 = ~new_R1165_U182;
  assign new_R1165_U313 = ~new_R1165_U498 | ~new_R1165_U54;
  assign new_R1165_U314 = ~new_R1165_U313 | ~new_R1165_U182;
  assign new_R1165_U315 = ~new_R1165_U132 | ~new_R1165_U314;
  assign new_R1165_U316 = ~new_R1165_U133 | ~new_R1165_U311;
  assign new_R1165_U317 = ~new_U3152 | ~new_R1165_U87;
  assign new_R1165_U318 = ~new_R1165_U134 | ~new_R1165_U316;
  assign new_R1165_U319 = ~new_R1165_U498 | ~new_R1165_U54;
  assign new_R1165_U320 = ~new_R1165_U284 | ~new_R1165_U190;
  assign new_R1165_U321 = ~new_R1165_U59;
  assign new_R1165_U322 = ~new_R1165_U483 | ~new_R1165_U48;
  assign new_R1165_U323 = ~new_R1165_U322 | ~new_R1165_U59;
  assign new_R1165_U324 = ~new_R1165_U135 | ~new_R1165_U323;
  assign new_R1165_U325 = ~new_R1165_U321 | ~new_R1165_U204;
  assign new_R1165_U326 = ~new_U3157 | ~new_R1165_U82;
  assign new_R1165_U327 = ~new_R1165_U136 | ~new_R1165_U325;
  assign new_R1165_U328 = ~new_R1165_U483 | ~new_R1165_U48;
  assign new_R1165_U329 = ~new_R1165_U474 | ~new_R1165_U36;
  assign new_R1165_U330 = ~new_R1165_U329 | ~new_R1165_U60;
  assign new_R1165_U331 = ~new_R1165_U137 | ~new_R1165_U330;
  assign new_R1165_U332 = ~new_R1165_U266 | ~new_R1165_U37;
  assign new_R1165_U333 = ~new_U3161 | ~new_R1165_U73;
  assign new_R1165_U334 = ~new_R1165_U138 | ~new_R1165_U332;
  assign new_R1165_U335 = ~new_R1165_U474 | ~new_R1165_U36;
  assign new_R1165_U336 = ~new_R1165_U256 | ~new_R1165_U197;
  assign new_R1165_U337 = ~new_R1165_U61;
  assign new_R1165_U338 = ~new_R1165_U459 | ~new_R1165_U39;
  assign new_R1165_U339 = ~new_R1165_U338 | ~new_R1165_U61;
  assign new_R1165_U340 = ~new_R1165_U139 | ~new_R1165_U339;
  assign new_R1165_U341 = ~new_R1165_U337 | ~new_R1165_U203;
  assign new_R1165_U342 = ~new_U3165 | ~new_R1165_U75;
  assign new_R1165_U343 = ~new_R1165_U140 | ~new_R1165_U341;
  assign new_R1165_U344 = ~new_R1165_U459 | ~new_R1165_U39;
  assign new_R1165_U345 = ~new_R1165_U239 | ~new_R1165_U21;
  assign new_R1165_U346 = ~new_R1165_U246 | ~new_R1165_U27;
  assign new_R1165_U347 = ~new_R1165_U319 | ~new_R1165_U205;
  assign new_R1165_U348 = ~new_R1165_U302 | ~new_R1165_U56;
  assign new_R1165_U349 = ~new_R1165_U328 | ~new_R1165_U204;
  assign new_R1165_U350 = ~new_R1165_U284 | ~new_R1165_U50;
  assign new_R1165_U351 = ~new_R1165_U335 | ~new_R1165_U37;
  assign new_R1165_U352 = ~new_R1165_U344 | ~new_R1165_U203;
  assign new_R1165_U353 = ~new_R1165_U256 | ~new_R1165_U41;
  assign new_R1165_U354 = ~new_U3174 | ~new_R1165_U67;
  assign new_R1165_U355 = ~new_U3169 | ~new_R1165_U62;
  assign new_R1165_U356 = ~new_R1165_U130 | ~new_R1165_U304;
  assign new_R1165_U357 = ~new_R1165_U114 | ~new_R1165_U359;
  assign new_R1165_U358 = ~new_R1165_U211 | ~new_R1165_U359;
  assign new_R1165_U359 = ~new_R1165_U389 | ~new_R1165_U29;
  assign new_R1165_U360 = ~new_R1165_U224 | ~new_R1165_U5;
  assign new_R1165_U361 = ~new_R1165_U33;
  assign new_R1165_U362 = ~new_R1165_U33 | ~new_R1165_U231;
  assign new_R1165_U363 = ~new_R1165_U250 | ~new_R1165_U10;
  assign new_R1165_U364 = ~new_R1165_U223 | ~new_R1165_U157;
  assign new_R1165_U365 = ~new_R1165_U34;
  assign new_R1165_U366 = ~new_R1165_U11 | ~new_R1165_U157;
  assign new_R1165_U367 = ~new_R1165_U155;
  assign new_R1165_U368 = ~new_R1165_U116 | ~new_R1165_U157;
  assign new_R1165_U369 = ~new_R1165_U153;
  assign new_R1165_U370 = ~new_R1165_U222 | ~new_R1165_U159;
  assign new_R1165_U371 = ~new_R1165_U157;
  assign new_R1165_U372 = ~new_R1165_U249 | ~new_R1165_U199;
  assign new_R1165_U373 = ~new_R1165_U197;
  assign new_R1165_U374 = ~new_R1165_U123 | ~new_R1165_U199;
  assign new_R1165_U375 = ~new_R1165_U196;
  assign new_R1165_U376 = ~new_U3208 | ~new_R1165_U142;
  assign new_R1165_U377 = ~new_U3198 | ~new_R1165_U18;
  assign new_R1165_U378 = ~new_R1165_U62;
  assign new_R1165_U379 = ~new_R1165_U378 | ~new_U3169;
  assign new_R1165_U380 = ~new_R1165_U62 | ~new_R1165_U32;
  assign new_R1165_U381 = ~new_R1165_U378 | ~new_U3169;
  assign new_R1165_U382 = ~new_R1165_U62 | ~new_R1165_U32;
  assign new_R1165_U383 = ~new_R1165_U382 | ~new_R1165_U381;
  assign new_R1165_U384 = ~new_U3208 | ~new_R1165_U144;
  assign new_R1165_U385 = ~new_U3203 | ~new_R1165_U18;
  assign new_R1165_U386 = ~new_R1165_U67;
  assign new_R1165_U387 = ~new_U3208 | ~new_R1165_U145;
  assign new_R1165_U388 = ~new_U3206 | ~new_R1165_U18;
  assign new_R1165_U389 = ~new_R1165_U70;
  assign new_R1165_U390 = ~new_U3208 | ~new_R1165_U146;
  assign new_R1165_U391 = ~new_U3207 | ~new_R1165_U18;
  assign new_R1165_U392 = ~new_R1165_U71;
  assign new_R1165_U393 = ~new_U3208 | ~new_R1165_U147;
  assign new_R1165_U394 = ~new_U3204 | ~new_R1165_U18;
  assign new_R1165_U395 = ~new_R1165_U69;
  assign new_R1165_U396 = ~new_U3208 | ~new_R1165_U148;
  assign new_R1165_U397 = ~new_U3205 | ~new_R1165_U18;
  assign new_R1165_U398 = ~new_R1165_U68;
  assign new_R1165_U399 = ~new_U3208 | ~new_R1165_U149;
  assign new_R1165_U400 = ~new_U3199 | ~new_R1165_U18;
  assign new_R1165_U401 = ~new_R1165_U63;
  assign new_R1165_U402 = ~new_U3208 | ~new_R1165_U150;
  assign new_R1165_U403 = ~new_U3202 | ~new_R1165_U18;
  assign new_R1165_U404 = ~new_R1165_U66;
  assign new_R1165_U405 = ~new_U3208 | ~new_R1165_U151;
  assign new_R1165_U406 = ~new_U3200 | ~new_R1165_U18;
  assign new_R1165_U407 = ~new_R1165_U65;
  assign new_R1165_U408 = ~new_U3208 | ~new_R1165_U152;
  assign new_R1165_U409 = ~new_U3201 | ~new_R1165_U18;
  assign new_R1165_U410 = ~new_R1165_U64;
  assign new_R1165_U411 = ~new_R1165_U143 | ~new_R1165_U153;
  assign new_R1165_U412 = ~new_R1165_U369 | ~new_R1165_U383;
  assign new_R1165_U413 = ~new_R1165_U401 | ~new_U3170;
  assign new_R1165_U414 = ~new_R1165_U63 | ~new_R1165_U19;
  assign new_R1165_U415 = ~new_R1165_U401 | ~new_U3170;
  assign new_R1165_U416 = ~new_R1165_U63 | ~new_R1165_U19;
  assign new_R1165_U417 = ~new_R1165_U416 | ~new_R1165_U415;
  assign new_R1165_U418 = ~new_R1165_U154 | ~new_R1165_U155;
  assign new_R1165_U419 = ~new_R1165_U367 | ~new_R1165_U417;
  assign new_R1165_U420 = ~new_R1165_U407 | ~new_U3171;
  assign new_R1165_U421 = ~new_R1165_U65 | ~new_R1165_U22;
  assign new_R1165_U422 = ~new_R1165_U410 | ~new_U3172;
  assign new_R1165_U423 = ~new_R1165_U64 | ~new_R1165_U20;
  assign new_R1165_U424 = ~new_R1165_U423 | ~new_R1165_U422;
  assign new_R1165_U425 = ~new_R1165_U34 | ~new_R1165_U345;
  assign new_R1165_U426 = ~new_R1165_U424 | ~new_R1165_U365;
  assign new_R1165_U427 = ~new_R1165_U404 | ~new_U3173;
  assign new_R1165_U428 = ~new_R1165_U66 | ~new_R1165_U23;
  assign new_R1165_U429 = ~new_R1165_U404 | ~new_U3173;
  assign new_R1165_U430 = ~new_R1165_U66 | ~new_R1165_U23;
  assign new_R1165_U431 = ~new_R1165_U430 | ~new_R1165_U429;
  assign new_R1165_U432 = ~new_R1165_U156 | ~new_R1165_U157;
  assign new_R1165_U433 = ~new_R1165_U371 | ~new_R1165_U431;
  assign new_R1165_U434 = ~new_R1165_U386 | ~new_U3174;
  assign new_R1165_U435 = ~new_R1165_U67 | ~new_R1165_U25;
  assign new_R1165_U436 = ~new_R1165_U386 | ~new_U3174;
  assign new_R1165_U437 = ~new_R1165_U67 | ~new_R1165_U25;
  assign new_R1165_U438 = ~new_R1165_U437 | ~new_R1165_U436;
  assign new_R1165_U439 = ~new_R1165_U158 | ~new_R1165_U159;
  assign new_R1165_U440 = ~new_R1165_U221 | ~new_R1165_U438;
  assign new_R1165_U441 = ~new_R1165_U395 | ~new_U3175;
  assign new_R1165_U442 = ~new_R1165_U69 | ~new_R1165_U28;
  assign new_R1165_U443 = ~new_R1165_U398 | ~new_U3176;
  assign new_R1165_U444 = ~new_R1165_U68 | ~new_R1165_U26;
  assign new_R1165_U445 = ~new_R1165_U444 | ~new_R1165_U443;
  assign new_R1165_U446 = ~new_R1165_U346 | ~new_R1165_U35;
  assign new_R1165_U447 = ~new_R1165_U445 | ~new_R1165_U214;
  assign new_R1165_U448 = ~new_U3208 | ~new_R1165_U160;
  assign new_R1165_U449 = ~new_U3180 | ~new_R1165_U18;
  assign new_R1165_U450 = ~new_R1165_U89;
  assign new_R1165_U451 = ~new_U3208 | ~new_R1165_U161;
  assign new_R1165_U452 = ~new_U3196 | ~new_R1165_U18;
  assign new_R1165_U453 = ~new_R1165_U76;
  assign new_R1165_U454 = ~new_U3208 | ~new_R1165_U162;
  assign new_R1165_U455 = ~new_U3194 | ~new_R1165_U18;
  assign new_R1165_U456 = ~new_R1165_U75;
  assign new_R1165_U457 = ~new_U3208 | ~new_R1165_U163;
  assign new_R1165_U458 = ~new_U3195 | ~new_R1165_U18;
  assign new_R1165_U459 = ~new_R1165_U74;
  assign new_R1165_U460 = ~new_U3208 | ~new_R1165_U164;
  assign new_R1165_U461 = ~new_U3197 | ~new_R1165_U18;
  assign new_R1165_U462 = ~new_R1165_U77;
  assign new_R1165_U463 = ~new_U3208 | ~new_R1165_U165;
  assign new_R1165_U464 = ~new_U3193 | ~new_R1165_U18;
  assign new_R1165_U465 = ~new_R1165_U78;
  assign new_R1165_U466 = ~new_U3208 | ~new_R1165_U166;
  assign new_R1165_U467 = ~new_U3192 | ~new_R1165_U18;
  assign new_R1165_U468 = ~new_R1165_U79;
  assign new_R1165_U469 = ~new_U3208 | ~new_R1165_U167;
  assign new_R1165_U470 = ~new_U3190 | ~new_R1165_U18;
  assign new_R1165_U471 = ~new_R1165_U73;
  assign new_R1165_U472 = ~new_U3208 | ~new_R1165_U168;
  assign new_R1165_U473 = ~new_U3191 | ~new_R1165_U18;
  assign new_R1165_U474 = ~new_R1165_U72;
  assign new_R1165_U475 = ~new_U3208 | ~new_R1165_U169;
  assign new_R1165_U476 = ~new_U3189 | ~new_R1165_U18;
  assign new_R1165_U477 = ~new_R1165_U80;
  assign new_R1165_U478 = ~new_U3208 | ~new_R1165_U170;
  assign new_R1165_U479 = ~new_U3186 | ~new_R1165_U18;
  assign new_R1165_U480 = ~new_R1165_U82;
  assign new_R1165_U481 = ~new_U3208 | ~new_R1165_U171;
  assign new_R1165_U482 = ~new_U3187 | ~new_R1165_U18;
  assign new_R1165_U483 = ~new_R1165_U83;
  assign new_R1165_U484 = ~new_U3208 | ~new_R1165_U172;
  assign new_R1165_U485 = ~new_U3188 | ~new_R1165_U18;
  assign new_R1165_U486 = ~new_R1165_U81;
  assign new_R1165_U487 = ~new_U3208 | ~new_R1165_U173;
  assign new_R1165_U488 = ~new_U3185 | ~new_R1165_U18;
  assign new_R1165_U489 = ~new_R1165_U84;
  assign new_R1165_U490 = ~new_U3208 | ~new_R1165_U174;
  assign new_R1165_U491 = ~new_U3184 | ~new_R1165_U18;
  assign new_R1165_U492 = ~new_R1165_U85;
  assign new_R1165_U493 = ~new_U3208 | ~new_R1165_U175;
  assign new_R1165_U494 = ~new_U3181 | ~new_R1165_U18;
  assign new_R1165_U495 = ~new_R1165_U87;
  assign new_R1165_U496 = ~new_U3208 | ~new_R1165_U176;
  assign new_R1165_U497 = ~new_U3182 | ~new_R1165_U18;
  assign new_R1165_U498 = ~new_R1165_U88;
  assign new_R1165_U499 = ~new_U3208 | ~new_R1165_U177;
  assign new_R1165_U500 = ~new_U3183 | ~new_R1165_U18;
  assign new_R1165_U501 = ~new_R1165_U86;
  assign new_R1165_U502 = ~new_U3208 | ~new_R1165_U178;
  assign new_R1165_U503 = ~new_U3150 | ~new_R1165_U18;
  assign new_R1165_U504 = ~new_R1165_U131;
  assign new_R1165_U505 = ~new_U3179 | ~new_R1165_U504;
  assign new_R1165_U506 = ~new_R1165_U131 | ~new_R1165_U179;
  assign new_R1165_U507 = ~new_R1165_U90;
  assign new_R1165_U508 = ~new_R1165_U507 | ~new_R1165_U356 | ~new_R1165_U307;
  assign new_R1165_U509 = ~new_R1165_U90 | ~new_R1165_U309 | ~new_R1165_U200;
  assign new_R1165_U510 = ~new_R1165_U450 | ~new_U3151;
  assign new_R1165_U511 = ~new_R1165_U89 | ~new_R1165_U58;
  assign new_R1165_U512 = ~new_R1165_U450 | ~new_U3151;
  assign new_R1165_U513 = ~new_R1165_U89 | ~new_R1165_U58;
  assign new_R1165_U514 = ~new_R1165_U513 | ~new_R1165_U512;
  assign new_R1165_U515 = ~new_R1165_U180 | ~new_R1165_U181;
  assign new_R1165_U516 = ~new_R1165_U306 | ~new_R1165_U514;
  assign new_R1165_U517 = ~new_R1165_U495 | ~new_U3152;
  assign new_R1165_U518 = ~new_R1165_U87 | ~new_R1165_U57;
  assign new_R1165_U519 = ~new_R1165_U498 | ~new_U3153;
  assign new_R1165_U520 = ~new_R1165_U88 | ~new_R1165_U54;
  assign new_R1165_U521 = ~new_R1165_U520 | ~new_R1165_U519;
  assign new_R1165_U522 = ~new_R1165_U347 | ~new_R1165_U182;
  assign new_R1165_U523 = ~new_R1165_U312 | ~new_R1165_U521;
  assign new_R1165_U524 = ~new_R1165_U501 | ~new_U3154;
  assign new_R1165_U525 = ~new_R1165_U86 | ~new_R1165_U55;
  assign new_R1165_U526 = ~new_R1165_U525 | ~new_R1165_U524;
  assign new_R1165_U527 = ~new_R1165_U348 | ~new_R1165_U183;
  assign new_R1165_U528 = ~new_R1165_U296 | ~new_R1165_U526;
  assign new_R1165_U529 = ~new_R1165_U492 | ~new_U3155;
  assign new_R1165_U530 = ~new_R1165_U85 | ~new_R1165_U53;
  assign new_R1165_U531 = ~new_R1165_U492 | ~new_U3155;
  assign new_R1165_U532 = ~new_R1165_U85 | ~new_R1165_U53;
  assign new_R1165_U533 = ~new_R1165_U532 | ~new_R1165_U531;
  assign new_R1165_U534 = ~new_R1165_U184 | ~new_R1165_U185;
  assign new_R1165_U535 = ~new_R1165_U292 | ~new_R1165_U533;
  assign new_R1165_U536 = ~new_R1165_U489 | ~new_U3156;
  assign new_R1165_U537 = ~new_R1165_U84 | ~new_R1165_U52;
  assign new_R1165_U538 = ~new_R1165_U489 | ~new_U3156;
  assign new_R1165_U539 = ~new_R1165_U84 | ~new_R1165_U52;
  assign new_R1165_U540 = ~new_R1165_U539 | ~new_R1165_U538;
  assign new_R1165_U541 = ~new_R1165_U186 | ~new_R1165_U187;
  assign new_R1165_U542 = ~new_R1165_U288 | ~new_R1165_U540;
  assign new_R1165_U543 = ~new_R1165_U480 | ~new_U3157;
  assign new_R1165_U544 = ~new_R1165_U82 | ~new_R1165_U51;
  assign new_R1165_U545 = ~new_R1165_U483 | ~new_U3158;
  assign new_R1165_U546 = ~new_R1165_U83 | ~new_R1165_U48;
  assign new_R1165_U547 = ~new_R1165_U546 | ~new_R1165_U545;
  assign new_R1165_U548 = ~new_R1165_U349 | ~new_R1165_U59;
  assign new_R1165_U549 = ~new_R1165_U547 | ~new_R1165_U321;
  assign new_R1165_U550 = ~new_R1165_U389 | ~new_U3177;
  assign new_R1165_U551 = ~new_R1165_U70 | ~new_R1165_U29;
  assign new_R1165_U552 = ~new_R1165_U389 | ~new_U3177;
  assign new_R1165_U553 = ~new_R1165_U70 | ~new_R1165_U29;
  assign new_R1165_U554 = ~new_R1165_U553 | ~new_R1165_U552;
  assign new_R1165_U555 = ~new_R1165_U188 | ~new_R1165_U189;
  assign new_R1165_U556 = ~new_R1165_U212 | ~new_R1165_U554;
  assign new_R1165_U557 = ~new_R1165_U486 | ~new_U3159;
  assign new_R1165_U558 = ~new_R1165_U81 | ~new_R1165_U49;
  assign new_R1165_U559 = ~new_R1165_U558 | ~new_R1165_U557;
  assign new_R1165_U560 = ~new_R1165_U350 | ~new_R1165_U190;
  assign new_R1165_U561 = ~new_R1165_U278 | ~new_R1165_U559;
  assign new_R1165_U562 = ~new_R1165_U477 | ~new_U3160;
  assign new_R1165_U563 = ~new_R1165_U80 | ~new_R1165_U47;
  assign new_R1165_U564 = ~new_R1165_U477 | ~new_U3160;
  assign new_R1165_U565 = ~new_R1165_U80 | ~new_R1165_U47;
  assign new_R1165_U566 = ~new_R1165_U565 | ~new_R1165_U564;
  assign new_R1165_U567 = ~new_R1165_U191 | ~new_R1165_U192;
  assign new_R1165_U568 = ~new_R1165_U274 | ~new_R1165_U566;
  assign new_R1165_U569 = ~new_R1165_U471 | ~new_U3161;
  assign new_R1165_U570 = ~new_R1165_U73 | ~new_R1165_U38;
  assign new_R1165_U571 = ~new_R1165_U474 | ~new_U3162;
  assign new_R1165_U572 = ~new_R1165_U72 | ~new_R1165_U36;
  assign new_R1165_U573 = ~new_R1165_U572 | ~new_R1165_U571;
  assign new_R1165_U574 = ~new_R1165_U351 | ~new_R1165_U60;
  assign new_R1165_U575 = ~new_R1165_U573 | ~new_R1165_U266;
  assign new_R1165_U576 = ~new_R1165_U468 | ~new_U3163;
  assign new_R1165_U577 = ~new_R1165_U79 | ~new_R1165_U46;
  assign new_R1165_U578 = ~new_R1165_U468 | ~new_U3163;
  assign new_R1165_U579 = ~new_R1165_U79 | ~new_R1165_U46;
  assign new_R1165_U580 = ~new_R1165_U579 | ~new_R1165_U578;
  assign new_R1165_U581 = ~new_R1165_U193 | ~new_R1165_U194;
  assign new_R1165_U582 = ~new_R1165_U262 | ~new_R1165_U580;
  assign new_R1165_U583 = ~new_R1165_U465 | ~new_U3164;
  assign new_R1165_U584 = ~new_R1165_U78 | ~new_R1165_U45;
  assign new_R1165_U585 = ~new_R1165_U465 | ~new_U3164;
  assign new_R1165_U586 = ~new_R1165_U78 | ~new_R1165_U45;
  assign new_R1165_U587 = ~new_R1165_U586 | ~new_R1165_U585;
  assign new_R1165_U588 = ~new_R1165_U195 | ~new_R1165_U196;
  assign new_R1165_U589 = ~new_R1165_U375 | ~new_R1165_U587;
  assign new_R1165_U590 = ~new_R1165_U456 | ~new_U3165;
  assign new_R1165_U591 = ~new_R1165_U75 | ~new_R1165_U42;
  assign new_R1165_U592 = ~new_R1165_U459 | ~new_U3166;
  assign new_R1165_U593 = ~new_R1165_U74 | ~new_R1165_U39;
  assign new_R1165_U594 = ~new_R1165_U593 | ~new_R1165_U592;
  assign new_R1165_U595 = ~new_R1165_U352 | ~new_R1165_U61;
  assign new_R1165_U596 = ~new_R1165_U594 | ~new_R1165_U337;
  assign new_R1165_U597 = ~new_R1165_U453 | ~new_U3167;
  assign new_R1165_U598 = ~new_R1165_U76 | ~new_R1165_U40;
  assign new_R1165_U599 = ~new_R1165_U598 | ~new_R1165_U597;
  assign new_R1165_U600 = ~new_R1165_U197 | ~new_R1165_U353;
  assign new_R1165_U601 = ~new_R1165_U373 | ~new_R1165_U599;
  assign new_R1165_U602 = ~new_R1165_U462 | ~new_U3168;
  assign new_R1165_U603 = ~new_R1165_U77 | ~new_R1165_U43;
  assign new_R1165_U604 = ~new_R1165_U462 | ~new_U3168;
  assign new_R1165_U605 = ~new_R1165_U77 | ~new_R1165_U43;
  assign new_R1165_U606 = ~new_R1165_U605 | ~new_R1165_U604;
  assign new_R1165_U607 = ~new_R1165_U198 | ~new_R1165_U199;
  assign new_R1165_U608 = ~new_R1165_U248 | ~new_R1165_U606;
  assign new_R1165_U609 = ~new_U3178 | ~new_R1165_U18;
  assign new_R1165_U610 = ~new_U3208 | ~new_R1165_U30;
  assign new_R1165_U611 = ~new_R1165_U141;
  assign new_R1165_U612 = ~new_R1165_U71 | ~new_R1165_U611;
  assign new_R1165_U613 = ~new_R1165_U141 | ~new_R1165_U392;
  assign new_R1150_U6 = new_R1150_U224 & new_R1150_U223;
  assign new_R1150_U7 = new_R1150_U204 & new_R1150_U257;
  assign new_R1150_U8 = new_R1150_U259 & new_R1150_U258;
  assign new_R1150_U9 = new_R1150_U205 & new_R1150_U268;
  assign new_R1150_U10 = new_R1150_U270 & new_R1150_U269;
  assign new_R1150_U11 = new_R1150_U206 & new_R1150_U286;
  assign new_R1150_U12 = new_R1150_U288 & new_R1150_U287;
  assign new_R1150_U13 = new_R1150_U227 & new_R1150_U222 & new_R1150_U209;
  assign new_R1150_U14 = new_R1150_U232 & new_R1150_U210;
  assign new_R1150_U15 = new_R1150_U7 & new_R1150_U237;
  assign new_R1150_U16 = new_R1150_U9 & new_R1150_U273;
  assign new_R1150_U17 = new_R1150_U11 & new_R1150_U291;
  assign new_R1150_U18 = new_R1150_U15 & new_R1150_U264;
  assign new_R1150_U19 = new_R1150_U284 & new_R1150_U282;
  assign new_R1150_U20 = new_R1150_U19 & new_R1150_U17;
  assign new_R1150_U21 = new_R1150_U20 & new_R1150_U294;
  assign new_R1150_U22 = new_R1150_U418 & new_R1150_U417;
  assign new_R1150_U23 = ~new_R1150_U335 | ~new_R1150_U338;
  assign new_R1150_U24 = ~new_R1150_U326 | ~new_R1150_U329;
  assign new_R1150_U25 = ~new_R1150_U315 | ~new_R1150_U318;
  assign new_R1150_U26 = ~new_R1150_U307 | ~new_R1150_U309;
  assign new_R1150_U27 = ~new_R1150_U344 | ~new_R1150_U179 | ~new_R1150_U199;
  assign new_R1150_U28 = ~new_R1150_U255 | ~new_R1150_U380;
  assign new_R1150_U29 = ~new_R1150_U248 | ~new_R1150_U251;
  assign new_R1150_U30 = ~new_R1150_U240 | ~new_R1150_U242;
  assign new_R1150_U31 = ~new_R1150_U189 | ~new_R1150_U341;
  assign new_R1150_U32 = ~new_U3067;
  assign new_R1150_U33 = ~new_U3067 | ~new_R1150_U38;
  assign new_R1150_U34 = ~new_U3081;
  assign new_R1150_U35 = ~new_U3476;
  assign new_R1150_U36 = ~new_U3478;
  assign new_R1150_U37 = ~new_U3474;
  assign new_R1150_U38 = ~new_U3480;
  assign new_R1150_U39 = ~new_U3482;
  assign new_R1150_U40 = ~new_U3065;
  assign new_R1150_U41 = ~new_U3065 | ~new_R1150_U43;
  assign new_R1150_U42 = ~new_U3061;
  assign new_R1150_U43 = ~new_U3470;
  assign new_R1150_U44 = ~new_U3464;
  assign new_R1150_U45 = ~new_U3075;
  assign new_R1150_U46 = ~new_U3472;
  assign new_R1150_U47 = ~new_U3068;
  assign new_R1150_U48 = ~new_U3064;
  assign new_R1150_U49 = ~new_U3057;
  assign new_R1150_U50 = ~new_U3057 | ~new_R1150_U37;
  assign new_R1150_U51 = ~new_R1150_U228 | ~new_R1150_U226;
  assign new_R1150_U52 = ~new_U3484;
  assign new_R1150_U53 = ~new_U3080;
  assign new_R1150_U54 = ~new_R1150_U51 | ~new_R1150_U229;
  assign new_R1150_U55 = ~new_R1150_U50 | ~new_R1150_U244;
  assign new_R1150_U56 = ~new_R1150_U342 | ~new_R1150_U216 | ~new_R1150_U200;
  assign new_R1150_U57 = ~new_U4031;
  assign new_R1150_U58 = ~new_U4030;
  assign new_R1150_U59 = ~new_U3055;
  assign new_R1150_U60 = ~new_U4032;
  assign new_R1150_U61 = ~new_U3062;
  assign new_R1150_U62 = ~new_U4033;
  assign new_R1150_U63 = ~new_U3063;
  assign new_R1150_U64 = ~new_U3058;
  assign new_R1150_U65 = ~new_U3072;
  assign new_R1150_U66 = ~new_U4034;
  assign new_R1150_U67 = ~new_U4035;
  assign new_R1150_U68 = ~new_U3072 | ~new_R1150_U69;
  assign new_R1150_U69 = ~new_U4036;
  assign new_R1150_U70 = ~new_U3073;
  assign new_R1150_U71 = ~new_U3078;
  assign new_R1150_U72 = ~new_U4037;
  assign new_R1150_U73 = ~new_U3078 | ~new_R1150_U74;
  assign new_R1150_U74 = ~new_U3504;
  assign new_R1150_U75 = ~new_U3079;
  assign new_R1150_U76 = ~new_U3066;
  assign new_R1150_U77 = ~new_U3500;
  assign new_R1150_U78 = ~new_U3498;
  assign new_R1150_U79 = ~new_U3496;
  assign new_R1150_U80 = ~new_U3494;
  assign new_R1150_U81 = ~new_U3077;
  assign new_R1150_U82 = ~new_U3492;
  assign new_R1150_U83 = ~new_U3490;
  assign new_R1150_U84 = ~new_U3060;
  assign new_R1150_U85 = ~new_U3059;
  assign new_R1150_U86 = ~new_U3488;
  assign new_R1150_U87 = ~new_U3486;
  assign new_R1150_U88 = ~new_U3080 | ~new_R1150_U52;
  assign new_R1150_U89 = ~new_U3069;
  assign new_R1150_U90 = ~new_R1150_U347 | ~new_R1150_U264;
  assign new_R1150_U91 = ~new_U3070;
  assign new_R1150_U92 = ~new_U3071;
  assign new_R1150_U93 = ~new_U3076;
  assign new_R1150_U94 = ~new_U3076 | ~new_R1150_U80;
  assign new_R1150_U95 = ~new_R1150_U274 | ~new_R1150_U272;
  assign new_R1150_U96 = ~new_U3502;
  assign new_R1150_U97 = ~new_U3054;
  assign new_R1150_U98 = ~new_U3054 | ~new_R1150_U57;
  assign new_R1150_U99 = ~new_U3050;
  assign new_R1150_U100 = ~new_U4029;
  assign new_R1150_U101 = ~new_U3051;
  assign new_R1150_U102 = ~new_R1150_U146 | ~new_R1150_U367;
  assign new_R1150_U103 = ~new_R1150_U356 | ~new_R1150_U295;
  assign new_R1150_U104 = ~new_R1150_U354 | ~new_R1150_U293;
  assign new_R1150_U105 = ~new_R1150_U352 | ~new_R1150_U285;
  assign new_R1150_U106 = ~new_R1150_U68 | ~new_R1150_U311;
  assign new_R1150_U107 = ~new_R1150_U94 | ~new_R1150_U322;
  assign new_R1150_U108 = ~new_R1150_U369 | ~new_R1150_U88;
  assign new_R1150_U109 = ~new_U3074;
  assign new_R1150_U110 = ~new_R1150_U428 | ~new_R1150_U427;
  assign new_R1150_U111 = ~new_R1150_U442 | ~new_R1150_U441;
  assign new_R1150_U112 = ~new_R1150_U447 | ~new_R1150_U446;
  assign new_R1150_U113 = ~new_R1150_U463 | ~new_R1150_U462;
  assign new_R1150_U114 = ~new_R1150_U468 | ~new_R1150_U467;
  assign new_R1150_U115 = ~new_R1150_U473 | ~new_R1150_U472;
  assign new_R1150_U116 = ~new_R1150_U478 | ~new_R1150_U477;
  assign new_R1150_U117 = ~new_R1150_U483 | ~new_R1150_U482;
  assign new_R1150_U118 = ~new_R1150_U499 | ~new_R1150_U498;
  assign new_R1150_U119 = ~new_R1150_U504 | ~new_R1150_U503;
  assign new_R1150_U120 = ~new_R1150_U387 | ~new_R1150_U386;
  assign new_R1150_U121 = ~new_R1150_U396 | ~new_R1150_U395;
  assign new_R1150_U122 = ~new_R1150_U403 | ~new_R1150_U402;
  assign new_R1150_U123 = ~new_R1150_U407 | ~new_R1150_U406;
  assign new_R1150_U124 = ~new_R1150_U416 | ~new_R1150_U415;
  assign new_R1150_U125 = ~new_R1150_U437 | ~new_R1150_U436;
  assign new_R1150_U126 = ~new_R1150_U454 | ~new_R1150_U453;
  assign new_R1150_U127 = ~new_R1150_U458 | ~new_R1150_U457;
  assign new_R1150_U128 = ~new_R1150_U490 | ~new_R1150_U489;
  assign new_R1150_U129 = ~new_R1150_U494 | ~new_R1150_U493;
  assign new_R1150_U130 = ~new_R1150_U511 | ~new_R1150_U510;
  assign new_R1150_U131 = new_R1150_U218 & new_R1150_U208;
  assign new_R1150_U132 = new_R1150_U221 & new_R1150_U220;
  assign new_R1150_U133 = new_R1150_U14 & new_R1150_U13;
  assign new_R1150_U134 = new_R1150_U235 & new_R1150_U234;
  assign new_R1150_U135 = new_R1150_U346 & new_R1150_U134;
  assign new_R1150_U136 = new_R1150_U33 & new_R1150_U389 & new_R1150_U388;
  assign new_R1150_U137 = new_R1150_U392 & new_R1150_U210;
  assign new_R1150_U138 = new_R1150_U250 & new_R1150_U6;
  assign new_R1150_U139 = new_R1150_U399 & new_R1150_U209;
  assign new_R1150_U140 = new_R1150_U41 & new_R1150_U409 & new_R1150_U408;
  assign new_R1150_U141 = new_R1150_U412 & new_R1150_U208;
  assign new_R1150_U142 = new_R1150_U266 & new_R1150_U18;
  assign new_R1150_U143 = new_R1150_U16 & new_R1150_U278;
  assign new_R1150_U144 = new_R1150_U351 & new_R1150_U279;
  assign new_R1150_U145 = new_R1150_U21 & new_R1150_U296;
  assign new_R1150_U146 = new_R1150_U358 & new_R1150_U297;
  assign new_R1150_U147 = new_R1150_U298 & new_R1150_U207;
  assign new_R1150_U148 = new_R1150_U301 & new_R1150_U302;
  assign new_R1150_U149 = new_R1150_U304 & new_R1150_U421;
  assign new_R1150_U150 = new_R1150_U301 & new_R1150_U302;
  assign new_R1150_U151 = new_R1150_U22 & new_R1150_U305;
  assign new_R1150_U152 = ~new_R1150_U425 | ~new_R1150_U424;
  assign new_R1150_U153 = new_R1150_U98 & new_R1150_U430 & new_R1150_U429;
  assign new_R1150_U154 = new_R1150_U433 & new_R1150_U207;
  assign new_R1150_U155 = ~new_R1150_U439 | ~new_R1150_U438;
  assign new_R1150_U156 = ~new_R1150_U444 | ~new_R1150_U443;
  assign new_R1150_U157 = new_R1150_U317 & new_R1150_U12;
  assign new_R1150_U158 = new_R1150_U450 & new_R1150_U206;
  assign new_R1150_U159 = ~new_R1150_U460 | ~new_R1150_U459;
  assign new_R1150_U160 = ~new_R1150_U465 | ~new_R1150_U464;
  assign new_R1150_U161 = ~new_R1150_U470 | ~new_R1150_U469;
  assign new_R1150_U162 = ~new_R1150_U475 | ~new_R1150_U474;
  assign new_R1150_U163 = ~new_R1150_U480 | ~new_R1150_U479;
  assign new_R1150_U164 = new_R1150_U328 & new_R1150_U10;
  assign new_R1150_U165 = new_R1150_U486 & new_R1150_U205;
  assign new_R1150_U166 = ~new_R1150_U496 | ~new_R1150_U495;
  assign new_R1150_U167 = ~new_R1150_U501 | ~new_R1150_U500;
  assign new_R1150_U168 = new_R1150_U337 & new_R1150_U8;
  assign new_R1150_U169 = new_R1150_U507 & new_R1150_U204;
  assign new_R1150_U170 = new_R1150_U385 & new_R1150_U384;
  assign new_R1150_U171 = ~new_R1150_U135 | ~new_R1150_U345;
  assign new_R1150_U172 = new_R1150_U394 & new_R1150_U393;
  assign new_R1150_U173 = new_R1150_U401 & new_R1150_U400;
  assign new_R1150_U174 = new_R1150_U405 & new_R1150_U404;
  assign new_R1150_U175 = ~new_R1150_U132 | ~new_R1150_U377;
  assign new_R1150_U176 = new_R1150_U414 & new_R1150_U413;
  assign new_R1150_U177 = ~new_U4040;
  assign new_R1150_U178 = ~new_U3052;
  assign new_R1150_U179 = new_R1150_U423 & new_R1150_U422;
  assign new_R1150_U180 = ~new_R1150_U148 | ~new_R1150_U299;
  assign new_R1150_U181 = new_R1150_U435 & new_R1150_U434;
  assign new_R1150_U182 = ~new_R1150_U357 | ~new_R1150_U365;
  assign new_R1150_U183 = ~new_R1150_U355 | ~new_R1150_U363;
  assign new_R1150_U184 = new_R1150_U452 & new_R1150_U451;
  assign new_R1150_U185 = new_R1150_U456 & new_R1150_U455;
  assign new_R1150_U186 = ~new_R1150_U353 | ~new_R1150_U361;
  assign new_R1150_U187 = ~new_R1150_U359 | ~new_R1150_U73;
  assign new_R1150_U188 = ~new_U3468;
  assign new_R1150_U189 = ~new_U3464 | ~new_R1150_U109;
  assign new_R1150_U190 = ~new_R1150_U382 | ~new_R1150_U343;
  assign new_R1150_U191 = ~new_R1150_U144 | ~new_R1150_U350;
  assign new_R1150_U192 = ~new_R1150_U95 | ~new_R1150_U275;
  assign new_R1150_U193 = new_R1150_U488 & new_R1150_U487;
  assign new_R1150_U194 = new_R1150_U492 & new_R1150_U491;
  assign new_R1150_U195 = ~new_R1150_U375 | ~new_R1150_U349 | ~new_R1150_U267;
  assign new_R1150_U196 = ~new_R1150_U373 | ~new_R1150_U90;
  assign new_R1150_U197 = ~new_R1150_U371 | ~new_R1150_U263;
  assign new_R1150_U198 = new_R1150_U509 & new_R1150_U508;
  assign new_R1150_U199 = ~new_R1150_U149 | ~new_R1150_U180;
  assign new_R1150_U200 = ~new_R1150_U189 | ~new_R1150_U188;
  assign new_R1150_U201 = ~new_R1150_U98;
  assign new_R1150_U202 = ~new_R1150_U41;
  assign new_R1150_U203 = ~new_R1150_U33;
  assign new_R1150_U204 = ~new_U3486 | ~new_R1150_U85;
  assign new_R1150_U205 = ~new_U3496 | ~new_R1150_U92;
  assign new_R1150_U206 = ~new_U4035 | ~new_R1150_U64;
  assign new_R1150_U207 = ~new_U4031 | ~new_R1150_U97;
  assign new_R1150_U208 = ~new_U3470 | ~new_R1150_U40;
  assign new_R1150_U209 = ~new_U3476 | ~new_R1150_U48;
  assign new_R1150_U210 = ~new_U3480 | ~new_R1150_U32;
  assign new_R1150_U211 = ~new_R1150_U94;
  assign new_R1150_U212 = ~new_R1150_U68;
  assign new_R1150_U213 = ~new_R1150_U50;
  assign new_R1150_U214 = ~new_R1150_U88;
  assign new_R1150_U215 = ~new_R1150_U189;
  assign new_R1150_U216 = ~new_U3075 | ~new_R1150_U189;
  assign new_R1150_U217 = ~new_R1150_U56;
  assign new_R1150_U218 = ~new_U3472 | ~new_R1150_U42;
  assign new_R1150_U219 = ~new_R1150_U42 | ~new_R1150_U41;
  assign new_R1150_U220 = ~new_R1150_U219 | ~new_R1150_U46;
  assign new_R1150_U221 = ~new_U3061 | ~new_R1150_U202;
  assign new_R1150_U222 = ~new_U3478 | ~new_R1150_U47;
  assign new_R1150_U223 = ~new_U3068 | ~new_R1150_U36;
  assign new_R1150_U224 = ~new_U3064 | ~new_R1150_U35;
  assign new_R1150_U225 = ~new_R1150_U213 | ~new_R1150_U209;
  assign new_R1150_U226 = ~new_R1150_U6 | ~new_R1150_U225;
  assign new_R1150_U227 = ~new_U3474 | ~new_R1150_U49;
  assign new_R1150_U228 = ~new_U3478 | ~new_R1150_U47;
  assign new_R1150_U229 = ~new_R1150_U13 | ~new_R1150_U175;
  assign new_R1150_U230 = ~new_R1150_U51;
  assign new_R1150_U231 = ~new_R1150_U54;
  assign new_R1150_U232 = ~new_U3482 | ~new_R1150_U34;
  assign new_R1150_U233 = ~new_R1150_U34 | ~new_R1150_U33;
  assign new_R1150_U234 = ~new_R1150_U233 | ~new_R1150_U39;
  assign new_R1150_U235 = ~new_U3081 | ~new_R1150_U203;
  assign new_R1150_U236 = ~new_R1150_U171;
  assign new_R1150_U237 = ~new_U3484 | ~new_R1150_U53;
  assign new_R1150_U238 = ~new_R1150_U237 | ~new_R1150_U88;
  assign new_R1150_U239 = ~new_R1150_U231 | ~new_R1150_U33;
  assign new_R1150_U240 = ~new_R1150_U137 | ~new_R1150_U239;
  assign new_R1150_U241 = ~new_R1150_U54 | ~new_R1150_U210;
  assign new_R1150_U242 = ~new_R1150_U136 | ~new_R1150_U241;
  assign new_R1150_U243 = ~new_R1150_U33 | ~new_R1150_U210;
  assign new_R1150_U244 = ~new_R1150_U227 | ~new_R1150_U175;
  assign new_R1150_U245 = ~new_R1150_U55;
  assign new_R1150_U246 = ~new_U3064 | ~new_R1150_U35;
  assign new_R1150_U247 = ~new_R1150_U245 | ~new_R1150_U246;
  assign new_R1150_U248 = ~new_R1150_U139 | ~new_R1150_U247;
  assign new_R1150_U249 = ~new_R1150_U55 | ~new_R1150_U209;
  assign new_R1150_U250 = ~new_U3478 | ~new_R1150_U47;
  assign new_R1150_U251 = ~new_R1150_U138 | ~new_R1150_U249;
  assign new_R1150_U252 = ~new_U3064 | ~new_R1150_U35;
  assign new_R1150_U253 = ~new_R1150_U209 | ~new_R1150_U252;
  assign new_R1150_U254 = ~new_R1150_U227 | ~new_R1150_U50;
  assign new_R1150_U255 = ~new_R1150_U141 | ~new_R1150_U381;
  assign new_R1150_U256 = ~new_R1150_U41 | ~new_R1150_U208;
  assign new_R1150_U257 = ~new_U3488 | ~new_R1150_U84;
  assign new_R1150_U258 = ~new_U3060 | ~new_R1150_U86;
  assign new_R1150_U259 = ~new_U3059 | ~new_R1150_U87;
  assign new_R1150_U260 = ~new_R1150_U214 | ~new_R1150_U7;
  assign new_R1150_U261 = ~new_R1150_U8 | ~new_R1150_U260;
  assign new_R1150_U262 = ~new_U3488 | ~new_R1150_U84;
  assign new_R1150_U263 = ~new_R1150_U262 | ~new_R1150_U261;
  assign new_R1150_U264 = ~new_U3490 | ~new_R1150_U89;
  assign new_R1150_U265 = ~new_U3069 | ~new_R1150_U83;
  assign new_R1150_U266 = ~new_U3492 | ~new_R1150_U81;
  assign new_R1150_U267 = ~new_U3077 | ~new_R1150_U82;
  assign new_R1150_U268 = ~new_U3498 | ~new_R1150_U91;
  assign new_R1150_U269 = ~new_U3070 | ~new_R1150_U78;
  assign new_R1150_U270 = ~new_U3071 | ~new_R1150_U79;
  assign new_R1150_U271 = ~new_R1150_U211 | ~new_R1150_U9;
  assign new_R1150_U272 = ~new_R1150_U10 | ~new_R1150_U271;
  assign new_R1150_U273 = ~new_U3494 | ~new_R1150_U93;
  assign new_R1150_U274 = ~new_U3498 | ~new_R1150_U91;
  assign new_R1150_U275 = ~new_R1150_U16 | ~new_R1150_U195;
  assign new_R1150_U276 = ~new_R1150_U95;
  assign new_R1150_U277 = ~new_R1150_U192;
  assign new_R1150_U278 = ~new_U3500 | ~new_R1150_U76;
  assign new_R1150_U279 = ~new_U3066 | ~new_R1150_U77;
  assign new_R1150_U280 = ~new_R1150_U191;
  assign new_R1150_U281 = ~new_U3502 | ~new_R1150_U75;
  assign new_R1150_U282 = ~new_U3504 | ~new_R1150_U71;
  assign new_R1150_U283 = ~new_R1150_U73;
  assign new_R1150_U284 = ~new_U4037 | ~new_R1150_U70;
  assign new_R1150_U285 = ~new_U3073 | ~new_R1150_U72;
  assign new_R1150_U286 = ~new_U4034 | ~new_R1150_U63;
  assign new_R1150_U287 = ~new_U3063 | ~new_R1150_U66;
  assign new_R1150_U288 = ~new_U3058 | ~new_R1150_U67;
  assign new_R1150_U289 = ~new_R1150_U212 | ~new_R1150_U11;
  assign new_R1150_U290 = ~new_R1150_U12 | ~new_R1150_U289;
  assign new_R1150_U291 = ~new_U4036 | ~new_R1150_U65;
  assign new_R1150_U292 = ~new_U4034 | ~new_R1150_U63;
  assign new_R1150_U293 = ~new_R1150_U292 | ~new_R1150_U290;
  assign new_R1150_U294 = ~new_U4033 | ~new_R1150_U61;
  assign new_R1150_U295 = ~new_U3062 | ~new_R1150_U62;
  assign new_R1150_U296 = ~new_U4032 | ~new_R1150_U59;
  assign new_R1150_U297 = ~new_U3055 | ~new_R1150_U60;
  assign new_R1150_U298 = ~new_U4030 | ~new_R1150_U99;
  assign new_R1150_U299 = ~new_R1150_U147 | ~new_R1150_U102;
  assign new_R1150_U300 = ~new_R1150_U99 | ~new_R1150_U98;
  assign new_R1150_U301 = ~new_R1150_U300 | ~new_R1150_U58;
  assign new_R1150_U302 = ~new_U3050 | ~new_R1150_U201;
  assign new_R1150_U303 = ~new_R1150_U180;
  assign new_R1150_U304 = ~new_U4029 | ~new_R1150_U101;
  assign new_R1150_U305 = ~new_U3051 | ~new_R1150_U100;
  assign new_R1150_U306 = ~new_R1150_U368 | ~new_R1150_U98;
  assign new_R1150_U307 = ~new_R1150_U154 | ~new_R1150_U306;
  assign new_R1150_U308 = ~new_R1150_U102 | ~new_R1150_U207;
  assign new_R1150_U309 = ~new_R1150_U153 | ~new_R1150_U308;
  assign new_R1150_U310 = ~new_R1150_U98 | ~new_R1150_U207;
  assign new_R1150_U311 = ~new_R1150_U291 | ~new_R1150_U186;
  assign new_R1150_U312 = ~new_R1150_U106;
  assign new_R1150_U313 = ~new_U3058 | ~new_R1150_U67;
  assign new_R1150_U314 = ~new_R1150_U312 | ~new_R1150_U313;
  assign new_R1150_U315 = ~new_R1150_U158 | ~new_R1150_U314;
  assign new_R1150_U316 = ~new_R1150_U106 | ~new_R1150_U206;
  assign new_R1150_U317 = ~new_U4034 | ~new_R1150_U63;
  assign new_R1150_U318 = ~new_R1150_U157 | ~new_R1150_U316;
  assign new_R1150_U319 = ~new_U3058 | ~new_R1150_U67;
  assign new_R1150_U320 = ~new_R1150_U206 | ~new_R1150_U319;
  assign new_R1150_U321 = ~new_R1150_U291 | ~new_R1150_U68;
  assign new_R1150_U322 = ~new_R1150_U273 | ~new_R1150_U195;
  assign new_R1150_U323 = ~new_R1150_U107;
  assign new_R1150_U324 = ~new_U3071 | ~new_R1150_U79;
  assign new_R1150_U325 = ~new_R1150_U323 | ~new_R1150_U324;
  assign new_R1150_U326 = ~new_R1150_U165 | ~new_R1150_U325;
  assign new_R1150_U327 = ~new_R1150_U107 | ~new_R1150_U205;
  assign new_R1150_U328 = ~new_U3498 | ~new_R1150_U91;
  assign new_R1150_U329 = ~new_R1150_U164 | ~new_R1150_U327;
  assign new_R1150_U330 = ~new_U3071 | ~new_R1150_U79;
  assign new_R1150_U331 = ~new_R1150_U205 | ~new_R1150_U330;
  assign new_R1150_U332 = ~new_R1150_U273 | ~new_R1150_U94;
  assign new_R1150_U333 = ~new_U3059 | ~new_R1150_U87;
  assign new_R1150_U334 = ~new_R1150_U370 | ~new_R1150_U333;
  assign new_R1150_U335 = ~new_R1150_U169 | ~new_R1150_U334;
  assign new_R1150_U336 = ~new_R1150_U108 | ~new_R1150_U204;
  assign new_R1150_U337 = ~new_U3488 | ~new_R1150_U84;
  assign new_R1150_U338 = ~new_R1150_U168 | ~new_R1150_U336;
  assign new_R1150_U339 = ~new_U3059 | ~new_R1150_U87;
  assign new_R1150_U340 = ~new_R1150_U204 | ~new_R1150_U339;
  assign new_R1150_U341 = ~new_U3074 | ~new_R1150_U44;
  assign new_R1150_U342 = ~new_U3075 | ~new_R1150_U188;
  assign new_R1150_U343 = ~new_U3079 | ~new_R1150_U96;
  assign new_R1150_U344 = ~new_R1150_U151 | ~new_R1150_U150 | ~new_R1150_U299;
  assign new_R1150_U345 = ~new_R1150_U133 | ~new_R1150_U175;
  assign new_R1150_U346 = ~new_R1150_U230 | ~new_R1150_U14;
  assign new_R1150_U347 = ~new_R1150_U265 | ~new_R1150_U263;
  assign new_R1150_U348 = ~new_R1150_U90;
  assign new_R1150_U349 = ~new_R1150_U348 | ~new_R1150_U266;
  assign new_R1150_U350 = ~new_R1150_U143 | ~new_R1150_U195;
  assign new_R1150_U351 = ~new_R1150_U276 | ~new_R1150_U278;
  assign new_R1150_U352 = ~new_R1150_U283 | ~new_R1150_U284;
  assign new_R1150_U353 = ~new_R1150_U105;
  assign new_R1150_U354 = ~new_R1150_U17 | ~new_R1150_U105;
  assign new_R1150_U355 = ~new_R1150_U104;
  assign new_R1150_U356 = ~new_R1150_U104 | ~new_R1150_U294;
  assign new_R1150_U357 = ~new_R1150_U103;
  assign new_R1150_U358 = ~new_R1150_U103 | ~new_R1150_U296;
  assign new_R1150_U359 = ~new_R1150_U282 | ~new_R1150_U190;
  assign new_R1150_U360 = ~new_R1150_U187;
  assign new_R1150_U361 = ~new_R1150_U19 | ~new_R1150_U190;
  assign new_R1150_U362 = ~new_R1150_U186;
  assign new_R1150_U363 = ~new_R1150_U20 | ~new_R1150_U190;
  assign new_R1150_U364 = ~new_R1150_U183;
  assign new_R1150_U365 = ~new_R1150_U21 | ~new_R1150_U190;
  assign new_R1150_U366 = ~new_R1150_U182;
  assign new_R1150_U367 = ~new_R1150_U145 | ~new_R1150_U190;
  assign new_R1150_U368 = ~new_R1150_U102;
  assign new_R1150_U369 = ~new_R1150_U237 | ~new_R1150_U171;
  assign new_R1150_U370 = ~new_R1150_U108;
  assign new_R1150_U371 = ~new_R1150_U15 | ~new_R1150_U171;
  assign new_R1150_U372 = ~new_R1150_U197;
  assign new_R1150_U373 = ~new_R1150_U18 | ~new_R1150_U171;
  assign new_R1150_U374 = ~new_R1150_U196;
  assign new_R1150_U375 = ~new_R1150_U142 | ~new_R1150_U171;
  assign new_R1150_U376 = ~new_R1150_U195;
  assign new_R1150_U377 = ~new_R1150_U131 | ~new_R1150_U56;
  assign new_R1150_U378 = ~new_R1150_U175;
  assign new_R1150_U379 = ~new_R1150_U208 | ~new_R1150_U56;
  assign new_R1150_U380 = ~new_R1150_U140 | ~new_R1150_U379;
  assign new_R1150_U381 = ~new_R1150_U217 | ~new_R1150_U41;
  assign new_R1150_U382 = ~new_R1150_U281 | ~new_R1150_U191;
  assign new_R1150_U383 = ~new_R1150_U190;
  assign new_R1150_U384 = ~new_U3484 | ~new_R1150_U53;
  assign new_R1150_U385 = ~new_U3080 | ~new_R1150_U52;
  assign new_R1150_U386 = ~new_R1150_U238 | ~new_R1150_U171;
  assign new_R1150_U387 = ~new_R1150_U236 | ~new_R1150_U170;
  assign new_R1150_U388 = ~new_U3482 | ~new_R1150_U34;
  assign new_R1150_U389 = ~new_U3081 | ~new_R1150_U39;
  assign new_R1150_U390 = ~new_U3482 | ~new_R1150_U34;
  assign new_R1150_U391 = ~new_U3081 | ~new_R1150_U39;
  assign new_R1150_U392 = ~new_R1150_U391 | ~new_R1150_U390;
  assign new_R1150_U393 = ~new_U3480 | ~new_R1150_U32;
  assign new_R1150_U394 = ~new_U3067 | ~new_R1150_U38;
  assign new_R1150_U395 = ~new_R1150_U243 | ~new_R1150_U54;
  assign new_R1150_U396 = ~new_R1150_U172 | ~new_R1150_U231;
  assign new_R1150_U397 = ~new_U3478 | ~new_R1150_U47;
  assign new_R1150_U398 = ~new_U3068 | ~new_R1150_U36;
  assign new_R1150_U399 = ~new_R1150_U398 | ~new_R1150_U397;
  assign new_R1150_U400 = ~new_U3476 | ~new_R1150_U48;
  assign new_R1150_U401 = ~new_U3064 | ~new_R1150_U35;
  assign new_R1150_U402 = ~new_R1150_U253 | ~new_R1150_U55;
  assign new_R1150_U403 = ~new_R1150_U173 | ~new_R1150_U245;
  assign new_R1150_U404 = ~new_U3474 | ~new_R1150_U49;
  assign new_R1150_U405 = ~new_U3057 | ~new_R1150_U37;
  assign new_R1150_U406 = ~new_R1150_U175 | ~new_R1150_U254;
  assign new_R1150_U407 = ~new_R1150_U378 | ~new_R1150_U174;
  assign new_R1150_U408 = ~new_U3472 | ~new_R1150_U42;
  assign new_R1150_U409 = ~new_U3061 | ~new_R1150_U46;
  assign new_R1150_U410 = ~new_U3472 | ~new_R1150_U42;
  assign new_R1150_U411 = ~new_U3061 | ~new_R1150_U46;
  assign new_R1150_U412 = ~new_R1150_U411 | ~new_R1150_U410;
  assign new_R1150_U413 = ~new_U3470 | ~new_R1150_U40;
  assign new_R1150_U414 = ~new_U3065 | ~new_R1150_U43;
  assign new_R1150_U415 = ~new_R1150_U256 | ~new_R1150_U56;
  assign new_R1150_U416 = ~new_R1150_U176 | ~new_R1150_U217;
  assign new_R1150_U417 = ~new_U4040 | ~new_R1150_U178;
  assign new_R1150_U418 = ~new_U3052 | ~new_R1150_U177;
  assign new_R1150_U419 = ~new_U4040 | ~new_R1150_U178;
  assign new_R1150_U420 = ~new_U3052 | ~new_R1150_U177;
  assign new_R1150_U421 = ~new_R1150_U420 | ~new_R1150_U419;
  assign new_R1150_U422 = ~new_R1150_U100 | ~new_U3051 | ~new_R1150_U421;
  assign new_R1150_U423 = ~new_U4029 | ~new_R1150_U22 | ~new_R1150_U101;
  assign new_R1150_U424 = ~new_U4029 | ~new_R1150_U101;
  assign new_R1150_U425 = ~new_U3051 | ~new_R1150_U100;
  assign new_R1150_U426 = ~new_R1150_U152;
  assign new_R1150_U427 = ~new_R1150_U303 | ~new_R1150_U426;
  assign new_R1150_U428 = ~new_R1150_U152 | ~new_R1150_U180;
  assign new_R1150_U429 = ~new_U4030 | ~new_R1150_U99;
  assign new_R1150_U430 = ~new_U3050 | ~new_R1150_U58;
  assign new_R1150_U431 = ~new_U4030 | ~new_R1150_U99;
  assign new_R1150_U432 = ~new_U3050 | ~new_R1150_U58;
  assign new_R1150_U433 = ~new_R1150_U432 | ~new_R1150_U431;
  assign new_R1150_U434 = ~new_U4031 | ~new_R1150_U97;
  assign new_R1150_U435 = ~new_U3054 | ~new_R1150_U57;
  assign new_R1150_U436 = ~new_R1150_U102 | ~new_R1150_U310;
  assign new_R1150_U437 = ~new_R1150_U181 | ~new_R1150_U368;
  assign new_R1150_U438 = ~new_U4032 | ~new_R1150_U59;
  assign new_R1150_U439 = ~new_U3055 | ~new_R1150_U60;
  assign new_R1150_U440 = ~new_R1150_U155;
  assign new_R1150_U441 = ~new_R1150_U366 | ~new_R1150_U440;
  assign new_R1150_U442 = ~new_R1150_U155 | ~new_R1150_U182;
  assign new_R1150_U443 = ~new_U4033 | ~new_R1150_U61;
  assign new_R1150_U444 = ~new_U3062 | ~new_R1150_U62;
  assign new_R1150_U445 = ~new_R1150_U156;
  assign new_R1150_U446 = ~new_R1150_U364 | ~new_R1150_U445;
  assign new_R1150_U447 = ~new_R1150_U156 | ~new_R1150_U183;
  assign new_R1150_U448 = ~new_U4034 | ~new_R1150_U63;
  assign new_R1150_U449 = ~new_U3063 | ~new_R1150_U66;
  assign new_R1150_U450 = ~new_R1150_U449 | ~new_R1150_U448;
  assign new_R1150_U451 = ~new_U4035 | ~new_R1150_U64;
  assign new_R1150_U452 = ~new_U3058 | ~new_R1150_U67;
  assign new_R1150_U453 = ~new_R1150_U320 | ~new_R1150_U106;
  assign new_R1150_U454 = ~new_R1150_U184 | ~new_R1150_U312;
  assign new_R1150_U455 = ~new_U4036 | ~new_R1150_U65;
  assign new_R1150_U456 = ~new_U3072 | ~new_R1150_U69;
  assign new_R1150_U457 = ~new_R1150_U186 | ~new_R1150_U321;
  assign new_R1150_U458 = ~new_R1150_U362 | ~new_R1150_U185;
  assign new_R1150_U459 = ~new_U4037 | ~new_R1150_U70;
  assign new_R1150_U460 = ~new_U3073 | ~new_R1150_U72;
  assign new_R1150_U461 = ~new_R1150_U159;
  assign new_R1150_U462 = ~new_R1150_U360 | ~new_R1150_U461;
  assign new_R1150_U463 = ~new_R1150_U159 | ~new_R1150_U187;
  assign new_R1150_U464 = ~new_U3468 | ~new_R1150_U45;
  assign new_R1150_U465 = ~new_U3075 | ~new_R1150_U188;
  assign new_R1150_U466 = ~new_R1150_U160;
  assign new_R1150_U467 = ~new_R1150_U215 | ~new_R1150_U466;
  assign new_R1150_U468 = ~new_R1150_U160 | ~new_R1150_U189;
  assign new_R1150_U469 = ~new_U3504 | ~new_R1150_U71;
  assign new_R1150_U470 = ~new_U3078 | ~new_R1150_U74;
  assign new_R1150_U471 = ~new_R1150_U161;
  assign new_R1150_U472 = ~new_R1150_U383 | ~new_R1150_U471;
  assign new_R1150_U473 = ~new_R1150_U161 | ~new_R1150_U190;
  assign new_R1150_U474 = ~new_U3502 | ~new_R1150_U75;
  assign new_R1150_U475 = ~new_U3079 | ~new_R1150_U96;
  assign new_R1150_U476 = ~new_R1150_U162;
  assign new_R1150_U477 = ~new_R1150_U280 | ~new_R1150_U476;
  assign new_R1150_U478 = ~new_R1150_U162 | ~new_R1150_U191;
  assign new_R1150_U479 = ~new_U3500 | ~new_R1150_U76;
  assign new_R1150_U480 = ~new_U3066 | ~new_R1150_U77;
  assign new_R1150_U481 = ~new_R1150_U163;
  assign new_R1150_U482 = ~new_R1150_U277 | ~new_R1150_U481;
  assign new_R1150_U483 = ~new_R1150_U163 | ~new_R1150_U192;
  assign new_R1150_U484 = ~new_U3498 | ~new_R1150_U91;
  assign new_R1150_U485 = ~new_U3070 | ~new_R1150_U78;
  assign new_R1150_U486 = ~new_R1150_U485 | ~new_R1150_U484;
  assign new_R1150_U487 = ~new_U3496 | ~new_R1150_U92;
  assign new_R1150_U488 = ~new_U3071 | ~new_R1150_U79;
  assign new_R1150_U489 = ~new_R1150_U331 | ~new_R1150_U107;
  assign new_R1150_U490 = ~new_R1150_U193 | ~new_R1150_U323;
  assign new_R1150_U491 = ~new_U3494 | ~new_R1150_U93;
  assign new_R1150_U492 = ~new_U3076 | ~new_R1150_U80;
  assign new_R1150_U493 = ~new_R1150_U195 | ~new_R1150_U332;
  assign new_R1150_U494 = ~new_R1150_U376 | ~new_R1150_U194;
  assign new_R1150_U495 = ~new_U3492 | ~new_R1150_U81;
  assign new_R1150_U496 = ~new_U3077 | ~new_R1150_U82;
  assign new_R1150_U497 = ~new_R1150_U166;
  assign new_R1150_U498 = ~new_R1150_U374 | ~new_R1150_U497;
  assign new_R1150_U499 = ~new_R1150_U166 | ~new_R1150_U196;
  assign new_R1150_U500 = ~new_U3490 | ~new_R1150_U89;
  assign new_R1150_U501 = ~new_U3069 | ~new_R1150_U83;
  assign new_R1150_U502 = ~new_R1150_U167;
  assign new_R1150_U503 = ~new_R1150_U372 | ~new_R1150_U502;
  assign new_R1150_U504 = ~new_R1150_U167 | ~new_R1150_U197;
  assign new_R1150_U505 = ~new_U3488 | ~new_R1150_U84;
  assign new_R1150_U506 = ~new_U3060 | ~new_R1150_U86;
  assign new_R1150_U507 = ~new_R1150_U506 | ~new_R1150_U505;
  assign new_R1150_U508 = ~new_U3486 | ~new_R1150_U85;
  assign new_R1150_U509 = ~new_U3059 | ~new_R1150_U87;
  assign new_R1150_U510 = ~new_R1150_U108 | ~new_R1150_U340;
  assign new_R1150_U511 = ~new_R1150_U198 | ~new_R1150_U370;
  assign new_R1192_U6 = new_R1192_U231 & new_R1192_U230;
  assign new_R1192_U7 = new_R1192_U211 & new_R1192_U264;
  assign new_R1192_U8 = new_R1192_U266 & new_R1192_U265;
  assign new_R1192_U9 = new_R1192_U212 & new_R1192_U275;
  assign new_R1192_U10 = new_R1192_U277 & new_R1192_U276;
  assign new_R1192_U11 = new_R1192_U106 & new_R1192_U293;
  assign new_R1192_U12 = new_R1192_U295 & new_R1192_U294;
  assign new_R1192_U13 = new_R1192_U234 & new_R1192_U229 & new_R1192_U216;
  assign new_R1192_U14 = new_R1192_U239 & new_R1192_U217;
  assign new_R1192_U15 = new_R1192_U7 & new_R1192_U244;
  assign new_R1192_U16 = new_R1192_U9 & new_R1192_U280;
  assign new_R1192_U17 = new_R1192_U11 & new_R1192_U298;
  assign new_R1192_U18 = new_R1192_U15 & new_R1192_U271;
  assign new_R1192_U19 = new_R1192_U291 & new_R1192_U289;
  assign new_R1192_U20 = new_R1192_U19 & new_R1192_U17;
  assign new_R1192_U21 = new_R1192_U20 & new_R1192_U301;
  assign new_R1192_U22 = new_R1192_U457 & new_R1192_U106;
  assign new_R1192_U23 = new_R1192_U423 & new_R1192_U422;
  assign new_R1192_U24 = ~new_R1192_U334 | ~new_R1192_U337;
  assign new_R1192_U25 = ~new_R1192_U325 | ~new_R1192_U328;
  assign new_R1192_U26 = ~new_R1192_U359 | ~new_R1192_U387 | ~new_R1192_U388 | ~new_R1192_U459 | ~new_R1192_U458;
  assign new_R1192_U27 = new_R1192_U344 & new_R1192_U313;
  assign new_R1192_U28 = ~new_R1192_U343 | ~new_R1192_U182 | ~new_R1192_U206;
  assign new_R1192_U29 = ~new_R1192_U262 | ~new_R1192_U383;
  assign new_R1192_U30 = ~new_R1192_U255 | ~new_R1192_U258;
  assign new_R1192_U31 = ~new_R1192_U247 | ~new_R1192_U249;
  assign new_R1192_U32 = ~new_R1192_U195 | ~new_R1192_U340;
  assign new_R1192_U33 = ~new_U3067;
  assign new_R1192_U34 = ~new_U3067 | ~new_R1192_U39;
  assign new_R1192_U35 = ~new_U3081;
  assign new_R1192_U36 = ~new_U3476;
  assign new_R1192_U37 = ~new_U3478;
  assign new_R1192_U38 = ~new_U3474;
  assign new_R1192_U39 = ~new_U3480;
  assign new_R1192_U40 = ~new_U3482;
  assign new_R1192_U41 = ~new_U3065;
  assign new_R1192_U42 = ~new_U3065 | ~new_R1192_U44;
  assign new_R1192_U43 = ~new_U3061;
  assign new_R1192_U44 = ~new_U3470;
  assign new_R1192_U45 = ~new_U3464;
  assign new_R1192_U46 = ~new_U3075;
  assign new_R1192_U47 = ~new_U3472;
  assign new_R1192_U48 = ~new_U3068;
  assign new_R1192_U49 = ~new_U3064;
  assign new_R1192_U50 = ~new_U3057;
  assign new_R1192_U51 = ~new_U3057 | ~new_R1192_U38;
  assign new_R1192_U52 = ~new_R1192_U235 | ~new_R1192_U233;
  assign new_R1192_U53 = ~new_U3484;
  assign new_R1192_U54 = ~new_U3080;
  assign new_R1192_U55 = ~new_R1192_U52 | ~new_R1192_U236;
  assign new_R1192_U56 = ~new_R1192_U51 | ~new_R1192_U251;
  assign new_R1192_U57 = ~new_R1192_U341 | ~new_R1192_U223 | ~new_R1192_U207;
  assign new_R1192_U58 = ~new_U4031;
  assign new_R1192_U59 = ~new_U4030;
  assign new_R1192_U60 = ~new_U3055;
  assign new_R1192_U61 = ~new_U4032;
  assign new_R1192_U62 = ~new_U3062;
  assign new_R1192_U63 = ~new_U4033;
  assign new_R1192_U64 = ~new_U3063;
  assign new_R1192_U65 = ~new_U3058;
  assign new_R1192_U66 = ~new_U3072;
  assign new_R1192_U67 = ~new_U4034;
  assign new_R1192_U68 = ~new_U4035;
  assign new_R1192_U69 = ~new_U3072 | ~new_R1192_U70;
  assign new_R1192_U70 = ~new_U4036;
  assign new_R1192_U71 = ~new_U3073;
  assign new_R1192_U72 = ~new_U3078;
  assign new_R1192_U73 = ~new_U4037;
  assign new_R1192_U74 = ~new_U3078 | ~new_R1192_U75;
  assign new_R1192_U75 = ~new_U3504;
  assign new_R1192_U76 = ~new_U3079;
  assign new_R1192_U77 = ~new_U3066;
  assign new_R1192_U78 = ~new_U3500;
  assign new_R1192_U79 = ~new_U3498;
  assign new_R1192_U80 = ~new_U3496;
  assign new_R1192_U81 = ~new_U3494;
  assign new_R1192_U82 = ~new_U3077;
  assign new_R1192_U83 = ~new_U3492;
  assign new_R1192_U84 = ~new_U3490;
  assign new_R1192_U85 = ~new_U3060;
  assign new_R1192_U86 = ~new_U3059;
  assign new_R1192_U87 = ~new_U3488;
  assign new_R1192_U88 = ~new_U3486;
  assign new_R1192_U89 = ~new_U3080 | ~new_R1192_U53;
  assign new_R1192_U90 = ~new_U3069;
  assign new_R1192_U91 = ~new_R1192_U347 | ~new_R1192_U271;
  assign new_R1192_U92 = ~new_U3070;
  assign new_R1192_U93 = ~new_U3071;
  assign new_R1192_U94 = ~new_U3076;
  assign new_R1192_U95 = ~new_U3076 | ~new_R1192_U81;
  assign new_R1192_U96 = ~new_R1192_U281 | ~new_R1192_U279;
  assign new_R1192_U97 = ~new_U3502;
  assign new_R1192_U98 = ~new_U3054;
  assign new_R1192_U99 = ~new_U3054 | ~new_R1192_U58;
  assign new_R1192_U100 = ~new_U3050;
  assign new_R1192_U101 = ~new_U4029;
  assign new_R1192_U102 = ~new_U3051;
  assign new_R1192_U103 = ~new_R1192_U356 | ~new_R1192_U302;
  assign new_R1192_U104 = ~new_R1192_U354 | ~new_R1192_U300;
  assign new_R1192_U105 = ~new_R1192_U352 | ~new_R1192_U292;
  assign new_R1192_U106 = ~new_U4035 | ~new_R1192_U65;
  assign new_R1192_U107 = ~new_R1192_U95 | ~new_R1192_U321;
  assign new_R1192_U108 = ~new_R1192_U372 | ~new_R1192_U89;
  assign new_R1192_U109 = ~new_U3074;
  assign new_R1192_U110 = ~new_R1192_U433 | ~new_R1192_U432;
  assign new_R1192_U111 = ~new_R1192_U449 | ~new_R1192_U448;
  assign new_R1192_U112 = ~new_R1192_U454 | ~new_R1192_U453;
  assign new_R1192_U113 = ~new_R1192_U472 | ~new_R1192_U471;
  assign new_R1192_U114 = ~new_R1192_U477 | ~new_R1192_U476;
  assign new_R1192_U115 = ~new_R1192_U482 | ~new_R1192_U481;
  assign new_R1192_U116 = ~new_R1192_U487 | ~new_R1192_U486;
  assign new_R1192_U117 = ~new_R1192_U492 | ~new_R1192_U491;
  assign new_R1192_U118 = ~new_R1192_U508 | ~new_R1192_U507;
  assign new_R1192_U119 = ~new_R1192_U513 | ~new_R1192_U512;
  assign new_R1192_U120 = ~new_R1192_U392 | ~new_R1192_U391;
  assign new_R1192_U121 = ~new_R1192_U401 | ~new_R1192_U400;
  assign new_R1192_U122 = ~new_R1192_U408 | ~new_R1192_U407;
  assign new_R1192_U123 = ~new_R1192_U412 | ~new_R1192_U411;
  assign new_R1192_U124 = ~new_R1192_U421 | ~new_R1192_U420;
  assign new_R1192_U125 = ~new_R1192_U444 | ~new_R1192_U443;
  assign new_R1192_U126 = ~new_R1192_U463 | ~new_R1192_U462;
  assign new_R1192_U127 = ~new_R1192_U467 | ~new_R1192_U466;
  assign new_R1192_U128 = ~new_R1192_U499 | ~new_R1192_U498;
  assign new_R1192_U129 = ~new_R1192_U503 | ~new_R1192_U502;
  assign new_R1192_U130 = ~new_R1192_U520 | ~new_R1192_U519;
  assign new_R1192_U131 = new_R1192_U225 & new_R1192_U215;
  assign new_R1192_U132 = new_R1192_U228 & new_R1192_U227;
  assign new_R1192_U133 = new_R1192_U14 & new_R1192_U13;
  assign new_R1192_U134 = new_R1192_U242 & new_R1192_U241;
  assign new_R1192_U135 = new_R1192_U346 & new_R1192_U134;
  assign new_R1192_U136 = new_R1192_U34 & new_R1192_U394 & new_R1192_U393;
  assign new_R1192_U137 = new_R1192_U397 & new_R1192_U217;
  assign new_R1192_U138 = new_R1192_U257 & new_R1192_U6;
  assign new_R1192_U139 = new_R1192_U404 & new_R1192_U216;
  assign new_R1192_U140 = new_R1192_U42 & new_R1192_U414 & new_R1192_U413;
  assign new_R1192_U141 = new_R1192_U417 & new_R1192_U215;
  assign new_R1192_U142 = new_R1192_U273 & new_R1192_U18;
  assign new_R1192_U143 = new_R1192_U16 & new_R1192_U285;
  assign new_R1192_U144 = new_R1192_U351 & new_R1192_U286;
  assign new_R1192_U145 = new_R1192_U21 & new_R1192_U303;
  assign new_R1192_U146 = new_R1192_U358 & new_R1192_U304;
  assign new_R1192_U147 = new_R1192_U305 & new_R1192_U214;
  assign new_R1192_U148 = new_R1192_U308 & new_R1192_U309;
  assign new_R1192_U149 = new_R1192_U311 & new_R1192_U426;
  assign new_R1192_U150 = new_R1192_U308 & new_R1192_U309;
  assign new_R1192_U151 = new_R1192_U23 & new_R1192_U312;
  assign new_R1192_U152 = ~new_R1192_U430 | ~new_R1192_U429;
  assign new_R1192_U153 = new_R1192_U436 & new_R1192_U214;
  assign new_R1192_U154 = new_R1192_U214 & new_R1192_U186;
  assign new_R1192_U155 = ~new_R1192_U446 | ~new_R1192_U445;
  assign new_R1192_U156 = ~new_R1192_U451 | ~new_R1192_U450;
  assign new_R1192_U157 = new_R1192_U22 & new_R1192_U298;
  assign new_R1192_U158 = new_R1192_U213 & new_R1192_U317;
  assign new_R1192_U159 = new_U3058 & new_R1192_U68;
  assign new_R1192_U160 = new_R1192_U19 & new_R1192_U298;
  assign new_R1192_U161 = new_R1192_U12 & new_R1192_U360 & new_R1192_U317;
  assign new_R1192_U162 = ~new_R1192_U469 | ~new_R1192_U468;
  assign new_R1192_U163 = ~new_R1192_U474 | ~new_R1192_U473;
  assign new_R1192_U164 = ~new_R1192_U479 | ~new_R1192_U478;
  assign new_R1192_U165 = ~new_R1192_U484 | ~new_R1192_U483;
  assign new_R1192_U166 = ~new_R1192_U489 | ~new_R1192_U488;
  assign new_R1192_U167 = new_R1192_U327 & new_R1192_U10;
  assign new_R1192_U168 = new_R1192_U495 & new_R1192_U212;
  assign new_R1192_U169 = ~new_R1192_U505 | ~new_R1192_U504;
  assign new_R1192_U170 = ~new_R1192_U510 | ~new_R1192_U509;
  assign new_R1192_U171 = new_R1192_U336 & new_R1192_U8;
  assign new_R1192_U172 = new_R1192_U516 & new_R1192_U211;
  assign new_R1192_U173 = new_R1192_U390 & new_R1192_U389;
  assign new_R1192_U174 = ~new_R1192_U135 | ~new_R1192_U345;
  assign new_R1192_U175 = new_R1192_U399 & new_R1192_U398;
  assign new_R1192_U176 = new_R1192_U406 & new_R1192_U405;
  assign new_R1192_U177 = new_R1192_U410 & new_R1192_U409;
  assign new_R1192_U178 = ~new_R1192_U132 | ~new_R1192_U380;
  assign new_R1192_U179 = new_R1192_U419 & new_R1192_U418;
  assign new_R1192_U180 = ~new_U4040;
  assign new_R1192_U181 = ~new_U3052;
  assign new_R1192_U182 = new_R1192_U428 & new_R1192_U427;
  assign new_R1192_U183 = ~new_R1192_U148 | ~new_R1192_U306;
  assign new_R1192_U184 = new_R1192_U440 & new_R1192_U439;
  assign new_R1192_U185 = new_R1192_U442 & new_R1192_U441;
  assign new_R1192_U186 = ~new_R1192_U146 | ~new_R1192_U370;
  assign new_R1192_U187 = ~new_R1192_U357 | ~new_R1192_U367;
  assign new_R1192_U188 = ~new_R1192_U355 | ~new_R1192_U365;
  assign new_R1192_U189 = new_R1192_U461 & new_R1192_U460;
  assign new_R1192_U190 = ~new_R1192_U69 | ~new_R1192_U315;
  assign new_R1192_U191 = new_R1192_U465 & new_R1192_U464;
  assign new_R1192_U192 = ~new_R1192_U353 | ~new_R1192_U363;
  assign new_R1192_U193 = ~new_R1192_U361 | ~new_R1192_U74;
  assign new_R1192_U194 = ~new_U3468;
  assign new_R1192_U195 = ~new_U3464 | ~new_R1192_U109;
  assign new_R1192_U196 = ~new_R1192_U385 | ~new_R1192_U342;
  assign new_R1192_U197 = ~new_R1192_U144 | ~new_R1192_U350;
  assign new_R1192_U198 = ~new_R1192_U96 | ~new_R1192_U282;
  assign new_R1192_U199 = new_R1192_U497 & new_R1192_U496;
  assign new_R1192_U200 = new_R1192_U501 & new_R1192_U500;
  assign new_R1192_U201 = ~new_R1192_U378 | ~new_R1192_U349 | ~new_R1192_U274;
  assign new_R1192_U202 = ~new_R1192_U376 | ~new_R1192_U91;
  assign new_R1192_U203 = ~new_R1192_U374 | ~new_R1192_U270;
  assign new_R1192_U204 = new_R1192_U518 & new_R1192_U517;
  assign new_R1192_U205 = ~new_R1192_U153 | ~new_R1192_U186;
  assign new_R1192_U206 = ~new_R1192_U149 | ~new_R1192_U183;
  assign new_R1192_U207 = ~new_R1192_U195 | ~new_R1192_U194;
  assign new_R1192_U208 = ~new_R1192_U99;
  assign new_R1192_U209 = ~new_R1192_U42;
  assign new_R1192_U210 = ~new_R1192_U34;
  assign new_R1192_U211 = ~new_U3486 | ~new_R1192_U86;
  assign new_R1192_U212 = ~new_U3496 | ~new_R1192_U93;
  assign new_R1192_U213 = ~new_R1192_U106;
  assign new_R1192_U214 = ~new_U4031 | ~new_R1192_U98;
  assign new_R1192_U215 = ~new_U3470 | ~new_R1192_U41;
  assign new_R1192_U216 = ~new_U3476 | ~new_R1192_U49;
  assign new_R1192_U217 = ~new_U3480 | ~new_R1192_U33;
  assign new_R1192_U218 = ~new_R1192_U95;
  assign new_R1192_U219 = ~new_R1192_U69;
  assign new_R1192_U220 = ~new_R1192_U51;
  assign new_R1192_U221 = ~new_R1192_U89;
  assign new_R1192_U222 = ~new_R1192_U195;
  assign new_R1192_U223 = ~new_U3075 | ~new_R1192_U195;
  assign new_R1192_U224 = ~new_R1192_U57;
  assign new_R1192_U225 = ~new_U3472 | ~new_R1192_U43;
  assign new_R1192_U226 = ~new_R1192_U43 | ~new_R1192_U42;
  assign new_R1192_U227 = ~new_R1192_U226 | ~new_R1192_U47;
  assign new_R1192_U228 = ~new_U3061 | ~new_R1192_U209;
  assign new_R1192_U229 = ~new_U3478 | ~new_R1192_U48;
  assign new_R1192_U230 = ~new_U3068 | ~new_R1192_U37;
  assign new_R1192_U231 = ~new_U3064 | ~new_R1192_U36;
  assign new_R1192_U232 = ~new_R1192_U220 | ~new_R1192_U216;
  assign new_R1192_U233 = ~new_R1192_U6 | ~new_R1192_U232;
  assign new_R1192_U234 = ~new_U3474 | ~new_R1192_U50;
  assign new_R1192_U235 = ~new_U3478 | ~new_R1192_U48;
  assign new_R1192_U236 = ~new_R1192_U13 | ~new_R1192_U178;
  assign new_R1192_U237 = ~new_R1192_U52;
  assign new_R1192_U238 = ~new_R1192_U55;
  assign new_R1192_U239 = ~new_U3482 | ~new_R1192_U35;
  assign new_R1192_U240 = ~new_R1192_U35 | ~new_R1192_U34;
  assign new_R1192_U241 = ~new_R1192_U240 | ~new_R1192_U40;
  assign new_R1192_U242 = ~new_U3081 | ~new_R1192_U210;
  assign new_R1192_U243 = ~new_R1192_U174;
  assign new_R1192_U244 = ~new_U3484 | ~new_R1192_U54;
  assign new_R1192_U245 = ~new_R1192_U244 | ~new_R1192_U89;
  assign new_R1192_U246 = ~new_R1192_U238 | ~new_R1192_U34;
  assign new_R1192_U247 = ~new_R1192_U137 | ~new_R1192_U246;
  assign new_R1192_U248 = ~new_R1192_U55 | ~new_R1192_U217;
  assign new_R1192_U249 = ~new_R1192_U136 | ~new_R1192_U248;
  assign new_R1192_U250 = ~new_R1192_U34 | ~new_R1192_U217;
  assign new_R1192_U251 = ~new_R1192_U234 | ~new_R1192_U178;
  assign new_R1192_U252 = ~new_R1192_U56;
  assign new_R1192_U253 = ~new_U3064 | ~new_R1192_U36;
  assign new_R1192_U254 = ~new_R1192_U252 | ~new_R1192_U253;
  assign new_R1192_U255 = ~new_R1192_U139 | ~new_R1192_U254;
  assign new_R1192_U256 = ~new_R1192_U56 | ~new_R1192_U216;
  assign new_R1192_U257 = ~new_U3478 | ~new_R1192_U48;
  assign new_R1192_U258 = ~new_R1192_U138 | ~new_R1192_U256;
  assign new_R1192_U259 = ~new_U3064 | ~new_R1192_U36;
  assign new_R1192_U260 = ~new_R1192_U216 | ~new_R1192_U259;
  assign new_R1192_U261 = ~new_R1192_U234 | ~new_R1192_U51;
  assign new_R1192_U262 = ~new_R1192_U141 | ~new_R1192_U384;
  assign new_R1192_U263 = ~new_R1192_U42 | ~new_R1192_U215;
  assign new_R1192_U264 = ~new_U3488 | ~new_R1192_U85;
  assign new_R1192_U265 = ~new_U3060 | ~new_R1192_U87;
  assign new_R1192_U266 = ~new_U3059 | ~new_R1192_U88;
  assign new_R1192_U267 = ~new_R1192_U221 | ~new_R1192_U7;
  assign new_R1192_U268 = ~new_R1192_U8 | ~new_R1192_U267;
  assign new_R1192_U269 = ~new_U3488 | ~new_R1192_U85;
  assign new_R1192_U270 = ~new_R1192_U269 | ~new_R1192_U268;
  assign new_R1192_U271 = ~new_U3490 | ~new_R1192_U90;
  assign new_R1192_U272 = ~new_U3069 | ~new_R1192_U84;
  assign new_R1192_U273 = ~new_U3492 | ~new_R1192_U82;
  assign new_R1192_U274 = ~new_U3077 | ~new_R1192_U83;
  assign new_R1192_U275 = ~new_U3498 | ~new_R1192_U92;
  assign new_R1192_U276 = ~new_U3070 | ~new_R1192_U79;
  assign new_R1192_U277 = ~new_U3071 | ~new_R1192_U80;
  assign new_R1192_U278 = ~new_R1192_U218 | ~new_R1192_U9;
  assign new_R1192_U279 = ~new_R1192_U10 | ~new_R1192_U278;
  assign new_R1192_U280 = ~new_U3494 | ~new_R1192_U94;
  assign new_R1192_U281 = ~new_U3498 | ~new_R1192_U92;
  assign new_R1192_U282 = ~new_R1192_U16 | ~new_R1192_U201;
  assign new_R1192_U283 = ~new_R1192_U96;
  assign new_R1192_U284 = ~new_R1192_U198;
  assign new_R1192_U285 = ~new_U3500 | ~new_R1192_U77;
  assign new_R1192_U286 = ~new_U3066 | ~new_R1192_U78;
  assign new_R1192_U287 = ~new_R1192_U197;
  assign new_R1192_U288 = ~new_U3502 | ~new_R1192_U76;
  assign new_R1192_U289 = ~new_U3504 | ~new_R1192_U72;
  assign new_R1192_U290 = ~new_R1192_U74;
  assign new_R1192_U291 = ~new_U4037 | ~new_R1192_U71;
  assign new_R1192_U292 = ~new_U3073 | ~new_R1192_U73;
  assign new_R1192_U293 = ~new_U4034 | ~new_R1192_U64;
  assign new_R1192_U294 = ~new_U3063 | ~new_R1192_U67;
  assign new_R1192_U295 = ~new_U3058 | ~new_R1192_U68;
  assign new_R1192_U296 = ~new_R1192_U219 | ~new_R1192_U11;
  assign new_R1192_U297 = ~new_R1192_U12 | ~new_R1192_U296;
  assign new_R1192_U298 = ~new_U4036 | ~new_R1192_U66;
  assign new_R1192_U299 = ~new_U4034 | ~new_R1192_U64;
  assign new_R1192_U300 = ~new_R1192_U299 | ~new_R1192_U297;
  assign new_R1192_U301 = ~new_U4033 | ~new_R1192_U62;
  assign new_R1192_U302 = ~new_U3062 | ~new_R1192_U63;
  assign new_R1192_U303 = ~new_U4032 | ~new_R1192_U60;
  assign new_R1192_U304 = ~new_U3055 | ~new_R1192_U61;
  assign new_R1192_U305 = ~new_U4030 | ~new_R1192_U100;
  assign new_R1192_U306 = ~new_R1192_U147 | ~new_R1192_U186;
  assign new_R1192_U307 = ~new_R1192_U100 | ~new_R1192_U99;
  assign new_R1192_U308 = ~new_R1192_U307 | ~new_R1192_U59;
  assign new_R1192_U309 = ~new_U3050 | ~new_R1192_U208;
  assign new_R1192_U310 = ~new_R1192_U183;
  assign new_R1192_U311 = ~new_U4029 | ~new_R1192_U102;
  assign new_R1192_U312 = ~new_U3051 | ~new_R1192_U101;
  assign new_R1192_U313 = ~new_R1192_U154 | ~new_R1192_U205;
  assign new_R1192_U314 = ~new_R1192_U99 | ~new_R1192_U214;
  assign new_R1192_U315 = ~new_R1192_U298 | ~new_R1192_U192;
  assign new_R1192_U316 = ~new_R1192_U190;
  assign new_R1192_U317 = ~new_U4034 | ~new_R1192_U64;
  assign new_R1192_U318 = ~new_U3058 | ~new_R1192_U68;
  assign new_R1192_U319 = ~new_R1192_U106 | ~new_R1192_U318;
  assign new_R1192_U320 = ~new_R1192_U298 | ~new_R1192_U69;
  assign new_R1192_U321 = ~new_R1192_U280 | ~new_R1192_U201;
  assign new_R1192_U322 = ~new_R1192_U107;
  assign new_R1192_U323 = ~new_U3071 | ~new_R1192_U80;
  assign new_R1192_U324 = ~new_R1192_U322 | ~new_R1192_U323;
  assign new_R1192_U325 = ~new_R1192_U168 | ~new_R1192_U324;
  assign new_R1192_U326 = ~new_R1192_U107 | ~new_R1192_U212;
  assign new_R1192_U327 = ~new_U3498 | ~new_R1192_U92;
  assign new_R1192_U328 = ~new_R1192_U167 | ~new_R1192_U326;
  assign new_R1192_U329 = ~new_U3071 | ~new_R1192_U80;
  assign new_R1192_U330 = ~new_R1192_U212 | ~new_R1192_U329;
  assign new_R1192_U331 = ~new_R1192_U280 | ~new_R1192_U95;
  assign new_R1192_U332 = ~new_U3059 | ~new_R1192_U88;
  assign new_R1192_U333 = ~new_R1192_U373 | ~new_R1192_U332;
  assign new_R1192_U334 = ~new_R1192_U172 | ~new_R1192_U333;
  assign new_R1192_U335 = ~new_R1192_U108 | ~new_R1192_U211;
  assign new_R1192_U336 = ~new_U3488 | ~new_R1192_U85;
  assign new_R1192_U337 = ~new_R1192_U171 | ~new_R1192_U335;
  assign new_R1192_U338 = ~new_U3059 | ~new_R1192_U88;
  assign new_R1192_U339 = ~new_R1192_U211 | ~new_R1192_U338;
  assign new_R1192_U340 = ~new_U3074 | ~new_R1192_U45;
  assign new_R1192_U341 = ~new_U3075 | ~new_R1192_U194;
  assign new_R1192_U342 = ~new_U3079 | ~new_R1192_U97;
  assign new_R1192_U343 = ~new_R1192_U151 | ~new_R1192_U150 | ~new_R1192_U306;
  assign new_R1192_U344 = ~new_R1192_U184 | ~new_R1192_U205;
  assign new_R1192_U345 = ~new_R1192_U133 | ~new_R1192_U178;
  assign new_R1192_U346 = ~new_R1192_U237 | ~new_R1192_U14;
  assign new_R1192_U347 = ~new_R1192_U272 | ~new_R1192_U270;
  assign new_R1192_U348 = ~new_R1192_U91;
  assign new_R1192_U349 = ~new_R1192_U348 | ~new_R1192_U273;
  assign new_R1192_U350 = ~new_R1192_U143 | ~new_R1192_U201;
  assign new_R1192_U351 = ~new_R1192_U283 | ~new_R1192_U285;
  assign new_R1192_U352 = ~new_R1192_U290 | ~new_R1192_U291;
  assign new_R1192_U353 = ~new_R1192_U105;
  assign new_R1192_U354 = ~new_R1192_U17 | ~new_R1192_U105;
  assign new_R1192_U355 = ~new_R1192_U104;
  assign new_R1192_U356 = ~new_R1192_U104 | ~new_R1192_U301;
  assign new_R1192_U357 = ~new_R1192_U103;
  assign new_R1192_U358 = ~new_R1192_U103 | ~new_R1192_U303;
  assign new_R1192_U359 = ~new_R1192_U157 | ~new_R1192_U192;
  assign new_R1192_U360 = ~new_R1192_U105 | ~new_R1192_U298;
  assign new_R1192_U361 = ~new_R1192_U289 | ~new_R1192_U196;
  assign new_R1192_U362 = ~new_R1192_U193;
  assign new_R1192_U363 = ~new_R1192_U19 | ~new_R1192_U196;
  assign new_R1192_U364 = ~new_R1192_U192;
  assign new_R1192_U365 = ~new_R1192_U20 | ~new_R1192_U196;
  assign new_R1192_U366 = ~new_R1192_U188;
  assign new_R1192_U367 = ~new_R1192_U21 | ~new_R1192_U196;
  assign new_R1192_U368 = ~new_R1192_U187;
  assign new_R1192_U369 = ~new_R1192_U160 | ~new_R1192_U196;
  assign new_R1192_U370 = ~new_R1192_U145 | ~new_R1192_U196;
  assign new_R1192_U371 = ~new_R1192_U186;
  assign new_R1192_U372 = ~new_R1192_U244 | ~new_R1192_U174;
  assign new_R1192_U373 = ~new_R1192_U108;
  assign new_R1192_U374 = ~new_R1192_U15 | ~new_R1192_U174;
  assign new_R1192_U375 = ~new_R1192_U203;
  assign new_R1192_U376 = ~new_R1192_U18 | ~new_R1192_U174;
  assign new_R1192_U377 = ~new_R1192_U202;
  assign new_R1192_U378 = ~new_R1192_U142 | ~new_R1192_U174;
  assign new_R1192_U379 = ~new_R1192_U201;
  assign new_R1192_U380 = ~new_R1192_U131 | ~new_R1192_U57;
  assign new_R1192_U381 = ~new_R1192_U178;
  assign new_R1192_U382 = ~new_R1192_U215 | ~new_R1192_U57;
  assign new_R1192_U383 = ~new_R1192_U140 | ~new_R1192_U382;
  assign new_R1192_U384 = ~new_R1192_U224 | ~new_R1192_U42;
  assign new_R1192_U385 = ~new_R1192_U288 | ~new_R1192_U197;
  assign new_R1192_U386 = ~new_R1192_U196;
  assign new_R1192_U387 = ~new_R1192_U158 | ~new_R1192_U12;
  assign new_R1192_U388 = ~new_R1192_U159 | ~new_R1192_U457;
  assign new_R1192_U389 = ~new_U3484 | ~new_R1192_U54;
  assign new_R1192_U390 = ~new_U3080 | ~new_R1192_U53;
  assign new_R1192_U391 = ~new_R1192_U245 | ~new_R1192_U174;
  assign new_R1192_U392 = ~new_R1192_U243 | ~new_R1192_U173;
  assign new_R1192_U393 = ~new_U3482 | ~new_R1192_U35;
  assign new_R1192_U394 = ~new_U3081 | ~new_R1192_U40;
  assign new_R1192_U395 = ~new_U3482 | ~new_R1192_U35;
  assign new_R1192_U396 = ~new_U3081 | ~new_R1192_U40;
  assign new_R1192_U397 = ~new_R1192_U396 | ~new_R1192_U395;
  assign new_R1192_U398 = ~new_U3480 | ~new_R1192_U33;
  assign new_R1192_U399 = ~new_U3067 | ~new_R1192_U39;
  assign new_R1192_U400 = ~new_R1192_U250 | ~new_R1192_U55;
  assign new_R1192_U401 = ~new_R1192_U175 | ~new_R1192_U238;
  assign new_R1192_U402 = ~new_U3478 | ~new_R1192_U48;
  assign new_R1192_U403 = ~new_U3068 | ~new_R1192_U37;
  assign new_R1192_U404 = ~new_R1192_U403 | ~new_R1192_U402;
  assign new_R1192_U405 = ~new_U3476 | ~new_R1192_U49;
  assign new_R1192_U406 = ~new_U3064 | ~new_R1192_U36;
  assign new_R1192_U407 = ~new_R1192_U260 | ~new_R1192_U56;
  assign new_R1192_U408 = ~new_R1192_U176 | ~new_R1192_U252;
  assign new_R1192_U409 = ~new_U3474 | ~new_R1192_U50;
  assign new_R1192_U410 = ~new_U3057 | ~new_R1192_U38;
  assign new_R1192_U411 = ~new_R1192_U178 | ~new_R1192_U261;
  assign new_R1192_U412 = ~new_R1192_U381 | ~new_R1192_U177;
  assign new_R1192_U413 = ~new_U3472 | ~new_R1192_U43;
  assign new_R1192_U414 = ~new_U3061 | ~new_R1192_U47;
  assign new_R1192_U415 = ~new_U3472 | ~new_R1192_U43;
  assign new_R1192_U416 = ~new_U3061 | ~new_R1192_U47;
  assign new_R1192_U417 = ~new_R1192_U416 | ~new_R1192_U415;
  assign new_R1192_U418 = ~new_U3470 | ~new_R1192_U41;
  assign new_R1192_U419 = ~new_U3065 | ~new_R1192_U44;
  assign new_R1192_U420 = ~new_R1192_U263 | ~new_R1192_U57;
  assign new_R1192_U421 = ~new_R1192_U179 | ~new_R1192_U224;
  assign new_R1192_U422 = ~new_U4040 | ~new_R1192_U181;
  assign new_R1192_U423 = ~new_U3052 | ~new_R1192_U180;
  assign new_R1192_U424 = ~new_U4040 | ~new_R1192_U181;
  assign new_R1192_U425 = ~new_U3052 | ~new_R1192_U180;
  assign new_R1192_U426 = ~new_R1192_U425 | ~new_R1192_U424;
  assign new_R1192_U427 = ~new_R1192_U102 | ~new_U4029 | ~new_R1192_U23;
  assign new_R1192_U428 = ~new_U3051 | ~new_R1192_U426 | ~new_R1192_U101;
  assign new_R1192_U429 = ~new_U4029 | ~new_R1192_U102;
  assign new_R1192_U430 = ~new_U3051 | ~new_R1192_U101;
  assign new_R1192_U431 = ~new_R1192_U152;
  assign new_R1192_U432 = ~new_R1192_U310 | ~new_R1192_U431;
  assign new_R1192_U433 = ~new_R1192_U152 | ~new_R1192_U183;
  assign new_R1192_U434 = ~new_U4030 | ~new_R1192_U100;
  assign new_R1192_U435 = ~new_U3050 | ~new_R1192_U59;
  assign new_R1192_U436 = ~new_R1192_U435 | ~new_R1192_U434;
  assign new_R1192_U437 = ~new_U4030 | ~new_R1192_U100;
  assign new_R1192_U438 = ~new_U3050 | ~new_R1192_U59;
  assign new_R1192_U439 = ~new_R1192_U99 | ~new_R1192_U438 | ~new_R1192_U437;
  assign new_R1192_U440 = ~new_R1192_U436 | ~new_R1192_U208;
  assign new_R1192_U441 = ~new_U4031 | ~new_R1192_U98;
  assign new_R1192_U442 = ~new_U3054 | ~new_R1192_U58;
  assign new_R1192_U443 = ~new_R1192_U186 | ~new_R1192_U314;
  assign new_R1192_U444 = ~new_R1192_U371 | ~new_R1192_U185;
  assign new_R1192_U445 = ~new_U4032 | ~new_R1192_U60;
  assign new_R1192_U446 = ~new_U3055 | ~new_R1192_U61;
  assign new_R1192_U447 = ~new_R1192_U155;
  assign new_R1192_U448 = ~new_R1192_U368 | ~new_R1192_U447;
  assign new_R1192_U449 = ~new_R1192_U155 | ~new_R1192_U187;
  assign new_R1192_U450 = ~new_U4033 | ~new_R1192_U62;
  assign new_R1192_U451 = ~new_U3062 | ~new_R1192_U63;
  assign new_R1192_U452 = ~new_R1192_U156;
  assign new_R1192_U453 = ~new_R1192_U366 | ~new_R1192_U452;
  assign new_R1192_U454 = ~new_R1192_U156 | ~new_R1192_U188;
  assign new_R1192_U455 = ~new_U4034 | ~new_R1192_U64;
  assign new_R1192_U456 = ~new_U3063 | ~new_R1192_U67;
  assign new_R1192_U457 = ~new_R1192_U456 | ~new_R1192_U455;
  assign new_R1192_U458 = ~new_R1192_U69 | ~new_R1192_U161 | ~new_R1192_U369;
  assign new_R1192_U459 = ~new_R1192_U22 | ~new_R1192_U219;
  assign new_R1192_U460 = ~new_U4035 | ~new_R1192_U65;
  assign new_R1192_U461 = ~new_U3058 | ~new_R1192_U68;
  assign new_R1192_U462 = ~new_R1192_U319 | ~new_R1192_U190;
  assign new_R1192_U463 = ~new_R1192_U316 | ~new_R1192_U189;
  assign new_R1192_U464 = ~new_U4036 | ~new_R1192_U66;
  assign new_R1192_U465 = ~new_U3072 | ~new_R1192_U70;
  assign new_R1192_U466 = ~new_R1192_U192 | ~new_R1192_U320;
  assign new_R1192_U467 = ~new_R1192_U364 | ~new_R1192_U191;
  assign new_R1192_U468 = ~new_U4037 | ~new_R1192_U71;
  assign new_R1192_U469 = ~new_U3073 | ~new_R1192_U73;
  assign new_R1192_U470 = ~new_R1192_U162;
  assign new_R1192_U471 = ~new_R1192_U362 | ~new_R1192_U470;
  assign new_R1192_U472 = ~new_R1192_U162 | ~new_R1192_U193;
  assign new_R1192_U473 = ~new_U3468 | ~new_R1192_U46;
  assign new_R1192_U474 = ~new_U3075 | ~new_R1192_U194;
  assign new_R1192_U475 = ~new_R1192_U163;
  assign new_R1192_U476 = ~new_R1192_U222 | ~new_R1192_U475;
  assign new_R1192_U477 = ~new_R1192_U163 | ~new_R1192_U195;
  assign new_R1192_U478 = ~new_U3504 | ~new_R1192_U72;
  assign new_R1192_U479 = ~new_U3078 | ~new_R1192_U75;
  assign new_R1192_U480 = ~new_R1192_U164;
  assign new_R1192_U481 = ~new_R1192_U386 | ~new_R1192_U480;
  assign new_R1192_U482 = ~new_R1192_U164 | ~new_R1192_U196;
  assign new_R1192_U483 = ~new_U3502 | ~new_R1192_U76;
  assign new_R1192_U484 = ~new_U3079 | ~new_R1192_U97;
  assign new_R1192_U485 = ~new_R1192_U165;
  assign new_R1192_U486 = ~new_R1192_U287 | ~new_R1192_U485;
  assign new_R1192_U487 = ~new_R1192_U165 | ~new_R1192_U197;
  assign new_R1192_U488 = ~new_U3500 | ~new_R1192_U77;
  assign new_R1192_U489 = ~new_U3066 | ~new_R1192_U78;
  assign new_R1192_U490 = ~new_R1192_U166;
  assign new_R1192_U491 = ~new_R1192_U284 | ~new_R1192_U490;
  assign new_R1192_U492 = ~new_R1192_U166 | ~new_R1192_U198;
  assign new_R1192_U493 = ~new_U3498 | ~new_R1192_U92;
  assign new_R1192_U494 = ~new_U3070 | ~new_R1192_U79;
  assign new_R1192_U495 = ~new_R1192_U494 | ~new_R1192_U493;
  assign new_R1192_U496 = ~new_U3496 | ~new_R1192_U93;
  assign new_R1192_U497 = ~new_U3071 | ~new_R1192_U80;
  assign new_R1192_U498 = ~new_R1192_U330 | ~new_R1192_U107;
  assign new_R1192_U499 = ~new_R1192_U199 | ~new_R1192_U322;
  assign new_R1192_U500 = ~new_U3494 | ~new_R1192_U94;
  assign new_R1192_U501 = ~new_U3076 | ~new_R1192_U81;
  assign new_R1192_U502 = ~new_R1192_U201 | ~new_R1192_U331;
  assign new_R1192_U503 = ~new_R1192_U379 | ~new_R1192_U200;
  assign new_R1192_U504 = ~new_U3492 | ~new_R1192_U82;
  assign new_R1192_U505 = ~new_U3077 | ~new_R1192_U83;
  assign new_R1192_U506 = ~new_R1192_U169;
  assign new_R1192_U507 = ~new_R1192_U377 | ~new_R1192_U506;
  assign new_R1192_U508 = ~new_R1192_U169 | ~new_R1192_U202;
  assign new_R1192_U509 = ~new_U3490 | ~new_R1192_U90;
  assign new_R1192_U510 = ~new_U3069 | ~new_R1192_U84;
  assign new_R1192_U511 = ~new_R1192_U170;
  assign new_R1192_U512 = ~new_R1192_U375 | ~new_R1192_U511;
  assign new_R1192_U513 = ~new_R1192_U170 | ~new_R1192_U203;
  assign new_R1192_U514 = ~new_U3488 | ~new_R1192_U85;
  assign new_R1192_U515 = ~new_U3060 | ~new_R1192_U87;
  assign new_R1192_U516 = ~new_R1192_U515 | ~new_R1192_U514;
  assign new_R1192_U517 = ~new_U3486 | ~new_R1192_U86;
  assign new_R1192_U518 = ~new_U3059 | ~new_R1192_U88;
  assign new_R1192_U519 = ~new_R1192_U108 | ~new_R1192_U339;
  assign new_R1192_U520 = ~new_R1192_U204 | ~new_R1192_U373;
  assign new_R1347_U6 = new_R1347_U139 & new_R1347_U141 & new_R1347_U143 & new_R1347_U142;
  assign new_R1347_U7 = new_R1347_U84 & new_R1347_U6;
  assign new_R1347_U8 = new_R1347_U7 & new_R1347_U147;
  assign new_R1347_U9 = new_R1347_U181 & new_R1347_U180;
  assign new_R1347_U10 = new_R1347_U83 & new_R1347_U11;
  assign new_R1347_U11 = new_R1347_U79 & new_R1347_U78 & new_R1347_U183;
  assign new_R1347_U12 = new_R1347_U209 & new_R1347_U132;
  assign new_R1347_U13 = new_R1347_U198 & new_R1347_U118;
  assign new_R1347_U14 = ~new_U3596;
  assign new_R1347_U15 = ~new_U3486;
  assign new_R1347_U16 = ~new_U3484;
  assign new_R1347_U17 = ~new_U3480;
  assign new_R1347_U18 = ~new_U3482;
  assign new_R1347_U19 = ~new_U3478;
  assign new_R1347_U20 = ~new_U3476;
  assign new_R1347_U21 = ~new_U3474;
  assign new_R1347_U22 = ~new_U3472;
  assign new_R1347_U23 = ~new_U3612;
  assign new_R1347_U24 = ~new_U3470;
  assign new_R1347_U25 = ~new_U3468;
  assign new_R1347_U26 = ~new_U3498;
  assign new_R1347_U27 = ~new_U3496;
  assign new_R1347_U28 = ~new_U3608;
  assign new_R1347_U29 = ~new_U3490;
  assign new_R1347_U30 = ~new_U3609;
  assign new_R1347_U31 = ~new_R1347_U153 | ~new_R1347_U152;
  assign new_R1347_U32 = ~new_U3488;
  assign new_R1347_U33 = ~new_U3492;
  assign new_R1347_U34 = ~new_U3494;
  assign new_R1347_U35 = ~new_U4036;
  assign new_R1347_U36 = ~new_U4035;
  assign new_R1347_U37 = ~new_U3602;
  assign new_R1347_U38 = ~new_U3502;
  assign new_R1347_U39 = ~new_U3603;
  assign new_R1347_U40 = ~new_R1347_U135 | ~new_R1347_U136;
  assign new_R1347_U41 = ~new_U3500;
  assign new_R1347_U42 = ~new_U3504;
  assign new_R1347_U43 = ~new_U4037;
  assign new_R1347_U44 = ~new_U3601;
  assign new_R1347_U45 = ~new_U3590;
  assign new_R1347_U46 = ~new_U3587;
  assign new_R1347_U47 = ~new_U3586;
  assign new_R1347_U48 = ~new_U3585;
  assign new_R1347_U49 = ~new_U3584;
  assign new_R1347_U50 = ~new_U3583;
  assign new_R1347_U51 = ~new_U3582;
  assign new_R1347_U52 = ~new_U3611;
  assign new_R1347_U53 = ~new_U3610;
  assign new_R1347_U54 = ~new_U3607;
  assign new_R1347_U55 = ~new_U3606;
  assign new_R1347_U56 = ~new_U3605;
  assign new_R1347_U57 = ~new_U3604;
  assign new_R1347_U58 = ~new_U3600;
  assign new_R1347_U59 = ~new_U3599;
  assign new_R1347_U60 = ~new_U3598;
  assign new_R1347_U61 = ~new_U3597;
  assign new_R1347_U62 = ~new_U4034;
  assign new_R1347_U63 = ~new_U4033;
  assign new_R1347_U64 = ~new_U4031;
  assign new_R1347_U65 = ~new_U4030;
  assign new_R1347_U66 = ~new_U3588;
  assign new_R1347_U67 = ~new_U4039;
  assign new_R1347_U68 = ~new_U3589;
  assign new_R1347_U69 = ~new_U4038;
  assign new_R1347_U70 = ~new_U3592;
  assign new_R1347_U71 = ~new_U3593;
  assign new_R1347_U72 = ~new_U3594;
  assign new_R1347_U73 = new_U3464 & new_R1347_U121;
  assign new_R1347_U74 = new_U3490 & new_R1347_U30;
  assign new_R1347_U75 = new_U3488 & new_R1347_U53;
  assign new_R1347_U76 = new_U3502 & new_R1347_U39;
  assign new_R1347_U77 = new_U3500 & new_R1347_U57;
  assign new_R1347_U78 = new_R1347_U184 & new_R1347_U182;
  assign new_R1347_U79 = new_R1347_U9 & new_R1347_U185;
  assign new_R1347_U80 = new_R1347_U138 & new_R1347_U134;
  assign new_R1347_U81 = new_R1347_U80 & new_R1347_U172;
  assign new_R1347_U82 = new_R1347_U175 & new_R1347_U174;
  assign new_R1347_U83 = new_R1347_U82 & new_R1347_U81 & new_R1347_U173;
  assign new_R1347_U84 = new_R1347_U146 & new_R1347_U145 & new_R1347_U144;
  assign new_R1347_U85 = new_R1347_U149 & new_R1347_U150;
  assign new_R1347_U86 = new_R1347_U85 & new_R1347_U148;
  assign new_R1347_U87 = new_U3590 & new_R1347_U22;
  assign new_R1347_U88 = new_R1347_U7 & new_R1347_U87;
  assign new_R1347_U89 = new_R1347_U145 & new_R1347_U144;
  assign new_R1347_U90 = new_R1347_U162 & new_R1347_U163;
  assign new_R1347_U91 = new_R1347_U6 & new_R1347_U164;
  assign new_R1347_U92 = new_R1347_U141 & new_R1347_U139;
  assign new_R1347_U93 = new_R1347_U92 & new_R1347_U157;
  assign new_R1347_U94 = new_U3611 & new_R1347_U15;
  assign new_R1347_U95 = new_U3610 & new_R1347_U32;
  assign new_R1347_U96 = new_R1347_U138 & new_U3607 & new_R1347_U134 & new_R1347_U34;
  assign new_R1347_U97 = new_U3606 & new_R1347_U27;
  assign new_R1347_U98 = new_R1347_U134 & new_R1347_U97;
  assign new_R1347_U99 = new_U3605 & new_R1347_U26;
  assign new_R1347_U100 = new_U3604 & new_R1347_U41;
  assign new_R1347_U101 = new_U3600 & new_R1347_U43;
  assign new_R1347_U102 = new_U3599 & new_R1347_U35;
  assign new_R1347_U103 = new_R1347_U165 & new_R1347_U151 & new_R1347_U133;
  assign new_R1347_U104 = new_R1347_U167 & new_R1347_U166;
  assign new_R1347_U105 = new_R1347_U168 & new_R1347_U169 & new_R1347_U176 & new_R1347_U170;
  assign new_R1347_U106 = new_R1347_U178 & new_R1347_U177;
  assign new_R1347_U107 = new_R1347_U108 & new_R1347_U179;
  assign new_R1347_U108 = new_R1347_U188 & new_R1347_U186;
  assign new_R1347_U109 = new_R1347_U190 & new_R1347_U189;
  assign new_R1347_U110 = new_R1347_U109 & new_R1347_U206;
  assign new_R1347_U111 = new_R1347_U107 & new_R1347_U106 & new_R1347_U110 & new_R1347_U207;
  assign new_R1347_U112 = new_U4034 & new_R1347_U61;
  assign new_R1347_U113 = new_R1347_U192 & new_R1347_U193;
  assign new_R1347_U114 = new_R1347_U132 & new_R1347_U123;
  assign new_R1347_U115 = new_R1347_U12 & new_R1347_U197;
  assign new_R1347_U116 = new_R1347_U115 & new_R1347_U210;
  assign new_R1347_U117 = new_U3589 & new_R1347_U67;
  assign new_R1347_U118 = new_R1347_U212 & new_R1347_U120;
  assign new_R1347_U119 = new_R1347_U204 & new_R1347_U199 & new_R1347_U201;
  assign new_R1347_U120 = new_R1347_U119 & new_R1347_U205;
  assign new_R1347_U121 = ~new_U3613;
  assign new_R1347_U122 = ~new_U4040;
  assign new_R1347_U123 = ~new_U4029;
  assign new_R1347_U124 = ~new_U3595;
  assign new_R1347_U125 = ~new_R1347_U203 | ~new_R1347_U202;
  assign new_R1347_U126 = ~new_R1347_U208 | ~new_R1347_U131;
  assign new_R1347_U127 = ~new_U4032 | ~new_R1347_U194;
  assign new_R1347_U128 = ~new_U3588 | ~new_R1347_U69;
  assign new_R1347_U129 = ~new_R1347_U128 | ~new_R1347_U130 | ~new_R1347_U122;
  assign new_R1347_U130 = ~new_U4039 | ~new_R1347_U68;
  assign new_R1347_U131 = ~new_R1347_U114 | ~new_R1347_U209;
  assign new_R1347_U132 = ~new_U4030 | ~new_R1347_U71;
  assign new_R1347_U133 = ~new_U3596 | ~new_R1347_U63;
  assign new_R1347_U134 = ~new_U3498 | ~new_R1347_U56;
  assign new_R1347_U135 = ~new_U3602 | ~new_R1347_U42;
  assign new_R1347_U136 = ~new_U3603 | ~new_R1347_U38;
  assign new_R1347_U137 = ~new_R1347_U40;
  assign new_R1347_U138 = ~new_U3496 | ~new_R1347_U55;
  assign new_R1347_U139 = ~new_U3486 | ~new_R1347_U52;
  assign new_R1347_U140 = ~new_U3612 | ~new_R1347_U25;
  assign new_R1347_U141 = ~new_U3484 | ~new_R1347_U51;
  assign new_R1347_U142 = ~new_U3480 | ~new_R1347_U49;
  assign new_R1347_U143 = ~new_U3482 | ~new_R1347_U50;
  assign new_R1347_U144 = ~new_U3478 | ~new_R1347_U48;
  assign new_R1347_U145 = ~new_U3476 | ~new_R1347_U47;
  assign new_R1347_U146 = ~new_U3474 | ~new_R1347_U46;
  assign new_R1347_U147 = ~new_U3472 | ~new_R1347_U45;
  assign new_R1347_U148 = ~new_R1347_U73 | ~new_R1347_U140;
  assign new_R1347_U149 = ~new_U3470 | ~new_R1347_U44;
  assign new_R1347_U150 = ~new_U3468 | ~new_R1347_U23;
  assign new_R1347_U151 = ~new_R1347_U10 | ~new_R1347_U8 | ~new_R1347_U86;
  assign new_R1347_U152 = ~new_U3609 | ~new_R1347_U29;
  assign new_R1347_U153 = ~new_U3608 | ~new_R1347_U33;
  assign new_R1347_U154 = ~new_R1347_U31;
  assign new_R1347_U155 = ~new_U3583 | ~new_R1347_U18;
  assign new_R1347_U156 = ~new_U3582 | ~new_R1347_U16;
  assign new_R1347_U157 = ~new_R1347_U156 | ~new_R1347_U155;
  assign new_R1347_U158 = ~new_U3587 | ~new_R1347_U21;
  assign new_R1347_U159 = ~new_U3586 | ~new_R1347_U20;
  assign new_R1347_U160 = ~new_R1347_U159 | ~new_R1347_U158;
  assign new_R1347_U161 = ~new_R1347_U89 | ~new_R1347_U160;
  assign new_R1347_U162 = ~new_U3585 | ~new_R1347_U19;
  assign new_R1347_U163 = ~new_U3584 | ~new_R1347_U17;
  assign new_R1347_U164 = ~new_R1347_U90 | ~new_R1347_U161;
  assign new_R1347_U165 = ~new_R1347_U24 | ~new_R1347_U10 | ~new_U3601 | ~new_R1347_U8;
  assign new_R1347_U166 = ~new_R1347_U88 | ~new_R1347_U10;
  assign new_R1347_U167 = ~new_R1347_U91 | ~new_R1347_U10;
  assign new_R1347_U168 = ~new_R1347_U93 | ~new_R1347_U10;
  assign new_R1347_U169 = ~new_R1347_U94 | ~new_R1347_U10;
  assign new_R1347_U170 = ~new_R1347_U95 | ~new_R1347_U10;
  assign new_R1347_U171 = ~new_U3608 | ~new_R1347_U33;
  assign new_R1347_U172 = ~new_R1347_U74 | ~new_R1347_U171;
  assign new_R1347_U173 = ~new_R1347_U75 | ~new_R1347_U154;
  assign new_R1347_U174 = ~new_U3492 | ~new_R1347_U28;
  assign new_R1347_U175 = ~new_U3494 | ~new_R1347_U54;
  assign new_R1347_U176 = ~new_R1347_U96 | ~new_R1347_U11;
  assign new_R1347_U177 = ~new_R1347_U98 | ~new_R1347_U11;
  assign new_R1347_U178 = ~new_R1347_U99 | ~new_R1347_U11;
  assign new_R1347_U179 = ~new_R1347_U100 | ~new_R1347_U11;
  assign new_R1347_U180 = ~new_U4036 | ~new_R1347_U59;
  assign new_R1347_U181 = ~new_U4035 | ~new_R1347_U60;
  assign new_R1347_U182 = ~new_R1347_U76 | ~new_R1347_U135;
  assign new_R1347_U183 = ~new_R1347_U77 | ~new_R1347_U137;
  assign new_R1347_U184 = ~new_U3504 | ~new_R1347_U37;
  assign new_R1347_U185 = ~new_U4037 | ~new_R1347_U58;
  assign new_R1347_U186 = ~new_R1347_U101 | ~new_R1347_U9;
  assign new_R1347_U187 = ~new_U4035 | ~new_R1347_U60;
  assign new_R1347_U188 = ~new_R1347_U102 | ~new_R1347_U187;
  assign new_R1347_U189 = ~new_U3598 | ~new_R1347_U36;
  assign new_R1347_U190 = ~new_U3597 | ~new_R1347_U62;
  assign new_R1347_U191 = ~new_R1347_U111 | ~new_R1347_U105 | ~new_R1347_U104 | ~new_R1347_U103;
  assign new_R1347_U192 = ~new_R1347_U112 | ~new_R1347_U133;
  assign new_R1347_U193 = ~new_U4033 | ~new_R1347_U14;
  assign new_R1347_U194 = ~new_R1347_U113 | ~new_R1347_U191;
  assign new_R1347_U195 = ~new_U4032 | ~new_R1347_U124;
  assign new_R1347_U196 = ~new_R1347_U194 | ~new_R1347_U124;
  assign new_R1347_U197 = ~new_U4031 | ~new_R1347_U72;
  assign new_R1347_U198 = ~new_R1347_U196 | ~new_R1347_U116 | ~new_R1347_U195 | ~new_R1347_U127;
  assign new_R1347_U199 = ~new_R1347_U117 | ~new_R1347_U128;
  assign new_R1347_U200 = ~new_U4039 | ~new_R1347_U68;
  assign new_R1347_U201 = ~new_U3591 | ~new_R1347_U128 | ~new_R1347_U200 | ~new_R1347_U122;
  assign new_R1347_U202 = ~new_U3593 | ~new_R1347_U65;
  assign new_R1347_U203 = ~new_U3594 | ~new_R1347_U64;
  assign new_R1347_U204 = ~new_U4038 | ~new_R1347_U66;
  assign new_R1347_U205 = ~new_U3592 | ~new_R1347_U209 | ~new_R1347_U123;
  assign new_R1347_U206 = ~new_R1347_U11 | ~new_R1347_U40;
  assign new_R1347_U207 = ~new_R1347_U10 | ~new_R1347_U31;
  assign new_R1347_U208 = ~new_U3592 | ~new_R1347_U12;
  assign new_R1347_U209 = ~new_R1347_U129 | ~new_R1347_U211;
  assign new_R1347_U210 = ~new_R1347_U131 | ~new_R1347_U70;
  assign new_R1347_U211 = ~new_U3591 | ~new_R1347_U130 | ~new_R1347_U128;
  assign new_R1347_U212 = ~new_R1347_U126 | ~new_R1347_U125;
  assign new_R1171_U4 = new_R1171_U196 & new_R1171_U195;
  assign new_R1171_U5 = new_R1171_U197 & new_R1171_U198;
  assign new_R1171_U6 = new_R1171_U210 & new_R1171_U209;
  assign new_R1171_U7 = new_R1171_U250 & new_R1171_U249;
  assign new_R1171_U8 = new_R1171_U258 & new_R1171_U257;
  assign new_R1171_U9 = new_R1171_U274 & new_R1171_U273;
  assign new_R1171_U10 = new_R1171_U282 & new_R1171_U281;
  assign new_R1171_U11 = new_R1171_U10 & new_R1171_U283;
  assign new_R1171_U12 = new_R1171_U7 & new_R1171_U217;
  assign new_R1171_U13 = new_R1171_U8 & new_R1171_U262;
  assign new_R1171_U14 = new_R1171_U11 & new_R1171_U292;
  assign new_R1171_U15 = new_R1171_U13 & new_R1171_U267;
  assign new_R1171_U16 = new_R1171_U9 & new_R1171_U14;
  assign new_R1171_U17 = new_R1171_U299 & new_R1171_U305;
  assign new_R1171_U18 = new_R1171_U359 & new_R1171_U356;
  assign new_R1171_U19 = new_R1171_U352 & new_R1171_U349;
  assign new_R1171_U20 = new_R1171_U343 & new_R1171_U340;
  assign new_R1171_U21 = new_R1171_U334 & new_R1171_U331;
  assign new_R1171_U22 = new_R1171_U328 & new_R1171_U326;
  assign new_R1171_U23 = new_R1171_U321 & new_R1171_U318;
  assign new_R1171_U24 = new_R1171_U248 & new_R1171_U245;
  assign new_R1171_U25 = new_R1171_U240 & new_R1171_U237;
  assign new_R1171_U26 = new_R1171_U226 & new_R1171_U223;
  assign new_R1171_U27 = ~new_U3470;
  assign new_R1171_U28 = ~new_U3065;
  assign new_R1171_U29 = ~new_U3472;
  assign new_R1171_U30 = ~new_U3061;
  assign new_R1171_U31 = ~new_U3474;
  assign new_R1171_U32 = ~new_U3057;
  assign new_R1171_U33 = ~new_U3064;
  assign new_R1171_U34 = ~new_U3057 | ~new_U3474;
  assign new_R1171_U35 = ~new_U3476;
  assign new_R1171_U36 = ~new_U3468 | ~new_U3075;
  assign new_R1171_U37 = ~new_U3464;
  assign new_R1171_U38 = ~new_U3074;
  assign new_R1171_U39 = ~new_R1171_U131 | ~new_R1171_U200;
  assign new_R1171_U40 = ~new_U3478;
  assign new_R1171_U41 = ~new_U3068;
  assign new_R1171_U42 = ~new_U3067;
  assign new_R1171_U43 = ~new_U3068 | ~new_U3478;
  assign new_R1171_U44 = ~new_U3480;
  assign new_R1171_U45 = ~new_R1171_U214 | ~new_R1171_U213;
  assign new_R1171_U46 = ~new_U3482;
  assign new_R1171_U47 = ~new_U3081;
  assign new_R1171_U48 = ~new_U3080;
  assign new_R1171_U49 = ~new_U3484;
  assign new_R1171_U50 = ~new_R1171_U65 | ~new_R1171_U218;
  assign new_R1171_U51 = ~new_R1171_U133 | ~new_R1171_U132;
  assign new_R1171_U52 = ~new_R1171_U136 | ~new_R1171_U232;
  assign new_R1171_U53 = ~new_R1171_U229 | ~new_R1171_U228;
  assign new_R1171_U54 = ~new_U4030;
  assign new_R1171_U55 = ~new_U3050;
  assign new_R1171_U56 = ~new_U3054;
  assign new_R1171_U57 = ~new_U4031;
  assign new_R1171_U58 = ~new_U4033;
  assign new_R1171_U59 = ~new_U3062;
  assign new_R1171_U60 = ~new_U3062 | ~new_U4033;
  assign new_R1171_U61 = ~new_U4035;
  assign new_R1171_U62 = ~new_U3058;
  assign new_R1171_U63 = ~new_U3496;
  assign new_R1171_U64 = ~new_U3071;
  assign new_R1171_U65 = ~new_U3081 | ~new_U3482;
  assign new_R1171_U66 = ~new_U3486;
  assign new_R1171_U67 = ~new_U3059;
  assign new_R1171_U68 = ~new_U3490;
  assign new_R1171_U69 = ~new_U3069;
  assign new_R1171_U70 = ~new_U3488;
  assign new_R1171_U71 = ~new_U3060;
  assign new_R1171_U72 = ~new_U3060 | ~new_U3488;
  assign new_R1171_U73 = ~new_U3492;
  assign new_R1171_U74 = ~new_U3077;
  assign new_R1171_U75 = ~new_U3494;
  assign new_R1171_U76 = ~new_U3076;
  assign new_R1171_U77 = ~new_R1171_U380 | ~new_R1171_U267;
  assign new_R1171_U78 = ~new_U3504;
  assign new_R1171_U79 = ~new_U3078;
  assign new_R1171_U80 = ~new_U3078 | ~new_U3504;
  assign new_R1171_U81 = ~new_U4037;
  assign new_R1171_U82 = ~new_U3502;
  assign new_R1171_U83 = ~new_U3079;
  assign new_R1171_U84 = ~new_U3079 | ~new_U3502;
  assign new_R1171_U85 = ~new_U4036;
  assign new_R1171_U86 = ~new_U3072;
  assign new_R1171_U87 = ~new_U3498;
  assign new_R1171_U88 = ~new_U3070;
  assign new_R1171_U89 = ~new_U3066;
  assign new_R1171_U90 = ~new_U3070 | ~new_U3498;
  assign new_R1171_U91 = ~new_U3500;
  assign new_R1171_U92 = ~new_U4034;
  assign new_R1171_U93 = ~new_U3063;
  assign new_R1171_U94 = ~new_R1171_U146 | ~new_R1171_U388;
  assign new_R1171_U95 = ~new_U4032;
  assign new_R1171_U96 = ~new_U3055;
  assign new_R1171_U97 = ~new_R1171_U397 | ~new_R1171_U396 | ~new_R1171_U306;
  assign new_R1171_U98 = ~new_U3051;
  assign new_R1171_U99 = ~new_U4029;
  assign new_R1171_U100 = ~new_R1171_U60 | ~new_R1171_U314;
  assign new_R1171_U101 = ~new_R1171_U385 | ~new_R1171_U294;
  assign new_R1171_U102 = ~new_R1171_U278 | ~new_R1171_U277;
  assign new_R1171_U103 = ~new_U3073;
  assign new_R1171_U104 = ~new_R1171_U84 | ~new_R1171_U323;
  assign new_R1171_U105 = ~new_R1171_U382 | ~new_R1171_U383 | ~new_R1171_U271;
  assign new_R1171_U106 = ~new_R1171_U72 | ~new_R1171_U345;
  assign new_R1171_U107 = ~new_R1171_U484 | ~new_R1171_U483;
  assign new_R1171_U108 = ~new_R1171_U531 | ~new_R1171_U530;
  assign new_R1171_U109 = ~new_R1171_U402 | ~new_R1171_U401;
  assign new_R1171_U110 = ~new_R1171_U407 | ~new_R1171_U406;
  assign new_R1171_U111 = ~new_R1171_U414 | ~new_R1171_U413;
  assign new_R1171_U112 = ~new_R1171_U421 | ~new_R1171_U420;
  assign new_R1171_U113 = ~new_R1171_U426 | ~new_R1171_U425;
  assign new_R1171_U114 = ~new_R1171_U435 | ~new_R1171_U434;
  assign new_R1171_U115 = ~new_R1171_U442 | ~new_R1171_U441;
  assign new_R1171_U116 = ~new_R1171_U449 | ~new_R1171_U448;
  assign new_R1171_U117 = ~new_R1171_U456 | ~new_R1171_U455;
  assign new_R1171_U118 = ~new_R1171_U461 | ~new_R1171_U460;
  assign new_R1171_U119 = ~new_R1171_U468 | ~new_R1171_U467;
  assign new_R1171_U120 = ~new_R1171_U475 | ~new_R1171_U474;
  assign new_R1171_U121 = ~new_R1171_U489 | ~new_R1171_U488;
  assign new_R1171_U122 = ~new_R1171_U494 | ~new_R1171_U493;
  assign new_R1171_U123 = ~new_R1171_U501 | ~new_R1171_U500;
  assign new_R1171_U124 = ~new_R1171_U508 | ~new_R1171_U507;
  assign new_R1171_U125 = ~new_R1171_U515 | ~new_R1171_U514;
  assign new_R1171_U126 = ~new_R1171_U522 | ~new_R1171_U521;
  assign new_R1171_U127 = ~new_R1171_U527 | ~new_R1171_U526;
  assign new_R1171_U128 = new_R1171_U129 & new_R1171_U197;
  assign new_R1171_U129 = new_U3065 & new_U3470;
  assign new_R1171_U130 = new_U3472 & new_U3061;
  assign new_R1171_U131 = new_U3464 & new_U3074;
  assign new_R1171_U132 = new_R1171_U203 & new_R1171_U204 & new_R1171_U206;
  assign new_R1171_U133 = new_R1171_U374 & new_R1171_U373 & new_R1171_U207;
  assign new_R1171_U134 = new_R1171_U43 & new_R1171_U409 & new_R1171_U408;
  assign new_R1171_U135 = new_R1171_U225 & new_R1171_U6;
  assign new_R1171_U136 = new_R1171_U233 & new_R1171_U231;
  assign new_R1171_U137 = new_R1171_U34 & new_R1171_U416 & new_R1171_U415;
  assign new_R1171_U138 = new_R1171_U239 & new_R1171_U4;
  assign new_R1171_U139 = new_R1171_U247 & new_R1171_U198;
  assign new_R1171_U140 = new_R1171_U252 & new_R1171_U188;
  assign new_R1171_U141 = new_R1171_U6 & new_R1171_U12;
  assign new_R1171_U142 = new_R1171_U378 & new_R1171_U255;
  assign new_R1171_U143 = new_R1171_U270 & new_R1171_U15;
  assign new_R1171_U144 = new_R1171_U260 & new_R1171_U189;
  assign new_R1171_U145 = new_R1171_U296 & new_R1171_U16;
  assign new_R1171_U146 = new_R1171_U389 & new_R1171_U297;
  assign new_R1171_U147 = new_R1171_U309 & new_R1171_U185;
  assign new_R1171_U148 = new_R1171_U395 & new_R1171_U393 & new_R1171_U310;
  assign new_R1171_U149 = new_R1171_U17 & new_R1171_U185;
  assign new_R1171_U150 = new_R1171_U97 & new_R1171_U304;
  assign new_R1171_U151 = new_R1171_U190 & new_R1171_U451 & new_R1171_U450;
  assign new_R1171_U152 = new_R1171_U320 & new_R1171_U185;
  assign new_R1171_U153 = new_R1171_U176 & new_R1171_U288;
  assign new_R1171_U154 = new_R1171_U80 & new_R1171_U482 & new_R1171_U481;
  assign new_R1171_U155 = new_R1171_U333 & new_R1171_U10;
  assign new_R1171_U156 = new_R1171_U90 & new_R1171_U496 & new_R1171_U495;
  assign new_R1171_U157 = new_R1171_U342 & new_R1171_U9;
  assign new_R1171_U158 = new_R1171_U189 & new_R1171_U517 & new_R1171_U516;
  assign new_R1171_U159 = new_R1171_U351 & new_R1171_U8;
  assign new_R1171_U160 = new_R1171_U188 & new_R1171_U529 & new_R1171_U528;
  assign new_R1171_U161 = new_R1171_U358 & new_R1171_U7;
  assign new_R1171_U162 = ~new_R1171_U375 | ~new_R1171_U215;
  assign new_R1171_U163 = ~new_R1171_U230 | ~new_R1171_U242;
  assign new_R1171_U164 = ~new_U3052;
  assign new_R1171_U165 = ~new_U4040;
  assign new_R1171_U166 = new_R1171_U430 & new_R1171_U429;
  assign new_R1171_U167 = ~new_R1171_U372 | ~new_R1171_U312 | ~new_R1171_U186;
  assign new_R1171_U168 = new_R1171_U437 & new_R1171_U436;
  assign new_R1171_U169 = ~new_R1171_U148 | ~new_R1171_U394;
  assign new_R1171_U170 = new_R1171_U444 & new_R1171_U443;
  assign new_R1171_U171 = ~new_R1171_U150 | ~new_R1171_U307;
  assign new_R1171_U172 = ~new_R1171_U301 | ~new_R1171_U300;
  assign new_R1171_U173 = new_R1171_U463 & new_R1171_U462;
  assign new_R1171_U174 = new_R1171_U470 & new_R1171_U469;
  assign new_R1171_U175 = ~new_R1171_U386 | ~new_R1171_U384;
  assign new_R1171_U176 = new_R1171_U477 & new_R1171_U476;
  assign new_R1171_U177 = ~new_U3074 | ~new_U3464;
  assign new_R1171_U178 = ~new_R1171_U36 | ~new_R1171_U335;
  assign new_R1171_U179 = ~new_R1171_U376 | ~new_R1171_U279;
  assign new_R1171_U180 = new_R1171_U503 & new_R1171_U502;
  assign new_R1171_U181 = ~new_R1171_U77 | ~new_R1171_U379;
  assign new_R1171_U182 = new_R1171_U510 & new_R1171_U509;
  assign new_R1171_U183 = ~new_R1171_U265 | ~new_R1171_U264;
  assign new_R1171_U184 = ~new_R1171_U142 | ~new_R1171_U377;
  assign new_R1171_U185 = ~new_R1171_U391 | ~new_R1171_U390;
  assign new_R1171_U186 = ~new_U3051 | ~new_R1171_U169;
  assign new_R1171_U187 = ~new_R1171_U34;
  assign new_R1171_U188 = ~new_U3484 | ~new_U3080;
  assign new_R1171_U189 = ~new_U3069 | ~new_U3490;
  assign new_R1171_U190 = ~new_U3055 | ~new_U4032;
  assign new_R1171_U191 = ~new_R1171_U72;
  assign new_R1171_U192 = ~new_R1171_U84;
  assign new_R1171_U193 = ~new_R1171_U60;
  assign new_R1171_U194 = ~new_R1171_U65;
  assign new_R1171_U195 = new_U3064 | new_U3476;
  assign new_R1171_U196 = new_U3057 | new_U3474;
  assign new_R1171_U197 = new_U3472 | new_U3061;
  assign new_R1171_U198 = new_U3470 | new_U3065;
  assign new_R1171_U199 = ~new_R1171_U177;
  assign new_R1171_U200 = new_U3468 | new_U3075;
  assign new_R1171_U201 = ~new_R1171_U39;
  assign new_R1171_U202 = ~new_R1171_U36;
  assign new_R1171_U203 = ~new_R1171_U4 | ~new_R1171_U128;
  assign new_R1171_U204 = ~new_R1171_U130 | ~new_R1171_U4;
  assign new_R1171_U205 = ~new_R1171_U35 | ~new_R1171_U34;
  assign new_R1171_U206 = ~new_U3064 | ~new_R1171_U205;
  assign new_R1171_U207 = ~new_U3476 | ~new_R1171_U187;
  assign new_R1171_U208 = ~new_R1171_U51;
  assign new_R1171_U209 = new_U3067 | new_U3480;
  assign new_R1171_U210 = new_U3068 | new_U3478;
  assign new_R1171_U211 = ~new_R1171_U43;
  assign new_R1171_U212 = ~new_R1171_U44 | ~new_R1171_U43;
  assign new_R1171_U213 = ~new_U3067 | ~new_R1171_U212;
  assign new_R1171_U214 = ~new_U3480 | ~new_R1171_U211;
  assign new_R1171_U215 = ~new_R1171_U6 | ~new_R1171_U51;
  assign new_R1171_U216 = ~new_R1171_U162;
  assign new_R1171_U217 = new_U3482 | new_U3081;
  assign new_R1171_U218 = ~new_R1171_U217 | ~new_R1171_U162;
  assign new_R1171_U219 = ~new_R1171_U50;
  assign new_R1171_U220 = new_U3080 | new_U3484;
  assign new_R1171_U221 = new_U3478 | new_U3068;
  assign new_R1171_U222 = ~new_R1171_U221 | ~new_R1171_U51;
  assign new_R1171_U223 = ~new_R1171_U134 | ~new_R1171_U222;
  assign new_R1171_U224 = ~new_R1171_U208 | ~new_R1171_U43;
  assign new_R1171_U225 = ~new_U3480 | ~new_U3067;
  assign new_R1171_U226 = ~new_R1171_U135 | ~new_R1171_U224;
  assign new_R1171_U227 = new_U3068 | new_U3478;
  assign new_R1171_U228 = ~new_R1171_U202 | ~new_R1171_U198;
  assign new_R1171_U229 = ~new_U3065 | ~new_U3470;
  assign new_R1171_U230 = ~new_R1171_U53;
  assign new_R1171_U231 = ~new_R1171_U201 | ~new_R1171_U5;
  assign new_R1171_U232 = ~new_R1171_U53 | ~new_R1171_U197;
  assign new_R1171_U233 = ~new_U3061 | ~new_U3472;
  assign new_R1171_U234 = ~new_R1171_U52;
  assign new_R1171_U235 = new_U3474 | new_U3057;
  assign new_R1171_U236 = ~new_R1171_U235 | ~new_R1171_U52;
  assign new_R1171_U237 = ~new_R1171_U137 | ~new_R1171_U236;
  assign new_R1171_U238 = ~new_R1171_U234 | ~new_R1171_U34;
  assign new_R1171_U239 = ~new_U3476 | ~new_U3064;
  assign new_R1171_U240 = ~new_R1171_U138 | ~new_R1171_U238;
  assign new_R1171_U241 = new_U3057 | new_U3474;
  assign new_R1171_U242 = ~new_R1171_U201 | ~new_R1171_U198;
  assign new_R1171_U243 = ~new_R1171_U163;
  assign new_R1171_U244 = ~new_U3061 | ~new_U3472;
  assign new_R1171_U245 = ~new_R1171_U39 | ~new_R1171_U36 | ~new_R1171_U428 | ~new_R1171_U427;
  assign new_R1171_U246 = ~new_R1171_U36 | ~new_R1171_U39;
  assign new_R1171_U247 = ~new_U3065 | ~new_U3470;
  assign new_R1171_U248 = ~new_R1171_U139 | ~new_R1171_U246;
  assign new_R1171_U249 = new_U3080 | new_U3484;
  assign new_R1171_U250 = new_U3059 | new_U3486;
  assign new_R1171_U251 = ~new_R1171_U194 | ~new_R1171_U7;
  assign new_R1171_U252 = ~new_U3059 | ~new_U3486;
  assign new_R1171_U253 = ~new_R1171_U140 | ~new_R1171_U251;
  assign new_R1171_U254 = new_U3486 | new_U3059;
  assign new_R1171_U255 = ~new_R1171_U254 | ~new_R1171_U253;
  assign new_R1171_U256 = ~new_R1171_U184;
  assign new_R1171_U257 = new_U3077 | new_U3492;
  assign new_R1171_U258 = new_U3069 | new_U3490;
  assign new_R1171_U259 = ~new_R1171_U191 | ~new_R1171_U8;
  assign new_R1171_U260 = ~new_U3077 | ~new_U3492;
  assign new_R1171_U261 = ~new_R1171_U144 | ~new_R1171_U259;
  assign new_R1171_U262 = new_U3488 | new_U3060;
  assign new_R1171_U263 = new_U3492 | new_U3077;
  assign new_R1171_U264 = ~new_R1171_U13 | ~new_R1171_U184;
  assign new_R1171_U265 = ~new_R1171_U263 | ~new_R1171_U261;
  assign new_R1171_U266 = ~new_R1171_U183;
  assign new_R1171_U267 = new_U3494 | new_U3076;
  assign new_R1171_U268 = ~new_U3076 | ~new_U3494;
  assign new_R1171_U269 = ~new_R1171_U181;
  assign new_R1171_U270 = new_U3496 | new_U3071;
  assign new_R1171_U271 = ~new_U3071 | ~new_U3496;
  assign new_R1171_U272 = ~new_R1171_U105;
  assign new_R1171_U273 = new_U3066 | new_U3500;
  assign new_R1171_U274 = new_U3070 | new_U3498;
  assign new_R1171_U275 = ~new_R1171_U90;
  assign new_R1171_U276 = ~new_R1171_U91 | ~new_R1171_U90;
  assign new_R1171_U277 = ~new_U3066 | ~new_R1171_U276;
  assign new_R1171_U278 = ~new_U3500 | ~new_R1171_U275;
  assign new_R1171_U279 = ~new_R1171_U9 | ~new_R1171_U105;
  assign new_R1171_U280 = ~new_R1171_U179;
  assign new_R1171_U281 = new_U3073 | new_U4037;
  assign new_R1171_U282 = new_U3078 | new_U3504;
  assign new_R1171_U283 = new_U3072 | new_U4036;
  assign new_R1171_U284 = ~new_R1171_U80;
  assign new_R1171_U285 = ~new_U4037 | ~new_R1171_U284;
  assign new_R1171_U286 = ~new_R1171_U285 | ~new_R1171_U103;
  assign new_R1171_U287 = ~new_R1171_U80 | ~new_R1171_U81;
  assign new_R1171_U288 = ~new_R1171_U287 | ~new_R1171_U286;
  assign new_R1171_U289 = ~new_R1171_U192 | ~new_R1171_U11;
  assign new_R1171_U290 = ~new_U3072 | ~new_U4036;
  assign new_R1171_U291 = ~new_R1171_U290 | ~new_R1171_U289 | ~new_R1171_U288;
  assign new_R1171_U292 = new_U3502 | new_U3079;
  assign new_R1171_U293 = new_U4036 | new_U3072;
  assign new_R1171_U294 = ~new_R1171_U293 | ~new_R1171_U291;
  assign new_R1171_U295 = ~new_R1171_U175;
  assign new_R1171_U296 = new_U4035 | new_U3058;
  assign new_R1171_U297 = ~new_U3058 | ~new_U4035;
  assign new_R1171_U298 = ~new_R1171_U94;
  assign new_R1171_U299 = new_U4034 | new_U3063;
  assign new_R1171_U300 = ~new_R1171_U299 | ~new_R1171_U94;
  assign new_R1171_U301 = ~new_U3063 | ~new_U4034;
  assign new_R1171_U302 = ~new_R1171_U172;
  assign new_R1171_U303 = new_U3055 | new_U4032;
  assign new_R1171_U304 = ~new_R1171_U193 | ~new_R1171_U185;
  assign new_R1171_U305 = new_U4033 | new_U3062;
  assign new_R1171_U306 = new_U4031 | new_U3054;
  assign new_R1171_U307 = ~new_R1171_U149 | ~new_R1171_U392;
  assign new_R1171_U308 = ~new_R1171_U171;
  assign new_R1171_U309 = new_U4030 | new_U3050;
  assign new_R1171_U310 = ~new_U3050 | ~new_U4030;
  assign new_R1171_U311 = ~new_R1171_U169;
  assign new_R1171_U312 = ~new_U4029 | ~new_R1171_U169;
  assign new_R1171_U313 = ~new_R1171_U167;
  assign new_R1171_U314 = ~new_R1171_U305 | ~new_R1171_U172;
  assign new_R1171_U315 = ~new_R1171_U100;
  assign new_R1171_U316 = new_U4032 | new_U3055;
  assign new_R1171_U317 = ~new_R1171_U316 | ~new_R1171_U100;
  assign new_R1171_U318 = ~new_R1171_U151 | ~new_R1171_U317;
  assign new_R1171_U319 = ~new_R1171_U315 | ~new_R1171_U190;
  assign new_R1171_U320 = ~new_U4031 | ~new_U3054;
  assign new_R1171_U321 = ~new_R1171_U152 | ~new_R1171_U319;
  assign new_R1171_U322 = new_U3055 | new_U4032;
  assign new_R1171_U323 = ~new_R1171_U292 | ~new_R1171_U179;
  assign new_R1171_U324 = ~new_R1171_U104;
  assign new_R1171_U325 = ~new_R1171_U10 | ~new_R1171_U104;
  assign new_R1171_U326 = ~new_R1171_U153 | ~new_R1171_U325;
  assign new_R1171_U327 = ~new_R1171_U325 | ~new_R1171_U288;
  assign new_R1171_U328 = ~new_R1171_U480 | ~new_R1171_U327;
  assign new_R1171_U329 = new_U3504 | new_U3078;
  assign new_R1171_U330 = ~new_R1171_U329 | ~new_R1171_U104;
  assign new_R1171_U331 = ~new_R1171_U154 | ~new_R1171_U330;
  assign new_R1171_U332 = ~new_R1171_U324 | ~new_R1171_U80;
  assign new_R1171_U333 = ~new_U3073 | ~new_U4037;
  assign new_R1171_U334 = ~new_R1171_U155 | ~new_R1171_U332;
  assign new_R1171_U335 = new_U3468 | new_U3075;
  assign new_R1171_U336 = ~new_R1171_U178;
  assign new_R1171_U337 = new_U3078 | new_U3504;
  assign new_R1171_U338 = new_U3498 | new_U3070;
  assign new_R1171_U339 = ~new_R1171_U338 | ~new_R1171_U105;
  assign new_R1171_U340 = ~new_R1171_U156 | ~new_R1171_U339;
  assign new_R1171_U341 = ~new_R1171_U272 | ~new_R1171_U90;
  assign new_R1171_U342 = ~new_U3500 | ~new_U3066;
  assign new_R1171_U343 = ~new_R1171_U157 | ~new_R1171_U341;
  assign new_R1171_U344 = new_U3070 | new_U3498;
  assign new_R1171_U345 = ~new_R1171_U262 | ~new_R1171_U184;
  assign new_R1171_U346 = ~new_R1171_U106;
  assign new_R1171_U347 = new_U3490 | new_U3069;
  assign new_R1171_U348 = ~new_R1171_U347 | ~new_R1171_U106;
  assign new_R1171_U349 = ~new_R1171_U158 | ~new_R1171_U348;
  assign new_R1171_U350 = ~new_R1171_U346 | ~new_R1171_U189;
  assign new_R1171_U351 = ~new_U3077 | ~new_U3492;
  assign new_R1171_U352 = ~new_R1171_U159 | ~new_R1171_U350;
  assign new_R1171_U353 = new_U3069 | new_U3490;
  assign new_R1171_U354 = new_U3484 | new_U3080;
  assign new_R1171_U355 = ~new_R1171_U354 | ~new_R1171_U50;
  assign new_R1171_U356 = ~new_R1171_U160 | ~new_R1171_U355;
  assign new_R1171_U357 = ~new_R1171_U219 | ~new_R1171_U188;
  assign new_R1171_U358 = ~new_U3059 | ~new_U3486;
  assign new_R1171_U359 = ~new_R1171_U161 | ~new_R1171_U357;
  assign new_R1171_U360 = ~new_R1171_U220 | ~new_R1171_U188;
  assign new_R1171_U361 = ~new_R1171_U217 | ~new_R1171_U65;
  assign new_R1171_U362 = ~new_R1171_U227 | ~new_R1171_U43;
  assign new_R1171_U363 = ~new_R1171_U241 | ~new_R1171_U34;
  assign new_R1171_U364 = ~new_R1171_U244 | ~new_R1171_U197;
  assign new_R1171_U365 = ~new_R1171_U322 | ~new_R1171_U190;
  assign new_R1171_U366 = ~new_R1171_U305 | ~new_R1171_U60;
  assign new_R1171_U367 = ~new_R1171_U337 | ~new_R1171_U80;
  assign new_R1171_U368 = ~new_R1171_U292 | ~new_R1171_U84;
  assign new_R1171_U369 = ~new_R1171_U344 | ~new_R1171_U90;
  assign new_R1171_U370 = ~new_R1171_U353 | ~new_R1171_U189;
  assign new_R1171_U371 = ~new_R1171_U262 | ~new_R1171_U72;
  assign new_R1171_U372 = ~new_U4029 | ~new_U3051;
  assign new_R1171_U373 = ~new_R1171_U5 | ~new_R1171_U202 | ~new_R1171_U4;
  assign new_R1171_U374 = ~new_R1171_U201 | ~new_R1171_U5 | ~new_R1171_U4;
  assign new_R1171_U375 = ~new_R1171_U45;
  assign new_R1171_U376 = ~new_R1171_U102;
  assign new_R1171_U377 = ~new_R1171_U141 | ~new_R1171_U51;
  assign new_R1171_U378 = ~new_R1171_U12 | ~new_R1171_U45;
  assign new_R1171_U379 = ~new_R1171_U15 | ~new_R1171_U184;
  assign new_R1171_U380 = ~new_R1171_U268 | ~new_R1171_U265;
  assign new_R1171_U381 = ~new_R1171_U77;
  assign new_R1171_U382 = ~new_R1171_U143 | ~new_R1171_U184;
  assign new_R1171_U383 = ~new_R1171_U381 | ~new_R1171_U270;
  assign new_R1171_U384 = ~new_R1171_U16 | ~new_R1171_U105;
  assign new_R1171_U385 = ~new_R1171_U14 | ~new_R1171_U102;
  assign new_R1171_U386 = ~new_R1171_U101;
  assign new_R1171_U387 = ~new_R1171_U97;
  assign new_R1171_U388 = ~new_R1171_U145 | ~new_R1171_U105;
  assign new_R1171_U389 = ~new_R1171_U101 | ~new_R1171_U296;
  assign new_R1171_U390 = ~new_U3054 | ~new_R1171_U303;
  assign new_R1171_U391 = ~new_U4031 | ~new_R1171_U303;
  assign new_R1171_U392 = ~new_R1171_U298 | ~new_R1171_U301;
  assign new_R1171_U393 = ~new_R1171_U309 | ~new_R1171_U193 | ~new_R1171_U185;
  assign new_R1171_U394 = ~new_R1171_U147 | ~new_R1171_U17 | ~new_R1171_U392;
  assign new_R1171_U395 = ~new_R1171_U387 | ~new_R1171_U309;
  assign new_R1171_U396 = ~new_R1171_U57 | ~new_R1171_U190;
  assign new_R1171_U397 = ~new_R1171_U56 | ~new_R1171_U190;
  assign new_R1171_U398 = ~new_U3080 | ~new_R1171_U49;
  assign new_R1171_U399 = ~new_U3484 | ~new_R1171_U48;
  assign new_R1171_U400 = ~new_R1171_U399 | ~new_R1171_U398;
  assign new_R1171_U401 = ~new_R1171_U360 | ~new_R1171_U50;
  assign new_R1171_U402 = ~new_R1171_U400 | ~new_R1171_U219;
  assign new_R1171_U403 = ~new_U3081 | ~new_R1171_U46;
  assign new_R1171_U404 = ~new_U3482 | ~new_R1171_U47;
  assign new_R1171_U405 = ~new_R1171_U404 | ~new_R1171_U403;
  assign new_R1171_U406 = ~new_R1171_U361 | ~new_R1171_U162;
  assign new_R1171_U407 = ~new_R1171_U216 | ~new_R1171_U405;
  assign new_R1171_U408 = ~new_U3067 | ~new_R1171_U44;
  assign new_R1171_U409 = ~new_U3480 | ~new_R1171_U42;
  assign new_R1171_U410 = ~new_U3068 | ~new_R1171_U40;
  assign new_R1171_U411 = ~new_U3478 | ~new_R1171_U41;
  assign new_R1171_U412 = ~new_R1171_U411 | ~new_R1171_U410;
  assign new_R1171_U413 = ~new_R1171_U362 | ~new_R1171_U51;
  assign new_R1171_U414 = ~new_R1171_U412 | ~new_R1171_U208;
  assign new_R1171_U415 = ~new_U3064 | ~new_R1171_U35;
  assign new_R1171_U416 = ~new_U3476 | ~new_R1171_U33;
  assign new_R1171_U417 = ~new_U3057 | ~new_R1171_U31;
  assign new_R1171_U418 = ~new_U3474 | ~new_R1171_U32;
  assign new_R1171_U419 = ~new_R1171_U418 | ~new_R1171_U417;
  assign new_R1171_U420 = ~new_R1171_U363 | ~new_R1171_U52;
  assign new_R1171_U421 = ~new_R1171_U419 | ~new_R1171_U234;
  assign new_R1171_U422 = ~new_U3061 | ~new_R1171_U29;
  assign new_R1171_U423 = ~new_U3472 | ~new_R1171_U30;
  assign new_R1171_U424 = ~new_R1171_U423 | ~new_R1171_U422;
  assign new_R1171_U425 = ~new_R1171_U364 | ~new_R1171_U163;
  assign new_R1171_U426 = ~new_R1171_U243 | ~new_R1171_U424;
  assign new_R1171_U427 = ~new_U3065 | ~new_R1171_U27;
  assign new_R1171_U428 = ~new_U3470 | ~new_R1171_U28;
  assign new_R1171_U429 = ~new_U3052 | ~new_R1171_U165;
  assign new_R1171_U430 = ~new_U4040 | ~new_R1171_U164;
  assign new_R1171_U431 = ~new_U3052 | ~new_R1171_U165;
  assign new_R1171_U432 = ~new_U4040 | ~new_R1171_U164;
  assign new_R1171_U433 = ~new_R1171_U432 | ~new_R1171_U431;
  assign new_R1171_U434 = ~new_R1171_U166 | ~new_R1171_U167;
  assign new_R1171_U435 = ~new_R1171_U313 | ~new_R1171_U433;
  assign new_R1171_U436 = ~new_U3051 | ~new_R1171_U99;
  assign new_R1171_U437 = ~new_U4029 | ~new_R1171_U98;
  assign new_R1171_U438 = ~new_U3051 | ~new_R1171_U99;
  assign new_R1171_U439 = ~new_U4029 | ~new_R1171_U98;
  assign new_R1171_U440 = ~new_R1171_U439 | ~new_R1171_U438;
  assign new_R1171_U441 = ~new_R1171_U168 | ~new_R1171_U169;
  assign new_R1171_U442 = ~new_R1171_U311 | ~new_R1171_U440;
  assign new_R1171_U443 = ~new_U3050 | ~new_R1171_U54;
  assign new_R1171_U444 = ~new_U4030 | ~new_R1171_U55;
  assign new_R1171_U445 = ~new_U3050 | ~new_R1171_U54;
  assign new_R1171_U446 = ~new_U4030 | ~new_R1171_U55;
  assign new_R1171_U447 = ~new_R1171_U446 | ~new_R1171_U445;
  assign new_R1171_U448 = ~new_R1171_U170 | ~new_R1171_U171;
  assign new_R1171_U449 = ~new_R1171_U308 | ~new_R1171_U447;
  assign new_R1171_U450 = ~new_U3054 | ~new_R1171_U57;
  assign new_R1171_U451 = ~new_U4031 | ~new_R1171_U56;
  assign new_R1171_U452 = ~new_U3055 | ~new_R1171_U95;
  assign new_R1171_U453 = ~new_U4032 | ~new_R1171_U96;
  assign new_R1171_U454 = ~new_R1171_U453 | ~new_R1171_U452;
  assign new_R1171_U455 = ~new_R1171_U365 | ~new_R1171_U100;
  assign new_R1171_U456 = ~new_R1171_U454 | ~new_R1171_U315;
  assign new_R1171_U457 = ~new_U3062 | ~new_R1171_U58;
  assign new_R1171_U458 = ~new_U4033 | ~new_R1171_U59;
  assign new_R1171_U459 = ~new_R1171_U458 | ~new_R1171_U457;
  assign new_R1171_U460 = ~new_R1171_U366 | ~new_R1171_U172;
  assign new_R1171_U461 = ~new_R1171_U302 | ~new_R1171_U459;
  assign new_R1171_U462 = ~new_U3063 | ~new_R1171_U92;
  assign new_R1171_U463 = ~new_U4034 | ~new_R1171_U93;
  assign new_R1171_U464 = ~new_U3063 | ~new_R1171_U92;
  assign new_R1171_U465 = ~new_U4034 | ~new_R1171_U93;
  assign new_R1171_U466 = ~new_R1171_U465 | ~new_R1171_U464;
  assign new_R1171_U467 = ~new_R1171_U173 | ~new_R1171_U94;
  assign new_R1171_U468 = ~new_R1171_U466 | ~new_R1171_U298;
  assign new_R1171_U469 = ~new_U3058 | ~new_R1171_U61;
  assign new_R1171_U470 = ~new_U4035 | ~new_R1171_U62;
  assign new_R1171_U471 = ~new_U3058 | ~new_R1171_U61;
  assign new_R1171_U472 = ~new_U4035 | ~new_R1171_U62;
  assign new_R1171_U473 = ~new_R1171_U472 | ~new_R1171_U471;
  assign new_R1171_U474 = ~new_R1171_U174 | ~new_R1171_U175;
  assign new_R1171_U475 = ~new_R1171_U295 | ~new_R1171_U473;
  assign new_R1171_U476 = ~new_U3072 | ~new_R1171_U85;
  assign new_R1171_U477 = ~new_U4036 | ~new_R1171_U86;
  assign new_R1171_U478 = ~new_U3072 | ~new_R1171_U85;
  assign new_R1171_U479 = ~new_U4036 | ~new_R1171_U86;
  assign new_R1171_U480 = ~new_R1171_U479 | ~new_R1171_U478;
  assign new_R1171_U481 = ~new_U3073 | ~new_R1171_U81;
  assign new_R1171_U482 = ~new_U4037 | ~new_R1171_U103;
  assign new_R1171_U483 = ~new_R1171_U199 | ~new_R1171_U178;
  assign new_R1171_U484 = ~new_R1171_U336 | ~new_R1171_U177;
  assign new_R1171_U485 = ~new_U3078 | ~new_R1171_U78;
  assign new_R1171_U486 = ~new_U3504 | ~new_R1171_U79;
  assign new_R1171_U487 = ~new_R1171_U486 | ~new_R1171_U485;
  assign new_R1171_U488 = ~new_R1171_U367 | ~new_R1171_U104;
  assign new_R1171_U489 = ~new_R1171_U487 | ~new_R1171_U324;
  assign new_R1171_U490 = ~new_U3079 | ~new_R1171_U82;
  assign new_R1171_U491 = ~new_U3502 | ~new_R1171_U83;
  assign new_R1171_U492 = ~new_R1171_U491 | ~new_R1171_U490;
  assign new_R1171_U493 = ~new_R1171_U368 | ~new_R1171_U179;
  assign new_R1171_U494 = ~new_R1171_U280 | ~new_R1171_U492;
  assign new_R1171_U495 = ~new_U3066 | ~new_R1171_U91;
  assign new_R1171_U496 = ~new_U3500 | ~new_R1171_U89;
  assign new_R1171_U497 = ~new_U3070 | ~new_R1171_U87;
  assign new_R1171_U498 = ~new_U3498 | ~new_R1171_U88;
  assign new_R1171_U499 = ~new_R1171_U498 | ~new_R1171_U497;
  assign new_R1171_U500 = ~new_R1171_U369 | ~new_R1171_U105;
  assign new_R1171_U501 = ~new_R1171_U499 | ~new_R1171_U272;
  assign new_R1171_U502 = ~new_U3071 | ~new_R1171_U63;
  assign new_R1171_U503 = ~new_U3496 | ~new_R1171_U64;
  assign new_R1171_U504 = ~new_U3071 | ~new_R1171_U63;
  assign new_R1171_U505 = ~new_U3496 | ~new_R1171_U64;
  assign new_R1171_U506 = ~new_R1171_U505 | ~new_R1171_U504;
  assign new_R1171_U507 = ~new_R1171_U180 | ~new_R1171_U181;
  assign new_R1171_U508 = ~new_R1171_U269 | ~new_R1171_U506;
  assign new_R1171_U509 = ~new_U3076 | ~new_R1171_U75;
  assign new_R1171_U510 = ~new_U3494 | ~new_R1171_U76;
  assign new_R1171_U511 = ~new_U3076 | ~new_R1171_U75;
  assign new_R1171_U512 = ~new_U3494 | ~new_R1171_U76;
  assign new_R1171_U513 = ~new_R1171_U512 | ~new_R1171_U511;
  assign new_R1171_U514 = ~new_R1171_U182 | ~new_R1171_U183;
  assign new_R1171_U515 = ~new_R1171_U266 | ~new_R1171_U513;
  assign new_R1171_U516 = ~new_U3077 | ~new_R1171_U73;
  assign new_R1171_U517 = ~new_U3492 | ~new_R1171_U74;
  assign new_R1171_U518 = ~new_U3069 | ~new_R1171_U68;
  assign new_R1171_U519 = ~new_U3490 | ~new_R1171_U69;
  assign new_R1171_U520 = ~new_R1171_U519 | ~new_R1171_U518;
  assign new_R1171_U521 = ~new_R1171_U370 | ~new_R1171_U106;
  assign new_R1171_U522 = ~new_R1171_U520 | ~new_R1171_U346;
  assign new_R1171_U523 = ~new_U3060 | ~new_R1171_U70;
  assign new_R1171_U524 = ~new_U3488 | ~new_R1171_U71;
  assign new_R1171_U525 = ~new_R1171_U524 | ~new_R1171_U523;
  assign new_R1171_U526 = ~new_R1171_U371 | ~new_R1171_U184;
  assign new_R1171_U527 = ~new_R1171_U256 | ~new_R1171_U525;
  assign new_R1171_U528 = ~new_U3059 | ~new_R1171_U66;
  assign new_R1171_U529 = ~new_U3486 | ~new_R1171_U67;
  assign new_R1171_U530 = ~new_U3074 | ~new_R1171_U37;
  assign new_R1171_U531 = ~new_U3464 | ~new_R1171_U38;
  assign new_R1138_U4 = new_R1138_U196 & new_R1138_U195;
  assign new_R1138_U5 = new_R1138_U197 & new_R1138_U198;
  assign new_R1138_U6 = new_R1138_U210 & new_R1138_U209;
  assign new_R1138_U7 = new_R1138_U250 & new_R1138_U249;
  assign new_R1138_U8 = new_R1138_U258 & new_R1138_U257;
  assign new_R1138_U9 = new_R1138_U274 & new_R1138_U273;
  assign new_R1138_U10 = new_R1138_U282 & new_R1138_U281;
  assign new_R1138_U11 = new_R1138_U10 & new_R1138_U283;
  assign new_R1138_U12 = new_R1138_U7 & new_R1138_U217;
  assign new_R1138_U13 = new_R1138_U8 & new_R1138_U262;
  assign new_R1138_U14 = new_R1138_U11 & new_R1138_U292;
  assign new_R1138_U15 = new_R1138_U13 & new_R1138_U267;
  assign new_R1138_U16 = new_R1138_U9 & new_R1138_U14;
  assign new_R1138_U17 = new_R1138_U299 & new_R1138_U305;
  assign new_R1138_U18 = new_R1138_U359 & new_R1138_U356;
  assign new_R1138_U19 = new_R1138_U352 & new_R1138_U349;
  assign new_R1138_U20 = new_R1138_U343 & new_R1138_U340;
  assign new_R1138_U21 = new_R1138_U334 & new_R1138_U331;
  assign new_R1138_U22 = new_R1138_U328 & new_R1138_U326;
  assign new_R1138_U23 = new_R1138_U321 & new_R1138_U318;
  assign new_R1138_U24 = new_R1138_U248 & new_R1138_U245;
  assign new_R1138_U25 = new_R1138_U240 & new_R1138_U237;
  assign new_R1138_U26 = new_R1138_U226 & new_R1138_U223;
  assign new_R1138_U27 = ~new_U3470;
  assign new_R1138_U28 = ~new_U3065;
  assign new_R1138_U29 = ~new_U3472;
  assign new_R1138_U30 = ~new_U3061;
  assign new_R1138_U31 = ~new_U3474;
  assign new_R1138_U32 = ~new_U3057;
  assign new_R1138_U33 = ~new_U3064;
  assign new_R1138_U34 = ~new_U3057 | ~new_U3474;
  assign new_R1138_U35 = ~new_U3476;
  assign new_R1138_U36 = ~new_U3468 | ~new_U3075;
  assign new_R1138_U37 = ~new_U3464;
  assign new_R1138_U38 = ~new_U3074;
  assign new_R1138_U39 = ~new_R1138_U131 | ~new_R1138_U200;
  assign new_R1138_U40 = ~new_U3478;
  assign new_R1138_U41 = ~new_U3068;
  assign new_R1138_U42 = ~new_U3067;
  assign new_R1138_U43 = ~new_U3068 | ~new_U3478;
  assign new_R1138_U44 = ~new_U3480;
  assign new_R1138_U45 = ~new_R1138_U214 | ~new_R1138_U213;
  assign new_R1138_U46 = ~new_U3482;
  assign new_R1138_U47 = ~new_U3081;
  assign new_R1138_U48 = ~new_U3080;
  assign new_R1138_U49 = ~new_U3484;
  assign new_R1138_U50 = ~new_R1138_U65 | ~new_R1138_U218;
  assign new_R1138_U51 = ~new_R1138_U133 | ~new_R1138_U132;
  assign new_R1138_U52 = ~new_R1138_U136 | ~new_R1138_U232;
  assign new_R1138_U53 = ~new_R1138_U229 | ~new_R1138_U228;
  assign new_R1138_U54 = ~new_U4030;
  assign new_R1138_U55 = ~new_U3050;
  assign new_R1138_U56 = ~new_U3054;
  assign new_R1138_U57 = ~new_U4031;
  assign new_R1138_U58 = ~new_U4033;
  assign new_R1138_U59 = ~new_U3062;
  assign new_R1138_U60 = ~new_U3062 | ~new_U4033;
  assign new_R1138_U61 = ~new_U4035;
  assign new_R1138_U62 = ~new_U3058;
  assign new_R1138_U63 = ~new_U3496;
  assign new_R1138_U64 = ~new_U3071;
  assign new_R1138_U65 = ~new_U3081 | ~new_U3482;
  assign new_R1138_U66 = ~new_U3486;
  assign new_R1138_U67 = ~new_U3059;
  assign new_R1138_U68 = ~new_U3490;
  assign new_R1138_U69 = ~new_U3069;
  assign new_R1138_U70 = ~new_U3488;
  assign new_R1138_U71 = ~new_U3060;
  assign new_R1138_U72 = ~new_U3060 | ~new_U3488;
  assign new_R1138_U73 = ~new_U3492;
  assign new_R1138_U74 = ~new_U3077;
  assign new_R1138_U75 = ~new_U3494;
  assign new_R1138_U76 = ~new_U3076;
  assign new_R1138_U77 = ~new_R1138_U380 | ~new_R1138_U267;
  assign new_R1138_U78 = ~new_U3504;
  assign new_R1138_U79 = ~new_U3078;
  assign new_R1138_U80 = ~new_U3078 | ~new_U3504;
  assign new_R1138_U81 = ~new_U4037;
  assign new_R1138_U82 = ~new_U3502;
  assign new_R1138_U83 = ~new_U3079;
  assign new_R1138_U84 = ~new_U3079 | ~new_U3502;
  assign new_R1138_U85 = ~new_U4036;
  assign new_R1138_U86 = ~new_U3072;
  assign new_R1138_U87 = ~new_U3498;
  assign new_R1138_U88 = ~new_U3070;
  assign new_R1138_U89 = ~new_U3066;
  assign new_R1138_U90 = ~new_U3070 | ~new_U3498;
  assign new_R1138_U91 = ~new_U3500;
  assign new_R1138_U92 = ~new_U4034;
  assign new_R1138_U93 = ~new_U3063;
  assign new_R1138_U94 = ~new_R1138_U146 | ~new_R1138_U388;
  assign new_R1138_U95 = ~new_U4032;
  assign new_R1138_U96 = ~new_U3055;
  assign new_R1138_U97 = ~new_R1138_U397 | ~new_R1138_U396 | ~new_R1138_U306;
  assign new_R1138_U98 = ~new_U3051;
  assign new_R1138_U99 = ~new_U4029;
  assign new_R1138_U100 = ~new_R1138_U60 | ~new_R1138_U314;
  assign new_R1138_U101 = ~new_R1138_U385 | ~new_R1138_U294;
  assign new_R1138_U102 = ~new_R1138_U278 | ~new_R1138_U277;
  assign new_R1138_U103 = ~new_U3073;
  assign new_R1138_U104 = ~new_R1138_U84 | ~new_R1138_U323;
  assign new_R1138_U105 = ~new_R1138_U382 | ~new_R1138_U383 | ~new_R1138_U271;
  assign new_R1138_U106 = ~new_R1138_U72 | ~new_R1138_U345;
  assign new_R1138_U107 = ~new_R1138_U484 | ~new_R1138_U483;
  assign new_R1138_U108 = ~new_R1138_U531 | ~new_R1138_U530;
  assign new_R1138_U109 = ~new_R1138_U402 | ~new_R1138_U401;
  assign new_R1138_U110 = ~new_R1138_U407 | ~new_R1138_U406;
  assign new_R1138_U111 = ~new_R1138_U414 | ~new_R1138_U413;
  assign new_R1138_U112 = ~new_R1138_U421 | ~new_R1138_U420;
  assign new_R1138_U113 = ~new_R1138_U426 | ~new_R1138_U425;
  assign new_R1138_U114 = ~new_R1138_U435 | ~new_R1138_U434;
  assign new_R1138_U115 = ~new_R1138_U442 | ~new_R1138_U441;
  assign new_R1138_U116 = ~new_R1138_U449 | ~new_R1138_U448;
  assign new_R1138_U117 = ~new_R1138_U456 | ~new_R1138_U455;
  assign new_R1138_U118 = ~new_R1138_U461 | ~new_R1138_U460;
  assign new_R1138_U119 = ~new_R1138_U468 | ~new_R1138_U467;
  assign new_R1138_U120 = ~new_R1138_U475 | ~new_R1138_U474;
  assign new_R1138_U121 = ~new_R1138_U489 | ~new_R1138_U488;
  assign new_R1138_U122 = ~new_R1138_U494 | ~new_R1138_U493;
  assign new_R1138_U123 = ~new_R1138_U501 | ~new_R1138_U500;
  assign new_R1138_U124 = ~new_R1138_U508 | ~new_R1138_U507;
  assign new_R1138_U125 = ~new_R1138_U515 | ~new_R1138_U514;
  assign new_R1138_U126 = ~new_R1138_U522 | ~new_R1138_U521;
  assign new_R1138_U127 = ~new_R1138_U527 | ~new_R1138_U526;
  assign new_R1138_U128 = new_R1138_U129 & new_R1138_U197;
  assign new_R1138_U129 = new_U3065 & new_U3470;
  assign new_R1138_U130 = new_U3472 & new_U3061;
  assign new_R1138_U131 = new_U3464 & new_U3074;
  assign new_R1138_U132 = new_R1138_U203 & new_R1138_U204 & new_R1138_U206;
  assign new_R1138_U133 = new_R1138_U374 & new_R1138_U373 & new_R1138_U207;
  assign new_R1138_U134 = new_R1138_U43 & new_R1138_U409 & new_R1138_U408;
  assign new_R1138_U135 = new_R1138_U225 & new_R1138_U6;
  assign new_R1138_U136 = new_R1138_U233 & new_R1138_U231;
  assign new_R1138_U137 = new_R1138_U34 & new_R1138_U416 & new_R1138_U415;
  assign new_R1138_U138 = new_R1138_U239 & new_R1138_U4;
  assign new_R1138_U139 = new_R1138_U247 & new_R1138_U198;
  assign new_R1138_U140 = new_R1138_U252 & new_R1138_U188;
  assign new_R1138_U141 = new_R1138_U6 & new_R1138_U12;
  assign new_R1138_U142 = new_R1138_U378 & new_R1138_U255;
  assign new_R1138_U143 = new_R1138_U270 & new_R1138_U15;
  assign new_R1138_U144 = new_R1138_U260 & new_R1138_U189;
  assign new_R1138_U145 = new_R1138_U296 & new_R1138_U16;
  assign new_R1138_U146 = new_R1138_U389 & new_R1138_U297;
  assign new_R1138_U147 = new_R1138_U309 & new_R1138_U185;
  assign new_R1138_U148 = new_R1138_U395 & new_R1138_U393 & new_R1138_U310;
  assign new_R1138_U149 = new_R1138_U17 & new_R1138_U185;
  assign new_R1138_U150 = new_R1138_U97 & new_R1138_U304;
  assign new_R1138_U151 = new_R1138_U190 & new_R1138_U451 & new_R1138_U450;
  assign new_R1138_U152 = new_R1138_U320 & new_R1138_U185;
  assign new_R1138_U153 = new_R1138_U176 & new_R1138_U288;
  assign new_R1138_U154 = new_R1138_U80 & new_R1138_U482 & new_R1138_U481;
  assign new_R1138_U155 = new_R1138_U333 & new_R1138_U10;
  assign new_R1138_U156 = new_R1138_U90 & new_R1138_U496 & new_R1138_U495;
  assign new_R1138_U157 = new_R1138_U342 & new_R1138_U9;
  assign new_R1138_U158 = new_R1138_U189 & new_R1138_U517 & new_R1138_U516;
  assign new_R1138_U159 = new_R1138_U351 & new_R1138_U8;
  assign new_R1138_U160 = new_R1138_U188 & new_R1138_U529 & new_R1138_U528;
  assign new_R1138_U161 = new_R1138_U358 & new_R1138_U7;
  assign new_R1138_U162 = ~new_R1138_U375 | ~new_R1138_U215;
  assign new_R1138_U163 = ~new_R1138_U230 | ~new_R1138_U242;
  assign new_R1138_U164 = ~new_U3052;
  assign new_R1138_U165 = ~new_U4040;
  assign new_R1138_U166 = new_R1138_U430 & new_R1138_U429;
  assign new_R1138_U167 = ~new_R1138_U372 | ~new_R1138_U312 | ~new_R1138_U186;
  assign new_R1138_U168 = new_R1138_U437 & new_R1138_U436;
  assign new_R1138_U169 = ~new_R1138_U148 | ~new_R1138_U394;
  assign new_R1138_U170 = new_R1138_U444 & new_R1138_U443;
  assign new_R1138_U171 = ~new_R1138_U150 | ~new_R1138_U307;
  assign new_R1138_U172 = ~new_R1138_U301 | ~new_R1138_U300;
  assign new_R1138_U173 = new_R1138_U463 & new_R1138_U462;
  assign new_R1138_U174 = new_R1138_U470 & new_R1138_U469;
  assign new_R1138_U175 = ~new_R1138_U386 | ~new_R1138_U384;
  assign new_R1138_U176 = new_R1138_U477 & new_R1138_U476;
  assign new_R1138_U177 = ~new_U3074 | ~new_U3464;
  assign new_R1138_U178 = ~new_R1138_U36 | ~new_R1138_U335;
  assign new_R1138_U179 = ~new_R1138_U376 | ~new_R1138_U279;
  assign new_R1138_U180 = new_R1138_U503 & new_R1138_U502;
  assign new_R1138_U181 = ~new_R1138_U77 | ~new_R1138_U379;
  assign new_R1138_U182 = new_R1138_U510 & new_R1138_U509;
  assign new_R1138_U183 = ~new_R1138_U265 | ~new_R1138_U264;
  assign new_R1138_U184 = ~new_R1138_U142 | ~new_R1138_U377;
  assign new_R1138_U185 = ~new_R1138_U391 | ~new_R1138_U390;
  assign new_R1138_U186 = ~new_U3051 | ~new_R1138_U169;
  assign new_R1138_U187 = ~new_R1138_U34;
  assign new_R1138_U188 = ~new_U3484 | ~new_U3080;
  assign new_R1138_U189 = ~new_U3069 | ~new_U3490;
  assign new_R1138_U190 = ~new_U3055 | ~new_U4032;
  assign new_R1138_U191 = ~new_R1138_U72;
  assign new_R1138_U192 = ~new_R1138_U84;
  assign new_R1138_U193 = ~new_R1138_U60;
  assign new_R1138_U194 = ~new_R1138_U65;
  assign new_R1138_U195 = new_U3064 | new_U3476;
  assign new_R1138_U196 = new_U3057 | new_U3474;
  assign new_R1138_U197 = new_U3472 | new_U3061;
  assign new_R1138_U198 = new_U3470 | new_U3065;
  assign new_R1138_U199 = ~new_R1138_U177;
  assign new_R1138_U200 = new_U3468 | new_U3075;
  assign new_R1138_U201 = ~new_R1138_U39;
  assign new_R1138_U202 = ~new_R1138_U36;
  assign new_R1138_U203 = ~new_R1138_U4 | ~new_R1138_U128;
  assign new_R1138_U204 = ~new_R1138_U130 | ~new_R1138_U4;
  assign new_R1138_U205 = ~new_R1138_U35 | ~new_R1138_U34;
  assign new_R1138_U206 = ~new_U3064 | ~new_R1138_U205;
  assign new_R1138_U207 = ~new_U3476 | ~new_R1138_U187;
  assign new_R1138_U208 = ~new_R1138_U51;
  assign new_R1138_U209 = new_U3067 | new_U3480;
  assign new_R1138_U210 = new_U3068 | new_U3478;
  assign new_R1138_U211 = ~new_R1138_U43;
  assign new_R1138_U212 = ~new_R1138_U44 | ~new_R1138_U43;
  assign new_R1138_U213 = ~new_U3067 | ~new_R1138_U212;
  assign new_R1138_U214 = ~new_U3480 | ~new_R1138_U211;
  assign new_R1138_U215 = ~new_R1138_U6 | ~new_R1138_U51;
  assign new_R1138_U216 = ~new_R1138_U162;
  assign new_R1138_U217 = new_U3482 | new_U3081;
  assign new_R1138_U218 = ~new_R1138_U217 | ~new_R1138_U162;
  assign new_R1138_U219 = ~new_R1138_U50;
  assign new_R1138_U220 = new_U3080 | new_U3484;
  assign new_R1138_U221 = new_U3478 | new_U3068;
  assign new_R1138_U222 = ~new_R1138_U221 | ~new_R1138_U51;
  assign new_R1138_U223 = ~new_R1138_U134 | ~new_R1138_U222;
  assign new_R1138_U224 = ~new_R1138_U208 | ~new_R1138_U43;
  assign new_R1138_U225 = ~new_U3480 | ~new_U3067;
  assign new_R1138_U226 = ~new_R1138_U135 | ~new_R1138_U224;
  assign new_R1138_U227 = new_U3068 | new_U3478;
  assign new_R1138_U228 = ~new_R1138_U202 | ~new_R1138_U198;
  assign new_R1138_U229 = ~new_U3065 | ~new_U3470;
  assign new_R1138_U230 = ~new_R1138_U53;
  assign new_R1138_U231 = ~new_R1138_U201 | ~new_R1138_U5;
  assign new_R1138_U232 = ~new_R1138_U53 | ~new_R1138_U197;
  assign new_R1138_U233 = ~new_U3061 | ~new_U3472;
  assign new_R1138_U234 = ~new_R1138_U52;
  assign new_R1138_U235 = new_U3474 | new_U3057;
  assign new_R1138_U236 = ~new_R1138_U235 | ~new_R1138_U52;
  assign new_R1138_U237 = ~new_R1138_U137 | ~new_R1138_U236;
  assign new_R1138_U238 = ~new_R1138_U234 | ~new_R1138_U34;
  assign new_R1138_U239 = ~new_U3476 | ~new_U3064;
  assign new_R1138_U240 = ~new_R1138_U138 | ~new_R1138_U238;
  assign new_R1138_U241 = new_U3057 | new_U3474;
  assign new_R1138_U242 = ~new_R1138_U201 | ~new_R1138_U198;
  assign new_R1138_U243 = ~new_R1138_U163;
  assign new_R1138_U244 = ~new_U3061 | ~new_U3472;
  assign new_R1138_U245 = ~new_R1138_U39 | ~new_R1138_U36 | ~new_R1138_U428 | ~new_R1138_U427;
  assign new_R1138_U246 = ~new_R1138_U36 | ~new_R1138_U39;
  assign new_R1138_U247 = ~new_U3065 | ~new_U3470;
  assign new_R1138_U248 = ~new_R1138_U139 | ~new_R1138_U246;
  assign new_R1138_U249 = new_U3080 | new_U3484;
  assign new_R1138_U250 = new_U3059 | new_U3486;
  assign new_R1138_U251 = ~new_R1138_U194 | ~new_R1138_U7;
  assign new_R1138_U252 = ~new_U3059 | ~new_U3486;
  assign new_R1138_U253 = ~new_R1138_U140 | ~new_R1138_U251;
  assign new_R1138_U254 = new_U3486 | new_U3059;
  assign new_R1138_U255 = ~new_R1138_U254 | ~new_R1138_U253;
  assign new_R1138_U256 = ~new_R1138_U184;
  assign new_R1138_U257 = new_U3077 | new_U3492;
  assign new_R1138_U258 = new_U3069 | new_U3490;
  assign new_R1138_U259 = ~new_R1138_U191 | ~new_R1138_U8;
  assign new_R1138_U260 = ~new_U3077 | ~new_U3492;
  assign new_R1138_U261 = ~new_R1138_U144 | ~new_R1138_U259;
  assign new_R1138_U262 = new_U3488 | new_U3060;
  assign new_R1138_U263 = new_U3492 | new_U3077;
  assign new_R1138_U264 = ~new_R1138_U13 | ~new_R1138_U184;
  assign new_R1138_U265 = ~new_R1138_U263 | ~new_R1138_U261;
  assign new_R1138_U266 = ~new_R1138_U183;
  assign new_R1138_U267 = new_U3494 | new_U3076;
  assign new_R1138_U268 = ~new_U3076 | ~new_U3494;
  assign new_R1138_U269 = ~new_R1138_U181;
  assign new_R1138_U270 = new_U3496 | new_U3071;
  assign new_R1138_U271 = ~new_U3071 | ~new_U3496;
  assign new_R1138_U272 = ~new_R1138_U105;
  assign new_R1138_U273 = new_U3066 | new_U3500;
  assign new_R1138_U274 = new_U3070 | new_U3498;
  assign new_R1138_U275 = ~new_R1138_U90;
  assign new_R1138_U276 = ~new_R1138_U91 | ~new_R1138_U90;
  assign new_R1138_U277 = ~new_U3066 | ~new_R1138_U276;
  assign new_R1138_U278 = ~new_U3500 | ~new_R1138_U275;
  assign new_R1138_U279 = ~new_R1138_U9 | ~new_R1138_U105;
  assign new_R1138_U280 = ~new_R1138_U179;
  assign new_R1138_U281 = new_U3073 | new_U4037;
  assign new_R1138_U282 = new_U3078 | new_U3504;
  assign new_R1138_U283 = new_U3072 | new_U4036;
  assign new_R1138_U284 = ~new_R1138_U80;
  assign new_R1138_U285 = ~new_U4037 | ~new_R1138_U284;
  assign new_R1138_U286 = ~new_R1138_U285 | ~new_R1138_U103;
  assign new_R1138_U287 = ~new_R1138_U80 | ~new_R1138_U81;
  assign new_R1138_U288 = ~new_R1138_U287 | ~new_R1138_U286;
  assign new_R1138_U289 = ~new_R1138_U192 | ~new_R1138_U11;
  assign new_R1138_U290 = ~new_U3072 | ~new_U4036;
  assign new_R1138_U291 = ~new_R1138_U290 | ~new_R1138_U289 | ~new_R1138_U288;
  assign new_R1138_U292 = new_U3502 | new_U3079;
  assign new_R1138_U293 = new_U4036 | new_U3072;
  assign new_R1138_U294 = ~new_R1138_U293 | ~new_R1138_U291;
  assign new_R1138_U295 = ~new_R1138_U175;
  assign new_R1138_U296 = new_U4035 | new_U3058;
  assign new_R1138_U297 = ~new_U3058 | ~new_U4035;
  assign new_R1138_U298 = ~new_R1138_U94;
  assign new_R1138_U299 = new_U4034 | new_U3063;
  assign new_R1138_U300 = ~new_R1138_U299 | ~new_R1138_U94;
  assign new_R1138_U301 = ~new_U3063 | ~new_U4034;
  assign new_R1138_U302 = ~new_R1138_U172;
  assign new_R1138_U303 = new_U3055 | new_U4032;
  assign new_R1138_U304 = ~new_R1138_U193 | ~new_R1138_U185;
  assign new_R1138_U305 = new_U4033 | new_U3062;
  assign new_R1138_U306 = new_U4031 | new_U3054;
  assign new_R1138_U307 = ~new_R1138_U149 | ~new_R1138_U392;
  assign new_R1138_U308 = ~new_R1138_U171;
  assign new_R1138_U309 = new_U4030 | new_U3050;
  assign new_R1138_U310 = ~new_U3050 | ~new_U4030;
  assign new_R1138_U311 = ~new_R1138_U169;
  assign new_R1138_U312 = ~new_U4029 | ~new_R1138_U169;
  assign new_R1138_U313 = ~new_R1138_U167;
  assign new_R1138_U314 = ~new_R1138_U305 | ~new_R1138_U172;
  assign new_R1138_U315 = ~new_R1138_U100;
  assign new_R1138_U316 = new_U4032 | new_U3055;
  assign new_R1138_U317 = ~new_R1138_U316 | ~new_R1138_U100;
  assign new_R1138_U318 = ~new_R1138_U151 | ~new_R1138_U317;
  assign new_R1138_U319 = ~new_R1138_U315 | ~new_R1138_U190;
  assign new_R1138_U320 = ~new_U4031 | ~new_U3054;
  assign new_R1138_U321 = ~new_R1138_U152 | ~new_R1138_U319;
  assign new_R1138_U322 = new_U3055 | new_U4032;
  assign new_R1138_U323 = ~new_R1138_U292 | ~new_R1138_U179;
  assign new_R1138_U324 = ~new_R1138_U104;
  assign new_R1138_U325 = ~new_R1138_U10 | ~new_R1138_U104;
  assign new_R1138_U326 = ~new_R1138_U153 | ~new_R1138_U325;
  assign new_R1138_U327 = ~new_R1138_U325 | ~new_R1138_U288;
  assign new_R1138_U328 = ~new_R1138_U480 | ~new_R1138_U327;
  assign new_R1138_U329 = new_U3504 | new_U3078;
  assign new_R1138_U330 = ~new_R1138_U329 | ~new_R1138_U104;
  assign new_R1138_U331 = ~new_R1138_U154 | ~new_R1138_U330;
  assign new_R1138_U332 = ~new_R1138_U324 | ~new_R1138_U80;
  assign new_R1138_U333 = ~new_U3073 | ~new_U4037;
  assign new_R1138_U334 = ~new_R1138_U155 | ~new_R1138_U332;
  assign new_R1138_U335 = new_U3468 | new_U3075;
  assign new_R1138_U336 = ~new_R1138_U178;
  assign new_R1138_U337 = new_U3078 | new_U3504;
  assign new_R1138_U338 = new_U3498 | new_U3070;
  assign new_R1138_U339 = ~new_R1138_U338 | ~new_R1138_U105;
  assign new_R1138_U340 = ~new_R1138_U156 | ~new_R1138_U339;
  assign new_R1138_U341 = ~new_R1138_U272 | ~new_R1138_U90;
  assign new_R1138_U342 = ~new_U3500 | ~new_U3066;
  assign new_R1138_U343 = ~new_R1138_U157 | ~new_R1138_U341;
  assign new_R1138_U344 = new_U3070 | new_U3498;
  assign new_R1138_U345 = ~new_R1138_U262 | ~new_R1138_U184;
  assign new_R1138_U346 = ~new_R1138_U106;
  assign new_R1138_U347 = new_U3490 | new_U3069;
  assign new_R1138_U348 = ~new_R1138_U347 | ~new_R1138_U106;
  assign new_R1138_U349 = ~new_R1138_U158 | ~new_R1138_U348;
  assign new_R1138_U350 = ~new_R1138_U346 | ~new_R1138_U189;
  assign new_R1138_U351 = ~new_U3077 | ~new_U3492;
  assign new_R1138_U352 = ~new_R1138_U159 | ~new_R1138_U350;
  assign new_R1138_U353 = new_U3069 | new_U3490;
  assign new_R1138_U354 = new_U3484 | new_U3080;
  assign new_R1138_U355 = ~new_R1138_U354 | ~new_R1138_U50;
  assign new_R1138_U356 = ~new_R1138_U160 | ~new_R1138_U355;
  assign new_R1138_U357 = ~new_R1138_U219 | ~new_R1138_U188;
  assign new_R1138_U358 = ~new_U3059 | ~new_U3486;
  assign new_R1138_U359 = ~new_R1138_U161 | ~new_R1138_U357;
  assign new_R1138_U360 = ~new_R1138_U220 | ~new_R1138_U188;
  assign new_R1138_U361 = ~new_R1138_U217 | ~new_R1138_U65;
  assign new_R1138_U362 = ~new_R1138_U227 | ~new_R1138_U43;
  assign new_R1138_U363 = ~new_R1138_U241 | ~new_R1138_U34;
  assign new_R1138_U364 = ~new_R1138_U244 | ~new_R1138_U197;
  assign new_R1138_U365 = ~new_R1138_U322 | ~new_R1138_U190;
  assign new_R1138_U366 = ~new_R1138_U305 | ~new_R1138_U60;
  assign new_R1138_U367 = ~new_R1138_U337 | ~new_R1138_U80;
  assign new_R1138_U368 = ~new_R1138_U292 | ~new_R1138_U84;
  assign new_R1138_U369 = ~new_R1138_U344 | ~new_R1138_U90;
  assign new_R1138_U370 = ~new_R1138_U353 | ~new_R1138_U189;
  assign new_R1138_U371 = ~new_R1138_U262 | ~new_R1138_U72;
  assign new_R1138_U372 = ~new_U4029 | ~new_U3051;
  assign new_R1138_U373 = ~new_R1138_U5 | ~new_R1138_U202 | ~new_R1138_U4;
  assign new_R1138_U374 = ~new_R1138_U201 | ~new_R1138_U5 | ~new_R1138_U4;
  assign new_R1138_U375 = ~new_R1138_U45;
  assign new_R1138_U376 = ~new_R1138_U102;
  assign new_R1138_U377 = ~new_R1138_U141 | ~new_R1138_U51;
  assign new_R1138_U378 = ~new_R1138_U12 | ~new_R1138_U45;
  assign new_R1138_U379 = ~new_R1138_U15 | ~new_R1138_U184;
  assign new_R1138_U380 = ~new_R1138_U268 | ~new_R1138_U265;
  assign new_R1138_U381 = ~new_R1138_U77;
  assign new_R1138_U382 = ~new_R1138_U143 | ~new_R1138_U184;
  assign new_R1138_U383 = ~new_R1138_U381 | ~new_R1138_U270;
  assign new_R1138_U384 = ~new_R1138_U16 | ~new_R1138_U105;
  assign new_R1138_U385 = ~new_R1138_U14 | ~new_R1138_U102;
  assign new_R1138_U386 = ~new_R1138_U101;
  assign new_R1138_U387 = ~new_R1138_U97;
  assign new_R1138_U388 = ~new_R1138_U145 | ~new_R1138_U105;
  assign new_R1138_U389 = ~new_R1138_U101 | ~new_R1138_U296;
  assign new_R1138_U390 = ~new_U3054 | ~new_R1138_U303;
  assign new_R1138_U391 = ~new_U4031 | ~new_R1138_U303;
  assign new_R1138_U392 = ~new_R1138_U298 | ~new_R1138_U301;
  assign new_R1138_U393 = ~new_R1138_U309 | ~new_R1138_U193 | ~new_R1138_U185;
  assign new_R1138_U394 = ~new_R1138_U147 | ~new_R1138_U17 | ~new_R1138_U392;
  assign new_R1138_U395 = ~new_R1138_U387 | ~new_R1138_U309;
  assign new_R1138_U396 = ~new_R1138_U57 | ~new_R1138_U190;
  assign new_R1138_U397 = ~new_R1138_U56 | ~new_R1138_U190;
  assign new_R1138_U398 = ~new_U3080 | ~new_R1138_U49;
  assign new_R1138_U399 = ~new_U3484 | ~new_R1138_U48;
  assign new_R1138_U400 = ~new_R1138_U399 | ~new_R1138_U398;
  assign new_R1138_U401 = ~new_R1138_U360 | ~new_R1138_U50;
  assign new_R1138_U402 = ~new_R1138_U400 | ~new_R1138_U219;
  assign new_R1138_U403 = ~new_U3081 | ~new_R1138_U46;
  assign new_R1138_U404 = ~new_U3482 | ~new_R1138_U47;
  assign new_R1138_U405 = ~new_R1138_U404 | ~new_R1138_U403;
  assign new_R1138_U406 = ~new_R1138_U361 | ~new_R1138_U162;
  assign new_R1138_U407 = ~new_R1138_U216 | ~new_R1138_U405;
  assign new_R1138_U408 = ~new_U3067 | ~new_R1138_U44;
  assign new_R1138_U409 = ~new_U3480 | ~new_R1138_U42;
  assign new_R1138_U410 = ~new_U3068 | ~new_R1138_U40;
  assign new_R1138_U411 = ~new_U3478 | ~new_R1138_U41;
  assign new_R1138_U412 = ~new_R1138_U411 | ~new_R1138_U410;
  assign new_R1138_U413 = ~new_R1138_U362 | ~new_R1138_U51;
  assign new_R1138_U414 = ~new_R1138_U412 | ~new_R1138_U208;
  assign new_R1138_U415 = ~new_U3064 | ~new_R1138_U35;
  assign new_R1138_U416 = ~new_U3476 | ~new_R1138_U33;
  assign new_R1138_U417 = ~new_U3057 | ~new_R1138_U31;
  assign new_R1138_U418 = ~new_U3474 | ~new_R1138_U32;
  assign new_R1138_U419 = ~new_R1138_U418 | ~new_R1138_U417;
  assign new_R1138_U420 = ~new_R1138_U363 | ~new_R1138_U52;
  assign new_R1138_U421 = ~new_R1138_U419 | ~new_R1138_U234;
  assign new_R1138_U422 = ~new_U3061 | ~new_R1138_U29;
  assign new_R1138_U423 = ~new_U3472 | ~new_R1138_U30;
  assign new_R1138_U424 = ~new_R1138_U423 | ~new_R1138_U422;
  assign new_R1138_U425 = ~new_R1138_U364 | ~new_R1138_U163;
  assign new_R1138_U426 = ~new_R1138_U243 | ~new_R1138_U424;
  assign new_R1138_U427 = ~new_U3065 | ~new_R1138_U27;
  assign new_R1138_U428 = ~new_U3470 | ~new_R1138_U28;
  assign new_R1138_U429 = ~new_U3052 | ~new_R1138_U165;
  assign new_R1138_U430 = ~new_U4040 | ~new_R1138_U164;
  assign new_R1138_U431 = ~new_U3052 | ~new_R1138_U165;
  assign new_R1138_U432 = ~new_U4040 | ~new_R1138_U164;
  assign new_R1138_U433 = ~new_R1138_U432 | ~new_R1138_U431;
  assign new_R1138_U434 = ~new_R1138_U166 | ~new_R1138_U167;
  assign new_R1138_U435 = ~new_R1138_U313 | ~new_R1138_U433;
  assign new_R1138_U436 = ~new_U3051 | ~new_R1138_U99;
  assign new_R1138_U437 = ~new_U4029 | ~new_R1138_U98;
  assign new_R1138_U438 = ~new_U3051 | ~new_R1138_U99;
  assign new_R1138_U439 = ~new_U4029 | ~new_R1138_U98;
  assign new_R1138_U440 = ~new_R1138_U439 | ~new_R1138_U438;
  assign new_R1138_U441 = ~new_R1138_U168 | ~new_R1138_U169;
  assign new_R1138_U442 = ~new_R1138_U311 | ~new_R1138_U440;
  assign new_R1138_U443 = ~new_U3050 | ~new_R1138_U54;
  assign new_R1138_U444 = ~new_U4030 | ~new_R1138_U55;
  assign new_R1138_U445 = ~new_U3050 | ~new_R1138_U54;
  assign new_R1138_U446 = ~new_U4030 | ~new_R1138_U55;
  assign new_R1138_U447 = ~new_R1138_U446 | ~new_R1138_U445;
  assign new_R1138_U448 = ~new_R1138_U170 | ~new_R1138_U171;
  assign new_R1138_U449 = ~new_R1138_U308 | ~new_R1138_U447;
  assign new_R1138_U450 = ~new_U3054 | ~new_R1138_U57;
  assign new_R1138_U451 = ~new_U4031 | ~new_R1138_U56;
  assign new_R1138_U452 = ~new_U3055 | ~new_R1138_U95;
  assign new_R1138_U453 = ~new_U4032 | ~new_R1138_U96;
  assign new_R1138_U454 = ~new_R1138_U453 | ~new_R1138_U452;
  assign new_R1138_U455 = ~new_R1138_U365 | ~new_R1138_U100;
  assign new_R1138_U456 = ~new_R1138_U454 | ~new_R1138_U315;
  assign new_R1138_U457 = ~new_U3062 | ~new_R1138_U58;
  assign new_R1138_U458 = ~new_U4033 | ~new_R1138_U59;
  assign new_R1138_U459 = ~new_R1138_U458 | ~new_R1138_U457;
  assign new_R1138_U460 = ~new_R1138_U366 | ~new_R1138_U172;
  assign new_R1138_U461 = ~new_R1138_U302 | ~new_R1138_U459;
  assign new_R1138_U462 = ~new_U3063 | ~new_R1138_U92;
  assign new_R1138_U463 = ~new_U4034 | ~new_R1138_U93;
  assign new_R1138_U464 = ~new_U3063 | ~new_R1138_U92;
  assign new_R1138_U465 = ~new_U4034 | ~new_R1138_U93;
  assign new_R1138_U466 = ~new_R1138_U465 | ~new_R1138_U464;
  assign new_R1138_U467 = ~new_R1138_U173 | ~new_R1138_U94;
  assign new_R1138_U468 = ~new_R1138_U466 | ~new_R1138_U298;
  assign new_R1138_U469 = ~new_U3058 | ~new_R1138_U61;
  assign new_R1138_U470 = ~new_U4035 | ~new_R1138_U62;
  assign new_R1138_U471 = ~new_U3058 | ~new_R1138_U61;
  assign new_R1138_U472 = ~new_U4035 | ~new_R1138_U62;
  assign new_R1138_U473 = ~new_R1138_U472 | ~new_R1138_U471;
  assign new_R1138_U474 = ~new_R1138_U174 | ~new_R1138_U175;
  assign new_R1138_U475 = ~new_R1138_U295 | ~new_R1138_U473;
  assign new_R1138_U476 = ~new_U3072 | ~new_R1138_U85;
  assign new_R1138_U477 = ~new_U4036 | ~new_R1138_U86;
  assign new_R1138_U478 = ~new_U3072 | ~new_R1138_U85;
  assign new_R1138_U479 = ~new_U4036 | ~new_R1138_U86;
  assign new_R1138_U480 = ~new_R1138_U479 | ~new_R1138_U478;
  assign new_R1138_U481 = ~new_U3073 | ~new_R1138_U81;
  assign new_R1138_U482 = ~new_U4037 | ~new_R1138_U103;
  assign new_R1138_U483 = ~new_R1138_U199 | ~new_R1138_U178;
  assign new_R1138_U484 = ~new_R1138_U336 | ~new_R1138_U177;
  assign new_R1138_U485 = ~new_U3078 | ~new_R1138_U78;
  assign new_R1138_U486 = ~new_U3504 | ~new_R1138_U79;
  assign new_R1138_U487 = ~new_R1138_U486 | ~new_R1138_U485;
  assign new_R1138_U488 = ~new_R1138_U367 | ~new_R1138_U104;
  assign new_R1138_U489 = ~new_R1138_U487 | ~new_R1138_U324;
  assign new_R1138_U490 = ~new_U3079 | ~new_R1138_U82;
  assign new_R1138_U491 = ~new_U3502 | ~new_R1138_U83;
  assign new_R1138_U492 = ~new_R1138_U491 | ~new_R1138_U490;
  assign new_R1138_U493 = ~new_R1138_U368 | ~new_R1138_U179;
  assign new_R1138_U494 = ~new_R1138_U280 | ~new_R1138_U492;
  assign new_R1138_U495 = ~new_U3066 | ~new_R1138_U91;
  assign new_R1138_U496 = ~new_U3500 | ~new_R1138_U89;
  assign new_R1138_U497 = ~new_U3070 | ~new_R1138_U87;
  assign new_R1138_U498 = ~new_U3498 | ~new_R1138_U88;
  assign new_R1138_U499 = ~new_R1138_U498 | ~new_R1138_U497;
  assign new_R1138_U500 = ~new_R1138_U369 | ~new_R1138_U105;
  assign new_R1138_U501 = ~new_R1138_U499 | ~new_R1138_U272;
  assign new_R1138_U502 = ~new_U3071 | ~new_R1138_U63;
  assign new_R1138_U503 = ~new_U3496 | ~new_R1138_U64;
  assign new_R1138_U504 = ~new_U3071 | ~new_R1138_U63;
  assign new_R1138_U505 = ~new_U3496 | ~new_R1138_U64;
  assign new_R1138_U506 = ~new_R1138_U505 | ~new_R1138_U504;
  assign new_R1138_U507 = ~new_R1138_U180 | ~new_R1138_U181;
  assign new_R1138_U508 = ~new_R1138_U269 | ~new_R1138_U506;
  assign new_R1138_U509 = ~new_U3076 | ~new_R1138_U75;
  assign new_R1138_U510 = ~new_U3494 | ~new_R1138_U76;
  assign new_R1138_U511 = ~new_U3076 | ~new_R1138_U75;
  assign new_R1138_U512 = ~new_U3494 | ~new_R1138_U76;
  assign new_R1138_U513 = ~new_R1138_U512 | ~new_R1138_U511;
  assign new_R1138_U514 = ~new_R1138_U182 | ~new_R1138_U183;
  assign new_R1138_U515 = ~new_R1138_U266 | ~new_R1138_U513;
  assign new_R1138_U516 = ~new_U3077 | ~new_R1138_U73;
  assign new_R1138_U517 = ~new_U3492 | ~new_R1138_U74;
  assign new_R1138_U518 = ~new_U3069 | ~new_R1138_U68;
  assign new_R1138_U519 = ~new_U3490 | ~new_R1138_U69;
  assign new_R1138_U520 = ~new_R1138_U519 | ~new_R1138_U518;
  assign new_R1138_U521 = ~new_R1138_U370 | ~new_R1138_U106;
  assign new_R1138_U522 = ~new_R1138_U520 | ~new_R1138_U346;
  assign new_R1138_U523 = ~new_U3060 | ~new_R1138_U70;
  assign new_R1138_U524 = ~new_U3488 | ~new_R1138_U71;
  assign new_R1138_U525 = ~new_R1138_U524 | ~new_R1138_U523;
  assign new_R1138_U526 = ~new_R1138_U371 | ~new_R1138_U184;
  assign new_R1138_U527 = ~new_R1138_U256 | ~new_R1138_U525;
  assign new_R1138_U528 = ~new_U3059 | ~new_R1138_U66;
  assign new_R1138_U529 = ~new_U3486 | ~new_R1138_U67;
  assign new_R1138_U530 = ~new_U3074 | ~new_R1138_U37;
  assign new_R1138_U531 = ~new_U3464 | ~new_R1138_U38;
  assign new_R1222_U4 = new_R1222_U190 & new_R1222_U189;
  assign new_R1222_U5 = new_R1222_U191 & new_R1222_U192;
  assign new_R1222_U6 = new_R1222_U204 & new_R1222_U203;
  assign new_R1222_U7 = new_R1222_U239 & new_R1222_U238;
  assign new_R1222_U8 = new_R1222_U246 & new_R1222_U245;
  assign new_R1222_U9 = new_R1222_U262 & new_R1222_U261;
  assign new_R1222_U10 = new_R1222_U268 & new_R1222_U267;
  assign new_R1222_U11 = new_R1222_U10 & new_R1222_U269;
  assign new_R1222_U12 = new_R1222_U290 & new_R1222_U289;
  assign new_R1222_U13 = new_R1222_U7 & new_R1222_U209;
  assign new_R1222_U14 = new_R1222_U8 & new_R1222_U250;
  assign new_R1222_U15 = new_R1222_U11 & new_R1222_U278;
  assign new_R1222_U16 = new_R1222_U14 & new_R1222_U255;
  assign new_R1222_U17 = new_R1222_U347 & new_R1222_U344;
  assign new_R1222_U18 = new_R1222_U340 & new_R1222_U337;
  assign new_R1222_U19 = new_R1222_U331 & new_R1222_U383;
  assign new_R1222_U20 = new_R1222_U325 & new_R1222_U322;
  assign new_R1222_U21 = new_R1222_U319 & new_R1222_U317;
  assign new_R1222_U22 = new_R1222_U312 & new_R1222_U309;
  assign new_R1222_U23 = new_R1222_U237 & new_R1222_U234;
  assign new_R1222_U24 = new_R1222_U229 & new_R1222_U226;
  assign new_R1222_U25 = new_R1222_U215 & new_R1222_U376;
  assign new_R1222_U26 = ~new_U3478;
  assign new_R1222_U27 = ~new_U3068;
  assign new_R1222_U28 = ~new_U3067;
  assign new_R1222_U29 = ~new_U3068 | ~new_U3478;
  assign new_R1222_U30 = ~new_U3480;
  assign new_R1222_U31 = ~new_U3470;
  assign new_R1222_U32 = ~new_U3065;
  assign new_R1222_U33 = ~new_U3472;
  assign new_R1222_U34 = ~new_U3061;
  assign new_R1222_U35 = ~new_U3474;
  assign new_R1222_U36 = ~new_U3057;
  assign new_R1222_U37 = ~new_U3064;
  assign new_R1222_U38 = ~new_U3057 | ~new_U3474;
  assign new_R1222_U39 = ~new_U3476;
  assign new_R1222_U40 = ~new_U3468 | ~new_U3075;
  assign new_R1222_U41 = ~new_U3464;
  assign new_R1222_U42 = ~new_U3074;
  assign new_R1222_U43 = ~new_R1222_U127 | ~new_R1222_U194;
  assign new_R1222_U44 = ~new_R1222_U208 | ~new_R1222_U207;
  assign new_R1222_U45 = ~new_U3482;
  assign new_R1222_U46 = ~new_U3081;
  assign new_R1222_U47 = ~new_U3080;
  assign new_R1222_U48 = ~new_U3484;
  assign new_R1222_U49 = ~new_R1222_U69 | ~new_R1222_U210;
  assign new_R1222_U50 = ~new_R1222_U129 | ~new_R1222_U128;
  assign new_R1222_U51 = ~new_R1222_U132 | ~new_R1222_U221;
  assign new_R1222_U52 = ~new_R1222_U218 | ~new_R1222_U217;
  assign new_R1222_U53 = ~new_U3504;
  assign new_R1222_U54 = ~new_U3078;
  assign new_R1222_U55 = ~new_U3078 | ~new_U3504;
  assign new_R1222_U56 = ~new_U4037;
  assign new_R1222_U57 = ~new_U3502;
  assign new_R1222_U58 = ~new_U3079;
  assign new_R1222_U59 = ~new_U3079 | ~new_U3502;
  assign new_R1222_U60 = ~new_U4036;
  assign new_R1222_U61 = ~new_U3072;
  assign new_R1222_U62 = ~new_U3498;
  assign new_R1222_U63 = ~new_U3070;
  assign new_R1222_U64 = ~new_U3066;
  assign new_R1222_U65 = ~new_U3070 | ~new_U3498;
  assign new_R1222_U66 = ~new_U3500;
  assign new_R1222_U67 = ~new_U3496;
  assign new_R1222_U68 = ~new_U3071;
  assign new_R1222_U69 = ~new_U3081 | ~new_U3482;
  assign new_R1222_U70 = ~new_U3486;
  assign new_R1222_U71 = ~new_U3059;
  assign new_R1222_U72 = ~new_U3490;
  assign new_R1222_U73 = ~new_U3069;
  assign new_R1222_U74 = ~new_U3488;
  assign new_R1222_U75 = ~new_U3060;
  assign new_R1222_U76 = ~new_U3060 | ~new_U3488;
  assign new_R1222_U77 = ~new_U3492;
  assign new_R1222_U78 = ~new_U3077;
  assign new_R1222_U79 = ~new_U3494;
  assign new_R1222_U80 = ~new_U3076;
  assign new_R1222_U81 = ~new_R1222_U367 | ~new_R1222_U255;
  assign new_R1222_U82 = ~new_U4035;
  assign new_R1222_U83 = ~new_U3058;
  assign new_R1222_U84 = ~new_U4034;
  assign new_R1222_U85 = ~new_U3063;
  assign new_R1222_U86 = ~new_U4032;
  assign new_R1222_U87 = ~new_U3055;
  assign new_R1222_U88 = ~new_U4033;
  assign new_R1222_U89 = ~new_U3062;
  assign new_R1222_U90 = ~new_U3062 | ~new_U4033;
  assign new_R1222_U91 = ~new_U4031;
  assign new_R1222_U92 = ~new_U3054;
  assign new_R1222_U93 = ~new_U4030;
  assign new_R1222_U94 = ~new_U3050;
  assign new_R1222_U95 = ~new_U3051;
  assign new_R1222_U96 = ~new_U4029;
  assign new_R1222_U97 = ~new_R1222_U90 | ~new_R1222_U305;
  assign new_R1222_U98 = ~new_R1222_U266 | ~new_R1222_U265;
  assign new_R1222_U99 = ~new_U3073;
  assign new_R1222_U100 = ~new_R1222_U59 | ~new_R1222_U314;
  assign new_R1222_U101 = ~new_R1222_U369 | ~new_R1222_U370 | ~new_R1222_U259;
  assign new_R1222_U102 = ~new_R1222_U76 | ~new_R1222_U333;
  assign new_R1222_U103 = ~new_R1222_U472 | ~new_R1222_U471;
  assign new_R1222_U104 = ~new_R1222_U519 | ~new_R1222_U518;
  assign new_R1222_U105 = ~new_R1222_U390 | ~new_R1222_U389;
  assign new_R1222_U106 = ~new_R1222_U395 | ~new_R1222_U394;
  assign new_R1222_U107 = ~new_R1222_U402 | ~new_R1222_U401;
  assign new_R1222_U108 = ~new_R1222_U409 | ~new_R1222_U408;
  assign new_R1222_U109 = ~new_R1222_U414 | ~new_R1222_U413;
  assign new_R1222_U110 = ~new_R1222_U423 | ~new_R1222_U422;
  assign new_R1222_U111 = ~new_R1222_U430 | ~new_R1222_U429;
  assign new_R1222_U112 = ~new_R1222_U437 | ~new_R1222_U436;
  assign new_R1222_U113 = ~new_R1222_U444 | ~new_R1222_U443;
  assign new_R1222_U114 = ~new_R1222_U449 | ~new_R1222_U448;
  assign new_R1222_U115 = ~new_R1222_U456 | ~new_R1222_U455;
  assign new_R1222_U116 = ~new_R1222_U463 | ~new_R1222_U462;
  assign new_R1222_U117 = ~new_R1222_U477 | ~new_R1222_U476;
  assign new_R1222_U118 = ~new_R1222_U482 | ~new_R1222_U481;
  assign new_R1222_U119 = ~new_R1222_U489 | ~new_R1222_U488;
  assign new_R1222_U120 = ~new_R1222_U496 | ~new_R1222_U495;
  assign new_R1222_U121 = ~new_R1222_U503 | ~new_R1222_U502;
  assign new_R1222_U122 = ~new_R1222_U510 | ~new_R1222_U509;
  assign new_R1222_U123 = ~new_R1222_U515 | ~new_R1222_U514;
  assign new_R1222_U124 = new_R1222_U125 & new_R1222_U191;
  assign new_R1222_U125 = new_U3065 & new_U3470;
  assign new_R1222_U126 = new_U3472 & new_U3061;
  assign new_R1222_U127 = new_U3464 & new_U3074;
  assign new_R1222_U128 = new_R1222_U197 & new_R1222_U198 & new_R1222_U200;
  assign new_R1222_U129 = new_R1222_U362 & new_R1222_U361 & new_R1222_U201;
  assign new_R1222_U130 = new_R1222_U29 & new_R1222_U397 & new_R1222_U396;
  assign new_R1222_U131 = new_R1222_U6 & new_R1222_U214;
  assign new_R1222_U132 = new_R1222_U222 & new_R1222_U220;
  assign new_R1222_U133 = new_R1222_U38 & new_R1222_U404 & new_R1222_U403;
  assign new_R1222_U134 = new_R1222_U228 & new_R1222_U4;
  assign new_R1222_U135 = new_R1222_U236 & new_R1222_U192;
  assign new_R1222_U136 = new_R1222_U241 & new_R1222_U182;
  assign new_R1222_U137 = new_R1222_U6 & new_R1222_U13;
  assign new_R1222_U138 = new_R1222_U365 & new_R1222_U244;
  assign new_R1222_U139 = new_R1222_U16 & new_R1222_U258;
  assign new_R1222_U140 = new_R1222_U248 & new_R1222_U183;
  assign new_R1222_U141 = new_R1222_U15 & new_R1222_U9;
  assign new_R1222_U142 = new_R1222_U371 & new_R1222_U280;
  assign new_R1222_U143 = new_R1222_U294 & new_R1222_U12;
  assign new_R1222_U144 = new_R1222_U292 & new_R1222_U184;
  assign new_R1222_U145 = new_R1222_U184 & new_R1222_U439 & new_R1222_U438;
  assign new_R1222_U146 = new_R1222_U311 & new_R1222_U12;
  assign new_R1222_U147 = new_R1222_U171 & new_R1222_U274;
  assign new_R1222_U148 = new_R1222_U55 & new_R1222_U470 & new_R1222_U469;
  assign new_R1222_U149 = new_R1222_U324 & new_R1222_U10;
  assign new_R1222_U150 = new_R1222_U65 & new_R1222_U484 & new_R1222_U483;
  assign new_R1222_U151 = new_R1222_U9 & new_R1222_U330;
  assign new_R1222_U152 = new_R1222_U183 & new_R1222_U505 & new_R1222_U504;
  assign new_R1222_U153 = new_R1222_U339 & new_R1222_U8;
  assign new_R1222_U154 = new_R1222_U182 & new_R1222_U517 & new_R1222_U516;
  assign new_R1222_U155 = new_R1222_U346 & new_R1222_U7;
  assign new_R1222_U156 = ~new_R1222_U363 | ~new_R1222_U373;
  assign new_R1222_U157 = ~new_R1222_U219 | ~new_R1222_U231;
  assign new_R1222_U158 = ~new_U3052;
  assign new_R1222_U159 = ~new_U4040;
  assign new_R1222_U160 = new_R1222_U418 & new_R1222_U417;
  assign new_R1222_U161 = ~new_R1222_U360 | ~new_R1222_U303 | ~new_R1222_U180;
  assign new_R1222_U162 = new_R1222_U425 & new_R1222_U424;
  assign new_R1222_U163 = ~new_R1222_U301 | ~new_R1222_U300;
  assign new_R1222_U164 = new_R1222_U432 & new_R1222_U431;
  assign new_R1222_U165 = ~new_R1222_U297 | ~new_R1222_U296;
  assign new_R1222_U166 = ~new_R1222_U287 | ~new_R1222_U286;
  assign new_R1222_U167 = new_R1222_U451 & new_R1222_U450;
  assign new_R1222_U168 = ~new_R1222_U283 | ~new_R1222_U282;
  assign new_R1222_U169 = new_R1222_U458 & new_R1222_U457;
  assign new_R1222_U170 = ~new_R1222_U142 | ~new_R1222_U384;
  assign new_R1222_U171 = new_R1222_U465 & new_R1222_U464;
  assign new_R1222_U172 = ~new_U3074 | ~new_U3464;
  assign new_R1222_U173 = ~new_R1222_U40 | ~new_R1222_U326;
  assign new_R1222_U174 = ~new_R1222_U364 | ~new_R1222_U380;
  assign new_R1222_U175 = new_R1222_U491 & new_R1222_U490;
  assign new_R1222_U176 = ~new_R1222_U81 | ~new_R1222_U366;
  assign new_R1222_U177 = new_R1222_U498 & new_R1222_U497;
  assign new_R1222_U178 = ~new_R1222_U253 | ~new_R1222_U252;
  assign new_R1222_U179 = ~new_R1222_U138 | ~new_R1222_U377;
  assign new_R1222_U180 = ~new_U3051 | ~new_R1222_U163;
  assign new_R1222_U181 = ~new_R1222_U38;
  assign new_R1222_U182 = ~new_U3484 | ~new_U3080;
  assign new_R1222_U183 = ~new_U3069 | ~new_U3490;
  assign new_R1222_U184 = ~new_U3055 | ~new_U4032;
  assign new_R1222_U185 = ~new_R1222_U76;
  assign new_R1222_U186 = ~new_R1222_U59;
  assign new_R1222_U187 = ~new_R1222_U90;
  assign new_R1222_U188 = ~new_R1222_U69;
  assign new_R1222_U189 = new_U3064 | new_U3476;
  assign new_R1222_U190 = new_U3057 | new_U3474;
  assign new_R1222_U191 = new_U3472 | new_U3061;
  assign new_R1222_U192 = new_U3470 | new_U3065;
  assign new_R1222_U193 = ~new_R1222_U172;
  assign new_R1222_U194 = new_U3468 | new_U3075;
  assign new_R1222_U195 = ~new_R1222_U43;
  assign new_R1222_U196 = ~new_R1222_U40;
  assign new_R1222_U197 = ~new_R1222_U4 | ~new_R1222_U124;
  assign new_R1222_U198 = ~new_R1222_U126 | ~new_R1222_U4;
  assign new_R1222_U199 = ~new_R1222_U39 | ~new_R1222_U38;
  assign new_R1222_U200 = ~new_U3064 | ~new_R1222_U199;
  assign new_R1222_U201 = ~new_U3476 | ~new_R1222_U181;
  assign new_R1222_U202 = ~new_R1222_U50;
  assign new_R1222_U203 = new_U3067 | new_U3480;
  assign new_R1222_U204 = new_U3068 | new_U3478;
  assign new_R1222_U205 = ~new_R1222_U29;
  assign new_R1222_U206 = ~new_R1222_U30 | ~new_R1222_U29;
  assign new_R1222_U207 = ~new_U3067 | ~new_R1222_U206;
  assign new_R1222_U208 = ~new_U3480 | ~new_R1222_U205;
  assign new_R1222_U209 = new_U3482 | new_U3081;
  assign new_R1222_U210 = ~new_R1222_U209 | ~new_R1222_U156;
  assign new_R1222_U211 = ~new_R1222_U49;
  assign new_R1222_U212 = new_U3080 | new_U3484;
  assign new_R1222_U213 = new_U3478 | new_U3068;
  assign new_R1222_U214 = ~new_U3480 | ~new_U3067;
  assign new_R1222_U215 = ~new_R1222_U131 | ~new_R1222_U372;
  assign new_R1222_U216 = new_U3068 | new_U3478;
  assign new_R1222_U217 = ~new_R1222_U196 | ~new_R1222_U192;
  assign new_R1222_U218 = ~new_U3065 | ~new_U3470;
  assign new_R1222_U219 = ~new_R1222_U52;
  assign new_R1222_U220 = ~new_R1222_U195 | ~new_R1222_U5;
  assign new_R1222_U221 = ~new_R1222_U52 | ~new_R1222_U191;
  assign new_R1222_U222 = ~new_U3061 | ~new_U3472;
  assign new_R1222_U223 = ~new_R1222_U51;
  assign new_R1222_U224 = new_U3474 | new_U3057;
  assign new_R1222_U225 = ~new_R1222_U224 | ~new_R1222_U51;
  assign new_R1222_U226 = ~new_R1222_U133 | ~new_R1222_U225;
  assign new_R1222_U227 = ~new_R1222_U223 | ~new_R1222_U38;
  assign new_R1222_U228 = ~new_U3476 | ~new_U3064;
  assign new_R1222_U229 = ~new_R1222_U134 | ~new_R1222_U227;
  assign new_R1222_U230 = new_U3057 | new_U3474;
  assign new_R1222_U231 = ~new_R1222_U195 | ~new_R1222_U192;
  assign new_R1222_U232 = ~new_R1222_U157;
  assign new_R1222_U233 = ~new_U3061 | ~new_U3472;
  assign new_R1222_U234 = ~new_R1222_U43 | ~new_R1222_U40 | ~new_R1222_U416 | ~new_R1222_U415;
  assign new_R1222_U235 = ~new_R1222_U40 | ~new_R1222_U43;
  assign new_R1222_U236 = ~new_U3065 | ~new_U3470;
  assign new_R1222_U237 = ~new_R1222_U135 | ~new_R1222_U235;
  assign new_R1222_U238 = new_U3080 | new_U3484;
  assign new_R1222_U239 = new_U3059 | new_U3486;
  assign new_R1222_U240 = ~new_R1222_U188 | ~new_R1222_U7;
  assign new_R1222_U241 = ~new_U3059 | ~new_U3486;
  assign new_R1222_U242 = ~new_R1222_U136 | ~new_R1222_U240;
  assign new_R1222_U243 = new_U3486 | new_U3059;
  assign new_R1222_U244 = ~new_R1222_U243 | ~new_R1222_U242;
  assign new_R1222_U245 = new_U3077 | new_U3492;
  assign new_R1222_U246 = new_U3069 | new_U3490;
  assign new_R1222_U247 = ~new_R1222_U185 | ~new_R1222_U8;
  assign new_R1222_U248 = ~new_U3077 | ~new_U3492;
  assign new_R1222_U249 = ~new_R1222_U140 | ~new_R1222_U247;
  assign new_R1222_U250 = new_U3488 | new_U3060;
  assign new_R1222_U251 = new_U3492 | new_U3077;
  assign new_R1222_U252 = ~new_R1222_U14 | ~new_R1222_U179;
  assign new_R1222_U253 = ~new_R1222_U251 | ~new_R1222_U249;
  assign new_R1222_U254 = ~new_R1222_U178;
  assign new_R1222_U255 = new_U3494 | new_U3076;
  assign new_R1222_U256 = ~new_U3076 | ~new_U3494;
  assign new_R1222_U257 = ~new_R1222_U176;
  assign new_R1222_U258 = new_U3496 | new_U3071;
  assign new_R1222_U259 = ~new_U3071 | ~new_U3496;
  assign new_R1222_U260 = ~new_R1222_U101;
  assign new_R1222_U261 = new_U3066 | new_U3500;
  assign new_R1222_U262 = new_U3070 | new_U3498;
  assign new_R1222_U263 = ~new_R1222_U65;
  assign new_R1222_U264 = ~new_R1222_U66 | ~new_R1222_U65;
  assign new_R1222_U265 = ~new_U3066 | ~new_R1222_U264;
  assign new_R1222_U266 = ~new_U3500 | ~new_R1222_U263;
  assign new_R1222_U267 = new_U3073 | new_U4037;
  assign new_R1222_U268 = new_U3078 | new_U3504;
  assign new_R1222_U269 = new_U3072 | new_U4036;
  assign new_R1222_U270 = ~new_R1222_U55;
  assign new_R1222_U271 = ~new_U4037 | ~new_R1222_U270;
  assign new_R1222_U272 = ~new_R1222_U271 | ~new_R1222_U99;
  assign new_R1222_U273 = ~new_R1222_U55 | ~new_R1222_U56;
  assign new_R1222_U274 = ~new_R1222_U273 | ~new_R1222_U272;
  assign new_R1222_U275 = ~new_R1222_U186 | ~new_R1222_U11;
  assign new_R1222_U276 = ~new_U3072 | ~new_U4036;
  assign new_R1222_U277 = ~new_R1222_U276 | ~new_R1222_U275 | ~new_R1222_U274;
  assign new_R1222_U278 = new_U3502 | new_U3079;
  assign new_R1222_U279 = new_U4036 | new_U3072;
  assign new_R1222_U280 = ~new_R1222_U279 | ~new_R1222_U277;
  assign new_R1222_U281 = new_U4035 | new_U3058;
  assign new_R1222_U282 = ~new_R1222_U281 | ~new_R1222_U170;
  assign new_R1222_U283 = ~new_U3058 | ~new_U4035;
  assign new_R1222_U284 = ~new_R1222_U168;
  assign new_R1222_U285 = new_U4034 | new_U3063;
  assign new_R1222_U286 = ~new_R1222_U285 | ~new_R1222_U168;
  assign new_R1222_U287 = ~new_U3063 | ~new_U4034;
  assign new_R1222_U288 = ~new_R1222_U166;
  assign new_R1222_U289 = new_U3054 | new_U4031;
  assign new_R1222_U290 = new_U3055 | new_U4032;
  assign new_R1222_U291 = ~new_R1222_U187 | ~new_R1222_U12;
  assign new_R1222_U292 = ~new_U3054 | ~new_U4031;
  assign new_R1222_U293 = ~new_R1222_U144 | ~new_R1222_U291;
  assign new_R1222_U294 = new_U4033 | new_U3062;
  assign new_R1222_U295 = new_U4031 | new_U3054;
  assign new_R1222_U296 = ~new_R1222_U143 | ~new_R1222_U166;
  assign new_R1222_U297 = ~new_R1222_U295 | ~new_R1222_U293;
  assign new_R1222_U298 = ~new_R1222_U165;
  assign new_R1222_U299 = new_U4030 | new_U3050;
  assign new_R1222_U300 = ~new_R1222_U299 | ~new_R1222_U165;
  assign new_R1222_U301 = ~new_U3050 | ~new_U4030;
  assign new_R1222_U302 = ~new_R1222_U163;
  assign new_R1222_U303 = ~new_U4029 | ~new_R1222_U163;
  assign new_R1222_U304 = ~new_R1222_U161;
  assign new_R1222_U305 = ~new_R1222_U294 | ~new_R1222_U166;
  assign new_R1222_U306 = ~new_R1222_U97;
  assign new_R1222_U307 = new_U4032 | new_U3055;
  assign new_R1222_U308 = ~new_R1222_U307 | ~new_R1222_U97;
  assign new_R1222_U309 = ~new_R1222_U145 | ~new_R1222_U308;
  assign new_R1222_U310 = ~new_R1222_U306 | ~new_R1222_U184;
  assign new_R1222_U311 = ~new_U3054 | ~new_U4031;
  assign new_R1222_U312 = ~new_R1222_U146 | ~new_R1222_U310;
  assign new_R1222_U313 = new_U3055 | new_U4032;
  assign new_R1222_U314 = ~new_R1222_U278 | ~new_R1222_U174;
  assign new_R1222_U315 = ~new_R1222_U100;
  assign new_R1222_U316 = ~new_R1222_U10 | ~new_R1222_U100;
  assign new_R1222_U317 = ~new_R1222_U147 | ~new_R1222_U316;
  assign new_R1222_U318 = ~new_R1222_U316 | ~new_R1222_U274;
  assign new_R1222_U319 = ~new_R1222_U468 | ~new_R1222_U318;
  assign new_R1222_U320 = new_U3504 | new_U3078;
  assign new_R1222_U321 = ~new_R1222_U320 | ~new_R1222_U100;
  assign new_R1222_U322 = ~new_R1222_U148 | ~new_R1222_U321;
  assign new_R1222_U323 = ~new_R1222_U315 | ~new_R1222_U55;
  assign new_R1222_U324 = ~new_U3073 | ~new_U4037;
  assign new_R1222_U325 = ~new_R1222_U149 | ~new_R1222_U323;
  assign new_R1222_U326 = new_U3468 | new_U3075;
  assign new_R1222_U327 = ~new_R1222_U173;
  assign new_R1222_U328 = new_U3078 | new_U3504;
  assign new_R1222_U329 = new_U3498 | new_U3070;
  assign new_R1222_U330 = ~new_U3500 | ~new_U3066;
  assign new_R1222_U331 = ~new_R1222_U151 | ~new_R1222_U379;
  assign new_R1222_U332 = new_U3070 | new_U3498;
  assign new_R1222_U333 = ~new_R1222_U250 | ~new_R1222_U179;
  assign new_R1222_U334 = ~new_R1222_U102;
  assign new_R1222_U335 = new_U3490 | new_U3069;
  assign new_R1222_U336 = ~new_R1222_U335 | ~new_R1222_U102;
  assign new_R1222_U337 = ~new_R1222_U152 | ~new_R1222_U336;
  assign new_R1222_U338 = ~new_R1222_U334 | ~new_R1222_U183;
  assign new_R1222_U339 = ~new_U3077 | ~new_U3492;
  assign new_R1222_U340 = ~new_R1222_U153 | ~new_R1222_U338;
  assign new_R1222_U341 = new_U3069 | new_U3490;
  assign new_R1222_U342 = new_U3484 | new_U3080;
  assign new_R1222_U343 = ~new_R1222_U342 | ~new_R1222_U49;
  assign new_R1222_U344 = ~new_R1222_U154 | ~new_R1222_U343;
  assign new_R1222_U345 = ~new_R1222_U211 | ~new_R1222_U182;
  assign new_R1222_U346 = ~new_U3059 | ~new_U3486;
  assign new_R1222_U347 = ~new_R1222_U155 | ~new_R1222_U345;
  assign new_R1222_U348 = ~new_R1222_U212 | ~new_R1222_U182;
  assign new_R1222_U349 = ~new_R1222_U209 | ~new_R1222_U69;
  assign new_R1222_U350 = ~new_R1222_U216 | ~new_R1222_U29;
  assign new_R1222_U351 = ~new_R1222_U230 | ~new_R1222_U38;
  assign new_R1222_U352 = ~new_R1222_U233 | ~new_R1222_U191;
  assign new_R1222_U353 = ~new_R1222_U313 | ~new_R1222_U184;
  assign new_R1222_U354 = ~new_R1222_U294 | ~new_R1222_U90;
  assign new_R1222_U355 = ~new_R1222_U328 | ~new_R1222_U55;
  assign new_R1222_U356 = ~new_R1222_U278 | ~new_R1222_U59;
  assign new_R1222_U357 = ~new_R1222_U332 | ~new_R1222_U65;
  assign new_R1222_U358 = ~new_R1222_U341 | ~new_R1222_U183;
  assign new_R1222_U359 = ~new_R1222_U250 | ~new_R1222_U76;
  assign new_R1222_U360 = ~new_U4029 | ~new_U3051;
  assign new_R1222_U361 = ~new_R1222_U5 | ~new_R1222_U196 | ~new_R1222_U4;
  assign new_R1222_U362 = ~new_R1222_U195 | ~new_R1222_U5 | ~new_R1222_U4;
  assign new_R1222_U363 = ~new_R1222_U44;
  assign new_R1222_U364 = ~new_R1222_U98;
  assign new_R1222_U365 = ~new_R1222_U13 | ~new_R1222_U44;
  assign new_R1222_U366 = ~new_R1222_U16 | ~new_R1222_U179;
  assign new_R1222_U367 = ~new_R1222_U256 | ~new_R1222_U253;
  assign new_R1222_U368 = ~new_R1222_U81;
  assign new_R1222_U369 = ~new_R1222_U139 | ~new_R1222_U179;
  assign new_R1222_U370 = ~new_R1222_U368 | ~new_R1222_U258;
  assign new_R1222_U371 = ~new_R1222_U15 | ~new_R1222_U98;
  assign new_R1222_U372 = ~new_R1222_U202 | ~new_R1222_U29;
  assign new_R1222_U373 = ~new_R1222_U6 | ~new_R1222_U50;
  assign new_R1222_U374 = ~new_R1222_U156;
  assign new_R1222_U375 = ~new_R1222_U213 | ~new_R1222_U50;
  assign new_R1222_U376 = ~new_R1222_U130 | ~new_R1222_U375;
  assign new_R1222_U377 = ~new_R1222_U137 | ~new_R1222_U50;
  assign new_R1222_U378 = ~new_R1222_U179;
  assign new_R1222_U379 = ~new_R1222_U260 | ~new_R1222_U65;
  assign new_R1222_U380 = ~new_R1222_U9 | ~new_R1222_U101;
  assign new_R1222_U381 = ~new_R1222_U174;
  assign new_R1222_U382 = ~new_R1222_U329 | ~new_R1222_U101;
  assign new_R1222_U383 = ~new_R1222_U150 | ~new_R1222_U382;
  assign new_R1222_U384 = ~new_R1222_U141 | ~new_R1222_U101;
  assign new_R1222_U385 = ~new_R1222_U170;
  assign new_R1222_U386 = ~new_U3080 | ~new_R1222_U48;
  assign new_R1222_U387 = ~new_U3484 | ~new_R1222_U47;
  assign new_R1222_U388 = ~new_R1222_U387 | ~new_R1222_U386;
  assign new_R1222_U389 = ~new_R1222_U348 | ~new_R1222_U49;
  assign new_R1222_U390 = ~new_R1222_U388 | ~new_R1222_U211;
  assign new_R1222_U391 = ~new_U3081 | ~new_R1222_U45;
  assign new_R1222_U392 = ~new_U3482 | ~new_R1222_U46;
  assign new_R1222_U393 = ~new_R1222_U392 | ~new_R1222_U391;
  assign new_R1222_U394 = ~new_R1222_U156 | ~new_R1222_U349;
  assign new_R1222_U395 = ~new_R1222_U374 | ~new_R1222_U393;
  assign new_R1222_U396 = ~new_U3067 | ~new_R1222_U30;
  assign new_R1222_U397 = ~new_U3480 | ~new_R1222_U28;
  assign new_R1222_U398 = ~new_U3068 | ~new_R1222_U26;
  assign new_R1222_U399 = ~new_U3478 | ~new_R1222_U27;
  assign new_R1222_U400 = ~new_R1222_U399 | ~new_R1222_U398;
  assign new_R1222_U401 = ~new_R1222_U350 | ~new_R1222_U50;
  assign new_R1222_U402 = ~new_R1222_U400 | ~new_R1222_U202;
  assign new_R1222_U403 = ~new_U3064 | ~new_R1222_U39;
  assign new_R1222_U404 = ~new_U3476 | ~new_R1222_U37;
  assign new_R1222_U405 = ~new_U3057 | ~new_R1222_U35;
  assign new_R1222_U406 = ~new_U3474 | ~new_R1222_U36;
  assign new_R1222_U407 = ~new_R1222_U406 | ~new_R1222_U405;
  assign new_R1222_U408 = ~new_R1222_U351 | ~new_R1222_U51;
  assign new_R1222_U409 = ~new_R1222_U407 | ~new_R1222_U223;
  assign new_R1222_U410 = ~new_U3061 | ~new_R1222_U33;
  assign new_R1222_U411 = ~new_U3472 | ~new_R1222_U34;
  assign new_R1222_U412 = ~new_R1222_U411 | ~new_R1222_U410;
  assign new_R1222_U413 = ~new_R1222_U352 | ~new_R1222_U157;
  assign new_R1222_U414 = ~new_R1222_U232 | ~new_R1222_U412;
  assign new_R1222_U415 = ~new_U3065 | ~new_R1222_U31;
  assign new_R1222_U416 = ~new_U3470 | ~new_R1222_U32;
  assign new_R1222_U417 = ~new_U3052 | ~new_R1222_U159;
  assign new_R1222_U418 = ~new_U4040 | ~new_R1222_U158;
  assign new_R1222_U419 = ~new_U3052 | ~new_R1222_U159;
  assign new_R1222_U420 = ~new_U4040 | ~new_R1222_U158;
  assign new_R1222_U421 = ~new_R1222_U420 | ~new_R1222_U419;
  assign new_R1222_U422 = ~new_R1222_U160 | ~new_R1222_U161;
  assign new_R1222_U423 = ~new_R1222_U304 | ~new_R1222_U421;
  assign new_R1222_U424 = ~new_U3051 | ~new_R1222_U96;
  assign new_R1222_U425 = ~new_U4029 | ~new_R1222_U95;
  assign new_R1222_U426 = ~new_U3051 | ~new_R1222_U96;
  assign new_R1222_U427 = ~new_U4029 | ~new_R1222_U95;
  assign new_R1222_U428 = ~new_R1222_U427 | ~new_R1222_U426;
  assign new_R1222_U429 = ~new_R1222_U162 | ~new_R1222_U163;
  assign new_R1222_U430 = ~new_R1222_U302 | ~new_R1222_U428;
  assign new_R1222_U431 = ~new_U3050 | ~new_R1222_U93;
  assign new_R1222_U432 = ~new_U4030 | ~new_R1222_U94;
  assign new_R1222_U433 = ~new_U3050 | ~new_R1222_U93;
  assign new_R1222_U434 = ~new_U4030 | ~new_R1222_U94;
  assign new_R1222_U435 = ~new_R1222_U434 | ~new_R1222_U433;
  assign new_R1222_U436 = ~new_R1222_U164 | ~new_R1222_U165;
  assign new_R1222_U437 = ~new_R1222_U298 | ~new_R1222_U435;
  assign new_R1222_U438 = ~new_U3054 | ~new_R1222_U91;
  assign new_R1222_U439 = ~new_U4031 | ~new_R1222_U92;
  assign new_R1222_U440 = ~new_U3055 | ~new_R1222_U86;
  assign new_R1222_U441 = ~new_U4032 | ~new_R1222_U87;
  assign new_R1222_U442 = ~new_R1222_U441 | ~new_R1222_U440;
  assign new_R1222_U443 = ~new_R1222_U353 | ~new_R1222_U97;
  assign new_R1222_U444 = ~new_R1222_U442 | ~new_R1222_U306;
  assign new_R1222_U445 = ~new_U3062 | ~new_R1222_U88;
  assign new_R1222_U446 = ~new_U4033 | ~new_R1222_U89;
  assign new_R1222_U447 = ~new_R1222_U446 | ~new_R1222_U445;
  assign new_R1222_U448 = ~new_R1222_U354 | ~new_R1222_U166;
  assign new_R1222_U449 = ~new_R1222_U288 | ~new_R1222_U447;
  assign new_R1222_U450 = ~new_U3063 | ~new_R1222_U84;
  assign new_R1222_U451 = ~new_U4034 | ~new_R1222_U85;
  assign new_R1222_U452 = ~new_U3063 | ~new_R1222_U84;
  assign new_R1222_U453 = ~new_U4034 | ~new_R1222_U85;
  assign new_R1222_U454 = ~new_R1222_U453 | ~new_R1222_U452;
  assign new_R1222_U455 = ~new_R1222_U167 | ~new_R1222_U168;
  assign new_R1222_U456 = ~new_R1222_U284 | ~new_R1222_U454;
  assign new_R1222_U457 = ~new_U3058 | ~new_R1222_U82;
  assign new_R1222_U458 = ~new_U4035 | ~new_R1222_U83;
  assign new_R1222_U459 = ~new_U3058 | ~new_R1222_U82;
  assign new_R1222_U460 = ~new_U4035 | ~new_R1222_U83;
  assign new_R1222_U461 = ~new_R1222_U460 | ~new_R1222_U459;
  assign new_R1222_U462 = ~new_R1222_U169 | ~new_R1222_U170;
  assign new_R1222_U463 = ~new_R1222_U385 | ~new_R1222_U461;
  assign new_R1222_U464 = ~new_U3072 | ~new_R1222_U60;
  assign new_R1222_U465 = ~new_U4036 | ~new_R1222_U61;
  assign new_R1222_U466 = ~new_U3072 | ~new_R1222_U60;
  assign new_R1222_U467 = ~new_U4036 | ~new_R1222_U61;
  assign new_R1222_U468 = ~new_R1222_U467 | ~new_R1222_U466;
  assign new_R1222_U469 = ~new_U3073 | ~new_R1222_U56;
  assign new_R1222_U470 = ~new_U4037 | ~new_R1222_U99;
  assign new_R1222_U471 = ~new_R1222_U193 | ~new_R1222_U173;
  assign new_R1222_U472 = ~new_R1222_U327 | ~new_R1222_U172;
  assign new_R1222_U473 = ~new_U3078 | ~new_R1222_U53;
  assign new_R1222_U474 = ~new_U3504 | ~new_R1222_U54;
  assign new_R1222_U475 = ~new_R1222_U474 | ~new_R1222_U473;
  assign new_R1222_U476 = ~new_R1222_U355 | ~new_R1222_U100;
  assign new_R1222_U477 = ~new_R1222_U475 | ~new_R1222_U315;
  assign new_R1222_U478 = ~new_U3079 | ~new_R1222_U57;
  assign new_R1222_U479 = ~new_U3502 | ~new_R1222_U58;
  assign new_R1222_U480 = ~new_R1222_U479 | ~new_R1222_U478;
  assign new_R1222_U481 = ~new_R1222_U174 | ~new_R1222_U356;
  assign new_R1222_U482 = ~new_R1222_U381 | ~new_R1222_U480;
  assign new_R1222_U483 = ~new_U3066 | ~new_R1222_U66;
  assign new_R1222_U484 = ~new_U3500 | ~new_R1222_U64;
  assign new_R1222_U485 = ~new_U3070 | ~new_R1222_U62;
  assign new_R1222_U486 = ~new_U3498 | ~new_R1222_U63;
  assign new_R1222_U487 = ~new_R1222_U486 | ~new_R1222_U485;
  assign new_R1222_U488 = ~new_R1222_U357 | ~new_R1222_U101;
  assign new_R1222_U489 = ~new_R1222_U487 | ~new_R1222_U260;
  assign new_R1222_U490 = ~new_U3071 | ~new_R1222_U67;
  assign new_R1222_U491 = ~new_U3496 | ~new_R1222_U68;
  assign new_R1222_U492 = ~new_U3071 | ~new_R1222_U67;
  assign new_R1222_U493 = ~new_U3496 | ~new_R1222_U68;
  assign new_R1222_U494 = ~new_R1222_U493 | ~new_R1222_U492;
  assign new_not_keyinput0 = ~keyinput0;
  assign new_not_keyinput1 = ~keyinput1;
  assign new_not_keyinput2 = ~keyinput2;
  assign new_not_keyinput3 = ~keyinput3;
  assign new_not_keyinput4 = ~keyinput4;
  assign new_not_0 = ~Q_1;
  assign new_and_1 = new_not_0 & Q_3;
  assign new_not_2 = ~Q_2;
  assign new_and_3 = new_not_2 & Q_3;
  assign new_not_4 = ~Q_0;
  assign new_and_5 = new_not_4 & Q_3;
  assign new_not_6 = ~Q_3;
  assign new_and_7 = new_not_6 & Q_2 & Q_0 & Q_1;
  assign n20711 = new_and_7 | new_and_5 | new_and_1 | new_and_3;
  assign new_not_9 = ~Q_2;
  assign new_and_10 = new_not_9 & Q_0 & Q_1;
  assign new_not_11 = ~Q_0;
  assign new_and_12 = new_not_11 & Q_2;
  assign new_not_13 = ~Q_1;
  assign new_and_14 = new_not_13 & Q_2;
  assign n20708 = new_and_14 | new_and_10 | new_and_12;
  assign new_not_16 = ~Q_1;
  assign new_and_17 = Q_0 & new_not_16;
  assign new_not_18 = ~Q_0;
  assign new_and_19 = new_not_18 & Q_1;
  assign n20705 = new_and_17 | new_and_19;
  assign n20702 = ~Q_0;
  assign new_not_Q_0 = ~Q_0;
  assign new_not_Q_1 = ~Q_1;
  assign new_not_Q_2 = ~Q_2;
  assign new_not_Q_3 = ~Q_3;
  assign new_count_state_1 = Q_0 & new_not_Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_2 = new_not_Q_0 & Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_3 = Q_0 & Q_1 & new_not_Q_3 & new_not_Q_2;
  assign new_count_state_4 = new_not_Q_0 & new_not_Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_5 = Q_0 & new_not_Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_6 = new_not_Q_0 & Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_7 = Q_0 & Q_1 & new_not_Q_3 & Q_2;
  assign new_count_state_8 = new_not_Q_0 & new_not_Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_9 = Q_0 & new_not_Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_10 = new_not_Q_0 & Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_11 = Q_0 & Q_1 & Q_3 & new_not_Q_2;
  assign new_count_state_12 = new_not_Q_0 & new_not_Q_1 & Q_3 & Q_2;
  assign new_count_state_13 = Q_0 & new_not_Q_1 & Q_3 & Q_2;
  assign new_count_state_14 = new_not_Q_0 & Q_1 & Q_3 & Q_2;
  assign new_count_state_15 = Q_0 & Q_1 & Q_3 & Q_2;
  assign new_y_mux_key0_and_0 = n194 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_1 = new_U3352 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0 = new_y_mux_key0_and_0 | new_y_mux_key0_and_1;
  assign new_y_mux_key1_and_0 = n194 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key1_and_1 = new_U3352 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1 = new_y_mux_key1_and_0 | new_y_mux_key1_and_1;
  assign new_y_mux_key2_and_0 = n194 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key2_and_1 = new_U3352 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2 = new_y_mux_key2_and_0 | new_y_mux_key2_and_1;
  assign new_y_mux_key3_and_0 = n194 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3_and_1 = new_U3352 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3 = new_y_mux_key3_and_0 | new_y_mux_key3_and_1;
  assign new_y_mux_key4_and_0 = n194 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key4_and_1 = new_U3352 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key4 = new_y_mux_key4_and_0 | new_y_mux_key4_and_1;
  assign new_y_mux_key5_and_0 = n194 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key5_and_1 = new_U3352 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key5 = new_y_mux_key5_and_0 | new_y_mux_key5_and_1;
  assign new_y_mux_key6_and_0 = n194 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key6_and_1 = new_U3352 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key6 = new_y_mux_key6_and_0 | new_y_mux_key6_and_1;
  assign new_y_mux_key7_and_0 = n194 & keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key7_and_1 = new_U3352 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key7 = new_y_mux_key7_and_0 | new_y_mux_key7_and_1;
  assign new_y_mux_key8_and_0 = n194 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8_and_1 = new_U3352 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key8 = new_y_mux_key8_and_0 | new_y_mux_key8_and_1;
  assign new_y_mux_key9_and_0 = n194 & keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key9_and_1 = new_U3352 & keyinput4 & keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key9 = new_y_mux_key9_and_0 | new_y_mux_key9_and_1;
  assign new_y_mux_key10_and_0 = n194 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10_and_1 = new_U3352 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key10 = new_y_mux_key10_and_0 | new_y_mux_key10_and_1;
  assign new_y_mux_key11_and_0 = n194 & new_not_keyinput4 & keyinput3 & new_not_keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key11_and_1 = new_U3352 & keyinput4 & new_not_keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key11 = new_y_mux_key11_and_0 | new_y_mux_key11_and_1;
  assign new_y_mux_key12_and_0 = n194 & new_not_keyinput4 & new_not_keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key12_and_1 = new_U3352 & new_not_keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key12 = new_y_mux_key12_and_0 | new_y_mux_key12_and_1;
  assign new_y_mux_key13_and_0 = n194 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key13_and_1 = new_U3352 & keyinput4 & keyinput3 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key13 = new_y_mux_key13_and_0 | new_y_mux_key13_and_1;
  assign new_y_mux_key14_and_0 = n194 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & keyinput1;
  assign new_y_mux_key14_and_1 = new_U3352 & new_not_keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key14 = new_y_mux_key14_and_0 | new_y_mux_key14_and_1;
  assign new_y_mux_key15_and_0 = n194 & new_not_keyinput4 & keyinput3 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15_and_1 = new_U3352 & keyinput4 & new_not_keyinput3 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key15 = new_y_mux_key15_and_0 | new_y_mux_key15_and_1;
  assign new__state_1 = new_count_state_1;
  assign new__state_2 = new_count_state_2;
  assign new__state_3 = new_count_state_3;
  assign new__state_4 = new_count_state_4;
  assign new__state_5 = new_count_state_5;
  assign new__state_6 = new_count_state_6;
  assign new__state_7 = new_count_state_7;
  assign new__state_8 = new_count_state_8;
  assign new__state_9 = new_count_state_9;
  assign new__state_10 = new_count_state_10;
  assign new__state_11 = new_count_state_11;
  assign new__state_12 = new_count_state_12;
  assign new__state_13 = new_count_state_13;
  assign new__state_14 = new_count_state_14;
  assign new__state_15 = new_count_state_15;
  assign new__state_17 = new__state_2 | new__state_3;
  assign new__state_18 = new__state_4 | new__state_5;
  assign new__state_19 = new__state_6 | new__state_7;
  assign new__state_20 = new__state_8 | new__state_9;
  assign new__state_21 = new__state_10 | new__state_11;
  assign new__state_22 = new__state_12 | new__state_13;
  assign new__state_23 = new__state_14 | new__state_15;
  assign new__state_25 = new__state_18 | new__state_19;
  assign new__state_26 = new__state_20 | new__state_21;
  assign new__state_27 = new__state_22 | new__state_23;
  assign new__state_29 = new__state_26 | new__state_27;
  assign new_s__state_1 = new__state_1;
  assign new_not_s__state_1 = ~new_s__state_1;
  assign new_I0__state_1 = new_y_mux_key0;
  assign new_I1__state_1 = new_y_mux_key1;
  assign new_and_mux__state_1 = new_not_s__state_1 & new_I0__state_1;
  assign new_and_mux__state_1_2 = new_s__state_1 & new_I1__state_1;
  assign new_y_mux_16 = new_and_mux__state_1 | new_and_mux__state_1_2;
  assign new_s__state_3 = new__state_3;
  assign new_not_s__state_3 = ~new_s__state_3;
  assign new_I0__state_3 = new_y_mux_key2;
  assign new_I1__state_3 = new_y_mux_key3;
  assign new_and_mux__state_3 = new_not_s__state_3 & new_I0__state_3;
  assign new_and_mux__state_3_2 = new_s__state_3 & new_I1__state_3;
  assign new_y_mux_17 = new_and_mux__state_3 | new_and_mux__state_3_2;
  assign new_s__state_5 = new__state_5;
  assign new_not_s__state_5 = ~new_s__state_5;
  assign new_I0__state_5 = new_y_mux_key4;
  assign new_I1__state_5 = new_y_mux_key5;
  assign new_and_mux__state_5 = new_not_s__state_5 & new_I0__state_5;
  assign new_and_mux__state_5_2 = new_s__state_5 & new_I1__state_5;
  assign new_y_mux_18 = new_and_mux__state_5 | new_and_mux__state_5_2;
  assign new_s__state_7 = new__state_7;
  assign new_not_s__state_7 = ~new_s__state_7;
  assign new_I0__state_7 = new_y_mux_key6;
  assign new_I1__state_7 = new_y_mux_key7;
  assign new_and_mux__state_7 = new_not_s__state_7 & new_I0__state_7;
  assign new_and_mux__state_7_2 = new_s__state_7 & new_I1__state_7;
  assign new_y_mux_19 = new_and_mux__state_7 | new_and_mux__state_7_2;
  assign new_s__state_9 = new__state_9;
  assign new_not_s__state_9 = ~new_s__state_9;
  assign new_I0__state_9 = new_y_mux_key8;
  assign new_I1__state_9 = new_y_mux_key9;
  assign new_and_mux__state_9 = new_not_s__state_9 & new_I0__state_9;
  assign new_and_mux__state_9_2 = new_s__state_9 & new_I1__state_9;
  assign new_y_mux_20 = new_and_mux__state_9 | new_and_mux__state_9_2;
  assign new_s__state_11 = new__state_11;
  assign new_not_s__state_11 = ~new_s__state_11;
  assign new_I0__state_11 = new_y_mux_key10;
  assign new_I1__state_11 = new_y_mux_key11;
  assign new_and_mux__state_11 = new_not_s__state_11 & new_I0__state_11;
  assign new_and_mux__state_11_2 = new_s__state_11 & new_I1__state_11;
  assign new_y_mux_21 = new_and_mux__state_11 | new_and_mux__state_11_2;
  assign new_s__state_13 = new__state_13;
  assign new_not_s__state_13 = ~new_s__state_13;
  assign new_I0__state_13 = new_y_mux_key12;
  assign new_I1__state_13 = new_y_mux_key13;
  assign new_and_mux__state_13 = new_not_s__state_13 & new_I0__state_13;
  assign new_and_mux__state_13_2 = new_s__state_13 & new_I1__state_13;
  assign new_y_mux_22 = new_and_mux__state_13 | new_and_mux__state_13_2;
  assign new_s__state_15 = new__state_15;
  assign new_not_s__state_15 = ~new_s__state_15;
  assign new_I0__state_15 = new_y_mux_key14;
  assign new_I1__state_15 = new_y_mux_key15;
  assign new_and_mux__state_15 = new_not_s__state_15 & new_I0__state_15;
  assign new_and_mux__state_15_2 = new_s__state_15 & new_I1__state_15;
  assign new_y_mux_23 = new_and_mux__state_15 | new_and_mux__state_15_2;
  assign new_s__state_17 = new__state_17;
  assign new_not_s__state_17 = ~new_s__state_17;
  assign new_I0__state_17 = new_y_mux_16;
  assign new_I1__state_17 = new_y_mux_17;
  assign new_and_mux__state_17 = new_not_s__state_17 & new_I0__state_17;
  assign new_and_mux__state_17_2 = new_s__state_17 & new_I1__state_17;
  assign new_y_mux_24 = new_and_mux__state_17 | new_and_mux__state_17_2;
  assign new_s__state_19 = new__state_19;
  assign new_not_s__state_19 = ~new_s__state_19;
  assign new_I0__state_19 = new_y_mux_18;
  assign new_I1__state_19 = new_y_mux_19;
  assign new_and_mux__state_19 = new_not_s__state_19 & new_I0__state_19;
  assign new_and_mux__state_19_2 = new_s__state_19 & new_I1__state_19;
  assign new_y_mux_25 = new_and_mux__state_19 | new_and_mux__state_19_2;
  assign new_s__state_21 = new__state_21;
  assign new_not_s__state_21 = ~new_s__state_21;
  assign new_I0__state_21 = new_y_mux_20;
  assign new_I1__state_21 = new_y_mux_21;
  assign new_and_mux__state_21 = new_not_s__state_21 & new_I0__state_21;
  assign new_and_mux__state_21_2 = new_s__state_21 & new_I1__state_21;
  assign new_y_mux_26 = new_and_mux__state_21 | new_and_mux__state_21_2;
  assign new_s__state_23 = new__state_23;
  assign new_not_s__state_23 = ~new_s__state_23;
  assign new_I0__state_23 = new_y_mux_22;
  assign new_I1__state_23 = new_y_mux_23;
  assign new_and_mux__state_23 = new_not_s__state_23 & new_I0__state_23;
  assign new_and_mux__state_23_2 = new_s__state_23 & new_I1__state_23;
  assign new_y_mux_27 = new_and_mux__state_23 | new_and_mux__state_23_2;
  assign new_s__state_25 = new__state_25;
  assign new_not_s__state_25 = ~new_s__state_25;
  assign new_I0__state_25 = new_y_mux_24;
  assign new_I1__state_25 = new_y_mux_25;
  assign new_and_mux__state_25 = new_not_s__state_25 & new_I0__state_25;
  assign new_and_mux__state_25_2 = new_s__state_25 & new_I1__state_25;
  assign new_y_mux_28 = new_and_mux__state_25 | new_and_mux__state_25_2;
  assign new_s__state_27 = new__state_27;
  assign new_not_s__state_27 = ~new_s__state_27;
  assign new_I0__state_27 = new_y_mux_26;
  assign new_I1__state_27 = new_y_mux_27;
  assign new_and_mux__state_27 = new_not_s__state_27 & new_I0__state_27;
  assign new_and_mux__state_27_2 = new_s__state_27 & new_I1__state_27;
  assign new_y_mux_29 = new_and_mux__state_27 | new_and_mux__state_27_2;
  assign new_s__state_29 = new__state_29;
  assign new_not_s__state_29 = ~new_s__state_29;
  assign new_I0__state_29 = new_y_mux_28;
  assign new_I1__state_29 = new_y_mux_29;
  assign new_and_mux__state_29 = new_not_s__state_29 & new_I0__state_29;
  assign new_and_mux__state_29_2 = new_s__state_29 & new_I1__state_29;
  assign n184 = new_and_mux__state_29 | new_and_mux__state_29_2;
  always @ (posedge clock) begin
    IR_REG_0_ <= n184;
    IR_REG_1_ <= n189;
    IR_REG_2_ <= n194;
    IR_REG_3_ <= n199;
    IR_REG_4_ <= n204;
    IR_REG_5_ <= n209;
    IR_REG_6_ <= n214;
    IR_REG_7_ <= n219;
    IR_REG_8_ <= n224;
    IR_REG_9_ <= n229;
    IR_REG_10_ <= n234;
    IR_REG_11_ <= n239;
    IR_REG_12_ <= n244;
    IR_REG_13_ <= n249;
    IR_REG_14_ <= n254;
    IR_REG_15_ <= n259;
    IR_REG_16_ <= n264;
    IR_REG_17_ <= n269;
    IR_REG_18_ <= n274;
    IR_REG_19_ <= n279;
    IR_REG_20_ <= n284;
    IR_REG_21_ <= n289;
    IR_REG_22_ <= n294;
    IR_REG_23_ <= n299;
    IR_REG_24_ <= n304;
    IR_REG_25_ <= n309;
    IR_REG_26_ <= n314;
    IR_REG_27_ <= n319;
    IR_REG_28_ <= n324;
    IR_REG_29_ <= n329;
    IR_REG_30_ <= n334;
    IR_REG_31_ <= n339;
    D_REG_0_ <= n344;
    D_REG_1_ <= n349;
    D_REG_2_ <= n354;
    D_REG_3_ <= n359;
    D_REG_4_ <= n364;
    D_REG_5_ <= n369;
    D_REG_6_ <= n374;
    D_REG_7_ <= n379;
    D_REG_8_ <= n384;
    D_REG_9_ <= n389;
    D_REG_10_ <= n394;
    D_REG_11_ <= n399;
    D_REG_12_ <= n404;
    D_REG_13_ <= n409;
    D_REG_14_ <= n414;
    D_REG_15_ <= n419;
    D_REG_16_ <= n424;
    D_REG_17_ <= n429;
    D_REG_18_ <= n434;
    D_REG_19_ <= n439;
    D_REG_20_ <= n444;
    D_REG_21_ <= n449;
    D_REG_22_ <= n454;
    D_REG_23_ <= n459;
    D_REG_24_ <= n464;
    D_REG_25_ <= n469;
    D_REG_26_ <= n474;
    D_REG_27_ <= n479;
    D_REG_28_ <= n484;
    D_REG_29_ <= n489;
    D_REG_30_ <= n494;
    D_REG_31_ <= n499;
    REG0_REG_0_ <= n504;
    REG0_REG_1_ <= n509;
    REG0_REG_2_ <= n514;
    REG0_REG_3_ <= n519;
    REG0_REG_4_ <= n524;
    REG0_REG_5_ <= n529;
    REG0_REG_6_ <= n534;
    REG0_REG_7_ <= n539;
    REG0_REG_8_ <= n544;
    REG0_REG_9_ <= n549;
    REG0_REG_10_ <= n554;
    REG0_REG_11_ <= n559;
    REG0_REG_12_ <= n564;
    REG0_REG_13_ <= n569;
    REG0_REG_14_ <= n574;
    REG0_REG_15_ <= n579;
    REG0_REG_16_ <= n584;
    REG0_REG_17_ <= n589;
    REG0_REG_18_ <= n594;
    REG0_REG_19_ <= n599;
    REG0_REG_20_ <= n604;
    REG0_REG_21_ <= n609;
    REG0_REG_22_ <= n614;
    REG0_REG_23_ <= n619;
    REG0_REG_24_ <= n624;
    REG0_REG_25_ <= n629;
    REG0_REG_26_ <= n634;
    REG0_REG_27_ <= n639;
    REG0_REG_28_ <= n644;
    REG0_REG_29_ <= n649;
    REG0_REG_30_ <= n654;
    REG0_REG_31_ <= n659;
    REG1_REG_0_ <= n664;
    REG1_REG_1_ <= n669;
    REG1_REG_2_ <= n674;
    REG1_REG_3_ <= n679;
    REG1_REG_4_ <= n684;
    REG1_REG_5_ <= n689;
    REG1_REG_6_ <= n694;
    REG1_REG_7_ <= n699;
    REG1_REG_8_ <= n704;
    REG1_REG_9_ <= n709;
    REG1_REG_10_ <= n714;
    REG1_REG_11_ <= n719;
    REG1_REG_12_ <= n724;
    REG1_REG_13_ <= n729;
    REG1_REG_14_ <= n734;
    REG1_REG_15_ <= n739;
    REG1_REG_16_ <= n744;
    REG1_REG_17_ <= n749;
    REG1_REG_18_ <= n754;
    REG1_REG_19_ <= n759;
    REG1_REG_20_ <= n764;
    REG1_REG_21_ <= n769;
    REG1_REG_22_ <= n774;
    REG1_REG_23_ <= n779;
    REG1_REG_24_ <= n784;
    REG1_REG_25_ <= n789;
    REG1_REG_26_ <= n794;
    REG1_REG_27_ <= n799;
    REG1_REG_28_ <= n804;
    REG1_REG_29_ <= n809;
    REG1_REG_30_ <= n814;
    REG1_REG_31_ <= n819;
    REG2_REG_0_ <= n824;
    REG2_REG_1_ <= n829;
    REG2_REG_2_ <= n834;
    REG2_REG_3_ <= n839;
    REG2_REG_4_ <= n844;
    REG2_REG_5_ <= n849;
    REG2_REG_6_ <= n854;
    REG2_REG_7_ <= n859;
    REG2_REG_8_ <= n864;
    REG2_REG_9_ <= n869;
    REG2_REG_10_ <= n874;
    REG2_REG_11_ <= n879;
    REG2_REG_12_ <= n884;
    REG2_REG_13_ <= n889;
    REG2_REG_14_ <= n894;
    REG2_REG_15_ <= n899;
    REG2_REG_16_ <= n904;
    REG2_REG_17_ <= n909;
    REG2_REG_18_ <= n914;
    REG2_REG_19_ <= n919;
    REG2_REG_20_ <= n924;
    REG2_REG_21_ <= n929;
    REG2_REG_22_ <= n934;
    REG2_REG_23_ <= n939;
    REG2_REG_24_ <= n944;
    REG2_REG_25_ <= n949;
    REG2_REG_26_ <= n954;
    REG2_REG_27_ <= n959;
    REG2_REG_28_ <= n964;
    REG2_REG_29_ <= n969;
    REG2_REG_30_ <= n974;
    REG2_REG_31_ <= n979;
    ADDR_REG_19_ <= n984;
    ADDR_REG_18_ <= n988;
    ADDR_REG_17_ <= n992;
    ADDR_REG_16_ <= n996;
    ADDR_REG_15_ <= n1000;
    ADDR_REG_14_ <= n1004;
    ADDR_REG_13_ <= n1008;
    ADDR_REG_12_ <= n1012;
    ADDR_REG_11_ <= n1016;
    ADDR_REG_10_ <= n1020;
    ADDR_REG_9_ <= n1024;
    ADDR_REG_8_ <= n1028;
    ADDR_REG_7_ <= n1032;
    ADDR_REG_6_ <= n1036;
    ADDR_REG_5_ <= n1040;
    ADDR_REG_4_ <= n1044;
    ADDR_REG_3_ <= n1048;
    ADDR_REG_2_ <= n1052;
    ADDR_REG_1_ <= n1056;
    ADDR_REG_0_ <= n1060;
    DATAO_REG_0_ <= n1064;
    DATAO_REG_1_ <= n1068;
    DATAO_REG_2_ <= n1072;
    DATAO_REG_3_ <= n1076;
    DATAO_REG_4_ <= n1080;
    DATAO_REG_5_ <= n1084;
    DATAO_REG_6_ <= n1088;
    DATAO_REG_7_ <= n1092;
    DATAO_REG_8_ <= n1096;
    DATAO_REG_9_ <= n1100;
    DATAO_REG_10_ <= n1104;
    DATAO_REG_11_ <= n1108;
    DATAO_REG_12_ <= n1112;
    DATAO_REG_13_ <= n1116;
    DATAO_REG_14_ <= n1120;
    DATAO_REG_15_ <= n1124;
    DATAO_REG_16_ <= n1128;
    DATAO_REG_17_ <= n1132;
    DATAO_REG_18_ <= n1136;
    DATAO_REG_19_ <= n1140;
    DATAO_REG_20_ <= n1144;
    DATAO_REG_21_ <= n1148;
    DATAO_REG_22_ <= n1152;
    DATAO_REG_23_ <= n1156;
    DATAO_REG_24_ <= n1160;
    DATAO_REG_25_ <= n1164;
    DATAO_REG_26_ <= n1168;
    DATAO_REG_27_ <= n1172;
    DATAO_REG_28_ <= n1176;
    DATAO_REG_29_ <= n1180;
    DATAO_REG_30_ <= n1184;
    DATAO_REG_31_ <= n1188;
    B_REG <= n1192;
    REG3_REG_15_ <= n1197;
    REG3_REG_26_ <= n1202;
    REG3_REG_6_ <= n1207;
    REG3_REG_18_ <= n1212;
    REG3_REG_2_ <= n1217;
    REG3_REG_11_ <= n1222;
    REG3_REG_22_ <= n1227;
    REG3_REG_13_ <= n1232;
    REG3_REG_20_ <= n1237;
    REG3_REG_0_ <= n1242;
    REG3_REG_9_ <= n1247;
    REG3_REG_4_ <= n1252;
    REG3_REG_24_ <= n1257;
    REG3_REG_17_ <= n1262;
    REG3_REG_5_ <= n1267;
    REG3_REG_16_ <= n1272;
    REG3_REG_25_ <= n1277;
    REG3_REG_12_ <= n1282;
    REG3_REG_21_ <= n1287;
    REG3_REG_1_ <= n1292;
    REG3_REG_8_ <= n1297;
    REG3_REG_28_ <= n1302;
    REG3_REG_19_ <= n1307;
    REG3_REG_3_ <= n1312;
    REG3_REG_10_ <= n1317;
    REG3_REG_23_ <= n1322;
    REG3_REG_14_ <= n1327;
    REG3_REG_27_ <= n1332;
    REG3_REG_7_ <= n1337;
    STATE_REG <= n1342;
    RD_REG <= n1347;
    WR_REG <= n1351;
    Q_0 <= n20702;
    Q_1 <= n20705;
    Q_2 <= n20708;
    Q_3 <= n20711;
  end
endmodule
