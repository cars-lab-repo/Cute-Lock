library ieee;
use ieee.std_logic_1164.all;

entity knot2 is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9 : out std_logic );
end knot2;

architecture ARC of knot2 is

   type states_knot2 is ( s1,s2,s3,s4,s5,s6,s7,s8,s9 );
   signal current_knot2 : states_knot2;

begin
   process (clk , rst)
   procedure proc_knot2 is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;

   case current_knot2 is
   when s1 =>
      if ( x1 and x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( x1 and not x2 and x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_knot2 <= s3;

      elsif ( x1 and not x2 and x3 and not x6 and x7 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         current_knot2 <= s3;

      elsif ( x1 and not x2 and x3 and not x6 and not x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_knot2 <= s3;

      elsif ( x1 and not x2 and not x3 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         current_knot2 <= s4;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         current_knot2 <= s5;

      end if;

   when s2 =>
      if ( x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_knot2 <= s6;

      elsif ( x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_knot2 <= s2;

      else
         y3 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s7;

      end if;

   when s3 =>
      if ( x6 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( x6 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_knot2 <= s6;

      elsif ( x6 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_knot2 <= s2;

      elsif ( x6 and not x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_knot2 <= s8;

      else
         y6 <= '1' ;
         current_knot2 <= s2;

      end if;

   when s4 =>
      if ( x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_knot2 <= s6;

      elsif ( x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_knot2 <= s2;

      else
         y6 <= '1' ;
         current_knot2 <= s2;

      end if;

   when s5 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         current_knot2 <= s9;

      elsif ( not x3 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( not x3 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_knot2 <= s6;

      elsif ( not x3 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_knot2 <= s2;

      else
         y6 <= '1' ;
         current_knot2 <= s2;

      end if;

   when s6 =>
      if ( x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s7;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         current_knot2 <= s1;

      end if;

   when s7 =>
      if ( x2 ) = '1' then
         y5 <= '1' ;
         current_knot2 <= s9;

      elsif ( not x2 and x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_knot2 <= s1;

      else
         y2 <= '1' ;
         y5 <= '1' ;
         current_knot2 <= s1;

      end if;

   when s8 =>
      if ( x3 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y4 <= '1' ;
         current_knot2 <= s3;

      elsif ( x3 and not x6 ) = '1' then
         y6 <= '1' ;
         current_knot2 <= s2;

      elsif ( not x3 and x4 and x5 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( not x3 and x4 and x5 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_knot2 <= s6;

      elsif ( not x3 and x4 and not x5 ) = '1' then
         y6 <= '1' ;
         current_knot2 <= s2;

      else
         y6 <= '1' ;
         current_knot2 <= s2;

      end if;

   when s9 =>
      if ( x6 and x3 ) = '1' then
         y4 <= '1' ;
         current_knot2 <= s9;

      elsif ( x6 and not x3 and x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_knot2 <= s2;

      elsif ( x6 and not x3 and not x1 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_knot2 <= s6;

      else
         y1 <= '1' ;
         y3 <= '1' ;
         current_knot2 <= s3;

      end if;

   end case;
   end proc_knot2;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;
	current_knot2 <= s1;
      elsif (clk'event and clk ='1') then
        proc_knot2;
      end if;
   end process;
end ARC;
